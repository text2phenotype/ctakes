C0010419|T201|COMP|20997-3|LNC|Cryptosporidium|Cryptosporidium
C0344390|T201|COMP|4690-4|LNC|Viscosity|Viscosity
C0362090|T201|COMP|1-8|LNC|Acyclovir|Acyclovir
C0362092|T201|COMP|3-4|LNC|Almecillin|Almecillin
C0362093|T201|COMP|4-2|LNC|Almecillin|Almecillin
C0362094|T201|COMP|5-9|LNC|Almecillin|Almecillin
C0362095|T201|COMP|6-7|LNC|Amantadine|Amantadine
C0362097|T201|COMP|8-3|LNC|Amdinocillin|Amdinocillin
C0362098|T201|COMP|9-1|LNC|Amdinocillin|Amdinocillin
C0362099|T201|COMP|10-9|LNC|Amdinocillin|Amdinocillin
C0362101|T201|COMP|12-5|LNC|Amikacin|Amikacin
C0362102|T201|COMP|13-3|LNC|Amikacin|Amikacin
C0362103|T201|COMP|14-1|LNC|Amikacin|Amikacin
C0362105|T201|COMP|16-6|LNC|Amoxicillin|Amoxicillin
C0362106|T201|COMP|17-4|LNC|Amoxicillin|Amoxicillin
C0362107|T201|COMP|18-2|LNC|Amoxicillin|Amoxicillin
C0362109|T201|COMP|20-8|LNC|Amoxicillin+Clavulanate|Amoxicillin+Clavulanate
C0362110|T201|COMP|21-6|LNC|Amoxicillin+Clavulanate|Amoxicillin+Clavulanate
C0362111|T201|COMP|22-4|LNC|Amoxicillin+Clavulanate|Amoxicillin+Clavulanate
C0362113|T201|COMP|24-0|LNC|Amphotericin B|Amphotericin B
C0362114|T201|COMP|25-7|LNC|Amphotericin B|Amphotericin B
C0362115|T201|COMP|26-5|LNC|Amphotericin B|Amphotericin B
C0362117|T201|COMP|28-1|LNC|Ampicillin|Ampicillin
C0362118|T201|COMP|29-9|LNC|Ampicillin|Ampicillin
C0362119|T201|COMP|30-7|LNC|Ampicillin|Ampicillin
C0362121|T201|COMP|32-3|LNC|Ampicillin+Sulbactam|Ampicillin+Sulbactam
C0362122|T201|COMP|33-1|LNC|Ampicillin+Sulbactam|Ampicillin+Sulbactam
C0362123|T201|COMP|34-9|LNC|Ampicillin+Sulbactam|Ampicillin+Sulbactam
C0362125|T201|COMP|36-4|LNC|Azithromycin|Azithromycin
C0362126|T201|COMP|37-2|LNC|Azithromycin|Azithromycin
C0362127|T201|COMP|38-0|LNC|Azithromycin|Azithromycin
C0362129|T201|COMP|40-6|LNC|Azlocillin|Azlocillin
C0362130|T201|COMP|41-4|LNC|Azlocillin|Azlocillin
C0362131|T201|COMP|42-2|LNC|Azlocillin|Azlocillin
C0362133|T201|COMP|44-8|LNC|Aztreonam|Aztreonam
C0362134|T201|COMP|45-5|LNC|Aztreonam|Aztreonam
C0362135|T201|COMP|46-3|LNC|Aztreonam|Aztreonam
C0362137|T201|COMP|48-9|LNC|Bacampicillin|Bacampicillin
C0362138|T201|COMP|49-7|LNC|Bacampicillin|Bacampicillin
C0362139|T201|COMP|50-5|LNC|Bacampicillin|Bacampicillin
C0362141|T201|COMP|52-1|LNC|Butirosin|Butirosin
C0362142|T201|COMP|53-9|LNC|Butirosin|Butirosin
C0362143|T201|COMP|54-7|LNC|Butirosin|Butirosin
C0362145|T201|COMP|56-2|LNC|Capreomycin|Capreomycin
C0362146|T201|COMP|57-0|LNC|Capreomycin|Capreomycin
C0362147|T201|COMP|58-8|LNC|Capreomycin|Capreomycin
C0362149|T201|COMP|60-4|LNC|Carbenicillin|Carbenicillin
C0362150|T201|COMP|61-2|LNC|Carbenicillin|Carbenicillin
C0362151|T201|COMP|62-0|LNC|Carbenicillin|Carbenicillin
C0362153|T201|COMP|64-6|LNC|Cefadroxil|Cefadroxil
C0362154|T201|COMP|65-3|LNC|Cefadroxil|Cefadroxil
C0362157|T201|COMP|68-7|LNC|Cefamandole|Cefamandole
C0362158|T201|COMP|69-5|LNC|Cefamandole|Cefamandole
C0362159|T201|COMP|70-3|LNC|Cefamandole|Cefamandole
C0362161|T201|COMP|72-9|LNC|Cefatrizine|Cefatrizine
C0362162|T201|COMP|73-7|LNC|Cefatrizine|Cefatrizine
C0362163|T201|COMP|74-5|LNC|Cefatrizine|Cefatrizine
C0362165|T201|COMP|76-0|LNC|ceFAZolin|ceFAZolin
C0362166|T201|COMP|77-8|LNC|ceFAZolin|ceFAZolin
C0362167|T201|COMP|78-6|LNC|ceFAZolin|ceFAZolin
C0362169|T201|COMP|80-2|LNC|Cefixime|Cefixime
C0362170|T201|COMP|81-0|LNC|Cefixime|Cefixime
C0362171|T201|COMP|82-8|LNC|Cefixime|Cefixime
C0362177|T201|COMP|88-5|LNC|Cefmetazole|Cefmetazole
C0362178|T201|COMP|89-3|LNC|Cefmetazole|Cefmetazole
C0362179|T201|COMP|90-1|LNC|Cefmetazole|Cefmetazole
C0362181|T201|COMP|92-7|LNC|Cefodizime|Cefodizime
C0362182|T201|COMP|93-5|LNC|Cefodizime|Cefodizime
C0362183|T201|COMP|94-3|LNC|Cefodizime|Cefodizime
C0362185|T201|COMP|96-8|LNC|Cefonicid|Cefonicid
C0362186|T201|COMP|97-6|LNC|Cefonicid|Cefonicid
C0362187|T201|COMP|98-4|LNC|Cefonicid|Cefonicid
C0362189|T201|COMP|100-8|LNC|Cefoperazone|Cefoperazone
C0362190|T201|COMP|101-6|LNC|Cefoperazone|Cefoperazone
C0362191|T201|COMP|102-4|LNC|Cefoperazone|Cefoperazone
C0362193|T201|COMP|104-0|LNC|Ceforanide|Ceforanide
C0362194|T201|COMP|105-7|LNC|Ceforanide|Ceforanide
C0362195|T201|COMP|106-5|LNC|Ceforanide|Ceforanide
C0362197|T201|COMP|108-1|LNC|Cefotaxime|Cefotaxime
C0362198|T201|COMP|109-9|LNC|Cefotaxime|Cefotaxime
C0362199|T201|COMP|110-7|LNC|Cefotaxime|Cefotaxime
C0362201|T201|COMP|112-3|LNC|cefoTEtan|cefoTEtan
C0362202|T201|COMP|113-1|LNC|cefoTEtan|cefoTEtan
C0362203|T201|COMP|114-9|LNC|cefoTEtan|cefoTEtan
C0362205|T201|COMP|116-4|LNC|cefOXitin|cefOXitin
C0362206|T201|COMP|117-2|LNC|cefOXitin|cefOXitin
C0362207|T201|COMP|118-0|LNC|cefOXitin|cefOXitin
C0362209|T201|COMP|120-6|LNC|Cefpodoxime|Cefpodoxime
C0362210|T201|COMP|121-4|LNC|Cefpodoxime|Cefpodoxime
C0362211|T201|COMP|122-2|LNC|Cefpodoxime|Cefpodoxime
C0362213|T201|COMP|124-8|LNC|Cefprozil|Cefprozil
C0362214|T201|COMP|125-5|LNC|Cefprozil|Cefprozil
C0362215|T201|COMP|126-3|LNC|Cefprozil|Cefprozil
C0362217|T201|COMP|128-9|LNC|Cefsulodin|Cefsulodin
C0362218|T201|COMP|129-7|LNC|Cefsulodin|Cefsulodin
C0362219|T201|COMP|130-5|LNC|Cefsulodin|Cefsulodin
C0362220|T201|COMP|131-3|LNC|Cefsulodin|Cefsulodin
C0362222|T201|COMP|133-9|LNC|cefTAZidime|cefTAZidime
C0362223|T201|COMP|134-7|LNC|cefTAZidime|cefTAZidime
C0362224|T201|COMP|135-4|LNC|cefTAZidime|cefTAZidime
C0362226|T201|COMP|137-0|LNC|Ceftizoxime|Ceftizoxime
C0362227|T201|COMP|138-8|LNC|Ceftizoxime|Ceftizoxime
C0362228|T201|COMP|139-6|LNC|Ceftizoxime|Ceftizoxime
C0362230|T201|COMP|141-2|LNC|cefTRIAXone|cefTRIAXone
C0362231|T201|COMP|142-0|LNC|cefTRIAXone|cefTRIAXone
C0362232|T201|COMP|143-8|LNC|cefTRIAXone|cefTRIAXone
C0362234|T201|COMP|145-3|LNC|Cefuroxime.parenteral|Cefuroxime.parenteral
C0362235|T201|COMP|146-1|LNC|Cefuroxime.parenteral|Cefuroxime.parenteral
C0362236|T201|COMP|147-9|LNC|Cefuroxime.parenteral|Cefuroxime.parenteral
C0362238|T201|COMP|149-5|LNC|Cephalexin|Cephalexin
C0362239|T201|COMP|150-3|LNC|Cephalexin|Cephalexin
C0362240|T201|COMP|151-1|LNC|Cephalexin|Cephalexin
C0362242|T201|COMP|153-7|LNC|Cephaloglycin|Cephaloglycin
C0362243|T201|COMP|154-5|LNC|Cephaloglycin|Cephaloglycin
C0362244|T201|COMP|155-2|LNC|Cephaloglycin|Cephaloglycin
C0362246|T201|COMP|157-8|LNC|Cephaloridine|Cephaloridine
C0362247|T201|COMP|158-6|LNC|Cephaloridine|Cephaloridine
C0362248|T201|COMP|159-4|LNC|Cephaloridine|Cephaloridine
C0362250|T201|COMP|161-0|LNC|Cephalothin|Cephalothin
C0362251|T201|COMP|162-8|LNC|Cephalothin|Cephalothin
C0362252|T201|COMP|163-6|LNC|Cephalothin|Cephalothin
C0362254|T201|COMP|165-1|LNC|Cephapirin|Cephapirin
C0362255|T201|COMP|166-9|LNC|Cephapirin|Cephapirin
C0362256|T201|COMP|167-7|LNC|Cephapirin|Cephapirin
C0362258|T201|COMP|169-3|LNC|Cephradine|Cephradine
C0362259|T201|COMP|170-1|LNC|Cephradine|Cephradine
C0362260|T201|COMP|171-9|LNC|Cephradine|Cephradine
C0362262|T201|COMP|173-5|LNC|Chloramphenicol|Chloramphenicol
C0362263|T201|COMP|174-3|LNC|Chloramphenicol|Chloramphenicol
C0362264|T201|COMP|175-0|LNC|Chloramphenicol|Chloramphenicol
C0362266|T201|COMP|177-6|LNC|Chlortetracycline|Chlortetracycline
C0362267|T201|COMP|178-4|LNC|Chlortetracycline|Chlortetracycline
C0362268|T201|COMP|179-2|LNC|Chlortetracycline|Chlortetracycline
C0362270|T201|COMP|181-8|LNC|Cinoxacin|Cinoxacin
C0362271|T201|COMP|182-6|LNC|Cinoxacin|Cinoxacin
C0362272|T201|COMP|183-4|LNC|Cinoxacin|Cinoxacin
C0362274|T201|COMP|185-9|LNC|Ciprofloxacin|Ciprofloxacin
C0362275|T201|COMP|186-7|LNC|Ciprofloxacin|Ciprofloxacin
C0362276|T201|COMP|187-5|LNC|Ciprofloxacin|Ciprofloxacin
C0362278|T201|COMP|189-1|LNC|Clarithromycin|Clarithromycin
C0362279|T201|COMP|190-9|LNC|Clarithromycin|Clarithromycin
C0362280|T201|COMP|191-7|LNC|Clarithromycin|Clarithromycin
C0362282|T201|COMP|193-3|LNC|Clindamycin|Clindamycin
C0362283|T201|COMP|194-1|LNC|Clindamycin|Clindamycin
C0362284|T201|COMP|195-8|LNC|Clindamycin|Clindamycin
C0362286|T201|COMP|197-4|LNC|Cloxacillin|Cloxacillin
C0362287|T201|COMP|198-2|LNC|Cloxacillin|Cloxacillin
C0362288|T201|COMP|199-0|LNC|Cloxacillin|Cloxacillin
C0362290|T201|COMP|201-4|LNC|Colistimethate|Colistimethate
C0362291|T201|COMP|202-2|LNC|Colistimethate|Colistimethate
C0362292|T201|COMP|203-0|LNC|Colistimethate|Colistimethate
C0362294|T201|COMP|205-5|LNC|Colistin|Colistin
C0362295|T201|COMP|206-3|LNC|Colistin|Colistin
C0362296|T201|COMP|207-1|LNC|Colistin|Colistin
C0362298|T201|COMP|209-7|LNC|Cyclacillin|Cyclacillin
C0362299|T201|COMP|210-5|LNC|Cyclacillin|Cyclacillin
C0362300|T201|COMP|211-3|LNC|Cyclacillin|Cyclacillin
C0362302|T201|COMP|213-9|LNC|cycloSERINE|cycloSERINE
C0362303|T201|COMP|214-7|LNC|cycloSERINE|cycloSERINE
C0362304|T201|COMP|215-4|LNC|cycloSERINE|cycloSERINE
C0362306|T201|COMP|217-0|LNC|Demeclocycline|Demeclocycline
C0362307|T201|COMP|218-8|LNC|Demeclocycline|Demeclocycline
C0362308|T201|COMP|219-6|LNC|Demeclocycline|Demeclocycline
C0362310|T201|COMP|221-2|LNC|Dicloxacillin|Dicloxacillin
C0362311|T201|COMP|222-0|LNC|Dicloxacillin|Dicloxacillin
C0362312|T201|COMP|223-8|LNC|Dicloxacillin|Dicloxacillin
C0362314|T201|COMP|225-3|LNC|Doxycycline|Doxycycline
C0362315|T201|COMP|226-1|LNC|Doxycycline|Doxycycline
C0362316|T201|COMP|227-9|LNC|Doxycycline|Doxycycline
C0362318|T201|COMP|229-5|LNC|Enoxacin|Enoxacin
C0362319|T201|COMP|230-3|LNC|Enoxacin|Enoxacin
C0362320|T201|COMP|231-1|LNC|Enoxacin|Enoxacin
C0362322|T201|COMP|233-7|LNC|Erythromycin|Erythromycin
C0362323|T201|COMP|234-5|LNC|Erythromycin|Erythromycin
C0362324|T201|COMP|235-2|LNC|Erythromycin|Erythromycin
C0362326|T201|COMP|237-8|LNC|Erythromycin+sulfiSOXAZOLE|Erythromycin+sulfiSOXAZOLE
C0362327|T201|COMP|238-6|LNC|Erythromycin+sulfiSOXAZOLE|Erythromycin+sulfiSOXAZOLE
C0362328|T201|COMP|239-4|LNC|Erythromycin+sulfiSOXAZOLE|Erythromycin+sulfiSOXAZOLE
C0362330|T201|COMP|241-0|LNC|Ethambutol|Ethambutol
C0362331|T201|COMP|242-8|LNC|Ethambutol|Ethambutol
C0362332|T201|COMP|243-6|LNC|Ethambutol|Ethambutol
C0362334|T201|COMP|245-1|LNC|Floxacillin|Floxacillin
C0362335|T201|COMP|246-9|LNC|Floxacillin|Floxacillin
C0362336|T201|COMP|247-7|LNC|Floxacillin|Floxacillin
C0362338|T201|COMP|249-3|LNC|Fluconazole|Fluconazole
C0362339|T201|COMP|250-1|LNC|Fluconazole|Fluconazole
C0362340|T201|COMP|251-9|LNC|Fluconazole|Fluconazole
C0362342|T201|COMP|253-5|LNC|5-Fluorocytosine|5-Fluorocytosine
C0362343|T201|COMP|254-3|LNC|5-Fluorocytosine|5-Fluorocytosine
C0362344|T201|COMP|255-0|LNC|5-Fluorocytosine|5-Fluorocytosine
C0362345|T201|COMP|256-8|LNC|Foscarnet|Foscarnet
C0362347|T201|COMP|258-4|LNC|Framycetin|Framycetin
C0362348|T201|COMP|259-2|LNC|Framycetin|Framycetin
C0362349|T201|COMP|260-0|LNC|Framycetin|Framycetin
C0362351|T201|COMP|262-6|LNC|Fusidate|Fusidate
C0362352|T201|COMP|263-4|LNC|Fusidate|Fusidate
C0362353|T201|COMP|264-2|LNC|Fusidate|Fusidate
C0362354|T201|COMP|265-9|LNC|Ganciclovir|Ganciclovir
C0362356|T201|COMP|267-5|LNC|Gentamicin|Gentamicin
C0362357|T201|COMP|268-3|LNC|Gentamicin|Gentamicin
C0362358|T201|COMP|269-1|LNC|Gentamicin|Gentamicin
C0362360|T201|COMP|271-7|LNC|Gramicidin D|Gramicidin D
C0362361|T201|COMP|272-5|LNC|Gramicidin D|Gramicidin D
C0362362|T201|COMP|273-3|LNC|Gramicidin D|Gramicidin D
C0362364|T201|COMP|275-8|LNC|Hetacillin|Hetacillin
C0362365|T201|COMP|276-6|LNC|Hetacillin|Hetacillin
C0362366|T201|COMP|277-4|LNC|Hetacillin|Hetacillin
C0362368|T201|COMP|279-0|LNC|Imipenem|Imipenem
C0362369|T201|COMP|280-8|LNC|Imipenem|Imipenem
C0362370|T201|COMP|281-6|LNC|Imipenem|Imipenem
C0362372|T201|COMP|283-2|LNC|Imipenem+Cilastatin|Imipenem+Cilastatin
C0362373|T201|COMP|284-0|LNC|Imipenem+Cilastatin|Imipenem+Cilastatin
C0362374|T201|COMP|285-7|LNC|Imipenem+Cilastatin|Imipenem+Cilastatin
C0362376|T201|COMP|287-3|LNC|Isoniazid|Isoniazid
C0362377|T201|COMP|288-1|LNC|Isoniazid|Isoniazid
C0362378|T201|COMP|289-9|LNC|Isoniazid|Isoniazid
C0362380|T201|COMP|291-5|LNC|Kanamycin|Kanamycin
C0362381|T201|COMP|292-3|LNC|Kanamycin|Kanamycin
C0362382|T201|COMP|293-1|LNC|Kanamycin|Kanamycin
C0362384|T201|COMP|295-6|LNC|Ketoconazole|Ketoconazole
C0362385|T201|COMP|296-4|LNC|Ketoconazole|Ketoconazole
C0362386|T201|COMP|297-2|LNC|Ketoconazole|Ketoconazole
C0362388|T201|COMP|299-8|LNC|Lincomycin|Lincomycin
C0362389|T201|COMP|300-4|LNC|Lincomycin|Lincomycin
C0362390|T201|COMP|301-2|LNC|Lincomycin|Lincomycin
C0362392|T201|COMP|303-8|LNC|Lomefloxacin|Lomefloxacin
C0362393|T201|COMP|304-6|LNC|Lomefloxacin|Lomefloxacin
C0362394|T201|COMP|305-3|LNC|Lomefloxacin|Lomefloxacin
C0362396|T201|COMP|307-9|LNC|Loracarbef|Loracarbef
C0362397|T201|COMP|308-7|LNC|Loracarbef|Loracarbef
C0362398|T201|COMP|309-5|LNC|Loracarbef|Loracarbef
C0362400|T201|COMP|311-1|LNC|Lymecycline|Lymecycline
C0362401|T201|COMP|312-9|LNC|Lymecycline|Lymecycline
C0362402|T201|COMP|313-7|LNC|Lymecycline|Lymecycline
C0362404|T201|COMP|315-2|LNC|Meclocycline|Meclocycline
C0362405|T201|COMP|316-0|LNC|Meclocycline|Meclocycline
C0362406|T201|COMP|317-8|LNC|Meclocycline|Meclocycline
C0362408|T201|COMP|319-4|LNC|Methacycline|Methacycline
C0362409|T201|COMP|320-2|LNC|Methacycline|Methacycline
C0362410|T201|COMP|321-0|LNC|Methacycline|Methacycline
C0362412|T201|COMP|323-6|LNC|Methicillin|Methicillin
C0362413|T201|COMP|324-4|LNC|Methicillin|Methicillin
C0362414|T201|COMP|325-1|LNC|Methicillin|Methicillin
C0362416|T201|COMP|327-7|LNC|metroNIDAZOLE|metroNIDAZOLE
C0362417|T201|COMP|328-5|LNC|metroNIDAZOLE|metroNIDAZOLE
C0362418|T201|COMP|329-3|LNC|metroNIDAZOLE|metroNIDAZOLE
C0362420|T201|COMP|331-9|LNC|Mezlocillin|Mezlocillin
C0362421|T201|COMP|332-7|LNC|Mezlocillin|Mezlocillin
C0362422|T201|COMP|333-5|LNC|Mezlocillin|Mezlocillin
C0362424|T201|COMP|335-0|LNC|Minocycline|Minocycline
C0362425|T201|COMP|336-8|LNC|Minocycline|Minocycline
C0362426|T201|COMP|337-6|LNC|Minocycline|Minocycline
C0362428|T201|COMP|339-2|LNC|Miocamycin|Miocamycin
C0362429|T201|COMP|340-0|LNC|Miocamycin|Miocamycin
C0362430|T201|COMP|341-8|LNC|Miocamycin|Miocamycin
C0362432|T201|COMP|343-4|LNC|Moxalactam|Moxalactam
C0362433|T201|COMP|344-2|LNC|Moxalactam|Moxalactam
C0362434|T201|COMP|345-9|LNC|Moxalactam|Moxalactam
C0362436|T201|COMP|347-5|LNC|Nafcillin|Nafcillin
C0362437|T201|COMP|348-3|LNC|Nafcillin|Nafcillin
C0362438|T201|COMP|349-1|LNC|Nafcillin|Nafcillin
C0362440|T201|COMP|351-7|LNC|Nalidixate|Nalidixate
C0362441|T201|COMP|352-5|LNC|Nalidixate|Nalidixate
C0362442|T201|COMP|353-3|LNC|Nalidixate|Nalidixate
C0362444|T201|COMP|355-8|LNC|Neomycin|Neomycin
C0362445|T201|COMP|356-6|LNC|Neomycin|Neomycin
C0362446|T201|COMP|357-4|LNC|Neomycin|Neomycin
C0362448|T201|COMP|359-0|LNC|Netilmicin|Netilmicin
C0362449|T201|COMP|360-8|LNC|Netilmicin|Netilmicin
C0362450|T201|COMP|361-6|LNC|Netilmicin|Netilmicin
C0362452|T201|COMP|363-2|LNC|Nitrofurantoin|Nitrofurantoin
C0362453|T201|COMP|364-0|LNC|Nitrofurantoin|Nitrofurantoin
C0362454|T201|COMP|365-7|LNC|Nitrofurantoin|Nitrofurantoin
C0362456|T201|COMP|367-3|LNC|Norfloxacin|Norfloxacin
C0362457|T201|COMP|368-1|LNC|Norfloxacin|Norfloxacin
C0362458|T201|COMP|369-9|LNC|Norfloxacin|Norfloxacin
C0362460|T201|COMP|371-5|LNC|Novobiocin|Novobiocin
C0362461|T201|COMP|372-3|LNC|Novobiocin|Novobiocin
C0362462|T201|COMP|373-1|LNC|Novobiocin|Novobiocin
C0362464|T201|COMP|375-6|LNC|Ofloxacin|Ofloxacin
C0362465|T201|COMP|376-4|LNC|Ofloxacin|Ofloxacin
C0362466|T201|COMP|377-2|LNC|Ofloxacin|Ofloxacin
C0362468|T201|COMP|379-8|LNC|Oleandomycin|Oleandomycin
C0362469|T201|COMP|380-6|LNC|Oleandomycin|Oleandomycin
C0362470|T201|COMP|381-4|LNC|Oleandomycin|Oleandomycin
C0362472|T201|COMP|383-0|LNC|Oxacillin|Oxacillin
C0362473|T201|COMP|384-8|LNC|Oxacillin|Oxacillin
C0362474|T201|COMP|385-5|LNC|Oxacillin|Oxacillin
C0362476|T201|COMP|387-1|LNC|Oxytetracycline|Oxytetracycline
C0362477|T201|COMP|388-9|LNC|Oxytetracycline|Oxytetracycline
C0362478|T201|COMP|389-7|LNC|Oxytetracycline|Oxytetracycline
C0362479|T201|COMP|390-5|LNC|Pefloxacin|Pefloxacin
C0362481|T201|COMP|392-1|LNC|Penicillin G|Penicillin G
C0362482|T201|COMP|393-9|LNC|Penicillin G|Penicillin G
C0362483|T201|COMP|394-7|LNC|Penicillin G|Penicillin G
C0362485|T201|COMP|396-2|LNC|Penicillin V|Penicillin V
C0362486|T201|COMP|397-0|LNC|Penicillin V|Penicillin V
C0362487|T201|COMP|398-8|LNC|Penicillin V|Penicillin V
C0362489|T201|COMP|400-2|LNC|Phenethicillin|Phenethicillin
C0362490|T201|COMP|401-0|LNC|Phenethicillin|Phenethicillin
C0362491|T201|COMP|402-8|LNC|Phenethicillin|Phenethicillin
C0362493|T201|COMP|404-4|LNC|Pipemidate|Pipemidate
C0362494|T201|COMP|405-1|LNC|Pipemidate|Pipemidate
C0362495|T201|COMP|406-9|LNC|Pipemidate|Pipemidate
C0362497|T201|COMP|408-5|LNC|Piperacillin|Piperacillin
C0362498|T201|COMP|409-3|LNC|Piperacillin|Piperacillin
C0362499|T201|COMP|410-1|LNC|Piperacillin|Piperacillin
C0362501|T201|COMP|412-7|LNC|Piperacillin+Tazobactam|Piperacillin+Tazobactam
C0362502|T201|COMP|413-5|LNC|Piperacillin+Tazobactam|Piperacillin+Tazobactam
C0362503|T201|COMP|414-3|LNC|Piperacillin+Tazobactam|Piperacillin+Tazobactam
C0362505|T201|COMP|416-8|LNC|Pivampicillin|Pivampicillin
C0362506|T201|COMP|417-6|LNC|Pivampicillin|Pivampicillin
C0362507|T201|COMP|418-4|LNC|Pivampicillin|Pivampicillin
C0362509|T201|COMP|420-0|LNC|Polymyxin B|Polymyxin B
C0362510|T201|COMP|421-8|LNC|Polymyxin B|Polymyxin B
C0362511|T201|COMP|422-6|LNC|Polymyxin B|Polymyxin B
C0362513|T201|COMP|424-2|LNC|Pyrazinamide|Pyrazinamide
C0362514|T201|COMP|425-9|LNC|Pyrazinamide|Pyrazinamide
C0362515|T201|COMP|426-7|LNC|Pyrazinamide|Pyrazinamide
C0362517|T201|COMP|428-3|LNC|rifAMPin|rifAMPin
C0362518|T201|COMP|429-1|LNC|rifAMPin|rifAMPin
C0362519|T201|COMP|430-9|LNC|rifAMPin|rifAMPin
C0362521|T201|COMP|432-5|LNC|Ristocetin|Ristocetin
C0362522|T201|COMP|433-3|LNC|Ristocetin|Ristocetin
C0362523|T201|COMP|434-1|LNC|Ristocetin|Ristocetin
C0362525|T201|COMP|436-6|LNC|Rolitetracycline|Rolitetracycline
C0362526|T201|COMP|437-4|LNC|Rolitetracycline|Rolitetracycline
C0362527|T201|COMP|438-2|LNC|Rolitetracycline|Rolitetracycline
C0362529|T201|COMP|440-8|LNC|Rosoxacin|Rosoxacin
C0362530|T201|COMP|441-6|LNC|Rosoxacin|Rosoxacin
C0362531|T201|COMP|442-4|LNC|Rosoxacin|Rosoxacin
C0362533|T201|COMP|444-0|LNC|Roxithromycin|Roxithromycin
C0362534|T201|COMP|445-7|LNC|Roxithromycin|Roxithromycin
C0362535|T201|COMP|446-5|LNC|Roxithromycin|Roxithromycin
C0362537|T201|COMP|448-1|LNC|Sisomicin|Sisomicin
C0362538|T201|COMP|449-9|LNC|Sisomicin|Sisomicin
C0362539|T201|COMP|450-7|LNC|Sisomicin|Sisomicin
C0362541|T201|COMP|452-3|LNC|Spectinomycin|Spectinomycin
C0362542|T201|COMP|453-1|LNC|Spectinomycin|Spectinomycin
C0362543|T201|COMP|454-9|LNC|Spectinomycin|Spectinomycin
C0362545|T201|COMP|456-4|LNC|Spiramycin|Spiramycin
C0362546|T201|COMP|457-2|LNC|Spiramycin|Spiramycin
C0362547|T201|COMP|458-0|LNC|Spiramycin|Spiramycin
C0362549|T201|COMP|460-6|LNC|Streptomycin|Streptomycin
C0362550|T201|COMP|461-4|LNC|Streptomycin|Streptomycin
C0362551|T201|COMP|462-2|LNC|Streptomycin|Streptomycin
C0362553|T201|COMP|464-8|LNC|sulfADIAZINE|sulfADIAZINE
C0362554|T201|COMP|465-5|LNC|sulfADIAZINE|sulfADIAZINE
C0362555|T201|COMP|466-3|LNC|sulfADIAZINE|sulfADIAZINE
C0362557|T201|COMP|468-9|LNC|Sulfamethoxazole|Sulfamethoxazole
C0362558|T201|COMP|469-7|LNC|Sulfamethoxazole|Sulfamethoxazole
C0362559|T201|COMP|470-5|LNC|Sulfamethoxazole|Sulfamethoxazole
C0362561|T201|COMP|472-1|LNC|sulfiSOXAZOLE|sulfiSOXAZOLE
C0362562|T201|COMP|473-9|LNC|sulfiSOXAZOLE|sulfiSOXAZOLE
C0362563|T201|COMP|474-7|LNC|sulfiSOXAZOLE|sulfiSOXAZOLE
C0362565|T201|COMP|476-2|LNC|Sulfonamide|Sulfonamide
C0362566|T201|COMP|477-0|LNC|Sulfonamide|Sulfonamide
C0362567|T201|COMP|478-8|LNC|Sulfonamide|Sulfonamide
C0362569|T201|COMP|480-4|LNC|Talampicillin|Talampicillin
C0362570|T201|COMP|481-2|LNC|Talampicillin|Talampicillin
C0362571|T201|COMP|482-0|LNC|Talampicillin|Talampicillin
C0362573|T201|COMP|484-6|LNC|Teicoplanin|Teicoplanin
C0362574|T201|COMP|485-3|LNC|Teicoplanin|Teicoplanin
C0362575|T201|COMP|486-1|LNC|Teicoplanin|Teicoplanin
C0362577|T201|COMP|488-7|LNC|Temafloxacin|Temafloxacin
C0362578|T201|COMP|489-5|LNC|Temafloxacin|Temafloxacin
C0362579|T201|COMP|490-3|LNC|Temafloxacin|Temafloxacin
C0362581|T201|COMP|492-9|LNC|Temocillin|Temocillin
C0362582|T201|COMP|493-7|LNC|Temocillin|Temocillin
C0362583|T201|COMP|494-5|LNC|Temocillin|Temocillin
C0362585|T201|COMP|496-0|LNC|Tetracycline|Tetracycline
C0362586|T201|COMP|497-8|LNC|Tetracycline|Tetracycline
C0362587|T201|COMP|498-6|LNC|Tetracycline|Tetracycline
C0362589|T201|COMP|500-9|LNC|Ticarcillin|Ticarcillin
C0362590|T201|COMP|501-7|LNC|Ticarcillin|Ticarcillin
C0362591|T201|COMP|502-5|LNC|Ticarcillin|Ticarcillin
C0362593|T201|COMP|504-1|LNC|Ticarcillin+Clavulanate|Ticarcillin+Clavulanate
C0362594|T201|COMP|505-8|LNC|Ticarcillin+Clavulanate|Ticarcillin+Clavulanate
C0362595|T201|COMP|506-6|LNC|Ticarcillin+Clavulanate|Ticarcillin+Clavulanate
C0362597|T201|COMP|508-2|LNC|Tobramycin|Tobramycin
C0362598|T201|COMP|509-0|LNC|Tobramycin|Tobramycin
C0362599|T201|COMP|510-8|LNC|Tobramycin|Tobramycin
C0362601|T201|COMP|512-4|LNC|Trimethoprim|Trimethoprim
C0362602|T201|COMP|513-2|LNC|Trimethoprim|Trimethoprim
C0362603|T201|COMP|514-0|LNC|Trimethoprim|Trimethoprim
C0362605|T201|COMP|516-5|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0362606|T201|COMP|517-3|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0362607|T201|COMP|518-1|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0362609|T201|COMP|520-7|LNC|Troleandomycin|Troleandomycin
C0362610|T201|COMP|521-5|LNC|Troleandomycin|Troleandomycin
C0362611|T201|COMP|522-3|LNC|Troleandomycin|Troleandomycin
C0362613|T201|COMP|524-9|LNC|Vancomycin|Vancomycin
C0362614|T201|COMP|525-6|LNC|Vancomycin|Vancomycin
C0362615|T201|COMP|526-4|LNC|Vancomycin|Vancomycin
C0362617|T201|COMP|528-0|LNC|Viomycin|Viomycin
C0362618|T201|COMP|529-8|LNC|Viomycin|Viomycin
C0362619|T201|COMP|530-6|LNC|Viomycin|Viomycin
C0362620|T201|COMP|531-4|LNC|Zidovudine|Zidovudine
C0362621|T201|COMP|6015-2|LNC|Acacia longifolia Ab.IgE|Acacia longifolia Ab.IgE
C0362623|T201|COMP|6017-8|LNC|Alder Ab.IgE|Alder Ab.IgE
C0362624|T201|COMP|6018-6|LNC|House dust Allergopharma Ab.IgE|House dust Allergopharma Ab.IgE
C0362625|T201|COMP|6019-4|LNC|Prunus dulcis Ab.IgE|Prunus dulcis Ab.IgE
C0362627|T201|COMP|6021-0|LNC|Malus sylvestris Ab.IgE|Malus sylvestris Ab.IgE
C0362628|T201|COMP|6022-8|LNC|Ascaris sp Ab.IgE|Ascaris sp Ab.IgE
C0362629|T201|COMP|6023-6|LNC|Aspergillus amstelodami Ab.IgE|Aspergillus amstelodami Ab.IgE
C0362630|T201|COMP|6024-4|LNC|Aspergillus flavus Ab.IgE|Aspergillus flavus Ab.IgE
C0362631|T201|COMP|6025-1|LNC|Aspergillus fumigatus Ab.IgE|Aspergillus fumigatus Ab.IgE
C0362632|T201|COMP|6026-9|LNC|Aspergillus terreus Ab.IgE|Aspergillus terreus Ab.IgE
C0362633|T201|COMP|6027-7|LNC|Aspergillus versicolor Ab.IgE|Aspergillus versicolor Ab.IgE
C0362634|T201|COMP|6029-3|LNC|Aureobasidium pullulans Ab.IgE|Aureobasidium pullulans Ab.IgE
C0362635|T201|COMP|6304-0|LNC|Budgerigar droppings Ab.IgE|Budgerigar droppings Ab.IgE
C0362636|T201|COMP|6030-1|LNC|Budgerigar feather Ab.IgE|Budgerigar feather Ab.IgE
C0362637|T201|COMP|6031-9|LNC|Budgerigar serum proteins Ab.IgE|Budgerigar serum proteins Ab.IgE
C0362638|T201|COMP|6032-7|LNC|Casuarina equisetifolia Ab.IgE|Casuarina equisetifolia Ab.IgE
C0362639|T201|COMP|6033-5|LNC|Persea americana Ab.IgE|Persea americana Ab.IgE
C0362640|T201|COMP|6034-3|LNC|Paspalum notatum Ab.IgE|Paspalum notatum Ab.IgE
C0362641|T201|COMP|6035-0|LNC|Musa spp Ab.IgE|Musa spp Ab.IgE
C0362642|T201|COMP|6037-6|LNC|Hordeum vulgare Ab.IgE|Hordeum vulgare Ab.IgE
C0362644|T201|COMP|6038-4|LNC|Fagus grandifolia Ab.IgE|Fagus grandifolia Ab.IgE
C0362645|T201|COMP|6039-2|LNC|Beef Ab.IgE|Beef Ab.IgE
C0362646|T201|COMP|6040-0|LNC|House dust Bencard Ab.IgE|House dust Bencard Ab.IgE
C0362647|T201|COMP|6041-8|LNC|Cynodon dactylon Ab.IgE|Cynodon dactylon Ab.IgE
C0362648|T201|COMP|6042-6|LNC|Beta lactoglobulin MF77 Ab.IgE|Beta lactoglobulin MF77 Ab.IgE
C0362649|T201|COMP|6043-4|LNC|Birch Ab.IgE|Birch Ab.IgE
C0362650|T201|COMP|6044-2|LNC|Monomorium minimum Ab.IgE|Monomorium minimum Ab.IgE
C0362651|T201|COMP|6045-9|LNC|Piper nigrum Ab.IgE|Piper nigrum Ab.IgE
C0362653|T201|COMP|6047-5|LNC|Chironomus thummi Ab.IgE|Chironomus thummi Ab.IgE
C0362654|T201|COMP|6048-3|LNC|Mytilus edulis Ab.IgE|Mytilus edulis Ab.IgE
C0362655|T201|COMP|6049-1|LNC|Botrytis cinerea Ab.IgE|Botrytis cinerea Ab.IgE
C0362656|T201|COMP|6050-9|LNC|Bertholletia excelsa Ab.IgE|Bertholletia excelsa Ab.IgE
C0362657|T201|COMP|6051-7|LNC|Yeast brewer's Ab.IgE|Yeast brewer's Ab.IgE
C0362658|T201|COMP|6052-5|LNC|Brassica oleracea var italica Ab.IgE|Brassica oleracea var italica Ab.IgE
C0362659|T201|COMP|6053-3|LNC|Bromus inermis Ab.IgE|Bromus inermis Ab.IgE
C0362660|T201|COMP|6054-1|LNC|Fagopyrum esculentum Ab.IgE|Fagopyrum esculentum Ab.IgE
C0362661|T201|COMP|6055-8|LNC|Budgerigar feather Ab.IgE|Budgerigar feather Ab.IgE
C0362662|T201|COMP|6056-6|LNC|Bombus terrestris Ab.IgE|Bombus terrestris Ab.IgE
C0362663|T201|COMP|6057-4|LNC|Matricaria chamomilla Ab.IgE|Matricaria chamomilla Ab.IgE
C0362664|T201|COMP|6058-2|LNC|Phalaris arundinacea Ab.IgE|Phalaris arundinacea Ab.IgE
C0362665|T201|COMP|6059-0|LNC|Candida albicans Ab.IgE|Candida albicans Ab.IgE
C0362667|T201|COMP|6061-6|LNC|Daucus carota Ab.IgE|Daucus carota Ab.IgE
C0362668|T201|COMP|6062-4|LNC|Casein Ab.IgE|Casein Ab.IgE
C0362669|T201|COMP|6063-2|LNC|Ricinus communis Ab.IgE|Ricinus communis Ab.IgE
C0362671|T201|COMP|6065-7|LNC|Apium graveolens Ab.IgE|Apium graveolens Ab.IgE
C0362672|T201|COMP|6066-5|LNC|Acremonium sp Ab.IgE|Acremonium sp Ab.IgE
C0362673|T201|COMP|6067-3|LNC|Cheese cheddar type Ab.IgE|Cheese cheddar type Ab.IgE
C0362674|T201|COMP|6068-1|LNC|Cheese mold type Ab.IgE|Cheese mold type Ab.IgE
C0362675|T201|COMP|6069-9|LNC|Castanea sativa pollen Ab.IgE|Castanea sativa pollen Ab.IgE
C0362676|T201|COMP|6070-7|LNC|Chicken feather Ab.IgE|Chicken feather Ab.IgE
C0362677|T201|COMP|6071-5|LNC|Chicken meat Ab.IgE|Chicken meat Ab.IgE
C0362678|T201|COMP|6072-3|LNC|Chloramin T Ab.IgE|Chloramin T Ab.IgE
C0362679|T201|COMP|6073-1|LNC|Chocolate Ab.IgE|Chocolate Ab.IgE
C0362680|T201|COMP|6074-9|LNC|Chymopapain Ab.IgE|Chymopapain Ab.IgE
C0362681|T201|COMP|6075-6|LNC|Cladosporium herbarum Ab.IgE|Cladosporium herbarum Ab.IgE
C0362682|T201|COMP|6076-4|LNC|Ruditapes spp Ab.IgE|Ruditapes spp Ab.IgE
C0362683|T201|COMP|6077-2|LNC|Xanthium commune Ab.IgE|Xanthium commune Ab.IgE
C0362684|T201|COMP|6078-0|LNC|Blatella germanica Ab.IgE|Blatella germanica Ab.IgE
C0362685|T201|COMP|6080-6|LNC|Theobroma cacao Ab.IgE|Theobroma cacao Ab.IgE
C0362686|T201|COMP|6081-4|LNC|Cocos nucifera Ab.IgE|Cocos nucifera Ab.IgE
C0362687|T201|COMP|6082-2|LNC|Gadus morhua Ab.IgE|Gadus morhua Ab.IgE
C0362688|T201|COMP|6083-0|LNC|Coffea spp Ab.IgE|Coffea spp Ab.IgE
C0362689|T201|COMP|6084-8|LNC|Colza Ab.IgE|Colza Ab.IgE
C0362690|T201|COMP|6085-5|LNC|Ambrosia elatior Ab.IgE|Ambrosia elatior Ab.IgE
C0362691|T201|COMP|6087-1|LNC|Zea mays Ab.IgE|Zea mays Ab.IgE
C0362692|T201|COMP|6088-9|LNC|Cotton cultivated Ab.IgE|Cotton cultivated Ab.IgE
C0362693|T201|COMP|6089-7|LNC|Cottonseed Ab.IgE|Cottonseed Ab.IgE
C0362694|T201|COMP|6090-5|LNC|Populus deltoides Ab.IgE|Populus deltoides Ab.IgE
C0362695|T201|COMP|6091-3|LNC|Cow dander Ab.IgE|Cow dander Ab.IgE
C0362696|T201|COMP|6092-1|LNC|Cancer pagurus Ab.IgE|Cancer pagurus Ab.IgE
C0362697|T201|COMP|6094-7|LNC|Curvularia lunata Ab.IgE|Curvularia lunata Ab.IgE
C0362698|T201|COMP|6097-0|LNC|Taraxacum vulgare Ab.IgE|Taraxacum vulgare Ab.IgE
C0362699|T201|COMP|6095-4|LNC|Dermatophagoides farinae Ab.IgE|Dermatophagoides farinae Ab.IgE
C0362700|T201|COMP|6096-2|LNC|Dermatophagoides pteronyssinus Ab.IgE|Dermatophagoides pteronyssinus Ab.IgE
C0362701|T201|COMP|6098-8|LNC|Dog dander Ab.IgE|Dog dander Ab.IgE
C0362702|T201|COMP|6099-6|LNC|Dog epithelium Ab.IgE|Dog epithelium Ab.IgE
C0362703|T201|COMP|6100-2|LNC|Duck feather Ab.IgE|Duck feather Ab.IgE
C0362704|T201|COMP|6101-0|LNC|Duck meat Ab.IgE|Duck meat Ab.IgE
C0362705|T201|COMP|6102-8|LNC|Dust profile Ab.IgE|Dust profile Ab.IgE
C0362706|T201|COMP|6103-6|LNC|Echinococcus sp Ab.IgE|Echinococcus sp Ab.IgE
C0362707|T201|COMP|6105-1|LNC|Anguilla anguilla Ab.IgE|Anguilla anguilla Ab.IgE
C0362708|T201|COMP|6106-9|LNC|Egg white Ab.IgE|Egg white Ab.IgE
C0362709|T201|COMP|6107-7|LNC|Egg yolk Ab.IgE|Egg yolk Ab.IgE
C0362712|T201|COMP|6110-1|LNC|Plantago lanceolata Ab.IgE|Plantago lanceolata Ab.IgE
C0362714|T201|COMP|6112-7|LNC|Ethylene oxide Ab.IgE|Ethylene oxide Ab.IgE
C0362715|T201|COMP|6113-5|LNC|Eucalyptus spp Ab.IgE|Eucalyptus spp Ab.IgE
C0362716|T201|COMP|6114-3|LNC|Euroglyphus maynei Ab.IgE|Euroglyphus maynei Ab.IgE
C0362717|T201|COMP|6115-0|LNC|Franseria acanthicarpa Ab.IgE|Franseria acanthicarpa Ab.IgE
C0362718|T201|COMP|6116-8|LNC|Ficus sp Ab.IgE|Ficus sp Ab.IgE
C0362721|T201|COMP|6119-2|LNC|Formaldehyde Ab.IgE|Formaldehyde Ab.IgE
C0362722|T201|COMP|6120-0|LNC|Fusarium culmorum Ab.IgE|Fusarium culmorum Ab.IgE
C0362724|T201|COMP|6122-6|LNC|Allium sativum Ab.IgE|Allium sativum Ab.IgE
C0362725|T201|COMP|6123-4|LNC|Pelargonium sp Ab.IgE|Pelargonium sp Ab.IgE
C0362727|T201|COMP|6125-9|LNC|Gluten Ab.IgE|Gluten Ab.IgE
C0362728|T201|COMP|6126-7|LNC|Glycyphagus domesticus Ab.IgE|Glycyphagus domesticus Ab.IgE
C0362729|T201|COMP|6127-5|LNC|Goat epithelium Ab.IgE|Goat epithelium Ab.IgE
C0362730|T201|COMP|6128-3|LNC|Solidago virgaurea Ab.IgE|Solidago virgaurea Ab.IgE
C0362731|T201|COMP|6129-1|LNC|Goose feather Ab.IgE|Goose feather Ab.IgE
C0362732|T201|COMP|6130-9|LNC|Goose meat Ab.IgE|Goose meat Ab.IgE
C0362733|T201|COMP|6131-7|LNC|Citrus paradisis Ab.IgE|Citrus paradisis Ab.IgE
C0362734|T201|COMP|6132-5|LNC|Coffee bean green Ab.IgE|Coffee bean green Ab.IgE
C0362735|T201|COMP|6133-3|LNC|Cladotanytarsus lewisi Ab.IgE|Cladotanytarsus lewisi Ab.IgE
C0362736|T201|COMP|6134-1|LNC|Guinea pig epithelium Ab.IgE|Guinea pig epithelium Ab.IgE
C0362737|T201|COMP|6135-8|LNC|Hamster epithelium Ab.IgE|Hamster epithelium Ab.IgE
C0362738|T201|COMP|6136-6|LNC|Corylus avellana Ab.IgE|Corylus avellana Ab.IgE
C0362739|T201|COMP|6137-4|LNC|Corylus avellana pollen Ab.IgE|Corylus avellana pollen Ab.IgE
C0362740|T201|COMP|6138-2|LNC|Setomelanomma rostrata Ab.IgE|Setomelanomma rostrata Ab.IgE
C0362741|T201|COMP|6139-0|LNC|Clupea harengus Ab.IgE|Clupea harengus Ab.IgE
C0362742|T201|COMP|6140-8|LNC|Hickory Ab.IgE|Hickory Ab.IgE
C0362743|T201|COMP|6141-6|LNC|Humulus lupus Ab.IgE|Humulus lupus Ab.IgE
C0362744|T201|COMP|6142-4|LNC|Hornet venom Ab.IgE|Hornet venom Ab.IgE
C0362745|T201|COMP|6143-2|LNC|Horse dander Ab.IgE|Horse dander Ab.IgE
C0362747|T201|COMP|6145-7|LNC|House dust Ab.IgE|House dust Ab.IgE
C0362748|T201|COMP|6147-3|LNC|Insulin bovine Ab.IgE|Insulin bovine Ab.IgE
C0362749|T201|COMP|6148-1|LNC|Insulin human Ab.IgE|Insulin human Ab.IgE
C0362750|T201|COMP|6149-9|LNC|Insulin porcine Ab.IgE|Insulin porcine Ab.IgE
C0362751|T201|COMP|6150-7|LNC|Ispaghula laxative Ab.IgE|Ispaghula laxative Ab.IgE
C0362752|T201|COMP|6151-5|LNC|Cupressus sempervirens Ab.IgE|Cupressus sempervirens Ab.IgE
C0362753|T201|COMP|6152-3|LNC|Sorghum halepense Ab.IgE|Sorghum halepense Ab.IgE
C0362754|T201|COMP|6153-1|LNC|Poa pratensis Ab.IgE|Poa pratensis Ab.IgE
C0362755|T201|COMP|6154-9|LNC|Actinidia chinensis Ab.IgE|Actinidia chinensis Ab.IgE
C0362756|T201|COMP|6155-6|LNC|Lamb Ab.IgE|Lamb Ab.IgE
C0362757|T201|COMP|6157-2|LNC|Mutton Ab.IgE|Mutton Ab.IgE
C0362758|T201|COMP|6156-4|LNC|Chenopodium album Ab.IgE|Chenopodium album Ab.IgE
C0362759|T201|COMP|6158-0|LNC|Latex Ab.IgE|Latex Ab.IgE
C0362760|T201|COMP|6159-8|LNC|Citrus limon Ab.IgE|Citrus limon Ab.IgE
C0362762|T201|COMP|6161-4|LNC|Lactuca sativa Ab.IgE|Lactuca sativa Ab.IgE
C0362763|T201|COMP|6162-2|LNC|Syringa vulgaris Ab.IgE|Syringa vulgaris Ab.IgE
C0362764|T201|COMP|6163-0|LNC|Citrus aurantifolia tree Ab.IgE|Citrus aurantifolia tree Ab.IgE
C0362766|T201|COMP|6165-5|LNC|Homarus gammarus Ab.IgE|Homarus gammarus Ab.IgE
C0362767|T201|COMP|6166-3|LNC|Malt Ab.IgE|Malt Ab.IgE
C0362768|T201|COMP|6167-1|LNC|Mangifera indica Ab.IgE|Mangifera indica Ab.IgE
C0362769|T201|COMP|6168-9|LNC|Maple Ab.IgE|Maple Ab.IgE
C0362771|T201|COMP|6170-5|LNC|Alopercurus pratensis Ab.IgE|Alopercurus pratensis Ab.IgE
C0362772|T201|COMP|6171-3|LNC|Melaleuca leucadendron Ab.IgE|Melaleuca leucadendron Ab.IgE
C0362774|T201|COMP|6173-9|LNC|Prosopis juliflora Ab.IgE|Prosopis juliflora Ab.IgE
C0362775|T201|COMP|6174-7|LNC|Milk Ab.IgE|Milk Ab.IgE
C0362776|T201|COMP|6175-4|LNC|Panicum milliaceum Ab.IgE|Panicum milliaceum Ab.IgE
C0362777|T201|COMP|6176-2|LNC|Mimosa spp Ab.IgE|Mimosa spp Ab.IgE
C0362778|T201|COMP|6177-0|LNC|Aedes communis Ab.IgE|Aedes communis Ab.IgE
C0362779|T201|COMP|6178-8|LNC|Juniperus sabinoides Ab.IgE|Juniperus sabinoides Ab.IgE
C0362780|T201|COMP|6179-6|LNC|Mouse epithelium Ab.IgE|Mouse epithelium Ab.IgE
C0362781|T201|COMP|6180-4|LNC|Mouse serum proteins Ab.IgE|Mouse serum proteins Ab.IgE
C0362782|T201|COMP|6181-2|LNC|Mouse urine proteins Ab.IgE|Mouse urine proteins Ab.IgE
C0362783|T201|COMP|6182-0|LNC|Mucor racemosus Ab.IgE|Mucor racemosus Ab.IgE
C0362784|T201|COMP|6183-8|LNC|Artemisia vulgaris Ab.IgE|Artemisia vulgaris Ab.IgE
C0362785|T201|COMP|6184-6|LNC|Mussel Ab.IgE|Mussel Ab.IgE
C0362786|T201|COMP|6185-3|LNC|Mustard Ab.IgE|Mustard Ab.IgE
C0362787|T201|COMP|6186-1|LNC|Urtica dioica Ab.IgE|Urtica dioica Ab.IgE
C0362788|T201|COMP|6187-9|LNC|Neurospora sitophila Ab.IgE|Neurospora sitophila Ab.IgE
C0362789|T201|COMP|6188-7|LNC|Nutmeg Ab.IgE|Nutmeg Ab.IgE
C0362792|T201|COMP|6093-9|LNC|Avena sativa cultivated Ab.IgE|Avena sativa cultivated Ab.IgE
C0362793|T201|COMP|6192-9|LNC|Olea europaea pollen Ab.IgE|Olea europaea pollen Ab.IgE
C0362794|T201|COMP|6193-7|LNC|Allium cepa Ab.IgE|Allium cepa Ab.IgE
C0362795|T201|COMP|6194-5|LNC|Citrus sinensis Ab.IgE|Citrus sinensis Ab.IgE
C0362796|T201|COMP|6195-2|LNC|Dactylis glomerata Ab.IgE|Dactylis glomerata Ab.IgE
C0362797|T201|COMP|6196-0|LNC|Chrysanthemum leucanthemum Ab.IgE|Chrysanthemum leucanthemum Ab.IgE
C0362798|T201|COMP|6197-8|LNC|Paecilomyces sp Ab.IgE|Paecilomyces sp Ab.IgE
C0362800|T201|COMP|6199-4|LNC|Parietaria judaica Ab.IgE|Parietaria judaica Ab.IgE
C0362801|T201|COMP|6200-0|LNC|Parietaria officinalis Ab.IgE|Parietaria officinalis Ab.IgE
C0362802|T201|COMP|6201-8|LNC|Parrot droppings Ab.IgE|Parrot droppings Ab.IgE
C0362803|T201|COMP|6202-6|LNC|Parrot feather Ab.IgE|Parrot feather Ab.IgE
C0362804|T201|COMP|6203-4|LNC|Petroselinum crispum Ab.IgE|Petroselinum crispum Ab.IgE
C0362805|T201|COMP|6204-2|LNC|Pisum sativum Ab.IgE|Pisum sativum Ab.IgE
C0362806|T201|COMP|6205-9|LNC|Prunus persica Ab.IgE|Prunus persica Ab.IgE
C0362807|T201|COMP|6206-7|LNC|Arachis hypogaea Ab.IgE|Arachis hypogaea Ab.IgE
C0362808|T201|COMP|6207-5|LNC|Pyrus communis Ab.IgE|Pyrus communis Ab.IgE
C0362811|T201|COMP|6210-9|LNC|Penicillin V Ab.IgE|Penicillin V Ab.IgE
C0362812|T201|COMP|6211-7|LNC|Penicillium brevicompactum Ab.IgE|Penicillium brevicompactum Ab.IgE
C0362813|T201|COMP|6212-5|LNC|Penicillium notatum Ab.IgE|Penicillium notatum Ab.IgE
C0362814|T201|COMP|6213-3|LNC|Schinus molle Ab.IgE|Schinus molle Ab.IgE
C0362815|T201|COMP|6214-1|LNC|Perca spp Ab.IgE|Perca spp Ab.IgE
C0362816|T201|COMP|6215-8|LNC|Lolium perenne Ab.IgE|Lolium perenne Ab.IgE
C0362816|T201|COMP|7371-8|LNC|Lolium perenne Ab.IgE|Lolium perenne Ab.IgE
C0362816|T201|COMP|7372-6|LNC|Lolium perenne Ab.IgE|Lolium perenne Ab.IgE
C0362817|T201|COMP|6216-6|LNC|Phoma betae Ab.IgE|Phoma betae Ab.IgE
C0362818|T201|COMP|6217-4|LNC|Pigeon droppings Ab.IgE|Pigeon droppings Ab.IgE
C0362819|T201|COMP|6218-2|LNC|Ananas comosus Ab.IgE|Ananas comosus Ab.IgE
C0362820|T201|COMP|6219-0|LNC|Pork Ab.IgE|Pork Ab.IgE
C0362822|T201|COMP|6221-6|LNC|Primrose Ab.IgE|Primrose Ab.IgE
C0362823|T201|COMP|6222-4|LNC|Syagrus romanzoffianum Ab.IgE|Syagrus romanzoffianum Ab.IgE
C0362824|T201|COMP|6223-2|LNC|Rabbit epithelium Ab.IgE|Rabbit epithelium Ab.IgE
C0362825|T201|COMP|6224-0|LNC|Rat epithelium Ab.IgE|Rat epithelium Ab.IgE
C0362826|T201|COMP|6225-7|LNC|Rat serum proteins Ab.IgE|Rat serum proteins Ab.IgE
C0362827|T201|COMP|6226-5|LNC|Rat urine proteins Ab.IgE|Rat urine proteins Ab.IgE
C0362828|T201|COMP|6227-3|LNC|Pepper red Ab.IgE|Pepper red Ab.IgE
C0362830|T201|COMP|6229-9|LNC|Rhizopus nigricans Ab.IgE|Rhizopus nigricans Ab.IgE
C0362831|T201|COMP|6230-7|LNC|Oryza sativa Ab.IgE|Oryza sativa Ab.IgE
C0362832|T201|COMP|6231-5|LNC|Rosa spp hip Ab.IgE|Rosa spp hip Ab.IgE
C0362833|T201|COMP|6232-3|LNC|Iva ciliata Ab.IgE|Iva ciliata Ab.IgE
C0362834|T201|COMP|6233-1|LNC|Pigweed rough Ab.IgE|Pigweed rough Ab.IgE
C0362835|T201|COMP|6234-9|LNC|Salsola kali Ab.IgE|Salsola kali Ab.IgE
C0362836|T201|COMP|7674-5|LNC|Secale cereale Ab.IgE|Secale cereale Ab.IgE
C0362838|T201|COMP|6237-2|LNC|Salmo salar Ab.IgE|Salmo salar Ab.IgE
C0362839|T201|COMP|6238-0|LNC|Distichlis spicata Ab.IgE|Distichlis spicata Ab.IgE
C0362841|T201|COMP|6240-6|LNC|Seminal fluid Ab.IgE|Seminal fluid Ab.IgE
C0362842|T201|COMP|6241-4|LNC|Serpula lacrymans Ab.IgE|Serpula lacrymans Ab.IgE
C0362843|T201|COMP|6242-2|LNC|Sesamum indicum Ab.IgE|Sesamum indicum Ab.IgE
C0362844|T201|COMP|6243-0|LNC|Sheep epithelium Ab.IgE|Sheep epithelium Ab.IgE
C0362845|T201|COMP|6244-8|LNC|Rumex acetosella Ab.IgE|Rumex acetosella Ab.IgE
C0362846|T201|COMP|6245-5|LNC|Sheep wool Ab.IgE|Sheep wool Ab.IgE
C0362847|T201|COMP|6246-3|LNC|Pandalus borealis Ab.IgE|Pandalus borealis Ab.IgE
C0362848|T201|COMP|6247-1|LNC|Silk Ab.IgE|Silk Ab.IgE
C0362850|T201|COMP|6249-7|LNC|Palinurus spp Ab.IgE|Palinurus spp Ab.IgE
C0362851|T201|COMP|6250-5|LNC|Pigweed spiny Ab.IgE|Pigweed spiny Ab.IgE
C0362852|T201|COMP|6251-3|LNC|Sporobolomyces roseus Ab.IgE|Sporobolomyces roseus Ab.IgE
C0362853|T201|COMP|6252-1|LNC|Stemphylium botryosum Ab.IgE|Stemphylium botryosum Ab.IgE
C0362855|T201|COMP|6254-7|LNC|Acarus siro Ab.IgE|Acarus siro Ab.IgE
C0362856|T201|COMP|6160-6|LNC|Lepidoglyphus destructor Ab.IgE|Lepidoglyphus destructor Ab.IgE
C0362857|T201|COMP|6256-2|LNC|Tyrophagus putrescentiae Ab.IgE|Tyrophagus putrescentiae Ab.IgE
C0362858|T201|COMP|6257-0|LNC|Fragaria vesca Ab.IgE|Fragaria vesca Ab.IgE
C0362862|T201|COMP|6261-2|LNC|Anthoxanthum odoratum Ab.IgE|Anthoxanthum odoratum Ab.IgE
C0362863|T201|COMP|6262-0|LNC|Swine epithelium Ab.IgE|Swine epithelium Ab.IgE
C0362865|T201|COMP|6264-6|LNC|Camellia sinensis Ab.IgE|Camellia sinensis Ab.IgE
C0362866|T201|COMP|6265-3|LNC|Phleum pratense Ab.IgE|Phleum pratense Ab.IgE
C0362867|T201|COMP|6266-1|LNC|Lycopersicon lycopersicum Ab.IgE|Lycopersicon lycopersicum Ab.IgE
C0362868|T201|COMP|6267-9|LNC|Trichoderma viride Ab.IgE|Trichoderma viride Ab.IgE
C0362869|T201|COMP|6268-7|LNC|Oncorhynchus mykiss Ab.IgE|Oncorhynchus mykiss Ab.IgE
C0362870|T201|COMP|6269-5|LNC|Tulipa spp Ab.IgE|Tulipa spp Ab.IgE
C0362871|T201|COMP|6270-3|LNC|Thunnus albacares Ab.IgE|Thunnus albacares Ab.IgE
C0362872|T201|COMP|6271-1|LNC|Turkey meat Ab.IgE|Turkey meat Ab.IgE
C0362873|T201|COMP|6272-9|LNC|Holcus lanatus Ab.IgE|Holcus lanatus Ab.IgE
C0362874|T201|COMP|6273-7|LNC|Juglans spp Ab.IgE|Juglans spp Ab.IgE
C0362875|T201|COMP|6274-5|LNC|Juglans california Ab.IgE|Juglans california Ab.IgE
C0362876|T201|COMP|6275-2|LNC|Ambrosia psilostachya Ab.IgE|Ambrosia psilostachya Ab.IgE
C0362877|T201|COMP|6276-0|LNC|Triticum aestivum Ab.IgE|Triticum aestivum Ab.IgE
C0362879|T201|COMP|6278-6|LNC|Fraxinus americana Ab.IgE|Fraxinus americana Ab.IgE
C0362880|T201|COMP|6279-4|LNC|Bean white Ab.IgE|Bean white Ab.IgE
C0362881|T201|COMP|6280-2|LNC|Dolichovespula maculata Ab.IgE|Dolichovespula maculata Ab.IgE
C0362884|T201|COMP|16922-7|LNC|Elymus triticoides Ab.IgE|Elymus triticoides Ab.IgE
C0362885|T201|COMP|6284-4|LNC|Silk wild Ab.IgE|Silk wild Ab.IgE
C0362886|T201|COMP|6285-1|LNC|Salix caprea Ab.IgE|Salix caprea Ab.IgE
C0362887|T201|COMP|6286-9|LNC|Artemisia absinthium Ab.IgE|Artemisia absinthium Ab.IgE
C0362888|T201|COMP|6287-7|LNC|Saccharomyces cerevisiae Ab.IgE|Saccharomyces cerevisiae Ab.IgE
C0362889|T201|COMP|6288-5|LNC|Dolichovespula arenaria Ab.IgE|Dolichovespula arenaria Ab.IgE
C0362890|T201|COMP|702-1|LNC|Anisocytosis|Anisocytosis
C0362891|T201|COMP|703-9|LNC|Basophilic stippling|Basophilic stippling
C0362892|T201|COMP|704-7|LNC|Basophils|Basophils
C0362893|T201|COMP|705-4|LNC|Basophils|Basophils
C0362894|T201|COMP|706-2|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0362895|T201|COMP|707-0|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0362896|T201|COMP|708-8|LNC|Blasts|Blasts
C0362897|T201|COMP|709-6|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C0362898|T201|COMP|5909-7|LNC|Blood smear finding|Blood smear finding
C0362899|T201|COMP|710-4|LNC|Blood smear finding positive|Blood smear finding positive
C0362900|T201|COMP|711-2|LNC|Eosinophils|Eosinophils
C0362901|T201|COMP|712-0|LNC|Eosinophils|Eosinophils
C0362902|T201|COMP|713-8|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0362903|T201|COMP|714-6|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0362904|T201|COMP|715-3|LNC|Normoblasts|Normoblasts
C0362905|T201|COMP|784-9|LNC|Erythrocyte mean corpuscular diameter|Erythrocyte mean corpuscular diameter
C0362906|T201|COMP|785-6|LNC|Erythrocyte mean corpuscular hemoglobin|Erythrocyte mean corpuscular hemoglobin
C0362908|T201|COMP|787-2|LNC|Erythrocyte mean corpuscular volume|Erythrocyte mean corpuscular volume
C0362909|T201|COMP|788-0|LNC|Erythrocyte distribution width|Erythrocyte distribution width
C0362910|T201|COMP|789-8|LNC|Erythrocytes|Erythrocytes
C0362911|T201|COMP|790-6|LNC|Erythrocytes|Erythrocytes
C0362912|T201|COMP|791-4|LNC|Erythrocytes|Erythrocytes
C0362913|T201|COMP|792-2|LNC|Erythrocytes|Erythrocytes
C0362914|T201|COMP|794-8|LNC|Erythrocytes|Erythrocytes
C0362915|T201|COMP|793-0|LNC|Erythrocytes|Erythrocytes
C0362916|T201|COMP|795-5|LNC|Erythrocytes|Erythrocytes
C0362917|T201|COMP|796-3|LNC|Erythrocytes|Erythrocytes
C0362918|T201|COMP|797-1|LNC|Erythrocytes|Erythrocytes
C0362919|T201|COMP|798-9|LNC|Erythrocytes|Erythrocytes
C0362920|T201|COMP|799-7|LNC|Erythrocytes|Erythrocytes
C0362921|T201|COMP|716-1|LNC|Heinz bodies|Heinz bodies
C0362922|T201|COMP|717-9|LNC|Hemoglobin|Hemoglobin
C0362923|T201|COMP|718-7|LNC|Hemoglobin|Hemoglobin
C0362924|T201|COMP|719-5|LNC|Hemoglobin|Hemoglobin
C0362925|T201|COMP|720-3|LNC|Hemoglobin.free|Hemoglobin.free
C0362926|T201|COMP|721-1|LNC|Hemoglobin.free|Hemoglobin.free
C0362927|T201|COMP|722-9|LNC|Hemoglobin|Hemoglobin
C0362928|T201|COMP|723-7|LNC|Hemoglobin|Hemoglobin
C0362929|T201|COMP|724-5|LNC|Hemoglobin|Hemoglobin
C0362930|T201|COMP|725-2|LNC|Hemoglobin|Hemoglobin
C0362931|T201|COMP|726-0|LNC|Hemoglobin|Hemoglobin
C0362932|T201|COMP|727-8|LNC|Hemoglobin distribution width|Hemoglobin distribution width
C0362933|T201|COMP|728-6|LNC|Hypochromia|Hypochromia
C0362934|T201|COMP|804-5|LNC|Leukocytes|Leukocytes
C0362935|T201|COMP|805-2|LNC|Leukocytes|Leukocytes
C0362936|T201|COMP|806-0|LNC|Leukocytes|Leukocytes
C0362937|T201|COMP|807-8|LNC|Leukocytes|Leukocytes
C0362938|T201|COMP|808-6|LNC|Leukocytes|Leukocytes
C0362939|T201|COMP|809-4|LNC|Leukocytes|Leukocytes
C0362940|T201|COMP|810-2|LNC|Leukocytes|Leukocytes
C0362941|T201|COMP|811-0|LNC|Leukocytes|Leukocytes
C0362942|T201|COMP|812-8|LNC|Leukocytes|Leukocytes
C0362943|T201|COMP|813-6|LNC|Leukocytes|Leukocytes
C0362944|T201|COMP|814-4|LNC|Leukocytes|Leukocytes
C0362945|T201|COMP|729-4|LNC|Leukocytes other|Leukocytes other
C0362946|T201|COMP|730-2|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0362947|T201|COMP|731-0|LNC|Lymphocytes|Lymphocytes
C0362948|T201|COMP|732-8|LNC|Lymphocytes|Lymphocytes
C0362949|T201|COMP|733-6|LNC|Lymphocytes.variant|Lymphocytes.variant
C0362950|T201|COMP|734-4|LNC|Lymphocytes.variant|Lymphocytes.variant
C0362951|T201|COMP|735-1|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C0362952|T201|COMP|736-9|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0362953|T201|COMP|737-7|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0362954|T201|COMP|738-5|LNC|Macrocytes|Macrocytes
C0362955|T201|COMP|739-3|LNC|Metamyelocytes|Metamyelocytes
C0362956|T201|COMP|740-1|LNC|Metamyelocytes/100 leukocytes|Metamyelocytes/100 leukocytes
C0362957|T201|COMP|741-9|LNC|Microcytes|Microcytes
C0362958|T201|COMP|742-7|LNC|Monocytes|Monocytes
C0362959|T201|COMP|743-5|LNC|Monocytes|Monocytes
C0362960|T201|COMP|5905-5|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0362961|T201|COMP|744-3|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0362962|T201|COMP|745-0|LNC|Myeloblasts|Myeloblasts
C0362963|T201|COMP|746-8|LNC|Myeloblasts|Myeloblasts
C0362964|T201|COMP|747-6|LNC|Myeloblasts/100 leukocytes|Myeloblasts/100 leukocytes
C0362965|T201|COMP|748-4|LNC|Myelocytes|Myelocytes
C0362966|T201|COMP|750-0|LNC|Myelocytes/100 leukocytes|Myelocytes/100 leukocytes
C0362967|T201|COMP|749-2|LNC|Myelocytes/100 leukocytes|Myelocytes/100 leukocytes
C0362968|T201|COMP|751-8|LNC|Neutrophils|Neutrophils
C0362969|T201|COMP|753-4|LNC|Neutrophils|Neutrophils
C0362970|T201|COMP|754-2|LNC|Neutrophils|Neutrophils
C0362971|T201|COMP|755-9|LNC|Neutrophils|Neutrophils
C0362972|T201|COMP|756-7|LNC|Neutrophils|Neutrophils
C0362973|T201|COMP|757-5|LNC|Neutrophils|Neutrophils
C0362974|T201|COMP|758-3|LNC|Neutrophils|Neutrophils
C0362975|T201|COMP|759-1|LNC|Neutrophils|Neutrophils
C0362976|T201|COMP|5906-3|LNC|Neutrophils|Neutrophils
C0362977|T201|COMP|760-9|LNC|Neutrophils|Neutrophils
C0362978|T201|COMP|761-7|LNC|Neutrophils|Neutrophils
C0362979|T201|COMP|762-5|LNC|Neutrophils|Neutrophils
C0362980|T201|COMP|763-3|LNC|Neutrophils.band form|Neutrophils.band form
C0362981|T201|COMP|764-1|LNC|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0362982|T201|COMP|765-8|LNC|Neutrophils.hypersegmented|Neutrophils.hypersegmented
C0362983|T201|COMP|766-6|LNC|Neutrophils.hypersegmented|Neutrophils.hypersegmented
C0362984|T201|COMP|767-4|LNC|Neutrophils.hypersegmented/100 leukocytes|Neutrophils.hypersegmented/100 leukocytes
C0362985|T201|COMP|768-2|LNC|Neutrophils.segmented|Neutrophils.segmented
C0362986|T201|COMP|769-0|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C0362987|T201|COMP|770-8|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0362988|T201|COMP|771-6|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C0362989|T201|COMP|772-4|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C0362990|T201|COMP|773-2|LNC|Erythrocytes.nucleated/100 erythrocytes|Erythrocytes.nucleated/100 erythrocytes
C0362991|T201|COMP|774-0|LNC|Ovalocytes|Ovalocytes
C0362992|T201|COMP|775-7|LNC|Platelet mean diameter|Platelet mean diameter
C0362993|T201|COMP|776-5|LNC|Platelet mean volume|Platelet mean volume
C0362994|T201|COMP|777-3|LNC|Platelets|Platelets
C0362995|T201|COMP|778-1|LNC|Platelets|Platelets
C0362996|T201|COMP|5908-9|LNC|Platelets.giant|Platelets.giant
C0362997|T201|COMP|7791-7|LNC|Dacryocytes|Dacryocytes
C0362998|T201|COMP|780-7|LNC|Promyelocytes|Promyelocytes
C0362999|T201|COMP|781-5|LNC|Promyelocytes|Promyelocytes
C0363000|T201|COMP|782-3|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C0363002|T201|COMP|800-3|LNC|Schistocytes|Schistocytes
C0363003|T201|COMP|801-1|LNC|Sickle cells|Sickle cells
C0363004|T201|COMP|802-9|LNC|Spherocytes|Spherocytes
C0363005|T201|COMP|803-7|LNC|Toxic granules|Toxic granules
C0363075|T201|COMP|884-7|LNC|ABO & Rh group|ABO & Rh group
C0363081|T201|COMP|890-4|LNC|Blood group antibody screen|Blood group antibody screen
C0363084|T201|COMP|893-8|LNC|Blood group antibody screen.autologous|Blood group antibody screen.autologous
C0363085|T201|COMP|894-6|LNC|Blood group antibody screen.cell II|Blood group antibody screen.cell II
C0363086|T201|COMP|895-3|LNC|Blood group antibody screen.cells I+II+III|Blood group antibody screen.cells I+II+III
C0363087|T201|COMP|896-1|LNC|Blood group antibody screen|Blood group antibody screen
C0363088|T201|COMP|897-9|LNC|Blood group antibody screen|Blood group antibody screen
C0363089|T201|COMP|898-7|LNC|Blood group antibody screen.cell I|Blood group antibody screen.cell I
C0363090|T201|COMP|899-5|LNC|Blood group antibody screen.cell II|Blood group antibody screen.cell II
C0363091|T201|COMP|900-1|LNC|Blood group antibody screen.cell III|Blood group antibody screen.cell III
C0363092|T201|COMP|901-9|LNC|Blood group antibody screen.cells I+II+III|Blood group antibody screen.cells I+II+III
C0363093|T201|COMP|902-7|LNC|Blood group antibody screen.autologous|Blood group antibody screen.autologous
C0363094|T201|COMP|903-5|LNC|Blood group antibody screen|Blood group antibody screen
C0363095|T201|COMP|904-3|LNC|Blood group antibody screen|Blood group antibody screen
C0363115|T201|COMP|923-3|LNC|Blood collection bag lot identifier|Blood collection bag lot identifier
C0363116|T201|COMP|924-1|LNC|Blood product dispensed|Blood product dispensed
C0363117|T201|COMP|925-8|LNC|Blood product disposition|Blood product disposition
C0363118|T201|COMP|926-6|LNC|Blood product.other given|Blood product.other given
C0363119|T201|COMP|927-4|LNC|Blood product identifier.pooled|Blood product identifier.pooled
C0363120|T201|COMP|928-2|LNC|Blood product reaction|Blood product reaction
C0363121|T201|COMP|929-0|LNC|Blood product release time|Blood product release time
C0363122|T201|COMP|930-8|LNC|Blood product reservation|Blood product reservation
C0363123|T201|COMP|931-6|LNC|Blood product source|Blood product source
C0363124|T201|COMP|932-4|LNC|Blood product type|Blood product type
C0363126|T201|COMP|934-0|LNC|Blood product unit ID|Blood product unit ID
C0363127|T201|COMP|935-7|LNC|Blood product unit expiration|Blood product unit expiration
C0363128|T201|COMP|936-5|LNC|Blood product unit identifier|Blood product unit identifier
C0363153|T201|COMP|943-1|LNC|C Ab|C Ab
C0363154|T201|COMP|944-9|LNC|C Ab|C Ab
C0363155|T201|COMP|945-6|LNC|C Ab|C Ab
C0363156|T201|COMP|946-4|LNC|C Ag|C Ag
C0363157|T201|COMP|947-2|LNC|C Ag|C Ag
C0363158|T201|COMP|948-0|LNC|C Ag|C Ag
C0363183|T201|COMP|1304-5|LNC|D Ab|D Ab
C0363184|T201|COMP|1305-2|LNC|D Ag|D Ag
C0363229|T201|COMP|1034-8|LNC|Fetal cell screen|Fetal cell screen
C0363230|T201|COMP|1035-5|LNC|Fresh frozen plasma given|Fresh frozen plasma given
C0363243|T201|COMP|1051-2|LNC|Hemolytic disease of newborn screen|Hemolytic disease of newborn screen
C0363341|T201|COMP|1154-4|LNC|little c Ab|little c Ab
C0363342|T201|COMP|1155-1|LNC|little c Ab|little c Ab
C0363343|T201|COMP|1156-9|LNC|little c Ab|little c Ab
C0363344|T201|COMP|1157-7|LNC|little c Ag|little c Ag
C0363345|T201|COMP|1158-5|LNC|little c Ag|little c Ag
C0363346|T201|COMP|1159-3|LNC|little c Ag|little c Ag
C0363413|T201|COMP|1250-0|LNC|Major crossmatch|Major crossmatch
C0363414|T201|COMP|1251-8|LNC|Major crossmatch|Major crossmatch
C0363415|T201|COMP|1252-6|LNC|Major crossmatch^post immediate spin|Major crossmatch^post immediate spin
C0363416|T201|COMP|1253-4|LNC|Major crossmatch|Major crossmatch
C0363417|T201|COMP|1254-2|LNC|Major crossmatch.re-crossmatch|Major crossmatch.re-crossmatch
C0363418|T201|COMP|1255-9|LNC|Minor crossmatch|Minor crossmatch
C0363449|T201|COMP|1298-9|LNC|Packed erythrocytes given|Packed erythrocytes given
C0363450|T201|COMP|1299-7|LNC|Platelets given|Platelets given
C0363454|T201|COMP|1303-7|LNC|Reverse ABO group|Reverse ABO group
C0363457|T201|COMP|1321-9|LNC|Transfusion duration|Transfusion duration
C0363458|T201|COMP|1322-7|LNC|Transfusion volume|Transfusion volume
C0363471|T201|COMP|1335-9|LNC|Whole blood given|Whole blood given
C0363492|T201|COMP|1356-5|LNC|11-Deoxycortisol^8H post 30 mg/kg metyraPONE PO|11-Deoxycortisol^8H post 30 mg/kg metyraPONE PO
C0363493|T201|COMP|1357-3|LNC|11-Deoxycortisol^post 750 mg metyraPONE Q4H X 6|11-Deoxycortisol^post 750 mg metyraPONE Q4H X 6
C0363494|T201|COMP|1358-1|LNC|Corticotropin^1.5H post dose insulin IV|Corticotropin^1.5H post dose insulin IV
C0363496|T201|COMP|1360-7|LNC|Corticotropin^1H post dose insulin IV|Corticotropin^1H post dose insulin IV
C0363499|T201|COMP|1363-1|LNC|Corticotropin^30M post dose insulin IV|Corticotropin^30M post dose insulin IV
C0363501|T201|COMP|1365-6|LNC|Corticotropin^45M post dose insulin IV|Corticotropin^45M post dose insulin IV
C0363505|T201|COMP|1369-8|LNC|Ascorbate^post dose PO|Ascorbate^post dose PO
C0363507|T201|COMP|1371-4|LNC|Bromsulphthalein|Bromsulphthalein
C0363509|T201|COMP|1373-0|LNC|Calcitonin^10M post 2.4 mg/kg calcium short IV|Calcitonin^10M post 2.4 mg/kg calcium short IV
C0363510|T201|COMP|1374-8|LNC|Calcitonin^3H post 15 mg/kg calcium gluconate IV|Calcitonin^3H post 15 mg/kg calcium gluconate IV
C0363511|T201|COMP|1375-5|LNC|Calcitonin^4H post 15 mg/kg calcium gluconate IV|Calcitonin^4H post 15 mg/kg calcium gluconate IV
C0363513|T201|COMP|1377-1|LNC|Calcitonin^5M post 2.4 mg/kg calcium short IV|Calcitonin^5M post 2.4 mg/kg calcium short IV
C0363516|T201|COMP|1380-5|LNC|Calcium/Phosphate parathyroid-challenge test|Calcium/Phosphate parathyroid-challenge test
C0363517|T201|COMP|1381-3|LNC|Calcium^10M post 2.4 mg/kg calcium short IV|Calcium^10M post 2.4 mg/kg calcium short IV
C0363518|T201|COMP|1382-1|LNC|Calcium^5M post 2.4 mg/kg calcium short IV|Calcium^5M post 2.4 mg/kg calcium short IV
C0363520|T201|COMP|1384-7|LNC|Calcium^post calcium infusion|Calcium^post calcium infusion
C0363534|T201|COMP|1398-7|LNC|Cortisol^1.5H post dose insulin IV|Cortisol^1.5H post dose insulin IV
C0363540|T201|COMP|1404-3|LNC|Cortisol^1H post dose insulin IV|Cortisol^1H post dose insulin IV
C0363554|T201|COMP|1419-1|LNC|Cortisol^30M post dose insulin IV|Cortisol^30M post dose insulin IV
C0363558|T201|COMP|1424-1|LNC|Cortisol^45M post dose insulin IV|Cortisol^45M post dose insulin IV
C0363568|T201|COMP|1434-0|LNC|Cortisol^8H post 1 mg dexamethasone PO overnight|Cortisol^8H post 1 mg dexamethasone PO overnight
C0363570|T201|COMP|1436-5|LNC|Cortisol^8H post 30 mg/kg metyraPONE PO|Cortisol^8H post 30 mg/kg metyraPONE PO
C0363574|T201|COMP|1440-7|LNC|Cortisol^9H post 1 mg dexamethasone PO overnight|Cortisol^9H post 1 mg dexamethasone PO overnight
C0363575|T201|COMP|1441-5|LNC|Cortisol^9H post 3 g metyraPONE PO overnight|Cortisol^9H post 3 g metyraPONE PO overnight
C0363594|T201|COMP|1460-5|LNC|Cobalamins^post dose cyanocobalamin|Cobalamins^post dose cyanocobalamin
C0363599|T201|COMP|1465-4|LNC|EPINEPHrine^supine|EPINEPHrine^supine
C0363600|T201|COMP|1466-2|LNC|Follitropin^1.5H post 100 g lutropin IV|Follitropin^1.5H post 100 g lutropin IV
C0363611|T201|COMP|1477-9|LNC|Follitropin^baseline|Follitropin^baseline
C0363613|T201|COMP|1479-5|LNC|Galactose^1.5H post 40 g galactose PO|Galactose^1.5H post 40 g galactose PO
C0363614|T201|COMP|1480-3|LNC|Galactose^1H post 40 g galactose PO|Galactose^1H post 40 g galactose PO
C0363615|T201|COMP|1481-1|LNC|Galactose^2H post 40 g galactose PO|Galactose^2H post 40 g galactose PO
C0363616|T201|COMP|1482-9|LNC|Galactose^30M post 40 g galactose PO|Galactose^30M post 40 g galactose PO
C0363617|T201|COMP|1483-7|LNC|Galactose^post 40 g dose PO|Galactose^post 40 g dose PO
C0363618|T201|COMP|1484-5|LNC|Gastrin^10M post 0.2 U/kg secretin|Gastrin^10M post 0.2 U/kg secretin
C0363619|T201|COMP|1485-2|LNC|Gastrin^15M post 0.2 U/kg secretin|Gastrin^15M post 0.2 U/kg secretin
C0363620|T201|COMP|1486-0|LNC|Gastrin^20M post 0.2 U/kg secretin|Gastrin^20M post 0.2 U/kg secretin
C0363621|T201|COMP|1487-8|LNC|Gastrin^25M post 0.2 U/kg secretin|Gastrin^25M post 0.2 U/kg secretin
C0363622|T201|COMP|1488-6|LNC|Gastrin^30M post 0.2 U/kg secretin|Gastrin^30M post 0.2 U/kg secretin
C0363623|T201|COMP|1489-4|LNC|Gastrin^5M post 0.2 U/kg secretin|Gastrin^5M post 0.2 U/kg secretin
C0363625|T201|COMP|1491-0|LNC|Glucose^30M post 100 g glucose PO|Glucose^30M post 100 g glucose PO
C0363626|T201|COMP|1492-8|LNC|Glucose^1.5H post 0.5 g/kg glucose IV|Glucose^1.5H post 0.5 g/kg glucose IV
C0363628|T201|COMP|1494-4|LNC|Glucose^1.5H post 100 g glucose PO|Glucose^1.5H post 100 g glucose PO
C0363629|T201|COMP|1495-1|LNC|Glucose^1.5H post 100 g glucose PO|Glucose^1.5H post 100 g glucose PO
C0363631|T201|COMP|1497-7|LNC|Glucose^1.5H post dose insulin IV|Glucose^1.5H post dose insulin IV
C0363632|T201|COMP|1498-5|LNC|Glucose^10M post 0.5 g/kg glucose IV|Glucose^10M post 0.5 g/kg glucose IV
C0363633|T201|COMP|1499-3|LNC|Glucose^1H post 0.5 g/kg glucose IV|Glucose^1H post 0.5 g/kg glucose IV
C0363635|T201|COMP|1501-6|LNC|Glucose^1H post 100 g glucose PO|Glucose^1H post 100 g glucose PO
C0363636|T201|COMP|1502-4|LNC|Glucose^1H post 100 g glucose PO|Glucose^1H post 100 g glucose PO
C0363637|T201|COMP|1503-2|LNC|Glucose^1H post 100 g glucose PO|Glucose^1H post 100 g glucose PO
C0363638|T201|COMP|1504-0|LNC|Glucose^1H post 50 g glucose PO|Glucose^1H post 50 g glucose PO
C0363639|T201|COMP|1505-7|LNC|Glucose^1H post 50 g glucose PO|Glucose^1H post 50 g glucose PO
C0363640|T201|COMP|1506-5|LNC|Glucose^1H post 50 g lactose PO|Glucose^1H post 50 g lactose PO
C0363641|T201|COMP|1507-3|LNC|Glucose^1H post 75 g glucose PO|Glucose^1H post 75 g glucose PO
C0363642|T201|COMP|1508-1|LNC|Glucose^1H post 75 g glucose PO|Glucose^1H post 75 g glucose PO
C0363643|T201|COMP|1509-9|LNC|Glucose^1H post 75 g glucose PO|Glucose^1H post 75 g glucose PO
C0363644|T201|COMP|1510-7|LNC|Glucose^1H post dose insulin IV|Glucose^1H post dose insulin IV
C0363645|T201|COMP|1512-3|LNC|Glucose^1M post 0.5 g/kg glucose IV|Glucose^1M post 0.5 g/kg glucose IV
C0363646|T201|COMP|1513-1|LNC|Glucose^20M post 0.5 g/kg glucose IV|Glucose^20M post 0.5 g/kg glucose IV
C0363647|T201|COMP|1514-9|LNC|Glucose^2H post 100 g glucose PO|Glucose^2H post 100 g glucose PO
C0363648|T201|COMP|1515-6|LNC|Glucose^2H post 100 g glucose PO|Glucose^2H post 100 g glucose PO
C0363649|T201|COMP|1516-4|LNC|Glucose^2H post 100 g glucose PO|Glucose^2H post 100 g glucose PO
C0363650|T201|COMP|1517-2|LNC|Glucose^2H post 50 g lactose PO|Glucose^2H post 50 g lactose PO
C0363651|T201|COMP|1518-0|LNC|Glucose^2H post 75 g glucose PO|Glucose^2H post 75 g glucose PO
C0363652|T201|COMP|1519-8|LNC|Glucose^2H post 75 g glucose PO|Glucose^2H post 75 g glucose PO
C0363653|T201|COMP|1520-6|LNC|Glucose^2H post 75 g glucose PO|Glucose^2H post 75 g glucose PO
C0363655|T201|COMP|1522-2|LNC|Glucose^30M post 0.5 g/kg glucose IV|Glucose^30M post 0.5 g/kg glucose IV
C0363658|T201|COMP|1525-5|LNC|Glucose^30M post 100 g glucose PO|Glucose^30M post 100 g glucose PO
C0363659|T201|COMP|1526-3|LNC|Glucose^30M post 50 g lactose PO|Glucose^30M post 50 g lactose PO
C0363661|T201|COMP|1528-9|LNC|Glucose^30M post dose insulin IV|Glucose^30M post dose insulin IV
C0363662|T201|COMP|1530-5|LNC|Glucose^3H post 100 g glucose PO|Glucose^3H post 100 g glucose PO
C0363663|T201|COMP|1531-3|LNC|Glucose^3H post 100 g glucose PO|Glucose^3H post 100 g glucose PO
C0363664|T201|COMP|1532-1|LNC|Glucose^3H post 100 g glucose PO|Glucose^3H post 100 g glucose PO
C0363665|T201|COMP|1533-9|LNC|Glucose^3H post 75 g glucose PO|Glucose^3H post 75 g glucose PO
C0363666|T201|COMP|1534-7|LNC|Glucose^3M post 0.5 g/kg glucose IV|Glucose^3M post 0.5 g/kg glucose IV
C0363667|T201|COMP|1535-4|LNC|Glucose^40M post 0.5 g/kg glucose IV|Glucose^40M post 0.5 g/kg glucose IV
C0363668|T201|COMP|1536-2|LNC|Glucose^45M post dose insulin IV|Glucose^45M post dose insulin IV
C0363669|T201|COMP|1537-0|LNC|Glucose^4H post 100 g glucose PO|Glucose^4H post 100 g glucose PO
C0363670|T201|COMP|1538-8|LNC|Glucose^4H post 100 g glucose PO|Glucose^4H post 100 g glucose PO
C0363671|T201|COMP|1539-6|LNC|Glucose^4H post 75 g glucose PO|Glucose^4H post 75 g glucose PO
C0363672|T201|COMP|1540-4|LNC|Glucose^5H post 100 g glucose PO|Glucose^5H post 100 g glucose PO
C0363673|T201|COMP|1541-2|LNC|Glucose^5H post 100 g glucose PO|Glucose^5H post 100 g glucose PO
C0363674|T201|COMP|1542-0|LNC|Glucose^5H post 75 g glucose PO|Glucose^5H post 75 g glucose PO
C0363675|T201|COMP|1543-8|LNC|Glucose^5M post 0.5 g/kg glucose IV|Glucose^5M post 0.5 g/kg glucose IV
C0363676|T201|COMP|1545-3|LNC|Glucose^6H post 100 g glucose PO|Glucose^6H post 100 g glucose PO
C0363677|T201|COMP|1546-1|LNC|Glucose^6H post 100 g glucose PO|Glucose^6H post 100 g glucose PO
C0363678|T201|COMP|1547-9|LNC|Glucose^baseline|Glucose^baseline
C0363685|T201|COMP|1554-5|LNC|Glucose^post 12H CFst|Glucose^post 12H CFst
C0363686|T201|COMP|1555-2|LNC|Glucose^post 12H CFst|Glucose^post 12H CFst
C0363687|T201|COMP|1556-0|LNC|Glucose^post CFst|Glucose^post CFst
C0363688|T201|COMP|1557-8|LNC|Glucose^post CFst|Glucose^post CFst
C0363693|T201|COMP|1561-0|LNC|Insulin^1H post 75 g glucose PO|Insulin^1H post 75 g glucose PO
C0363696|T201|COMP|1564-4|LNC|Insulin^2H post 75 g glucose PO|Insulin^2H post 75 g glucose PO
C0363699|T201|COMP|1567-7|LNC|Insulin^3H post 75 g glucose PO|Insulin^3H post 75 g glucose PO
C0363700|T201|COMP|1568-5|LNC|Insulin^4H post 75 g glucose PO|Insulin^4H post 75 g glucose PO
C0363701|T201|COMP|1569-3|LNC|Insulin^5H post 75 g glucose PO|Insulin^5H post 75 g glucose PO
C0363702|T201|COMP|1570-1|LNC|Insulin^baseline|Insulin^baseline
C0363705|T201|COMP|1573-5|LNC|Insulin^post 12H CFst|Insulin^post 12H CFst
C0363714|T201|COMP|1582-6|LNC|Lactose^1H post 50 g lactose PO|Lactose^1H post 50 g lactose PO
C0363715|T201|COMP|1583-4|LNC|Lactose^2H post 50 g lactose PO|Lactose^2H post 50 g lactose PO
C0363716|T201|COMP|1584-2|LNC|Lactose^30M post 50 g lactose PO|Lactose^30M post 50 g lactose PO
C0363718|T201|COMP|1586-7|LNC|Lead^post EDTA therapy|Lead^post EDTA therapy
C0363719|T201|COMP|1587-5|LNC|Lutropin^1.5H post 100 g lutropin IV|Lutropin^1.5H post 100 g lutropin IV
C0363721|T201|COMP|1589-1|LNC|Lutropin^105M post 100 g lutropin IV|Lutropin^105M post 100 g lutropin IV
C0363722|T201|COMP|1590-9|LNC|Lutropin^15M post 100 g lutropin IV|Lutropin^15M post 100 g lutropin IV
C0363723|T201|COMP|1591-7|LNC|Lutropin^1H post 100 g lutropin IV|Lutropin^1H post 100 g lutropin IV
C0363725|T201|COMP|1593-3|LNC|Lutropin^2H post 100 g lutropin IV|Lutropin^2H post 100 g lutropin IV
C0363727|T201|COMP|1595-8|LNC|Lutropin^30M post 100 g lutropin IV|Lutropin^30M post 100 g lutropin IV
C0363729|T201|COMP|1597-4|LNC|Lutropin^45M post 100 g lutropin IV|Lutropin^45M post 100 g lutropin IV
C0363730|T201|COMP|1598-2|LNC|Lutropin^75M post 100 g lutropin IV|Lutropin^75M post 100 g lutropin IV
C0363731|T201|COMP|1599-0|LNC|Lutropin^baseline|Lutropin^baseline
C0363733|T201|COMP|1601-4|LNC|Norepinephrine^supine|Norepinephrine^supine
C0363734|T201|COMP|1602-2|LNC|Norepinephrine^10M post standing|Norepinephrine^10M post standing
C0363739|T201|COMP|1607-1|LNC|Osmolality^post 12H FFst|Osmolality^post 12H FFst
C0363740|T201|COMP|1608-9|LNC|Osmolality^post 8H FFst|Osmolality^post 8H FFst
C0363753|T201|COMP|1622-0|LNC|Renin^5H post 600 ug furosemide PO|Renin^5H post 600 ug furosemide PO
C0363755|T201|COMP|1624-6|LNC|Retinol^3H post 5000 units|Retinol^3H post 5000 units
C0363756|T201|COMP|1625-3|LNC|Retinol^6H post 5000 units|Retinol^6H post 5000 units
C0363757|T201|COMP|1626-1|LNC|Retinol^pre 5000 units|Retinol^pre 5000 units
C0363758|T201|COMP|1627-9|LNC|Somatotropin^1.5H post dose insulin IV|Somatotropin^1.5H post dose insulin IV
C0363759|T201|COMP|1628-7|LNC|Somatotropin^1H post 1 g/kg glucose PO|Somatotropin^1H post 1 g/kg glucose PO
C0363760|T201|COMP|1629-5|LNC|Somatotropin^1H post dose insulin IV|Somatotropin^1H post dose insulin IV
C0363761|T201|COMP|1630-3|LNC|Somatotropin^2H post 1 g/kg glucose PO|Somatotropin^2H post 1 g/kg glucose PO
C0363762|T201|COMP|1631-1|LNC|Somatotropin^30M post dose insulin IV|Somatotropin^30M post dose insulin IV
C0363763|T201|COMP|1632-9|LNC|Somatotropin^3H post 1 g/kg glucose PO|Somatotropin^3H post 1 g/kg glucose PO
C0363764|T201|COMP|1633-7|LNC|Somatotropin^45M post dose insulin IV|Somatotropin^45M post dose insulin IV
C0363769|T201|COMP|1638-6|LNC|Testosterone^96H post 5000 U HCG IM|Testosterone^96H post 5000 U HCG IM
C0363773|T201|COMP|1642-8|LNC|Thyrotropin^baseline|Thyrotropin^baseline
C0363775|T201|COMP|1644-4|LNC|Triglyceride^post 12H CFst|Triglyceride^post 12H CFst
C0363776|T201|COMP|1645-1|LNC|Xylose^2H post 25 g xylose PO|Xylose^2H post 25 g xylose PO
C0363777|T201|COMP|1646-9|LNC|Xylose^post dose PO|Xylose^post dose PO
C0363778|T201|COMP|1647-7|LNC|Tuberculosis reaction wheal^3D post 25 TU ID|Tuberculosis reaction wheal^3D post 25 TU ID
C0363779|T201|COMP|1648-5|LNC|Tuberculosis reaction wheal^3D post 5 TU ID|Tuberculosis reaction wheal^3D post 5 TU ID
C0363780|T201|COMP|5930-3|LNC|Mumps reaction wheal^3D post 0.1 mL mumps ID|Mumps reaction wheal^3D post 0.1 mL mumps ID
C0363783|T201|COMP|1649-3|LNC|Calcitriol|Calcitriol
C0363784|T201|COMP|1650-1|LNC|1,4-Alpha glucan branching enzyme|1,4-Alpha glucan branching enzyme
C0363785|T201|COMP|1651-9|LNC|1-Methylhistidine|1-Methylhistidine
C0363786|T201|COMP|1652-7|LNC|1-Methylhistidine|1-Methylhistidine
C0363787|T201|COMP|1653-5|LNC|1-Methylhistidine|1-Methylhistidine
C0363788|T201|COMP|1654-3|LNC|1-Naphthalene|1-Naphthalene
C0363789|T201|COMP|1655-0|LNC|11-Deoxy/11-Oxy steroids|11-Deoxy/11-Oxy steroids
C0363790|T201|COMP|1656-8|LNC|11-Deoxycorticosterone|11-Deoxycorticosterone
C0363791|T201|COMP|1657-6|LNC|11-Deoxycortisol|11-Deoxycortisol
C0363792|T201|COMP|1658-4|LNC|11-Hydroxyandrostenedione|11-Hydroxyandrostenedione
C0363793|T201|COMP|1659-2|LNC|11-Hydroxyandrosterone|11-Hydroxyandrosterone
C0363794|T201|COMP|1660-0|LNC|11-Hydroxyetiocholanolone|11-Hydroxyetiocholanolone
C0363795|T201|COMP|1661-8|LNC|11-Ketoandrosterone|11-Ketoandrosterone
C0363796|T201|COMP|1662-6|LNC|11-Ketoetiocholanolone|11-Ketoetiocholanolone
C0363797|T201|COMP|1663-4|LNC|11-Oxycorticosterone|11-Oxycorticosterone
C0363798|T201|COMP|1664-2|LNC|17-Hydroxycorticosteroids|17-Hydroxycorticosteroids
C0363799|T201|COMP|1665-9|LNC|17-Hydroxycorticosteroids|17-Hydroxycorticosteroids
C0363800|T201|COMP|1666-7|LNC|17-Hydroxycorticosteroids|17-Hydroxycorticosteroids
C0363801|T201|COMP|1667-5|LNC|17-Hydroxyketosteroids|17-Hydroxyketosteroids
C0363802|T201|COMP|1668-3|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C0363803|T201|COMP|1669-1|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C0363804|T201|COMP|1670-9|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C0363806|T201|COMP|1671-7|LNC|17-Ketogenic steroids|17-Ketogenic steroids
C0363807|T201|COMP|1673-3|LNC|17-Ketogenic steroids|17-Ketogenic steroids
C0363808|T201|COMP|1674-1|LNC|18-Hydroxycorticosterone|18-Hydroxycorticosterone
C0363809|T201|COMP|1675-8|LNC|2,3-Diphosphoglycerate|2,3-Diphosphoglycerate
C0363810|T201|COMP|1676-6|LNC|2,3-Diphosphoglycerate|2,3-Diphosphoglycerate
C0363811|T201|COMP|1677-4|LNC|Alpha hydroxybutyrate dehydrogenase|Alpha hydroxybutyrate dehydrogenase
C0363812|T201|COMP|1678-2|LNC|20-Hydroxyprogesterone|20-Hydroxyprogesterone
C0363813|T201|COMP|1679-0|LNC|24r-Hydroxycalcidiol|24r-Hydroxycalcidiol
C0363814|T201|COMP|1680-8|LNC|3-Alpha-Androstanediol glucuronide|3-Alpha-Androstanediol glucuronide
C0363815|T201|COMP|1681-6|LNC|Beta hydroxybutyrate dehydrogenase|Beta hydroxybutyrate dehydrogenase
C0363817|T201|COMP|1683-2|LNC|3-Hydroxyisovalerate|3-Hydroxyisovalerate
C0363818|T201|COMP|1684-0|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C0363819|T201|COMP|1685-7|LNC|3-Methylhistidine|3-Methylhistidine
C0363820|T201|COMP|1686-5|LNC|3-Methylhistidine|3-Methylhistidine
C0363821|T201|COMP|1687-3|LNC|3-Methylhistidine|3-Methylhistidine
C0363822|T201|COMP|1688-1|LNC|4-Pyridoxate|4-Pyridoxate
C0363823|T201|COMP|1689-9|LNC|5'-Nucleotidase|5'-Nucleotidase
C0363824|T201|COMP|1690-7|LNC|5'-Nucleotidase|5'-Nucleotidase
C0363825|T201|COMP|1691-5|LNC|5,10-Methylenetetrahydrofolate reductase|5,10-Methylenetetrahydrofolate reductase
C0363826|T201|COMP|1692-3|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C0363827|T201|COMP|1693-1|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C0363828|T201|COMP|1694-9|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C0363829|T201|COMP|1695-6|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C0363831|T201|COMP|1697-2|LNC|6-Phosphogluconate dehydrogenase|6-Phosphogluconate dehydrogenase
C0363832|T201|COMP|1698-0|LNC|8-Hydroxyamoxapine|8-Hydroxyamoxapine
C0363833|T201|COMP|1699-8|LNC|Alpha-L-iduronidase|Alpha-L-iduronidase
C0363834|T201|COMP|1700-4|LNC|Acetaldehyde|Acetaldehyde
C0363835|T201|COMP|1701-2|LNC|Acetaldehyde|Acetaldehyde
C0363836|T201|COMP|1702-0|LNC|Acetoacetate|Acetoacetate
C0363837|T201|COMP|1703-8|LNC|Acetoacetate|Acetoacetate
C0363838|T201|COMP|1704-6|LNC|Acetoacetate|Acetoacetate
C0363839|T201|COMP|1705-3|LNC|Acetoacetate|Acetoacetate
C0363840|T201|COMP|1706-1|LNC|Acetonitrile|Acetonitrile
C0363841|T201|COMP|1707-9|LNC|Acetylcholine|Acetylcholine
C0363842|T201|COMP|1708-7|LNC|Acetylcholinesterase|Acetylcholinesterase
C0363843|T201|COMP|1709-5|LNC|Acetylcholinesterase|Acetylcholinesterase
C0363844|T201|COMP|1710-3|LNC|Acetylcholinesterase|Acetylcholinesterase
C0363845|T201|COMP|1711-1|LNC|Acid phosphatase|Acid phosphatase
C0363846|T201|COMP|1712-9|LNC|Acid phosphatase.prostatic|Acid phosphatase.prostatic
C0363847|T201|COMP|1713-7|LNC|Acid phosphatase.prostatic|Acid phosphatase.prostatic
C0363848|T201|COMP|1714-5|LNC|Acid phosphatase.prostatic|Acid phosphatase.prostatic
C0363849|T201|COMP|1715-2|LNC|Acid phosphatase|Acid phosphatase
C0363850|T201|COMP|1716-0|LNC|Acidity.titratable|Acidity.titratable
C0363851|T201|COMP|1717-8|LNC|Acylcarnitine|Acylcarnitine
C0363852|T201|COMP|1718-6|LNC|Acyl CoA dehydrogenase|Acyl CoA dehydrogenase
C0363853|T201|COMP|1719-4|LNC|Adenine|Adenine
C0363854|T201|COMP|1720-2|LNC|Adenine phosphoribosyltransferase|Adenine phosphoribosyltransferase
C0363856|T201|COMP|1722-8|LNC|Adenosine deaminase|Adenosine deaminase
C0363857|T201|COMP|1723-6|LNC|Adenosine deaminase binding protein|Adenosine deaminase binding protein
C0363858|T201|COMP|1724-4|LNC|Adenosine diphosphate|Adenosine diphosphate
C0363859|T201|COMP|1725-1|LNC|Adenosine monophosphate deaminase|Adenosine monophosphate deaminase
C0363860|T201|COMP|1726-9|LNC|Adenosine monophosphate.cyclic|Adenosine monophosphate.cyclic
C0363861|T201|COMP|1727-7|LNC|Adenosine monophosphate.cyclic|Adenosine monophosphate.cyclic
C0363862|T201|COMP|1728-5|LNC|Adenosine monophosphate.cyclic/Creatinine|Adenosine monophosphate.cyclic/Creatinine
C0363863|T201|COMP|1729-3|LNC|Adenosine triphosphatase|Adenosine triphosphatase
C0363864|T201|COMP|1730-1|LNC|Adenosine triphosphatase|Adenosine triphosphatase
C0363865|T201|COMP|1731-9|LNC|Adenylate kinase|Adenylate kinase
C0363866|T201|COMP|1732-7|LNC|Adenylosuccinate lyase|Adenylosuccinate lyase
C0363867|T201|COMP|1733-5|LNC|Adipate|Adipate
C0363869|T201|COMP|1735-0|LNC|Alanine|Alanine
C0363870|T201|COMP|1736-8|LNC|Alanine|Alanine
C0363871|T201|COMP|1737-6|LNC|Alanine|Alanine
C0363872|T201|COMP|1738-4|LNC|Alanine|Alanine
C0363873|T201|COMP|1739-2|LNC|Alanine|Alanine
C0363874|T201|COMP|1740-0|LNC|Alanine aminopeptidase|Alanine aminopeptidase
C0363875|T201|COMP|1741-8|LNC|Alanine aminotransferase|Alanine aminotransferase
C0363876|T201|COMP|1742-6|LNC|Alanine aminotransferase|Alanine aminotransferase
C0363877|T201|COMP|1743-4|LNC|Alanine aminotransferase|Alanine aminotransferase
C0363878|T201|COMP|1744-2|LNC|Alanine aminotransferase|Alanine aminotransferase
C0363879|T201|COMP|1745-9|LNC|Albumin|Albumin
C0363880|T201|COMP|1746-7|LNC|Albumin|Albumin
C0363881|T201|COMP|1747-5|LNC|Albumin|Albumin
C0363882|T201|COMP|1748-3|LNC|Albumin|Albumin
C0363883|T201|COMP|1749-1|LNC|Albumin|Albumin
C0363884|T201|COMP|1750-9|LNC|Albumin|Albumin
C0363885|T201|COMP|1751-7|LNC|Albumin|Albumin
C0363886|T201|COMP|1752-5|LNC|Albumin|Albumin
C0363887|T201|COMP|1753-3|LNC|Albumin|Albumin
C0363888|T201|COMP|1754-1|LNC|Albumin|Albumin
C0363889|T201|COMP|1755-8|LNC|Albumin|Albumin
C0363890|T201|COMP|1756-6|LNC|Albumin.CSF/Albumin.SerPl|Albumin.CSF/Albumin.SerPl
C0363891|T201|COMP|1757-4|LNC|Albumin renal clearance|Albumin renal clearance
C0363892|T201|COMP|1758-2|LNC|Albumin.glycated|Albumin.glycated
C0363893|T201|COMP|1759-0|LNC|Albumin/Globulin|Albumin/Globulin
C0363894|T201|COMP|1760-8|LNC|Alcohol dehydrogenase|Alcohol dehydrogenase
C0363895|T201|COMP|1761-6|LNC|Aldolase|Aldolase
C0363896|T201|COMP|1762-4|LNC|Aldosterone|Aldosterone
C0363897|T201|COMP|1763-2|LNC|Aldosterone|Aldosterone
C0363898|T201|COMP|1764-0|LNC|Aldosterone|Aldosterone
C0363899|T201|COMP|1765-7|LNC|Aldosterone|Aldosterone
C0363900|T201|COMP|1766-5|LNC|Aldosterone receptors|Aldosterone receptors
C0363901|T201|COMP|1767-3|LNC|Aldosterone^supine|Aldosterone^supine
C0363902|T201|COMP|1768-1|LNC|Aldosterone^upright|Aldosterone^upright
C0363904|T201|COMP|1770-7|LNC|Aliphatic carboxylate C14-C26.absorption|Aliphatic carboxylate C14-C26.absorption
C0363905|T201|COMP|1771-5|LNC|Aliphatic carboxylate C14-C26.esters|Aliphatic carboxylate C14-C26.esters
C0363906|T201|COMP|1772-3|LNC|Aliphatic carboxylate C14-C26.esters|Aliphatic carboxylate C14-C26.esters
C0363907|T201|COMP|1773-1|LNC|Fatty acids.very long chain.C24:0/C22:0|Fatty acids.very long chain.C24:0/C22:0
C0363908|T201|COMP|1774-9|LNC|Fatty acids.very long chain.C26:0/C22:0|Fatty acids.very long chain.C26:0/C22:0
C0363909|T201|COMP|1775-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363910|T201|COMP|1776-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363911|T201|COMP|1777-2|LNC|Alkaline phosphatase.bone|Alkaline phosphatase.bone
C0363912|T201|COMP|1778-0|LNC|Alkaline phosphatase.intestinal|Alkaline phosphatase.intestinal
C0363913|T201|COMP|1779-8|LNC|Alkaline phosphatase.liver|Alkaline phosphatase.liver
C0363914|T201|COMP|1780-6|LNC|Alkaline phosphatase.placental|Alkaline phosphatase.placental
C0363915|T201|COMP|1781-4|LNC|Alkaline phosphatase.regan|Alkaline phosphatase.regan
C0363916|T201|COMP|1782-2|LNC|Alkaline phosphatase.renal|Alkaline phosphatase.renal
C0363917|T201|COMP|1783-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363918|T201|COMP|1784-8|LNC|Alpha amino acid nitrogen|Alpha amino acid nitrogen
C0363919|T201|COMP|1785-5|LNC|Alpha amino acid nitrogen|Alpha amino acid nitrogen
C0363920|T201|COMP|1786-3|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0363921|T201|COMP|1787-1|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0363922|T201|COMP|1788-9|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0363923|T201|COMP|1789-7|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0363924|T201|COMP|1790-5|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0363925|T201|COMP|1791-3|LNC|Alpha aminoadipate|Alpha aminoadipate
C0363926|T201|COMP|1792-1|LNC|Alpha aminoadipate|Alpha aminoadipate
C0363927|T201|COMP|1793-9|LNC|Alpha aminoadipate|Alpha aminoadipate
C0363928|T201|COMP|1794-7|LNC|Amylase|Amylase
C0363929|T201|COMP|1795-4|LNC|Amylase|Amylase
C0363930|T201|COMP|1796-2|LNC|Amylase|Amylase
C0363931|T201|COMP|1797-0|LNC|Amylase|Amylase
C0363933|T201|COMP|1799-6|LNC|Amylase|Amylase
C0363934|T201|COMP|1800-2|LNC|Amylase|Amylase
C0363935|T201|COMP|1801-0|LNC|Amylase renal clearance|Amylase renal clearance
C0363936|T201|COMP|1802-8|LNC|Amylase.P1|Amylase.P1
C0363937|T201|COMP|1803-6|LNC|Amylase.P2|Amylase.P2
C0363938|T201|COMP|1804-4|LNC|Amylase.P3|Amylase.P3
C0363939|T201|COMP|1805-1|LNC|Amylase.pancreatic|Amylase.pancreatic
C0363940|T201|COMP|1806-9|LNC|Amylase.S1|Amylase.S1
C0363941|T201|COMP|1807-7|LNC|Amylase.S2|Amylase.S2
C0363942|T201|COMP|1808-5|LNC|Amylase.S3|Amylase.S3
C0363943|T201|COMP|1809-3|LNC|Amylase.salivary|Amylase.salivary
C0363944|T201|COMP|1810-1|LNC|Amylase/Creatinine|Amylase/Creatinine
C0363945|T201|COMP|1811-9|LNC|Amylase/Creatinine renal clearance|Amylase/Creatinine renal clearance
C0363946|T201|COMP|1812-7|LNC|Alpha fucosidase|Alpha fucosidase
C0363947|T201|COMP|1813-5|LNC|Alpha galactosidase A|Alpha galactosidase A
C0363948|T201|COMP|1814-3|LNC|Acid alpha glucosidase|Acid alpha glucosidase
C0363949|T201|COMP|1815-0|LNC|Acid alpha glucosidase|Acid alpha glucosidase
C0363950|T201|COMP|1816-8|LNC|Acid alpha glucosidase|Acid alpha glucosidase
C0363951|T201|COMP|1818-4|LNC|Alpha mannosidase|Alpha mannosidase
C0363952|T201|COMP|1819-2|LNC|Alpha mannosidase|Alpha mannosidase
C0363953|T201|COMP|1820-0|LNC|Alpha melanocyte stimulating hormone|Alpha melanocyte stimulating hormone
C0363954|T201|COMP|1821-8|LNC|Alpha naphthylesterase|Alpha naphthylesterase
C0363955|T201|COMP|1822-6|LNC|Alpha thymosin|Alpha thymosin
C0363956|T201|COMP|1823-4|LNC|Alpha tocopherol|Alpha tocopherol
C0363957|T201|COMP|2684-9|LNC|Alpha-1-Acid glycoprotein|Alpha-1-Acid glycoprotein
C0363958|T201|COMP|2685-6|LNC|Alpha-1-Acid glycoprotein|Alpha-1-Acid glycoprotein
C0363959|T201|COMP|1824-2|LNC|Alpha-1-Antichymotrypsin|Alpha-1-Antichymotrypsin
C0363960|T201|COMP|1826-7|LNC|Alpha 1 antitrypsin.MM|Alpha 1 antitrypsin.MM
C0363961|T201|COMP|1827-5|LNC|Alpha 1 antitrypsin.MS|Alpha 1 antitrypsin.MS
C0363962|T201|COMP|1828-3|LNC|Alpha 1 antitrypsin.MZ|Alpha 1 antitrypsin.MZ
C0363963|T201|COMP|1829-1|LNC|Alpha 1 antitrypsin.SS|Alpha 1 antitrypsin.SS
C0363964|T201|COMP|1830-9|LNC|Alpha 1 antitrypsin.SZ|Alpha 1 antitrypsin.SZ
C0363965|T201|COMP|1831-7|LNC|Alpha 1 antitrypsin.ZZ|Alpha 1 antitrypsin.ZZ
C0363966|T201|COMP|1832-5|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0363967|T201|COMP|1833-3|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0363968|T201|COMP|1834-1|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0363970|T201|COMP|1835-8|LNC|Alpha-2-Macroglobulin|Alpha-2-Macroglobulin
C0363971|T201|COMP|1836-6|LNC|Alpha-2-Retinol binding protein|Alpha-2-Retinol binding protein
C0363973|T201|COMP|1838-2|LNC|Alpha-N-acetylglucosaminidase|Alpha-N-acetylglucosaminidase
C0363974|T201|COMP|1839-0|LNC|Ammonia|Ammonia
C0363975|T201|COMP|1840-8|LNC|Ammonia|Ammonia
C0363976|T201|COMP|1841-6|LNC|Ammonia|Ammonia
C0363977|T201|COMP|1842-4|LNC|Ammonia|Ammonia
C0363978|T201|COMP|1843-2|LNC|Ammonia nitrogen|Ammonia nitrogen
C0363979|T201|COMP|1844-0|LNC|Ammonium ion|Ammonium ion
C0363980|T201|COMP|1845-7|LNC|Ammonium ion|Ammonium ion
C0363981|T201|COMP|1846-5|LNC|Amylo-alpha-1,6-glucosidase|Amylo-alpha-1,6-glucosidase
C0363982|T201|COMP|1847-3|LNC|Amyloid associated protein|Amyloid associated protein
C0363983|T201|COMP|1848-1|LNC|Androstanolone|Androstanolone
C0363984|T201|COMP|1849-9|LNC|Androstanolone|Androstanolone
C0363985|T201|COMP|1850-7|LNC|Androstanediol|Androstanediol
C0363986|T201|COMP|1851-5|LNC|Androstenedione|Androstenedione
C0363987|T201|COMP|1852-3|LNC|Androstenedione|Androstenedione
C0363988|T201|COMP|1853-1|LNC|Androstenedione|Androstenedione
C0363989|T201|COMP|1854-9|LNC|Androstenedione|Androstenedione
C0363990|T201|COMP|1855-6|LNC|Androstenedione|Androstenedione
C0363991|T201|COMP|1856-4|LNC|Androsterone|Androsterone
C0363992|T201|COMP|1857-2|LNC|Angiotensin converting enzyme|Angiotensin converting enzyme
C0363993|T201|COMP|1858-0|LNC|Angiotensin I|Angiotensin I
C0363994|T201|COMP|1859-8|LNC|Angiotensin II|Angiotensin II
C0363995|T201|COMP|1860-6|LNC|Angiotensin II|Angiotensin II
C0363996|T201|COMP|1861-4|LNC|Angiotensinogen|Angiotensinogen
C0363997|T201|COMP|1862-2|LNC|Aniline|Aniline
C0363998|T201|COMP|1863-0|LNC|Anion gap 4|Anion gap 4
C0363999|T201|COMP|1864-8|LNC|Anserine|Anserine
C0364000|T201|COMP|1865-5|LNC|Anserine|Anserine
C0364001|T201|COMP|1866-3|LNC|Anserine|Anserine
C0364002|T201|COMP|1867-1|LNC|Anserine|Anserine
C0364003|T201|COMP|1868-9|LNC|Antithrombin Ag|Antithrombin Ag
C0364005|T201|COMP|1870-5|LNC|Apolipoprotein A-II|Apolipoprotein A-II
C0364006|T201|COMP|1871-3|LNC|Apolipoprotein B-100|Apolipoprotein B-100
C0364007|T201|COMP|1872-1|LNC|Apolipoprotein B-150|Apolipoprotein B-150
C0364008|T201|COMP|1873-9|LNC|Apolipoprotein B-48|Apolipoprotein B-48
C0364010|T201|COMP|1875-4|LNC|Apolipoprotein C-I|Apolipoprotein C-I
C0364011|T201|COMP|1876-2|LNC|Apolipoprotein C-II|Apolipoprotein C-II
C0364012|T201|COMP|1877-0|LNC|Apolipoprotein C-III|Apolipoprotein C-III
C0364013|T201|COMP|1878-8|LNC|Apolipoprotein A-III|Apolipoprotein A-III
C0364014|T201|COMP|1879-6|LNC|Apolipoprotein E2|Apolipoprotein E2
C0364015|T201|COMP|1880-4|LNC|Beta 2 glycoprotein 1|Beta 2 glycoprotein 1
C0364016|T201|COMP|1881-2|LNC|Apolipoprotein LPA|Apolipoprotein LPA
C0364017|T201|COMP|1882-0|LNC|Apolipoprotein LPQ|Apolipoprotein LPQ
C0364018|T201|COMP|1883-8|LNC|Apolipoprotein A|Apolipoprotein A
C0364019|T201|COMP|1884-6|LNC|Apolipoprotein B|Apolipoprotein B
C0364020|T201|COMP|1885-3|LNC|Apolipoprotein C|Apolipoprotein C
C0364021|T201|COMP|1886-1|LNC|Apolipoprotein E|Apolipoprotein E
C0364022|T201|COMP|1887-9|LNC|Appearance|Appearance
C0364023|T201|COMP|1888-7|LNC|Aquacobalamin|Aquacobalamin
C0364024|T201|COMP|1889-5|LNC|Arachidonate|Arachidonate
C0364025|T201|COMP|1890-3|LNC|Arginase|Arginase
C0364026|T201|COMP|1891-1|LNC|Arginine|Arginine
C0364027|T201|COMP|1892-9|LNC|Arginine|Arginine
C0364028|T201|COMP|1893-7|LNC|Arginine|Arginine
C0364029|T201|COMP|1894-5|LNC|Arginine|Arginine
C0364030|T201|COMP|1895-2|LNC|Arginine|Arginine
C0364031|T201|COMP|1896-0|LNC|Argininosuccinate|Argininosuccinate
C0364032|T201|COMP|1897-8|LNC|Argininosuccinate|Argininosuccinate
C0364033|T201|COMP|1898-6|LNC|Argininosuccinate lyase|Argininosuccinate lyase
C0364034|T201|COMP|1899-4|LNC|Argininosuccinate synthase|Argininosuccinate synthase
C0364035|T201|COMP|1900-0|LNC|Arylamidase|Arylamidase
C0364036|T201|COMP|1901-8|LNC|Arylsulfatase|Arylsulfatase
C0364037|T201|COMP|1902-6|LNC|Ascorbate|Ascorbate
C0364039|T201|COMP|1904-2|LNC|Ascorbate|Ascorbate
C0364040|T201|COMP|1905-9|LNC|Ascorbate|Ascorbate
C0364041|T201|COMP|1906-7|LNC|Asparagine|Asparagine
C0364042|T201|COMP|1907-5|LNC|Asparagine|Asparagine
C0364043|T201|COMP|1908-3|LNC|Asparagine|Asparagine
C0364044|T201|COMP|1909-1|LNC|Asparagine|Asparagine
C0364045|T201|COMP|1910-9|LNC|Asparagine|Asparagine
C0364046|T201|COMP|1911-7|LNC|Aspartate|Aspartate
C0364047|T201|COMP|1912-5|LNC|Aspartate|Aspartate
C0364048|T201|COMP|1913-3|LNC|Aspartate|Aspartate
C0364049|T201|COMP|1914-1|LNC|Aspartate|Aspartate
C0364050|T201|COMP|1915-8|LNC|Aspartate|Aspartate
C0364052|T201|COMP|1917-4|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0364053|T201|COMP|1918-2|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0364054|T201|COMP|1919-0|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0364055|T201|COMP|1920-8|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0364056|T201|COMP|1921-6|LNC|Atrial natriuretic factor|Atrial natriuretic factor
C0364057|T201|COMP|1922-4|LNC|Base deficit|Base deficit
C0364058|T201|COMP|1923-2|LNC|Base deficit|Base deficit
C0364059|T201|COMP|1924-0|LNC|Base deficit|Base deficit
C0364060|T201|COMP|1925-7|LNC|Base excess|Base excess
C0364061|T201|COMP|1926-5|LNC|Base excess|Base excess
C0364062|T201|COMP|1927-3|LNC|Base excess|Base excess
C0364063|T201|COMP|1930-7|LNC|Benzoate|Benzoate
C0364064|T201|COMP|1931-5|LNC|Beta alanine|Beta alanine
C0364065|T201|COMP|1932-3|LNC|Beta alanine|Beta alanine
C0364066|T201|COMP|1933-1|LNC|Beta alanine|Beta alanine
C0364067|T201|COMP|1934-9|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0364068|T201|COMP|1935-6|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0364069|T201|COMP|1936-4|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0364070|T201|COMP|1937-2|LNC|Beta endorphin|Beta endorphin
C0364072|T201|COMP|1939-8|LNC|Beta fructofuranosidase|Beta fructofuranosidase
C0364073|T201|COMP|1940-6|LNC|Beta galactosidase|Beta galactosidase
C0364074|T201|COMP|1941-4|LNC|Beta galactosidase|Beta galactosidase
C0364075|T201|COMP|1942-2|LNC|Beta galactosidase|Beta galactosidase
C0364076|T201|COMP|1943-0|LNC|Glucosylceramidase|Glucosylceramidase
C0364077|T201|COMP|1944-8|LNC|Beta glucuronidase|Beta glucuronidase
C0364078|T201|COMP|1945-5|LNC|Beta glucuronidase|Beta glucuronidase
C0364079|T201|COMP|1946-3|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C0364080|T201|COMP|1947-1|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C0364081|T201|COMP|1682-4|LNC|Beta hydroxybutyrate dehydrogenase|Beta hydroxybutyrate dehydrogenase
C0364082|T201|COMP|1949-7|LNC|Beta lipotropin|Beta lipotropin
C0364083|T201|COMP|1950-5|LNC|Beta melanocyte stimulating hormone|Beta melanocyte stimulating hormone
C0364084|T201|COMP|1951-3|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C0364085|T201|COMP|1952-1|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C0364086|T201|COMP|1953-9|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C0364087|T201|COMP|1954-7|LNC|Beta-N-acetylhexosaminidase|Beta-N-acetylhexosaminidase
C0364088|T201|COMP|1955-4|LNC|Beta-N-acetylhexosaminidase|Beta-N-acetylhexosaminidase
C0364089|T201|COMP|1956-2|LNC|Beta-N-acetylhexosaminidase.A|Beta-N-acetylhexosaminidase.A
C0364090|T201|COMP|1957-0|LNC|Beta-N-acetylhexosaminidase.B|Beta-N-acetylhexosaminidase.B
C0364091|T201|COMP|1958-8|LNC|Beta-N-acetylhexosaminidase.I|Beta-N-acetylhexosaminidase.I
C0364092|T201|COMP|1959-6|LNC|Bicarbonate|Bicarbonate
C0364093|T201|COMP|1960-4|LNC|Bicarbonate|Bicarbonate
C0364094|T201|COMP|1961-2|LNC|Bicarbonate|Bicarbonate
C0364095|T201|COMP|1962-0|LNC|Bicarbonate|Bicarbonate
C0364096|T201|COMP|1963-8|LNC|Bicarbonate|Bicarbonate
C0364097|T201|COMP|1964-6|LNC|Bicarbonate|Bicarbonate
C0364098|T201|COMP|1965-3|LNC|Bile|Bile
C0364100|T201|COMP|1967-9|LNC|Bile acid|Bile acid
C0364101|T201|COMP|1968-7|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C0364102|T201|COMP|1969-5|LNC|Bilirubin renal clearance|Bilirubin renal clearance
C0364103|T201|COMP|1970-3|LNC|Bilirubin.albumin bound|Bilirubin.albumin bound
C0364104|T201|COMP|1971-1|LNC|Bilirubin.non-glucuronidated|Bilirubin.non-glucuronidated
C0364105|T201|COMP|1972-9|LNC|Bilirubin|Bilirubin
C0364106|T201|COMP|1973-7|LNC|Bilirubin|Bilirubin
C0364108|T201|COMP|1975-2|LNC|Bilirubin|Bilirubin
C0364109|T201|COMP|1976-0|LNC|Bilirubin|Bilirubin
C0364110|T201|COMP|1977-8|LNC|Bilirubin|Bilirubin
C0364111|T201|COMP|1978-6|LNC|Bilirubin|Bilirubin
C0364112|T201|COMP|1979-4|LNC|Biopterin|Biopterin
C0364113|T201|COMP|1980-2|LNC|Biotin|Biotin
C0364114|T201|COMP|1981-0|LNC|Biotinidase|Biotinidase
C0364115|T201|COMP|1982-8|LNC|Biotinidase|Biotinidase
C0364116|T201|COMP|1983-6|LNC|Bradykinin|Bradykinin
C0364117|T201|COMP|1984-4|LNC|Bromide|Bromide
C0364118|T201|COMP|1985-1|LNC|Bromide|Bromide
C0364119|T201|COMP|1986-9|LNC|C peptide|C peptide
C0364120|T201|COMP|1987-7|LNC|C peptide|C peptide
C0364121|T201|COMP|1988-5|LNC|C reactive protein|C reactive protein
C0364122|T201|COMP|1989-3|LNC|Calcidiol|Calcidiol
C0364123|T201|COMP|1990-1|LNC|Cholecalciferol|Cholecalciferol
C0364124|T201|COMP|1991-9|LNC|Calciferol binding proteins|Calciferol binding proteins
C0364125|T201|COMP|1992-7|LNC|Calcitonin|Calcitonin
C0364126|T201|COMP|1993-5|LNC|Calcium renal clearance|Calcium renal clearance
C0364127|T201|COMP|1994-3|LNC|Calcium.ionized|Calcium.ionized
C0364128|T201|COMP|1995-0|LNC|Calcium.ionized|Calcium.ionized
C0364129|T201|COMP|1996-8|LNC|Calcium|Calcium
C0364130|T201|COMP|1997-6|LNC|Calcium|Calcium
C0364131|T201|COMP|1998-4|LNC|Calcium|Calcium
C0364132|T201|COMP|1999-2|LNC|Calcium|Calcium
C0364133|T201|COMP|2000-8|LNC|Calcium|Calcium
C0364134|T201|COMP|2001-6|LNC|Calcium|Calcium
C0364135|T201|COMP|2002-4|LNC|Calcium|Calcium
C0364136|T201|COMP|2004-0|LNC|Calcium|Calcium
C0364137|T201|COMP|2003-2|LNC|Calcium|Calcium
C0364138|T201|COMP|2005-7|LNC|Calcium^post 12H CFst|Calcium^post 12H CFst
C0364139|T201|COMP|2006-5|LNC|Cancer Ag 125|Cancer Ag 125
C0364140|T201|COMP|2007-3|LNC|Cancer Ag 15-3|Cancer Ag 15-3
C0364141|T201|COMP|2008-1|LNC|Cancer Ag 19-5|Cancer Ag 19-5
C0364142|T201|COMP|2009-9|LNC|Cancer Ag 19-9|Cancer Ag 19-9
C0364143|T201|COMP|2011-5|LNC|Cancer Ag 242|Cancer Ag 242
C0364144|T201|COMP|2012-3|LNC|Cancer Ag 27-29|Cancer Ag 27-29
C0364145|T201|COMP|2013-1|LNC|Cancer Ag 50|Cancer Ag 50
C0364146|T201|COMP|2014-9|LNC|Cancer Ag 549|Cancer Ag 549
C0364147|T201|COMP|2015-6|LNC|Cancer Ag 72-4|Cancer Ag 72-4
C0364148|T201|COMP|2016-4|LNC|Carbamoyl phosphate synthetase|Carbamoyl phosphate synthetase
C0364149|T201|COMP|2017-2|LNC|Carbamoyl phosphate synthetase(ammonia)|Carbamoyl phosphate synthetase(ammonia)
C0364150|T201|COMP|2018-0|LNC|Carbon dioxide|Carbon dioxide
C0364151|T201|COMP|2019-8|LNC|Carbon dioxide|Carbon dioxide
C0364152|T201|COMP|2020-6|LNC|Carbon dioxide|Carbon dioxide
C0364153|T201|COMP|2021-4|LNC|Carbon dioxide|Carbon dioxide
C0364154|T201|COMP|2022-2|LNC|Carbon dioxide|Carbon dioxide
C0364155|T201|COMP|2023-0|LNC|Carbon dioxide|Carbon dioxide
C0364156|T201|COMP|2024-8|LNC|Carbon dioxide.dissolved|Carbon dioxide.dissolved
C0364157|T201|COMP|2025-5|LNC|Carbon dioxide.dissolved|Carbon dioxide.dissolved
C0364158|T201|COMP|2026-3|LNC|Carbon dioxide|Carbon dioxide
C0364159|T201|COMP|2027-1|LNC|Carbon dioxide|Carbon dioxide
C0364160|T201|COMP|2028-9|LNC|Carbon dioxide|Carbon dioxide
C0364162|T201|COMP|2030-5|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C0364163|T201|COMP|2031-3|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C0364164|T201|COMP|2032-1|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C0364165|T201|COMP|2033-9|LNC|Carbonate|Carbonate
C0364166|T201|COMP|2034-7|LNC|Carbonate|Carbonate
C0364167|T201|COMP|2035-4|LNC|Carbonate|Carbonate
C0364168|T201|COMP|2036-2|LNC|Carbonate dehydratase|Carbonate dehydratase
C0364169|T201|COMP|2037-0|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0364170|T201|COMP|2038-8|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0364171|T201|COMP|2039-6|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0364172|T201|COMP|2040-4|LNC|Cardiolipin|Cardiolipin
C0364173|T201|COMP|2041-2|LNC|Carnitine acyltransferase|Carnitine acyltransferase
C0364174|T201|COMP|2042-0|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C0364175|T201|COMP|2043-8|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C0364176|T201|COMP|2044-6|LNC|Carnitine|Carnitine
C0364177|T201|COMP|2045-3|LNC|Carnitine|Carnitine
C0364178|T201|COMP|2046-1|LNC|Carnitine|Carnitine
C0364179|T201|COMP|2047-9|LNC|Carnitine|Carnitine
C0364180|T201|COMP|2048-7|LNC|Carnitine/Creatinine|Carnitine/Creatinine
C0364181|T201|COMP|2049-5|LNC|Carnosine|Carnosine
C0364182|T201|COMP|2050-3|LNC|Carnosine|Carnosine
C0364183|T201|COMP|2051-1|LNC|Carnosine|Carnosine
C0364184|T201|COMP|2052-9|LNC|Carotene|Carotene
C0364185|T201|COMP|2053-7|LNC|Carotene|Carotene
C0364186|T201|COMP|2054-5|LNC|Catalase|Catalase
C0364187|T201|COMP|2055-2|LNC|Catecholamines|Catecholamines
C0364188|T201|COMP|2056-0|LNC|Catecholamines|Catecholamines
C0364189|T201|COMP|2057-8|LNC|Catecholamines|Catecholamines
C0364190|T201|COMP|2058-6|LNC|Catecholamines|Catecholamines
C0364191|T201|COMP|2059-4|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C0364192|T201|COMP|2060-2|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C0364193|T201|COMP|2061-0|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C0364194|T201|COMP|2062-8|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C0364195|T201|COMP|2063-6|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C0364196|T201|COMP|2064-4|LNC|Ceruloplasmin|Ceruloplasmin
C0364197|T201|COMP|2065-1|LNC|Chenodeoxycholate|Chenodeoxycholate
C0364198|T201|COMP|2066-9|LNC|Chenodeoxycholylglycine|Chenodeoxycholylglycine
C0364199|T201|COMP|2067-7|LNC|Chenodeoxycholylglycine.conjugated|Chenodeoxycholylglycine.conjugated
C0364200|T201|COMP|2068-5|LNC|Chloride|Chloride
C0364201|T201|COMP|2069-3|LNC|Chloride|Chloride
C0364202|T201|COMP|2070-1|LNC|Chloride|Chloride
C0364203|T201|COMP|2071-9|LNC|Chloride|Chloride
C0364204|T201|COMP|2072-7|LNC|Chloride|Chloride
C0364205|T201|COMP|2073-5|LNC|Chloride|Chloride
C0364206|T201|COMP|2074-3|LNC|Chloride|Chloride
C0364207|T201|COMP|2075-0|LNC|Chloride|Chloride
C0364208|T201|COMP|2076-8|LNC|Chloride|Chloride
C0364209|T201|COMP|2077-6|LNC|Chloride|Chloride
C0364210|T201|COMP|2078-4|LNC|Chloride|Chloride
C0364211|T201|COMP|2079-2|LNC|Chloride|Chloride
C0364212|T201|COMP|2080-0|LNC|Cholate|Cholate
C0364213|T201|COMP|2081-8|LNC|Cholecystokinin|Cholecystokinin
C0364214|T201|COMP|2082-6|LNC|Cholestanol|Cholestanol
C0364215|T201|COMP|5932-9|LNC|Cholesterol|Cholesterol
C0364216|T201|COMP|2083-4|LNC|Cholesterol esterase|Cholesterol esterase
C0364217|T201|COMP|2084-2|LNC|Cholesterol esters|Cholesterol esters
C0364218|T201|COMP|2094-1|LNC|Cholesterol.non-esterified|Cholesterol.non-esterified
C0364219|T201|COMP|2096-6|LNC|Cholesterol/Triglyceride|Cholesterol/Triglyceride
C0364221|T201|COMP|2085-9|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C0364223|T201|COMP|2087-5|LNC|Cholesterol.in IDL|Cholesterol.in IDL
C0364225|T201|COMP|2089-1|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C0364227|T201|COMP|2091-7|LNC|Cholesterol.in VLDL|Cholesterol.in VLDL
C0364229|T201|COMP|2097-4|LNC|Cholinesterase|Cholinesterase
C0364230|T201|COMP|2098-2|LNC|Cholinesterase|Cholinesterase
C0364231|T201|COMP|2099-0|LNC|Cholinesterase|Cholinesterase
C0364232|T201|COMP|2100-6|LNC|Cholylglycine|Cholylglycine
C0364233|T201|COMP|2101-4|LNC|Cholylglycine.conjugated|Cholylglycine.conjugated
C0364234|T201|COMP|2102-2|LNC|Chondroitin sulfate|Chondroitin sulfate
C0364235|T201|COMP|2105-5|LNC|Choriogonadotropin|Choriogonadotropin
C0364236|T201|COMP|2106-3|LNC|Choriogonadotropin (pregnancy test)|Choriogonadotropin (pregnancy test)
C0364237|T201|COMP|2107-1|LNC|Choriogonadotropin|Choriogonadotropin
C0364238|T201|COMP|2118-8|LNC|Choriogonadotropin (pregnancy test)|Choriogonadotropin (pregnancy test)
C0364239|T201|COMP|2119-6|LNC|Choriogonadotropin|Choriogonadotropin
C0364240|T201|COMP|2103-0|LNC|Choriomammotropin|Choriomammotropin
C0364241|T201|COMP|2104-8|LNC|Choriomammotropin|Choriomammotropin
C0364242|T201|COMP|2108-9|LNC|Choriogonadotropin.alpha subunit|Choriogonadotropin.alpha subunit
C0364243|T201|COMP|2109-7|LNC|Choriogonadotropin.alpha subunit|Choriogonadotropin.alpha subunit
C0364244|T201|COMP|2110-5|LNC|Choriogonadotropin.beta subunit (pregnancy test)|Choriogonadotropin.beta subunit (pregnancy test)
C0364245|T201|COMP|2111-3|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0364246|T201|COMP|2112-1|LNC|Choriogonadotropin.beta subunit (pregnancy test)|Choriogonadotropin.beta subunit (pregnancy test)
C0364247|T201|COMP|2113-9|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0364248|T201|COMP|2114-7|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0364249|T201|COMP|2115-4|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C0364250|T201|COMP|2116-2|LNC|Choriogonadotropin.intact|Choriogonadotropin.intact
C0364251|T201|COMP|2117-0|LNC|Choriogonadotropin.intact|Choriogonadotropin.intact
C0364252|T201|COMP|2120-4|LNC|Chylomicrons|Chylomicrons
C0364253|T201|COMP|2121-2|LNC|Chylomicrons|Chylomicrons
C0364254|T201|COMP|2122-0|LNC|Chymopapain|Chymopapain
C0364255|T201|COMP|2123-8|LNC|Chymotrypsin|Chymotrypsin
C0364256|T201|COMP|2124-6|LNC|Chymotrypsin|Chymotrypsin
C0364257|T201|COMP|2125-3|LNC|Chymotrypsin|Chymotrypsin
C0364258|T201|COMP|2126-1|LNC|Citrate|Citrate
C0364259|T201|COMP|2127-9|LNC|Citrate|Citrate
C0364260|T201|COMP|2128-7|LNC|Citrate|Citrate
C0364261|T201|COMP|2129-5|LNC|Citrulline|Citrulline
C0364262|T201|COMP|2130-3|LNC|Citrulline|Citrulline
C0364263|T201|COMP|2131-1|LNC|Citrulline|Citrulline
C0364264|T201|COMP|2132-9|LNC|Cobalamins|Cobalamins
C0364265|T201|COMP|2133-7|LNC|Collagenase|Collagenase
C0364266|T201|COMP|2134-5|LNC|Coproporphyrin|Coproporphyrin
C0364267|T201|COMP|2135-2|LNC|Coproporphyrin|Coproporphyrin
C0364268|T201|COMP|2136-0|LNC|Coproporphyrin|Coproporphyrin
C0364269|T201|COMP|2137-8|LNC|Coproporphyrin|Coproporphyrin
C0364270|T201|COMP|2138-6|LNC|Coproporphyrinogen oxidase|Coproporphyrinogen oxidase
C0364271|T201|COMP|2139-4|LNC|Corticosterone|Corticosterone
C0364272|T201|COMP|2140-2|LNC|Corticotropin|Corticotropin
C0364273|T201|COMP|2141-0|LNC|Corticotropin|Corticotropin
C0364274|T201|COMP|2142-8|LNC|Cortisol|Cortisol
C0364275|T201|COMP|2143-6|LNC|Cortisol|Cortisol
C0364276|T201|COMP|2144-4|LNC|Cortisol|Cortisol
C0364278|T201|COMP|2145-1|LNC|Cortisol.free|Cortisol.free
C0364279|T201|COMP|2147-7|LNC|Cortisol.free|Cortisol.free
C0364280|T201|COMP|2148-5|LNC|Creatine|Creatine
C0364281|T201|COMP|2149-3|LNC|Creatine|Creatine
C0364282|T201|COMP|2150-1|LNC|Creatine|Creatine
C0364283|T201|COMP|2151-9|LNC|Creatine kinase|Creatine kinase
C0364284|T201|COMP|5912-1|LNC|Creatine kinase isoenzymes|Creatine kinase isoenzymes
C0364285|T201|COMP|2152-7|LNC|Creatine kinase.BB|Creatine kinase.BB
C0364286|T201|COMP|2153-5|LNC|Creatine kinase.macromolecular|Creatine kinase.macromolecular
C0364287|T201|COMP|2154-3|LNC|Creatine kinase.MB|Creatine kinase.MB
C0364288|T201|COMP|2155-0|LNC|Creatine kinase.MM|Creatine kinase.MM
C0364289|T201|COMP|2156-8|LNC|Creatine kinase|Creatine kinase
C0364290|T201|COMP|2157-6|LNC|Creatine kinase|Creatine kinase
C0364291|T201|COMP|2158-4|LNC|Creatine kinase.total/Creatine kinase.MB|Creatine kinase.total/Creatine kinase.MB
C0364292|T201|COMP|2159-2|LNC|Creatinine|Creatinine
C0364293|T201|COMP|5919-6|LNC|Creatinine|Creatinine
C0364294|T201|COMP|2160-0|LNC|Creatinine|Creatinine
C0364295|T201|COMP|2161-8|LNC|Creatinine|Creatinine
C0364296|T201|COMP|2162-6|LNC|Creatinine|Creatinine
C0364297|T201|COMP|2163-4|LNC|Creatinine renal clearance|Creatinine renal clearance
C0364298|T201|COMP|2164-2|LNC|Creatinine renal clearance|Creatinine renal clearance
C0364299|T201|COMP|2165-9|LNC|Cryofibrinogen|Cryofibrinogen
C0364300|T201|COMP|2166-7|LNC|Cryoglobulin|Cryoglobulin
C0364301|T201|COMP|2167-5|LNC|Cryoglobulin|Cryoglobulin
C0364302|T201|COMP|2168-3|LNC|Cryoglobulin|Cryoglobulin
C0364303|T201|COMP|2169-1|LNC|Cobalamins renal clearance|Cobalamins renal clearance
C0364304|T201|COMP|2170-9|LNC|Cyanocobalamin.true|Cyanocobalamin.true
C0364305|T201|COMP|2171-7|LNC|Cobalamins.unsaturated binding capacity|Cobalamins.unsaturated binding capacity
C0364306|T201|COMP|2172-5|LNC|Cystathionine|Cystathionine
C0364307|T201|COMP|2173-3|LNC|Cystathionine|Cystathionine
C0364308|T201|COMP|2174-1|LNC|Cystathionine|Cystathionine
C0364309|T201|COMP|2175-8|LNC|Cystine|Cystine
C0364310|T201|COMP|2176-6|LNC|Cystine|Cystine
C0364311|T201|COMP|2177-4|LNC|Cystine|Cystine
C0364312|T201|COMP|2178-2|LNC|Cystine|Cystine
C0364313|T201|COMP|2179-0|LNC|Cystine|Cystine
C0364314|T201|COMP|2180-8|LNC|Cystine+Cysteine|Cystine+Cysteine
C0364315|T201|COMP|2181-6|LNC|Cystinyl aminopeptidase|Cystinyl aminopeptidase
C0364316|T201|COMP|2182-4|LNC|Cytochrome B reductase|Cytochrome B reductase
C0364317|T201|COMP|2183-2|LNC|Cytochrome B5 reductase|Cytochrome B5 reductase
C0364318|T201|COMP|2184-0|LNC|Cytochrome C oxidase|Cytochrome C oxidase
C0364319|T201|COMP|2185-7|LNC|Cytochrome C oxidase|Cytochrome C oxidase
C0364320|T201|COMP|2186-5|LNC|Cytochrome C oxidase|Cytochrome C oxidase
C0364321|T201|COMP|2187-3|LNC|Cytosol aminopeptidase|Cytosol aminopeptidase
C0364322|T201|COMP|2188-1|LNC|Cytosol aminopeptidase|Cytosol aminopeptidase
C0364323|T201|COMP|2189-9|LNC|Cytosol aminopeptidase|Cytosol aminopeptidase
C0364324|T201|COMP|2190-7|LNC|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C0364325|T201|COMP|2191-5|LNC|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C0364326|T201|COMP|2192-3|LNC|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C0364327|T201|COMP|2193-1|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C0364328|T201|COMP|2194-9|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C0364329|T201|COMP|2195-6|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C0364330|T201|COMP|2196-4|LNC|Dehydroepiandrosterone.unconjugated|Dehydroepiandrosterone.unconjugated
C0364331|T201|COMP|2197-2|LNC|Dehydroepiandrosterone.unconjugated|Dehydroepiandrosterone.unconjugated
C0364332|T201|COMP|2198-0|LNC|Delta aminolevulinate|Delta aminolevulinate
C0364333|T201|COMP|2199-8|LNC|Delta aminolevulinate|Delta aminolevulinate
C0364334|T201|COMP|2200-4|LNC|Delta aminolevulinate|Delta aminolevulinate
C0364335|T201|COMP|2201-2|LNC|Deoxycholate|Deoxycholate
C0364336|T201|COMP|2202-0|LNC|Deoxycholylglycine|Deoxycholylglycine
C0364337|T201|COMP|2203-8|LNC|Dermatan sulfate|Dermatan sulfate
C0364338|T201|COMP|2204-6|LNC|Dermatan sulfate|Dermatan sulfate
C0364339|T201|COMP|2205-3|LNC|Diacetate|Diacetate
C0364340|T201|COMP|2206-1|LNC|Dicarboxylate C6-C8-C10|Dicarboxylate C6-C8-C10
C0364341|T201|COMP|2207-9|LNC|Dicarboxylate C6-C8-C10|Dicarboxylate C6-C8-C10
C0364342|T201|COMP|2208-7|LNC|Diethyl ether|Diethyl ether
C0364343|T201|COMP|2209-5|LNC|Dihydrofolate|Dihydrofolate
C0364344|T201|COMP|2210-3|LNC|Dihydrolipoamide acetyl transferase|Dihydrolipoamide acetyl transferase
C0364345|T201|COMP|2211-1|LNC|Dihydrolipoamide dehydrogenase|Dihydrolipoamide dehydrogenase
C0364346|T201|COMP|2212-9|LNC|Dihydropteridine reductase|Dihydropteridine reductase
C0364347|T201|COMP|2213-7|LNC|Dimethadione|Dimethadione
C0364348|T201|COMP|2214-5|LNC|Dinitrobenzene|Dinitrobenzene
C0364349|T201|COMP|2215-2|LNC|Dipalmitoylphosphatidylcholine|Dipalmitoylphosphatidylcholine
C0364350|T201|COMP|2216-0|LNC|DOPamine|DOPamine
C0364351|T201|COMP|2217-8|LNC|DOPamine|DOPamine
C0364352|T201|COMP|2218-6|LNC|DOPamine|DOPamine
C0364353|T201|COMP|2219-4|LNC|DOPamine beta-hydroxylase|DOPamine beta-hydroxylase
C0364354|T201|COMP|2556-9|LNC|Lecithin phosphorus|Lecithin phosphorus
C0364355|T201|COMP|2220-2|LNC|Elastase.pancreatic.free|Elastase.pancreatic.free
C0364356|T201|COMP|2221-0|LNC|Elastase.pancreatic|Elastase.pancreatic
C0364357|T201|COMP|2222-8|LNC|Elastase.pancreatic 2|Elastase.pancreatic 2
C0364358|T201|COMP|2223-6|LNC|Elastase.leukocyte|Elastase.leukocyte
C0364359|T201|COMP|2224-4|LNC|Enolase|Enolase
C0364360|T201|COMP|2225-1|LNC|Enolase.neuron specific|Enolase.neuron specific
C0364361|T201|COMP|2226-9|LNC|Enteroglucagon|Enteroglucagon
C0364362|T201|COMP|2227-7|LNC|Enteropeptidase|Enteropeptidase
C0364363|T201|COMP|2228-5|LNC|Enterotoxin|Enterotoxin
C0364364|T201|COMP|2229-3|LNC|Epiandrosterone|Epiandrosterone
C0364365|T201|COMP|2230-1|LNC|EPINEPHrine|EPINEPHrine
C0364366|T201|COMP|2231-9|LNC|EPINEPHrine|EPINEPHrine
C0364367|T201|COMP|2232-7|LNC|EPINEPHrine|EPINEPHrine
C0364368|T201|COMP|2233-5|LNC|Epitestosterone|Epitestosterone
C0364369|T201|COMP|2234-3|LNC|Epitestosterone|Epitestosterone
C0364370|T201|COMP|2235-0|LNC|Epitestosterone|Epitestosterone
C0364371|T201|COMP|2236-8|LNC|Calciferol|Calciferol
C0364372|T201|COMP|2237-6|LNC|Erythropoietin|Erythropoietin
C0364374|T201|COMP|2239-2|LNC|Estradiol|Estradiol
C0364375|T201|COMP|2240-0|LNC|Estradiol.free|Estradiol.free
C0364376|T201|COMP|2241-8|LNC|Estradiol.free|Estradiol.free
C0364377|T201|COMP|2242-6|LNC|Estradiol.free|Estradiol.free
C0364378|T201|COMP|2243-4|LNC|Estradiol|Estradiol
C0364379|T201|COMP|2238-4|LNC|Estradiol|Estradiol
C0364380|T201|COMP|2245-9|LNC|Estradiol|Estradiol
C0364381|T201|COMP|2246-7|LNC|Estradiol.unconjugated|Estradiol.unconjugated
C0364382|T201|COMP|2247-5|LNC|Estriol.conjugated|Estriol.conjugated
C0364383|T201|COMP|2248-3|LNC|Estriol|Estriol
C0364384|T201|COMP|2249-1|LNC|Estriol.unconjugated|Estriol.unconjugated
C0364385|T201|COMP|2250-9|LNC|Estriol.unconjugated|Estriol.unconjugated
C0364386|T201|COMP|2251-7|LNC|Estriol|Estriol
C0364387|T201|COMP|2252-5|LNC|Estriol|Estriol
C0364388|T201|COMP|2253-3|LNC|Estriol|Estriol
C0364389|T201|COMP|2254-1|LNC|Estrogen|Estrogen
C0364390|T201|COMP|2255-8|LNC|Estrogen|Estrogen
C0364391|T201|COMP|2256-6|LNC|Estrogen|Estrogen
C0364392|T201|COMP|2257-4|LNC|Estrone|Estrone
C0364393|T201|COMP|2258-2|LNC|Estrone|Estrone
C0364394|T201|COMP|2259-0|LNC|Estrone|Estrone
C0364395|T201|COMP|2260-8|LNC|Estrone.unconjugated|Estrone.unconjugated
C0364396|T201|COMP|2261-6|LNC|Estrone.unconjugated|Estrone.unconjugated
C0364397|T201|COMP|2262-4|LNC|Estrone.unconjugated|Estrone.unconjugated
C0364398|T201|COMP|2263-2|LNC|Ethanolamine|Ethanolamine
C0364399|T201|COMP|2264-0|LNC|Ethanolamine|Ethanolamine
C0364400|T201|COMP|2265-7|LNC|Ethylmalonate|Ethylmalonate
C0364401|T201|COMP|2266-5|LNC|Etiocholanolone|Etiocholanolone
C0364402|T201|COMP|2267-3|LNC|Etiocholanolone|Etiocholanolone
C0364403|T201|COMP|2268-1|LNC|Etiocholanolone|Etiocholanolone
C0364404|T201|COMP|2269-9|LNC|Complement factor B|Complement factor B
C0364408|T201|COMP|2273-1|LNC|Fatty acids.esterified|Fatty acids.esterified
C0364409|T201|COMP|2274-9|LNC|Fatty acids.nonesterified|Fatty acids.nonesterified
C0364410|T201|COMP|2275-6|LNC|Fatty acids|Fatty acids
C0364411|T201|COMP|2276-4|LNC|Ferritin|Ferritin
C0364412|T201|COMP|2277-2|LNC|Ferrochelatase|Ferrochelatase
C0364413|T201|COMP|2279-8|LNC|Fibrinopeptide A|Fibrinopeptide A
C0364414|T201|COMP|2278-0|LNC|Fibrinopeptide B|Fibrinopeptide B
C0364415|T201|COMP|2280-6|LNC|Fibronectin|Fibronectin
C0364416|T201|COMP|2281-4|LNC|Flavin adenine dinucleotide|Flavin adenine dinucleotide
C0364417|T201|COMP|2282-2|LNC|Folate|Folate
C0364418|T201|COMP|2283-0|LNC|Folate|Folate
C0364419|T201|COMP|2284-8|LNC|Folate|Folate
C0364420|T201|COMP|2285-5|LNC|Follitropin|Follitropin
C0364421|T201|COMP|2286-3|LNC|Follitropin|Follitropin
C0364422|T201|COMP|2287-1|LNC|Follitropin|Follitropin
C0364423|T201|COMP|2288-9|LNC|Follitropin.alpha subunit|Follitropin.alpha subunit
C0364424|T201|COMP|2289-7|LNC|Follitropin.beta subunit|Follitropin.beta subunit
C0364425|T201|COMP|2290-5|LNC|Follitropin/Lutropin|Follitropin/Lutropin
C0364426|T201|COMP|2291-3|LNC|Formate|Formate
C0364427|T201|COMP|2292-1|LNC|Formate|Formate
C0364428|T201|COMP|2293-9|LNC|Fructokinase|Fructokinase
C0364429|T201|COMP|2294-7|LNC|Fructosamine|Fructosamine
C0364430|T201|COMP|2295-4|LNC|Fructose|Fructose
C0364431|T201|COMP|2296-2|LNC|Fructose|Fructose
C0364432|T201|COMP|2297-0|LNC|Fructose|Fructose
C0364435|T201|COMP|2298-8|LNC|Aldolase|Aldolase
C0364435|T201|COMP|2300-2|LNC|Aldolase|Aldolase
C0364435|T201|COMP|6698-5|LNC|Aldolase|Aldolase
C0364436|T201|COMP|2301-0|LNC|Aldolase|Aldolase
C0364437|T201|COMP|2302-8|LNC|Fumarase|Fumarase
C0364438|T201|COMP|2303-6|LNC|Fumarate|Fumarate
C0364439|T201|COMP|2304-4|LNC|Fumarylacetoacetate|Fumarylacetoacetate
C0364440|T201|COMP|2305-1|LNC|Galactokinase|Galactokinase
C0364441|T201|COMP|2306-9|LNC|Galactose|Galactose
C0364442|T201|COMP|2307-7|LNC|Galactose|Galactose
C0364443|T201|COMP|2308-5|LNC|Galactose|Galactose
C0364444|T201|COMP|2309-3|LNC|Galactose|Galactose
C0364445|T201|COMP|2310-1|LNC|Galactose|Galactose
C0364446|T201|COMP|2311-9|LNC|Galactose renal clearance|Galactose renal clearance
C0364447|T201|COMP|2312-7|LNC|Galactose 1 phosphate|Galactose 1 phosphate
C0364448|T201|COMP|2314-3|LNC|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C0364449|T201|COMP|2313-5|LNC|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C0364450|T201|COMP|2315-0|LNC|Galactosylceramidase|Galactosylceramidase
C0364451|T201|COMP|2316-8|LNC|Galactosylgalactosylglucosylceramidase|Galactosylgalactosylglucosylceramidase
C0364452|T201|COMP|2317-6|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0364453|T201|COMP|2318-4|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0364454|T201|COMP|2319-2|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0364455|T201|COMP|2320-0|LNC|Gamma glutamyl cysteine synthetase|Gamma glutamyl cysteine synthetase
C0364456|T201|COMP|2321-8|LNC|Gamma glutamyl cysteine synthetase|Gamma glutamyl cysteine synthetase
C0364457|T201|COMP|2322-6|LNC|Gamma glutamyl transferase|Gamma glutamyl transferase
C0364458|T201|COMP|2323-4|LNC|Gamma glutamyl transferase|Gamma glutamyl transferase
C0364459|T201|COMP|2324-2|LNC|Gamma glutamyl transferase|Gamma glutamyl transferase
C0364461|T201|COMP|5925-3|LNC|Gastric acid|Gastric acid
C0364462|T201|COMP|5923-8|LNC|Gastric acid.free|Gastric acid.free
C0364463|T201|COMP|5922-0|LNC|Gastric acid|Gastric acid
C0364464|T201|COMP|2326-7|LNC|Gastric inhibitory polypeptide|Gastric inhibitory polypeptide
C0364465|T201|COMP|2327-5|LNC|Gastrin releasing polypeptide|Gastrin releasing polypeptide
C0364466|T201|COMP|2328-3|LNC|Gastrin releasing polypeptide|Gastrin releasing polypeptide
C0364467|T201|COMP|2329-1|LNC|Gastrin releasing polypeptide|Gastrin releasing polypeptide
C0364468|T201|COMP|2331-7|LNC|Gastrin.17 residue fragment|Gastrin.17 residue fragment
C0364469|T201|COMP|2330-9|LNC|Gastrin.34 residue fragment|Gastrin.34 residue fragment
C0364470|T201|COMP|2332-5|LNC|Gastrin.14 residue fragment|Gastrin.14 residue fragment
C0364471|T201|COMP|2333-3|LNC|Gastrin|Gastrin
C0364472|T201|COMP|2334-1|LNC|Hemoglobin.gastrointestinal|Hemoglobin.gastrointestinal
C0364473|T201|COMP|2335-8|LNC|Hemoglobin.gastrointestinal|Hemoglobin.gastrointestinal
C0364474|T201|COMP|2336-6|LNC|Globulin|Globulin
C0364475|T201|COMP|2337-4|LNC|Glucagon|Glucagon
C0364476|T201|COMP|2338-2|LNC|Glucagon|Glucagon
C0364477|T201|COMP|6300-8|LNC|Glucose|Glucose
C0364478|T201|COMP|5914-7|LNC|Glucose|Glucose
C0364479|T201|COMP|2339-0|LNC|Glucose|Glucose
C0364480|T201|COMP|2340-8|LNC|Glucose|Glucose
C0364481|T201|COMP|2341-6|LNC|Glucose|Glucose
C0364482|T201|COMP|2342-4|LNC|Glucose|Glucose
C0364483|T201|COMP|2343-2|LNC|Glucose|Glucose
C0364484|T201|COMP|2344-0|LNC|Glucose|Glucose
C0364486|T201|COMP|2346-5|LNC|Glucose|Glucose
C0364487|T201|COMP|2347-3|LNC|Glucose|Glucose
C0364488|T201|COMP|2348-1|LNC|Glucose|Glucose
C0364489|T201|COMP|2349-9|LNC|Glucose|Glucose
C0364490|T201|COMP|2350-7|LNC|Glucose|Glucose
C0364491|T201|COMP|2351-5|LNC|Glucose|Glucose
C0364492|T201|COMP|2352-3|LNC|Glucose CSF/Glucose plas|Glucose CSF/Glucose plas
C0364493|T201|COMP|2353-1|LNC|Glucose phosphate isomerase|Glucose phosphate isomerase
C0364494|T201|COMP|2354-9|LNC|Glucose-6-Phosphatase|Glucose-6-Phosphatase
C0364495|T201|COMP|2355-6|LNC|Glucose-6-Phosphatase|Glucose-6-Phosphatase
C0364496|T201|COMP|2356-4|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C0364497|T201|COMP|2357-2|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C0364498|T201|COMP|2358-0|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C0364499|T201|COMP|2359-8|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C0364500|T201|COMP|2360-6|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C0364501|T201|COMP|2361-4|LNC|Glucosylceramidase|Glucosylceramidase
C0364502|T201|COMP|2362-2|LNC|Glutamate|Glutamate
C0364503|T201|COMP|2363-0|LNC|Glutamate|Glutamate
C0364504|T201|COMP|2364-8|LNC|Glutamate|Glutamate
C0364505|T201|COMP|2365-5|LNC|Glutamate|Glutamate
C0364506|T201|COMP|2366-3|LNC|Glutamate|Glutamate
C0364507|T201|COMP|2367-1|LNC|Glutamate dehydrogenase|Glutamate dehydrogenase
C0364508|T201|COMP|2368-9|LNC|Glutamate dehydrogenase.NAD|Glutamate dehydrogenase.NAD
C0364509|T201|COMP|2369-7|LNC|Glutamate dehydrogenase.NADP|Glutamate dehydrogenase.NADP
C0364510|T201|COMP|2370-5|LNC|Glutamine|Glutamine
C0364511|T201|COMP|2371-3|LNC|Glutamine|Glutamine
C0364512|T201|COMP|2372-1|LNC|Glutamine|Glutamine
C0364513|T201|COMP|2373-9|LNC|Glutamine|Glutamine
C0364514|T201|COMP|2374-7|LNC|Glutamine|Glutamine
C0364515|T201|COMP|2375-4|LNC|Glutaryl CoA dehydrogenase|Glutaryl CoA dehydrogenase
C0364516|T201|COMP|2376-2|LNC|Glutathione peroxidase|Glutathione peroxidase
C0364517|T201|COMP|2377-0|LNC|Glutathione peroxidase|Glutathione peroxidase
C0364518|T201|COMP|2378-8|LNC|Glutathione reductase|Glutathione reductase
C0364519|T201|COMP|2379-6|LNC|Glutathione S-transferase|Glutathione S-transferase
C0364520|T201|COMP|2380-4|LNC|Glutathione synthase|Glutathione synthase
C0364521|T201|COMP|2381-2|LNC|Glutathione.oxidized|Glutathione.oxidized
C0364522|T201|COMP|2382-0|LNC|Glutathione.reduced|Glutathione.reduced
C0364523|T201|COMP|2383-8|LNC|Glutathione|Glutathione
C0364524|T201|COMP|2384-6|LNC|Glyceraldehyde 3 phosphate dehydrogenase|Glyceraldehyde 3 phosphate dehydrogenase
C0364525|T201|COMP|2385-3|LNC|Glycerate|Glycerate
C0364526|T201|COMP|2386-1|LNC|Glycerate|Glycerate
C0364527|T201|COMP|2388-7|LNC|Glycerol|Glycerol
C0364528|T201|COMP|2387-9|LNC|Glycerol|Glycerol
C0364529|T201|COMP|2389-5|LNC|Glycine|Glycine
C0364530|T201|COMP|2390-3|LNC|Glycine|Glycine
C0364531|T201|COMP|2391-1|LNC|Glycine|Glycine
C0364532|T201|COMP|2392-9|LNC|Glycine|Glycine
C0364533|T201|COMP|2393-7|LNC|Glycine|Glycine
C0364534|T201|COMP|2394-5|LNC|Glycogen synthase|Glycogen synthase
C0364535|T201|COMP|2395-2|LNC|Glycolate|Glycolate
C0364536|T201|COMP|2396-0|LNC|Glycolate|Glycolate
C0364537|T201|COMP|2397-8|LNC|Glycoproteins|Glycoproteins
C0364538|T201|COMP|2398-6|LNC|Glycosaminoglycans|Glycosaminoglycans
C0364539|T201|COMP|2399-4|LNC|Glycosaminoglycans|Glycosaminoglycans
C0364540|T201|COMP|2400-0|LNC|Guanine deaminase|Guanine deaminase
C0364541|T201|COMP|2401-8|LNC|Guanine deaminase|Guanine deaminase
C0364542|T201|COMP|2402-6|LNC|Guanosine monophosphate.cyclic|Guanosine monophosphate.cyclic
C0364543|T201|COMP|2095-8|LNC|Cholesterol.in HDL/Cholesterol.total|Cholesterol.in HDL/Cholesterol.total
C0364545|T201|COMP|2404-2|LNC|Hemopexin|Hemopexin
C0364546|T201|COMP|2405-9|LNC|Heparan sulfate|Heparan sulfate
C0364547|T201|COMP|2406-7|LNC|Heparan sulfate|Heparan sulfate
C0364548|T201|COMP|2407-5|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C0364549|T201|COMP|2408-3|LNC|Hexachlorophene|Hexachlorophene
C0364550|T201|COMP|2409-1|LNC|Hexokinase|Hexokinase
C0364551|T201|COMP|2410-9|LNC|Hexokinase|Hexokinase
C0364552|T201|COMP|2411-7|LNC|Hexokinase 1/Hexokinase.total|Hexokinase 1/Hexokinase.total
C0364553|T201|COMP|2412-5|LNC|Hexokinase 3/Hexokinase.total|Hexokinase 3/Hexokinase.total
C0364554|T201|COMP|2413-3|LNC|Hippuran renal clearance|Hippuran renal clearance
C0364555|T201|COMP|2414-1|LNC|Hippurate|Hippurate
C0364556|T201|COMP|2415-8|LNC|Histamine|Histamine
C0364557|T201|COMP|2416-6|LNC|Histamine|Histamine
C0364558|T201|COMP|2417-4|LNC|Histamine|Histamine
C0364559|T201|COMP|2418-2|LNC|Histidine|Histidine
C0364560|T201|COMP|2419-0|LNC|Histidine|Histidine
C0364561|T201|COMP|2420-8|LNC|Histidine|Histidine
C0364562|T201|COMP|2421-6|LNC|Histidine|Histidine
C0364563|T201|COMP|2422-4|LNC|Histidine|Histidine
C0364564|T201|COMP|2423-2|LNC|Histidine|Histidine
C0364565|T201|COMP|2424-0|LNC|Histidine|Histidine
C0364566|T201|COMP|2425-7|LNC|Histidine ammonia lyase|Histidine ammonia lyase
C0364567|T201|COMP|2426-5|LNC|Homocarnosine|Homocarnosine
C0364568|T201|COMP|2427-3|LNC|Homocitrulline|Homocitrulline
C0364569|T201|COMP|2428-1|LNC|Homocysteine|Homocysteine
C0364570|T201|COMP|2429-9|LNC|Homocystine|Homocystine
C0364571|T201|COMP|2430-7|LNC|Homocystine|Homocystine
C0364572|T201|COMP|2431-5|LNC|Homocystine|Homocystine
C0364573|T201|COMP|2432-3|LNC|Homogentisate|Homogentisate
C0364574|T201|COMP|2433-1|LNC|Homogentisate|Homogentisate
C0364575|T201|COMP|2434-9|LNC|Homovanillate|Homovanillate
C0364576|T201|COMP|2435-6|LNC|Homovanillate|Homovanillate
C0364577|T201|COMP|2436-4|LNC|Homovanillate|Homovanillate
C0364578|T201|COMP|2438-0|LNC|Hydrogen sulfide|Hydrogen sulfide
C0364579|T201|COMP|2439-8|LNC|Hydroxycalcidiol|Hydroxycalcidiol
C0364580|T201|COMP|2440-6|LNC|Hydroxocobalamin|Hydroxocobalamin
C0364581|T201|COMP|2441-4|LNC|Hydroxylysine|Hydroxylysine
C0364582|T201|COMP|2442-2|LNC|Hydroxylysine|Hydroxylysine
C0364583|T201|COMP|2443-0|LNC|Hydroxylysine|Hydroxylysine
C0364584|T201|COMP|2444-8|LNC|Hydroxymethylglutaryl CoA lyase|Hydroxymethylglutaryl CoA lyase
C0364585|T201|COMP|2445-5|LNC|Hydroxyproline|Hydroxyproline
C0364586|T201|COMP|2446-3|LNC|Hydroxyproline|Hydroxyproline
C0364588|T201|COMP|2448-9|LNC|Hydroxyproline.free|Hydroxyproline.free
C0364589|T201|COMP|2449-7|LNC|Hydroxyproline.free|Hydroxyproline.free
C0364590|T201|COMP|2450-5|LNC|Hydroxyproline.free|Hydroxyproline.free
C0364591|T201|COMP|2451-3|LNC|Hydroxyproline|Hydroxyproline
C0364592|T201|COMP|2452-1|LNC|Hypoxanthine|Hypoxanthine
C0364593|T201|COMP|2453-9|LNC|Hypoxanthine|Hypoxanthine
C0364594|T201|COMP|2454-7|LNC|Hypoxanthine phosphoribosyltransferase|Hypoxanthine phosphoribosyltransferase
C0364595|T201|COMP|2455-4|LNC|Hypoxanthine phosphoribosyltransferase|Hypoxanthine phosphoribosyltransferase
C0364596|T201|COMP|2456-2|LNC|Iduronate-2-Sulfatase|Iduronate-2-Sulfatase
C0364597|T201|COMP|2457-0|LNC|IgA|IgA
C0364598|T201|COMP|2458-8|LNC|IgA|IgA
C0364599|T201|COMP|2459-6|LNC|IgA.monoclonal|IgA.monoclonal
C0364600|T201|COMP|2460-4|LNC|IgD|IgD
C0364601|T201|COMP|2461-2|LNC|IgD.monoclonal|IgD.monoclonal
C0364602|T201|COMP|2462-0|LNC|IgE|IgE
C0364603|T201|COMP|2463-8|LNC|IgE.monoclonal|IgE.monoclonal
C0364604|T201|COMP|2464-6|LNC|IgG|IgG
C0364605|T201|COMP|2465-3|LNC|IgG|IgG
C0364606|T201|COMP|2466-1|LNC|IgG subclass 1|IgG subclass 1
C0364607|T201|COMP|2467-9|LNC|IgG subclass 2|IgG subclass 2
C0364608|T201|COMP|2468-7|LNC|IgG subclass 3|IgG subclass 3
C0364609|T201|COMP|2469-5|LNC|IgG subclass 4|IgG subclass 4
C0364610|T201|COMP|2470-3|LNC|IgG/Albumin|IgG/Albumin
C0364611|T201|COMP|2471-1|LNC|IgM|IgM
C0364612|T201|COMP|2472-9|LNC|IgM|IgM
C0364613|T201|COMP|2473-7|LNC|IgM.monoclonal|IgM.monoclonal
C0364614|T201|COMP|1928-1|LNC|Immunoglobulin light chains|Immunoglobulin light chains
C0364615|T201|COMP|1929-9|LNC|Immunoglobulin light chains|Immunoglobulin light chains
C0364616|T201|COMP|2474-5|LNC|Indicans|Indicans
C0364617|T201|COMP|2475-2|LNC|Indicans|Indicans
C0364618|T201|COMP|2476-0|LNC|Indolamine|Indolamine
C0364619|T201|COMP|2477-8|LNC|Indole|Indole
C0364620|T201|COMP|2478-6|LNC|Inhibin|Inhibin
C0364621|T201|COMP|2479-4|LNC|Inosine|Inosine
C0364622|T201|COMP|2480-2|LNC|Inositol.free|Inositol.free
C0364623|T201|COMP|2481-0|LNC|Insulin Ab|Insulin Ab
C0364624|T201|COMP|2482-8|LNC|Insulin Ab|Insulin Ab
C0364625|T201|COMP|2483-6|LNC|Insulin-like growth factor binding protein 3|Insulin-like growth factor binding protein 3
C0364626|T201|COMP|2484-4|LNC|Insulin-like growth factor-I|Insulin-like growth factor-I
C0364627|T201|COMP|2485-1|LNC|Insulin-like growth factor-II|Insulin-like growth factor-II
C0364628|T201|COMP|2487-7|LNC|Inter alpha trypsin inhibitor|Inter alpha trypsin inhibitor
C0364629|T201|COMP|2488-5|LNC|Intrinsic factor|Intrinsic factor
C0364630|T201|COMP|2489-3|LNC|Intrinsic factor blocking Ab|Intrinsic factor blocking Ab
C0364631|T201|COMP|2490-1|LNC|Inulin|Inulin
C0364632|T201|COMP|2491-9|LNC|Inulin renal clearance|Inulin renal clearance
C0364633|T201|COMP|2492-7|LNC|Iodine|Iodine
C0364634|T201|COMP|2493-5|LNC|Iodine.free|Iodine.free
C0364635|T201|COMP|2494-3|LNC|Iodine|Iodine
C0364636|T201|COMP|2495-0|LNC|Iodine|Iodine
C0364637|T201|COMP|2496-8|LNC|Iodohippuran renal clearance|Iodohippuran renal clearance
C0364638|T201|COMP|2497-6|LNC|Iron|Iron
C0364639|T201|COMP|2498-4|LNC|Iron|Iron
C0364640|T201|COMP|2499-2|LNC|Iron|Iron
C0364641|T201|COMP|2500-7|LNC|Iron binding capacity|Iron binding capacity
C0364642|T201|COMP|2501-5|LNC|Iron binding capacity.unsaturated|Iron binding capacity.unsaturated
C0364643|T201|COMP|2502-3|LNC|Iron saturation|Iron saturation
C0364644|T201|COMP|2503-1|LNC|Iron.chelated|Iron.chelated
C0364645|T201|COMP|2504-9|LNC|Iron|Iron
C0364646|T201|COMP|2505-6|LNC|Iron/Iron binding capacity.total|Iron/Iron binding capacity.total
C0364647|T201|COMP|2506-4|LNC|Isocitrate dehydrogenase|Isocitrate dehydrogenase
C0364648|T201|COMP|2507-2|LNC|Isoleucine|Isoleucine
C0364649|T201|COMP|2508-0|LNC|Isoleucine|Isoleucine
C0364650|T201|COMP|2509-8|LNC|Isoleucine|Isoleucine
C0364651|T201|COMP|2510-6|LNC|Isoleucine|Isoleucine
C0364652|T201|COMP|2511-4|LNC|Keratan sulfate|Keratan sulfate
C0364653|T201|COMP|2512-2|LNC|Keratan sulfate|Keratan sulfate
C0364654|T201|COMP|2513-0|LNC|Ketones|Ketones
C0364655|T201|COMP|2514-8|LNC|Ketones|Ketones
C0364656|T201|COMP|2515-5|LNC|Kynurenate|Kynurenate
C0364657|T201|COMP|2516-3|LNC|L-iditol dehydrogenase|L-iditol dehydrogenase
C0364658|T201|COMP|2517-1|LNC|L-iditol dehydrogenase|L-iditol dehydrogenase
C0364659|T201|COMP|2518-9|LNC|Lactate|Lactate
C0364660|T201|COMP|2519-7|LNC|Lactate|Lactate
C0364661|T201|COMP|2520-5|LNC|Lactate|Lactate
C0364662|T201|COMP|2521-3|LNC|Lactate|Lactate
C0364663|T201|COMP|2522-1|LNC|Lactate|Lactate
C0364664|T201|COMP|2523-9|LNC|Lactate|Lactate
C0364665|T201|COMP|2524-7|LNC|Lactate|Lactate
C0364666|T201|COMP|2525-4|LNC|Lactate|Lactate
C0364667|T201|COMP|2526-2|LNC|Lactate|Lactate
C0364668|T201|COMP|2527-0|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0364669|T201|COMP|2528-8|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0364670|T201|COMP|5921-2|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0364671|T201|COMP|2529-6|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0364672|T201|COMP|2530-4|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0364673|T201|COMP|2531-2|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0364674|T201|COMP|2532-0|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0364675|T201|COMP|2533-8|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0364676|T201|COMP|2534-6|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0364677|T201|COMP|5910-5|LNC|Lactate dehydrogenase isoenzymes|Lactate dehydrogenase isoenzymes
C0364678|T201|COMP|2535-3|LNC|Lactate dehydrogenase 1|Lactate dehydrogenase 1
C0364680|T201|COMP|2537-9|LNC|Lactate dehydrogenase 1|Lactate dehydrogenase 1
C0364681|T201|COMP|2538-7|LNC|Lactate dehydrogenase 2|Lactate dehydrogenase 2
C0364683|T201|COMP|2540-3|LNC|Lactate dehydrogenase 2|Lactate dehydrogenase 2
C0364684|T201|COMP|2541-1|LNC|Lactate dehydrogenase 3|Lactate dehydrogenase 3
C0364686|T201|COMP|2543-7|LNC|Lactate dehydrogenase 3|Lactate dehydrogenase 3
C0364687|T201|COMP|2544-5|LNC|Lactate dehydrogenase 4|Lactate dehydrogenase 4
C0364689|T201|COMP|2546-0|LNC|Lactate dehydrogenase 4|Lactate dehydrogenase 4
C0364690|T201|COMP|2547-8|LNC|Lactate dehydrogenase 5|Lactate dehydrogenase 5
C0364692|T201|COMP|2549-4|LNC|Lactate dehydrogenase 5|Lactate dehydrogenase 5
C0364693|T201|COMP|2550-2|LNC|Lactate/Pyruvate|Lactate/Pyruvate
C0364694|T201|COMP|2551-0|LNC|Lactoferrin|Lactoferrin
C0364695|T201|COMP|2552-8|LNC|Lactose|Lactose
C0364696|T201|COMP|2553-6|LNC|Lactose|Lactose
C0364697|T201|COMP|2554-4|LNC|Lactose|Lactose
C0364698|T201|COMP|5933-7|LNC|Lead|Lead
C0364699|T201|COMP|2555-1|LNC|Lecithin cholesterol acyltransferase|Lecithin cholesterol acyltransferase
C0364700|T201|COMP|2557-7|LNC|Lecithin/Sphingomyelin|Lecithin/Sphingomyelin
C0364701|T201|COMP|2558-5|LNC|Leucine|Leucine
C0364702|T201|COMP|2559-3|LNC|Leucine|Leucine
C0364703|T201|COMP|2560-1|LNC|Leucine|Leucine
C0364704|T201|COMP|2561-9|LNC|Leucine|Leucine
C0364705|T201|COMP|2562-7|LNC|Leucine|Leucine
C0364706|T201|COMP|2563-5|LNC|Leukocyte esterase|Leukocyte esterase
C0364707|T201|COMP|2564-3|LNC|Linoleate|Linoleate
C0364708|T201|COMP|2093-3|LNC|Cholesterol|Cholesterol
C0364709|T201|COMP|1769-9|LNC|Fatty acids.nonesterified|Fatty acids.nonesterified
C0364710|T201|COMP|2567-6|LNC|Phospholipid phosphorus|Phospholipid phosphorus
C0364712|T201|COMP|2569-2|LNC|Lipids|Lipids
C0364714|T201|COMP|2571-8|LNC|Triglyceride|Triglyceride
C0364715|T201|COMP|5911-3|LNC|Lipoprotein pattern|Lipoprotein pattern
C0364716|T201|COMP|2572-6|LNC|Lipoprotein lipase|Lipoprotein lipase
C0364717|T201|COMP|2573-4|LNC|Lipoprotein.alpha|Lipoprotein.alpha
C0364718|T201|COMP|2574-2|LNC|Lipoprotein.beta|Lipoprotein.beta
C0364719|T201|COMP|2575-9|LNC|Lipoprotein.pre-beta|Lipoprotein.pre-beta
C0364720|T201|COMP|2576-7|LNC|Lipoprotein|Lipoprotein
C0364721|T201|COMP|2577-5|LNC|Lithocholate|Lithocholate
C0364722|T201|COMP|2578-3|LNC|Lutropin|Lutropin
C0364723|T201|COMP|2579-1|LNC|Lutropin|Lutropin
C0364724|T201|COMP|2580-9|LNC|Lutropin|Lutropin
C0364725|T201|COMP|2581-7|LNC|Gonadotropin releasing hormone|Gonadotropin releasing hormone
C0364726|T201|COMP|2582-5|LNC|Lutropin.alpha subunit|Lutropin.alpha subunit
C0364727|T201|COMP|2583-3|LNC|Lutropin.beta subunit|Lutropin.beta subunit
C0364728|T201|COMP|2584-1|LNC|Lysine|Lysine
C0364729|T201|COMP|2585-8|LNC|Lysine|Lysine
C0364730|T201|COMP|2586-6|LNC|Lysine|Lysine
C0364731|T201|COMP|2587-4|LNC|Lysine|Lysine
C0364732|T201|COMP|2588-2|LNC|Lysolecithin acyltransferase|Lysolecithin acyltransferase
C0364733|T201|COMP|2589-0|LNC|Lysozyme|Lysozyme
C0364734|T201|COMP|2590-8|LNC|Lysozyme|Lysozyme
C0364735|T201|COMP|2591-6|LNC|Macroamylase|Macroamylase
C0364736|T201|COMP|2592-4|LNC|Macroglobulin|Macroglobulin
C0364737|T201|COMP|2593-2|LNC|Magnesium|Magnesium
C0364738|T201|COMP|2594-0|LNC|Magnesium|Magnesium
C0364739|T201|COMP|2595-7|LNC|Magnesium|Magnesium
C0364740|T201|COMP|2596-5|LNC|Magnesium|Magnesium
C0364741|T201|COMP|2597-3|LNC|Magnesium|Magnesium
C0364742|T201|COMP|2598-1|LNC|Magnesium|Magnesium
C0364743|T201|COMP|2599-9|LNC|Magnesium|Magnesium
C0364744|T201|COMP|2600-5|LNC|Magnesium.ionized|Magnesium.ionized
C0364745|T201|COMP|2601-3|LNC|Magnesium|Magnesium
C0364746|T201|COMP|2602-1|LNC|Malate dehydrogenase|Malate dehydrogenase
C0364747|T201|COMP|2603-9|LNC|Malonate|Malonate
C0364748|T201|COMP|2604-7|LNC|Mannitol renal clearance|Mannitol renal clearance
C0364749|T201|COMP|2605-4|LNC|Meat fibers|Meat fibers
C0364750|T201|COMP|2606-2|LNC|Melanin|Melanin
C0364751|T201|COMP|2607-0|LNC|Melanin|Melanin
C0364752|T201|COMP|3129-4|LNC|Menadione|Menadione
C0364753|T201|COMP|11139-3|LNC|Metanephrine|Metanephrine
C0364756|T201|COMP|2611-2|LNC|Methcoproporphyrin|Methcoproporphyrin
C0364757|T201|COMP|2612-0|LNC|Methemalbumin|Methemalbumin
C0364758|T201|COMP|2613-8|LNC|Methemoglobin|Methemoglobin
C0364759|T201|COMP|2614-6|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C0364760|T201|COMP|2615-3|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C0364761|T201|COMP|2616-1|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C0364762|T201|COMP|2617-9|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C0364763|T201|COMP|2619-5|LNC|Methemoglobin|Methemoglobin
C0364764|T201|COMP|2618-7|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C0364765|T201|COMP|2620-3|LNC|Methionine|Methionine
C0364766|T201|COMP|2621-1|LNC|Methionine|Methionine
C0364767|T201|COMP|2622-9|LNC|Methionine|Methionine
C0364768|T201|COMP|2623-7|LNC|Methionine|Methionine
C0364769|T201|COMP|2624-5|LNC|Methionine|Methionine
C0364770|T201|COMP|2625-2|LNC|Methionine adenosyltransferase|Methionine adenosyltransferase
C0364771|T201|COMP|2626-0|LNC|Methoxyacetate|Methoxyacetate
C0364772|T201|COMP|2627-8|LNC|Methylenetetrahydrofolate dehydrogenase.NAD|Methylenetetrahydrofolate dehydrogenase.NAD
C0364773|T201|COMP|2628-6|LNC|Methylenetetrahydrofolate dehydrogenase.NADP|Methylenetetrahydrofolate dehydrogenase.NADP
C0364774|T201|COMP|2629-4|LNC|Methylmalonate|Methylmalonate
C0364775|T201|COMP|2630-2|LNC|Methylmalonate|Methylmalonate
C0364776|T201|COMP|2631-0|LNC|Methylmalonyl CoA mutase|Methylmalonyl CoA mutase
C0364777|T201|COMP|2632-8|LNC|methylTESTOSTERone|methylTESTOSTERone
C0364778|T201|COMP|2633-6|LNC|methylTESTOSTERone|methylTESTOSTERone
C0364779|T201|COMP|2634-4|LNC|methylTESTOSTERone|methylTESTOSTERone
C0364780|T201|COMP|2635-1|LNC|Mianserin|Mianserin
C0364781|T201|COMP|2636-9|LNC|Mianserin|Mianserin
C0364782|T201|COMP|2637-7|LNC|Mucoprotein|Mucoprotein
C0364783|T201|COMP|2638-5|LNC|Myelin basic protein|Myelin basic protein
C0364784|T201|COMP|2639-3|LNC|Myoglobin|Myoglobin
C0364785|T201|COMP|2640-1|LNC|Myoglobin|Myoglobin
C0364786|T201|COMP|2641-9|LNC|Myoglobin|Myoglobin
C0364787|T201|COMP|2642-7|LNC|Myoglobin|Myoglobin
C0364788|T201|COMP|2643-5|LNC|N-acetyl-beta-glucosaminidase|N-acetyl-beta-glucosaminidase
C0364789|T201|COMP|2644-3|LNC|Alpha-N-acetylglucosaminidase|Alpha-N-acetylglucosaminidase
C0364790|T201|COMP|2645-0|LNC|N-Acetylgalactosamine-4-Sulfatase|N-Acetylgalactosamine-4-Sulfatase
C0364791|T201|COMP|2646-8|LNC|N-Acetylgalactosamine-4-Sulfatase|N-Acetylgalactosamine-4-Sulfatase
C0364792|T201|COMP|2647-6|LNC|N-Acetylgalactosamine-4-Sulfatase|N-Acetylgalactosamine-4-Sulfatase
C0364793|T201|COMP|2648-4|LNC|N-Acetylgalactosamine-4-Sulfatase|N-Acetylgalactosamine-4-Sulfatase
C0364794|T201|COMP|2649-2|LNC|N-Acetylgalactosamine-6-Sulfatase|N-Acetylgalactosamine-6-Sulfatase
C0364795|T201|COMP|2650-0|LNC|N-Acetylglucosamine-6-Sulfatase|N-Acetylglucosamine-6-Sulfatase
C0364796|T201|COMP|2651-8|LNC|NADH dehydrogenase|NADH dehydrogenase
C0364797|T201|COMP|2652-6|LNC|NADH dehydrogenase|NADH dehydrogenase
C0364798|T201|COMP|2653-4|LNC|Cytochrome b5 reductase|Cytochrome b5 reductase
C0364799|T201|COMP|2654-2|LNC|Neurophysin|Neurophysin
C0364800|T201|COMP|2655-9|LNC|Neurotensin|Neurotensin
C0364801|T201|COMP|2656-7|LNC|Niacin|Niacin
C0364802|T201|COMP|2657-5|LNC|Nitrite|Nitrite
C0364805|T201|COMP|2660-9|LNC|Nitrogen|Nitrogen
C0364806|T201|COMP|2661-7|LNC|Nitrogen.nonprotein|Nitrogen.nonprotein
C0364807|T201|COMP|2662-5|LNC|Nitrogen.nonprotein|Nitrogen.nonprotein
C0364808|T201|COMP|2663-3|LNC|Nitrogen.nonprotein|Nitrogen.nonprotein
C0364809|T201|COMP|2659-1|LNC|Nitrogen|Nitrogen
C0364809|T201|COMP|2664-1|LNC|Nitrogen|Nitrogen
C0364810|T201|COMP|2665-8|LNC|Nitrogen|Nitrogen
C0364811|T201|COMP|2666-6|LNC|Norepinephrine|Norepinephrine
C0364812|T201|COMP|2667-4|LNC|Norepinephrine|Norepinephrine
C0364813|T201|COMP|2668-2|LNC|Norepinephrine|Norepinephrine
C0364814|T201|COMP|2669-0|LNC|Normetanephrine|Normetanephrine
C0364815|T201|COMP|2670-8|LNC|Normetanephrine|Normetanephrine
C0364816|T201|COMP|2671-6|LNC|Normetanephrine|Normetanephrine
C0364817|T201|COMP|2672-4|LNC|Octopamine|Octopamine
C0364818|T201|COMP|2673-2|LNC|Oleate|Oleate
C0364819|T201|COMP|2674-0|LNC|Ornithine|Ornithine
C0364820|T201|COMP|2675-7|LNC|Ornithine|Ornithine
C0364821|T201|COMP|2676-5|LNC|Organic acids|Organic acids
C0364822|T201|COMP|2677-3|LNC|Organochloride|Organochloride
C0364823|T201|COMP|2678-1|LNC|Ornithine|Ornithine
C0364824|T201|COMP|2679-9|LNC|Ornithine|Ornithine
C0364825|T201|COMP|2680-7|LNC|Ornithine|Ornithine
C0364826|T201|COMP|2681-5|LNC|Ornithine|Ornithine
C0364827|T201|COMP|2682-3|LNC|Ornithine carbamoyltransferase|Ornithine carbamoyltransferase
C0364828|T201|COMP|2683-1|LNC|Ornithine carbamoyltransferase|Ornithine carbamoyltransferase
C0364829|T201|COMP|2686-4|LNC|Orotate|Orotate
C0364830|T201|COMP|2687-2|LNC|Orotate phosphoribosyltransferase|Orotate phosphoribosyltransferase
C0364831|T201|COMP|2688-0|LNC|Orotidine-5'-Phosphate decarboxylase|Orotidine-5'-Phosphate decarboxylase
C0364832|T201|COMP|2689-8|LNC|Osmolality|Osmolality
C0364833|T201|COMP|2690-6|LNC|Osmolality|Osmolality
C0364834|T201|COMP|2691-4|LNC|Osmolality|Osmolality
C0364835|T201|COMP|2692-2|LNC|Osmolality|Osmolality
C0364836|T201|COMP|2693-0|LNC|Osmolality|Osmolality
C0364837|T201|COMP|2694-8|LNC|Osmolality|Osmolality
C0364838|T201|COMP|2695-5|LNC|Osmolality|Osmolality
C0364839|T201|COMP|2696-3|LNC|Osmolality|Osmolality
C0364840|T201|COMP|2697-1|LNC|Osteocalcin|Osteocalcin
C0364841|T201|COMP|2698-9|LNC|Osteonectin|Osteonectin
C0364842|T201|COMP|2699-7|LNC|Oxalate|Oxalate
C0364843|T201|COMP|2700-3|LNC|Oxalate|Oxalate
C0364844|T201|COMP|2701-1|LNC|Oxalate|Oxalate
C0364845|T201|COMP|2702-9|LNC|Oxalate renal clearance|Oxalate renal clearance
C0364846|T201|COMP|19255-9|LNC|Oxygen^^adjusted to patient's actual temperature|Oxygen^^adjusted to patient's actual temperature
C0364847|T201|COMP|19256-7|LNC|Oxygen^^adjusted to patient's actual temperature|Oxygen^^adjusted to patient's actual temperature
C0364848|T201|COMP|19258-3|LNC|Oxygen^^adjusted to patient's actual temperature|Oxygen^^adjusted to patient's actual temperature
C0364849|T201|COMP|2706-0|LNC|Oxygen|Oxygen
C0364850|T201|COMP|2707-8|LNC|Oxygen affinity|Oxygen affinity
C0364851|T201|COMP|2708-6|LNC|Oxygen saturation|Oxygen saturation
C0364856|T201|COMP|2713-6|LNC|Oxygen saturation|Oxygen saturation
C0364857|T201|COMP|2714-4|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C0364858|T201|COMP|2715-1|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C0364859|T201|COMP|2716-9|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C0364860|T201|COMP|2717-7|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C0364861|T201|COMP|2718-5|LNC|Oxytocin|Oxytocin
C0364862|T201|COMP|2719-3|LNC|Palmitate|Palmitate
C0364863|T201|COMP|2720-1|LNC|Palmitoylphosphatidyl choline|Palmitoylphosphatidyl choline
C0364864|T201|COMP|2721-9|LNC|Pancreatic polypeptide|Pancreatic polypeptide
C0364865|T201|COMP|2722-7|LNC|Pantothenate|Pantothenate
C0364867|T201|COMP|2724-3|LNC|Para aminohippurate|Para aminohippurate
C0364868|T201|COMP|2725-0|LNC|Para methylhippurate|Para methylhippurate
C0364869|T201|COMP|2726-8|LNC|Para nitrophenol|Para nitrophenol
C0364870|T201|COMP|2727-6|LNC|Para nitrophenol|Para nitrophenol
C0364871|T201|COMP|2728-4|LNC|Parathion|Parathion
C0364872|T201|COMP|2729-2|LNC|Parathyrin related protein|Parathyrin related protein
C0364873|T201|COMP|2730-0|LNC|Parathyrin.C-terminal|Parathyrin.C-terminal
C0364874|T201|COMP|2731-8|LNC|Parathyrin.intact|Parathyrin.intact
C0364875|T201|COMP|2732-6|LNC|Parathyrin.mid molecule|Parathyrin.mid molecule
C0364876|T201|COMP|2733-4|LNC|Parathyrin.N-terminal|Parathyrin.N-terminal
C0364877|T201|COMP|2734-2|LNC|Pentoses|Pentoses
C0364878|T201|COMP|2735-9|LNC|Pepsinogen|Pepsinogen
C0364879|T201|COMP|2736-7|LNC|Pepsinogen I|Pepsinogen I
C0364880|T201|COMP|2737-5|LNC|Pepsinogen I|Pepsinogen I
C0364881|T201|COMP|2738-3|LNC|Pepsinogen II|Pepsinogen II
C0364882|T201|COMP|2739-1|LNC|Pepsinogen|Pepsinogen
C0364883|T201|COMP|2740-9|LNC|Pepsins|Pepsins
C0364884|T201|COMP|2741-7|LNC|Pepsins|Pepsins
C0364885|T201|COMP|2742-5|LNC|Angiotensin converting enzyme|Angiotensin converting enzyme
C0364900|T201|COMP|2757-3|LNC|Phenol|Phenol
C0364901|T201|COMP|2759-9|LNC|Phenols|Phenols
C0364902|T201|COMP|2760-7|LNC|Phenolsulphonphthalein|Phenolsulphonphthalein
C0364903|T201|COMP|2762-3|LNC|Phenylalanine|Phenylalanine
C0364904|T201|COMP|2763-1|LNC|Phenylalanine|Phenylalanine
C0364905|T201|COMP|2764-9|LNC|Phenylalanine|Phenylalanine
C0364906|T201|COMP|2765-6|LNC|Phenylalanine|Phenylalanine
C0364907|T201|COMP|2766-4|LNC|Phenylalanine|Phenylalanine
C0364908|T201|COMP|2767-2|LNC|Phenylalanine|Phenylalanine
C0364909|T201|COMP|2768-0|LNC|Phenylalanine/Tyrosine|Phenylalanine/Tyrosine
C0364910|T201|COMP|2761-5|LNC|Phenylketones|Phenylketones
C0364911|T201|COMP|2769-8|LNC|Phenylketones|Phenylketones
C0364912|T201|COMP|2770-6|LNC|Phenylpyruvate|Phenylpyruvate
C0364913|T201|COMP|2771-4|LNC|Phenylpyruvate|Phenylpyruvate
C0364914|T201|COMP|2772-2|LNC|Phenylpyruvate|Phenylpyruvate
C0364915|T201|COMP|2773-0|LNC|Phenylpyruvate|Phenylpyruvate
C0364916|T201|COMP|2774-8|LNC|Phosphate|Phosphate
C0364917|T201|COMP|2775-5|LNC|Phosphate|Phosphate
C0364918|T201|COMP|2776-3|LNC|Phosphate renal clearance|Phosphate renal clearance
C0364922|T201|COMP|2780-5|LNC|Phosphate|Phosphate
C0364923|T201|COMP|2778-9|LNC|Phosphate|Phosphate
C0364924|T201|COMP|2779-7|LNC|Phosphate|Phosphate
C0364925|T201|COMP|2783-9|LNC|Lecithin|Lecithin
C0364926|T201|COMP|2784-7|LNC|Phosphatidylcholine.saturated|Phosphatidylcholine.saturated
C0364927|T201|COMP|2785-4|LNC|Phosphatidylglycerol|Phosphatidylglycerol
C0364928|T201|COMP|2786-2|LNC|Phosphatidylglycerol|Phosphatidylglycerol
C0364929|T201|COMP|2787-0|LNC|Phosphatidylinositol|Phosphatidylinositol
C0364930|T201|COMP|2788-8|LNC|Phosphoenolpyruvate carboxykinase|Phosphoenolpyruvate carboxykinase
C0364931|T201|COMP|2789-6|LNC|Phosphoethanolamine|Phosphoethanolamine
C0364932|T201|COMP|2790-4|LNC|Phosphoethanolamine|Phosphoethanolamine
C0364933|T201|COMP|2791-2|LNC|Phosphofructokinase|Phosphofructokinase
C0364934|T201|COMP|2792-0|LNC|Phosphofructokinase|Phosphofructokinase
C0364939|T201|COMP|2797-9|LNC|Phosphoglucomutase|Phosphoglucomutase
C0364940|T201|COMP|2798-7|LNC|Phosphoglycerate kinase|Phosphoglycerate kinase
C0364941|T201|COMP|2799-5|LNC|Phosphoglyceromutase|Phosphoglyceromutase
C0364942|T201|COMP|2800-1|LNC|Glucose phosphate isomerase|Glucose phosphate isomerase
C0364943|T201|COMP|2568-4|LNC|Phospholipid|Phospholipid
C0364944|T201|COMP|2802-7|LNC|Phosphoserine|Phosphoserine
C0364945|T201|COMP|2804-3|LNC|Phytanate|Phytanate
C0364947|T201|COMP|2805-0|LNC|Pipecolate|Pipecolate
C0364948|T201|COMP|2806-8|LNC|Pipecolate|Pipecolate
C0364949|T201|COMP|2807-6|LNC|Pipecolate|Pipecolate
C0364950|T201|COMP|2808-4|LNC|Porphobilin|Porphobilin
C0364951|T201|COMP|2809-2|LNC|Porphobilinogen|Porphobilinogen
C0364952|T201|COMP|2810-0|LNC|Porphobilinogen|Porphobilinogen
C0364953|T201|COMP|2811-8|LNC|Porphobilinogen|Porphobilinogen
C0364954|T201|COMP|2812-6|LNC|Porphobilinogen deaminase|Porphobilinogen deaminase
C0364955|T201|COMP|2813-4|LNC|Porphobilinogen synthase|Porphobilinogen synthase
C0364956|T201|COMP|2814-2|LNC|Porphyrins|Porphyrins
C0364957|T201|COMP|2815-9|LNC|Porphyrins|Porphyrins
C0364958|T201|COMP|2816-7|LNC|Porphyrins|Porphyrins
C0364959|T201|COMP|2817-5|LNC|Porphyrins|Porphyrins
C0364960|T201|COMP|2818-3|LNC|Porphyrins|Porphyrins
C0364961|T201|COMP|6298-4|LNC|Potassium|Potassium
C0364962|T201|COMP|2819-1|LNC|Potassium|Potassium
C0364963|T201|COMP|2820-9|LNC|Potassium|Potassium
C0364964|T201|COMP|2821-7|LNC|Potassium|Potassium
C0364965|T201|COMP|2822-5|LNC|Potassium|Potassium
C0364966|T201|COMP|2824-1|LNC|Potassium|Potassium
C0364967|T201|COMP|2825-8|LNC|Potassium|Potassium
C0364968|T201|COMP|2823-3|LNC|Potassium|Potassium
C0364969|T201|COMP|2826-6|LNC|Potassium|Potassium
C0364970|T201|COMP|2827-4|LNC|Potassium|Potassium
C0364971|T201|COMP|2828-2|LNC|Potassium|Potassium
C0364972|T201|COMP|2829-0|LNC|Potassium|Potassium
C0364973|T201|COMP|2830-8|LNC|Potassium renal clearance|Potassium renal clearance
C0364974|T201|COMP|2831-6|LNC|Pregnancy specific protein 1|Pregnancy specific protein 1
C0364975|T201|COMP|2832-4|LNC|Pregnanediol|Pregnanediol
C0364976|T201|COMP|2833-2|LNC|Pregnanediol|Pregnanediol
C0364977|T201|COMP|2834-0|LNC|Pregnanediol|Pregnanediol
C0364978|T201|COMP|2835-7|LNC|Pregnanetriol|Pregnanetriol
C0364979|T201|COMP|2836-5|LNC|Pregnanetriol|Pregnanetriol
C0364980|T201|COMP|2837-3|LNC|Pregnenolone|Pregnenolone
C0364981|T201|COMP|2838-1|LNC|Progesterone|Progesterone
C0364982|T201|COMP|2839-9|LNC|Progesterone|Progesterone
C0364983|T201|COMP|2840-7|LNC|Proinsulin|Proinsulin
C0364986|T201|COMP|2843-1|LNC|Proline|Proline
C0364987|T201|COMP|2844-9|LNC|Proline|Proline
C0364988|T201|COMP|2845-6|LNC|Proline|Proline
C0364989|T201|COMP|2846-4|LNC|Proline|Proline
C0364990|T201|COMP|2847-2|LNC|Proline|Proline
C0364991|T201|COMP|2848-0|LNC|Proline dipeptidase|Proline dipeptidase
C0364992|T201|COMP|2849-8|LNC|Propionate|Propionate
C0364993|T201|COMP|2850-6|LNC|Propionyl CO-A carboxylase|Propionyl CO-A carboxylase
C0364994|T201|COMP|2851-4|LNC|Prostaglandin E|Prostaglandin E
C0364995|T201|COMP|2852-2|LNC|Prostaglandin E1|Prostaglandin E1
C0364996|T201|COMP|2853-0|LNC|Prostaglandin E2|Prostaglandin E2
C0364997|T201|COMP|2854-8|LNC|Prostaglandin F|Prostaglandin F
C0364998|T201|COMP|2855-5|LNC|Prostaglandin F2|Prostaglandin F2
C0364999|T201|COMP|2856-3|LNC|Prostaglandin|Prostaglandin
C0365000|T201|COMP|2857-1|LNC|Prostate specific Ag|Prostate specific Ag
C0365001|T201|COMP|2858-9|LNC|Protein.CSF/Protein.serum|Protein.CSF/Protein.serum
C0365002|T201|COMP|2859-7|LNC|Protein kinase|Protein kinase
C0365003|T201|COMP|2860-5|LNC|Protein nitrogen|Protein nitrogen
C0365004|T201|COMP|2861-3|LNC|Albumin|Albumin
C0365005|T201|COMP|2862-1|LNC|Albumin|Albumin
C0365006|T201|COMP|2863-9|LNC|Albumin|Albumin
C0365007|T201|COMP|2864-7|LNC|Alpha 1 globulin|Alpha 1 globulin
C0365008|T201|COMP|2865-4|LNC|Alpha 1 globulin|Alpha 1 globulin
C0365009|T201|COMP|2866-2|LNC|Alpha 1 globulin|Alpha 1 globulin
C0365010|T201|COMP|2867-0|LNC|Alpha 2 globulin|Alpha 2 globulin
C0365011|T201|COMP|2868-8|LNC|Alpha 2 globulin|Alpha 2 globulin
C0365012|T201|COMP|2869-6|LNC|Alpha 2 globulin|Alpha 2 globulin
C0365013|T201|COMP|2870-4|LNC|Beta globulin|Beta globulin
C0365014|T201|COMP|2871-2|LNC|Beta globulin|Beta globulin
C0365015|T201|COMP|2872-0|LNC|Beta globulin|Beta globulin
C0365016|T201|COMP|2873-8|LNC|Gamma globulin|Gamma globulin
C0365017|T201|COMP|2874-6|LNC|Gamma globulin|Gamma globulin
C0365018|T201|COMP|2875-3|LNC|Gamma globulin|Gamma globulin
C0365019|T201|COMP|2876-1|LNC|Prealbumin|Prealbumin
C0365020|T201|COMP|2877-9|LNC|Prealbumin|Prealbumin
C0365021|T201|COMP|2878-7|LNC|Protein|Protein
C0365022|T201|COMP|2879-5|LNC|Protein|Protein
C0365023|T201|COMP|2880-3|LNC|Protein|Protein
C0365024|T201|COMP|5920-4|LNC|Protein|Protein
C0365025|T201|COMP|2881-1|LNC|Protein|Protein
C0365026|T201|COMP|2882-9|LNC|Protein|Protein
C0365027|T201|COMP|2883-7|LNC|Protein|Protein
C0365028|T201|COMP|2884-5|LNC|Protein|Protein
C0365029|T201|COMP|2885-2|LNC|Protein|Protein
C0365030|T201|COMP|2886-0|LNC|Protein|Protein
C0365031|T201|COMP|2887-8|LNC|Protein|Protein
C0365032|T201|COMP|2888-6|LNC|Protein|Protein
C0365033|T201|COMP|2889-4|LNC|Protein|Protein
C0365034|T201|COMP|2890-2|LNC|Protein/Creatinine|Protein/Creatinine
C0365035|T201|COMP|2891-0|LNC|Protoporphyrin|Protoporphyrin
C0365036|T201|COMP|2892-8|LNC|Protoporphyrin.free|Protoporphyrin.free
C0365037|T201|COMP|2893-6|LNC|Protoporphyrin.zinc|Protoporphyrin.zinc
C0365038|T201|COMP|2894-4|LNC|Protoporphyrin.zinc|Protoporphyrin.zinc
C0365039|T201|COMP|2895-1|LNC|Protoporphyrin.zinc|Protoporphyrin.zinc
C0365040|T201|COMP|2896-9|LNC|Protoporphyrin|Protoporphyrin
C0365041|T201|COMP|2897-7|LNC|Protoporphyrin|Protoporphyrin
C0365042|T201|COMP|2898-5|LNC|Protoporphyrin|Protoporphyrin
C0365043|T201|COMP|2899-3|LNC|Purine nucleoside phosphorylase|Purine nucleoside phosphorylase
C0365044|T201|COMP|2900-9|LNC|Pyridoxine|Pyridoxine
C0365045|T201|COMP|2901-7|LNC|Pyridoxine congeners|Pyridoxine congeners
C0365046|T201|COMP|2902-5|LNC|Pyrimidine-5'-Nucleotidase|Pyrimidine-5'-Nucleotidase
C0365047|T201|COMP|2903-3|LNC|Pyrimidine-5'-Nucleotidase|Pyrimidine-5'-Nucleotidase
C0365048|T201|COMP|2904-1|LNC|Pyrophosphate crystals|Pyrophosphate crystals
C0365049|T201|COMP|2905-8|LNC|Pyruvate|Pyruvate
C0365050|T201|COMP|2906-6|LNC|Pyruvate|Pyruvate
C0365051|T201|COMP|2907-4|LNC|Pyruvate|Pyruvate
C0365052|T201|COMP|2908-2|LNC|Pyruvate|Pyruvate
C0365053|T201|COMP|2909-0|LNC|Pyruvate carboxylase|Pyruvate carboxylase
C0365054|T201|COMP|2910-8|LNC|Pyruvate dehydrogenase.cytochrome|Pyruvate dehydrogenase.cytochrome
C0365055|T201|COMP|2911-6|LNC|Pyruvate dehydrogenase.lipoamide|Pyruvate dehydrogenase.lipoamide
C0365056|T201|COMP|2912-4|LNC|Pyruvate kinase|Pyruvate kinase
C0365057|T201|COMP|2913-2|LNC|Pyruvate kinase|Pyruvate kinase
C0365058|T201|COMP|2914-0|LNC|Pyruvate oxidase|Pyruvate oxidase
C0365059|T201|COMP|2915-7|LNC|Renin|Renin
C0365060|T201|COMP|2916-5|LNC|Renin renal clearance|Renin renal clearance
C0365061|T201|COMP|2917-3|LNC|Renin^supine|Renin^supine
C0365062|T201|COMP|2918-1|LNC|Renin^upright|Renin^upright
C0365063|T201|COMP|2919-9|LNC|Reticulin|Reticulin
C0365064|T201|COMP|2920-7|LNC|Retinal|Retinal
C0365065|T201|COMP|2921-5|LNC|Retinoate|Retinoate
C0365066|T201|COMP|2922-3|LNC|Retinol|Retinol
C0365067|T201|COMP|2923-1|LNC|Retinol|Retinol
C0365068|T201|COMP|2924-9|LNC|Riboflavin|Riboflavin
C0365069|T201|COMP|2925-6|LNC|Ribonuclease|Ribonuclease
C0365070|T201|COMP|2926-4|LNC|Ribose|Ribose
C0365071|T201|COMP|2927-2|LNC|Ribulose|Ribulose
C0365072|T201|COMP|1938-0|LNC|Beta fructofuranosidase|Beta fructofuranosidase
C0365073|T201|COMP|2929-8|LNC|Saccharides|Saccharides
C0365074|T201|COMP|2930-6|LNC|Sarcosine|Sarcosine
C0365075|T201|COMP|2931-4|LNC|Sarcosine|Sarcosine
C0365076|T201|COMP|2932-2|LNC|Sarcosine|Sarcosine
C0365077|T201|COMP|2933-0|LNC|Secretin|Secretin
C0365078|T201|COMP|2934-8|LNC|Serine|Serine
C0365079|T201|COMP|2935-5|LNC|Serine|Serine
C0365080|T201|COMP|2936-3|LNC|Serine|Serine
C0365081|T201|COMP|2937-1|LNC|Serine|Serine
C0365082|T201|COMP|2938-9|LNC|Serine|Serine
C0365083|T201|COMP|2939-7|LNC|Serotonin|Serotonin
C0365084|T201|COMP|2940-5|LNC|Serotonin|Serotonin
C0365085|T201|COMP|2941-3|LNC|Serotonin|Serotonin
C0365086|T201|COMP|2942-1|LNC|Sex hormone binding globulin|Sex hormone binding globulin
C0365087|T201|COMP|2943-9|LNC|Sialate|Sialate
C0365088|T201|COMP|2944-7|LNC|Sialate|Sialate
C0365089|T201|COMP|2945-4|LNC|Sialidase|Sialidase
C0365090|T201|COMP|2946-2|LNC|Sialidase|Sialidase
C0365091|T201|COMP|2947-0|LNC|Sodium|Sodium
C0365092|T201|COMP|2948-8|LNC|Sodium|Sodium
C0365093|T201|COMP|2949-6|LNC|Sodium|Sodium
C0365094|T201|COMP|2950-4|LNC|Sodium|Sodium
C0365095|T201|COMP|2951-2|LNC|Sodium|Sodium
C0365096|T201|COMP|2952-0|LNC|Sodium|Sodium
C0365097|T201|COMP|2953-8|LNC|Sodium|Sodium
C0365098|T201|COMP|2954-6|LNC|Sodium|Sodium
C0365099|T201|COMP|2955-3|LNC|Sodium|Sodium
C0365100|T201|COMP|2956-1|LNC|Sodium|Sodium
C0365101|T201|COMP|2957-9|LNC|Sodium renal clearance|Sodium renal clearance
C0365102|T201|COMP|2958-7|LNC|Sodium/Potassium|Sodium/Potassium
C0365103|T201|COMP|2959-5|LNC|Sodium/Potassium|Sodium/Potassium
C0365104|T201|COMP|2486-9|LNC|Somatomedins|Somatomedins
C0365105|T201|COMP|2960-3|LNC|Somatostatin|Somatostatin
C0365106|T201|COMP|2961-1|LNC|Somatostatin|Somatostatin
C0365107|T201|COMP|2962-9|LNC|Somatotropin|Somatotropin
C0365108|T201|COMP|2963-7|LNC|Somatotropin|Somatotropin
C0365109|T201|COMP|2964-5|LNC|Specific gravity|Specific gravity
C0365110|T201|COMP|2966-0|LNC|Specific gravity|Specific gravity
C0365111|T201|COMP|2965-2|LNC|Specific gravity|Specific gravity
C0365112|T201|COMP|2967-8|LNC|Starch granules|Starch granules
C0365113|T201|COMP|2968-6|LNC|Starch granules|Starch granules
C0365114|T201|COMP|2969-4|LNC|Stercobilin|Stercobilin
C0365115|T201|COMP|2970-2|LNC|Streptomyces proteinase|Streptomyces proteinase
C0365116|T201|COMP|2971-0|LNC|Substance P|Substance P
C0365117|T201|COMP|2972-8|LNC|Succinate|Succinate
C0365118|T201|COMP|2973-6|LNC|Succinylacetone|Succinylacetone
C0365119|T201|COMP|2974-4|LNC|Sucrose|Sucrose
C0365120|T201|COMP|2975-1|LNC|Sulfate|Sulfate
C0365121|T201|COMP|2976-9|LNC|Sulfate.inorganic|Sulfate.inorganic
C0365122|T201|COMP|2977-7|LNC|Sulfite oxidase|Sulfite oxidase
C0365123|T201|COMP|2978-5|LNC|Superoxide dismutase|Superoxide dismutase
C0365124|T201|COMP|2979-3|LNC|Taurine|Taurine
C0365125|T201|COMP|2980-1|LNC|Taurine|Taurine
C0365126|T201|COMP|2981-9|LNC|Taurine|Taurine
C0365127|T201|COMP|2982-7|LNC|Taurine|Taurine
C0365128|T201|COMP|2984-3|LNC|Testosterone|Testosterone
C0365129|T201|COMP|2985-0|LNC|Testosterone|Testosterone
C0365131|T201|COMP|2987-6|LNC|Testosterone|Testosterone
C0365132|T201|COMP|2988-4|LNC|Testosterone|Testosterone
C0365133|T201|COMP|2989-2|LNC|Testosterone|Testosterone
C0365134|T201|COMP|2990-0|LNC|Testosterone.free+weakly bound|Testosterone.free+weakly bound
C0365135|T201|COMP|2991-8|LNC|Testosterone.free|Testosterone.free
C0365136|T201|COMP|2992-6|LNC|Testosterone|Testosterone
C0365137|T201|COMP|2986-8|LNC|Testosterone|Testosterone
C0365138|T201|COMP|2994-2|LNC|Testosterone.free|Testosterone.free
C0365139|T201|COMP|2995-9|LNC|Tetrahydrocortisol|Tetrahydrocortisol
C0365140|T201|COMP|2996-7|LNC|Tetrahydrodeoxycortisol|Tetrahydrodeoxycortisol
C0365141|T201|COMP|2997-5|LNC|Tetrahydrofolate|Tetrahydrofolate
C0365142|T201|COMP|2998-3|LNC|Thiamine|Thiamine
C0365143|T201|COMP|2999-1|LNC|Thiamine|Thiamine
C0365144|T201|COMP|3000-7|LNC|Thiamine pyrophosphate|Thiamine pyrophosphate
C0365145|T201|COMP|3001-5|LNC|Thiocyanate|Thiocyanate
C0365146|T201|COMP|3002-3|LNC|Thiocyanate|Thiocyanate
C0365147|T201|COMP|3003-1|LNC|Thiocyanate|Thiocyanate
C0365148|T201|COMP|3004-9|LNC|Thiocyanate|Thiocyanate
C0365149|T201|COMP|3005-6|LNC|Thiosulfate renal clearance|Thiosulfate renal clearance
C0365150|T201|COMP|3006-4|LNC|Threonine|Threonine
C0365151|T201|COMP|3007-2|LNC|Threonine|Threonine
C0365152|T201|COMP|3008-0|LNC|Threonine|Threonine
C0365153|T201|COMP|3009-8|LNC|Threonine|Threonine
C0365154|T201|COMP|3010-6|LNC|Threonine|Threonine
C0365155|T201|COMP|3011-4|LNC|Thromboxane alpha 2|Thromboxane alpha 2
C0365156|T201|COMP|3012-2|LNC|Thromboxane beta 2|Thromboxane beta 2
C0365157|T201|COMP|3013-0|LNC|Thyroglobulin|Thyroglobulin
C0365158|T201|COMP|3014-8|LNC|Thyroid stimulating immunoglobulins|Thyroid stimulating immunoglobulins
C0365159|T201|COMP|3015-5|LNC|Thyrotropin|Thyrotropin
C0365160|T201|COMP|3016-3|LNC|Thyrotropin|Thyrotropin
C0365161|T201|COMP|3017-1|LNC|Thyrotropin binding inhibitory immunoglobulins|Thyrotropin binding inhibitory immunoglobulins
C0365162|T201|COMP|3018-9|LNC|Thyrotropin releasing hormone|Thyrotropin releasing hormone
C0365163|T201|COMP|3019-7|LNC|Thyrotropin.long acting|Thyrotropin.long acting
C0365164|T201|COMP|3020-5|LNC|Thyroxine binding globulin|Thyroxine binding globulin
C0365165|T201|COMP|3021-3|LNC|Thyroxine binding globulin|Thyroxine binding globulin
C0365166|T201|COMP|3022-1|LNC|Thyroxine free index|Thyroxine free index
C0365167|T201|COMP|3023-9|LNC|Thyroxine uptake|Thyroxine uptake
C0365168|T201|COMP|3024-7|LNC|Thyroxine.free|Thyroxine.free
C0365169|T201|COMP|3025-4|LNC|Thyroxine|Thyroxine
C0365170|T201|COMP|3026-2|LNC|Thyroxine|Thyroxine
C0365171|T201|COMP|3027-0|LNC|Thyroxine/Thyroxine binding globulin|Thyroxine/Thyroxine binding globulin
C0365172|T201|COMP|3028-8|LNC|Thyroxine/Triiodothyronine uptake index|Thyroxine/Triiodothyronine uptake index
C0365173|T201|COMP|3029-6|LNC|Transcobalamin I|Transcobalamin I
C0365174|T201|COMP|3030-4|LNC|Transcobalamin II|Transcobalamin II
C0365175|T201|COMP|3031-2|LNC|Transcobalamin III|Transcobalamin III
C0365176|T201|COMP|3032-0|LNC|Transcobalamin|Transcobalamin
C0365177|T201|COMP|3033-8|LNC|Transcortin|Transcortin
C0365178|T201|COMP|3034-6|LNC|Transferrin|Transferrin
C0365179|T201|COMP|3035-3|LNC|Transferrin|Transferrin
C0365180|T201|COMP|3036-1|LNC|Transketolase|Transketolase
C0365181|T201|COMP|3037-9|LNC|Prealbumin|Prealbumin
C0365182|T201|COMP|3038-7|LNC|Trehalase|Trehalase
C0365183|T201|COMP|3039-5|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C0365184|T201|COMP|3040-3|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C0365185|T201|COMP|3041-1|LNC|Trichloroacetate|Trichloroacetate
C0365187|T201|COMP|3043-7|LNC|Triglyceride|Triglyceride
C0365188|T201|COMP|3044-5|LNC|Triglyceride+ester.in HDL|Triglyceride+ester.in HDL
C0365189|T201|COMP|3045-2|LNC|Triglyceride+ester.in IDL|Triglyceride+ester.in IDL
C0365190|T201|COMP|3046-0|LNC|Triglyceride+ester.in LDL|Triglyceride+ester.in LDL
C0365191|T201|COMP|3047-8|LNC|Triglyceride+ester.in VLDL|Triglyceride+ester.in VLDL
C0365192|T201|COMP|3048-6|LNC|Triglyceride^post CFst|Triglyceride^post CFst
C0365193|T201|COMP|3049-4|LNC|Triglyceride|Triglyceride
C0365194|T201|COMP|3050-2|LNC|Triiodothyronine resin uptake (T3RU)|Triiodothyronine resin uptake (T3RU)
C0365195|T201|COMP|3051-0|LNC|Triiodothyronine.free|Triiodothyronine.free
C0365196|T201|COMP|3052-8|LNC|Triiodothyronine.reverse|Triiodothyronine.reverse
C0365197|T201|COMP|3053-6|LNC|Triiodothyronine|Triiodothyronine
C0365198|T201|COMP|3054-4|LNC|Triiodothyronine.true|Triiodothyronine.true
C0365199|T201|COMP|3055-1|LNC|Triiodothyronine/Triiodothyronine uptake index|Triiodothyronine/Triiodothyronine uptake index
C0365200|T201|COMP|3056-9|LNC|Trimethylamine|Trimethylamine
C0365201|T201|COMP|3057-7|LNC|Triokinase|Triokinase
C0365202|T201|COMP|3058-5|LNC|Triosephosphate isomerase|Triosephosphate isomerase
C0365203|T201|COMP|3059-3|LNC|Trypsin|Trypsin
C0365204|T201|COMP|3060-1|LNC|Trypsin|Trypsin
C0365205|T201|COMP|3063-5|LNC|Trypsin|Trypsin
C0365206|T201|COMP|3061-9|LNC|Trypsin|Trypsin
C0365207|T201|COMP|3062-7|LNC|Trypsin|Trypsin
C0365208|T201|COMP|3064-3|LNC|Trypsin+Trypsinogen|Trypsin+Trypsinogen
C0365209|T201|COMP|3065-0|LNC|Trypsinogen|Trypsinogen
C0365210|T201|COMP|3066-8|LNC|Trypsinogen|Trypsinogen
C0365211|T201|COMP|3067-6|LNC|Trypsinogen I.free|Trypsinogen I.free
C0365212|T201|COMP|3068-4|LNC|Tryptophan|Tryptophan
C0365213|T201|COMP|3069-2|LNC|Tryptophan|Tryptophan
C0365214|T201|COMP|3070-0|LNC|Tryptophan|Tryptophan
C0365215|T201|COMP|3071-8|LNC|Tryptophan|Tryptophan
C0365216|T201|COMP|3072-6|LNC|Tryptophan|Tryptophan
C0365217|T201|COMP|3073-4|LNC|Tryptophan.free|Tryptophan.free
C0365218|T201|COMP|3074-2|LNC|Tumor necrosis factor.alpha|Tumor necrosis factor.alpha
C0365219|T201|COMP|3075-9|LNC|Tyramine|Tyramine
C0365220|T201|COMP|3076-7|LNC|Tyramine|Tyramine
C0365221|T201|COMP|3077-5|LNC|Tyrosine|Tyrosine
C0365222|T201|COMP|3078-3|LNC|Tyrosine|Tyrosine
C0365223|T201|COMP|3079-1|LNC|Tyrosine|Tyrosine
C0365224|T201|COMP|3080-9|LNC|Tyrosine|Tyrosine
C0365225|T201|COMP|3081-7|LNC|Tyrosine|Tyrosine
C0365226|T201|COMP|3082-5|LNC|Tyrosine aminotransferase|Tyrosine aminotransferase
C0365227|T201|COMP|3083-3|LNC|Urate|Urate
C0365228|T201|COMP|3084-1|LNC|Urate|Urate
C0365229|T201|COMP|3085-8|LNC|Urate|Urate
C0365230|T201|COMP|3086-6|LNC|Urate|Urate
C0365231|T201|COMP|3087-4|LNC|Urate|Urate
C0365232|T201|COMP|3088-2|LNC|Urate renal clearance|Urate renal clearance
C0365233|T201|COMP|3089-0|LNC|Urate/Creatinine|Urate/Creatinine
C0365234|T201|COMP|3090-8|LNC|Urea|Urea
C0365235|T201|COMP|3091-6|LNC|Urea|Urea
C0365236|T201|COMP|3092-4|LNC|Urea|Urea
C0365237|T201|COMP|6299-2|LNC|Urea nitrogen|Urea nitrogen
C0365238|T201|COMP|5918-8|LNC|Urea nitrogen|Urea nitrogen
C0365239|T201|COMP|3093-2|LNC|Urea nitrogen|Urea nitrogen
C0365240|T201|COMP|3094-0|LNC|Urea nitrogen|Urea nitrogen
C0365241|T201|COMP|3095-7|LNC|Urea nitrogen|Urea nitrogen
C0365242|T201|COMP|3096-5|LNC|Urea nitrogen|Urea nitrogen
C0365243|T201|COMP|3097-3|LNC|Urea nitrogen/Creatinine|Urea nitrogen/Creatinine
C0365244|T201|COMP|3098-1|LNC|Urea renal clearance|Urea renal clearance
C0365245|T201|COMP|3099-9|LNC|Uridine diphosphate glucose-4-Epimerase|Uridine diphosphate glucose-4-Epimerase
C0365246|T201|COMP|3100-5|LNC|Uridyl transferase|Uridyl transferase
C0365247|T201|COMP|3101-3|LNC|Uridyl transferase|Uridyl transferase
C0365248|T201|COMP|3102-1|LNC|Urobilin|Urobilin
C0365249|T201|COMP|3103-9|LNC|Urobilin|Urobilin
C0365250|T201|COMP|3104-7|LNC|Urobilin|Urobilin
C0365251|T201|COMP|3105-4|LNC|Urobilinogen|Urobilinogen
C0365252|T201|COMP|3106-2|LNC|Urobilinogen|Urobilinogen
C0365253|T201|COMP|3107-0|LNC|Urobilinogen|Urobilinogen
C0365254|T201|COMP|3108-8|LNC|Urobilinogen|Urobilinogen
C0365255|T201|COMP|3109-6|LNC|Urobilinogen|Urobilinogen
C0365256|T201|COMP|3110-4|LNC|Uronate|Uronate
C0365257|T201|COMP|3112-0|LNC|Uroporphyrin|Uroporphyrin
C0365258|T201|COMP|3113-8|LNC|Uroporphyrin|Uroporphyrin
C0365259|T201|COMP|3111-2|LNC|Uroporphyrin 1 isomer|Uroporphyrin 1 isomer
C0365260|T201|COMP|3114-6|LNC|Uroporphyrinogen decarboxylase|Uroporphyrinogen decarboxylase
C0365261|T201|COMP|3115-3|LNC|Uroporphyrinogen III synthase|Uroporphyrinogen III synthase
C0365262|T201|COMP|3116-1|LNC|Valine|Valine
C0365263|T201|COMP|3117-9|LNC|Valine|Valine
C0365264|T201|COMP|3118-7|LNC|Valine|Valine
C0365265|T201|COMP|3119-5|LNC|Valine|Valine
C0365266|T201|COMP|3120-3|LNC|Valine|Valine
C0365267|T201|COMP|3121-1|LNC|Vanillylmandelate|Vanillylmandelate
C0365268|T201|COMP|3122-9|LNC|Vanillylmandelate|Vanillylmandelate
C0365269|T201|COMP|3123-7|LNC|Vanillylmandelate/Creatine|Vanillylmandelate/Creatine
C0365270|T201|COMP|3124-5|LNC|Vanillylmandelate/Creatinine|Vanillylmandelate/Creatinine
C0365271|T201|COMP|3125-2|LNC|Vasoactive intestinal peptide|Vasoactive intestinal peptide
C0365272|T201|COMP|3126-0|LNC|Vasopressin|Vasopressin
C0365273|T201|COMP|3127-8|LNC|Viscosity|Viscosity
C0365274|T201|COMP|3128-6|LNC|Viscosity|Viscosity
C0365275|T201|COMP|3130-2|LNC|Vitronectin|Vitronectin
C0365276|T201|COMP|3131-0|LNC|Xanthine|Xanthine
C0365277|T201|COMP|3132-8|LNC|Xanthine|Xanthine
C0365278|T201|COMP|3133-6|LNC|Xanthurenate|Xanthurenate
C0365279|T201|COMP|3134-4|LNC|Xylose|Xylose
C0365280|T201|COMP|3135-1|LNC|Xylose|Xylose
C0365281|T201|COMP|3136-9|LNC|Xylulose|Xylulose
C0365293|T201|COMP|3148-4|LNC|Oxygen|Oxygen
C0365294|T201|COMP|3149-2|LNC|Oxygen|Oxygen
C0365298|T201|COMP|3153-4|LNC|Specimen weight|Specimen weight
C0365299|T201|COMP|3154-2|LNC|Specimen weight|Specimen weight
C0365300|T201|COMP|3155-9|LNC|Specimen mass|Specimen mass
C0365301|T201|COMP|3156-7|LNC|Specimen volume|Specimen volume
C0365302|T201|COMP|3157-5|LNC|Specimen volume|Specimen volume
C0365303|T201|COMP|3158-3|LNC|Specimen volume|Specimen volume
C0365304|T201|COMP|3159-1|LNC|Specimen volume|Specimen volume
C0365305|T201|COMP|3160-9|LNC|Specimen volume|Specimen volume
C0365306|T201|COMP|3161-7|LNC|Specimen volume|Specimen volume
C0365307|T201|COMP|3162-5|LNC|Specimen volume|Specimen volume
C0365308|T201|COMP|3163-3|LNC|Specimen volume|Specimen volume
C0365309|T201|COMP|3164-1|LNC|Specimen volume|Specimen volume
C0365310|T201|COMP|3165-8|LNC|Specimen volume|Specimen volume
C0365311|T201|COMP|3166-6|LNC|Specimen volume|Specimen volume
C0365312|T201|COMP|3167-4|LNC|Specimen volume|Specimen volume
C0365313|T201|COMP|3168-2|LNC|Specimen volume|Specimen volume
C0365314|T201|COMP|3169-0|LNC|Specimen volume|Specimen volume
C0365315|T201|COMP|3170-8|LNC|Specimen volume|Specimen volume
C0365316|T201|COMP|3171-6|LNC|Specimen.dry weight|Specimen.dry weight
C0365322|T201|COMP|3178-1|LNC|Bleeding time|Bleeding time
C0365323|T201|COMP|3179-9|LNC|Bleeding time|Bleeding time
C0365324|T201|COMP|3180-7|LNC|Cardiolipin Ab|Cardiolipin Ab
C0365325|T201|COMP|3181-5|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C0365326|T201|COMP|3182-3|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C0365327|T201|COMP|3183-1|LNC|Clotting time|Clotting time
C0365329|T201|COMP|6303-2|LNC|Coagulation dilute Russell viper venom induced|Coagulation dilute Russell viper venom induced
C0365392|T201|COMP|3173-2|LNC|Coagulation surface induced|Coagulation surface induced
C0365393|T201|COMP|5898-2|LNC|Coagulation surface induced|Coagulation surface induced
C0365405|T201|COMP|5964-2|LNC|Coagulation tissue factor induced|Coagulation tissue factor induced
C0365422|T201|COMP|3245-8|LNC|Coagulum retraction|Coagulum retraction
C0365429|T201|COMP|3252-4|LNC|Fibrin+Fibrinogen fragments|Fibrin+Fibrinogen fragments
C0365431|T201|COMP|3254-0|LNC|Fibrin.soluble|Fibrin.soluble
C0365444|T201|COMP|3267-2|LNC|Heparin Ab|Heparin Ab
C0365449|T201|COMP|3272-2|LNC|Heparin.low molecular weight|Heparin.low molecular weight
C0365452|T201|COMP|3275-5|LNC|Heparin.unfractionated|Heparin.unfractionated
C0365457|T201|COMP|3280-5|LNC|Kininogen.low molecular weight|Kininogen.low molecular weight
C0365462|T201|COMP|3285-4|LNC|Phospholipid Ab|Phospholipid Ab
C0365463|T201|COMP|3286-2|LNC|Phospholipid Ab.IgG|Phospholipid Ab.IgG
C0365464|T201|COMP|3287-0|LNC|Phospholipid Ab.IgM|Phospholipid Ab.IgM
C0365471|T201|COMP|5971-7|LNC|Plasminogen activator tissue type Ag|Plasminogen activator tissue type Ag
C0365475|T201|COMP|5976-6|LNC|Plasminogen activator inhibitor 1|Plasminogen activator inhibitor 1
C0365485|T201|COMP|5984-0|LNC|Plasminogen activator urokinase type|Plasminogen activator urokinase type
C0365493|T201|COMP|5993-1|LNC|Platelet aggregation.arachidonate induced|Platelet aggregation.arachidonate induced
C0365494|T201|COMP|5994-9|LNC|Platelet aggregation.calcium ionophore induced|Platelet aggregation.calcium ionophore induced
C0365495|T201|COMP|5995-6|LNC|Platelet aggregation.collagen induced|Platelet aggregation.collagen induced
C0365496|T201|COMP|5996-4|LNC|Platelet aggregation.EPINEPHrine induced|Platelet aggregation.EPINEPHrine induced
C0365497|T201|COMP|5997-2|LNC|Platelet aggregation.norepinephrine induced|Platelet aggregation.norepinephrine induced
C0365498|T201|COMP|5998-0|LNC|Platelet aggregation.ristocetin induced|Platelet aggregation.ristocetin induced
C0365499|T201|COMP|5999-8|LNC|Platelet aggregation.serotonin induced|Platelet aggregation.serotonin induced
C0365500|T201|COMP|6000-4|LNC|Platelet aggregation.thrombin induced|Platelet aggregation.thrombin induced
C0365516|T201|COMP|4678-9|LNC|Protein S|Protein S
C0365519|T201|COMP|5900-6|LNC|Prothrombin fragment 1+2|Prothrombin fragment 1+2
C0365524|T201|COMP|3290-4|LNC|2-Oxoisocaproate|2-Oxoisocaproate
C0365525|T201|COMP|3291-2|LNC|2-Pyridone|2-Pyridone
C0365526|T201|COMP|3292-0|LNC|2-Pyridone/N'-Methylnicotinamide|2-Pyridone/N'-Methylnicotinamide
C0365527|T201|COMP|3293-8|LNC|Acebutolol|Acebutolol
C0365528|T201|COMP|3294-6|LNC|Acebutolol|Acebutolol
C0365529|T201|COMP|3295-3|LNC|Acebutolol|Acebutolol
C0365530|T201|COMP|3296-1|LNC|Acepromazine|Acepromazine
C0365531|T201|COMP|3297-9|LNC|Acetaminophen|Acetaminophen
C0365532|T201|COMP|3298-7|LNC|Acetaminophen|Acetaminophen
C0365533|T201|COMP|3299-5|LNC|Acetaminophen|Acetaminophen
C0365534|T201|COMP|3300-1|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C0365535|T201|COMP|3301-9|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C0365536|T201|COMP|3302-7|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C0365537|T201|COMP|3303-5|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C0365538|T201|COMP|3304-3|LNC|Acetyldigitoxin|Acetyldigitoxin
C0365539|T201|COMP|3305-0|LNC|Acetylsalicylate|Acetylsalicylate
C0365540|T201|COMP|3306-8|LNC|Acetylsalicylate|Acetylsalicylate
C0365541|T201|COMP|3307-6|LNC|Alfentanil|Alfentanil
C0365542|T201|COMP|3308-4|LNC|Alphaprodine|Alphaprodine
C0365543|T201|COMP|3309-2|LNC|Alphaprodine|Alphaprodine
C0365544|T201|COMP|3310-0|LNC|Alphaprodine|Alphaprodine
C0365545|T201|COMP|3311-8|LNC|Alphaprodine|Alphaprodine
C0365547|T201|COMP|3313-4|LNC|ALPRAZolam|ALPRAZolam
C0365548|T201|COMP|3314-2|LNC|Alprenolol|Alprenolol
C0365549|T201|COMP|3315-9|LNC|Alprenolol|Alprenolol
C0365550|T201|COMP|3316-7|LNC|Alprenolol|Alprenolol
C0365551|T201|COMP|3317-5|LNC|Amantadine|Amantadine
C0365552|T201|COMP|3318-3|LNC|Amdinocillin|Amdinocillin
C0365553|T201|COMP|3319-1|LNC|Amikacin^peak|Amikacin^peak
C0365554|T201|COMP|3320-9|LNC|Amikacin^random|Amikacin^random
C0365555|T201|COMP|3321-7|LNC|Amikacin^trough|Amikacin^trough
C0365556|T201|COMP|3322-5|LNC|aMILoride|aMILoride
C0365557|T201|COMP|3323-3|LNC|aMILoride|aMILoride
C0365558|T201|COMP|3324-1|LNC|aMILoride|aMILoride
C0365559|T201|COMP|3325-8|LNC|aMILoride|aMILoride
C0365560|T201|COMP|3326-6|LNC|Aminocaproate^trough|Aminocaproate^trough
C0365562|T201|COMP|3328-2|LNC|Aminopyrine|Aminopyrine
C0365563|T201|COMP|3329-0|LNC|Aminosalicylate|Aminosalicylate
C0365564|T201|COMP|3330-8|LNC|Amiodarone|Amiodarone
C0365565|T201|COMP|3331-6|LNC|Amiodarone+Desethylamiodarone|Amiodarone+Desethylamiodarone
C0365566|T201|COMP|3332-4|LNC|Amitriptyline|Amitriptyline
C0365567|T201|COMP|3333-2|LNC|Amitriptyline|Amitriptyline
C0365568|T201|COMP|3334-0|LNC|Amitriptyline|Amitriptyline
C0365569|T201|COMP|3335-7|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C0365570|T201|COMP|3336-5|LNC|Amitriptyline^trough >12h post dose|Amitriptyline^trough >12h post dose
C0365571|T201|COMP|3337-3|LNC|Amobarbital|Amobarbital
C0365572|T201|COMP|3338-1|LNC|Amobarbital|Amobarbital
C0365573|T201|COMP|3339-9|LNC|Amobarbital|Amobarbital
C0365574|T201|COMP|3340-7|LNC|Amoxapine|Amoxapine
C0365575|T201|COMP|3341-5|LNC|Amoxapine|Amoxapine
C0365576|T201|COMP|3342-3|LNC|Amoxapine|Amoxapine
C0365577|T201|COMP|3343-1|LNC|Amoxapine|Amoxapine
C0365578|T201|COMP|3344-9|LNC|Amoxicillin|Amoxicillin
C0365579|T201|COMP|3345-6|LNC|Diethylpropion|Diethylpropion
C0365580|T201|COMP|3346-4|LNC|Diethylpropion|Diethylpropion
C0365581|T201|COMP|3347-2|LNC|Diethylpropion|Diethylpropion
C0365582|T201|COMP|3348-0|LNC|Amphetamines|Amphetamines
C0365583|T201|COMP|3349-8|LNC|Amphetamines|Amphetamines
C0365584|T201|COMP|3350-6|LNC|Amphetaminil|Amphetaminil
C0365585|T201|COMP|3351-4|LNC|Amphetaminil|Amphetaminil
C0365586|T201|COMP|3352-2|LNC|Amphetaminil|Amphetaminil
C0365587|T201|COMP|3353-0|LNC|Amphotericin B|Amphotericin B
C0365588|T201|COMP|3354-8|LNC|Amphotericin B|Amphotericin B
C0365589|T201|COMP|3355-5|LNC|Ampicillin|Ampicillin
C0365590|T201|COMP|3356-3|LNC|Anileridine|Anileridine
C0365591|T201|COMP|3357-1|LNC|Anileridine|Anileridine
C0365592|T201|COMP|3358-9|LNC|Anileridine|Anileridine
C0365593|T201|COMP|3359-7|LNC|Anileridine|Anileridine
C0365594|T201|COMP|3363-9|LNC|Anthraquinone|Anthraquinone
C0365595|T201|COMP|3364-7|LNC|Antipyrine|Antipyrine
C0365596|T201|COMP|3365-4|LNC|Antipyrine renal clearance|Antipyrine renal clearance
C0365597|T201|COMP|3366-2|LNC|Atenolol|Atenolol
C0365598|T201|COMP|3360-5|LNC|Atenolol|Atenolol
C0365599|T201|COMP|3361-3|LNC|Atenolol|Atenolol
C0365600|T201|COMP|3362-1|LNC|Atenolol|Atenolol
C0365601|T201|COMP|3367-0|LNC|Atropine|Atropine
C0365602|T201|COMP|3368-8|LNC|Azlocillin|Azlocillin
C0365603|T201|COMP|3369-6|LNC|Aztreonam|Aztreonam
C0365604|T201|COMP|3370-4|LNC|Barbital|Barbital
C0365605|T201|COMP|3371-2|LNC|Barbital|Barbital
C0365606|T201|COMP|3372-0|LNC|Barbiturate screen absent|Barbiturate screen absent
C0365607|T201|COMP|3374-6|LNC|Barbiturate screen present|Barbiturate screen present
C0365608|T201|COMP|3376-1|LNC|Barbiturates|Barbiturates
C0365609|T201|COMP|3377-9|LNC|Barbiturates|Barbiturates
C0365610|T201|COMP|3378-7|LNC|Bendroflumethiazide|Bendroflumethiazide
C0365611|T201|COMP|3379-5|LNC|Bendroflumethiazide|Bendroflumethiazide
C0365612|T201|COMP|3380-3|LNC|Bendroflumethiazide|Bendroflumethiazide
C0365613|T201|COMP|3381-1|LNC|Benzfetamine|Benzfetamine
C0365614|T201|COMP|3382-9|LNC|Benzfetamine|Benzfetamine
C0365615|T201|COMP|3383-7|LNC|Benzfetamine|Benzfetamine
C0365616|T201|COMP|3384-5|LNC|Benzfetamine|Benzfetamine
C0365617|T201|COMP|3385-2|LNC|Benzodiazepines negative|Benzodiazepines negative
C0365618|T201|COMP|3387-8|LNC|Benzodiazepines positive|Benzodiazepines positive
C0365619|T201|COMP|3389-4|LNC|Benzodiazepines|Benzodiazepines
C0365620|T201|COMP|3390-2|LNC|Benzodiazepines|Benzodiazepines
C0365621|T201|COMP|3391-0|LNC|Benzoylecgonine|Benzoylecgonine
C0365622|T201|COMP|3392-8|LNC|Benzoylecgonine|Benzoylecgonine
C0365627|T201|COMP|3397-7|LNC|Cocaine|Cocaine
C0365629|T201|COMP|3399-3|LNC|Benzthiazide|Benzthiazide
C0365630|T201|COMP|3400-9|LNC|Benzthiazide|Benzthiazide
C0365631|T201|COMP|3401-7|LNC|Benzthiazide|Benzthiazide
C0365632|T201|COMP|3402-5|LNC|Bolasterone|Bolasterone
C0365633|T201|COMP|3403-3|LNC|Bolasterone|Bolasterone
C0365634|T201|COMP|3404-1|LNC|Bolasterone|Bolasterone
C0365635|T201|COMP|3405-8|LNC|Bromazepam|Bromazepam
C0365636|T201|COMP|3406-6|LNC|Bromazepam|Bromazepam
C0365637|T201|COMP|3407-4|LNC|Brompheniramine|Brompheniramine
C0365638|T201|COMP|3408-2|LNC|Brompheniramine|Brompheniramine
C0365639|T201|COMP|3409-0|LNC|Bumetanide|Bumetanide
C0365640|T201|COMP|3410-8|LNC|Bumetanide|Bumetanide
C0365641|T201|COMP|3411-6|LNC|Bumetanide|Bumetanide
C0365642|T201|COMP|3412-4|LNC|Bupivacaine|Bupivacaine
C0365643|T201|COMP|3413-2|LNC|Buprenorphine|Buprenorphine
C0365644|T201|COMP|3414-0|LNC|Buprenorphine|Buprenorphine
C0365645|T201|COMP|3415-7|LNC|Buprenorphine|Buprenorphine
C0365646|T201|COMP|3416-5|LNC|Buprenorphine|Buprenorphine
C0365647|T201|COMP|3417-3|LNC|Butabarbital|Butabarbital
C0365648|T201|COMP|3418-1|LNC|Butabarbital|Butabarbital
C0365649|T201|COMP|3419-9|LNC|Butabarbital|Butabarbital
C0365650|T201|COMP|3420-7|LNC|Butalbital|Butalbital
C0365651|T201|COMP|3421-5|LNC|Butalbital|Butalbital
C0365652|T201|COMP|3422-3|LNC|Caffeine|Caffeine
C0365653|T201|COMP|3423-1|LNC|Caffeine|Caffeine
C0365654|T201|COMP|3424-9|LNC|Caffeine|Caffeine
C0365655|T201|COMP|3425-6|LNC|Cannabinoids|Cannabinoids
C0365656|T201|COMP|3426-4|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0365657|T201|COMP|3428-0|LNC|Canrenone|Canrenone
C0365658|T201|COMP|3429-8|LNC|Canrenone|Canrenone
C0365659|T201|COMP|3430-6|LNC|Canrenone|Canrenone
C0365660|T201|COMP|3431-4|LNC|carBAMazepine|carBAMazepine
C0365661|T201|COMP|3432-2|LNC|carBAMazepine|carBAMazepine
C0365662|T201|COMP|3433-0|LNC|carBAMazepine.free|carBAMazepine.free
C0365663|T201|COMP|3434-8|LNC|Carbenicillin|Carbenicillin
C0365664|T201|COMP|3435-5|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0365665|T201|COMP|3436-3|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0365666|T201|COMP|3437-1|LNC|Carisoprodol|Carisoprodol
C0365667|T201|COMP|3438-9|LNC|Cathine|Cathine
C0365668|T201|COMP|3439-7|LNC|Cathine|Cathine
C0365669|T201|COMP|3440-5|LNC|Cathine|Cathine
C0365670|T201|COMP|3441-3|LNC|Cefamandole|Cefamandole
C0365672|T201|COMP|3443-9|LNC|ceFAZolin|ceFAZolin
C0365673|T201|COMP|3444-7|LNC|Cefonicid|Cefonicid
C0365674|T201|COMP|3445-4|LNC|Cefoperazone|Cefoperazone
C0365675|T201|COMP|3446-2|LNC|Cefotaxime|Cefotaxime
C0365676|T201|COMP|3447-0|LNC|cefoTEtan|cefoTEtan
C0365677|T201|COMP|3448-8|LNC|cefOXitin|cefOXitin
C0365678|T201|COMP|3449-6|LNC|cefTAZidime|cefTAZidime
C0365679|T201|COMP|3450-4|LNC|Ceftizoxime|Ceftizoxime
C0365680|T201|COMP|3451-2|LNC|cefTRIAXone|cefTRIAXone
C0365681|T201|COMP|3452-0|LNC|Cefuroxime.parenteral|Cefuroxime.parenteral
C0365682|T201|COMP|3453-8|LNC|Cephalexin|Cephalexin
C0365683|T201|COMP|3454-6|LNC|Cephalothin|Cephalothin
C0365684|T201|COMP|3455-3|LNC|Chloramphenicol|Chloramphenicol
C0365685|T201|COMP|3456-1|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0365686|T201|COMP|3457-9|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0365687|T201|COMP|3458-7|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0365688|T201|COMP|3459-5|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0365689|T201|COMP|3460-3|LNC|Chlormerodrin|Chlormerodrin
C0365690|T201|COMP|3461-1|LNC|Chlormerodrin|Chlormerodrin
C0365691|T201|COMP|3462-9|LNC|Chlormerodrin|Chlormerodrin
C0365692|T201|COMP|3463-7|LNC|Chloroquine|Chloroquine
C0365693|T201|COMP|3464-5|LNC|Chlorothiazide|Chlorothiazide
C0365694|T201|COMP|3465-2|LNC|Chlorpheniramine|Chlorpheniramine
C0365695|T201|COMP|3466-0|LNC|Chlorpheniramine|Chlorpheniramine
C0365696|T201|COMP|3467-8|LNC|Chlorpheniramine|Chlorpheniramine
C0365697|T201|COMP|3468-6|LNC|Chlorphentermine|Chlorphentermine
C0365698|T201|COMP|3469-4|LNC|Chlorphentermine|Chlorphentermine
C0365699|T201|COMP|3470-2|LNC|Chlorphentermine|Chlorphentermine
C0365700|T201|COMP|3471-0|LNC|chlorproMAZINE|chlorproMAZINE
C0365701|T201|COMP|3472-8|LNC|chlorproMAZINE|chlorproMAZINE
C0365702|T201|COMP|3473-6|LNC|chlorproMAZINE|chlorproMAZINE
C0365703|T201|COMP|3474-4|LNC|chlorproPAMIDE|chlorproPAMIDE
C0365704|T201|COMP|3475-1|LNC|Chlorprothixene|Chlorprothixene
C0365705|T201|COMP|3476-9|LNC|Chlorprothixene|Chlorprothixene
C0365706|T201|COMP|3477-7|LNC|Chlorprothixene|Chlorprothixene
C0365707|T201|COMP|3478-5|LNC|Chlorthalidone|Chlorthalidone
C0365708|T201|COMP|3479-3|LNC|Chlorthalidone|Chlorthalidone
C0365709|T201|COMP|3480-1|LNC|Chlorthalidone|Chlorthalidone
C0365710|T201|COMP|3481-9|LNC|Cimetidine|Cimetidine
C0365711|T201|COMP|3482-7|LNC|Cimetidine|Cimetidine
C0365712|T201|COMP|3483-5|LNC|Cimetidine|Cimetidine
C0365713|T201|COMP|3484-3|LNC|Ciprofloxacin|Ciprofloxacin
C0365714|T201|COMP|3485-0|LNC|CISplatin|CISplatin
C0365715|T201|COMP|3486-8|LNC|Clindamycin|Clindamycin
C0365716|T201|COMP|3487-6|LNC|cloBAZam|cloBAZam
C0365717|T201|COMP|3488-4|LNC|Clobenzorex|Clobenzorex
C0365718|T201|COMP|3489-2|LNC|Clobenzorex|Clobenzorex
C0365719|T201|COMP|3490-0|LNC|Clofibrate|Clofibrate
C0365720|T201|COMP|3491-8|LNC|clomiPRAMINE|clomiPRAMINE
C0365721|T201|COMP|3492-6|LNC|clomiPRAMINE|clomiPRAMINE
C0365722|T201|COMP|3493-4|LNC|Clomipramine+Norclomipramine|Clomipramine+Norclomipramine
C0365723|T201|COMP|3494-2|LNC|clonazePAM|clonazePAM
C0365724|T201|COMP|3495-9|LNC|cloNIDine|cloNIDine
C0365725|T201|COMP|3496-7|LNC|Clopenthixol|Clopenthixol
C0365726|T201|COMP|3497-5|LNC|Clopenthixol|Clopenthixol
C0365727|T201|COMP|3498-3|LNC|Clorazepate|Clorazepate
C0365728|T201|COMP|3499-1|LNC|Clorprenaline|Clorprenaline
C0365729|T201|COMP|3500-6|LNC|Clorprenaline|Clorprenaline
C0365730|T201|COMP|3501-4|LNC|Clorprenaline|Clorprenaline
C0365731|T201|COMP|3502-2|LNC|Clostebol|Clostebol
C0365732|T201|COMP|3503-0|LNC|Clostebol|Clostebol
C0365733|T201|COMP|3504-8|LNC|Clostebol|Clostebol
C0365734|T201|COMP|3505-5|LNC|Codeine|Codeine
C0365735|T201|COMP|3506-3|LNC|Codeine|Codeine
C0365736|T201|COMP|3507-1|LNC|Codeine|Codeine
C0365738|T201|COMP|3509-7|LNC|Prochlorperazine|Prochlorperazine
C0365739|T201|COMP|3510-5|LNC|Prochlorperazine|Prochlorperazine
C0365740|T201|COMP|3511-3|LNC|Cropropamide|Cropropamide
C0365741|T201|COMP|3512-1|LNC|Cropropamide|Cropropamide
C0365742|T201|COMP|3513-9|LNC|Cropropamide|Cropropamide
C0365743|T201|COMP|3514-7|LNC|Crotetamide|Crotetamide
C0365744|T201|COMP|3515-4|LNC|Crotetamide|Crotetamide
C0365745|T201|COMP|3516-2|LNC|Crotetamide|Crotetamide
C0365746|T201|COMP|3517-0|LNC|Cyclacillin|Cyclacillin
C0365747|T201|COMP|3518-8|LNC|Cyclizine|Cyclizine
C0365748|T201|COMP|3519-6|LNC|cycloSERINE|cycloSERINE
C0365749|T201|COMP|3520-4|LNC|cycloSPORINE|cycloSPORINE
C0365750|T201|COMP|3521-2|LNC|cycloSPORINE|cycloSPORINE
C0365751|T201|COMP|3522-0|LNC|cycloSPORINE+Metabolites|cycloSPORINE+Metabolites
C0365752|T201|COMP|3523-8|LNC|cycloSPORINE^12H post dose|cycloSPORINE^12H post dose
C0365753|T201|COMP|3524-6|LNC|cycloSPORINE^12H post dose|cycloSPORINE^12H post dose
C0365754|T201|COMP|3525-3|LNC|cycloSPORINE^24H post dose|cycloSPORINE^24H post dose
C0365755|T201|COMP|3526-1|LNC|cycloSPORINE^24H post dose|cycloSPORINE^24H post dose
C0365756|T201|COMP|3527-9|LNC|Dantron|Dantron
C0365757|T201|COMP|3528-7|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0365758|T201|COMP|3529-5|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0365759|T201|COMP|3530-3|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0365760|T201|COMP|3531-1|LNC|Desipramine|Desipramine
C0365761|T201|COMP|3532-9|LNC|Desipramine|Desipramine
C0365762|T201|COMP|3533-7|LNC|Desipramine|Desipramine
C0365763|T201|COMP|3534-5|LNC|Desipramine|Desipramine
C0365764|T201|COMP|3535-2|LNC|Desipramine^trough|Desipramine^trough
C0365766|T201|COMP|3537-8|LNC|Nordiazepam|Nordiazepam
C0365767|T201|COMP|3538-6|LNC|Dextromethorphan|Dextromethorphan
C0365768|T201|COMP|3539-4|LNC|Dextromethorphan|Dextromethorphan
C0365769|T201|COMP|3540-2|LNC|Dextromoramide|Dextromoramide
C0365770|T201|COMP|3541-0|LNC|Dextromoramide|Dextromoramide
C0365771|T201|COMP|3542-8|LNC|Propoxyphene|Propoxyphene
C0365772|T201|COMP|3543-6|LNC|Propoxyphene|Propoxyphene
C0365773|T201|COMP|19141-1|LNC|Propoxyphene|Propoxyphene
C0365774|T201|COMP|3545-1|LNC|Propoxyphene|Propoxyphene
C0365775|T201|COMP|3546-9|LNC|Diamorphine|Diamorphine
C0365776|T201|COMP|3547-7|LNC|Diamorphine|Diamorphine
C0365777|T201|COMP|3548-5|LNC|diazePAM|diazePAM
C0365778|T201|COMP|3549-3|LNC|diazePAM|diazePAM
C0365779|T201|COMP|3550-1|LNC|diazePAM|diazePAM
C0365780|T201|COMP|3551-9|LNC|diazePAM|diazePAM
C0365781|T201|COMP|3552-7|LNC|diazePAM^trough|diazePAM^trough
C0365782|T201|COMP|3553-5|LNC|Dibenzepin|Dibenzepin
C0365783|T201|COMP|3554-3|LNC|Dibucaine number|Dibucaine number
C0365784|T201|COMP|3555-0|LNC|Dichlorphenamide|Dichlorphenamide
C0365785|T201|COMP|3556-8|LNC|Dichlorphenamide|Dichlorphenamide
C0365786|T201|COMP|3557-6|LNC|Dichlorphenamide|Dichlorphenamide
C0365787|T201|COMP|3558-4|LNC|Dicoumarol|Dicoumarol
C0365788|T201|COMP|3559-2|LNC|Digitoxin|Digitoxin
C0365789|T201|COMP|3560-0|LNC|Digitoxin|Digitoxin
C0365790|T201|COMP|3561-8|LNC|Digitoxin>6H post dose|Digitoxin>6H post dose
C0365791|T201|COMP|3562-6|LNC|Digoxin.free|Digoxin.free
C0365792|T201|COMP|3563-4|LNC|Digoxin>12H post dose|Digoxin>12H post dose
C0365793|T201|COMP|3564-2|LNC|Dimetamphetamine|Dimetamphetamine
C0365794|T201|COMP|3565-9|LNC|Dimetamphetamine|Dimetamphetamine
C0365795|T201|COMP|3566-7|LNC|Dimetamphetamine|Dimetamphetamine
C0365796|T201|COMP|3567-5|LNC|Dimethyltryptamine|Dimethyltryptamine
C0365797|T201|COMP|3568-3|LNC|Dimethyltryptamine|Dimethyltryptamine
C0365798|T201|COMP|3569-1|LNC|diphenhydrAMINE|diphenhydrAMINE
C0365799|T201|COMP|3570-9|LNC|diphenhydrAMINE|diphenhydrAMINE
C0365800|T201|COMP|3571-7|LNC|diphenhydrAMINE|diphenhydrAMINE
C0365801|T201|COMP|3572-5|LNC|diphenhydrAMINE|diphenhydrAMINE
C0365802|T201|COMP|3573-3|LNC|Dipipanone|Dipipanone
C0365803|T201|COMP|3574-1|LNC|Dipipanone|Dipipanone
C0365804|T201|COMP|3575-8|LNC|Dipipanone|Dipipanone
C0365805|T201|COMP|3576-6|LNC|Disopyramide|Disopyramide
C0365806|T201|COMP|3577-4|LNC|Disulfiram|Disulfiram
C0365807|T201|COMP|3578-2|LNC|Doxepin|Doxepin
C0365808|T201|COMP|3579-0|LNC|Doxepin|Doxepin
C0365809|T201|COMP|3580-8|LNC|Doxepin|Doxepin
C0365810|T201|COMP|3581-6|LNC|Doxepin|Doxepin
C0365811|T201|COMP|3582-4|LNC|Doxepin+Nordoxepin|Doxepin+Nordoxepin
C0365812|T201|COMP|3583-2|LNC|Doxepin+Metabolites|Doxepin+Metabolites
C0365813|T201|COMP|3584-0|LNC|Doxepin^trough|Doxepin^trough
C0365814|T201|COMP|3585-7|LNC|Doxylamine|Doxylamine
C0365815|T201|COMP|3586-5|LNC|Doxylamine|Doxylamine
C0365816|T201|COMP|3587-3|LNC|Dyphylline|Dyphylline
C0365817|T201|COMP|3588-1|LNC|Emetine|Emetine
C0365818|T201|COMP|3589-9|LNC|Encainide|Encainide
C0365819|T201|COMP|3590-7|LNC|Enoxacin|Enoxacin
C0365820|T201|COMP|3591-5|LNC|ePHEDrine|ePHEDrine
C0365821|T201|COMP|3592-3|LNC|ePHEDrine|ePHEDrine
C0365822|T201|COMP|3593-1|LNC|ePHEDrine|ePHEDrine
C0365823|T201|COMP|3594-9|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C0365824|T201|COMP|3595-6|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C0365825|T201|COMP|3596-4|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C0365826|T201|COMP|3597-2|LNC|Erythromycin|Erythromycin
C0365827|T201|COMP|3598-0|LNC|Estazolam|Estazolam
C0365828|T201|COMP|3599-8|LNC|Etafedrine|Etafedrine
C0365829|T201|COMP|3600-4|LNC|Etafedrine|Etafedrine
C0365830|T201|COMP|3601-2|LNC|Etafedrine|Etafedrine
C0365831|T201|COMP|3602-0|LNC|Etamivan|Etamivan
C0365832|T201|COMP|3603-8|LNC|Etamivan|Etamivan
C0365833|T201|COMP|3604-6|LNC|Etamivan|Etamivan
C0365834|T201|COMP|3605-3|LNC|Ethacrynate|Ethacrynate
C0365835|T201|COMP|3606-1|LNC|Ethacrynate|Ethacrynate
C0365836|T201|COMP|3607-9|LNC|Ethambutol|Ethambutol
C0365837|T201|COMP|3608-7|LNC|Ethchlorvynol|Ethchlorvynol
C0365838|T201|COMP|3609-5|LNC|Ethchlorvynol|Ethchlorvynol
C0365839|T201|COMP|3610-3|LNC|Ethchlorvynol|Ethchlorvynol
C0365840|T201|COMP|3611-1|LNC|Ethchlorvynol|Ethchlorvynol
C0365841|T201|COMP|3612-9|LNC|Ethchlorvynol|Ethchlorvynol
C0365842|T201|COMP|3613-7|LNC|Ethoheptazine|Ethoheptazine
C0365843|T201|COMP|3614-5|LNC|Ethoheptazine|Ethoheptazine
C0365844|T201|COMP|3615-2|LNC|Ethoheptazine|Ethoheptazine
C0365845|T201|COMP|3616-0|LNC|Ethosuximide|Ethosuximide
C0365846|T201|COMP|3617-8|LNC|Ethotoin|Ethotoin
C0365847|T201|COMP|3618-6|LNC|Ethylmorphine|Ethylmorphine
C0365848|T201|COMP|3619-4|LNC|Ethylmorphine|Ethylmorphine
C0365850|T201|COMP|3621-0|LNC|Etilefrine|Etilefrine
C0365851|T201|COMP|3622-8|LNC|Etilefrine|Etilefrine
C0365852|T201|COMP|3623-6|LNC|Etilefrine|Etilefrine
C0365853|T201|COMP|3624-4|LNC|Fencamfamin|Fencamfamin
C0365854|T201|COMP|3625-1|LNC|Fencamfamin|Fencamfamin
C0365855|T201|COMP|3626-9|LNC|Fencamfamin|Fencamfamin
C0365856|T201|COMP|3627-7|LNC|Fenetylline|Fenetylline
C0365857|T201|COMP|3628-5|LNC|Fenetylline|Fenetylline
C0365858|T201|COMP|3629-3|LNC|Fenetylline|Fenetylline
C0365859|T201|COMP|3630-1|LNC|Fenfluramine|Fenfluramine
C0365860|T201|COMP|3631-9|LNC|Fenfluramine|Fenfluramine
C0365861|T201|COMP|3632-7|LNC|Fenoprofen|Fenoprofen
C0365862|T201|COMP|3633-5|LNC|Fenproporex|Fenproporex
C0365863|T201|COMP|3634-3|LNC|Fenproporex|Fenproporex
C0365864|T201|COMP|3635-0|LNC|Fenproporex|Fenproporex
C0365865|T201|COMP|3636-8|LNC|fentaNYL|fentaNYL
C0365866|T201|COMP|3637-6|LNC|fentaNYL|fentaNYL
C0365867|T201|COMP|3638-4|LNC|Flecainide|Flecainide
C0365868|T201|COMP|3639-2|LNC|5-Fluorocytosine|5-Fluorocytosine
C0365869|T201|COMP|3640-0|LNC|Flunitrazepam|Flunitrazepam
C0365870|T201|COMP|3641-8|LNC|Flunitrazepam|Flunitrazepam
C0365871|T201|COMP|3642-6|LNC|Fluorouracil|Fluorouracil
C0365872|T201|COMP|3643-4|LNC|FLUoxetine|FLUoxetine
C0365873|T201|COMP|3644-2|LNC|FLUoxetine|FLUoxetine
C0365874|T201|COMP|3645-9|LNC|FLUoxetine|FLUoxetine
C0365875|T201|COMP|3646-7|LNC|Fluoxymesterone|Fluoxymesterone
C0365876|T201|COMP|3647-5|LNC|Fluoxymesterone|Fluoxymesterone
C0365877|T201|COMP|3648-3|LNC|Fluoxymesterone|Fluoxymesterone
C0365878|T201|COMP|3649-1|LNC|Flupenthixol|Flupenthixol
C0365879|T201|COMP|3650-9|LNC|fluPHENAZine|fluPHENAZine
C0365880|T201|COMP|3651-7|LNC|fluPHENAZine|fluPHENAZine
C0365881|T201|COMP|3652-5|LNC|Flurazepam|Flurazepam
C0365882|T201|COMP|3653-3|LNC|Flurazepam|Flurazepam
C0365883|T201|COMP|3654-1|LNC|Flurazepam|Flurazepam
C0365884|T201|COMP|3655-8|LNC|Flurazepam|Flurazepam
C0365885|T201|COMP|3656-6|LNC|Furfenorex|Furfenorex
C0365886|T201|COMP|3657-4|LNC|Furfenorex|Furfenorex
C0365887|T201|COMP|3658-2|LNC|Furfenorex|Furfenorex
C0365888|T201|COMP|3659-0|LNC|Furosemide|Furosemide
C0365889|T201|COMP|3660-8|LNC|Furosemide|Furosemide
C0365890|T201|COMP|3661-6|LNC|Furosemide|Furosemide
C0365891|T201|COMP|3662-4|LNC|Furosemide|Furosemide
C0365892|T201|COMP|3663-2|LNC|Gentamicin^peak|Gentamicin^peak
C0365893|T201|COMP|3664-0|LNC|Gentamicin^random|Gentamicin^random
C0365894|T201|COMP|3665-7|LNC|Gentamicin^trough|Gentamicin^trough
C0365895|T201|COMP|3666-5|LNC|Glutethimide|Glutethimide
C0365896|T201|COMP|3667-3|LNC|Glutethimide|Glutethimide
C0365897|T201|COMP|3668-1|LNC|Glutethimide|Glutethimide
C0365898|T201|COMP|3669-9|LNC|Haloperidol|Haloperidol
C0365899|T201|COMP|3670-7|LNC|Haloperidol|Haloperidol
C0365900|T201|COMP|3671-5|LNC|Haloperidol|Haloperidol
C0365901|T201|COMP|3672-3|LNC|Heptaminol|Heptaminol
C0365902|T201|COMP|3673-1|LNC|Heptaminol|Heptaminol
C0365903|T201|COMP|3674-9|LNC|Heptaminol|Heptaminol
C0365904|T201|COMP|3675-6|LNC|hydroCHLOROthiazide|hydroCHLOROthiazide
C0365905|T201|COMP|3676-4|LNC|hydroCHLOROthiazide|hydroCHLOROthiazide
C0365906|T201|COMP|3677-2|LNC|hydroCHLOROthiazide|hydroCHLOROthiazide
C0365907|T201|COMP|3678-0|LNC|hydroCHLOROthiazide|hydroCHLOROthiazide
C0365908|T201|COMP|3679-8|LNC|HYDROcodone|HYDROcodone
C0365909|T201|COMP|3680-6|LNC|HYDROcodone|HYDROcodone
C0365910|T201|COMP|3681-4|LNC|HYDROcodone|HYDROcodone
C0365911|T201|COMP|3682-2|LNC|HYDROmorphone|HYDROmorphone
C0365912|T201|COMP|3683-0|LNC|HYDROmorphone|HYDROmorphone
C0365913|T201|COMP|3684-8|LNC|Hydroxychloroquine|Hydroxychloroquine
C0365914|T201|COMP|3685-5|LNC|Hydroxymethoxyphenamine|Hydroxymethoxyphenamine
C0365915|T201|COMP|3686-3|LNC|hydrOXYzine|hydrOXYzine
C0365916|T201|COMP|3687-1|LNC|Ibuprofen|Ibuprofen
C0365917|T201|COMP|3688-9|LNC|Imipenem+Cilastatin|Imipenem+Cilastatin
C0365918|T201|COMP|3689-7|LNC|Imipramine|Imipramine
C0365919|T201|COMP|3690-5|LNC|Imipramine|Imipramine
C0365920|T201|COMP|3691-3|LNC|Imipramine|Imipramine
C0365921|T201|COMP|3692-1|LNC|Imipramine|Imipramine
C0365922|T201|COMP|3693-9|LNC|Imipramine^trough|Imipramine^trough
C0365923|T201|COMP|3694-7|LNC|Indomethacin|Indomethacin
C0365924|T201|COMP|3696-2|LNC|Insulin renal clearance|Insulin renal clearance
C0365925|T201|COMP|3695-4|LNC|Insulin|Insulin
C0365926|T201|COMP|3697-0|LNC|Isoniazid|Isoniazid
C0365927|T201|COMP|3698-8|LNC|Kanamycin^peak|Kanamycin^peak
C0365928|T201|COMP|3699-6|LNC|Kanamycin^random|Kanamycin^random
C0365929|T201|COMP|3700-2|LNC|Kanamycin^trough|Kanamycin^trough
C0365930|T201|COMP|3701-0|LNC|Ketamine|Ketamine
C0365931|T201|COMP|3702-8|LNC|Ketobemidone|Ketobemidone
C0365932|T201|COMP|3703-6|LNC|Ketobemidone|Ketobemidone
C0365933|T201|COMP|3704-4|LNC|Labetalol|Labetalol
C0365934|T201|COMP|3705-1|LNC|Labetalol|Labetalol
C0365935|T201|COMP|3706-9|LNC|Labetalol|Labetalol
C0365936|T201|COMP|3707-7|LNC|Labetalol|Labetalol
C0365937|T201|COMP|3708-5|LNC|Methotrimeprazine|Methotrimeprazine
C0365938|T201|COMP|3709-3|LNC|Levomepromazine|Levomepromazine
C0365939|T201|COMP|3710-1|LNC|Levorphanol|Levorphanol
C0365940|T201|COMP|3711-9|LNC|Levorphanol|Levorphanol
C0365941|T201|COMP|3712-7|LNC|Levorphanol|Levorphanol
C0365942|T201|COMP|3713-5|LNC|Levorphanol|Levorphanol
C0365943|T201|COMP|3714-3|LNC|Lidocaine|Lidocaine
C0365944|T201|COMP|3715-0|LNC|Lidocaine|Lidocaine
C0365945|T201|COMP|3716-8|LNC|Lidocaine|Lidocaine
C0365946|T201|COMP|3717-6|LNC|Lidocaine^>45m post bolus dose|Lidocaine^>45m post bolus dose
C0365947|T201|COMP|3718-4|LNC|Lithium|Lithium
C0365948|T201|COMP|3719-2|LNC|Lithium|Lithium
C0365949|T201|COMP|3720-0|LNC|Lithium|Lithium
C0365950|T201|COMP|3721-8|LNC|Lithium|Lithium
C0365951|T201|COMP|3722-6|LNC|Lithium renal clearance|Lithium renal clearance
C0365952|T201|COMP|3723-4|LNC|Lithium^trough|Lithium^trough
C0365953|T201|COMP|3724-2|LNC|LORazepam|LORazepam
C0365954|T201|COMP|3725-9|LNC|LORazepam|LORazepam
C0365955|T201|COMP|3726-7|LNC|Lormetazepam|Lormetazepam
C0365956|T201|COMP|3727-5|LNC|Loxapine|Loxapine
C0365957|T201|COMP|3728-3|LNC|Loxapine|Loxapine
C0365958|T201|COMP|3729-1|LNC|Loxapine|Loxapine
C0365959|T201|COMP|3730-9|LNC|Lysergate diethylamide|Lysergate diethylamide
C0365960|T201|COMP|3731-7|LNC|Lysergate diethylamide|Lysergate diethylamide
C0365961|T201|COMP|3732-5|LNC|Lysergate diethylamide|Lysergate diethylamide
C0365962|T201|COMP|5679-6|LNC|Lysergate diethylamide|Lysergate diethylamide
C0365963|T201|COMP|3734-1|LNC|Maprotiline|Maprotiline
C0365964|T201|COMP|3735-8|LNC|Maprotiline|Maprotiline
C0365965|T201|COMP|3737-4|LNC|Maprotiline|Maprotiline
C0365966|T201|COMP|3738-2|LNC|Maprotiline|Maprotiline
C0365967|T201|COMP|3739-0|LNC|Medazepam|Medazepam
C0365968|T201|COMP|3740-8|LNC|Medazepam|Medazepam
C0365969|T201|COMP|3741-6|LNC|Mefenorex|Mefenorex
C0365970|T201|COMP|3742-4|LNC|Mefenorex|Mefenorex
C0365971|T201|COMP|3743-2|LNC|Mefenorex|Mefenorex
C0365972|T201|COMP|3744-0|LNC|Meperidine|Meperidine
C0365973|T201|COMP|3745-7|LNC|Meperidine|Meperidine
C0365974|T201|COMP|3746-5|LNC|Meperidine|Meperidine
C0365975|T201|COMP|3747-3|LNC|Meperidine|Meperidine
C0365976|T201|COMP|3748-1|LNC|Meperidine|Meperidine
C0365977|T201|COMP|3749-9|LNC|Mephenytoin|Mephenytoin
C0365978|T201|COMP|3750-7|LNC|Mephobarbital|Mephobarbital
C0365979|T201|COMP|3752-3|LNC|Meprobamate|Meprobamate
C0365980|T201|COMP|3753-1|LNC|Meprobamate|Meprobamate
C0365981|T201|COMP|3754-9|LNC|Meprobamate|Meprobamate
C0365982|T201|COMP|3755-6|LNC|Meprobamate|Meprobamate
C0365983|T201|COMP|3756-4|LNC|Mersalyl|Mersalyl
C0365984|T201|COMP|3757-2|LNC|Mersalyl|Mersalyl
C0365985|T201|COMP|3758-0|LNC|Mersalyl|Mersalyl
C0365986|T201|COMP|3759-8|LNC|Mesantoin|Mesantoin
C0365988|T201|COMP|3761-4|LNC|Mesterolone|Mesterolone
C0365989|T201|COMP|3762-2|LNC|Mesterolone|Mesterolone
C0365990|T201|COMP|3763-0|LNC|Mesterolone|Mesterolone
C0365991|T201|COMP|3764-8|LNC|Metandienone|Metandienone
C0365992|T201|COMP|3765-5|LNC|Metandienone|Metandienone
C0365993|T201|COMP|3766-3|LNC|Metandienone|Metandienone
C0365994|T201|COMP|3767-1|LNC|Metaraminol|Metaraminol
C0365995|T201|COMP|3768-9|LNC|Metenolone|Metenolone
C0365996|T201|COMP|3769-7|LNC|Metenolone|Metenolone
C0365997|T201|COMP|3770-5|LNC|Metenolone|Metenolone
C0365998|T201|COMP|3771-3|LNC|Methadone|Methadone
C0365999|T201|COMP|3772-1|LNC|Methadone|Methadone
C0366000|T201|COMP|3773-9|LNC|Methadone|Methadone
C0366001|T201|COMP|3774-7|LNC|Methadone|Methadone
C0366002|T201|COMP|3775-4|LNC|Methadone|Methadone
C0366003|T201|COMP|3776-2|LNC|Methamphetamine|Methamphetamine
C0366004|T201|COMP|3777-0|LNC|Methamphetamine|Methamphetamine
C0366005|T201|COMP|3778-8|LNC|Methamphetamine|Methamphetamine
C0366006|T201|COMP|3779-6|LNC|Methamphetamine|Methamphetamine
C0366007|T201|COMP|3780-4|LNC|Methamphetamine|Methamphetamine
C0366008|T201|COMP|3781-2|LNC|Methapyrilene|Methapyrilene
C0366009|T201|COMP|3782-0|LNC|Methapyrilene|Methapyrilene
C0366010|T201|COMP|3783-8|LNC|Methapyrilene|Methapyrilene
C0366011|T201|COMP|3784-6|LNC|Methaqualone|Methaqualone
C0366012|T201|COMP|3785-3|LNC|Methaqualone|Methaqualone
C0366013|T201|COMP|3786-1|LNC|Methaqualone|Methaqualone
C0366014|T201|COMP|3787-9|LNC|Methaqualone|Methaqualone
C0366015|T201|COMP|3788-7|LNC|Methicillin|Methicillin
C0366016|T201|COMP|3789-5|LNC|Methocarbamol|Methocarbamol
C0366017|T201|COMP|3790-3|LNC|Methocarbamol|Methocarbamol
C0366018|T201|COMP|3791-1|LNC|Methocarbamol|Methocarbamol
C0366019|T201|COMP|3792-9|LNC|Methotrexate|Methotrexate
C0366020|T201|COMP|3793-7|LNC|Methotrexate|Methotrexate
C0366021|T201|COMP|3794-5|LNC|Methotrexate^1-2w post dose|Methotrexate^1-2w post dose
C0366022|T201|COMP|3795-2|LNC|Methotrexate^24H post dose|Methotrexate^24H post dose
C0366023|T201|COMP|3796-0|LNC|Methotrexate^48H post dose|Methotrexate^48H post dose
C0366024|T201|COMP|3797-8|LNC|Methotrexate^72H post dose|Methotrexate^72H post dose
C0366025|T201|COMP|3798-6|LNC|Methoxyphenamine|Methoxyphenamine
C0366026|T201|COMP|3799-4|LNC|Methoxyphenamine|Methoxyphenamine
C0366027|T201|COMP|3800-0|LNC|Methoxyphenamine|Methoxyphenamine
C0366028|T201|COMP|3801-8|LNC|Methsuximide|Methsuximide
C0366029|T201|COMP|3802-6|LNC|Methyldopa|Methyldopa
C0366030|T201|COMP|3803-4|LNC|MethylePHEDrine|MethylePHEDrine
C0366031|T201|COMP|3804-2|LNC|MethylePHEDrine|MethylePHEDrine
C0366032|T201|COMP|3805-9|LNC|MethylePHEDrine|MethylePHEDrine
C0366033|T201|COMP|3806-7|LNC|Methylphenidate|Methylphenidate
C0366034|T201|COMP|3807-5|LNC|Methylphenidate|Methylphenidate
C0366035|T201|COMP|3808-3|LNC|Methylphenidate|Methylphenidate
C0366036|T201|COMP|3809-1|LNC|Methylphenidate|Methylphenidate
C0366037|T201|COMP|3810-9|LNC|Methylphenidate|Methylphenidate
C0366038|T201|COMP|3811-7|LNC|Methyprylon|Methyprylon
C0366039|T201|COMP|3812-5|LNC|Methyprylon|Methyprylon
C0366040|T201|COMP|3813-3|LNC|Methyprylon|Methyprylon
C0366041|T201|COMP|3814-1|LNC|Methyprylon|Methyprylon
C0366042|T201|COMP|3815-8|LNC|Metoprolol|Metoprolol
C0366043|T201|COMP|3816-6|LNC|Metoprolol|Metoprolol
C0366044|T201|COMP|3817-4|LNC|Metoprolol|Metoprolol
C0366045|T201|COMP|3818-2|LNC|Metoprolol|Metoprolol
C0366046|T201|COMP|3819-0|LNC|Mexiletine|Mexiletine
C0366047|T201|COMP|3820-8|LNC|Mezlocillin|Mezlocillin
C0366048|T201|COMP|3821-6|LNC|Midazolam|Midazolam
C0366049|T201|COMP|3822-4|LNC|Minocycline|Minocycline
C0366050|T201|COMP|3823-2|LNC|Morazone|Morazone
C0366051|T201|COMP|3824-0|LNC|Morazone|Morazone
C0366052|T201|COMP|3825-7|LNC|Morazone|Morazone
C0366053|T201|COMP|3826-5|LNC|Morphine|Morphine
C0366054|T201|COMP|3827-3|LNC|Morphine|Morphine
C0366055|T201|COMP|3828-1|LNC|Morphine.free|Morphine.free
C0366056|T201|COMP|3829-9|LNC|Morphine.free|Morphine.free
C0366057|T201|COMP|3830-7|LNC|Morphine|Morphine
C0366058|T201|COMP|3831-5|LNC|Morphine|Morphine
C0366059|T201|COMP|3832-3|LNC|Morphine|Morphine
C0366060|T201|COMP|3833-1|LNC|Moxalactam|Moxalactam
C0366061|T201|COMP|3834-9|LNC|N-acetylprocainamide|N-acetylprocainamide
C0366062|T201|COMP|3620-2|LNC|N-ethylnicotinamide|N-ethylnicotinamide
C0366063|T201|COMP|3836-4|LNC|Nadolol|Nadolol
C0366064|T201|COMP|3837-2|LNC|Nadolol|Nadolol
C0366065|T201|COMP|3838-0|LNC|Nadolol|Nadolol
C0366066|T201|COMP|3839-8|LNC|Nalbuphine|Nalbuphine
C0366067|T201|COMP|3840-6|LNC|Nalbuphine|Nalbuphine
C0366068|T201|COMP|3841-4|LNC|Nalbuphine|Nalbuphine
C0366069|T201|COMP|3842-2|LNC|Nalorphine|Nalorphine
C0366070|T201|COMP|3843-0|LNC|Nandrolone|Nandrolone
C0366071|T201|COMP|3844-8|LNC|Nandrolone|Nandrolone
C0366072|T201|COMP|3845-5|LNC|Nandrolone|Nandrolone
C0366073|T201|COMP|3846-3|LNC|Naproxen|Naproxen
C0366074|T201|COMP|3847-1|LNC|Neopterin|Neopterin
C0366075|T201|COMP|3848-9|LNC|Netilmicin^peak|Netilmicin^peak
C0366076|T201|COMP|3849-7|LNC|Netilmicin^random|Netilmicin^random
C0366077|T201|COMP|3850-5|LNC|Netilmicin^trough|Netilmicin^trough
C0366078|T201|COMP|3851-3|LNC|Nicomorphine|Nicomorphine
C0366079|T201|COMP|3852-1|LNC|Nicotinamide|Nicotinamide
C0366080|T201|COMP|3853-9|LNC|Nicotine|Nicotine
C0366081|T201|COMP|3854-7|LNC|Nicotine|Nicotine
C0366082|T201|COMP|3855-4|LNC|Nikethamide|Nikethamide
C0366083|T201|COMP|3856-2|LNC|Nikethamide|Nikethamide
C0366084|T201|COMP|3857-0|LNC|Nikethamide|Nikethamide
C0366085|T201|COMP|3858-8|LNC|Nitrazepam|Nitrazepam
C0366086|T201|COMP|3859-6|LNC|Nitrazepam|Nitrazepam
C0366087|T201|COMP|3860-4|LNC|Nitrofurantoin|Nitrofurantoin
C0366088|T201|COMP|3861-2|LNC|Nordiazepam|Nordiazepam
C0366089|T201|COMP|3862-0|LNC|Nordoxepin|Nordoxepin
C0366090|T201|COMP|3863-8|LNC|Norethandrolone|Norethandrolone
C0366091|T201|COMP|3864-6|LNC|Norethandrolone|Norethandrolone
C0366092|T201|COMP|3865-3|LNC|Norethandrolone|Norethandrolone
C0366093|T201|COMP|3866-1|LNC|Norfenefrine|Norfenefrine
C0366094|T201|COMP|3867-9|LNC|Norfloxacin|Norfloxacin
C0366095|T201|COMP|3868-7|LNC|Norfluoxetine|Norfluoxetine
C0366096|T201|COMP|3869-5|LNC|Normeperidine|Normeperidine
C0366097|T201|COMP|3870-3|LNC|Norpropoxyphene|Norpropoxyphene
C0366098|T201|COMP|3871-1|LNC|Norpropoxyphene|Norpropoxyphene
C0366099|T201|COMP|3872-9|LNC|Nortriptyline|Nortriptyline
C0366100|T201|COMP|3873-7|LNC|Nortriptyline|Nortriptyline
C0366101|T201|COMP|3874-5|LNC|Nortriptyline|Nortriptyline
C0366102|T201|COMP|3875-2|LNC|Nortriptyline|Nortriptyline
C0366103|T201|COMP|3876-0|LNC|Nortriptyline^trough >12h post dose|Nortriptyline^trough >12h post dose
C0366104|T201|COMP|3877-8|LNC|Ofloxacin|Ofloxacin
C0366105|T201|COMP|3878-6|LNC|Opiates|Opiates
C0366106|T201|COMP|3879-4|LNC|Opiates|Opiates
C0366107|T201|COMP|3880-2|LNC|Orphenadrine|Orphenadrine
C0366108|T201|COMP|3881-0|LNC|Ouabain|Ouabain
C0366109|T201|COMP|3882-8|LNC|Oxacillin|Oxacillin
C0366110|T201|COMP|3883-6|LNC|Oxandrolone|Oxandrolone
C0366111|T201|COMP|3884-4|LNC|Oxandrolone|Oxandrolone
C0366112|T201|COMP|3885-1|LNC|Oxandrolone|Oxandrolone
C0366113|T201|COMP|3886-9|LNC|Oxazepam|Oxazepam
C0366114|T201|COMP|3887-7|LNC|Oxazepam|Oxazepam
C0366115|T201|COMP|3888-5|LNC|Oxedrine|Oxedrine
C0366116|T201|COMP|3889-3|LNC|Oxprenolol|Oxprenolol
C0366117|T201|COMP|3890-1|LNC|Oxprenolol|Oxprenolol
C0366118|T201|COMP|3891-9|LNC|Oxprenolol|Oxprenolol
C0366119|T201|COMP|3892-7|LNC|Oxprenolol|Oxprenolol
C0366120|T201|COMP|3893-5|LNC|oxyCODONE|oxyCODONE
C0366121|T201|COMP|3894-3|LNC|Oxymesterone|Oxymesterone
C0366122|T201|COMP|3895-0|LNC|Oxymesterone|Oxymesterone
C0366123|T201|COMP|3896-8|LNC|Oxymesterone|Oxymesterone
C0366124|T201|COMP|3897-6|LNC|Oxymetholone|Oxymetholone
C0366125|T201|COMP|3898-4|LNC|Oxymetholone|Oxymetholone
C0366126|T201|COMP|3899-2|LNC|Oxymetholone|Oxymetholone
C0366127|T201|COMP|3900-8|LNC|Oxyphenbutazone|Oxyphenbutazone
C0366128|T201|COMP|3901-6|LNC|Para hydroxyamphetamine|Para hydroxyamphetamine
C0366129|T201|COMP|3902-4|LNC|Para hydroxyamphetamine|Para hydroxyamphetamine
C0366130|T201|COMP|3903-2|LNC|Para hydroxyamphetamine|Para hydroxyamphetamine
C0366131|T201|COMP|3904-0|LNC|Paraldehyde|Paraldehyde
C0366132|T201|COMP|3905-7|LNC|Paraldehyde|Paraldehyde
C0366133|T201|COMP|3906-5|LNC|Pefloxacin|Pefloxacin
C0366134|T201|COMP|3907-3|LNC|Pemoline|Pemoline
C0366135|T201|COMP|3908-1|LNC|Pemoline|Pemoline
C0366136|T201|COMP|3909-9|LNC|Pemoline|Pemoline
C0366137|T201|COMP|3910-7|LNC|Pemoline|Pemoline
C0366138|T201|COMP|3911-5|LNC|Penicillin|Penicillin
C0366139|T201|COMP|3912-3|LNC|Penicillin|Penicillin
C0366140|T201|COMP|3913-1|LNC|Penicillin G|Penicillin G
C0366141|T201|COMP|3914-9|LNC|Penicillin V|Penicillin V
C0366142|T201|COMP|3915-6|LNC|Pentazocine|Pentazocine
C0366143|T201|COMP|3916-4|LNC|Pentazocine|Pentazocine
C0366144|T201|COMP|3917-2|LNC|Pentazocine|Pentazocine
C0366145|T201|COMP|3918-0|LNC|Pentazocine|Pentazocine
C0366146|T201|COMP|3919-8|LNC|Pentazocine|Pentazocine
C0366147|T201|COMP|3920-6|LNC|Pentetrazol|Pentetrazol
C0366148|T201|COMP|3921-4|LNC|Pentetrazol|Pentetrazol
C0366149|T201|COMP|3922-2|LNC|Pentetrazol|Pentetrazol
C0366150|T201|COMP|3923-0|LNC|PENTobarbital|PENTobarbital
C0366151|T201|COMP|3924-8|LNC|PENTobarbital|PENTobarbital
C0366152|T201|COMP|3925-5|LNC|PENTobarbital|PENTobarbital
C0366153|T201|COMP|3926-3|LNC|PENTobarbital|PENTobarbital
C0366154|T201|COMP|3927-1|LNC|Perphenazine|Perphenazine
C0366155|T201|COMP|3928-9|LNC|Perphenazine|Perphenazine
C0366156|T201|COMP|3929-7|LNC|Phenacetin|Phenacetin
C0366157|T201|COMP|3930-5|LNC|Phenacetin|Phenacetin
C0366158|T201|COMP|3931-3|LNC|Phenazocine|Phenazocine
C0366159|T201|COMP|3932-1|LNC|Phenazocine|Phenazocine
C0366160|T201|COMP|3933-9|LNC|Phenazocine|Phenazocine
C0366161|T201|COMP|3934-7|LNC|Phencyclidine|Phencyclidine
C0366162|T201|COMP|3935-4|LNC|Phencyclidine|Phencyclidine
C0366163|T201|COMP|3936-2|LNC|Phencyclidine|Phencyclidine
C0366164|T201|COMP|3937-0|LNC|Phencyclidine|Phencyclidine
C0366165|T201|COMP|3938-8|LNC|Phendimetrazine|Phendimetrazine
C0366166|T201|COMP|3939-6|LNC|Phendimetrazine|Phendimetrazine
C0366167|T201|COMP|3940-4|LNC|Phendimetrazine|Phendimetrazine
C0366168|T201|COMP|3941-2|LNC|Phendimetrazine|Phendimetrazine
C0366169|T201|COMP|3942-0|LNC|Pheniramine|Pheniramine
C0366170|T201|COMP|3943-8|LNC|Phenmetrazine|Phenmetrazine
C0366171|T201|COMP|3944-6|LNC|Phenmetrazine|Phenmetrazine
C0366172|T201|COMP|3945-3|LNC|Phenmetrazine|Phenmetrazine
C0366173|T201|COMP|3946-1|LNC|Phenmetrazine|Phenmetrazine
C0366174|T201|COMP|3947-9|LNC|PHENobarbital|PHENobarbital
C0366175|T201|COMP|3948-7|LNC|PHENobarbital|PHENobarbital
C0366176|T201|COMP|3949-5|LNC|PHENobarbital|PHENobarbital
C0366177|T201|COMP|3950-3|LNC|PHENobarbital|PHENobarbital
C0366178|T201|COMP|3951-1|LNC|PHENobarbital.free|PHENobarbital.free
C0366179|T201|COMP|3952-9|LNC|Phenothiazines|Phenothiazines
C0366180|T201|COMP|3953-7|LNC|Phenothiazines|Phenothiazines
C0366181|T201|COMP|3954-5|LNC|Phenothiazines|Phenothiazines
C0366182|T201|COMP|3955-2|LNC|Phensuximide|Phensuximide
C0366183|T201|COMP|3956-0|LNC|Phentermine|Phentermine
C0366184|T201|COMP|3957-8|LNC|Phentermine|Phentermine
C0366185|T201|COMP|3958-6|LNC|Phentermine|Phentermine
C0366186|T201|COMP|3959-4|LNC|Phentermine|Phentermine
C0366187|T201|COMP|3960-2|LNC|Phenylbutazone|Phenylbutazone
C0366188|T201|COMP|3961-0|LNC|Phenylbutazone|Phenylbutazone
C0366189|T201|COMP|3962-8|LNC|Phenylephrine|Phenylephrine
C0366190|T201|COMP|3963-6|LNC|Phenylpropanolamine|Phenylpropanolamine
C0366191|T201|COMP|3964-4|LNC|Phenylpropanolamine|Phenylpropanolamine
C0366192|T201|COMP|3965-1|LNC|Phenylpropanolamine|Phenylpropanolamine
C0366193|T201|COMP|3966-9|LNC|Phenylpropanolamine|Phenylpropanolamine
C0366194|T201|COMP|3967-7|LNC|Phenytoin|Phenytoin
C0366195|T201|COMP|3968-5|LNC|Phenytoin|Phenytoin
C0366196|T201|COMP|3969-3|LNC|Phenytoin.free|Phenytoin.free
C0366197|T201|COMP|3970-1|LNC|Pholedrine|Pholedrine
C0366198|T201|COMP|3971-9|LNC|Pindolol|Pindolol
C0366199|T201|COMP|3972-7|LNC|Piperacillin|Piperacillin
C0366200|T201|COMP|3973-5|LNC|Pipradrol|Pipradrol
C0366201|T201|COMP|3974-3|LNC|Pipradrol|Pipradrol
C0366202|T201|COMP|3975-0|LNC|Pipradrol|Pipradrol
C0366203|T201|COMP|3976-8|LNC|Practolol|Practolol
C0366204|T201|COMP|3977-6|LNC|Prazepam|Prazepam
C0366205|T201|COMP|3978-4|LNC|Primidone|Primidone
C0366206|T201|COMP|3979-2|LNC|Probenecid|Probenecid
C0366207|T201|COMP|3980-0|LNC|Probenecid|Probenecid
C0366208|T201|COMP|3981-8|LNC|Probenecid|Probenecid
C0366209|T201|COMP|3982-6|LNC|Procainamide|Procainamide
C0366210|T201|COMP|3983-4|LNC|Procainamide+N-acetylprocainamide|Procainamide+N-acetylprocainamide
C0366211|T201|COMP|3984-2|LNC|Prolintane|Prolintane
C0366212|T201|COMP|3985-9|LNC|Prolintane|Prolintane
C0366213|T201|COMP|3986-7|LNC|Prolintane|Prolintane
C0366214|T201|COMP|3987-5|LNC|Promazine|Promazine
C0366215|T201|COMP|3988-3|LNC|Promethazine|Promethazine
C0366216|T201|COMP|3989-1|LNC|Promethazine|Promethazine
C0366217|T201|COMP|3991-7|LNC|Propranolol|Propranolol
C0366218|T201|COMP|3992-5|LNC|Propranolol|Propranolol
C0366219|T201|COMP|3993-3|LNC|Propranolol|Propranolol
C0366220|T201|COMP|3994-1|LNC|Propranolol|Propranolol
C0366221|T201|COMP|3990-9|LNC|Propranolol|Propranolol
C0366222|T201|COMP|3995-8|LNC|Propylhexedrine|Propylhexedrine
C0366223|T201|COMP|3996-6|LNC|Propylhexedrine|Propylhexedrine
C0366224|T201|COMP|3997-4|LNC|Propylhexedrine|Propylhexedrine
C0366225|T201|COMP|3998-2|LNC|Propylhexedrine|Propylhexedrine
C0366226|T201|COMP|3999-0|LNC|Protriptyline|Protriptyline
C0366227|T201|COMP|4000-6|LNC|Protriptyline|Protriptyline
C0366228|T201|COMP|4001-4|LNC|Protriptyline|Protriptyline
C0366229|T201|COMP|4002-2|LNC|Protriptyline^trough|Protriptyline^trough
C0366230|T201|COMP|4003-0|LNC|Pseudoephedrine|Pseudoephedrine
C0366231|T201|COMP|4004-8|LNC|Pseudoephedrine|Pseudoephedrine
C0366232|T201|COMP|4005-5|LNC|Pseudoephedrine|Pseudoephedrine
C0366233|T201|COMP|4006-3|LNC|Pyrilamine|Pyrilamine
C0366234|T201|COMP|4007-1|LNC|Pyrilamine|Pyrilamine
C0366235|T201|COMP|4008-9|LNC|Pyrilamine|Pyrilamine
C0366236|T201|COMP|4009-7|LNC|Pyrilamine|Pyrilamine
C0366237|T201|COMP|4010-5|LNC|Pyrilamine|Pyrilamine
C0366238|T201|COMP|4011-3|LNC|Pyrovalerone|Pyrovalerone
C0366239|T201|COMP|4012-1|LNC|Pyrovalerone|Pyrovalerone
C0366240|T201|COMP|4013-9|LNC|Pyrovalerone|Pyrovalerone
C0366241|T201|COMP|4014-7|LNC|quiNIDine|quiNIDine
C0366242|T201|COMP|4015-4|LNC|quiNIDine|quiNIDine
C0366243|T201|COMP|4016-2|LNC|quiNIDine+Quinine|quiNIDine+Quinine
C0366244|T201|COMP|4017-0|LNC|quiNIDine^trough|quiNIDine^trough
C0366245|T201|COMP|4018-8|LNC|quiNINE|quiNINE
C0366246|T201|COMP|4019-6|LNC|quiNINE|quiNINE
C0366247|T201|COMP|4020-4|LNC|quiNINE|quiNINE
C0366248|T201|COMP|4021-2|LNC|rifAMPin|rifAMPin
C0366249|T201|COMP|4022-0|LNC|Salicylamide|Salicylamide
C0366250|T201|COMP|4023-8|LNC|Salicylates|Salicylates
C0366251|T201|COMP|4024-6|LNC|Salicylates|Salicylates
C0366252|T201|COMP|4025-3|LNC|Salicylates|Salicylates
C0366253|T201|COMP|4026-1|LNC|Salicylates|Salicylates
C0366254|T201|COMP|4027-9|LNC|Secobarbital|Secobarbital
C0366255|T201|COMP|4028-7|LNC|Secobarbital|Secobarbital
C0366256|T201|COMP|4029-5|LNC|Secobarbital|Secobarbital
C0366257|T201|COMP|4030-3|LNC|Sotalol|Sotalol
C0366258|T201|COMP|4031-1|LNC|Sotalol|Sotalol
C0366259|T201|COMP|4032-9|LNC|Sotalol|Sotalol
C0366260|T201|COMP|4034-5|LNC|Spironolactone|Spironolactone
C0366261|T201|COMP|4035-2|LNC|Spironolactone|Spironolactone
C0366262|T201|COMP|4036-0|LNC|Stanozolol|Stanozolol
C0366263|T201|COMP|4037-8|LNC|Stanozolol|Stanozolol
C0366264|T201|COMP|4038-6|LNC|Stanozolol|Stanozolol
C0366265|T201|COMP|4039-4|LNC|Streptomycin|Streptomycin
C0366266|T201|COMP|4040-2|LNC|Sulfonamide|Sulfonamide
C0366267|T201|COMP|4041-0|LNC|Sulfonamide|Sulfonamide
C0366268|T201|COMP|4042-8|LNC|Sulfonamide|Sulfonamide
C0366269|T201|COMP|4043-6|LNC|Teicoplanin|Teicoplanin
C0366270|T201|COMP|4044-4|LNC|Tetracaine|Tetracaine
C0366271|T201|COMP|4045-1|LNC|Tetracycline|Tetracycline
C0366272|T201|COMP|4046-9|LNC|Tetrahydrocortisone|Tetrahydrocortisone
C0366273|T201|COMP|4047-7|LNC|Theophylline|Theophylline
C0366274|T201|COMP|4048-5|LNC|Theophylline|Theophylline
C0366275|T201|COMP|4049-3|LNC|Theophylline|Theophylline
C0366276|T201|COMP|4050-1|LNC|Thiopental|Thiopental
C0366277|T201|COMP|4051-9|LNC|Thioridazine|Thioridazine
C0366278|T201|COMP|4052-7|LNC|Thioridazine|Thioridazine
C0366279|T201|COMP|4053-5|LNC|Thioridazine|Thioridazine
C0366280|T201|COMP|4054-3|LNC|Ticarcillin|Ticarcillin
C0366281|T201|COMP|4055-0|LNC|Ticarcillin+Clavulanate|Ticarcillin+Clavulanate
C0366282|T201|COMP|4056-8|LNC|Timolol|Timolol
C0366283|T201|COMP|4057-6|LNC|Tobramycin^peak|Tobramycin^peak
C0366284|T201|COMP|4058-4|LNC|Tobramycin^random|Tobramycin^random
C0366285|T201|COMP|4059-2|LNC|Tobramycin^trough|Tobramycin^trough
C0366286|T201|COMP|4060-0|LNC|Tocainide|Tocainide
C0366287|T201|COMP|4061-8|LNC|TOLBUTamide|TOLBUTamide
C0366288|T201|COMP|4062-6|LNC|Tranylcypromine|Tranylcypromine
C0366289|T201|COMP|4063-4|LNC|traZODone|traZODone
C0366290|T201|COMP|4064-2|LNC|traZODone|traZODone
C0366291|T201|COMP|4065-9|LNC|traZODone|traZODone
C0366292|T201|COMP|4066-7|LNC|Triamterene|Triamterene
C0366293|T201|COMP|4067-5|LNC|Triamterene|Triamterene
C0366294|T201|COMP|4068-3|LNC|Triamterene|Triamterene
C0366295|T201|COMP|4069-1|LNC|Triazolam|Triazolam
C0366296|T201|COMP|4070-9|LNC|Triazolam|Triazolam
C0366297|T201|COMP|4071-7|LNC|Chloral hydrate|Chloral hydrate
C0366298|T201|COMP|4072-5|LNC|Chloral hydrate|Chloral hydrate
C0366299|T201|COMP|4073-3|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0366300|T201|COMP|4074-1|LNC|Trifluoperazine|Trifluoperazine
C0366301|T201|COMP|4075-8|LNC|Trimeperidine|Trimeperidine
C0366302|T201|COMP|4076-6|LNC|Trimeperidine|Trimeperidine
C0366303|T201|COMP|4077-4|LNC|Trimeperidine|Trimeperidine
C0366304|T201|COMP|4078-2|LNC|Trimethadione|Trimethadione
C0366305|T201|COMP|4079-0|LNC|Trimethoprim|Trimethoprim
C0366306|T201|COMP|4080-8|LNC|Trimethoprim|Trimethoprim
C0366307|T201|COMP|4081-6|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0366308|T201|COMP|4082-4|LNC|Trimipramine|Trimipramine
C0366309|T201|COMP|4083-2|LNC|Trimipramine|Trimipramine
C0366310|T201|COMP|4084-0|LNC|Trimipramine|Trimipramine
C0366311|T201|COMP|4085-7|LNC|Tripelennamine|Tripelennamine
C0366312|T201|COMP|4086-5|LNC|Valproate|Valproate
C0366313|T201|COMP|4087-3|LNC|Valproate.free|Valproate.free
C0366314|T201|COMP|4088-1|LNC|Valproate^trough|Valproate^trough
C0366315|T201|COMP|4089-9|LNC|Vancomycin.free|Vancomycin.free
C0366316|T201|COMP|4090-7|LNC|Vancomycin^peak|Vancomycin^peak
C0366317|T201|COMP|4091-5|LNC|Vancomycin^random|Vancomycin^random
C0366318|T201|COMP|4092-3|LNC|Vancomycin^trough|Vancomycin^trough
C0366319|T201|COMP|4093-1|LNC|Verapamil|Verapamil
C0366320|T201|COMP|4094-9|LNC|Verapamil|Verapamil
C0366321|T201|COMP|4095-6|LNC|Verapamil|Verapamil
C0366322|T201|COMP|4096-4|LNC|Volatile drugs negative|Volatile drugs negative
C0366323|T201|COMP|4097-2|LNC|Volatile drugs positive|Volatile drugs positive
C0366324|T201|COMP|4098-0|LNC|Warfarin|Warfarin
C0366325|T201|COMP|4099-8|LNC|Zimelidine|Zimelidine
C0366326|T201|COMP|4100-4|LNC|2-Oxoisocaproate|2-Oxoisocaproate
C0366327|T201|COMP|4101-2|LNC|2-Pyridone|2-Pyridone
C0366329|T201|COMP|4103-8|LNC|Acebutolol|Acebutolol
C0366330|T201|COMP|4104-6|LNC|Acepromazine|Acepromazine
C0366331|T201|COMP|4105-3|LNC|Acetaminophen|Acetaminophen
C0366332|T201|COMP|4106-1|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C0366334|T201|COMP|4108-7|LNC|Adenine|Adenine
C0366335|T201|COMP|4109-5|LNC|Alfentanil|Alfentanil
C0366336|T201|COMP|4110-3|LNC|Alphaprodine|Alphaprodine
C0366337|T201|COMP|4111-1|LNC|ALPRAZolam|ALPRAZolam
C0366338|T201|COMP|4112-9|LNC|Alprenolol|Alprenolol
C0366339|T201|COMP|4113-7|LNC|Amantadine|Amantadine
C0366340|T201|COMP|4114-5|LNC|Amdinocillin|Amdinocillin
C0366341|T201|COMP|4115-2|LNC|Amikacin|Amikacin
C0366342|T201|COMP|4116-0|LNC|aMILoride|aMILoride
C0366343|T201|COMP|4117-8|LNC|Aminopyrine|Aminopyrine
C0366344|T201|COMP|4118-6|LNC|Aminosalicylate|Aminosalicylate
C0366345|T201|COMP|4119-4|LNC|Amiodarone|Amiodarone
C0366346|T201|COMP|4120-2|LNC|Amitriptyline|Amitriptyline
C0366347|T201|COMP|4121-0|LNC|Amobarbital|Amobarbital
C0366348|T201|COMP|4122-8|LNC|Amoxapine|Amoxapine
C0366350|T201|COMP|4124-4|LNC|Diethylpropion|Diethylpropion
C0366351|T201|COMP|4125-1|LNC|Amphetaminil|Amphetaminil
C0366352|T201|COMP|4126-9|LNC|Amphotericin B|Amphotericin B
C0366353|T201|COMP|4127-7|LNC|Ampicillin|Ampicillin
C0366354|T201|COMP|4128-5|LNC|Anileridine|Anileridine
C0366355|T201|COMP|4129-3|LNC|Anthraquinone|Anthraquinone
C0366356|T201|COMP|4130-1|LNC|Antipyrine|Antipyrine
C0366357|T201|COMP|4131-9|LNC|Ascorbate.PO|Ascorbate.PO
C0366360|T201|COMP|4134-3|LNC|Azlocillin|Azlocillin
C0366361|T201|COMP|4135-0|LNC|Aztreonam|Aztreonam
C0366362|T201|COMP|4136-8|LNC|Barbital|Barbital
C0366363|T201|COMP|4137-6|LNC|Barbiturates|Barbiturates
C0366364|T201|COMP|4138-4|LNC|Bendroflumethiazide|Bendroflumethiazide
C0366365|T201|COMP|4139-2|LNC|Benzfetamine|Benzfetamine
C0366366|T201|COMP|4140-0|LNC|Benzoylecgonine|Benzoylecgonine
C0366367|T201|COMP|4141-8|LNC|Benzthiazide|Benzthiazide
C0366368|T201|COMP|4142-6|LNC|Bisacodyl|Bisacodyl
C0366369|T201|COMP|4143-4|LNC|Bolasterone|Bolasterone
C0366370|T201|COMP|4144-2|LNC|Bromazepam|Bromazepam
C0366371|T201|COMP|4145-9|LNC|Brompheniramine|Brompheniramine
C0366372|T201|COMP|4146-7|LNC|Bumetanide|Bumetanide
C0366373|T201|COMP|4147-5|LNC|Buprenorphine|Buprenorphine
C0366374|T201|COMP|4148-3|LNC|Butabarbital|Butabarbital
C0366375|T201|COMP|4149-1|LNC|Butalbital|Butalbital
C0366377|T201|COMP|4151-7|LNC|Canrenone|Canrenone
C0366378|T201|COMP|4152-5|LNC|carBAMazepine|carBAMazepine
C0366379|T201|COMP|4153-3|LNC|Carbenicillin|Carbenicillin
C0366380|T201|COMP|4154-1|LNC|Carbromal|Carbromal
C0366381|T201|COMP|4155-8|LNC|Carisoprodol|Carisoprodol
C0366382|T201|COMP|4156-6|LNC|Cathine|Cathine
C0366383|T201|COMP|4157-4|LNC|Cefamandole|Cefamandole
C0366385|T201|COMP|4159-0|LNC|ceFAZolin|ceFAZolin
C0366386|T201|COMP|4160-8|LNC|Cefonicid|Cefonicid
C0366387|T201|COMP|4161-6|LNC|Cefoperazone|Cefoperazone
C0366388|T201|COMP|4162-4|LNC|Cefotaxime|Cefotaxime
C0366389|T201|COMP|4163-2|LNC|cefoTEtan|cefoTEtan
C0366390|T201|COMP|4164-0|LNC|cefOXitin|cefOXitin
C0366391|T201|COMP|4165-7|LNC|Cefsulodin|Cefsulodin
C0366392|T201|COMP|4166-5|LNC|cefTAZidime|cefTAZidime
C0366393|T201|COMP|4167-3|LNC|Ceftizoxime|Ceftizoxime
C0366394|T201|COMP|4168-1|LNC|cefTRIAXone|cefTRIAXone
C0366395|T201|COMP|4169-9|LNC|Cefuroxime.parenteral|Cefuroxime.parenteral
C0366397|T201|COMP|4171-5|LNC|Cephalothin|Cephalothin
C0366398|T201|COMP|4172-3|LNC|Chloral hydrate|Chloral hydrate
C0366399|T201|COMP|4173-1|LNC|Chloramphenicol|Chloramphenicol
C0366400|T201|COMP|4174-9|LNC|Clorazepate|Clorazepate
C0366401|T201|COMP|4175-6|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0366402|T201|COMP|4176-4|LNC|Chlormerodrin|Chlormerodrin
C0366403|T201|COMP|4177-2|LNC|Chlorothiazide|Chlorothiazide
C0366404|T201|COMP|4178-0|LNC|Chlorpheniramine|Chlorpheniramine
C0366405|T201|COMP|4179-8|LNC|chlorproMAZINE|chlorproMAZINE
C0366406|T201|COMP|4180-6|LNC|chlorproPAMIDE|chlorproPAMIDE
C0366407|T201|COMP|4181-4|LNC|Chlorprothixene|Chlorprothixene
C0366408|T201|COMP|4182-2|LNC|Chloroquine|Chloroquine
C0366409|T201|COMP|4183-0|LNC|Chlorthalidone|Chlorthalidone
C0366410|T201|COMP|4184-8|LNC|Cilastatin|Cilastatin
C0366411|T201|COMP|4185-5|LNC|Cimetidine|Cimetidine
C0366414|T201|COMP|4188-9|LNC|Clavulanate|Clavulanate
C0366416|T201|COMP|4190-5|LNC|cloBAZam|cloBAZam
C0366417|T201|COMP|4191-3|LNC|Clobenzorex|Clobenzorex
C0366418|T201|COMP|4192-1|LNC|Clofibrate|Clofibrate
C0366420|T201|COMP|4194-7|LNC|clonazePAM|clonazePAM
C0366421|T201|COMP|4195-4|LNC|cloNIDine|cloNIDine
C0366422|T201|COMP|4196-2|LNC|Clopenthixol|Clopenthixol
C0366423|T201|COMP|4197-0|LNC|Clorprenaline|Clorprenaline
C0366424|T201|COMP|4198-8|LNC|Clostebol|Clostebol
C0366426|T201|COMP|4200-2|LNC|Prochlorperazine|Prochlorperazine
C0366427|T201|COMP|4201-0|LNC|Cropropamide|Cropropamide
C0366428|T201|COMP|4202-8|LNC|Crotetamide|Crotetamide
C0366429|T201|COMP|4203-6|LNC|Cyanocobalamin.PO|Cyanocobalamin.PO
C0366430|T201|COMP|4204-4|LNC|Cyclacillin|Cyclacillin
C0366431|T201|COMP|4205-1|LNC|Cyclizine|Cyclizine
C0366432|T201|COMP|4206-9|LNC|cycloSERINE|cycloSERINE
C0366433|T201|COMP|4207-7|LNC|cycloSPORINE|cycloSPORINE
C0366434|T201|COMP|4208-5|LNC|Dantron|Dantron
C0366435|T201|COMP|4193-9|LNC|clomiPRAMINE|clomiPRAMINE
C0366437|T201|COMP|4211-9|LNC|Desethylamiodarone|Desethylamiodarone
C0366440|T201|COMP|4214-3|LNC|Dextromethorphan|Dextromethorphan
C0366441|T201|COMP|4215-0|LNC|Dextromoramide|Dextromoramide
C0366442|T201|COMP|4216-8|LNC|Diamorphine|Diamorphine
C0366443|T201|COMP|4217-6|LNC|diazePAM|diazePAM
C0366444|T201|COMP|4218-4|LNC|Dibenzepin|Dibenzepin
C0366445|T201|COMP|4219-2|LNC|Dibucaine nbr|Dibucaine nbr
C0366446|T201|COMP|4220-0|LNC|Dichlorphenamide|Dichlorphenamide
C0366447|T201|COMP|4221-8|LNC|Digitoxin|Digitoxin
C0366450|T201|COMP|4224-2|LNC|diphenhydrAMINE|diphenhydrAMINE
C0366452|T201|COMP|4226-7|LNC|Diphenylhydramine|Diphenylhydramine
C0366453|T201|COMP|4227-5|LNC|Dipipanone|Dipipanone
C0366454|T201|COMP|4228-3|LNC|Disopyramide|Disopyramide
C0366455|T201|COMP|4229-1|LNC|Disulfiram|Disulfiram
C0366456|T201|COMP|4230-9|LNC|Doxepin|Doxepin
C0366457|T201|COMP|4231-7|LNC|Doxylamine|Doxylamine
C0366458|T201|COMP|4232-5|LNC|Dyphylline|Dyphylline
C0366459|T201|COMP|4233-3|LNC|Emetine|Emetine
C0366460|T201|COMP|4234-1|LNC|Encainide|Encainide
C0366461|T201|COMP|4235-8|LNC|Enoxacin|Enoxacin
C0366462|T201|COMP|4236-6|LNC|ePHEDrine|ePHEDrine
C0366463|T201|COMP|4237-4|LNC|Erythromycin|Erythromycin
C0366464|T201|COMP|4238-2|LNC|Estazolam|Estazolam
C0366465|T201|COMP|4239-0|LNC|Etafedrine|Etafedrine
C0366466|T201|COMP|4240-8|LNC|Etamivan|Etamivan
C0366467|T201|COMP|4241-6|LNC|Ethacrynate|Ethacrynate
C0366468|T201|COMP|4242-4|LNC|Ethambutol|Ethambutol
C0366469|T201|COMP|4243-2|LNC|Ethchlorvynol|Ethchlorvynol
C0366470|T201|COMP|4244-0|LNC|Ethoheptazine|Ethoheptazine
C0366471|T201|COMP|4245-7|LNC|Ethosuximide|Ethosuximide
C0366472|T201|COMP|4246-5|LNC|Ethotoin|Ethotoin
C0366473|T201|COMP|4247-3|LNC|Ethylmorphine|Ethylmorphine
C0366475|T201|COMP|4249-9|LNC|Etilefrine|Etilefrine
C0366476|T201|COMP|4250-7|LNC|Fencamfamin|Fencamfamin
C0366477|T201|COMP|4251-5|LNC|Fenetylline|Fenetylline
C0366478|T201|COMP|4252-3|LNC|Fenfluramine|Fenfluramine
C0366479|T201|COMP|4253-1|LNC|Fenoprofen|Fenoprofen
C0366480|T201|COMP|4254-9|LNC|Fenproporex|Fenproporex
C0366481|T201|COMP|4255-6|LNC|fentaNYL|fentaNYL
C0366482|T201|COMP|4256-4|LNC|Flecainide|Flecainide
C0366483|T201|COMP|4102-0|LNC|5-Fluorocytosine|5-Fluorocytosine
C0366484|T201|COMP|4258-0|LNC|Flunitrazepam|Flunitrazepam
C0366485|T201|COMP|4259-8|LNC|Fluorouracil|Fluorouracil
C0366486|T201|COMP|4260-6|LNC|FLUoxetine|FLUoxetine
C0366487|T201|COMP|4261-4|LNC|Fluoxymesterone|Fluoxymesterone
C0366488|T201|COMP|4262-2|LNC|Flupenthixol|Flupenthixol
C0366489|T201|COMP|4263-0|LNC|fluPHENAZine|fluPHENAZine
C0366490|T201|COMP|4264-8|LNC|Flurazepam|Flurazepam
C0366491|T201|COMP|4265-5|LNC|Furfenorex|Furfenorex
C0366492|T201|COMP|4266-3|LNC|Furosemide|Furosemide
C0366493|T201|COMP|4267-1|LNC|Galactose.PO|Galactose.PO
C0366494|T201|COMP|4268-9|LNC|Gentamicin|Gentamicin
C0366495|T201|COMP|4269-7|LNC|Glucose.PO|Glucose.PO
C0366496|T201|COMP|4270-5|LNC|Glutethimide|Glutethimide
C0366497|T201|COMP|4271-3|LNC|Gonadotropin releasing hormone|Gonadotropin releasing hormone
C0366498|T201|COMP|4272-1|LNC|Haloperidol|Haloperidol
C0366499|T201|COMP|4273-9|LNC|Heptaminol|Heptaminol
C0366500|T201|COMP|4274-7|LNC|Hippurate|Hippurate
C0366501|T201|COMP|4275-4|LNC|hydroCHLOROthiazide|hydroCHLOROthiazide
C0366502|T201|COMP|4276-2|LNC|HYDROcodone|HYDROcodone
C0366503|T201|COMP|4223-4|LNC|HYDROmorphone|HYDROmorphone
C0366504|T201|COMP|4278-8|LNC|Hydroxychloroquine|Hydroxychloroquine
C0366505|T201|COMP|4279-6|LNC|Hydroxymethoxyphenamine|Hydroxymethoxyphenamine
C0366506|T201|COMP|4280-4|LNC|hydrOXYzine|hydrOXYzine
C0366508|T201|COMP|4282-0|LNC|Imipenem|Imipenem
C0366509|T201|COMP|4283-8|LNC|Imipramine|Imipramine
C0366510|T201|COMP|4284-6|LNC|Indomethacin|Indomethacin
C0366511|T201|COMP|4285-3|LNC|Insulin Lente|Insulin Lente
C0366512|T201|COMP|4286-1|LNC|Insulin NPH|Insulin NPH
C0366513|T201|COMP|4287-9|LNC|Insulin regular|Insulin regular
C0366514|T201|COMP|4288-7|LNC|Insulin semilente|Insulin semilente
C0366515|T201|COMP|4289-5|LNC|Insulin ultralente|Insulin ultralente
C0366516|T201|COMP|4290-3|LNC|Isoniazid|Isoniazid
C0366517|T201|COMP|4291-1|LNC|Kanamycin|Kanamycin
C0366518|T201|COMP|4292-9|LNC|Ketamine|Ketamine
C0366519|T201|COMP|4293-7|LNC|Ketobemidone|Ketobemidone
C0366520|T201|COMP|4294-5|LNC|Levodopa.PO|Levodopa.PO
C0366521|T201|COMP|4295-2|LNC|Labetalol|Labetalol
C0366522|T201|COMP|4296-0|LNC|Methotrimeprazine|Methotrimeprazine
C0366523|T201|COMP|4297-8|LNC|Levomepromazine|Levomepromazine
C0366524|T201|COMP|4298-6|LNC|Levorphanol|Levorphanol
C0366525|T201|COMP|4299-4|LNC|Lidocaine|Lidocaine
C0366527|T201|COMP|4301-8|LNC|LORazepam|LORazepam
C0366528|T201|COMP|4302-6|LNC|Lormetazepam|Lormetazepam
C0366529|T201|COMP|4303-4|LNC|Loxapine|Loxapine
C0366530|T201|COMP|4304-2|LNC|Maprotiline|Maprotiline
C0366531|T201|COMP|4305-9|LNC|Medazepam|Medazepam
C0366532|T201|COMP|4306-7|LNC|Mefenorex|Mefenorex
C0366535|T201|COMP|4309-1|LNC|Mephobarbital|Mephobarbital
C0366536|T201|COMP|4310-9|LNC|Meprobamate|Meprobamate
C0366537|T201|COMP|4311-7|LNC|Mersalyl|Mersalyl
C0366538|T201|COMP|4308-3|LNC|Mephenytoin|Mephenytoin
C0366539|T201|COMP|4313-3|LNC|Mesoridazine|Mesoridazine
C0366540|T201|COMP|4314-1|LNC|Mesterolone|Mesterolone
C0366541|T201|COMP|4315-8|LNC|Metandienone|Metandienone
C0366542|T201|COMP|4316-6|LNC|Metaraminol|Metaraminol
C0366543|T201|COMP|4317-4|LNC|Metenolone|Metenolone
C0366545|T201|COMP|4319-0|LNC|Methamphetamine|Methamphetamine
C0366546|T201|COMP|4320-8|LNC|Methapyrilene|Methapyrilene
C0366547|T201|COMP|4321-6|LNC|Methaqualone|Methaqualone
C0366548|T201|COMP|4322-4|LNC|Methicillin|Methicillin
C0366549|T201|COMP|4323-2|LNC|Methocarbamol|Methocarbamol
C0366550|T201|COMP|4324-0|LNC|Methotrexate|Methotrexate
C0366551|T201|COMP|4325-7|LNC|Methoxyphenamine|Methoxyphenamine
C0366552|T201|COMP|4326-5|LNC|Methsuximide|Methsuximide
C0366553|T201|COMP|4327-3|LNC|Methyldopa|Methyldopa
C0366554|T201|COMP|4328-1|LNC|MethylePHEDrine|MethylePHEDrine
C0366555|T201|COMP|4329-9|LNC|Methylphenidate|Methylphenidate
C0366556|T201|COMP|4330-7|LNC|Methyprylon|Methyprylon
C0366558|T201|COMP|4332-3|LNC|Mexiletine|Mexiletine
C0366559|T201|COMP|4333-1|LNC|Mezlocillin|Mezlocillin
C0366560|T201|COMP|4334-9|LNC|Midazolam|Midazolam
C0366561|T201|COMP|4335-6|LNC|Minocycline|Minocycline
C0366562|T201|COMP|4336-4|LNC|Morazone|Morazone
C0366564|T201|COMP|4338-0|LNC|Moxalactam|Moxalactam
C0366565|T201|COMP|4339-8|LNC|N-acetylprocainamide|N-acetylprocainamide
C0366566|T201|COMP|4248-1|LNC|N-ethylnicotinamide|N-ethylnicotinamide
C0366567|T201|COMP|4341-4|LNC|Nadolol|Nadolol
C0366568|T201|COMP|4342-2|LNC|Nalbuphine|Nalbuphine
C0366569|T201|COMP|4343-0|LNC|Nalorphine|Nalorphine
C0366570|T201|COMP|4344-8|LNC|Nandrolone|Nandrolone
C0366571|T201|COMP|4345-5|LNC|Naproxen|Naproxen
C0366572|T201|COMP|4346-3|LNC|Neopterin|Neopterin
C0366573|T201|COMP|4347-1|LNC|Netilmicin|Netilmicin
C0366574|T201|COMP|4348-9|LNC|Nicomorphine|Nicomorphine
C0366575|T201|COMP|4349-7|LNC|Nicotinamide|Nicotinamide
C0366576|T201|COMP|4350-5|LNC|Nicotine|Nicotine
C0366577|T201|COMP|4351-3|LNC|Nikethamide|Nikethamide
C0366578|T201|COMP|4352-1|LNC|Nitrazepam|Nitrazepam
C0366579|T201|COMP|4353-9|LNC|Nitrofurantoin|Nitrofurantoin
C0366580|T201|COMP|4213-5|LNC|Nordiazepam|Nordiazepam
C0366581|T201|COMP|4210-1|LNC|Nordoxepin|Nordoxepin
C0366582|T201|COMP|4356-2|LNC|Norepinephrine|Norepinephrine
C0366583|T201|COMP|4357-0|LNC|Norethandrolone|Norethandrolone
C0366584|T201|COMP|4358-8|LNC|Norfenefrine|Norfenefrine
C0366585|T201|COMP|4359-6|LNC|Norfloxacin|Norfloxacin
C0366586|T201|COMP|4360-4|LNC|Normetanephrine|Normetanephrine
C0366587|T201|COMP|4361-2|LNC|Nortriptyline|Nortriptyline
C0366588|T201|COMP|4362-0|LNC|Ofloxacin|Ofloxacin
C0366589|T201|COMP|4363-8|LNC|Orphenadrine|Orphenadrine
C0366590|T201|COMP|4364-6|LNC|Ouabain|Ouabain
C0366591|T201|COMP|4365-3|LNC|Oxacillin|Oxacillin
C0366592|T201|COMP|4366-1|LNC|Oxandrolone|Oxandrolone
C0366593|T201|COMP|4367-9|LNC|Oxazepam|Oxazepam
C0366594|T201|COMP|4368-7|LNC|Oxedrine|Oxedrine
C0366595|T201|COMP|4369-5|LNC|Oxprenolol|Oxprenolol
C0366597|T201|COMP|4371-1|LNC|Oxymesterone|Oxymesterone
C0366598|T201|COMP|4372-9|LNC|Oxymetholone|Oxymetholone
C0366599|T201|COMP|4373-7|LNC|Oxyphenbutazone|Oxyphenbutazone
C0366600|T201|COMP|4374-5|LNC|Para methylhippurate|Para methylhippurate
C0366601|T201|COMP|4375-2|LNC|Para hydroxyamphetamine|Para hydroxyamphetamine
C0366602|T201|COMP|4376-0|LNC|Paraldehyde|Paraldehyde
C0366603|T201|COMP|4377-8|LNC|Pefloxacin|Pefloxacin
C0366604|T201|COMP|4378-6|LNC|Pemoline|Pemoline
C0366605|T201|COMP|4379-4|LNC|Penicillin G benzathine|Penicillin G benzathine
C0366606|T201|COMP|4380-2|LNC|Penicillin G potassium|Penicillin G potassium
C0366607|T201|COMP|4381-0|LNC|Penicillin G procaine|Penicillin G procaine
C0366608|T201|COMP|4382-8|LNC|Penicillin V potassium|Penicillin V potassium
C0366609|T201|COMP|4383-6|LNC|Pentazocine|Pentazocine
C0366610|T201|COMP|4384-4|LNC|Pentetrazol|Pentetrazol
C0366611|T201|COMP|4385-1|LNC|PENTobarbital|PENTobarbital
C0366612|T201|COMP|4386-9|LNC|Perphenazine|Perphenazine
C0366613|T201|COMP|4387-7|LNC|Phenacetin|Phenacetin
C0366614|T201|COMP|4388-5|LNC|Phenazocine|Phenazocine
C0366615|T201|COMP|4389-3|LNC|Phencyclidine|Phencyclidine
C0366616|T201|COMP|4390-1|LNC|Phendimetrazine|Phendimetrazine
C0366617|T201|COMP|4391-9|LNC|Pheniramine|Pheniramine
C0366618|T201|COMP|4392-7|LNC|Phenmetrazine|Phenmetrazine
C0366619|T201|COMP|4393-5|LNC|PHENobarbital|PHENobarbital
C0366620|T201|COMP|4394-3|LNC|Phenothiazines|Phenothiazines
C0366621|T201|COMP|4395-0|LNC|Phensuximide|Phensuximide
C0366622|T201|COMP|4396-8|LNC|Phentermine|Phentermine
C0366623|T201|COMP|4397-6|LNC|Phenylbutazone|Phenylbutazone
C0366624|T201|COMP|4398-4|LNC|Phenylephrine|Phenylephrine
C0366625|T201|COMP|4399-2|LNC|Phenylpropanolamine|Phenylpropanolamine
C0366626|T201|COMP|4225-9|LNC|Phenytoin|Phenytoin
C0366627|T201|COMP|4401-6|LNC|Pholedrine|Pholedrine
C0366628|T201|COMP|4402-4|LNC|Pindolol|Pindolol
C0366629|T201|COMP|4403-2|LNC|Piperacillin|Piperacillin
C0366630|T201|COMP|4404-0|LNC|Pipradrol|Pipradrol
C0366631|T201|COMP|4405-7|LNC|Practolol|Practolol
C0366632|T201|COMP|4406-5|LNC|Prazepam|Prazepam
C0366633|T201|COMP|4407-3|LNC|Primidone|Primidone
C0366634|T201|COMP|4408-1|LNC|Probenecid|Probenecid
C0366635|T201|COMP|4409-9|LNC|Procainamide|Procainamide
C0366636|T201|COMP|4410-7|LNC|Prolintane|Prolintane
C0366637|T201|COMP|4411-5|LNC|Promazine|Promazine
C0366638|T201|COMP|4412-3|LNC|Promethazine|Promethazine
C0366639|T201|COMP|4413-1|LNC|Propanol|Propanol
C0366640|T201|COMP|4414-9|LNC|Propranolol|Propranolol
C0366641|T201|COMP|4415-6|LNC|Propylhexedrine|Propylhexedrine
C0366642|T201|COMP|4416-4|LNC|Protriptyline|Protriptyline
C0366643|T201|COMP|4417-2|LNC|Pseudoephedrine|Pseudoephedrine
C0366644|T201|COMP|4418-0|LNC|Pyrilamine|Pyrilamine
C0366645|T201|COMP|4419-8|LNC|quiNIDine|quiNIDine
C0366646|T201|COMP|4420-6|LNC|quiNINE|quiNINE
C0366647|T201|COMP|4421-4|LNC|rifAMPin|rifAMPin
C0366648|T201|COMP|4422-2|LNC|Salicylamide|Salicylamide
C0366649|T201|COMP|4423-0|LNC|Salicylates|Salicylates
C0366650|T201|COMP|4424-8|LNC|Secobarbital|Secobarbital
C0366651|T201|COMP|4425-5|LNC|Sotalol|Sotalol
C0366652|T201|COMP|4426-3|LNC|Spironolactone|Spironolactone
C0366653|T201|COMP|4427-1|LNC|Stanozolol|Stanozolol
C0366654|T201|COMP|4428-9|LNC|Streptomycin|Streptomycin
C0366655|T201|COMP|4429-7|LNC|Sulbactam|Sulbactam
C0366656|T201|COMP|4430-5|LNC|sulfADIAZINE|sulfADIAZINE
C0366657|T201|COMP|4431-3|LNC|Sulfamethoxazole|Sulfamethoxazole
C0366658|T201|COMP|4432-1|LNC|sulfiSOXAZOLE|sulfiSOXAZOLE
C0366659|T201|COMP|4433-9|LNC|Sulfonamide|Sulfonamide
C0366660|T201|COMP|4435-4|LNC|Teicoplanin|Teicoplanin
C0366661|T201|COMP|4436-2|LNC|Tetracaine|Tetracaine
C0366662|T201|COMP|4437-0|LNC|Tetracycline|Tetracycline
C0366663|T201|COMP|4438-8|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0366664|T201|COMP|4439-6|LNC|Tetrahydrocortisone|Tetrahydrocortisone
C0366665|T201|COMP|4440-4|LNC|Theophylline|Theophylline
C0366666|T201|COMP|4441-2|LNC|Thiopental|Thiopental
C0366667|T201|COMP|4442-0|LNC|Thioridazine|Thioridazine
C0366668|T201|COMP|4443-8|LNC|Ticarcillin|Ticarcillin
C0366669|T201|COMP|4444-6|LNC|Timolol|Timolol
C0366671|T201|COMP|4446-1|LNC|Tocainide|Tocainide
C0366672|T201|COMP|4447-9|LNC|TOLBUTamide|TOLBUTamide
C0366673|T201|COMP|4448-7|LNC|TOLBUTamide.IV|TOLBUTamide.IV
C0366674|T201|COMP|4449-5|LNC|Tranylcypromine|Tranylcypromine
C0366675|T201|COMP|4450-3|LNC|traZODone|traZODone
C0366676|T201|COMP|4451-1|LNC|Triamterene|Triamterene
C0366677|T201|COMP|4452-9|LNC|Triazolam|Triazolam
C0366678|T201|COMP|4453-7|LNC|Trimeperidine|Trimeperidine
C0366679|T201|COMP|4454-5|LNC|Trimethadione|Trimethadione
C0366680|T201|COMP|4455-2|LNC|Trimethoprim|Trimethoprim
C0366681|T201|COMP|4456-0|LNC|Trimipramine|Trimipramine
C0366682|T201|COMP|4457-8|LNC|Tripelennamine|Tripelennamine
C0366683|T201|COMP|4458-6|LNC|Valproate|Valproate
C0366687|T201|COMP|4462-8|LNC|Xylose.PO|Xylose.PO
C0366688|T201|COMP|4463-6|LNC|Motility & count panel|Motility & count panel
C0366691|T201|COMP|4466-9|LNC|Stain.vital|Stain.vital
C0366693|T201|COMP|4468-5|LNC|Carbonyl hemoglobin/Hemoglobin.total|Carbonyl hemoglobin/Hemoglobin.total
C0366694|T201|COMP|4469-3|LNC|Cellano Ag|Cellano Ag
C0366695|T201|COMP|4470-1|LNC|Choleglobin/Hemoglobin.total|Choleglobin/Hemoglobin.total
C0366696|T201|COMP|4471-9|LNC|Complement activity.cell surface induced|Complement activity.cell surface induced
C0366697|T201|COMP|4472-7|LNC|Complement C'2 esterase|Complement C'2 esterase
C0366698|T201|COMP|4473-5|LNC|Complement C'3 esterase|Complement C'3 esterase
C0366699|T201|COMP|4474-3|LNC|Complement C'4 esterase|Complement C'4 esterase
C0366700|T201|COMP|4475-0|LNC|Complement C1|Complement C1
C0366701|T201|COMP|4476-8|LNC|Complement C1 esterase inhibitor.functional|Complement C1 esterase inhibitor.functional
C0366702|T201|COMP|4477-6|LNC|Complement C1 esterase inhibitor|Complement C1 esterase inhibitor
C0366703|T201|COMP|4478-4|LNC|Complement C1q|Complement C1q
C0366704|T201|COMP|6297-6|LNC|Complement C1q Ag|Complement C1q Ag
C0366705|T201|COMP|4479-2|LNC|Complement C1q Ag|Complement C1q Ag
C0366706|T201|COMP|4480-0|LNC|Complement C1q binding|Complement C1q binding
C0366707|T201|COMP|4481-8|LNC|Complement C1r|Complement C1r
C0366708|T201|COMP|4482-6|LNC|Complement C1r2+C1s2|Complement C1r2+C1s2
C0366709|T201|COMP|4483-4|LNC|Complement C1s|Complement C1s
C0366710|T201|COMP|4484-2|LNC|Complement C2|Complement C2
C0366711|T201|COMP|4485-9|LNC|Complement C3|Complement C3
C0366712|T201|COMP|4486-7|LNC|Complement C3 fragment|Complement C3 fragment
C0366713|T201|COMP|4487-5|LNC|Complement C3 fragment|Complement C3 fragment
C0366714|T201|COMP|4488-3|LNC|Complement C3a|Complement C3a
C0366715|T201|COMP|4489-1|LNC|Complement C3b|Complement C3b
C0366716|T201|COMP|6296-8|LNC|Complement C3b-C4b receptor|Complement C3b-C4b receptor
C0366717|T201|COMP|4490-9|LNC|Complement C3b-C4b receptor|Complement C3b-C4b receptor
C0366718|T201|COMP|4491-7|LNC|Complement C3c|Complement C3c
C0366719|T201|COMP|6295-0|LNC|Complement C3d|Complement C3d
C0366720|T201|COMP|4492-5|LNC|Complement C3d|Complement C3d
C0366721|T201|COMP|4493-3|LNC|Complement C3d+G|Complement C3d+G
C0366722|T201|COMP|4494-1|LNC|Complement C3d+G|Complement C3d+G
C0366723|T201|COMP|4495-8|LNC|Complement C3d+G|Complement C3d+G
C0366724|T201|COMP|4496-6|LNC|Complement C3d-C3d+Gg-IC3b receptors|Complement C3d-C3d+Gg-IC3b receptors
C0366725|T201|COMP|6294-3|LNC|Complement C3d-C3d+Gg-IC3b receptors|Complement C3d-C3d+Gg-IC3b receptors
C0366726|T201|COMP|4497-4|LNC|Complement C3PA|Complement C3PA
C0366727|T201|COMP|4498-2|LNC|Complement C4|Complement C4
C0366728|T201|COMP|4499-0|LNC|Complement C4 activated|Complement C4 activated
C0366729|T201|COMP|4500-5|LNC|Complement C4 CH50|Complement C4 CH50
C0366730|T201|COMP|4501-3|LNC|Complement C4a|Complement C4a
C0366731|T201|COMP|4502-1|LNC|Complement C4b binding protein|Complement C4b binding protein
C0366732|T201|COMP|4503-9|LNC|Complement C4b binding protein|Complement C4b binding protein
C0366733|T201|COMP|6293-5|LNC|Complement C4d|Complement C4d
C0366734|T201|COMP|4504-7|LNC|Complement C4d|Complement C4d
C0366735|T201|COMP|4505-4|LNC|Complement C5|Complement C5
C0366736|T201|COMP|4506-2|LNC|Complement C5a|Complement C5a
C0366737|T201|COMP|4507-0|LNC|Complement C6|Complement C6
C0366738|T201|COMP|4508-8|LNC|Complement C7|Complement C7
C0366739|T201|COMP|4509-6|LNC|Complement C8|Complement C8
C0366740|T201|COMP|4510-4|LNC|Complement C9|Complement C9
C0366741|T201|COMP|4512-0|LNC|Complement CH50|Complement CH50
C0366742|T201|COMP|4513-8|LNC|Complement C1r2+C1s2|Complement C1r2+C1s2
C0366743|T201|COMP|6292-7|LNC|Complement decay accelerating factor|Complement decay accelerating factor
C0366744|T201|COMP|4514-6|LNC|Complement decay accelerating factor|Complement decay accelerating factor
C0366745|T201|COMP|4515-3|LNC|Complement factor B|Complement factor B
C0366746|T201|COMP|4516-1|LNC|Complement factor Ba|Complement factor Ba
C0366747|T201|COMP|4517-9|LNC|Complement factor Bb|Complement factor Bb
C0366748|T201|COMP|4518-7|LNC|Complement factor D|Complement factor D
C0366749|T201|COMP|4519-5|LNC|Complement factor H|Complement factor H
C0366750|T201|COMP|4520-3|LNC|Complement factor I|Complement factor I
C0366751|T201|COMP|4521-1|LNC|Complement factor P|Complement factor P
C0366752|T201|COMP|4522-9|LNC|Complement iC3|Complement iC3
C0366753|T201|COMP|6291-9|LNC|Complement iC3b receptors|Complement iC3b receptors
C0366754|T201|COMP|4523-7|LNC|Complement iC3b receptors|Complement iC3b receptors
C0366756|T201|COMP|6290-1|LNC|Complement membrane C3b-C4b cofactor protein|Complement membrane C3b-C4b cofactor protein
C0366757|T201|COMP|4525-2|LNC|Complement membrane C3b-C4b cofactor protein|Complement membrane C3b-C4b cofactor protein
C0366758|T201|COMP|4526-0|LNC|Complement protein|Complement protein
C0366759|T201|COMP|4527-8|LNC|Complement receptor 1|Complement receptor 1
C0366760|T201|COMP|4528-6|LNC|Complement receptor 2|Complement receptor 2
C0366761|T201|COMP|4529-4|LNC|Complement receptor 3|Complement receptor 3
C0366762|T201|COMP|4530-2|LNC|Complement receptor 4|Complement receptor 4
C0366763|T201|COMP|4531-0|LNC|Complement total hemolytic|Complement total hemolytic
C0366764|T201|COMP|4511-2|LNC|Complement total hemolytic CH50|Complement total hemolytic CH50
C0366766|T201|COMP|4533-6|LNC|Complement+Immunoglobulin|Complement+Immunoglobulin
C0366767|T201|COMP|4534-4|LNC|Cyanmethemoglobin/Hemoglobin.total|Cyanmethemoglobin/Hemoglobin.total
C0366768|T201|COMP|4535-1|LNC|Cytotoxic percent reactive Ab|Cytotoxic percent reactive Ab
C0366769|T201|COMP|4536-9|LNC|Deoxyhemoglobin/Hemoglobin.total|Deoxyhemoglobin/Hemoglobin.total
C0366770|T201|COMP|4537-7|LNC|Erythrocyte sedimentation rate|Erythrocyte sedimentation rate
C0366771|T201|COMP|4538-5|LNC|Erythrocyte sedimentation rate|Erythrocyte sedimentation rate
C0366772|T201|COMP|4539-3|LNC|Erythrocyte sedimentation rate.Zeta|Erythrocyte sedimentation rate.Zeta
C0366773|T201|COMP|4540-1|LNC|Ethanol gelation|Ethanol gelation
C0366774|T201|COMP|4541-9|LNC|Euglobulin clot lysis|Euglobulin clot lysis
C0366775|T201|COMP|4542-7|LNC|Haptoglobin|Haptoglobin
C0366776|T201|COMP|4543-5|LNC|Haptoglobin|Haptoglobin
C0366777|T201|COMP|4544-3|LNC|Hematocrit|Hematocrit
C0366778|T201|COMP|4545-0|LNC|Hematocrit|Hematocrit
C0366779|T201|COMP|4546-8|LNC|Hemoglobin A/Hemoglobin.total|Hemoglobin A/Hemoglobin.total
C0366780|T201|COMP|4547-6|LNC|Hemoglobin A1/Hemoglobin.total|Hemoglobin A1/Hemoglobin.total
C0366781|T201|COMP|4548-4|LNC|Hemoglobin A1c/Hemoglobin.total|Hemoglobin A1c/Hemoglobin.total
C0366782|T201|COMP|4549-2|LNC|Hemoglobin A1c/Hemoglobin.total|Hemoglobin A1c/Hemoglobin.total
C0366783|T201|COMP|4550-0|LNC|Hemoglobin A2|Hemoglobin A2
C0366784|T201|COMP|4551-8|LNC|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C0366785|T201|COMP|4552-6|LNC|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C0366786|T201|COMP|4553-4|LNC|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C0366787|T201|COMP|4554-2|LNC|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C0366788|T201|COMP|4555-9|LNC|Hemoglobin A3/Hemoglobin.total|Hemoglobin A3/Hemoglobin.total
C0366789|T201|COMP|4556-7|LNC|Hemoglobin Abruzzo|Hemoglobin Abruzzo
C0366790|T201|COMP|4557-5|LNC|Hemoglobin Abruzzo|Hemoglobin Abruzzo
C0366791|T201|COMP|4558-3|LNC|Hemoglobin Barts|Hemoglobin Barts
C0366792|T201|COMP|4559-1|LNC|Hemoglobin Barts|Hemoglobin Barts
C0366793|T201|COMP|4560-9|LNC|Hemoglobin Bethesda|Hemoglobin Bethesda
C0366794|T201|COMP|4563-3|LNC|Hemoglobin C/Hemoglobin.total|Hemoglobin C/Hemoglobin.total
C0366795|T201|COMP|4561-7|LNC|Hemoglobin C/Hemoglobin.total|Hemoglobin C/Hemoglobin.total
C0366796|T201|COMP|4562-5|LNC|Hemoglobin C/Hemoglobin.total|Hemoglobin C/Hemoglobin.total
C0366797|T201|COMP|4564-1|LNC|Hemoglobin C-Harlem|Hemoglobin C-Harlem
C0366798|T201|COMP|4565-8|LNC|Hemoglobin Chesapeake|Hemoglobin Chesapeake
C0366799|T201|COMP|4566-6|LNC|Hemoglobin Chesapeake|Hemoglobin Chesapeake
C0366800|T201|COMP|4567-4|LNC|Hemoglobin Constant Spring|Hemoglobin Constant Spring
C0366801|T201|COMP|4568-2|LNC|Hemoglobin Constant Spring|Hemoglobin Constant Spring
C0366802|T201|COMP|4569-0|LNC|Hemoglobin D/Hemoglobin.total|Hemoglobin D/Hemoglobin.total
C0366803|T201|COMP|4571-6|LNC|Hemoglobin D-Punjab|Hemoglobin D-Punjab
C0366804|T201|COMP|4570-8|LNC|Hemoglobin D-Punjab|Hemoglobin D-Punjab
C0366805|T201|COMP|4572-4|LNC|Hemoglobin Denver|Hemoglobin Denver
C0366806|T201|COMP|4575-7|LNC|Hemoglobin E/Hemoglobin.total|Hemoglobin E/Hemoglobin.total
C0366807|T201|COMP|4573-2|LNC|Hemoglobin E/Hemoglobin.total|Hemoglobin E/Hemoglobin.total
C0366808|T201|COMP|4574-0|LNC|Hemoglobin E/Hemoglobin.total|Hemoglobin E/Hemoglobin.total
C0366809|T201|COMP|5913-9|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C0366810|T201|COMP|4632-6|LNC|Hemoglobin F|Hemoglobin F
C0366811|T201|COMP|4633-4|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C0366812|T201|COMP|4576-5|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C0366813|T201|COMP|4578-1|LNC|Hemoglobin F-Texas|Hemoglobin F-Texas
C0366814|T201|COMP|4577-3|LNC|Hemoglobin F-Texas|Hemoglobin F-Texas
C0366815|T201|COMP|4579-9|LNC|Hemoglobin F|Hemoglobin F
C0366816|T201|COMP|4580-7|LNC|Hemoglobin F1/Hemoglobin.total|Hemoglobin F1/Hemoglobin.total
C0366817|T201|COMP|4582-3|LNC|Hemoglobin G-Coushatta|Hemoglobin G-Coushatta
C0366818|T201|COMP|4581-5|LNC|Hemoglobin G-Coushatta|Hemoglobin G-Coushatta
C0366819|T201|COMP|4583-1|LNC|Hemoglobin G-Georgia|Hemoglobin G-Georgia
C0366820|T201|COMP|4584-9|LNC|Hemoglobin G-Georgia|Hemoglobin G-Georgia
C0366821|T201|COMP|4585-6|LNC|Hemoglobin G-Philadelphia|Hemoglobin G-Philadelphia
C0366822|T201|COMP|4586-4|LNC|Hemoglobin G-Philadelphia|Hemoglobin G-Philadelphia
C0366823|T201|COMP|4587-2|LNC|Hemoglobin H/Hemoglobin.total|Hemoglobin H/Hemoglobin.total
C0366824|T201|COMP|4588-0|LNC|Hemoglobin H/Hemoglobin.total|Hemoglobin H/Hemoglobin.total
C0366825|T201|COMP|4589-8|LNC|Hemoglobin Hasharon|Hemoglobin Hasharon
C0366826|T201|COMP|4590-6|LNC|Hemoglobin Hasharon|Hemoglobin Hasharon
C0366827|T201|COMP|4591-4|LNC|Hemoglobin Hope|Hemoglobin Hope
C0366828|T201|COMP|4592-2|LNC|Hemoglobin Hope|Hemoglobin Hope
C0366829|T201|COMP|4593-0|LNC|Hemoglobin I|Hemoglobin I
C0366830|T201|COMP|4594-8|LNC|Hemoglobin I|Hemoglobin I
C0366831|T201|COMP|4595-5|LNC|Hemoglobin J-Baltimore|Hemoglobin J-Baltimore
C0366832|T201|COMP|4596-3|LNC|Hemoglobin J-Baltimore|Hemoglobin J-Baltimore
C0366833|T201|COMP|4597-1|LNC|Hemoglobin J-Capetown|Hemoglobin J-Capetown
C0366834|T201|COMP|4598-9|LNC|Hemoglobin J-Oxford|Hemoglobin J-Oxford
C0366835|T201|COMP|4599-7|LNC|Hemoglobin J-Oxford|Hemoglobin J-Oxford
C0366836|T201|COMP|4600-3|LNC|Hemoglobin Kansas|Hemoglobin Kansas
C0366837|T201|COMP|4601-1|LNC|Hemoglobin Kempsey|Hemoglobin Kempsey
C0366838|T201|COMP|4602-9|LNC|Hemoglobin Kempsey|Hemoglobin Kempsey
C0366839|T201|COMP|4603-7|LNC|Hemoglobin Koln|Hemoglobin Koln
C0366840|T201|COMP|4604-5|LNC|Hemoglobin Lepore|Hemoglobin Lepore
C0366841|T201|COMP|4605-2|LNC|Hemoglobin Lepore|Hemoglobin Lepore
C0366842|T201|COMP|4606-0|LNC|Hemoglobin M-Boston|Hemoglobin M-Boston
C0366843|T201|COMP|4607-8|LNC|Hemoglobin M-Hyde park|Hemoglobin M-Hyde park
C0366844|T201|COMP|4608-6|LNC|Hemoglobin M-Iwate|Hemoglobin M-Iwate
C0366845|T201|COMP|4609-4|LNC|Hemoglobin M-Milwaukee|Hemoglobin M-Milwaukee
C0366846|T201|COMP|4610-2|LNC|Hemoglobin M-Saskatoon|Hemoglobin M-Saskatoon
C0366847|T201|COMP|4611-0|LNC|Hemoglobin Malmo|Hemoglobin Malmo
C0366848|T201|COMP|4612-8|LNC|Hemoglobin Malmo|Hemoglobin Malmo
C0366849|T201|COMP|4613-6|LNC|Hemoglobin N-Baltimore|Hemoglobin N-Baltimore
C0366850|T201|COMP|4614-4|LNC|Hemoglobin N-Baltimore|Hemoglobin N-Baltimore
C0366851|T201|COMP|4615-1|LNC|Hemoglobin N-Seattle|Hemoglobin N-Seattle
C0366852|T201|COMP|4616-9|LNC|Hemoglobin N-Seattle|Hemoglobin N-Seattle
C0366853|T201|COMP|4617-7|LNC|Hemoglobin O-Arab|Hemoglobin O-Arab
C0366854|T201|COMP|4618-5|LNC|Hemoglobin O-Arab|Hemoglobin O-Arab
C0366855|T201|COMP|4619-3|LNC|Hemoglobin Ranier|Hemoglobin Ranier
C0366856|T201|COMP|4621-9|LNC|Hemoglobin S|Hemoglobin S
C0366857|T201|COMP|4622-7|LNC|Hemoglobin S|Hemoglobin S
C0366858|T201|COMP|4623-5|LNC|Hemoglobin S|Hemoglobin S
C0366859|T201|COMP|4624-3|LNC|Hemoglobin S|Hemoglobin S
C0366860|T201|COMP|4625-0|LNC|Hemoglobin S/Hemoglobin.total|Hemoglobin S/Hemoglobin.total
C0366861|T201|COMP|4626-8|LNC|Hemoglobin Yakima|Hemoglobin Yakima
C0366862|T201|COMP|4627-6|LNC|Hemoglobin Yoshizuka|Hemoglobin Yoshizuka
C0366863|T201|COMP|4628-4|LNC|Hemoglobin Ypsilanti|Hemoglobin Ypsilanti
C0366864|T201|COMP|4629-2|LNC|Hemoglobin Zurich|Hemoglobin Zurich
C0366865|T201|COMP|4630-0|LNC|Hemoglobin Zurich|Hemoglobin Zurich
C0366866|T201|COMP|4631-8|LNC|Hemoglobin F|Hemoglobin F
C0366867|T201|COMP|4634-2|LNC|Hemoglobin.fetal|Hemoglobin.fetal
C0366869|T201|COMP|4636-7|LNC|Hemoglobin.free|Hemoglobin.free
C0366870|T201|COMP|4637-5|LNC|Hemoglobin.glycated|Hemoglobin.glycated
C0366871|T201|COMP|4638-3|LNC|Hemoglobin.thermolabile/Hemoglobin.total|Hemoglobin.thermolabile/Hemoglobin.total
C0366872|T201|COMP|4639-1|LNC|Hemoglobin.unstable|Hemoglobin.unstable
C0366873|T201|COMP|4640-9|LNC|Hemolysin.cold|Hemolysin.cold
C0366874|T201|COMP|4641-7|LNC|Hemolysin.warm|Hemolysin.warm
C0366875|T201|COMP|2403-4|LNC|Hemopexin|Hemopexin
C0366876|T201|COMP|4643-3|LNC|Hemosiderin|Hemosiderin
C0366877|T201|COMP|4645-8|LNC|Hemosiderin|Hemosiderin
C0366878|T201|COMP|4644-1|LNC|Hemosiderin|Hemosiderin
C0366879|T201|COMP|4646-6|LNC|Heparin|Heparin
C0366880|T201|COMP|4647-4|LNC|Heparin|Heparin
C0366881|T201|COMP|4648-2|LNC|Homologous restriction factor|Homologous restriction factor
C0366882|T201|COMP|4649-0|LNC|Interferon|Interferon
C0366883|T201|COMP|4650-8|LNC|Interleukin 1|Interleukin 1
C0366884|T201|COMP|4651-6|LNC|Interleukin 2|Interleukin 2
C0366885|T201|COMP|4652-4|LNC|Interleukin 3|Interleukin 3
C0366886|T201|COMP|4653-2|LNC|Interleukin 4|Interleukin 4
C0366887|T201|COMP|4654-0|LNC|Interleukin 5|Interleukin 5
C0366888|T201|COMP|4655-7|LNC|Interleukin 6|Interleukin 6
C0366889|T201|COMP|4656-5|LNC|Interleukin 7|Interleukin 7
C0366890|T201|COMP|4657-3|LNC|Kallikrein|Kallikrein
C0366891|T201|COMP|4658-1|LNC|Kallikrein.tissue type|Kallikrein.tissue type
C0366892|T201|COMP|4659-9|LNC|Phosphatase.leukocyte|Phosphatase.leukocyte
C0366893|T201|COMP|4660-7|LNC|Leukocyte.detection Ab|Leukocyte.detection Ab
C0366894|T201|COMP|4661-5|LNC|Lupus erythematosus factor|Lupus erythematosus factor
C0366896|T201|COMP|4663-1|LNC|Lymphocytotoxicity|Lymphocytotoxicity
C0366897|T201|COMP|4664-9|LNC|Lymphocytotoxicity|Lymphocytotoxicity
C0366898|T201|COMP|4665-6|LNC|Lysozyme|Lysozyme
C0366899|T201|COMP|6289-3|LNC|Lysozyme|Lysozyme
C0366900|T201|COMP|4667-2|LNC|Osmotic fragility|Osmotic fragility
C0366901|T201|COMP|4666-4|LNC|Osmotic fragility|Osmotic fragility
C0366902|T201|COMP|4668-0|LNC|Plasminogen Ag|Plasminogen Ag
C0366903|T201|COMP|4669-8|LNC|Prekallikrein|Prekallikrein
C0366904|T201|COMP|4670-6|LNC|Thrombomodulin factor B|Thrombomodulin factor B
C0366905|T201|COMP|4671-4|LNC|Protein C|Protein C
C0366906|T201|COMP|4672-2|LNC|Protein C Ag|Protein C Ag
C0366907|T201|COMP|4674-8|LNC|Protein C inhibitor.activated|Protein C inhibitor.activated
C0366908|T201|COMP|4679-7|LNC|Reticulocytes/100 erythrocytes|Reticulocytes/100 erythrocytes
C0366909|T201|COMP|4680-5|LNC|von Willebrand factor.ristocetin cofactor|von Willebrand factor.ristocetin cofactor
C0366910|T201|COMP|4681-3|LNC|Streptokinase|Streptokinase
C0366911|T201|COMP|4682-1|LNC|Streptokinase|Streptokinase
C0366912|T201|COMP|4684-7|LNC|Sulfhemoglobin|Sulfhemoglobin
C0366913|T201|COMP|4683-9|LNC|Sulfhemoglobin|Sulfhemoglobin
C0366914|T201|COMP|4685-4|LNC|Sulfhemoglobin/Hemoglobin.total|Sulfhemoglobin/Hemoglobin.total
C0366915|T201|COMP|4686-2|LNC|Thromboglobulin|Thromboglobulin
C0366916|T201|COMP|4687-0|LNC|Thromboglobulin beta|Thromboglobulin beta
C0366917|T201|COMP|4688-8|LNC|Thrombomodulin|Thrombomodulin
C0366918|T201|COMP|4689-6|LNC|Verdohemoglobin|Verdohemoglobin
C0366919|T201|COMP|4691-2|LNC|Viscosity|Viscosity
C0366920|T201|COMP|4692-0|LNC|HLA Ag|HLA Ag
C0366921|T201|COMP|4693-8|LNC|HLA Ag absent|HLA Ag absent
C0366922|T201|COMP|4694-6|LNC|HLA Ag present|HLA Ag present
C0367218|T201|COMP|5227-4|LNC|Streptococcal hyaluronidase Ab|Streptococcal hyaluronidase Ab
C0367219|T201|COMP|632-0|LNC|Bacteria identified|Bacteria identified
C0367220|T201|COMP|581-9|LNC|Streptococcus agalactiae|Streptococcus agalactiae
C0367221|T201|COMP|582-7|LNC|Streptococcus agalactiae|Streptococcus agalactiae
C0367222|T201|COMP|583-5|LNC|Streptococcus agalactiae|Streptococcus agalactiae
C0367223|T201|COMP|584-3|LNC|Streptococcus agalactiae|Streptococcus agalactiae
C0367224|T201|COMP|585-0|LNC|Streptococcus agalactiae|Streptococcus agalactiae
C0367225|T201|COMP|586-8|LNC|Streptococcus agalactiae|Streptococcus agalactiae
C0367226|T201|COMP|6551-6|LNC|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C0367227|T201|COMP|5034-4|LNC|Streptococcus agalactiae rRNA|Streptococcus agalactiae rRNA
C0367228|T201|COMP|6552-4|LNC|Streptococcus pneumoniae Ab|Streptococcus pneumoniae Ab
C0367229|T201|COMP|5368-6|LNC|Streptococcus pneumoniae Ab.IgG|Streptococcus pneumoniae Ab.IgG
C0367230|T201|COMP|6553-2|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C0367231|T201|COMP|6554-0|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C0367232|T201|COMP|6555-7|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C0367233|T201|COMP|5035-1|LNC|Streptococcus pneumoniae rRNA|Streptococcus pneumoniae rRNA
C0367234|T201|COMP|633-8|LNC|Bacteria identified|Bacteria identified
C0367235|T201|COMP|6462-6|LNC|Bacteria identified|Bacteria identified
C0367236|T201|COMP|6556-5|LNC|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C0367237|T201|COMP|634-6|LNC|Bacteria identified|Bacteria identified
C0367238|T201|COMP|635-3|LNC|Bacteria identified|Bacteria identified
C0367239|T201|COMP|6557-3|LNC|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C0367240|T201|COMP|6558-1|LNC|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C0367241|T201|COMP|6559-9|LNC|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C0367242|T201|COMP|5173-0|LNC|Streptococcus pyogenes enzyme Ab|Streptococcus pyogenes enzyme Ab
C0367243|T201|COMP|5172-2|LNC|Streptococcus pyogenes enzyme Ab|Streptococcus pyogenes enzyme Ab
C0367244|T201|COMP|6463-4|LNC|Bacteria identified|Bacteria identified
C0367245|T201|COMP|5036-9|LNC|Streptococcus pyogenes rRNA|Streptococcus pyogenes rRNA
C0367246|T201|COMP|546-2|LNC|Streptococcus.beta-hemolytic|Streptococcus.beta-hemolytic
C0367247|T201|COMP|547-0|LNC|Streptococcus.beta-hemolytic|Streptococcus.beta-hemolytic
C0367248|T201|COMP|5369-4|LNC|Streptokinase Ab|Streptokinase Ab
C0367249|T201|COMP|636-1|LNC|Bacteria identified|Bacteria identified
C0367250|T201|COMP|5370-2|LNC|Streptolysin O Ab|Streptolysin O Ab
C0367251|T201|COMP|5371-0|LNC|Streptolysin O Ab|Streptolysin O Ab
C0367252|T201|COMP|5246-4|LNC|Saccharopolyspora rectivirgula Ab|Saccharopolyspora rectivirgula Ab
C0367253|T201|COMP|5373-6|LNC|Strongyloides sp Ab|Strongyloides sp Ab
C0367254|T201|COMP|5374-4|LNC|Taenia saginata Ab|Taenia saginata Ab
C0367255|T201|COMP|5375-1|LNC|Taenia solium adult Ab|Taenia solium adult Ab
C0367256|T201|COMP|637-9|LNC|Plasmodium sp identified|Plasmodium sp identified
C0367257|T201|COMP|5376-9|LNC|Thermoactinomyces candidus Ab|Thermoactinomyces candidus Ab
C0367260|T201|COMP|5377-7|LNC|Thermoactinomyces sacchari Ab|Thermoactinomyces sacchari Ab
C0367264|T201|COMP|5378-5|LNC|Thermoactinomyces vulgaris Ab|Thermoactinomyces vulgaris Ab
C0367265|T201|COMP|5386-8|LNC|Toxocara canis Ab|Toxocara canis Ab
C0367266|T201|COMP|5387-6|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C0367268|T201|COMP|5388-4|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0367269|T201|COMP|5389-2|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0367271|T201|COMP|5390-0|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0367273|T201|COMP|5391-8|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0367275|T201|COMP|6580-7|LNC|Treponema identified|Treponema identified
C0367278|T201|COMP|5392-6|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0367281|T201|COMP|5393-4|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0367282|T201|COMP|5394-2|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0367283|T201|COMP|6561-5|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C0367284|T201|COMP|6562-3|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C0367286|T201|COMP|5395-9|LNC|Trichinella spiralis Ab|Trichinella spiralis Ab
C0367287|T201|COMP|6563-1|LNC|Trichinella spiralis Ab.IgG|Trichinella spiralis Ab.IgG
C0367288|T201|COMP|6564-9|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C0367289|T201|COMP|6565-6|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C0367297|T201|COMP|6566-4|LNC|Trichomonas vaginalis Ag|Trichomonas vaginalis Ag
C0367299|T201|COMP|6567-2|LNC|Trichomonas vaginalis Ag|Trichomonas vaginalis Ag
C0367301|T201|COMP|6568-0|LNC|Trichomonas vaginalis rRNA|Trichomonas vaginalis rRNA
C0367302|T201|COMP|5397-5|LNC|Trypanosoma brucei Ab|Trypanosoma brucei Ab
C0367303|T201|COMP|5398-3|LNC|Trypanosoma cruzi Ab|Trypanosoma cruzi Ab
C0367304|T201|COMP|5399-1|LNC|Trypanosoma sp Ab|Trypanosoma sp Ab
C0367305|T201|COMP|5400-7|LNC|Vaccinia virus Ab|Vaccinia virus Ab
C0367306|T201|COMP|5401-5|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C0367307|T201|COMP|5402-3|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C0367308|T201|COMP|5403-1|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0367313|T201|COMP|6569-8|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0367314|T201|COMP|5404-9|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0367315|T201|COMP|6570-6|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0367316|T201|COMP|5881-8|LNC|Varicella zoster virus Ag|Varicella zoster virus Ag
C0367317|T201|COMP|5882-6|LNC|Varicella zoster virus Ag|Varicella zoster virus Ag
C0367318|T201|COMP|6572-2|LNC|Venezuelan equine encephalitis virus Ag|Venezuelan equine encephalitis virus Ag
C0367320|T201|COMP|6571-4|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C0367321|T201|COMP|6573-0|LNC|Venezuelan equine encephalitis virus Ag|Venezuelan equine encephalitis virus Ag
C0367322|T201|COMP|6574-8|LNC|Escherichia coli verotoxin 1|Escherichia coli verotoxin 1
C0367329|T201|COMP|6576-3|LNC|Escherichia coli verotoxin 2|Escherichia coli verotoxin 2
C0367333|T201|COMP|5405-6|LNC|Vibrio cholerae Ab|Vibrio cholerae Ab
C0367334|T201|COMP|6578-9|LNC|Vibrio sp identified|Vibrio sp identified
C0367335|T201|COMP|6579-7|LNC|Vibrio sp identified|Vibrio sp identified
C0367345|T201|COMP|6580-5|LNC|Vibrio sp identified|Vibrio sp identified
C0367346|T201|COMP|6581-3|LNC|Vibrio sp identified|Vibrio sp identified
C0367350|T201|COMP|673-4|LNC|Ova & parasites identified|Ova & parasites identified
C0367351|T201|COMP|675-9|LNC|Enterobius vermicularis|Enterobius vermicularis
C0367356|T201|COMP|5883-4|LNC|Virus identified|Virus identified
C0367357|T201|COMP|5884-2|LNC|Virus identified|Virus identified
C0367359|T201|COMP|6583-9|LNC|Virus identified|Virus identified
C0367360|T201|COMP|5886-7|LNC|Virus identified|Virus identified
C0367361|T201|COMP|5885-9|LNC|Virus identified|Virus identified
C0367363|T201|COMP|5887-5|LNC|Virus identified|Virus identified
C0367364|T201|COMP|5888-3|LNC|Virus identified|Virus identified
C0367365|T201|COMP|17976-2|LNC|Virus identified^^^3|Virus identified^^^3
C0367366|T201|COMP|5406-4|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0367367|T201|COMP|6585-4|LNC|Western equine encephalitis virus Ag|Western equine encephalitis virus Ag
C0367368|T201|COMP|6586-2|LNC|Western equine encephalitis virus Ag|Western equine encephalitis virus Ag
C0367369|T201|COMP|6588-8|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C0367370|T201|COMP|6587-0|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C0367371|T201|COMP|6591-2|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C0367372|T201|COMP|6590-4|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C0367373|T201|COMP|6589-6|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C0367374|T201|COMP|6593-8|LNC|Yellow fever virus Ab.IgM|Yellow fever virus Ab.IgM
C0367375|T201|COMP|6592-0|LNC|Yellow fever virus Ab.IgG|Yellow fever virus Ab.IgG
C0367376|T201|COMP|5408-0|LNC|Yersinia enterocolitica O:8 Ab|Yersinia enterocolitica O:8 Ab
C0367377|T201|COMP|5407-2|LNC|Yersinia enterocolitica O:3 Ab|Yersinia enterocolitica O:3 Ab
C0367378|T201|COMP|5410-6|LNC|Yersinia pseudotuberculosis Ab|Yersinia pseudotuberculosis Ab
C0367379|T201|COMP|5409-8|LNC|Yersinia enterocolitica O:9 Ab|Yersinia enterocolitica O:9 Ab
C0367380|T201|COMP|701-3|LNC|Yersinia sp identified|Yersinia sp identified
C0367381|T201|COMP|5411-4|LNC|Yersinia sp Ab|Yersinia sp Ab
C0367382|T201|COMP|5037-7|LNC|Acetylcholine receptor binding Ab|Acetylcholine receptor binding Ab
C0367383|T201|COMP|5038-5|LNC|Acetylcholine receptor blocking Ab|Acetylcholine receptor blocking Ab
C0367385|T201|COMP|5039-3|LNC|Acetylcholine receptor modulation Ab|Acetylcholine receptor modulation Ab
C0367386|T201|COMP|5043-5|LNC|Adrenal Ab|Adrenal Ab
C0367387|T201|COMP|5044-3|LNC|Adrenal cortex Ab|Adrenal cortex Ab
C0367389|T201|COMP|6475-8|LNC|Mobiluncus sp rRNA|Mobiluncus sp rRNA
C0367390|T201|COMP|5248-0|LNC|Mucor sp Ab|Mucor sp Ab
C0367391|T201|COMP|5047-6|LNC|Nuclear Ab|Nuclear Ab
C0367392|T201|COMP|5249-8|LNC|Mumps virus Ab|Mumps virus Ab
C0367393|T201|COMP|5250-6|LNC|Mumps virus Ab|Mumps virus Ab
C0367394|T201|COMP|5048-4|LNC|Nuclear Ab|Nuclear Ab
C0367395|T201|COMP|5056-7|LNC|Basement membrane Ab|Basement membrane Ab
C0367396|T201|COMP|5076-5|LNC|Cardiolipin Ab.IgA|Cardiolipin Ab.IgA
C0367397|T201|COMP|5077-3|LNC|Centromere Ab|Centromere Ab
C0367398|T201|COMP|5091-4|LNC|Chymotrypsin Ab|Chymotrypsin Ab
C0367401|T201|COMP|5117-7|LNC|Cryoglobulin|Cryoglobulin
C0367402|T201|COMP|6476-6|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0367403|T201|COMP|6477-4|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0367404|T201|COMP|6478-2|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C0367405|T201|COMP|6479-0|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C0367406|T201|COMP|5022-9|LNC|Mycobacterium avium complex rRNA|Mycobacterium avium complex rRNA
C0367407|T201|COMP|6480-8|LNC|Mumps virus Ag|Mumps virus Ag
C0367408|T201|COMP|5023-7|LNC|Mycobacterium avium subspecies avium rRNA|Mycobacterium avium subspecies avium rRNA
C0367410|T201|COMP|5129-2|LNC|Deoxyribonuclease Ab|Deoxyribonuclease Ab
C0367411|T201|COMP|5130-0|LNC|DNA double strand Ab|DNA double strand Ab
C0367412|T201|COMP|5131-8|LNC|DNA double strand Ab|DNA double strand Ab
C0367413|T201|COMP|5132-6|LNC|DNA single strand Ab|DNA single strand Ab
C0367414|T201|COMP|5152-4|LNC|Epidermis Ab|Epidermis Ab
C0367415|T201|COMP|5161-5|LNC|Erythrocyte Ab|Erythrocyte Ab
C0367416|T201|COMP|5164-9|LNC|Fc fragment Ab|Fc fragment Ab
C0367417|T201|COMP|5168-0|LNC|Gall canaliculi Ab|Gall canaliculi Ab
C0367418|T201|COMP|5170-6|LNC|Gliadin Ab.IgG|Gliadin Ab.IgG
C0367419|T201|COMP|5024-5|LNC|Mycobacterium gordonae rRNA|Mycobacterium gordonae rRNA
C0367420|T201|COMP|532-2|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367421|T201|COMP|533-0|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367422|T201|COMP|534-8|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367423|T201|COMP|535-5|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367424|T201|COMP|536-3|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367426|T201|COMP|5217-5|LNC|Histone Ab|Histone Ab
C0367427|T201|COMP|5228-2|LNC|Immune complex|Immune complex
C0367428|T201|COMP|537-1|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367429|T201|COMP|538-9|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367430|T201|COMP|539-7|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367431|T201|COMP|540-5|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367432|T201|COMP|5232-4|LNC|Insulin Ab|Insulin Ab
C0367434|T201|COMP|5233-2|LNC|Intrinsic factor Ab|Intrinsic factor Ab
C0367435|T201|COMP|5247-2|LNC|Mitochondria Ab|Mitochondria Ab
C0367437|T201|COMP|5259-7|LNC|Myelin basic protein Ab|Myelin basic protein Ab
C0367438|T201|COMP|5251-4|LNC|Muscle sarcolemma Ab|Muscle sarcolemma Ab
C0367439|T201|COMP|542-1|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367440|T201|COMP|541-3|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367441|T201|COMP|5262-1|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C0367442|T201|COMP|5260-5|LNC|Myocardium Ab|Myocardium Ab
C0367443|T201|COMP|5025-2|LNC|Mycobacterium intracellulare rRNA|Mycobacterium intracellulare rRNA
C0367444|T201|COMP|543-9|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0367445|T201|COMP|5271-2|LNC|Parietal cell Ab|Parietal cell Ab
C0367446|T201|COMP|5265-4|LNC|Pancreatic islet cell Ab|Pancreatic islet cell Ab
C0367449|T201|COMP|5297-7|LNC|Rheumatoid factor|Rheumatoid factor
C0367450|T201|COMP|5296-9|LNC|Reticulin Ab|Reticulin Ab
C0367451|T201|COMP|5026-0|LNC|Mycobacterium kansasii rRNA|Mycobacterium kansasii rRNA
C0367452|T201|COMP|5298-5|LNC|Rheumatoid factor|Rheumatoid factor
C0367453|T201|COMP|5299-3|LNC|Rheumatoid factor|Rheumatoid factor
C0367454|T201|COMP|5027-8|LNC|Mycobacterium tuberculosis rRNA|Mycobacterium tuberculosis rRNA
C0367455|T201|COMP|5252-2|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C0367456|T201|COMP|5253-0|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C0367457|T201|COMP|5300-9|LNC|Rheumatoid factor|Rheumatoid factor
C0367460|T201|COMP|5337-1|LNC|Salivary gland Ab|Salivary gland Ab
C0367470|T201|COMP|5358-7|LNC|Smooth muscle Ab|Smooth muscle Ab
C0367471|T201|COMP|5359-5|LNC|Somatotropin Ab|Somatotropin Ab
C0367472|T201|COMP|5360-3|LNC|Spermatozoa Ab|Spermatozoa Ab
C0367474|T201|COMP|5362-9|LNC|Spermatozoa Ab|Spermatozoa Ab
C0367475|T201|COMP|5254-8|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C0367476|T201|COMP|5255-5|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C0367477|T201|COMP|6481-6|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C0367478|T201|COMP|5256-3|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C0367479|T201|COMP|5257-1|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C0367480|T201|COMP|5258-9|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C0367481|T201|COMP|5372-8|LNC|Striated muscle Ab|Striated muscle Ab
C0367484|T201|COMP|6482-4|LNC|Mycoplasma pneumoniae rRNA|Mycoplasma pneumoniae rRNA
C0367486|T201|COMP|5382-7|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C0367487|T201|COMP|6483-2|LNC|Mycoplasma pneumoniae rRNA|Mycoplasma pneumoniae rRNA
C0367488|T201|COMP|6484-0|LNC|Mycoplasma pneumoniae rRNA|Mycoplasma pneumoniae rRNA
C0367489|T201|COMP|5383-5|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C0367490|T201|COMP|5384-3|LNC|Thyrotropin Ab|Thyrotropin Ab
C0367491|T201|COMP|5385-0|LNC|Thyrotropin receptor Ab|Thyrotropin receptor Ab
C0367492|T201|COMP|5396-7|LNC|Triiodothyronine Ab|Triiodothyronine Ab
C0367493|T201|COMP|5412-2|LNC|B-B4|B-B4
C0367494|T201|COMP|5413-0|LNC|CD1|CD1
C0367495|T201|COMP|5414-8|LNC|CD10|CD10
C0367497|T201|COMP|5416-3|LNC|CD100|CD100
C0367498|T201|COMP|5417-1|LNC|CD102|CD102
C0367499|T201|COMP|6485-7|LNC|Mycoplasma pneumoniae rRNA|Mycoplasma pneumoniae rRNA
C0367500|T201|COMP|5418-9|LNC|CD103|CD103
C0367501|T201|COMP|5419-7|LNC|CD104|CD104
C0367502|T201|COMP|5420-5|LNC|CD105|CD105
C0367503|T201|COMP|6486-5|LNC|Mycoplasma sp identified|Mycoplasma sp identified
C0367504|T201|COMP|5421-3|LNC|CD106|CD106
C0367505|T201|COMP|683-3|LNC|Mycoplasma sp.genital identified|Mycoplasma sp.genital identified
C0367506|T201|COMP|684-1|LNC|Mycoplasma sp.respiratory identified|Mycoplasma sp.respiratory identified
C0367507|T201|COMP|685-8|LNC|Mycoplasma sp.respiratory identified|Mycoplasma sp.respiratory identified
C0367508|T201|COMP|5422-1|LNC|CD107a|CD107a
C0367509|T201|COMP|5423-9|LNC|CD107b|CD107b
C0367510|T201|COMP|686-6|LNC|Mycoplasma sp.respiratory identified|Mycoplasma sp.respiratory identified
C0367511|T201|COMP|687-4|LNC|Mycoplasma sp & Ureaplasma sp|Mycoplasma sp & Ureaplasma sp
C0367512|T201|COMP|688-2|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367513|T201|COMP|690-8|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367514|T201|COMP|5424-7|LNC|CD115|CD115
C0367515|T201|COMP|5425-4|LNC|CD117|CD117
C0367516|T201|COMP|5426-2|LNC|CD11a|CD11a
C0367517|T201|COMP|691-6|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367518|T201|COMP|5427-0|LNC|CD11b|CD11b
C0367519|T201|COMP|692-4|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367520|T201|COMP|5428-8|LNC|CD11c|CD11c
C0367521|T201|COMP|5429-6|LNC|CD120a|CD120a
C0367522|T201|COMP|5430-4|LNC|CD120b|CD120b
C0367523|T201|COMP|5431-2|LNC|CD122|CD122
C0367524|T201|COMP|5432-0|LNC|CD126|CD126
C0367525|T201|COMP|5433-8|LNC|CD128|CD128
C0367526|T201|COMP|5434-6|LNC|CD13|CD13
C0367527|T201|COMP|5435-3|LNC|CD14|CD14
C0367528|T201|COMP|5436-1|LNC|CD15|CD15
C0367529|T201|COMP|5437-9|LNC|CD16|CD16
C0367533|T201|COMP|5441-1|LNC|CD16-CD57-|CD16-CD57-
C0367534|T201|COMP|5442-9|LNC|CD16b|CD16b
C0367535|T201|COMP|5443-7|LNC|CD18|CD18
C0367536|T201|COMP|5444-5|LNC|CD19|CD19
C0367539|T201|COMP|693-2|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367540|T201|COMP|5447-8|LNC|CD2|CD2
C0367541|T201|COMP|5448-6|LNC|CD20|CD20
C0367542|T201|COMP|5449-4|LNC|CD21|CD21
C0367543|T201|COMP|5450-2|LNC|CD22|CD22
C0367545|T201|COMP|5452-8|LNC|CD23|CD23
C0367546|T201|COMP|5453-6|LNC|CD24|CD24
C0367547|T201|COMP|5454-4|LNC|CD25|CD25
C0367548|T201|COMP|5455-1|LNC|CD26|CD26
C0367549|T201|COMP|5456-9|LNC|CD27|CD27
C0367551|T201|COMP|5457-7|LNC|CD28|CD28
C0367552|T201|COMP|5458-5|LNC|CD29|CD29
C0367553|T201|COMP|5459-3|LNC|CD3|CD3
C0367555|T201|COMP|5461-9|LNC|CD30|CD30
C0367556|T201|COMP|5462-7|LNC|CD31|CD31
C0367557|T201|COMP|5463-5|LNC|CD32|CD32
C0367558|T201|COMP|5464-3|LNC|CD33|CD33
C0367560|T201|COMP|5467-6|LNC|CD35|CD35
C0367561|T201|COMP|5465-0|LNC|CD34|CD34
C0367562|T201|COMP|695-7|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367563|T201|COMP|5468-4|LNC|CD36|CD36
C0367564|T201|COMP|5469-2|LNC|CD37|CD37
C0367565|T201|COMP|5470-0|LNC|CD38|CD38
C0367566|T201|COMP|5471-8|LNC|CD39|CD39
C0367567|T201|COMP|5472-6|LNC|CD4|CD4
C0367569|T201|COMP|5474-2|LNC|CD4/CD8 ratio|CD4/CD8 ratio
C0367570|T201|COMP|5475-9|LNC|CD40|CD40
C0367571|T201|COMP|5476-7|LNC|CD41|CD41
C0367572|T201|COMP|5477-5|LNC|CD42a|CD42a
C0367573|T201|COMP|5478-3|LNC|CD42b|CD42b
C0367574|T201|COMP|5479-1|LNC|CD42c|CD42c
C0367575|T201|COMP|5480-9|LNC|CD42d|CD42d
C0367576|T201|COMP|5481-7|LNC|CD43|CD43
C0367577|T201|COMP|5482-5|LNC|CD44|CD44
C0367578|T201|COMP|5483-3|LNC|CD44R|CD44R
C0367579|T201|COMP|5484-1|LNC|CD45|CD45
C0367580|T201|COMP|5485-8|LNC|CD45RA|CD45RA
C0367581|T201|COMP|5486-6|LNC|CD45RB|CD45RB
C0367582|T201|COMP|5487-4|LNC|CD45RO|CD45RO
C0367583|T201|COMP|5488-2|LNC|CD46|CD46
C0367584|T201|COMP|697-3|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367585|T201|COMP|5489-0|LNC|CD47|CD47
C0367586|T201|COMP|5490-8|LNC|CD48|CD48
C0367587|T201|COMP|696-5|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367588|T201|COMP|5491-6|LNC|CD49a|CD49a
C0367589|T201|COMP|698-1|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367590|T201|COMP|5493-2|LNC|CD49c|CD49c
C0367591|T201|COMP|5261-3|LNC|Neisseria gonorrhoeae Ab|Neisseria gonorrhoeae Ab
C0367592|T201|COMP|5492-4|LNC|CD49B|CD49B
C0367593|T201|COMP|6487-3|LNC|Neisseria gonorrhoeae Ag|Neisseria gonorrhoeae Ag
C0367594|T201|COMP|5494-0|LNC|CD49d|CD49d
C0367595|T201|COMP|5495-7|LNC|CD49E|CD49E
C0367596|T201|COMP|5496-5|LNC|CD49f|CD49f
C0367597|T201|COMP|5497-3|LNC|CD5|CD5
C0367599|T201|COMP|5499-9|LNC|CD50|CD50
C0367600|T201|COMP|5500-4|LNC|CD51|CD51
C0367601|T201|COMP|5501-2|LNC|CD52|CD52
C0367602|T201|COMP|5502-0|LNC|CD53|CD53
C0367603|T201|COMP|5503-8|LNC|CD54|CD54
C0367604|T201|COMP|6488-1|LNC|Neisseria gonorrhoeae Ag|Neisseria gonorrhoeae Ag
C0367605|T201|COMP|6489-9|LNC|Neisseria gonorrhoeae Ag|Neisseria gonorrhoeae Ag
C0367606|T201|COMP|6490-7|LNC|Neisseria gonorrhoeae Ag|Neisseria gonorrhoeae Ag
C0367607|T201|COMP|5028-6|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C0367608|T201|COMP|5504-6|LNC|CD55|CD55
C0367609|T201|COMP|5505-3|LNC|CD56|CD56
C0367610|T201|COMP|5506-1|LNC|CD57|CD57
C0367611|T201|COMP|5507-9|LNC|CD58|CD58
C0367612|T201|COMP|5508-7|LNC|CD59|CD59
C0367613|T201|COMP|5509-5|LNC|CD6|CD6
C0367614|T201|COMP|5510-3|LNC|CD61|CD61
C0367615|T201|COMP|6492-3|LNC|Neisseria meningitidis Ag|Neisseria meningitidis Ag
C0367616|T201|COMP|6493-1|LNC|Neisseria meningitidis serogroup A Ag|Neisseria meningitidis serogroup A Ag
C0367617|T201|COMP|6494-9|LNC|Neisseria meningitidis serogroup A Ag|Neisseria meningitidis serogroup A Ag
C0367618|T201|COMP|6495-6|LNC|Neisseria meningitidis serogroup A Ag|Neisseria meningitidis serogroup A Ag
C0367619|T201|COMP|6496-4|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C0367620|T201|COMP|6497-2|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C0367621|T201|COMP|6498-0|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C0367622|T201|COMP|6499-8|LNC|Neisseria meningitidis serogroup C Ag|Neisseria meningitidis serogroup C Ag
C0367623|T201|COMP|6500-3|LNC|Neisseria meningitidis serogroup C Ag|Neisseria meningitidis serogroup C Ag
C0367624|T201|COMP|5511-1|LNC|CD62E|CD62E
C0367625|T201|COMP|5512-9|LNC|CD62L|CD62L
C0367626|T201|COMP|5513-7|LNC|CD62P|CD62P
C0367627|T201|COMP|5514-5|LNC|CD63|CD63
C0367628|T201|COMP|5515-2|LNC|CD64|CD64
C0367629|T201|COMP|5516-0|LNC|CD66a|CD66a
C0367630|T201|COMP|6501-1|LNC|Neisseria meningitidis serogroup C Ag|Neisseria meningitidis serogroup C Ag
C0367631|T201|COMP|6502-9|LNC|Neisseria meningitidis serogroup Y Ab|Neisseria meningitidis serogroup Y Ab
C0367632|T201|COMP|5517-8|LNC|CD66b|CD66b
C0367633|T201|COMP|5518-6|LNC|CD66c|CD66c
C0367634|T201|COMP|6503-7|LNC|Neisseria meningitidis serogroup Y Ag|Neisseria meningitidis serogroup Y Ag
C0367635|T201|COMP|6504-5|LNC|Neisseria meningitidis serogroup Y Ag|Neisseria meningitidis serogroup Y Ag
C0367636|T201|COMP|6505-2|LNC|Neisseria meningitidis serogroup Y Ag|Neisseria meningitidis serogroup Y Ag
C0367637|T201|COMP|6506-0|LNC|Neisseria meningitidis serogroup w135 Ag|Neisseria meningitidis serogroup w135 Ag
C0367638|T201|COMP|5519-4|LNC|CD66d|CD66d
C0367639|T201|COMP|6507-8|LNC|Neisseria meningitidis serogroup w135 Ag|Neisseria meningitidis serogroup w135 Ag
C0367640|T201|COMP|5520-2|LNC|CD66e|CD66e
C0367641|T201|COMP|5521-0|LNC|CD68|CD68
C0367642|T201|COMP|5522-8|LNC|CD69|CD69
C0367643|T201|COMP|5523-6|LNC|CD7|CD7
C0367645|T201|COMP|6508-6|LNC|Neisseria meningitidis Ag|Neisseria meningitidis Ag
C0367646|T201|COMP|6509-4|LNC|Neisseria meningitidis rRNA|Neisseria meningitidis rRNA
C0367647|T201|COMP|5525-1|LNC|CD71|CD71
C0367648|T201|COMP|5526-9|LNC|CD72|CD72
C0367649|T201|COMP|5527-7|LNC|CD73|CD73
C0367650|T201|COMP|5029-4|LNC|Neisseria meningitidis rRNA|Neisseria meningitidis rRNA
C0367651|T201|COMP|5263-9|LNC|Nocardia sp Ab|Nocardia sp Ab
C0367652|T201|COMP|5264-7|LNC|Onchocerca sp Ab|Onchocerca sp Ab
C0367653|T201|COMP|699-9|LNC|Organism count|Organism count
C0367654|T201|COMP|5528-5|LNC|CD74|CD74
C0367655|T201|COMP|5529-3|LNC|CD77|CD77
C0367656|T201|COMP|6510-2|LNC|Human papilloma virus Ab|Human papilloma virus Ab
C0367657|T201|COMP|5530-1|LNC|CD79a|CD79a
C0367658|T201|COMP|6511-0|LNC|Human papilloma virus Ab|Human papilloma virus Ab
C0367659|T201|COMP|5531-9|LNC|CD79b|CD79b
C0367660|T201|COMP|6512-8|LNC|Human papilloma virus Ab|Human papilloma virus Ab
C0367661|T201|COMP|5533-5|LNC|CD80|CD80
C0367662|T201|COMP|5532-7|LNC|CD8|CD8
C0367663|T201|COMP|5534-3|LNC|CD81|CD81
C0367664|T201|COMP|5535-0|LNC|CD82|CD82
C0367665|T201|COMP|5536-8|LNC|CD83|CD83
C0367666|T201|COMP|5537-6|LNC|CD85|CD85
C0367667|T201|COMP|5538-4|LNC|CD86|CD86
C0367668|T201|COMP|5539-2|LNC|CD87|CD87
C0367669|T201|COMP|5540-0|LNC|CD88|CD88
C0367670|T201|COMP|5541-8|LNC|CD89|CD89
C0367671|T201|COMP|5542-6|LNC|CD9|CD9
C0367672|T201|COMP|5543-4|LNC|CD91|CD91
C0367673|T201|COMP|5544-2|LNC|CD93|CD93
C0367674|T201|COMP|5545-9|LNC|CD94|CD94
C0367675|T201|COMP|5546-7|LNC|CD95|CD95
C0367676|T201|COMP|5547-5|LNC|CD96|CD96
C0367677|T201|COMP|5548-3|LNC|CD97|CD97
C0367678|T201|COMP|5549-1|LNC|CD98|CD98
C0367679|T201|COMP|5550-9|LNC|CD99|CD99
C0367680|T201|COMP|5551-7|LNC|CyCD3|CyCD3
C0367681|T201|COMP|5552-5|LNC|CyCD79|CyCD79
C0367682|T201|COMP|6513-6|LNC|Human papilloma virus Ab|Human papilloma virus Ab
C0367683|T201|COMP|5553-3|LNC|CyIg|CyIg
C0367684|T201|COMP|5554-1|LNC|CyIg mu|CyIg mu
C0367685|T201|COMP|5555-8|LNC|FMC7|FMC7
C0367686|T201|COMP|5556-6|LNC|GPA|GPA
C0367687|T201|COMP|5557-4|LNC|HLA-DR|HLA-DR
C0367688|T201|COMP|5558-2|LNC|Myeloperoxidase|Myeloperoxidase
C0367689|T201|COMP|5559-0|LNC|RFD9|RFD9
C0367690|T201|COMP|5560-8|LNC|SmIg|SmIg
C0367691|T201|COMP|5561-6|LNC|SmIg kappa|SmIg kappa
C0367692|T201|COMP|5562-4|LNC|SmIg lambda|SmIg lambda
C0367693|T201|COMP|5563-2|LNC|SmIg-CD79|SmIg-CD79
C0367694|T201|COMP|5564-0|LNC|TCR-CD3|TCR-CD3
C0367695|T201|COMP|5565-7|LNC|Terminal deoxyribonucleotidyl transferase|Terminal deoxyribonucleotidyl transferase
C0367696|T201|COMP|6514-4|LNC|Human papilloma virus rRNA|Human papilloma virus rRNA
C0367697|T201|COMP|6515-1|LNC|Human papilloma virus rRNA|Human papilloma virus rRNA
C0367699|T201|COMP|5567-3|LNC|Acetone|Acetone
C0367700|T201|COMP|5568-1|LNC|Acetone|Acetone
C0367701|T201|COMP|5569-9|LNC|Acetone|Acetone
C0367702|T201|COMP|5570-7|LNC|Acetone|Acetone
C0367703|T201|COMP|5571-5|LNC|Acrylonitrile|Acrylonitrile
C0367704|T201|COMP|5572-3|LNC|Aluminum|Aluminum
C0367705|T201|COMP|5573-1|LNC|Aluminum|Aluminum
C0367706|T201|COMP|5574-9|LNC|Aluminum|Aluminum
C0367707|T201|COMP|6516-9|LNC|Human papilloma virus rRNA|Human papilloma virus rRNA
C0367708|T201|COMP|5575-6|LNC|Aluminum|Aluminum
C0367709|T201|COMP|5576-4|LNC|Aluminum|Aluminum
C0367710|T201|COMP|5266-2|LNC|Paracoccidioides brasiliensis Ab|Paracoccidioides brasiliensis Ab
C0367711|T201|COMP|5577-2|LNC|Aluminum|Aluminum
C0367712|T201|COMP|5578-0|LNC|Antimony|Antimony
C0367713|T201|COMP|5579-8|LNC|Antimony|Antimony
C0367714|T201|COMP|5580-6|LNC|Antimony|Antimony
C0367715|T201|COMP|5581-4|LNC|Antimony|Antimony
C0367716|T201|COMP|5267-0|LNC|Paragonimus sp Ab|Paragonimus sp Ab
C0367717|T201|COMP|5268-8|LNC|Parainfluenza virus 1 Ab|Parainfluenza virus 1 Ab
C0367718|T201|COMP|5868-5|LNC|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C0367719|T201|COMP|5582-2|LNC|Arsenic|Arsenic
C0367720|T201|COMP|5583-0|LNC|Arsenic|Arsenic
C0367721|T201|COMP|5584-8|LNC|Arsenic|Arsenic
C0367722|T201|COMP|5869-3|LNC|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C0367723|T201|COMP|5585-5|LNC|Arsenic|Arsenic
C0367724|T201|COMP|5586-3|LNC|Arsenic|Arsenic
C0367725|T201|COMP|5587-1|LNC|Arsenic|Arsenic
C0367726|T201|COMP|5588-9|LNC|Barium|Barium
C0367727|T201|COMP|5589-7|LNC|Barium|Barium
C0367728|T201|COMP|5269-6|LNC|Parainfluenza virus 2 Ab|Parainfluenza virus 2 Ab
C0367729|T201|COMP|5590-5|LNC|Barium|Barium
C0367730|T201|COMP|5591-3|LNC|Benzene|Benzene
C0367731|T201|COMP|5870-1|LNC|Parainfluenza virus 2 Ag|Parainfluenza virus 2 Ag
C0367732|T201|COMP|5871-9|LNC|Parainfluenza virus 2 Ag|Parainfluenza virus 2 Ag
C0367733|T201|COMP|5270-4|LNC|Parainfluenza virus 3 Ab|Parainfluenza virus 3 Ab
C0367734|T201|COMP|5872-7|LNC|Parainfluenza virus 3 Ag|Parainfluenza virus 3 Ag
C0367735|T201|COMP|5873-5|LNC|Parainfluenza virus 3 Ag|Parainfluenza virus 3 Ag
C0367736|T201|COMP|5592-1|LNC|Benzene|Benzene
C0367737|T201|COMP|5593-9|LNC|Beryllium|Beryllium
C0367738|T201|COMP|5594-7|LNC|Beryllium|Beryllium
C0367739|T201|COMP|5595-4|LNC|Beryllium|Beryllium
C0367740|T201|COMP|6517-7|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0367741|T201|COMP|5596-2|LNC|Beryllium|Beryllium
C0367742|T201|COMP|5597-0|LNC|Bismuth|Bismuth
C0367743|T201|COMP|5598-8|LNC|Bismuth|Bismuth
C0367744|T201|COMP|5599-6|LNC|Boldenone|Boldenone
C0367745|T201|COMP|5600-2|LNC|Boldenone|Boldenone
C0367746|T201|COMP|5601-0|LNC|Boldenone|Boldenone
C0367747|T201|COMP|5602-8|LNC|Borate|Borate
C0367748|T201|COMP|5603-6|LNC|Borate|Borate
C0367749|T201|COMP|5604-4|LNC|Boron|Boron
C0367750|T201|COMP|5605-1|LNC|Boron|Boron
C0367751|T201|COMP|5606-9|LNC|Boron|Boron
C0367752|T201|COMP|5607-7|LNC|Boron|Boron
C0367753|T201|COMP|5608-5|LNC|Bufotenine|Bufotenine
C0367754|T201|COMP|5609-3|LNC|Cadmium|Cadmium
C0367755|T201|COMP|5610-1|LNC|Cadmium|Cadmium
C0367756|T201|COMP|5611-9|LNC|Cadmium|Cadmium
C0367757|T201|COMP|5612-7|LNC|Cadmium|Cadmium
C0367758|T201|COMP|5613-5|LNC|Carbon disulfide|Carbon disulfide
C0367759|T201|COMP|5614-3|LNC|Cesium|Cesium
C0367760|T201|COMP|5615-0|LNC|Cesium|Cesium
C0367761|T201|COMP|5616-8|LNC|Cesium|Cesium
C0367762|T201|COMP|5617-6|LNC|Cesium|Cesium
C0367763|T201|COMP|5618-4|LNC|Cesium|Cesium
C0367764|T201|COMP|5619-2|LNC|Chromium|Chromium
C0367765|T201|COMP|5620-0|LNC|Chromium|Chromium
C0367766|T201|COMP|5621-8|LNC|Chromium|Chromium
C0367767|T201|COMP|5622-6|LNC|Chromium|Chromium
C0367768|T201|COMP|5623-4|LNC|Chromium|Chromium
C0367769|T201|COMP|5624-2|LNC|Chromium|Chromium
C0367770|T201|COMP|5272-0|LNC|Parvovirus B19 Ab|Parvovirus B19 Ab
C0367771|T201|COMP|5625-9|LNC|Cobalt|Cobalt
C0367772|T201|COMP|5626-7|LNC|Cobalt|Cobalt
C0367773|T201|COMP|5627-5|LNC|Cobalt|Cobalt
C0367774|T201|COMP|5273-8|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0367775|T201|COMP|5274-6|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0367776|T201|COMP|5030-2|LNC|Parvovirus B19 RNA|Parvovirus B19 RNA
C0367777|T201|COMP|5031-0|LNC|Parvovirus B19 RNA|Parvovirus B19 RNA
C0367778|T201|COMP|5032-8|LNC|Parvovirus B19 RNA|Parvovirus B19 RNA
C0367779|T201|COMP|5628-3|LNC|Cobalt|Cobalt
C0367780|T201|COMP|5936-0|LNC|Benzoylecgonine|Benzoylecgonine
C0367781|T201|COMP|5938-6|LNC|Benzoylecgonine|Benzoylecgonine
C0367782|T201|COMP|3395-1|LNC|Cocaine|Cocaine
C0367783|T201|COMP|3396-9|LNC|Cocaine|Cocaine
C0367784|T201|COMP|3393-6|LNC|Benzoylecgonine|Benzoylecgonine
C0367786|T201|COMP|5629-1|LNC|Copper|Copper
C0367787|T201|COMP|5630-9|LNC|Copper|Copper
C0367788|T201|COMP|5631-7|LNC|Copper|Copper
C0367789|T201|COMP|5632-5|LNC|Copper|Copper
C0367790|T201|COMP|5633-3|LNC|Copper|Copper
C0367791|T201|COMP|5634-1|LNC|Cyanide|Cyanide
C0367792|T201|COMP|5635-8|LNC|Cyanide|Cyanide
C0367793|T201|COMP|5636-6|LNC|Cyanide|Cyanide
C0367794|T201|COMP|5637-4|LNC|Cyanide|Cyanide
C0367795|T201|COMP|5638-2|LNC|Diazinon|Diazinon
C0367797|T201|COMP|5640-8|LNC|Ethanol|Ethanol
C0367798|T201|COMP|5639-0|LNC|Ethanol|Ethanol
C0367799|T201|COMP|5642-4|LNC|Ethanol|Ethanol
C0367800|T201|COMP|5277-9|LNC|Penicillium roqueforti Ab|Penicillium roqueforti Ab
C0367801|T201|COMP|5643-2|LNC|Ethanol|Ethanol
C0367802|T201|COMP|5644-0|LNC|Ethanol|Ethanol
C0367803|T201|COMP|5645-7|LNC|Ethanol|Ethanol
C0367804|T201|COMP|5278-7|LNC|Plasmodium falciparum Ab|Plasmodium falciparum Ab
C0367805|T201|COMP|6305-7|LNC|Plasmodium malariae Ab|Plasmodium malariae Ab
C0367806|T201|COMP|6560-7|LNC|Plasmodium ovale Ab|Plasmodium ovale Ab
C0367807|T201|COMP|5279-5|LNC|Plasmodium sp Ab|Plasmodium sp Ab
C0367808|T201|COMP|5280-3|LNC|Plasmodium vivax Ab|Plasmodium vivax Ab
C0367809|T201|COMP|5646-5|LNC|Ethylene glycol|Ethylene glycol
C0367810|T201|COMP|5647-3|LNC|Ethylene glycol|Ethylene glycol
C0367811|T201|COMP|5648-1|LNC|Fluoride|Fluoride
C0367812|T201|COMP|5649-9|LNC|Fluoride|Fluoride
C0367813|T201|COMP|5650-7|LNC|Fluoride|Fluoride
C0367814|T201|COMP|5651-5|LNC|Fluoride|Fluoride
C0367815|T201|COMP|5652-3|LNC|Formaldehyde|Formaldehyde
C0367816|T201|COMP|5653-1|LNC|Formaldehyde|Formaldehyde
C0367817|T201|COMP|5654-9|LNC|Gallium|Gallium
C0367818|T201|COMP|5655-6|LNC|Germanium|Germanium
C0367819|T201|COMP|5656-4|LNC|Gold|Gold
C0367820|T201|COMP|5657-2|LNC|Gold|Gold
C0367821|T201|COMP|5658-0|LNC|Gold|Gold
C0367822|T201|COMP|5659-8|LNC|Gold|Gold
C0367823|T201|COMP|5660-6|LNC|Gold|Gold
C0367824|T201|COMP|5661-4|LNC|Gold|Gold
C0367825|T201|COMP|5662-2|LNC|Heavy metals|Heavy metals
C0367826|T201|COMP|6518-5|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0367827|T201|COMP|6519-3|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0367828|T201|COMP|700-5|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0367829|T201|COMP|6521-9|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C0367830|T201|COMP|5664-8|LNC|Heavy metals negative|Heavy metals negative
C0367831|T201|COMP|5281-1|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C0367832|T201|COMP|5282-9|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C0367833|T201|COMP|5283-7|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C0367834|T201|COMP|5284-5|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C0367835|T201|COMP|5285-2|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C0367836|T201|COMP|5286-0|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C0367837|T201|COMP|5287-8|LNC|Burkholderia pseudomallei Ab|Burkholderia pseudomallei Ab
C0367838|T201|COMP|6522-7|LNC|Rabies virus Ab|Rabies virus Ab
C0367839|T201|COMP|6523-5|LNC|Rabies virus Ab|Rabies virus Ab
C0367840|T201|COMP|5288-6|LNC|Rabies virus Ab|Rabies virus Ab
C0367841|T201|COMP|6524-3|LNC|Rabies virus Ab|Rabies virus Ab
C0367842|T201|COMP|6525-0|LNC|Rabies virus Ab|Rabies virus Ab
C0367843|T201|COMP|6526-8|LNC|Rabies virus Ab|Rabies virus Ab
C0367844|T201|COMP|6527-6|LNC|Rabies virus Ab|Rabies virus Ab
C0367845|T201|COMP|6529-2|LNC|Rabies virus Ag|Rabies virus Ag
C0367846|T201|COMP|6528-4|LNC|Rabies virus Ag|Rabies virus Ag
C0367847|T201|COMP|5663-0|LNC|Heavy metals positive|Heavy metals positive
C0367848|T201|COMP|5665-5|LNC|Indium|Indium
C0367849|T201|COMP|5666-3|LNC|Indium|Indium
C0367850|T201|COMP|5667-1|LNC|Isopropanol|Isopropanol
C0367851|T201|COMP|6533-4|LNC|Rabies virus Ag|Rabies virus Ag
C0367852|T201|COMP|6532-6|LNC|Rabies virus Ag|Rabies virus Ag
C0367853|T201|COMP|6536-7|LNC|Rabies virus identified|Rabies virus identified
C0367854|T201|COMP|5668-9|LNC|Isopropanol|Isopropanol
C0367855|T201|COMP|5669-7|LNC|Isopropanol|Isopropanol
C0367856|T201|COMP|5670-5|LNC|Isopropanol|Isopropanol
C0367857|T201|COMP|5671-3|LNC|Lead|Lead
C0367858|T201|COMP|5672-1|LNC|Lead|Lead
C0367859|T201|COMP|5673-9|LNC|Lead|Lead
C0367860|T201|COMP|5674-7|LNC|Lead|Lead
C0367861|T201|COMP|5675-4|LNC|Lead|Lead
C0367862|T201|COMP|5676-2|LNC|Lead|Lead
C0367863|T201|COMP|5677-0|LNC|Lead|Lead
C0367864|T201|COMP|5678-8|LNC|Lysergate diethylamide|Lysergate diethylamide
C0367865|T201|COMP|6539-1|LNC|Rabies virus identified|Rabies virus identified
C0367866|T201|COMP|5680-4|LNC|Malathion|Malathion
C0367867|T201|COMP|5681-2|LNC|Manganese|Manganese
C0367868|T201|COMP|5682-0|LNC|Manganese|Manganese
C0367869|T201|COMP|5683-8|LNC|Manganese|Manganese
C0367870|T201|COMP|5684-6|LNC|Manganese|Manganese
C0367871|T201|COMP|5685-3|LNC|Mercury|Mercury
C0367872|T201|COMP|5686-1|LNC|Mercury|Mercury
C0367873|T201|COMP|5687-9|LNC|Mercury|Mercury
C0367874|T201|COMP|5688-7|LNC|Mercury|Mercury
C0367875|T201|COMP|5689-5|LNC|Mercury|Mercury
C0367877|T201|COMP|5289-4|LNC|Reagin Ab|Reagin Ab
C0367879|T201|COMP|5290-2|LNC|Reagin Ab|Reagin Ab
C0367881|T201|COMP|5692-9|LNC|Methanol|Methanol
C0367882|T201|COMP|5695-2|LNC|Methanol|Methanol
C0367883|T201|COMP|5694-5|LNC|Methanol|Methanol
C0367884|T201|COMP|5697-8|LNC|Molybdenum|Molybdenum
C0367885|T201|COMP|5696-0|LNC|Molybdenum|Molybdenum
C0367886|T201|COMP|5698-6|LNC|Molybdenum|Molybdenum
C0367887|T201|COMP|5291-0|LNC|Reagin Ab|Reagin Ab
C0367888|T201|COMP|5292-8|LNC|Reagin Ab|Reagin Ab
C0367889|T201|COMP|5699-4|LNC|Molybdenum|Molybdenum
C0367890|T201|COMP|5293-6|LNC|Reovirus Ab|Reovirus Ab
C0367891|T201|COMP|5294-4|LNC|Respiratory syncytial virus Ab|Respiratory syncytial virus Ab
C0367892|T201|COMP|5295-1|LNC|Respiratory syncytial virus Ab|Respiratory syncytial virus Ab
C0367893|T201|COMP|5874-3|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C0367894|T201|COMP|5876-8|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C0367895|T201|COMP|5877-6|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C0367896|T201|COMP|5303-3|LNC|Rickettsia (Proteus OX19) Ab|Rickettsia (Proteus OX19) Ab
C0367897|T201|COMP|5875-0|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C0367898|T201|COMP|5305-8|LNC|Rickettsia (Proteus OXK) Ab|Rickettsia (Proteus OXK) Ab
C0367899|T201|COMP|5306-6|LNC|Rickettsia sp Ab|Rickettsia sp Ab
C0367900|T201|COMP|6542-5|LNC|Rickettsia prowazekii Ab|Rickettsia prowazekii Ab
C0367901|T201|COMP|5304-1|LNC|Rickettsia (Proteus OX2) Ab|Rickettsia (Proteus OX2) Ab
C0367908|T201|COMP|5700-0|LNC|Nickel|Nickel
C0367909|T201|COMP|5701-8|LNC|Nickel|Nickel
C0367911|T201|COMP|5703-4|LNC|Nickel|Nickel
C0367912|T201|COMP|5704-2|LNC|Nickel|Nickel
C0367913|T201|COMP|5705-9|LNC|Nickel|Nickel
C0367914|T201|COMP|5706-7|LNC|Opiates|Opiates
C0367915|T201|COMP|5708-3|LNC|Paraquat|Paraquat
C0367916|T201|COMP|5709-1|LNC|Paraquat|Paraquat
C0367917|T201|COMP|5710-9|LNC|Pentachlorophenol|Pentachlorophenol
C0367918|T201|COMP|5711-7|LNC|Pentachlorophenol|Pentachlorophenol
C0367919|T201|COMP|5713-3|LNC|Platinum|Platinum
C0367920|T201|COMP|5714-1|LNC|Platinum|Platinum
C0367922|T201|COMP|5715-8|LNC|Platinum|Platinum
C0367923|T201|COMP|5717-4|LNC|Polychlorinated biphenyl|Polychlorinated biphenyl
C0367924|T201|COMP|5716-6|LNC|Polychlorinated biphenyl|Polychlorinated biphenyl
C0367925|T201|COMP|5718-2|LNC|Rubidium|Rubidium
C0367926|T201|COMP|5719-0|LNC|Rubidium|Rubidium
C0367927|T201|COMP|5720-8|LNC|Rubidium|Rubidium
C0367928|T201|COMP|5721-6|LNC|Rubidium|Rubidium
C0367929|T201|COMP|5722-4|LNC|Selenium|Selenium
C0367930|T201|COMP|5724-0|LNC|Selenium|Selenium
C0367931|T201|COMP|5723-2|LNC|Selenium|Selenium
C0367932|T201|COMP|5725-7|LNC|Selenium|Selenium
C0367933|T201|COMP|5726-5|LNC|Selenium|Selenium
C0367934|T201|COMP|5727-3|LNC|Selenium|Selenium
C0367935|T201|COMP|5729-9|LNC|Silicate|Silicate
C0367936|T201|COMP|5730-7|LNC|Silicate|Silicate
C0367937|T201|COMP|5731-5|LNC|Silicate|Silicate
C0367939|T201|COMP|5728-1|LNC|Silicon|Silicon
C0367943|T201|COMP|5732-3|LNC|Silver|Silver
C0367944|T201|COMP|5733-1|LNC|Silver|Silver
C0367945|T201|COMP|5734-9|LNC|Silver|Silver
C0367946|T201|COMP|5735-6|LNC|Silver|Silver
C0367947|T201|COMP|5736-4|LNC|Strontium|Strontium
C0367948|T201|COMP|5737-2|LNC|Strychnine|Strychnine
C0367949|T201|COMP|5738-0|LNC|Strychnine|Strychnine
C0367950|T201|COMP|5739-8|LNC|Strychnine|Strychnine
C0367951|T201|COMP|5740-6|LNC|Strychnine|Strychnine
C0367953|T201|COMP|5741-4|LNC|Strychnine|Strychnine
C0367954|T201|COMP|5742-2|LNC|Tellurium|Tellurium
C0367955|T201|COMP|5743-0|LNC|Thallium|Thallium
C0367956|T201|COMP|5744-8|LNC|Thallium|Thallium
C0367957|T201|COMP|5745-5|LNC|Thallium|Thallium
C0367958|T201|COMP|5746-3|LNC|Thallium|Thallium
C0367960|T201|COMP|5747-1|LNC|Tin|Tin
C0367961|T201|COMP|5748-9|LNC|Tin|Tin
C0367963|T201|COMP|5749-7|LNC|Titanium|Titanium
C0367964|T201|COMP|5750-5|LNC|Toluene|Toluene
C0367965|T201|COMP|5751-3|LNC|Uranium|Uranium
C0367966|T201|COMP|5752-1|LNC|Uranium|Uranium
C0367967|T201|COMP|5753-9|LNC|Vanadium|Vanadium
C0367968|T201|COMP|5754-7|LNC|Vanadium|Vanadium
C0367969|T201|COMP|5755-4|LNC|Vanadium|Vanadium
C0367970|T201|COMP|5756-2|LNC|Vanadium|Vanadium
C0367971|T201|COMP|5757-0|LNC|Vanadium|Vanadium
C0367972|T201|COMP|5758-8|LNC|Dimethylbenzene|Dimethylbenzene
C0367973|T201|COMP|5759-6|LNC|Dimethylbenzene|Dimethylbenzene
C0367974|T201|COMP|5760-4|LNC|Zinc|Zinc
C0367975|T201|COMP|5761-2|LNC|Zinc|Zinc
C0367976|T201|COMP|5307-4|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C0367977|T201|COMP|5762-0|LNC|Zinc|Zinc
C0367978|T201|COMP|5763-8|LNC|Zinc|Zinc
C0367979|T201|COMP|5764-6|LNC|Zinc|Zinc
C0367980|T201|COMP|5765-3|LNC|Zinc|Zinc
C0367981|T201|COMP|5766-1|LNC|Ammonium urate crystals|Ammonium urate crystals
C0367982|T201|COMP|5767-9|LNC|Appearance|Appearance
C0367983|T201|COMP|5768-7|LNC|Ascorbate|Ascorbate
C0367984|T201|COMP|5769-5|LNC|Bacteria|Bacteria
C0367985|T201|COMP|5770-3|LNC|Bilirubin|Bilirubin
C0367986|T201|COMP|5771-1|LNC|Bilirubin crystals|Bilirubin crystals
C0367987|T201|COMP|5308-2|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C0367988|T201|COMP|5772-9|LNC|Calcium carbonate crystals|Calcium carbonate crystals
C0367989|T201|COMP|6543-3|LNC|Rickettsia rickettsii Ag|Rickettsia rickettsii Ag
C0367990|T201|COMP|5773-7|LNC|Calcium carbonate crystals|Calcium carbonate crystals
C0367991|T201|COMP|5878-4|LNC|Rickettsia sp identified|Rickettsia sp identified
C0367992|T201|COMP|6544-1|LNC|Rickettsia sp identified|Rickettsia sp identified
C0367993|T201|COMP|6545-8|LNC|Rickettsia sp identified|Rickettsia sp identified
C0367994|T201|COMP|5774-5|LNC|Calcium oxalate crystals|Calcium oxalate crystals
C0367995|T201|COMP|6546-6|LNC|Rickettsia sp identified|Rickettsia sp identified
C0367996|T201|COMP|5323-1|LNC|Orientia tsutsugamushi Ab|Orientia tsutsugamushi Ab
C0367997|T201|COMP|5324-9|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C0367998|T201|COMP|5325-6|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C0367999|T201|COMP|5775-2|LNC|Calcium phosphate crystals|Calcium phosphate crystals
C0368000|T201|COMP|5776-0|LNC|Calcium sulfate crystals|Calcium sulfate crystals
C0368001|T201|COMP|5777-8|LNC|Cholesterol crystals|Cholesterol crystals
C0368002|T201|COMP|5778-6|LNC|Color|Color
C0368003|T201|COMP|5779-4|LNC|Crystals|Crystals
C0368004|T201|COMP|5780-2|LNC|Crystals|Crystals
C0368005|T201|COMP|5781-0|LNC|Crystals|Crystals
C0368006|T201|COMP|5782-8|LNC|Crystals|Crystals
C0368007|T201|COMP|5783-6|LNC|Crystals.unidentified|Crystals.unidentified
C0368008|T201|COMP|5784-4|LNC|Cystine crystals|Cystine crystals
C0368009|T201|COMP|5785-1|LNC|Eosinophils|Eosinophils
C0368010|T201|COMP|5786-9|LNC|Epithelial casts|Epithelial casts
C0368011|T201|COMP|5787-7|LNC|Epithelial cells|Epithelial cells
C0368012|T201|COMP|5807-3|LNC|Erythrocyte casts|Erythrocyte casts
C0368013|T201|COMP|5808-1|LNC|Erythrocytes|Erythrocytes
C0368014|T201|COMP|5788-5|LNC|Oval fat bodies (globules)|Oval fat bodies (globules)
C0368015|T201|COMP|5789-3|LNC|Fatty casts|Fatty casts
C0368016|T201|COMP|5790-1|LNC|Fungi.filamentous|Fungi.filamentous
C0368017|T201|COMP|5791-9|LNC|Fungi.yeastlike|Fungi.yeastlike
C0368018|T201|COMP|5792-7|LNC|Glucose|Glucose
C0368020|T201|COMP|5794-3|LNC|Hemoglobin|Hemoglobin
C0368021|T201|COMP|5793-5|LNC|Granular casts|Granular casts
C0368022|T201|COMP|5795-0|LNC|Hippurate crystals|Hippurate crystals
C0368024|T201|COMP|5328-0|LNC|Rotavirus Ab|Rotavirus Ab
C0368025|T201|COMP|5796-8|LNC|Hyaline casts|Hyaline casts
C0368026|T201|COMP|5329-8|LNC|Rotavirus Ab|Rotavirus Ab
C0368027|T201|COMP|5879-2|LNC|Rotavirus Ag|Rotavirus Ag
C0368028|T201|COMP|5880-0|LNC|Rotavirus Ag|Rotavirus Ag
C0368029|T201|COMP|6547-4|LNC|Rotavirus identified|Rotavirus identified
C0368030|T201|COMP|5330-6|LNC|Rubella virus Ab|Rubella virus Ab
C0368031|T201|COMP|5331-4|LNC|Rubella virus Ab|Rubella virus Ab
C0368032|T201|COMP|5797-6|LNC|Ketones|Ketones
C0368033|T201|COMP|5798-4|LNC|Leucine crystals|Leucine crystals
C0368034|T201|COMP|5820-6|LNC|Leukocyte casts|Leukocyte casts
C0368035|T201|COMP|5799-2|LNC|Leukocyte esterase|Leukocyte esterase
C0368036|T201|COMP|5821-4|LNC|Leukocytes|Leukocytes
C0368037|T201|COMP|5800-8|LNC|Lipids|Lipids
C0368038|T201|COMP|5801-6|LNC|Magnesium ammonium phosphate crystals|Magnesium ammonium phosphate crystals
C0368039|T201|COMP|5332-2|LNC|Rubella virus Ab|Rubella virus Ab
C0368040|T201|COMP|5802-4|LNC|Nitrite|Nitrite
C0368041|T201|COMP|5333-0|LNC|Rubella virus Ab|Rubella virus Ab
C0368043|T201|COMP|5804-0|LNC|Protein|Protein
C0368044|T201|COMP|5334-8|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0368045|T201|COMP|5335-5|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C0368046|T201|COMP|6548-2|LNC|Rubella virus identified|Rubella virus identified
C0368048|T201|COMP|5365-2|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0368049|T201|COMP|6549-0|LNC|Saint Louis encephalitis virus Ag|Saint Louis encephalitis virus Ag
C0368050|T201|COMP|5338-9|LNC|Salmonella sp Ab|Salmonella sp Ab
C0368051|T201|COMP|5805-7|LNC|Pyrophosphate crystals|Pyrophosphate crystals
C0368052|T201|COMP|5339-7|LNC|Salmonella paratyphi A H Ab|Salmonella paratyphi A H Ab
C0368053|T201|COMP|5340-5|LNC|Salmonella paratyphi A O Ab|Salmonella paratyphi A O Ab
C0368054|T201|COMP|5341-3|LNC|Salmonella paratyphi B H Ab|Salmonella paratyphi B H Ab
C0368055|T201|COMP|5342-1|LNC|Salmonella paratyphi B O Ab|Salmonella paratyphi B O Ab
C0368056|T201|COMP|5343-9|LNC|Salmonella paratyphi C H Ab|Salmonella paratyphi C H Ab
C0368057|T201|COMP|5806-5|LNC|Pyrophosphate crystals|Pyrophosphate crystals
C0368058|T201|COMP|5809-9|LNC|Reducing substances|Reducing substances
C0368059|T201|COMP|5810-7|LNC|Specific gravity|Specific gravity
C0368060|T201|COMP|5344-7|LNC|Salmonella paratyphi C O Ab|Salmonella paratyphi C O Ab
C0368061|T201|COMP|5811-5|LNC|Specific gravity|Specific gravity
C0368062|T201|COMP|5812-3|LNC|Sulfonamide crystals|Sulfonamide crystals
C0368063|T201|COMP|5813-1|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C0368064|T201|COMP|5345-4|LNC|Salmonella typhi H Ab|Salmonella typhi H Ab
C0368065|T201|COMP|5814-9|LNC|Triple phosphate crystals|Triple phosphate crystals
C0368066|T201|COMP|5346-2|LNC|Salmonella typhi O Ab|Salmonella typhi O Ab
C0368067|T201|COMP|5347-0|LNC|Schistosoma sp Ab|Schistosoma sp Ab
C0368068|T201|COMP|5363-7|LNC|Spirillum minus Ab|Spirillum minus Ab
C0368069|T201|COMP|5033-6|LNC|Staphylococcus aureus rRNA|Staphylococcus aureus rRNA
C0368070|T201|COMP|5350-4|LNC|Shigella sp Ab|Shigella sp Ab
C0368071|T201|COMP|5364-5|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C0368072|T201|COMP|6550-8|LNC|Staphylococcus aureus Ab|Staphylococcus aureus Ab
C0368073|T201|COMP|5366-0|LNC|Staphylolysin Ab|Staphylolysin Ab
C0368074|T201|COMP|5367-8|LNC|Streptobacillus moniliformis Ab|Streptobacillus moniliformis Ab
C0368075|T201|COMP|5815-6|LNC|Tyrosine crystals|Tyrosine crystals
C0368076|T201|COMP|5816-4|LNC|Urate crystals|Urate crystals
C0368077|T201|COMP|5817-2|LNC|Urate crystals|Urate crystals
C0368078|T201|COMP|5818-0|LNC|Urobilinogen|Urobilinogen
C0368079|T201|COMP|5819-8|LNC|Waxy casts|Waxy casts
C0368080|T201|COMP|5822-2|LNC|Yeast|Yeast
C0368082|T201|COMP|6306-5|LNC|Adenovirus 40+41 Ag|Adenovirus 40+41 Ag
C0368083|T201|COMP|5041-9|LNC|Adenovirus Ab|Adenovirus Ab
C0368084|T201|COMP|5042-7|LNC|Adenovirus Ab.IgM|Adenovirus Ab.IgM
C0368085|T201|COMP|5823-0|LNC|Adenovirus Ag|Adenovirus Ag
C0368086|T201|COMP|5824-8|LNC|Adenovirus Ag|Adenovirus Ag
C0368087|T201|COMP|5825-5|LNC|Adenovirus Ag|Adenovirus Ag
C0368088|T201|COMP|5826-3|LNC|Adenovirus Ag|Adenovirus Ag
C0368089|T201|COMP|5827-1|LNC|Adenovirus Ag|Adenovirus Ag
C0368090|T201|COMP|5828-9|LNC|Adenovirus Ag|Adenovirus Ag
C0368091|T201|COMP|5829-7|LNC|Adenovirus Ag|Adenovirus Ag
C0368092|T201|COMP|5830-5|LNC|Adenovirus Ag|Adenovirus Ag
C0368093|T201|COMP|5831-3|LNC|Adenovirus Ag|Adenovirus Ag
C0368094|T201|COMP|5832-1|LNC|Adenovirus Ag|Adenovirus Ag
C0368095|T201|COMP|5833-9|LNC|Adenovirus Ag|Adenovirus Ag
C0368096|T201|COMP|5834-7|LNC|Adenovirus Ag|Adenovirus Ag
C0368097|T201|COMP|6307-3|LNC|Adenovirus rRNA|Adenovirus rRNA
C0368098|T201|COMP|6308-1|LNC|Adenovirus rRNA|Adenovirus rRNA
C0368099|T201|COMP|5045-0|LNC|Ancylostoma sp Ab|Ancylostoma sp Ab
C0368100|T201|COMP|6309-9|LNC|Arbovirus identified|Arbovirus identified
C0368101|T201|COMP|6310-7|LNC|Arbovirus identified|Arbovirus identified
C0368102|T201|COMP|5049-2|LNC|Ascaris lumbricoides Ab|Ascaris lumbricoides Ab
C0368103|T201|COMP|5050-0|LNC|Aspergillus fumigatus Ab|Aspergillus fumigatus Ab
C0368104|T201|COMP|5051-8|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C0368105|T201|COMP|5052-6|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C0368106|T201|COMP|5053-4|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C0368107|T201|COMP|6311-5|LNC|Babesia microti Ab|Babesia microti Ab
C0368108|T201|COMP|5054-2|LNC|Babesia sp Ab|Babesia sp Ab
C0368109|T201|COMP|5055-9|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0368110|T201|COMP|544-7|LNC|Bacteroides fragilis Ag|Bacteroides fragilis Ag
C0368111|T201|COMP|545-4|LNC|Bacteroides melaninogenicus Ag|Bacteroides melaninogenicus Ag
C0368112|T201|COMP|6312-3|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C0368113|T201|COMP|5057-5|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0368116|T201|COMP|4990-8|LNC|Blastomyces dermatitidis rRNA|Blastomyces dermatitidis rRNA
C0368117|T201|COMP|548-8|LNC|Bordetella pertussis|Bordetella pertussis
C0368118|T201|COMP|549-6|LNC|Bordetella pertussis|Bordetella pertussis
C0368121|T201|COMP|6315-6|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C0368122|T201|COMP|6316-4|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C0368123|T201|COMP|550-4|LNC|Bordetella pertussis Ag|Bordetella pertussis Ag
C0368124|T201|COMP|6317-2|LNC|Bordetella sp identified|Bordetella sp identified
C0368125|T201|COMP|6318-0|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0368126|T201|COMP|6319-8|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0368127|T201|COMP|5060-9|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0368128|T201|COMP|5061-7|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0368129|T201|COMP|5062-5|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0368130|T201|COMP|6320-6|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0368131|T201|COMP|5063-3|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0368132|T201|COMP|5064-1|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0368133|T201|COMP|6321-4|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0368134|T201|COMP|5065-8|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0368135|T201|COMP|6322-2|LNC|Borrelia burgdorferi Ag|Borrelia burgdorferi Ag
C0368136|T201|COMP|4991-6|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C0368137|T201|COMP|6323-0|LNC|Borrelia sp identified|Borrelia sp identified
C0368138|T201|COMP|5066-6|LNC|Brucella abortus Ab|Brucella abortus Ab
C0368139|T201|COMP|6324-8|LNC|Brucella abortus Ab|Brucella abortus Ab
C0368140|T201|COMP|6325-5|LNC|Brucella abortus Ab|Brucella abortus Ab
C0368141|T201|COMP|5067-4|LNC|Brucella abortus Ab|Brucella abortus Ab
C0368142|T201|COMP|6326-3|LNC|Brucella abortus Ab.IgM|Brucella abortus Ab.IgM
C0368143|T201|COMP|6327-1|LNC|Brucella canis Ab|Brucella canis Ab
C0368144|T201|COMP|5068-2|LNC|Brucella canis Ab|Brucella canis Ab
C0368145|T201|COMP|5069-0|LNC|Brucella melitensis Ab|Brucella melitensis Ab
C0368146|T201|COMP|551-2|LNC|Brucella sp identified|Brucella sp identified
C0368147|T201|COMP|552-0|LNC|Brucella sp identified|Brucella sp identified
C0368148|T201|COMP|6328-9|LNC|Brucella sp Ab|Brucella sp Ab
C0368149|T201|COMP|5070-8|LNC|Brucella sp Ab.IgM|Brucella sp Ab.IgM
C0368150|T201|COMP|5071-6|LNC|Brucella suis Ab|Brucella suis Ab
C0368151|T201|COMP|5072-4|LNC|Brush border Ab|Brush border Ab
C0368153|T201|COMP|6329-7|LNC|Campylobacter coli rRNA|Campylobacter coli rRNA
C0368154|T201|COMP|6330-5|LNC|Campylobacter sp identified|Campylobacter sp identified
C0368155|T201|COMP|6331-3|LNC|Campylobacter sp identified|Campylobacter sp identified
C0368157|T201|COMP|6333-9|LNC|Campylobacter jejuni rRNA|Campylobacter jejuni rRNA
C0368158|T201|COMP|6334-7|LNC|Campylobacter lari rRNA|Campylobacter lari rRNA
C0368159|T201|COMP|6332-1|LNC|Campylobacter sp identified|Campylobacter sp identified
C0368160|T201|COMP|4992-4|LNC|Campylobacter sp rRNA|Campylobacter sp rRNA
C0368161|T201|COMP|16537-3|LNC|Candida albicans Ab|Candida albicans Ab
C0368163|T201|COMP|6337-0|LNC|Candida albicans Ag|Candida albicans Ag
C0368164|T201|COMP|5075-7|LNC|Candida albicans Ag|Candida albicans Ag
C0368165|T201|COMP|553-8|LNC|Candida sp identified|Candida sp identified
C0368166|T201|COMP|554-6|LNC|Candida sp identified|Candida sp identified
C0368167|T201|COMP|555-3|LNC|Candida sp identified|Candida sp identified
C0368168|T201|COMP|5078-1|LNC|Chlamydophila pneumoniae Ab|Chlamydophila pneumoniae Ab
C0368169|T201|COMP|5079-9|LNC|Chlamydophila psittaci Ab|Chlamydophila psittaci Ab
C0368170|T201|COMP|5080-7|LNC|Chlamydophila psittaci Ab.IgG|Chlamydophila psittaci Ab.IgG
C0368171|T201|COMP|5081-5|LNC|Chlamydophila psittaci Ab.IgM|Chlamydophila psittaci Ab.IgM
C0368172|T201|COMP|6338-8|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C0368173|T201|COMP|6339-6|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C0368174|T201|COMP|6340-4|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C0368175|T201|COMP|6341-2|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C0368176|T201|COMP|556-1|LNC|Chlamydia sp identified|Chlamydia sp identified
C0368177|T201|COMP|557-9|LNC|Chlamydia sp identified|Chlamydia sp identified
C0368178|T201|COMP|558-7|LNC|Chlamydia sp identified|Chlamydia sp identified
C0368179|T201|COMP|559-5|LNC|Chlamydia sp identified|Chlamydia sp identified
C0368180|T201|COMP|560-3|LNC|Chlamydia sp identified|Chlamydia sp identified
C0368181|T201|COMP|5082-3|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0368182|T201|COMP|5083-1|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0368183|T201|COMP|5084-9|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0368184|T201|COMP|5085-6|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C0368185|T201|COMP|5086-4|LNC|Chlamydia sp Ab.IgM|Chlamydia sp Ab.IgM
C0368186|T201|COMP|6343-8|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0368187|T201|COMP|6344-6|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0368188|T201|COMP|6345-3|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0368189|T201|COMP|6346-1|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0368190|T201|COMP|6347-9|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0368191|T201|COMP|561-1|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0368192|T201|COMP|6348-7|LNC|Chlamydia sp identified|Chlamydia sp identified
C0368193|T201|COMP|6349-5|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C0368194|T201|COMP|5087-2|LNC|Chlamydia trachomatis Ab|Chlamydia trachomatis Ab
C0368195|T201|COMP|5088-0|LNC|Chlamydia trachomatis Ab|Chlamydia trachomatis Ab
C0368196|T201|COMP|5089-8|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C0368197|T201|COMP|5090-6|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C0368198|T201|COMP|6350-3|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0368199|T201|COMP|6351-1|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0368200|T201|COMP|6352-9|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0368201|T201|COMP|6353-7|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0368202|T201|COMP|6354-5|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0368203|T201|COMP|6355-2|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0368204|T201|COMP|6356-0|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0368205|T201|COMP|6357-8|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0368206|T201|COMP|4993-2|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C0368207|T201|COMP|562-9|LNC|Clostridioides difficile|Clostridioides difficile
C0368208|T201|COMP|563-7|LNC|Clostridioides difficile|Clostridioides difficile
C0368209|T201|COMP|6359-4|LNC|Clostridioides difficile toxin A|Clostridioides difficile toxin A
C0368210|T201|COMP|6360-2|LNC|Clostridioides difficile toxin A|Clostridioides difficile toxin A
C0368211|T201|COMP|6361-0|LNC|Clostridioides difficile toxin A+B|Clostridioides difficile toxin A+B
C0368212|T201|COMP|6363-6|LNC|Clostridioides difficile toxin A+B|Clostridioides difficile toxin A+B
C0368213|T201|COMP|6362-8|LNC|Clostridioides difficile toxin A+B|Clostridioides difficile toxin A+B
C0368214|T201|COMP|6364-4|LNC|Clostridioides difficile toxin A+B|Clostridioides difficile toxin A+B
C0368215|T201|COMP|6365-1|LNC|Clostridioides difficile toxin B|Clostridioides difficile toxin B
C0368216|T201|COMP|6366-9|LNC|Clostridioides difficile toxin B|Clostridioides difficile toxin B
C0368217|T201|COMP|5092-2|LNC|Clostridium tetani Ab|Clostridium tetani Ab
C0368218|T201|COMP|5093-0|LNC|Clostridium tetani Ab|Clostridium tetani Ab
C0368219|T201|COMP|6367-7|LNC|Clostridium tetani Ab.IgG|Clostridium tetani Ab.IgG
C0368220|T201|COMP|5094-8|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0368221|T201|COMP|5095-5|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0368222|T201|COMP|5096-3|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0368223|T201|COMP|6368-5|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0368224|T201|COMP|4994-0|LNC|Coccidioides immitis rRNA|Coccidioides immitis rRNA
C0368225|T201|COMP|564-5|LNC|Colony count|Colony count
C0368226|T201|COMP|565-2|LNC|Colony count|Colony count
C0368227|T201|COMP|5099-7|LNC|Coronavirus Ab|Coronavirus Ab
C0368229|T201|COMP|5101-1|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C0368230|T201|COMP|5102-9|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C0368231|T201|COMP|5103-7|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C0368232|T201|COMP|5104-5|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C0368233|T201|COMP|5105-2|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C0368234|T201|COMP|5106-0|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C0368235|T201|COMP|5107-8|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C0368236|T201|COMP|5108-6|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C0368237|T201|COMP|5109-4|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C0368238|T201|COMP|5110-2|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C0368239|T201|COMP|5111-0|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C0368240|T201|COMP|5112-8|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C0368241|T201|COMP|5113-6|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C0368242|T201|COMP|5114-4|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C0368245|T201|COMP|6369-3|LNC|Cryptococcus neoformans Ab|Cryptococcus neoformans Ab
C0368246|T201|COMP|5118-5|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C0368247|T201|COMP|5119-3|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C0368248|T201|COMP|4995-7|LNC|Cryptococcus neoformans rRNA|Cryptococcus neoformans rRNA
C0368249|T201|COMP|6370-1|LNC|Cryptococcus sp Ab|Cryptococcus sp Ab
C0368250|T201|COMP|6371-9|LNC|Cryptosporidium sp Ag|Cryptosporidium sp Ag
C0368251|T201|COMP|6372-7|LNC|Cryptosporidium sp Ag|Cryptosporidium sp Ag
C0368253|T201|COMP|6373-5|LNC|Taenia solium larva Ab.IgG|Taenia solium larva Ab.IgG
C0368254|T201|COMP|6374-3|LNC|Taenia solium larva Ab.IgG|Taenia solium larva Ab.IgG
C0368255|T201|COMP|5120-1|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C0368257|T201|COMP|5122-7|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0368258|T201|COMP|5121-9|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0368259|T201|COMP|5124-3|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0368260|T201|COMP|5125-0|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0368261|T201|COMP|5126-8|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0368262|T201|COMP|5127-6|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0368263|T201|COMP|6375-0|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0368264|T201|COMP|6376-8|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0368265|T201|COMP|6377-6|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0368266|T201|COMP|6378-4|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0368267|T201|COMP|6380-0|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0368268|T201|COMP|6379-2|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0368269|T201|COMP|6381-8|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0368270|T201|COMP|4996-5|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C0368271|T201|COMP|4997-3|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C0368272|T201|COMP|4998-1|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C0368273|T201|COMP|4999-9|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C0368274|T201|COMP|5000-5|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C0368275|T201|COMP|5835-4|LNC|Cytomegalovirus|Cytomegalovirus
C0368276|T201|COMP|5836-2|LNC|Cytomegalovirus|Cytomegalovirus
C0368277|T201|COMP|5837-0|LNC|Cytomegalovirus|Cytomegalovirus
C0368278|T201|COMP|5838-8|LNC|Cytomegalovirus|Cytomegalovirus
C0368281|T201|COMP|6384-2|LNC|Dengue virus Ag|Dengue virus Ag
C0368282|T201|COMP|6385-9|LNC|Dengue virus Ag|Dengue virus Ag
C0368283|T201|COMP|6386-7|LNC|Dengue virus DNA|Dengue virus DNA
C0368284|T201|COMP|6387-5|LNC|Dengue virus DNA|Dengue virus DNA
C0368285|T201|COMP|567-8|LNC|Diphtheria sp identified|Diphtheria sp identified
C0368286|T201|COMP|5133-4|LNC|DNAse B Ab.Streptococcal|DNAse B Ab.Streptococcal
C0368287|T201|COMP|5134-2|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0368288|T201|COMP|6388-3|LNC|Eastern equine encephalitis virus Ag|Eastern equine encephalitis virus Ag
C0368289|T201|COMP|6389-1|LNC|Eastern equine encephalitis virus Ag|Eastern equine encephalitis virus Ag
C0368290|T201|COMP|6390-9|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0368291|T201|COMP|6391-7|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0368292|T201|COMP|5135-9|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0368293|T201|COMP|5136-7|LNC|Echovirus 1 Ab|Echovirus 1 Ab
C0368294|T201|COMP|5137-5|LNC|Echovirus 1 Ab|Echovirus 1 Ab
C0368295|T201|COMP|5138-3|LNC|Echovirus 19 Ab|Echovirus 19 Ab
C0368296|T201|COMP|5139-1|LNC|Echovirus 19 Ab|Echovirus 19 Ab
C0368297|T201|COMP|5140-9|LNC|Echovirus 3 Ab|Echovirus 3 Ab
C0368298|T201|COMP|5141-7|LNC|Echovirus 3 Ab|Echovirus 3 Ab
C0368299|T201|COMP|6393-3|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C0368300|T201|COMP|6392-5|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C0368301|T201|COMP|5142-5|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C0368302|T201|COMP|5143-3|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C0368303|T201|COMP|6395-8|LNC|Echovirus 40 Ab|Echovirus 40 Ab
C0368304|T201|COMP|6394-1|LNC|Echovirus 40 Ab|Echovirus 40 Ab
C0368305|T201|COMP|5144-1|LNC|Echovirus 6 Ab|Echovirus 6 Ab
C0368306|T201|COMP|5145-8|LNC|Echovirus 6 Ab|Echovirus 6 Ab
C0368307|T201|COMP|5146-6|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C0368308|T201|COMP|5147-4|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C0368309|T201|COMP|5148-2|LNC|Echovirus NOS Ab|Echovirus NOS Ab
C0368310|T201|COMP|5149-0|LNC|Echovirus NOS Ab|Echovirus NOS Ab
C0368311|T201|COMP|6396-6|LNC|Entamoeba histolytica DNA|Entamoeba histolytica DNA
C0368312|T201|COMP|5150-8|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0368313|T201|COMP|5151-6|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0368314|T201|COMP|6397-4|LNC|Entamoeba histolytica Ag|Entamoeba histolytica Ag
C0368315|T201|COMP|6398-2|LNC|Entamoeba histolytica Ag|Entamoeba histolytica Ag
C0368316|T201|COMP|6399-0|LNC|Entamoeba histolytica Ag|Entamoeba histolytica Ag
C0368317|T201|COMP|5001-3|LNC|Enterococcus sp rRNA|Enterococcus sp rRNA
C0368318|T201|COMP|5839-6|LNC|Enterovirus identified|Enterovirus identified
C0368319|T201|COMP|5840-4|LNC|Enterovirus identified|Enterovirus identified
C0368320|T201|COMP|5841-2|LNC|Enterovirus identified|Enterovirus identified
C0368321|T201|COMP|5842-0|LNC|Enterovirus identified|Enterovirus identified
C0368322|T201|COMP|5843-8|LNC|Enterovirus identified|Enterovirus identified
C0368323|T201|COMP|5002-1|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C0368324|T201|COMP|5003-9|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C0368325|T201|COMP|5004-7|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C0368326|T201|COMP|5005-4|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C0368341|T201|COMP|5162-3|LNC|Fasciola hepatica Ab|Fasciola hepatica Ab
C0368342|T201|COMP|5163-1|LNC|Fasciola sp Ab|Fasciola sp Ab
C0368343|T201|COMP|5165-6|LNC|Filaria Ab|Filaria Ab
C0368344|T201|COMP|6406-3|LNC|Flavivirus identified|Flavivirus identified
C0368345|T201|COMP|5166-4|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C0368346|T201|COMP|5167-2|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C0368347|T201|COMP|6407-1|LNC|Francisella tularensis Ab.IgM|Francisella tularensis Ab.IgM
C0368348|T201|COMP|6408-9|LNC|Francisella tularensis Ag|Francisella tularensis Ag
C0368349|T201|COMP|568-6|LNC|Fungus identified|Fungus identified
C0368350|T201|COMP|569-4|LNC|Fungus identified|Fungus identified
C0368351|T201|COMP|570-2|LNC|Fungus identified|Fungus identified
C0368352|T201|COMP|571-0|LNC|Fungus identified|Fungus identified
C0368353|T201|COMP|572-8|LNC|Fungus identified|Fungus identified
C0368354|T201|COMP|573-6|LNC|Fungus identified|Fungus identified
C0368355|T201|COMP|574-4|LNC|Fungus identified|Fungus identified
C0368356|T201|COMP|575-1|LNC|Fungus identified|Fungus identified
C0368357|T201|COMP|576-9|LNC|Fungus identified|Fungus identified
C0368358|T201|COMP|577-7|LNC|Fungus identified|Fungus identified
C0368359|T201|COMP|6409-7|LNC|Fungus identified|Fungus identified
C0368360|T201|COMP|578-5|LNC|Fungus identified|Fungus identified
C0368361|T201|COMP|579-3|LNC|Fungus identified|Fungus identified
C0368362|T201|COMP|17949-9|LNC|Fungus identified^^^4|Fungus identified^^^4
C0368363|T201|COMP|6410-5|LNC|Gardnerella vaginalis rRNA|Gardnerella vaginalis rRNA
C0368364|T201|COMP|5169-8|LNC|Giardia lamblia Ab|Giardia lamblia Ab
C0368365|T201|COMP|6411-3|LNC|Giardia lamblia Ab.IgG|Giardia lamblia Ab.IgG
C0368366|T201|COMP|6412-1|LNC|Giardia lamblia Ag|Giardia lamblia Ag
C0368367|T201|COMP|6413-9|LNC|Giardia lamblia Ag|Giardia lamblia Ag
C0368368|T201|COMP|5178-9|LNC|Haemophilus influenzae Ab|Haemophilus influenzae Ab
C0368369|T201|COMP|5006-2|LNC|Haemophilus influenzae rRNA|Haemophilus influenzae rRNA
C0368375|T201|COMP|5046-8|LNC|Hantavirus Ab|Hantavirus Ab
C0368376|T201|COMP|587-6|LNC|Helicobacter pylori|Helicobacter pylori
C0368377|T201|COMP|5174-8|LNC|Helicobacter pylori Ab|Helicobacter pylori Ab
C0368378|T201|COMP|6419-6|LNC|Helicobacter pylori Ab|Helicobacter pylori Ab
C0368379|T201|COMP|5175-5|LNC|Helicobacter pylori Ab|Helicobacter pylori Ab
C0368380|T201|COMP|6420-4|LNC|Helicobacter pylori Ab.IgA|Helicobacter pylori Ab.IgA
C0368381|T201|COMP|5176-3|LNC|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C0368382|T201|COMP|5177-1|LNC|Helicobacter pylori Ab.IgM|Helicobacter pylori Ab.IgM
C0368383|T201|COMP|5179-7|LNC|Hepatitis A virus Ab.IgG|Hepatitis A virus Ab.IgG
C0368384|T201|COMP|5180-5|LNC|Hepatitis A virus Ab.IgG|Hepatitis A virus Ab.IgG
C0368385|T201|COMP|5181-3|LNC|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C0368386|T201|COMP|5182-1|LNC|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C0368387|T201|COMP|5183-9|LNC|Hepatitis A virus Ab|Hepatitis A virus Ab
C0368388|T201|COMP|5184-7|LNC|Hepatitis A virus Ab|Hepatitis A virus Ab
C0368389|T201|COMP|5185-4|LNC|Hepatitis B virus core Ab.IgM|Hepatitis B virus core Ab.IgM
C0368390|T201|COMP|5186-2|LNC|Hepatitis B virus core Ab.IgM|Hepatitis B virus core Ab.IgM
C0368391|T201|COMP|5187-0|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C0368392|T201|COMP|5188-8|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C0368393|T201|COMP|5007-0|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C0368394|T201|COMP|5008-8|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C0368395|T201|COMP|5009-6|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C0368400|T201|COMP|6421-2|LNC|Hepatitis B virus rRNA|Hepatitis B virus rRNA
C0368401|T201|COMP|5193-8|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0368402|T201|COMP|5194-6|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0368403|T201|COMP|5195-3|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C0368404|T201|COMP|5196-1|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C0368405|T201|COMP|5197-9|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C0368406|T201|COMP|5198-7|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C0368407|T201|COMP|5199-5|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C0368408|T201|COMP|5010-4|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C0368409|T201|COMP|5011-2|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C0368410|T201|COMP|5012-0|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C0368411|T201|COMP|6422-0|LNC|Hepatitis C virus rRNA|Hepatitis C virus rRNA
C0368412|T201|COMP|5200-1|LNC|Hepatitis D virus Ab|Hepatitis D virus Ab
C0368413|T201|COMP|5201-9|LNC|Hepatitis D virus Ab|Hepatitis D virus Ab
C0368414|T201|COMP|5844-6|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C0368415|T201|COMP|5845-3|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C0368416|T201|COMP|5846-1|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C0368417|T201|COMP|5847-9|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C0368418|T201|COMP|5848-7|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C0368419|T201|COMP|5849-5|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C0368420|T201|COMP|5202-7|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C0368421|T201|COMP|5203-5|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C0368422|T201|COMP|5204-3|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C0368423|T201|COMP|5850-3|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C0368424|T201|COMP|5851-1|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C0368425|T201|COMP|5852-9|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C0368426|T201|COMP|5853-7|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C0368427|T201|COMP|5854-5|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C0368428|T201|COMP|5855-2|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C0368429|T201|COMP|5013-8|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C0368430|T201|COMP|5014-6|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C0368431|T201|COMP|5856-0|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C0368432|T201|COMP|5857-8|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C0368433|T201|COMP|5858-6|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C0368434|T201|COMP|5859-4|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C0368435|T201|COMP|5205-0|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C0368436|T201|COMP|5207-6|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C0368437|T201|COMP|5208-4|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C0368438|T201|COMP|5209-2|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0368439|T201|COMP|5210-0|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C0368440|T201|COMP|5211-8|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C0368441|T201|COMP|5212-6|LNC|Herpes virus 6 Ab.IgM|Herpes virus 6 Ab.IgM
C0368443|T201|COMP|6425-3|LNC|Heterophile Ab|Heterophile Ab
C0368444|T201|COMP|5213-4|LNC|Heterophile Ab|Heterophile Ab
C0368445|T201|COMP|5215-9|LNC|Heterophile Ab|Heterophile Ab
C0368446|T201|COMP|6424-6|LNC|Heterophile Ab|Heterophile Ab
C0368447|T201|COMP|5216-7|LNC|Heterophile Ab after absorption|Heterophile Ab after absorption
C0368448|T201|COMP|6426-1|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0368449|T201|COMP|5218-3|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0368450|T201|COMP|6427-9|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0368451|T201|COMP|5219-1|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0368452|T201|COMP|6428-7|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C0368453|T201|COMP|5015-3|LNC|Histoplasma capsulatum DNA|Histoplasma capsulatum DNA
C0368454|T201|COMP|5016-1|LNC|Histoplasma capsulatum rRNA|Histoplasma capsulatum rRNA
C0368455|T201|COMP|5220-9|LNC|HIV 1 Ab|HIV 1 Ab
C0368456|T201|COMP|5221-7|LNC|HIV 1 Ab|HIV 1 Ab
C0368457|T201|COMP|5222-5|LNC|HIV 1 Ag|HIV 1 Ag
C0368458|T201|COMP|5017-9|LNC|HIV 1 RNA|HIV 1 RNA
C0368459|T201|COMP|5018-7|LNC|HIV 1 RNA|HIV 1 RNA
C0368460|T201|COMP|5223-3|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C0368461|T201|COMP|5224-1|LNC|HIV 2 Ab|HIV 2 Ab
C0368462|T201|COMP|5225-8|LNC|HIV 2 Ab|HIV 2 Ab
C0368463|T201|COMP|6429-5|LNC|HIV identified|HIV identified
C0368464|T201|COMP|6430-3|LNC|HIV identified|HIV identified
C0368465|T201|COMP|6431-1|LNC|HIV identified|HIV identified
C0368466|T201|COMP|6432-9|LNC|HTLV I Ab|HTLV I Ab
C0368467|T201|COMP|6433-7|LNC|HTLV I Ab.IgG|HTLV I Ab.IgG
C0368468|T201|COMP|5226-6|LNC|HTLV I+II Ab|HTLV I+II Ab
C0368469|T201|COMP|5019-5|LNC|HTLV I+II RNA|HTLV I+II RNA
C0368470|T201|COMP|5229-0|LNC|Influenza virus A Ab|Influenza virus A Ab
C0368471|T201|COMP|5860-2|LNC|Influenza virus A Ag|Influenza virus A Ag
C0368472|T201|COMP|5861-0|LNC|Influenza virus A Ag|Influenza virus A Ag
C0368473|T201|COMP|5862-8|LNC|Influenza virus A Ag|Influenza virus A Ag
C0368474|T201|COMP|5863-6|LNC|Influenza virus A Ag|Influenza virus A Ag
C0368475|T201|COMP|6434-5|LNC|Influenza virus A+B Ab|Influenza virus A+B Ab
C0368476|T201|COMP|6435-2|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C0368477|T201|COMP|6436-0|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C0368478|T201|COMP|6437-8|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C0368479|T201|COMP|6438-6|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C0368480|T201|COMP|6439-4|LNC|Influenza virus A+B+C Ag|Influenza virus A+B+C Ag
C0368481|T201|COMP|6440-2|LNC|Influenza virus A+B+C Ag|Influenza virus A+B+C Ag
C0368482|T201|COMP|6441-0|LNC|Influenza virus A+B+C Ag|Influenza virus A+B+C Ag
C0368483|T201|COMP|6442-8|LNC|Influenza virus A+B+C Ag|Influenza virus A+B+C Ag
C0368484|T201|COMP|5230-8|LNC|Influenza virus B Ab|Influenza virus B Ab
C0368485|T201|COMP|5864-4|LNC|Influenza virus B Ag|Influenza virus B Ag
C0368486|T201|COMP|5865-1|LNC|Influenza virus B Ag|Influenza virus B Ag
C0368487|T201|COMP|5866-9|LNC|Influenza virus B Ag|Influenza virus B Ag
C0368488|T201|COMP|5867-7|LNC|Influenza virus B Ag|Influenza virus B Ag
C0368489|T201|COMP|5231-6|LNC|Influenza virus C Ab|Influenza virus C Ab
C0368490|T201|COMP|6443-6|LNC|Lactoferrin|Lactoferrin
C0368491|T201|COMP|6444-4|LNC|Lactoferrin|Lactoferrin
C0368492|T201|COMP|5236-5|LNC|Legionella pneumophila Ab|Legionella pneumophila Ab
C0368493|T201|COMP|5237-3|LNC|Legionella pneumophila Ab|Legionella pneumophila Ab
C0368494|T201|COMP|6445-1|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C0368495|T201|COMP|6446-9|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C0368496|T201|COMP|6447-7|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C0368497|T201|COMP|6448-5|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C0368498|T201|COMP|588-4|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C0368499|T201|COMP|6449-3|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C0368500|T201|COMP|589-2|LNC|Legionella sp identified|Legionella sp identified
C0368501|T201|COMP|590-0|LNC|Legionella sp identified|Legionella sp identified
C0368502|T201|COMP|591-8|LNC|Legionella sp|Legionella sp
C0368503|T201|COMP|592-6|LNC|Legionella sp|Legionella sp
C0368504|T201|COMP|593-4|LNC|Legionella sp identified|Legionella sp identified
C0368505|T201|COMP|6450-1|LNC|Legionella sp Ab|Legionella sp Ab
C0368506|T201|COMP|6451-9|LNC|Legionella sp rRNA|Legionella sp rRNA
C0368507|T201|COMP|5020-3|LNC|Legionella sp rRNA|Legionella sp rRNA
C0368508|T201|COMP|5238-1|LNC|Leishmania sp Ab|Leishmania sp Ab
C0368509|T201|COMP|5239-9|LNC|Leptospira sp Ab|Leptospira sp Ab
C0368510|T201|COMP|6452-7|LNC|Leptospira interrogans Ag|Leptospira interrogans Ag
C0368511|T201|COMP|6453-5|LNC|Leptospira sp identified|Leptospira sp identified
C0368512|T201|COMP|6454-3|LNC|Leptospira sp identified|Leptospira sp identified
C0368513|T201|COMP|6455-0|LNC|Leptospira sp identified|Leptospira sp identified
C0368514|T201|COMP|594-2|LNC|Leptospira sp identified|Leptospira sp identified
C0368515|T201|COMP|5240-7|LNC|Listeria monocytogenes Ab|Listeria monocytogenes Ab
C0368516|T201|COMP|6456-8|LNC|Listeria monocytogenes Ab|Listeria monocytogenes Ab
C0368517|T201|COMP|5021-1|LNC|Listeria monocytogenes rRNA|Listeria monocytogenes rRNA
C0368519|T201|COMP|5241-5|LNC|Lymphocytic choriomeningitis virus Ab|Lymphocytic choriomeningitis virus Ab
C0368520|T201|COMP|6458-4|LNC|Lymphocytic choriomeningitis virus Ab|Lymphocytic choriomeningitis virus Ab
C0368521|T201|COMP|5242-3|LNC|Measles virus Ab|Measles virus Ab
C0368522|T201|COMP|5243-1|LNC|Measles virus Ab|Measles virus Ab
C0368523|T201|COMP|5244-9|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0368524|T201|COMP|5245-6|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C0368525|T201|COMP|595-9|LNC|Bacteria identified|Bacteria identified
C0368526|T201|COMP|596-7|LNC|Bacteria identified|Bacteria identified
C0368527|T201|COMP|597-5|LNC|Bacteria identified|Bacteria identified
C0368528|T201|COMP|598-3|LNC|Bacteria identified|Bacteria identified
C0368529|T201|COMP|599-1|LNC|Bacteria identified|Bacteria identified
C0368530|T201|COMP|600-7|LNC|Bacteria identified|Bacteria identified
C0368531|T201|COMP|601-5|LNC|Fungus identified|Fungus identified
C0368532|T201|COMP|17877-2|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0368533|T201|COMP|17941-6|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0368534|T201|COMP|17882-2|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0368535|T201|COMP|605-6|LNC|Bacteria identified|Bacteria identified
C0368536|T201|COMP|606-4|LNC|Bacteria identified|Bacteria identified
C0368537|T201|COMP|607-2|LNC|Bacteria identified|Bacteria identified
C0368538|T201|COMP|608-0|LNC|Bacteria identified|Bacteria identified
C0368539|T201|COMP|609-8|LNC|Bacteria identified|Bacteria identified
C0368540|T201|COMP|610-6|LNC|Bacteria identified|Bacteria identified
C0368541|T201|COMP|611-4|LNC|Bacteria identified|Bacteria identified
C0368542|T201|COMP|6459-2|LNC|Bacteria identified|Bacteria identified
C0368543|T201|COMP|612-2|LNC|Bacterial strain|Bacterial strain
C0368544|T201|COMP|613-0|LNC|Fungal strain|Fungal strain
C0368545|T201|COMP|614-8|LNC|Mycobacterial strain|Mycobacterial strain
C0368546|T201|COMP|615-5|LNC|Viral strain|Viral strain
C0368547|T201|COMP|17946-5|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0368548|T201|COMP|617-1|LNC|Bacteria identified|Bacteria identified
C0368549|T201|COMP|618-9|LNC|Bacteria identified|Bacteria identified
C0368550|T201|COMP|17963-0|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0368551|T201|COMP|620-5|LNC|Bacteria identified|Bacteria identified
C0368552|T201|COMP|621-3|LNC|Bacteria identified|Bacteria identified
C0368553|T201|COMP|17897-0|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0368555|T201|COMP|624-7|LNC|Bacteria identified|Bacteria identified
C0368556|T201|COMP|6460-0|LNC|Bacteria identified|Bacteria identified
C0368557|T201|COMP|6461-8|LNC|Bacteria identified|Bacteria identified
C0368558|T201|COMP|17968-9|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0368559|T201|COMP|626-2|LNC|Bacteria identified|Bacteria identified
C0368560|T201|COMP|17908-5|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0368561|T201|COMP|17924-2|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0368562|T201|COMP|629-6|LNC|Bacteria identified|Bacteria identified
C0368563|T201|COMP|630-4|LNC|Bacteria identified|Bacteria identified
C0368564|T201|COMP|631-2|LNC|Bacteria identified|Bacteria identified
C0368565|T201|COMP|1817-6|LNC|Alpha ketoglutarate|Alpha ketoglutarate
C0368566|T201|COMP|2983-5|LNC|Terminal deoxyribonucleotidyl transferase|Terminal deoxyribonucleotidyl transferase
C0368567|T201|COMP|5206-8|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C0369164|T201|COMP|12208-5|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0369741|T201|COMP|12238-2|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0481909|T201|COMP|1283-1|LNC|P NOS Ag|P NOS Ag
C0481910|T201|COMP|1284-9|LNC|P NOS Ag|P NOS Ag
C0481911|T201|COMP|1285-6|LNC|P NOS Ag|P NOS Ag
C0481912|T201|COMP|1317-7|LNC|S Ab|S Ab
C0481913|T201|COMP|1318-5|LNC|S Ag|S Ag
C0481914|T201|COMP|1319-3|LNC|S Ag|S Ag
C0481915|T201|COMP|1320-1|LNC|S Ag|S Ag
C0481916|T201|COMP|2-6|LNC|Almecillin|Almecillin
C0481917|T201|COMP|7-5|LNC|Amdinocillin|Amdinocillin
C0481918|T201|COMP|11-7|LNC|Amikacin|Amikacin
C0481919|T201|COMP|15-8|LNC|Amoxicillin|Amoxicillin
C0481920|T201|COMP|19-0|LNC|Amoxicillin+Clavulanate|Amoxicillin+Clavulanate
C0481921|T201|COMP|23-2|LNC|Amphotericin B|Amphotericin B
C0481922|T201|COMP|27-3|LNC|Ampicillin|Ampicillin
C0481923|T201|COMP|31-5|LNC|Ampicillin+Sulbactam|Ampicillin+Sulbactam
C0481924|T201|COMP|35-6|LNC|Azithromycin|Azithromycin
C0481925|T201|COMP|39-8|LNC|Azlocillin|Azlocillin
C0481926|T201|COMP|43-0|LNC|Aztreonam|Aztreonam
C0481927|T201|COMP|47-1|LNC|Bacampicillin|Bacampicillin
C0481928|T201|COMP|51-3|LNC|Butirosin|Butirosin
C0481929|T201|COMP|55-4|LNC|Capreomycin|Capreomycin
C0481930|T201|COMP|59-6|LNC|Carbenicillin|Carbenicillin
C0481931|T201|COMP|63-8|LNC|Cefadroxil|Cefadroxil
C0481932|T201|COMP|67-9|LNC|Cefamandole|Cefamandole
C0481933|T201|COMP|71-1|LNC|Cefatrizine|Cefatrizine
C0481934|T201|COMP|75-2|LNC|ceFAZolin|ceFAZolin
C0481935|T201|COMP|79-4|LNC|Cefixime|Cefixime
C0481936|T201|COMP|83-6|LNC|Cefaclor|Cefaclor
C0481937|T201|COMP|84-4|LNC|Cefaclor|Cefaclor
C0481938|T201|COMP|85-1|LNC|Cefaclor|Cefaclor
C0481939|T201|COMP|86-9|LNC|Cefaclor|Cefaclor
C0481940|T201|COMP|87-7|LNC|Cefmetazole|Cefmetazole
C0481941|T201|COMP|91-9|LNC|Cefodizime|Cefodizime
C0481942|T201|COMP|95-0|LNC|Cefonicid|Cefonicid
C0481943|T201|COMP|99-2|LNC|Cefoperazone|Cefoperazone
C0481944|T201|COMP|103-2|LNC|Ceforanide|Ceforanide
C0481945|T201|COMP|107-3|LNC|Cefotaxime|Cefotaxime
C0481946|T201|COMP|111-5|LNC|cefoTEtan|cefoTEtan
C0481947|T201|COMP|115-6|LNC|cefOXitin|cefOXitin
C0481948|T201|COMP|119-8|LNC|Cefpodoxime|Cefpodoxime
C0481949|T201|COMP|123-0|LNC|Cefprozil|Cefprozil
C0481950|T201|COMP|127-1|LNC|Cefsulodin|Cefsulodin
C0481951|T201|COMP|132-1|LNC|cefTAZidime|cefTAZidime
C0481952|T201|COMP|136-2|LNC|Ceftizoxime|Ceftizoxime
C0481953|T201|COMP|140-4|LNC|cefTRIAXone|cefTRIAXone
C0481954|T201|COMP|144-6|LNC|Cefuroxime.parenteral|Cefuroxime.parenteral
C0481955|T201|COMP|148-7|LNC|Cephalexin|Cephalexin
C0481956|T201|COMP|152-9|LNC|Cephaloglycin|Cephaloglycin
C0481957|T201|COMP|156-0|LNC|Cephaloridine|Cephaloridine
C0481958|T201|COMP|160-2|LNC|Cephalothin|Cephalothin
C0481959|T201|COMP|164-4|LNC|Cephapirin|Cephapirin
C0481960|T201|COMP|168-5|LNC|Cephradine|Cephradine
C0481961|T201|COMP|172-7|LNC|Chloramphenicol|Chloramphenicol
C0481962|T201|COMP|176-8|LNC|Chlortetracycline|Chlortetracycline
C0481963|T201|COMP|180-0|LNC|Cinoxacin|Cinoxacin
C0481964|T201|COMP|184-2|LNC|Ciprofloxacin|Ciprofloxacin
C0481965|T201|COMP|188-3|LNC|Clarithromycin|Clarithromycin
C0481966|T201|COMP|192-5|LNC|Clindamycin|Clindamycin
C0481967|T201|COMP|196-6|LNC|Cloxacillin|Cloxacillin
C0481968|T201|COMP|200-6|LNC|Colistimethate|Colistimethate
C0481969|T201|COMP|204-8|LNC|Colistin|Colistin
C0481970|T201|COMP|208-9|LNC|Cyclacillin|Cyclacillin
C0481971|T201|COMP|212-1|LNC|cycloSERINE|cycloSERINE
C0481972|T201|COMP|216-2|LNC|Demeclocycline|Demeclocycline
C0481973|T201|COMP|220-4|LNC|Dicloxacillin|Dicloxacillin
C0481974|T201|COMP|224-6|LNC|Doxycycline|Doxycycline
C0481975|T201|COMP|228-7|LNC|Enoxacin|Enoxacin
C0481976|T201|COMP|232-9|LNC|Erythromycin|Erythromycin
C0481977|T201|COMP|236-0|LNC|Erythromycin+sulfiSOXAZOLE|Erythromycin+sulfiSOXAZOLE
C0481978|T201|COMP|240-2|LNC|Ethambutol|Ethambutol
C0481979|T201|COMP|244-4|LNC|Floxacillin|Floxacillin
C0481980|T201|COMP|248-5|LNC|Fluconazole|Fluconazole
C0481981|T201|COMP|252-7|LNC|5-Fluorocytosine|5-Fluorocytosine
C0481982|T201|COMP|257-6|LNC|Framycetin|Framycetin
C0481983|T201|COMP|261-8|LNC|Fusidate|Fusidate
C0481984|T201|COMP|266-7|LNC|Gentamicin|Gentamicin
C0481985|T201|COMP|270-9|LNC|Gramicidin D|Gramicidin D
C0481986|T201|COMP|274-1|LNC|Hetacillin|Hetacillin
C0481987|T201|COMP|278-2|LNC|Imipenem|Imipenem
C0481988|T201|COMP|282-4|LNC|Imipenem+Cilastatin|Imipenem+Cilastatin
C0481989|T201|COMP|286-5|LNC|Isoniazid|Isoniazid
C0481990|T201|COMP|290-7|LNC|Kanamycin|Kanamycin
C0481991|T201|COMP|294-9|LNC|Ketoconazole|Ketoconazole
C0481992|T201|COMP|298-0|LNC|Lincomycin|Lincomycin
C0481993|T201|COMP|302-0|LNC|Lomefloxacin|Lomefloxacin
C0481994|T201|COMP|306-1|LNC|Loracarbef|Loracarbef
C0481995|T201|COMP|310-3|LNC|Lymecycline|Lymecycline
C0481996|T201|COMP|314-5|LNC|Meclocycline|Meclocycline
C0481997|T201|COMP|318-6|LNC|Methacycline|Methacycline
C0481998|T201|COMP|322-8|LNC|Methicillin|Methicillin
C0481999|T201|COMP|326-9|LNC|metroNIDAZOLE|metroNIDAZOLE
C0482000|T201|COMP|330-1|LNC|Mezlocillin|Mezlocillin
C0482001|T201|COMP|334-3|LNC|Minocycline|Minocycline
C0482002|T201|COMP|338-4|LNC|Miocamycin|Miocamycin
C0482003|T201|COMP|342-6|LNC|Moxalactam|Moxalactam
C0482004|T201|COMP|346-7|LNC|Nafcillin|Nafcillin
C0482005|T201|COMP|350-9|LNC|Nalidixate|Nalidixate
C0482006|T201|COMP|354-1|LNC|Neomycin|Neomycin
C0482007|T201|COMP|358-2|LNC|Netilmicin|Netilmicin
C0482008|T201|COMP|362-4|LNC|Nitrofurantoin|Nitrofurantoin
C0482009|T201|COMP|366-5|LNC|Norfloxacin|Norfloxacin
C0482010|T201|COMP|370-7|LNC|Novobiocin|Novobiocin
C0482011|T201|COMP|374-9|LNC|Ofloxacin|Ofloxacin
C0482012|T201|COMP|378-0|LNC|Oleandomycin|Oleandomycin
C0482013|T201|COMP|382-2|LNC|Oxacillin|Oxacillin
C0482014|T201|COMP|386-3|LNC|Oxytetracycline|Oxytetracycline
C0482015|T201|COMP|391-3|LNC|Penicillin G|Penicillin G
C0482016|T201|COMP|395-4|LNC|Penicillin V|Penicillin V
C0482017|T201|COMP|399-6|LNC|Phenethicillin|Phenethicillin
C0482018|T201|COMP|403-6|LNC|Pipemidate|Pipemidate
C0482019|T201|COMP|407-7|LNC|Piperacillin|Piperacillin
C0482020|T201|COMP|411-9|LNC|Piperacillin+Tazobactam|Piperacillin+Tazobactam
C0482021|T201|COMP|415-0|LNC|Pivampicillin|Pivampicillin
C0482022|T201|COMP|419-2|LNC|Polymyxin B|Polymyxin B
C0482023|T201|COMP|423-4|LNC|Pyrazinamide|Pyrazinamide
C0482024|T201|COMP|427-5|LNC|rifAMPin|rifAMPin
C0482025|T201|COMP|431-7|LNC|Ristocetin|Ristocetin
C0482026|T201|COMP|435-8|LNC|Rolitetracycline|Rolitetracycline
C0482027|T201|COMP|439-0|LNC|Rosoxacin|Rosoxacin
C0482028|T201|COMP|443-2|LNC|Roxithromycin|Roxithromycin
C0482029|T201|COMP|447-3|LNC|Sisomicin|Sisomicin
C0482030|T201|COMP|451-5|LNC|Spectinomycin|Spectinomycin
C0482031|T201|COMP|455-6|LNC|Spiramycin|Spiramycin
C0482032|T201|COMP|459-8|LNC|Streptomycin|Streptomycin
C0482033|T201|COMP|463-0|LNC|sulfADIAZINE|sulfADIAZINE
C0482034|T201|COMP|467-1|LNC|Sulfamethoxazole|Sulfamethoxazole
C0482035|T201|COMP|471-3|LNC|sulfiSOXAZOLE|sulfiSOXAZOLE
C0482036|T201|COMP|475-4|LNC|Sulfonamide|Sulfonamide
C0482037|T201|COMP|479-6|LNC|Talampicillin|Talampicillin
C0482038|T201|COMP|483-8|LNC|Teicoplanin|Teicoplanin
C0482039|T201|COMP|487-9|LNC|Temafloxacin|Temafloxacin
C0482040|T201|COMP|491-1|LNC|Temocillin|Temocillin
C0482041|T201|COMP|495-2|LNC|Tetracycline|Tetracycline
C0482042|T201|COMP|499-4|LNC|Ticarcillin|Ticarcillin
C0482043|T201|COMP|503-3|LNC|Ticarcillin+Clavulanate|Ticarcillin+Clavulanate
C0482044|T201|COMP|507-4|LNC|Tobramycin|Tobramycin
C0482045|T201|COMP|511-6|LNC|Trimethoprim|Trimethoprim
C0482046|T201|COMP|515-7|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0482047|T201|COMP|519-9|LNC|Troleandomycin|Troleandomycin
C0482048|T201|COMP|523-1|LNC|Vancomycin|Vancomycin
C0482049|T201|COMP|527-2|LNC|Viomycin|Viomycin
C0482050|T201|COMP|6016-0|LNC|Corticotropin Ab.IgE|Corticotropin Ab.IgE
C0482051|T201|COMP|6046-7|LNC|Juglans nigra pollen Ab.IgE|Juglans nigra pollen Ab.IgE
C0482052|T201|COMP|6064-0|LNC|Cat epithelium Ab.IgE|Cat epithelium Ab.IgE
C0482054|T201|COMP|6121-8|LNC|Fusarium moniliforme Ab.IgE|Fusarium moniliforme Ab.IgE
C0482055|T201|COMP|6124-2|LNC|Ambrosia trifida Ab.IgE|Ambrosia trifida Ab.IgE
C0482056|T201|COMP|6144-0|LNC|Tabanus spp Ab.IgE|Tabanus spp Ab.IgE
C0482057|T201|COMP|6208-3|LNC|Carya illinoinensis nut Ab.IgE|Carya illinoinensis nut Ab.IgE
C0482059|T201|COMP|6248-9|LNC|Glycine max Ab.IgE|Glycine max Ab.IgE
C0482060|T201|COMP|6253-9|LNC|Midge stinging Ab.IgE|Midge stinging Ab.IgE
C0482061|T201|COMP|6258-8|LNC|Helianthus annuus seed Ab.IgE|Helianthus annuus seed Ab.IgE
C0482062|T201|COMP|6260-4|LNC|Liquidambar styraciflua Ab.IgE|Liquidambar styraciflua Ab.IgE
C0482063|T201|COMP|815-1|LNC|A Ab|A Ab
C0482064|T201|COMP|816-9|LNC|A Ab|A Ab
C0482065|T201|COMP|817-7|LNC|A Ab|A Ab
C0482066|T201|COMP|818-5|LNC|A Ag|A Ag
C0482067|T201|COMP|819-3|LNC|A Ag|A Ag
C0482068|T201|COMP|820-1|LNC|A Ag|A Ag
C0482069|T201|COMP|821-9|LNC|A little u super little a Ab|A little u super little a Ab
C0482070|T201|COMP|822-7|LNC|A little u super little a Ab|A little u super little a Ab
C0482071|T201|COMP|823-5|LNC|A little u super little a Ab|A little u super little a Ab
C0482072|T201|COMP|824-3|LNC|A little u super little a Ag|A little u super little a Ag
C0482073|T201|COMP|825-0|LNC|A little u super little a Ag|A little u super little a Ag
C0482074|T201|COMP|826-8|LNC|A little u super little a Ag|A little u super little a Ag
C0482075|T201|COMP|827-6|LNC|Am Ag|Am Ag
C0482076|T201|COMP|828-4|LNC|Am Ag|Am Ag
C0482077|T201|COMP|829-2|LNC|Am Ag|Am Ag
C0482078|T201|COMP|830-0|LNC|A variant subtype|A variant subtype
C0482079|T201|COMP|831-8|LNC|A variant subtype|A variant subtype
C0482080|T201|COMP|832-6|LNC|A variant subtype|A variant subtype
C0482081|T201|COMP|833-4|LNC|A variant NOS Ag|A variant NOS Ag
C0482082|T201|COMP|834-2|LNC|A variant NOS Ag|A variant NOS Ag
C0482083|T201|COMP|835-9|LNC|A variant subtype|A variant subtype
C0482084|T201|COMP|836-7|LNC|Ax Ag|Ax Ag
C0482085|T201|COMP|837-5|LNC|Ax Ag|Ax Ag
C0482086|T201|COMP|838-3|LNC|Ax Ag|Ax Ag
C0482087|T201|COMP|839-1|LNC|A1 Ab|A1 Ab
C0482088|T201|COMP|840-9|LNC|A1 Ab|A1 Ab
C0482089|T201|COMP|841-7|LNC|A1 Ab|A1 Ab
C0482090|T201|COMP|842-5|LNC|A1 Ag|A1 Ag
C0482091|T201|COMP|843-3|LNC|A1 Ag|A1 Ag
C0482092|T201|COMP|844-1|LNC|A1 Ag|A1 Ag
C0482093|T201|COMP|845-8|LNC|A1 B Ab|A1 B Ab
C0482094|T201|COMP|846-6|LNC|A1 B Ab|A1 B Ab
C0482095|T201|COMP|847-4|LNC|A1 B Ab|A1 B Ab
C0482096|T201|COMP|848-2|LNC|A1 B Ag|A1 B Ag
C0482097|T201|COMP|849-0|LNC|A1 B Ag|A1 B Ag
C0482098|T201|COMP|850-8|LNC|A1 B Ag|A1 B Ag
C0482099|T201|COMP|851-6|LNC|A2 Ab|A2 Ab
C0482100|T201|COMP|852-4|LNC|A2 Ab|A2 Ab
C0482101|T201|COMP|853-2|LNC|A2 Ab|A2 Ab
C0482102|T201|COMP|854-0|LNC|A2 Ag|A2 Ag
C0482103|T201|COMP|855-7|LNC|A2 Ag|A2 Ag
C0482104|T201|COMP|856-5|LNC|A2 Ag|A2 Ag
C0482105|T201|COMP|857-3|LNC|A2 B Ab|A2 B Ab
C0482106|T201|COMP|858-1|LNC|A2 B Ab|A2 B Ab
C0482107|T201|COMP|859-9|LNC|A2 B Ab|A2 B Ab
C0482108|T201|COMP|860-7|LNC|A2 B Ag|A2 B Ag
C0482109|T201|COMP|861-5|LNC|A2 B Ag|A2 B Ag
C0482110|T201|COMP|862-3|LNC|A2 B Ag|A2 B Ag
C0482111|T201|COMP|863-1|LNC|A3 Ab|A3 Ab
C0482112|T201|COMP|864-9|LNC|A3 Ab|A3 Ab
C0482113|T201|COMP|865-6|LNC|A3 Ab|A3 Ab
C0482114|T201|COMP|866-4|LNC|A3 Ag|A3 Ag
C0482115|T201|COMP|867-2|LNC|A3 Ag|A3 Ag
C0482116|T201|COMP|868-0|LNC|A3 Ag|A3 Ag
C0482117|T201|COMP|869-8|LNC|A3 B Ab|A3 B Ab
C0482118|T201|COMP|870-6|LNC|A3 B Ab|A3 B Ab
C0482119|T201|COMP|871-4|LNC|A3 B Ab|A3 B Ab
C0482120|T201|COMP|872-2|LNC|A3 B Ag|A3 B Ag
C0482121|T201|COMP|873-0|LNC|A3 B Ag|A3 B Ag
C0482122|T201|COMP|874-8|LNC|A3 B Ag|A3 B Ag
C0482123|T201|COMP|875-5|LNC|A,B Ab|A,B Ab
C0482124|T201|COMP|876-3|LNC|A,B Ab|A,B Ab
C0482125|T201|COMP|877-1|LNC|A,B Ab|A,B Ab
C0482126|T201|COMP|878-9|LNC|A,B Ag|A,B Ag
C0482127|T201|COMP|879-7|LNC|A,B Ag|A,B Ag
C0482128|T201|COMP|880-5|LNC|A,B Ag|A,B Ag
C0482129|T201|COMP|881-3|LNC|ABO & Rh group|ABO & Rh group
C0482130|T201|COMP|882-1|LNC|ABO & Rh group|ABO & Rh group
C0482131|T201|COMP|883-9|LNC|ABO group|ABO group
C0482132|T201|COMP|885-4|LNC|Am Ab|Am Ab
C0482133|T201|COMP|886-2|LNC|Am Ab|Am Ab
C0482134|T201|COMP|887-0|LNC|Am Ab|Am Ab
C0482136|T201|COMP|889-6|LNC|Blood group antibodies identified|Blood group antibodies identified
C0482137|T201|COMP|891-2|LNC|Blood group antibody screen.cell I|Blood group antibody screen.cell I
C0482138|T201|COMP|892-0|LNC|Blood group antibody screen.cell III|Blood group antibody screen.cell III
C0482139|T201|COMP|905-0|LNC|Blood group antigens absent|Blood group antigens absent
C0482140|T201|COMP|5934-5|LNC|Blood group antigens absent|Blood group antigens absent
C0482141|T201|COMP|907-6|LNC|Blood group antigens present|Blood group antigens present
C0482142|T201|COMP|906-8|LNC|Blood group antigens present|Blood group antigens present
C0482143|T201|COMP|908-4|LNC|Ax Ab|Ax Ab
C0482144|T201|COMP|909-2|LNC|Ax Ab|Ax Ab
C0482145|T201|COMP|910-0|LNC|Ax Ab|Ax Ab
C0482146|T201|COMP|911-8|LNC|B Ab|B Ab
C0482147|T201|COMP|912-6|LNC|B Ab|B Ab
C0482148|T201|COMP|913-4|LNC|B Ab|B Ab
C0482149|T201|COMP|914-2|LNC|B Ag|B Ag
C0482150|T201|COMP|915-9|LNC|B Ag|B Ag
C0482151|T201|COMP|916-7|LNC|B Ag|B Ag
C0482152|T201|COMP|917-5|LNC|B variant subtype Ab|B variant subtype Ab
C0482153|T201|COMP|918-3|LNC|B variant subtype Ab|B variant subtype Ab
C0482154|T201|COMP|919-1|LNC|B variant subtype Ab|B variant subtype Ab
C0482155|T201|COMP|920-9|LNC|B variant NOS Ag|B variant NOS Ag
C0482156|T201|COMP|921-7|LNC|B variant NOS Ag|B variant NOS Ag
C0482157|T201|COMP|922-5|LNC|B variant NOS Ag|B variant NOS Ag
C0482158|T201|COMP|933-2|LNC|Blood product type|Blood product type
C0482159|T201|COMP|937-3|LNC|Bombay Ab|Bombay Ab
C0482160|T201|COMP|938-1|LNC|Bombay Ab|Bombay Ab
C0482161|T201|COMP|939-9|LNC|Bombay Ab|Bombay Ab
C0482162|T201|COMP|940-7|LNC|Bombay Ag|Bombay Ag
C0482163|T201|COMP|941-5|LNC|Bombay Ag|Bombay Ag
C0482164|T201|COMP|942-3|LNC|Bombay Ag|Bombay Ag
C0482165|T201|COMP|949-8|LNC|C little e Ab|C little e Ab
C0482166|T201|COMP|950-6|LNC|C little e Ab|C little e Ab
C0482167|T201|COMP|951-4|LNC|C little e Ab|C little e Ab
C0482168|T201|COMP|952-2|LNC|C little e Ag|C little e Ag
C0482169|T201|COMP|953-0|LNC|C little e Ag|C little e Ag
C0482170|T201|COMP|954-8|LNC|C little e Ag|C little e Ag
C0482171|T201|COMP|955-5|LNC|C little w Ab|C little w Ab
C0482172|T201|COMP|956-3|LNC|C little w Ab|C little w Ab
C0482173|T201|COMP|957-1|LNC|C little w Ab|C little w Ab
C0482174|T201|COMP|958-9|LNC|C little w Ag|C little w Ag
C0482175|T201|COMP|959-7|LNC|C little w Ag|C little w Ag
C0482176|T201|COMP|960-5|LNC|C little w Ag|C little w Ag
C0482177|T201|COMP|961-3|LNC|C little x Ab|C little x Ab
C0482178|T201|COMP|962-1|LNC|C little x Ab|C little x Ab
C0482179|T201|COMP|963-9|LNC|C little x Ab|C little x Ab
C0482180|T201|COMP|964-7|LNC|C little x Ag|C little x Ag
C0482181|T201|COMP|965-4|LNC|C little x Ag|C little x Ag
C0482182|T201|COMP|966-2|LNC|C little x Ag|C little x Ag
C0482183|T201|COMP|979-5|LNC|D little i super little a Ab|D little i super little a Ab
C0482184|T201|COMP|980-3|LNC|D little i super little a Ab|D little i super little a Ab
C0482185|T201|COMP|981-1|LNC|D little i super little a Ab|D little i super little a Ab
C0482186|T201|COMP|982-9|LNC|D little i super little a Ag|D little i super little a Ag
C0482187|T201|COMP|983-7|LNC|D little i super little a Ag|D little i super little a Ag
C0482188|T201|COMP|984-5|LNC|D little i super little a Ag|D little i super little a Ag
C0482189|T201|COMP|985-2|LNC|D little i super little b Ab|D little i super little b Ab
C0482190|T201|COMP|986-0|LNC|D little i super little b Ab|D little i super little b Ab
C0482191|T201|COMP|987-8|LNC|D little i super little b Ab|D little i super little b Ab
C0482192|T201|COMP|988-6|LNC|D little i super little b Ag|D little i super little b Ag
C0482193|T201|COMP|989-4|LNC|D little i super little b Ag|D little i super little b Ag
C0482194|T201|COMP|990-2|LNC|D little i super little b Ag|D little i super little b Ag
C0482195|T201|COMP|991-0|LNC|D little o super little a Ab|D little o super little a Ab
C0482196|T201|COMP|992-8|LNC|D little o super little a Ab|D little o super little a Ab
C0482197|T201|COMP|993-6|LNC|D little o super little a Ab|D little o super little a Ab
C0482198|T201|COMP|994-4|LNC|D little o super little a Ag|D little o super little a Ag
C0482199|T201|COMP|995-1|LNC|D little o super little a Ag|D little o super little a Ag
C0482200|T201|COMP|996-9|LNC|D little o super little a Ag|D little o super little a Ag
C0482201|T201|COMP|970-4|LNC|D little u Ag|D little u Ag
C0482202|T201|COMP|971-2|LNC|D little u Ag|D little u Ag
C0482203|T201|COMP|972-0|LNC|D little u Ag|D little u Ag
C0482204|T201|COMP|973-8|LNC|D Ab|D Ab
C0482205|T201|COMP|974-6|LNC|D Ab|D Ab
C0482206|T201|COMP|1306-0|LNC|D NOS Ab|D NOS Ab
C0482207|T201|COMP|976-1|LNC|D Ag|D Ag
C0482208|T201|COMP|977-9|LNC|D Ag|D Ag
C0482209|T201|COMP|978-7|LNC|D Ag|D Ag
C0482210|T201|COMP|997-7|LNC|DBG Ag|DBG Ag
C0482211|T201|COMP|998-5|LNC|DBG Ag|DBG Ag
C0482212|T201|COMP|999-3|LNC|DBG Ag|DBG Ag
C0482213|T201|COMP|1000-9|LNC|DBG Ab|DBG Ab
C0482214|T201|COMP|1001-7|LNC|DBG Ab|DBG Ab
C0482215|T201|COMP|1002-5|LNC|DBG Ab|DBG Ab
C0482217|T201|COMP|1006-6|LNC|Direct antiglobulin test.IgG specific reagent|Direct antiglobulin test.IgG specific reagent
C0482218|T201|COMP|1007-4|LNC|Direct antiglobulin test.poly specific reagent|Direct antiglobulin test.poly specific reagent
C0482219|T201|COMP|1010-8|LNC|E super little w Ab|E super little w Ab
C0482220|T201|COMP|1011-6|LNC|E super little w Ab|E super little w Ab
C0482221|T201|COMP|1012-4|LNC|E super little w Ab|E super little w Ab
C0482222|T201|COMP|1013-2|LNC|E super little w Ag|E super little w Ag
C0482223|T201|COMP|1014-0|LNC|E super little w Ag|E super little w Ag
C0482224|T201|COMP|1015-7|LNC|E super little w Ag|E super little w Ag
C0482225|T201|COMP|1022-3|LNC|F little y super little a Ab|F little y super little a Ab
C0482226|T201|COMP|1023-1|LNC|F little y super little a Ab|F little y super little a Ab
C0482227|T201|COMP|1024-9|LNC|F little y super little a Ab|F little y super little a Ab
C0482228|T201|COMP|1025-6|LNC|F little y super little a Ag|F little y super little a Ag
C0482229|T201|COMP|1026-4|LNC|F little y super little a Ag|F little y super little a Ag
C0482230|T201|COMP|1027-2|LNC|F little y super little a Ag|F little y super little a Ag
C0482231|T201|COMP|1028-0|LNC|F little y super little b Ab|F little y super little b Ab
C0482232|T201|COMP|1029-8|LNC|F little y super little b Ab|F little y super little b Ab
C0482233|T201|COMP|1030-6|LNC|F little y super little b Ab|F little y super little b Ab
C0482234|T201|COMP|1031-4|LNC|F little y super little b Ag|F little y super little b Ag
C0482235|T201|COMP|1032-2|LNC|F little y super little b Ag|F little y super little b Ag
C0482236|T201|COMP|1033-0|LNC|F little y super little b Ag|F little y super little b Ag
C0482237|T201|COMP|1036-3|LNC|G Ab|G Ab
C0482238|T201|COMP|1037-1|LNC|G Ab|G Ab
C0482239|T201|COMP|1038-9|LNC|G Ab|G Ab
C0482240|T201|COMP|1039-7|LNC|G Ag|G Ag
C0482241|T201|COMP|1040-5|LNC|G Ag|G Ag
C0482242|T201|COMP|1041-3|LNC|G Ag|G Ag
C0482243|T201|COMP|1042-1|LNC|H Ab|H Ab
C0482244|T201|COMP|1043-9|LNC|H Ab|H Ab
C0482245|T201|COMP|1044-7|LNC|H Ab|H Ab
C0482246|T201|COMP|1048-8|LNC|H NOS Ag|H NOS Ag
C0482247|T201|COMP|1049-6|LNC|H NOS Ag|H NOS Ag
C0482248|T201|COMP|1050-4|LNC|H NOS Ag|H NOS Ag
C0482249|T201|COMP|1052-0|LNC|I (int) subtype|I (int) subtype
C0482250|T201|COMP|1053-8|LNC|I (int) subtype|I (int) subtype
C0482251|T201|COMP|1054-6|LNC|I (int) subtype|I (int) subtype
C0482252|T201|COMP|1055-3|LNC|I (int) subtype|I (int) subtype
C0482253|T201|COMP|1056-1|LNC|I (int) subtype|I (int) subtype
C0482254|T201|COMP|1057-9|LNC|I (int) subtype|I (int) subtype
C0482255|T201|COMP|1067-8|LNC|J little k super little a Ab|J little k super little a Ab
C0482256|T201|COMP|1068-6|LNC|J little k super little a Ab|J little k super little a Ab
C0482257|T201|COMP|1069-4|LNC|J little k super little a Ab|J little k super little a Ab
C0482258|T201|COMP|1070-2|LNC|J little k super little a Ag|J little k super little a Ag
C0482259|T201|COMP|1071-0|LNC|J little k super little a Ag|J little k super little a Ag
C0482260|T201|COMP|1072-8|LNC|J little k super little a Ag|J little k super little a Ag
C0482261|T201|COMP|1073-6|LNC|J little k super little b Ab|J little k super little b Ab
C0482262|T201|COMP|1074-4|LNC|J little k super little b Ab|J little k super little b Ab
C0482263|T201|COMP|1075-1|LNC|J little k super little b Ab|J little k super little b Ab
C0482264|T201|COMP|1076-9|LNC|J little k super little b Ag|J little k super little b Ag
C0482265|T201|COMP|1077-7|LNC|J little k super little b Ag|J little k super little b Ag
C0482266|T201|COMP|1078-5|LNC|J little k super little b Ag|J little k super little b Ag
C0482267|T201|COMP|1079-3|LNC|J little s super little a Ab|J little s super little a Ab
C0482268|T201|COMP|1080-1|LNC|J little s super little a Ab|J little s super little a Ab
C0482269|T201|COMP|1081-9|LNC|J little s super little a Ab|J little s super little a Ab
C0482270|T201|COMP|1082-7|LNC|J little s super little a Ag|J little s super little a Ag
C0482271|T201|COMP|1083-5|LNC|J little s super little a Ag|J little s super little a Ag
C0482272|T201|COMP|1084-3|LNC|J little s super little a Ag|J little s super little a Ag
C0482273|T201|COMP|1085-0|LNC|J little s super little b Ab|J little s super little b Ab
C0482274|T201|COMP|1086-8|LNC|J little s super little b Ab|J little s super little b Ab
C0482275|T201|COMP|1087-6|LNC|J little s super little b Ab|J little s super little b Ab
C0482276|T201|COMP|1088-4|LNC|J little s super little b Ag|J little s super little b Ag
C0482277|T201|COMP|1089-2|LNC|J little s super little b Ag|J little s super little b Ag
C0482278|T201|COMP|1090-0|LNC|J little s super little b Ag|J little s super little b Ag
C0482279|T201|COMP|1097-5|LNC|K little p super little a Ab|K little p super little a Ab
C0482280|T201|COMP|1098-3|LNC|K little p super little a Ab|K little p super little a Ab
C0482281|T201|COMP|1099-1|LNC|K little p super little a Ab|K little p super little a Ab
C0482282|T201|COMP|1100-7|LNC|K little p super little a Ag|K little p super little a Ag
C0482283|T201|COMP|1101-5|LNC|K little p super little a Ag|K little p super little a Ag
C0482284|T201|COMP|1102-3|LNC|K little p super little a Ag|K little p super little a Ag
C0482285|T201|COMP|1103-1|LNC|K little p super little b Ab|K little p super little b Ab
C0482286|T201|COMP|1104-9|LNC|K little p super little b Ab|K little p super little b Ab
C0482287|T201|COMP|1105-6|LNC|K little p super little b Ab|K little p super little b Ab
C0482288|T201|COMP|1106-4|LNC|K little p super little b Ag|K little p super little b Ag
C0482289|T201|COMP|1107-2|LNC|K little p super little b Ag|K little p super little b Ag
C0482290|T201|COMP|1108-0|LNC|K little p super little b Ag|K little p super little b Ag
C0482291|T201|COMP|1109-8|LNC|L little b|L little b
C0482292|T201|COMP|1110-6|LNC|L little e super little a Ab|L little e super little a Ab
C0482293|T201|COMP|1111-4|LNC|L little e super little a Ab|L little e super little a Ab
C0482294|T201|COMP|1112-2|LNC|L little e super little a Ab|L little e super little a Ab
C0482295|T201|COMP|1113-0|LNC|L little e super little a Ag|L little e super little a Ag
C0482296|T201|COMP|1114-8|LNC|L little e super little a Ag|L little e super little a Ag
C0482297|T201|COMP|1115-5|LNC|L little e super little a Ag|L little e super little a Ag
C0482298|T201|COMP|1116-3|LNC|L little e super little b Ab|L little e super little b Ab
C0482299|T201|COMP|1117-1|LNC|L little e super little b Ab|L little e super little b Ab
C0482300|T201|COMP|1118-9|LNC|L little e super little b Ab|L little e super little b Ab
C0482301|T201|COMP|1119-7|LNC|L little e super little b Ag|L little e super little b Ag
C0482302|T201|COMP|1120-5|LNC|L little e super little b Ag|L little e super little b Ag
C0482303|T201|COMP|1121-3|LNC|L little e super little b Ag|L little e super little b Ag
C0482304|T201|COMP|1122-1|LNC|L little e super little x Ab|L little e super little x Ab
C0482305|T201|COMP|1123-9|LNC|L little e super little x Ab|L little e super little x Ab
C0482306|T201|COMP|1124-7|LNC|L little e super little x Ab|L little e super little x Ab
C0482307|T201|COMP|1125-4|LNC|L little e Ab|L little e Ab
C0482308|T201|COMP|1126-2|LNC|L little e Ab|L little e Ab
C0482309|T201|COMP|1129-6|LNC|L little e NOS Ab|L little e NOS Ab
C0482310|T201|COMP|1130-4|LNC|L little e NOS Ag|L little e NOS Ag
C0482311|T201|COMP|1131-2|LNC|L little e NOS Ag|L little e NOS Ag
C0482312|T201|COMP|1132-0|LNC|L little e NOS Ag|L little e NOS Ag
C0482313|T201|COMP|1133-8|LNC|L little u super little a Ab|L little u super little a Ab
C0482314|T201|COMP|1134-6|LNC|L little u super little a Ab|L little u super little a Ab
C0482315|T201|COMP|1135-3|LNC|L little u super little a Ab|L little u super little a Ab
C0482316|T201|COMP|1136-1|LNC|L little u super little a Ag|L little u super little a Ag
C0482317|T201|COMP|1137-9|LNC|L little u super little a Ag|L little u super little a Ag
C0482318|T201|COMP|1138-7|LNC|L little u super little a Ag|L little u super little a Ag
C0482319|T201|COMP|1139-5|LNC|L little u super little a super little b Ab|L little u super little a super little b Ab
C0482320|T201|COMP|1140-3|LNC|L little u super little a super little b Ab|L little u super little a super little b Ab
C0482321|T201|COMP|1141-1|LNC|L little u super little a super little b Ab|L little u super little a super little b Ab
C0482322|T201|COMP|1142-9|LNC|L little u super little b Ab|L little u super little b Ab
C0482323|T201|COMP|1143-7|LNC|L little u super little b Ab|L little u super little b Ab
C0482324|T201|COMP|1144-5|LNC|L little u super little b Ab|L little u super little b Ab
C0482325|T201|COMP|1145-2|LNC|L little u super little b Ag|L little u super little b Ag
C0482326|T201|COMP|1146-0|LNC|L little u super little b Ag|L little u super little b Ag
C0482327|T201|COMP|1147-8|LNC|L little u super little b Ag|L little u super little b Ag
C0482328|T201|COMP|1148-6|LNC|L little u NOS Ab|L little u NOS Ab
C0482329|T201|COMP|1149-4|LNC|L little u NOS Ab|L little u NOS Ab
C0482330|T201|COMP|1150-2|LNC|L little u NOS Ab|L little u NOS Ab
C0482331|T201|COMP|1151-0|LNC|L little u NOS Ag|L little u NOS Ag
C0482332|T201|COMP|1152-8|LNC|L little u NOS Ag|L little u NOS Ag
C0482333|T201|COMP|1153-6|LNC|L little u NOS Ag|L little u NOS Ag
C0482334|T201|COMP|1166-8|LNC|little f Ab|little f Ab
C0482335|T201|COMP|1167-6|LNC|little f Ab|little f Ab
C0482336|T201|COMP|1168-4|LNC|little f Ab|little f Ab
C0482337|T201|COMP|1169-2|LNC|little f Ag|little f Ag
C0482338|T201|COMP|1170-0|LNC|little f Ag|little f Ag
C0482339|T201|COMP|1171-8|LNC|little f Ag|little f Ag
C0482340|T201|COMP|1172-6|LNC|little i -1 Ab|little i -1 Ab
C0482341|T201|COMP|1173-4|LNC|little i -1 Ab|little i -1 Ab
C0482342|T201|COMP|1174-2|LNC|little i -1 Ab|little i -1 Ab
C0482343|T201|COMP|1175-9|LNC|little i -1 Ag|little i -1 Ag
C0482344|T201|COMP|1176-7|LNC|little i -1 Ag|little i -1 Ag
C0482345|T201|COMP|1177-5|LNC|little i -1 Ag|little i -1 Ag
C0482346|T201|COMP|1178-3|LNC|little i -2 Ab|little i -2 Ab
C0482347|T201|COMP|1179-1|LNC|little i -2 Ab|little i -2 Ab
C0482348|T201|COMP|1180-9|LNC|little i -2 Ab|little i -2 Ab
C0482349|T201|COMP|1181-7|LNC|little i -2 Ag|little i -2 Ag
C0482350|T201|COMP|1182-5|LNC|little i -2 Ag|little i -2 Ag
C0482351|T201|COMP|1183-3|LNC|little i -2 Ag|little i -2 Ag
C0482355|T201|COMP|1199-9|LNC|little p little k Ab|little p little k Ab
C0482356|T201|COMP|1200-5|LNC|little p little k Ab|little p little k Ab
C0482357|T201|COMP|1201-3|LNC|little p little k Ab|little p little k Ab
C0482358|T201|COMP|1202-1|LNC|little p little k Ag|little p little k Ag
C0482359|T201|COMP|1203-9|LNC|little p little k Ag|little p little k Ag
C0482360|T201|COMP|1204-7|LNC|little p little k Ag|little p little k Ag
C0482361|T201|COMP|1205-4|LNC|little p Ag|little p Ag
C0482362|T201|COMP|1206-2|LNC|little p Ag|little p Ag
C0482363|T201|COMP|1207-0|LNC|little p Ag|little p Ag
C0482364|T201|COMP|1214-6|LNC|LW Ab|LW Ab
C0482365|T201|COMP|1215-3|LNC|LW Ab|LW Ab
C0482366|T201|COMP|1216-1|LNC|LW Ab|LW Ab
C0482367|T201|COMP|1217-9|LNC|LW Ag|LW Ag
C0482368|T201|COMP|1218-7|LNC|LW Ag|LW Ag
C0482369|T201|COMP|1219-5|LNC|LW Ag|LW Ag
C0482370|T201|COMP|1220-3|LNC|M little g Ab|M little g Ab
C0482371|T201|COMP|1221-1|LNC|M little g Ab|M little g Ab
C0482372|T201|COMP|1222-9|LNC|M little g Ab|M little g Ab
C0482373|T201|COMP|1223-7|LNC|M little g Ag|M little g Ag
C0482374|T201|COMP|1224-5|LNC|M little g Ag|M little g Ag
C0482375|T201|COMP|1225-2|LNC|M little g Ag|M little g Ag
C0482376|T201|COMP|1235-1|LNC|M little i super little a Ab|M little i super little a Ab
C0482377|T201|COMP|1236-9|LNC|M little i super little a Ab|M little i super little a Ab
C0482378|T201|COMP|1237-7|LNC|M little i super little a Ab|M little i super little a Ab
C0482379|T201|COMP|1232-8|LNC|M little i super little a Ag|M little i super little a Ag
C0482380|T201|COMP|1233-6|LNC|M little i super little a Ag|M little i super little a Ag
C0482381|T201|COMP|1234-4|LNC|M little i super little a Ag|M little i super little a Ag
C0482382|T201|COMP|1226-0|LNC|M Ab|M Ab
C0482383|T201|COMP|1227-8|LNC|M Ab|M Ab
C0482384|T201|COMP|1228-6|LNC|M Ab|M Ab
C0482385|T201|COMP|1229-4|LNC|M Ag|M Ag
C0482386|T201|COMP|1230-2|LNC|M Ag|M Ag
C0482387|T201|COMP|1231-0|LNC|M Ag|M Ag
C0482388|T201|COMP|1244-3|LNC|M1 Ab|M1 Ab
C0482389|T201|COMP|1245-0|LNC|M1 Ab|M1 Ab
C0482390|T201|COMP|1246-8|LNC|M1 Ab|M1 Ab
C0482391|T201|COMP|1247-6|LNC|M1 Ag|M1 Ag
C0482392|T201|COMP|1248-4|LNC|M1 Ag|M1 Ag
C0482393|T201|COMP|1249-2|LNC|M1 Ag|M1 Ag
C0482394|T201|COMP|1256-7|LNC|N Ab|N Ab
C0482395|T201|COMP|1257-5|LNC|N Ab|N Ab
C0482396|T201|COMP|1258-3|LNC|N Ab|N Ab
C0482397|T201|COMP|1259-1|LNC|N Ag|N Ag
C0482398|T201|COMP|1260-9|LNC|N Ag|N Ag
C0482399|T201|COMP|1261-7|LNC|N Ag|N Ag
C0482400|T201|COMP|1268-2|LNC|NOS Ab|NOS Ab
C0482401|T201|COMP|1269-0|LNC|NOS Ab|NOS Ab
C0482402|T201|COMP|1270-8|LNC|Unidentified Ab|Unidentified Ab
C0482403|T201|COMP|1271-6|LNC|O NOS Ab|O NOS Ab
C0482404|T201|COMP|1272-4|LNC|O NOS Ab|O NOS Ab
C0482405|T201|COMP|1273-2|LNC|O NOS Ab|O NOS Ab
C0482406|T201|COMP|1274-0|LNC|O NOS Ag|O NOS Ag
C0482407|T201|COMP|1275-7|LNC|O NOS Ag|O NOS Ag
C0482408|T201|COMP|1276-5|LNC|O NOS Ag|O NOS Ag
C0482409|T201|COMP|1277-3|LNC|P Ab|P Ab
C0482410|T201|COMP|1278-1|LNC|P Ab|P Ab
C0482411|T201|COMP|1279-9|LNC|P Ab|P Ab
C0482412|T201|COMP|1286-4|LNC|P1 Ab|P1 Ab
C0482413|T201|COMP|1287-2|LNC|P1 Ab|P1 Ab
C0482414|T201|COMP|1288-0|LNC|P1 Ab|P1 Ab
C0482415|T201|COMP|1289-8|LNC|P1 Ag|P1 Ag
C0482416|T201|COMP|1290-6|LNC|P1 Ag|P1 Ag
C0482417|T201|COMP|1291-4|LNC|P1 Ag|P1 Ag
C0482418|T201|COMP|1292-2|LNC|P2 Ab|P2 Ab
C0482419|T201|COMP|1293-0|LNC|P2 Ab|P2 Ab
C0482420|T201|COMP|1294-8|LNC|P2 Ab|P2 Ab
C0482421|T201|COMP|1295-5|LNC|P2 Ag|P2 Ag
C0482422|T201|COMP|1296-3|LNC|P2 Ag|P2 Ag
C0482423|T201|COMP|1297-1|LNC|P2 Ag|P2 Ag
C0482424|T201|COMP|1300-3|LNC|PP1 Ab|PP1 Ab
C0482425|T201|COMP|1301-1|LNC|PP1 Ab|PP1 Ab
C0482426|T201|COMP|1302-9|LNC|PP1 Ab|PP1 Ab
C0482427|T201|COMP|1313-6|LNC|Rh immune globulin dosage.vials recommended|Rh immune globulin dosage.vials recommended
C0482428|T201|COMP|1314-4|LNC|Rh immune globulin screen|Rh immune globulin screen
C0482429|T201|COMP|1323-5|LNC|U Ab|U Ab
C0482430|T201|COMP|1324-3|LNC|U Ab|U Ab
C0482431|T201|COMP|1325-0|LNC|U Ab|U Ab
C0482432|T201|COMP|1326-8|LNC|U Ag|U Ag
C0482433|T201|COMP|1327-6|LNC|U Ag|U Ag
C0482434|T201|COMP|1328-4|LNC|U Ag|U Ag
C0482435|T201|COMP|1329-2|LNC|V Ab|V Ab
C0482436|T201|COMP|1330-0|LNC|V Ab|V Ab
C0482437|T201|COMP|1331-8|LNC|V Ab|V Ab
C0482438|T201|COMP|1332-6|LNC|V Ag|V Ag
C0482439|T201|COMP|1333-4|LNC|V Ag|V Ag
C0482440|T201|COMP|1334-2|LNC|V Ag|V Ag
C0482441|T201|COMP|1336-7|LNC|X little g super little a Ab|X little g super little a Ab
C0482442|T201|COMP|1337-5|LNC|X little g super little a Ab|X little g super little a Ab
C0482443|T201|COMP|1338-3|LNC|X little g super little a Ab|X little g super little a Ab
C0482444|T201|COMP|1339-1|LNC|X little g super little a Ag|X little g super little a Ag
C0482445|T201|COMP|1340-9|LNC|X little g super little a Ag|X little g super little a Ag
C0482446|T201|COMP|1341-7|LNC|X little g super little a Ag|X little g super little a Ag
C0482447|T201|COMP|1342-5|LNC|Y little t super little a Ab|Y little t super little a Ab
C0482448|T201|COMP|1343-3|LNC|Y little t super little a Ab|Y little t super little a Ab
C0482449|T201|COMP|1344-1|LNC|Y little t super little a Ab|Y little t super little a Ab
C0482450|T201|COMP|1345-8|LNC|Y little t super little a Ag|Y little t super little a Ag
C0482451|T201|COMP|1346-6|LNC|Y little t super little a Ag|Y little t super little a Ag
C0482452|T201|COMP|1347-4|LNC|Y little t super little a Ag|Y little t super little a Ag
C0482453|T201|COMP|1348-2|LNC|Y little t super little b Ab|Y little t super little b Ab
C0482454|T201|COMP|1349-0|LNC|Y little t super little b Ab|Y little t super little b Ab
C0482455|T201|COMP|1350-8|LNC|Y little t super little b Ab|Y little t super little b Ab
C0482456|T201|COMP|1351-6|LNC|Y little t super little b Ag|Y little t super little b Ag
C0482457|T201|COMP|1352-4|LNC|Y little t super little b Ag|Y little t super little b Ag
C0482458|T201|COMP|1353-2|LNC|Y little t super little b Ag|Y little t super little b Ag
C0482460|T201|COMP|1359-9|LNC|Corticotropin^1H post 1 ug/kg CRH IV|Corticotropin^1H post 1 ug/kg CRH IV
C0482461|T201|COMP|1361-5|LNC|Corticotropin^1M post 1 ug/kg CRH IV|Corticotropin^1M post 1 ug/kg CRH IV
C0482462|T201|COMP|1362-3|LNC|Corticotropin^30M post 1 ug/kg CRH IV|Corticotropin^30M post 1 ug/kg CRH IV
C0482463|T201|COMP|1364-9|LNC|Corticotropin^45M post 1 ug/kg CRH IV|Corticotropin^45M post 1 ug/kg CRH IV
C0482464|T201|COMP|1366-4|LNC|Corticotropin^5M post 1 ug/kg CRH IV|Corticotropin^5M post 1 ug/kg CRH IV
C0482465|T201|COMP|1367-2|LNC|Corticotropin^pre 1 ug/kg CRH IV|Corticotropin^pre 1 ug/kg CRH IV
C0482466|T201|COMP|1368-0|LNC|Corticotropin^pre dose insulin IV|Corticotropin^pre dose insulin IV
C0482467|T201|COMP|1370-6|LNC|Carotene^post 15000 U carotene QDx3 for 3D poly|Carotene^post 15000 U carotene QDx3 for 3D poly
C0482468|T201|COMP|1372-2|LNC|Calcitonin^90s post 0.5 ug/kg pentagastrin IV|Calcitonin^90s post 0.5 ug/kg pentagastrin IV
C0482469|T201|COMP|1376-3|LNC|Calcitonin^5M post 0.5 ug/kg pentagastrin IV|Calcitonin^5M post 0.5 ug/kg pentagastrin IV
C0482470|T201|COMP|1378-9|LNC|Calcitonin^pre 0.5 ug/kg pentagastrin IV|Calcitonin^pre 0.5 ug/kg pentagastrin IV
C0482471|T201|COMP|1379-7|LNC|Calcitonin^pre 2.4 mg/kg calcium short IV|Calcitonin^pre 2.4 mg/kg calcium short IV
C0482472|T201|COMP|1383-9|LNC|Calcium^pre 2.4 mg/kg calcium short IV|Calcium^pre 2.4 mg/kg calcium short IV
C0482481|T201|COMP|1394-6|LNC|Cortisol.free^pre 50 ug corticotropin IM 3 day|Cortisol.free^pre 50 ug corticotropin IM 3 day
C0482484|T201|COMP|1400-1|LNC|Cortisol^1H post 1 ug/kg CRH IV|Cortisol^1H post 1 ug/kg CRH IV
C0482485|T201|COMP|1401-9|LNC|Cortisol^1H post 250 ug corticotropin IM rapid|Cortisol^1H post 250 ug corticotropin IM rapid
C0482486|T201|COMP|1402-7|LNC|Cortisol^1H post 250 ug corticotropin IV rapid|Cortisol^1H post 250 ug corticotropin IV rapid
C0482487|T201|COMP|1403-5|LNC|Cortisol^1H post 250 ug corticotropin IM|Cortisol^1H post 250 ug corticotropin IM
C0482488|T201|COMP|1406-8|LNC|Cortisol^1M post 1 ug/kg CRH IV|Cortisol^1M post 1 ug/kg CRH IV
C0482490|T201|COMP|1409-2|LNC|Cortisol^24H post 500 ug corticotropin IM|Cortisol^24H post 500 ug corticotropin IM
C0482493|T201|COMP|1413-4|LNC|Cortisol^2D post 500 ug corticotropin IM|Cortisol^2D post 500 ug corticotropin IM
C0482494|T201|COMP|1415-9|LNC|Cortisol^30M post 1 ug/kg CRH IV|Cortisol^30M post 1 ug/kg CRH IV
C0482495|T201|COMP|1416-7|LNC|Cortisol^30M post 250 ug corticotropin IM rapid|Cortisol^30M post 250 ug corticotropin IM rapid
C0482496|T201|COMP|1417-5|LNC|Cortisol^30M post 250 ug corticotropin IV rapid|Cortisol^30M post 250 ug corticotropin IV rapid
C0482497|T201|COMP|1418-3|LNC|Cortisol^30M post 250 ug corticotropin IM|Cortisol^30M post 250 ug corticotropin IM
C0482499|T201|COMP|1422-5|LNC|Cortisol^3D post 500 ug corticotropin IM|Cortisol^3D post 500 ug corticotropin IM
C0482500|T201|COMP|1423-3|LNC|Cortisol^45M post 1 ug/kg CRH IV|Cortisol^45M post 1 ug/kg CRH IV
C0482505|T201|COMP|1431-6|LNC|Cortisol^5M post 1 ug/kg CRH IV|Cortisol^5M post 1 ug/kg CRH IV
C0482508|T201|COMP|1438-1|LNC|Cortisol^8H post 40 ug corticotropin IM BID 3 day|Cortisol^8H post 40 ug corticotropin IM BID 3 day
C0482509|T201|COMP|1443-1|LNC|Cortisol^pre 1 ug/kg CRH IV|Cortisol^pre 1 ug/kg CRH IV
C0482510|T201|COMP|1444-9|LNC|Cortisol^pre 12H CFst|Cortisol^pre 12H CFst
C0482511|T201|COMP|1445-6|LNC|Cortisol^pre 1 mg dexamethasone PO overnight|Cortisol^pre 1 mg dexamethasone PO overnight
C0482512|T201|COMP|1446-4|LNC|Cortisol^pre 3 g metyraPONE PO overnight|Cortisol^pre 3 g metyraPONE PO overnight
C0482513|T201|COMP|1447-2|LNC|Cortisol^pre 40 ug corticotropin IM 3 day|Cortisol^pre 40 ug corticotropin IM 3 day
C0482517|T201|COMP|1451-4|LNC|Cortisol^pre dose insulin IV|Cortisol^pre dose insulin IV
C0482522|T201|COMP|1457-1|LNC|Creatinine^pre 40 ug corticotropin IM 3 day|Creatinine^pre 40 ug corticotropin IM 3 day
C0482525|T201|COMP|1461-3|LNC|Epinephrine^1H post 300 ug cloNIDine PO|Epinephrine^1H post 300 ug cloNIDine PO
C0482526|T201|COMP|1462-1|LNC|Epinephrine^2H post 300 ug cloNIDine PO|Epinephrine^2H post 300 ug cloNIDine PO
C0482527|T201|COMP|1463-9|LNC|Epinephrine^3H post 300 ug cloNIDine PO|Epinephrine^3H post 300 ug cloNIDine PO
C0482528|T201|COMP|1464-7|LNC|Epinephrine^pre 300 ug cloNIDine PO|Epinephrine^pre 300 ug cloNIDine PO
C0482533|T201|COMP|1490-2|LNC|Gastrin^pre 0.2 U/kg secretin|Gastrin^pre 0.2 U/kg secretin
C0482534|T201|COMP|1496-9|LNC|Glucose^1.5H post 75 g glucose PO|Glucose^1.5H post 75 g glucose PO
C0482535|T201|COMP|1521-4|LNC|Glucose^2H post meal|Glucose^2H post meal
C0482536|T201|COMP|1524-8|LNC|Glucose^30M post 0.1 U/kg insulin|Glucose^30M post 0.1 U/kg insulin
C0482537|T201|COMP|1527-1|LNC|Glucose^30M post 75 g glucose PO|Glucose^30M post 75 g glucose PO
C0482538|T201|COMP|1548-7|LNC|Glucose^pre 0.5 g/kg glucose IV|Glucose^pre 0.5 g/kg glucose IV
C0482539|T201|COMP|1549-5|LNC|Glucose^pre 100 g glucose PO|Glucose^pre 100 g glucose PO
C0482540|T201|COMP|1550-3|LNC|Glucose^pre 12H CFst|Glucose^pre 12H CFst
C0482541|T201|COMP|1551-1|LNC|Glucose^pre 50 g lactose PO|Glucose^pre 50 g lactose PO
C0482542|T201|COMP|1552-9|LNC|Glucose^pre 75 g glucose PO|Glucose^pre 75 g glucose PO
C0482543|T201|COMP|1553-7|LNC|Glucose^pre dose insulin IV|Glucose^pre dose insulin IV
C0482544|T201|COMP|1558-6|LNC|Glucose^post CFst|Glucose^post CFst
C0482545|T201|COMP|2437-2|LNC|Hydrogen/Expired gas^post 50 g glucose PO|Hydrogen/Expired gas^post 50 g glucose PO
C0482546|T201|COMP|1559-4|LNC|Insulin^1.5H post dose TOLBUTamide IV|Insulin^1.5H post dose TOLBUTamide IV
C0482547|T201|COMP|1560-2|LNC|Insulin^1H post dose TOLBUTamide IV|Insulin^1H post dose TOLBUTamide IV
C0482548|T201|COMP|1562-8|LNC|Insulin^2.5H post dose TOLBUTamide IV|Insulin^2.5H post dose TOLBUTamide IV
C0482549|T201|COMP|1563-6|LNC|Insulin^2H post dose TOLBUTamide IV|Insulin^2H post dose TOLBUTamide IV
C0482550|T201|COMP|1565-1|LNC|Insulin^30M post dose TOLBUTamide IV|Insulin^30M post dose TOLBUTamide IV
C0482551|T201|COMP|1566-9|LNC|Insulin^3H post dose TOLBUTamide IV|Insulin^3H post dose TOLBUTamide IV
C0482552|T201|COMP|1571-9|LNC|Insulin^pre dose TOLBUTamide IV|Insulin^pre dose TOLBUTamide IV
C0482553|T201|COMP|1572-7|LNC|Insulin^pre 75 g glucose PO|Insulin^pre 75 g glucose PO
C0482561|T201|COMP|1585-9|LNC|Lactose^pre 12H CFst|Lactose^pre 12H CFst
C0482562|T201|COMP|1600-6|LNC|Lutropin^pre dose gonadotropin releasing hormone|Lutropin^pre dose gonadotropin releasing hormone
C0482563|T201|COMP|1603-0|LNC|Norepinephrine^1H post 300 ug clonidine PO|Norepinephrine^1H post 300 ug clonidine PO
C0482564|T201|COMP|1604-8|LNC|Norepinephrine^2H post 300 ug clonidine PO|Norepinephrine^2H post 300 ug clonidine PO
C0482565|T201|COMP|1605-5|LNC|Norepinephrine^3H post 300 ug clonidine PO|Norepinephrine^3H post 300 ug clonidine PO
C0482566|T201|COMP|1606-3|LNC|Norepinephrine^pre 300 ug clonidine PO|Norepinephrine^pre 300 ug clonidine PO
C0482567|T201|COMP|1609-7|LNC|Prolactin^1.5H post dose insulin IV|Prolactin^1.5H post dose insulin IV
C0482568|T201|COMP|1610-5|LNC|Prolactin^1H post dose L-Dopa PO|Prolactin^1H post dose L-Dopa PO
C0482569|T201|COMP|1611-3|LNC|Prolactin^1H post dose TRH IV|Prolactin^1H post dose TRH IV
C0482570|T201|COMP|1612-1|LNC|Prolactin^1H post dose insulin IV|Prolactin^1H post dose insulin IV
C0482571|T201|COMP|1613-9|LNC|Prolactin^2H post dose L-Dopa PO|Prolactin^2H post dose L-Dopa PO
C0482572|T201|COMP|1614-7|LNC|Prolactin^30M post dose TRH IV|Prolactin^30M post dose TRH IV
C0482573|T201|COMP|1615-4|LNC|Prolactin^30M post dose insulin IV|Prolactin^30M post dose insulin IV
C0482574|T201|COMP|1617-0|LNC|Prolactin^3H post dose L-Dopa PO|Prolactin^3H post dose L-Dopa PO
C0482575|T201|COMP|1618-8|LNC|Prolactin^45M post dose insulin IV|Prolactin^45M post dose insulin IV
C0482576|T201|COMP|1619-6|LNC|Prolactin^pre dose L-dopa PO|Prolactin^pre dose L-dopa PO
C0482577|T201|COMP|1620-4|LNC|Prolactin^pre dose TRH IV|Prolactin^pre dose TRH IV
C0482578|T201|COMP|1621-2|LNC|Prolactin^pre dose insulin IV|Prolactin^pre dose insulin IV
C0482579|T201|COMP|1623-8|LNC|Renin^pre 600 ug furosemide PO|Renin^pre 600 ug furosemide PO
C0482580|T201|COMP|1634-5|LNC|Somatotropin^52H post 250 ug L-Dopa TID 2day PO|Somatotropin^52H post 250 ug L-Dopa TID 2day PO
C0482581|T201|COMP|1635-2|LNC|Somatotropin^pre 1 g/kg glucose PO|Somatotropin^pre 1 g/kg glucose PO
C0482582|T201|COMP|1636-0|LNC|Somatotropin^pre 250 ug L-Dopa TID 2day PO|Somatotropin^pre 250 ug L-Dopa TID 2day PO
C0482583|T201|COMP|1637-8|LNC|Somatotropin^pre dose insulin IV|Somatotropin^pre dose insulin IV
C0482584|T201|COMP|1639-4|LNC|Testosterone^pre 5000 U HCG IM|Testosterone^pre 5000 U HCG IM
C0482585|T201|COMP|1640-2|LNC|Thyrotropin^30M post dose TRH IV|Thyrotropin^30M post dose TRH IV
C0482586|T201|COMP|1641-0|LNC|Thyrotropin^1H post dose TRH IV|Thyrotropin^1H post dose TRH IV
C0482587|T201|COMP|1643-6|LNC|Thyrotropin^pre dose TRH IV|Thyrotropin^pre dose TRH IV
C0482590|T201|COMP|1721-0|LNC|Adenosine triphosphate|Adenosine triphosphate
C0482591|T201|COMP|1734-3|LNC|Aldosterone renal clearance|Aldosterone renal clearance
C0482592|T201|COMP|1869-7|LNC|Apolipoprotein A-I|Apolipoprotein A-I
C0482593|T201|COMP|1966-1|LNC|Bile acid|Bile acid
C0482594|T201|COMP|2029-7|LNC|Carboxyhemoglobin|Carboxyhemoglobin
C0482595|T201|COMP|2610-4|LNC|Methane|Methane
C0482596|T201|COMP|2658-3|LNC|Nitrogen|Nitrogen
C0482597|T201|COMP|2723-5|LNC|Para aminohippurate renal clearance|Para aminohippurate renal clearance
C0482601|T201|COMP|2841-5|LNC|Prolactin|Prolactin
C0482602|T201|COMP|2842-3|LNC|Prolactin|Prolactin
C0482603|T201|COMP|3147-6|LNC|Oxygen|Oxygen
C0482604|T201|COMP|3174-0|LNC|Antithrombin|Antithrombin
C0482605|T201|COMP|3175-7|LNC|Antithrombin Ag|Antithrombin Ag
C0482606|T201|COMP|3176-5|LNC|Antithrombin|Antithrombin
C0482607|T201|COMP|3177-3|LNC|Antithrombin Ag|Antithrombin Ag
C0482608|T201|COMP|3184-9|LNC|Activated clotting time|Activated clotting time
C0482609|T201|COMP|3185-6|LNC|Coagulation factor IX inhibitor|Coagulation factor IX inhibitor
C0482610|T201|COMP|3186-4|LNC|Coagulation factor IX activated activity|Coagulation factor IX activated activity
C0482611|T201|COMP|3187-2|LNC|Coagulation factor IX activity actual/Normal|Coagulation factor IX activity actual/Normal
C0482612|T201|COMP|3188-0|LNC|Coagulation factor IX activity|Coagulation factor IX activity
C0482613|T201|COMP|3189-8|LNC|Coagulation factor IX Ag|Coagulation factor IX Ag
C0482614|T201|COMP|3190-6|LNC|Coagulation factor IX Ag actual/Normal|Coagulation factor IX Ag actual/Normal
C0482615|T201|COMP|3191-4|LNC|Coagulation factor V inhibitor|Coagulation factor V inhibitor
C0482616|T201|COMP|3192-2|LNC|Coagulation factor V activated activity|Coagulation factor V activated activity
C0482617|T201|COMP|3193-0|LNC|Coagulation factor V activity actual/Normal|Coagulation factor V activity actual/Normal
C0482618|T201|COMP|3194-8|LNC|Coagulation factor V Ag|Coagulation factor V Ag
C0482619|T201|COMP|3195-5|LNC|Coagulation factor V Ag actual/Normal|Coagulation factor V Ag actual/Normal
C0482620|T201|COMP|3196-3|LNC|Coagulation factor VII inhibitor|Coagulation factor VII inhibitor
C0482621|T201|COMP|3197-1|LNC|Coagulation factor VII activated activity|Coagulation factor VII activated activity
C0482622|T201|COMP|3198-9|LNC|Coagulation factor VII activity actual/Normal|Coagulation factor VII activity actual/Normal
C0482623|T201|COMP|3199-7|LNC|Coagulation factor VII activity|Coagulation factor VII activity
C0482624|T201|COMP|3200-3|LNC|Coagulation factor VII activity actual/Normal|Coagulation factor VII activity actual/Normal
C0482625|T201|COMP|3201-1|LNC|Coagulation factor VII Ag|Coagulation factor VII Ag
C0482626|T201|COMP|3202-9|LNC|Coagulation factor VII+Acarboxy Ag|Coagulation factor VII+Acarboxy Ag
C0482628|T201|COMP|3204-5|LNC|Coagulation factor VIII inhibitor|Coagulation factor VIII inhibitor
C0482629|T201|COMP|3205-2|LNC|Coagulation factor VIII Ab|Coagulation factor VIII Ab
C0482630|T201|COMP|3206-0|LNC|Coagulation factor VIII inhibitor|Coagulation factor VIII inhibitor
C0482631|T201|COMP|3207-8|LNC|Coagulation factor VIII inhibitor|Coagulation factor VIII inhibitor
C0482632|T201|COMP|3208-6|LNC|Coagulation factor VIII activated activity|Coagulation factor VIII activated activity
C0482633|T201|COMP|3209-4|LNC|Coagulation factor VIII activity actual/Normal|Coagulation factor VIII activity actual/Normal
C0482634|T201|COMP|3210-2|LNC|Coagulation factor VIII activity|Coagulation factor VIII activity
C0482635|T201|COMP|3211-0|LNC|Coagulation factor VIII activity actual/Normal|Coagulation factor VIII activity actual/Normal
C0482637|T201|COMP|3214-4|LNC|Coagulation factor VIII Ag|Coagulation factor VIII Ag
C0482638|T201|COMP|3215-1|LNC|Coagulation factor VIII Ag|Coagulation factor VIII Ag
C0482639|T201|COMP|3216-9|LNC|Coagulation factor X inhibitor|Coagulation factor X inhibitor
C0482640|T201|COMP|3217-7|LNC|Coagulation factor X activated activity|Coagulation factor X activated activity
C0482641|T201|COMP|3218-5|LNC|Coagulation factor X activity actual/Normal|Coagulation factor X activity actual/Normal
C0482642|T201|COMP|3219-3|LNC|Coagulation factor X activity|Coagulation factor X activity
C0482643|T201|COMP|3220-1|LNC|Coagulation factor X Ag|Coagulation factor X Ag
C0482644|T201|COMP|3221-9|LNC|Coagulation factor X Ag actual/Normal|Coagulation factor X Ag actual/Normal
C0482645|T201|COMP|3222-7|LNC|Coagulation factor X+Acarboxy Ag|Coagulation factor X+Acarboxy Ag
C0482646|T201|COMP|3223-5|LNC|Coagulation factor X+Acarboxy Ag actual/Normal|Coagulation factor X+Acarboxy Ag actual/Normal
C0482647|T201|COMP|3224-3|LNC|Coagulation factor XI inhibitor|Coagulation factor XI inhibitor
C0482648|T201|COMP|3225-0|LNC|Coagulation factor XI activated activity|Coagulation factor XI activated activity
C0482649|T201|COMP|3226-8|LNC|Coagulation factor XI activity actual/Normal|Coagulation factor XI activity actual/Normal
C0482650|T201|COMP|3227-6|LNC|Coagulation factor XI activity|Coagulation factor XI activity
C0482651|T201|COMP|3228-4|LNC|Coagulation factor XI Ag|Coagulation factor XI Ag
C0482652|T201|COMP|3229-2|LNC|Coagulation factor XI Ag actual/Normal|Coagulation factor XI Ag actual/Normal
C0482653|T201|COMP|3230-0|LNC|Coagulation factor XII inhibitor|Coagulation factor XII inhibitor
C0482654|T201|COMP|3231-8|LNC|Coagulation factor XII activated activity|Coagulation factor XII activated activity
C0482655|T201|COMP|3232-6|LNC|Coagulation factor XII activity actual/Normal|Coagulation factor XII activity actual/Normal
C0482656|T201|COMP|3233-4|LNC|Coagulation factor XII activity|Coagulation factor XII activity
C0482657|T201|COMP|3234-2|LNC|Coagulation factor XII Ag|Coagulation factor XII Ag
C0482658|T201|COMP|3235-9|LNC|Coagulation factor XII Ag actual/Normal|Coagulation factor XII Ag actual/Normal
C0482659|T201|COMP|3236-7|LNC|Coagulation factor XIII inhibitor|Coagulation factor XIII inhibitor
C0482660|T201|COMP|3237-5|LNC|Coagulation factor XIII activated activity|Coagulation factor XIII activated activity
C0482661|T201|COMP|3238-3|LNC|Coagulation factor XIII Ag|Coagulation factor XIII Ag
C0482662|T201|COMP|3239-1|LNC|Coagulation factor XIII Ag actual/Normal|Coagulation factor XIII Ag actual/Normal
C0482663|T201|COMP|3240-9|LNC|Coagulation factor XIII coagulum dissolution|Coagulation factor XIII coagulum dissolution
C0482665|T201|COMP|5942-8|LNC|Coagulation reptilase induced|Coagulation reptilase induced
C0482666|T201|COMP|5943-6|LNC|Coagulation reptilase induced|Coagulation reptilase induced
C0482667|T201|COMP|5903-0|LNC|Coagulation Russell viper venom induced|Coagulation Russell viper venom induced
C0482668|T201|COMP|5904-8|LNC|Coagulation Russell viper venom induced|Coagulation Russell viper venom induced
C0482669|T201|COMP|5944-4|LNC|Coagulation Russell viper venom induced|Coagulation Russell viper venom induced
C0482670|T201|COMP|5945-1|LNC|Coagulation Russell viper venom induced|Coagulation Russell viper venom induced
C0482679|T201|COMP|5899-0|LNC|Coagulation surface induced normal/Actual|Coagulation surface induced normal/Actual
C0482680|T201|COMP|5955-0|LNC|Coagulation thrombin induced|Coagulation thrombin induced
C0482681|T201|COMP|5954-3|LNC|Coagulation thrombin induced|Coagulation thrombin induced
C0482682|T201|COMP|5894-1|LNC|Coagulation tissue factor induced actual/Normal|Coagulation tissue factor induced actual/Normal
C0482691|T201|COMP|6301-6|LNC|Coagulation tissue factor induced.INR|Coagulation tissue factor induced.INR
C0482692|T201|COMP|6302-4|LNC|Coagulation tissue factor induced.normal/Actual|Coagulation tissue factor induced.normal/Actual
C0482693|T201|COMP|5901-4|LNC|Coagulation tissue factor induced|Coagulation tissue factor induced
C0482694|T201|COMP|5902-2|LNC|Coagulation tissue factor induced|Coagulation tissue factor induced
C0482695|T201|COMP|3242-5|LNC|Coagulation calcium ion induced|Coagulation calcium ion induced
C0482696|T201|COMP|3243-3|LNC|Coagulation thrombin induced|Coagulation thrombin induced
C0482697|T201|COMP|3244-1|LNC|Coagulum lysis|Coagulum lysis
C0482698|T201|COMP|3246-6|LNC|Fibrin D-dimer|Fibrin D-dimer
C0482699|T201|COMP|3247-4|LNC|Fibrin D-dimer|Fibrin D-dimer
C0482700|T201|COMP|3248-2|LNC|Fibrin fragments Ag|Fibrin fragments Ag
C0482701|T201|COMP|3249-0|LNC|Fibrin fragments|Fibrin fragments
C0482702|T201|COMP|3250-8|LNC|Fibrin monomer|Fibrin monomer
C0482703|T201|COMP|3251-6|LNC|Fibrin+Fibrinogen fragments|Fibrin+Fibrinogen fragments
C0482704|T201|COMP|3253-2|LNC|Fibrin.soluble|Fibrin.soluble
C0482705|T201|COMP|3255-7|LNC|Fibrinogen|Fibrinogen
C0482707|T201|COMP|3257-3|LNC|Fibrinogen|Fibrinogen
C0482708|T201|COMP|3256-5|LNC|Fibrinogen Ag|Fibrinogen Ag
C0482709|T201|COMP|3259-9|LNC|Fibrinogen fragments Ag|Fibrinogen fragments Ag
C0482710|T201|COMP|3260-7|LNC|Fibrinopeptide B beta (1-14) Ag|Fibrinopeptide B beta (1-14) Ag
C0482711|T201|COMP|3261-5|LNC|Fibrinopeptide B beta (1-42) Ag|Fibrinopeptide B beta (1-42) Ag
C0482712|T201|COMP|3262-3|LNC|Fibrinopeptide B beta (15-42) Ag|Fibrinopeptide B beta (15-42) Ag
C0482713|T201|COMP|3263-1|LNC|Fibrinopeptide B beta (43-47) Ag|Fibrinopeptide B beta (43-47) Ag
C0482714|T201|COMP|3264-9|LNC|Fibrinopeptide A Ag|Fibrinopeptide A Ag
C0482715|T201|COMP|3265-6|LNC|Fibrinopeptide B Ag|Fibrinopeptide B Ag
C0482716|T201|COMP|3266-4|LNC|Heparin Ab|Heparin Ab
C0482717|T201|COMP|3268-0|LNC|Heparin cofactor II Ag|Heparin cofactor II Ag
C0482718|T201|COMP|3269-8|LNC|Heparin neutralization|Heparin neutralization
C0482719|T201|COMP|3270-6|LNC|Heparin.low molecular weight|Heparin.low molecular weight
C0482720|T201|COMP|3271-4|LNC|Heparin.low molecular weight|Heparin.low molecular weight
C0482721|T201|COMP|3273-0|LNC|Heparin.unfractionated|Heparin.unfractionated
C0482722|T201|COMP|3274-8|LNC|Heparin.unfractionated|Heparin.unfractionated
C0482723|T201|COMP|3276-3|LNC|Kininogen.high molecular weight|Kininogen.high molecular weight
C0482724|T201|COMP|3277-1|LNC|Kininogen.high molecular weight|Kininogen.high molecular weight
C0482725|T201|COMP|3278-9|LNC|Kininogen.high molecular weight actual/Normal|Kininogen.high molecular weight actual/Normal
C0482726|T201|COMP|3279-7|LNC|Kininogen.low molecular weight|Kininogen.low molecular weight
C0482727|T201|COMP|3281-3|LNC|Lupus anticoagulant|Lupus anticoagulant
C0482730|T201|COMP|3284-7|LNC|Lupus anticoagulant neutralization.platelet|Lupus anticoagulant neutralization.platelet
C0482731|T201|COMP|5965-9|LNC|Plasmin inhibitor|Plasmin inhibitor
C0482732|T201|COMP|5967-5|LNC|Plasmin inhibitor Ag|Plasmin inhibitor Ag
C0482733|T201|COMP|5966-7|LNC|Plasmin inhibitor Ag|Plasmin inhibitor Ag
C0482734|T201|COMP|5969-1|LNC|Plasmin-plasmin inhibitor complex|Plasmin-plasmin inhibitor complex
C0482735|T201|COMP|5970-9|LNC|Plasminogen|Plasminogen
C0482738|T201|COMP|5974-1|LNC|Plasminogen activator inhibitor 1|Plasminogen activator inhibitor 1
C0482739|T201|COMP|5975-8|LNC|Plasminogen activator inhibitor 1 Ag|Plasminogen activator inhibitor 1 Ag
C0482740|T201|COMP|5978-2|LNC|Plasminogen activator inhibitor 2|Plasminogen activator inhibitor 2
C0482741|T201|COMP|5979-0|LNC|Plasminogen activator inhibitor 2 Ag|Plasminogen activator inhibitor 2 Ag
C0482742|T201|COMP|5977-4|LNC|Plasminogen activator inhibitor 2 Ag|Plasminogen activator inhibitor 2 Ag
C0482743|T201|COMP|5980-8|LNC|Plasminogen activator inhibitor Ag|Plasminogen activator inhibitor Ag
C0482747|T201|COMP|5985-7|LNC|Plasminogen activator urokinase type|Plasminogen activator urokinase type
C0482748|T201|COMP|5986-5|LNC|Plasminogen activator tissue type|Plasminogen activator tissue type
C0482749|T201|COMP|5987-3|LNC|Plasminogen activator tissue type|Plasminogen activator tissue type
C0482753|T201|COMP|5991-5|LNC|Plasminogen Ag|Plasminogen Ag
C0482754|T201|COMP|6001-2|LNC|Platelet factor 3|Platelet factor 3
C0482755|T201|COMP|6002-0|LNC|Platelet factor 4|Platelet factor 4
C0482756|T201|COMP|6003-8|LNC|Platelet factor 4 Ag|Platelet factor 4 Ag
C0482757|T201|COMP|6005-3|LNC|Prekallikrein|Prekallikrein
C0482758|T201|COMP|6004-6|LNC|Prekallikrein|Prekallikrein
C0482759|T201|COMP|6007-9|LNC|Protein C|Protein C
C0482760|T201|COMP|6006-1|LNC|Protein C|Protein C
C0482761|T201|COMP|6009-5|LNC|Protein C Ag|Protein C Ag
C0482762|T201|COMP|6008-7|LNC|Protein C+Acarboxy Ag|Protein C+Acarboxy Ag
C0482763|T201|COMP|6011-1|LNC|Protein C cofactor|Protein C cofactor
C0482764|T201|COMP|6010-3|LNC|Protein C inhibitor|Protein C inhibitor
C0482765|T201|COMP|5891-7|LNC|Protein S+Acarboxy Ag|Protein S+Acarboxy Ag
C0482766|T201|COMP|5890-9|LNC|Protein S+Acarboxy.free Ag|Protein S+Acarboxy.free Ag
C0482767|T201|COMP|5889-1|LNC|Protein S.free|Protein S.free
C0482768|T201|COMP|4677-1|LNC|Protein S.free Ag|Protein S.free Ag
C0482769|T201|COMP|5892-5|LNC|Protein S|Protein S
C0482770|T201|COMP|5893-3|LNC|Protein S|Protein S
C0482771|T201|COMP|3288-8|LNC|Prothrombin Ag|Prothrombin Ag
C0482772|T201|COMP|3289-6|LNC|Prothrombin.activity actual/Normal|Prothrombin.activity actual/Normal
C0482773|T201|COMP|6012-9|LNC|von Willebrand factor Ag|von Willebrand factor Ag
C0482774|T201|COMP|6013-7|LNC|von Willebrand factor multimers|von Willebrand factor multimers
C0482776|T201|COMP|3312-6|LNC|ALPRAZolam|ALPRAZolam
C0482777|T201|COMP|3327-4|LNC|Aminopyrine|Aminopyrine
C0482778|T201|COMP|3760-6|LNC|Mesoridazine|Mesoridazine
C0482780|T201|COMP|4532-8|LNC|Complement total hemolytic CH50|Complement total hemolytic CH50
C0482781|T201|COMP|4635-9|LNC|Hemoglobin.free|Hemoglobin.free
C0482782|T201|COMP|4662-3|LNC|Lymphocytes+Monocytes/100 leukocytes|Lymphocytes+Monocytes/100 leukocytes
C0482783|T201|COMP|4695-3|LNC|HLA-A19|HLA-A19
C0482784|T201|COMP|4696-1|LNC|HLA-A19|HLA-A19
C0482785|T201|COMP|4697-9|LNC|HLA-A33(19)|HLA-A33(19)
C0482786|T201|COMP|4698-7|LNC|HLA-A33(19)|HLA-A33(19)
C0482787|T201|COMP|4699-5|LNC|HLA-A34(10)|HLA-A34(10)
C0482788|T201|COMP|4700-1|LNC|HLA-A34(10)|HLA-A34(10)
C0482789|T201|COMP|4701-9|LNC|HLA-A36|HLA-A36
C0482790|T201|COMP|4702-7|LNC|HLA-A36|HLA-A36
C0482791|T201|COMP|4703-5|LNC|HLA-A43|HLA-A43
C0482792|T201|COMP|4704-3|LNC|HLA-A43|HLA-A43
C0482793|T201|COMP|4705-0|LNC|HLA-A66(10)|HLA-A66(10)
C0482794|T201|COMP|4706-8|LNC|HLA-A66(10)|HLA-A66(10)
C0482795|T201|COMP|4707-6|LNC|HLA-A68(28)|HLA-A68(28)
C0482796|T201|COMP|4708-4|LNC|HLA-A68(28)|HLA-A68(28)
C0482797|T201|COMP|4709-2|LNC|HLA-A69(28)|HLA-A69(28)
C0482798|T201|COMP|4710-0|LNC|HLA-A69(28)|HLA-A69(28)
C0482799|T201|COMP|4711-8|LNC|HLA-A74(19)|HLA-A74(19)
C0482800|T201|COMP|4712-6|LNC|HLA-A74(19)|HLA-A74(19)
C0482801|T201|COMP|4713-4|LNC|HLA-A10|HLA-A10
C0482802|T201|COMP|4714-2|LNC|HLA-A10|HLA-A10
C0482803|T201|COMP|4715-9|LNC|HLA-A11|HLA-A11
C0482804|T201|COMP|4716-7|LNC|HLA-A11|HLA-A11
C0482805|T201|COMP|4717-5|LNC|HLA-A1|HLA-A1
C0482806|T201|COMP|4718-3|LNC|HLA-A1|HLA-A1
C0482807|T201|COMP|4719-1|LNC|HLA-A23(9)|HLA-A23(9)
C0482808|T201|COMP|4720-9|LNC|HLA-A23(9)|HLA-A23(9)
C0482809|T201|COMP|4721-7|LNC|HLA-A24(9)|HLA-A24(9)
C0482810|T201|COMP|4722-5|LNC|HLA-A25(10)|HLA-A25(10)
C0482811|T201|COMP|4723-3|LNC|HLA-A25(10)|HLA-A25(10)
C0482812|T201|COMP|4724-1|LNC|HLA-A26(10)|HLA-A26(10)
C0482813|T201|COMP|4725-8|LNC|HLA-A26(10)|HLA-A26(10)
C0482814|T201|COMP|4726-6|LNC|HLA-A28|HLA-A28
C0482815|T201|COMP|4727-4|LNC|HLA-A28|HLA-A28
C0482816|T201|COMP|4728-2|LNC|HLA-A29(19)|HLA-A29(19)
C0482817|T201|COMP|4729-0|LNC|HLA-A29(19)|HLA-A29(19)
C0482818|T201|COMP|4730-8|LNC|HLA-A2|HLA-A2
C0482819|T201|COMP|4731-6|LNC|HLA-A2|HLA-A2
C0482820|T201|COMP|4732-4|LNC|HLA-A30(19)|HLA-A30(19)
C0482821|T201|COMP|4733-2|LNC|HLA-A30(19)|HLA-A30(19)
C0482822|T201|COMP|4734-0|LNC|HLA-A31(19)|HLA-A31(19)
C0482823|T201|COMP|4735-7|LNC|HLA-A31(19)|HLA-A31(19)
C0482824|T201|COMP|4736-5|LNC|HLA-A32(19)|HLA-A32(19)
C0482825|T201|COMP|4737-3|LNC|HLA-A32(19)|HLA-A32(19)
C0482826|T201|COMP|4738-1|LNC|HLA-A3|HLA-A3
C0482827|T201|COMP|4739-9|LNC|HLA-A3|HLA-A3
C0482828|T201|COMP|4740-7|LNC|HLA-A9|HLA-A9
C0482829|T201|COMP|4741-5|LNC|HLA-A9|HLA-A9
C0482830|T201|COMP|4742-3|LNC|HLA-B22|HLA-B22
C0482831|T201|COMP|4743-1|LNC|HLA-B22|HLA-B22
C0482832|T201|COMP|4744-9|LNC|HLA-B41|HLA-B41
C0482833|T201|COMP|4745-6|LNC|HLA-B41|HLA-B41
C0482834|T201|COMP|4746-4|LNC|HLA-B42|HLA-B42
C0482835|T201|COMP|4747-2|LNC|HLA-B42|HLA-B42
C0482836|T201|COMP|4748-0|LNC|HLA-B46|HLA-B46
C0482837|T201|COMP|4749-8|LNC|HLA-B46|HLA-B46
C0482838|T201|COMP|4750-6|LNC|HLA-B47|HLA-B47
C0482839|T201|COMP|4751-4|LNC|HLA-B47|HLA-B47
C0482840|T201|COMP|4752-2|LNC|HLA-B48|HLA-B48
C0482841|T201|COMP|4753-0|LNC|HLA-B48|HLA-B48
C0482842|T201|COMP|4754-8|LNC|HLA-B w4|HLA-B w4
C0482843|T201|COMP|4755-5|LNC|HLA-B w4|HLA-B w4
C0482844|T201|COMP|4756-3|LNC|HLA-B50(21)|HLA-B50(21)
C0482845|T201|COMP|4757-1|LNC|HLA-B50(21)|HLA-B50(21)
C0482846|T201|COMP|4758-9|LNC|HLA-B52(5)|HLA-B52(5)
C0482847|T201|COMP|4759-7|LNC|HLA-B52(5)|HLA-B52(5)
C0482848|T201|COMP|4760-5|LNC|HLA-B53|HLA-B53
C0482849|T201|COMP|4761-3|LNC|HLA-B53|HLA-B53
C0482850|T201|COMP|4762-1|LNC|HLA-B54(22)|HLA-B54(22)
C0482851|T201|COMP|4763-9|LNC|HLA-B54(22)|HLA-B54(22)
C0482852|T201|COMP|4764-7|LNC|HLA-B55(22)|HLA-B55(22)
C0482853|T201|COMP|4765-4|LNC|HLA-B55(22)|HLA-B55(22)
C0482854|T201|COMP|4766-2|LNC|HLA-B56(22)|HLA-B56(22)
C0482855|T201|COMP|4767-0|LNC|HLA-B56(22)|HLA-B56(22)
C0482856|T201|COMP|4768-8|LNC|HLA-B57(17)|HLA-B57(17)
C0482857|T201|COMP|4769-6|LNC|HLA-B57(17)|HLA-B57(17)
C0482858|T201|COMP|4770-4|LNC|HLA-B58(17)|HLA-B58(17)
C0482859|T201|COMP|4771-2|LNC|HLA-B58(17)|HLA-B58(17)
C0482860|T201|COMP|4772-0|LNC|HLA-B59|HLA-B59
C0482861|T201|COMP|4773-8|LNC|HLA-B59|HLA-B59
C0482862|T201|COMP|4774-6|LNC|HLA-B60(40)|HLA-B60(40)
C0482863|T201|COMP|4775-3|LNC|HLA-B60(40)|HLA-B60(40)
C0482864|T201|COMP|4776-1|LNC|HLA-B61(40)|HLA-B61(40)
C0482865|T201|COMP|4777-9|LNC|HLA-B61(40)|HLA-B61(40)
C0482866|T201|COMP|4778-7|LNC|HLA-B62(15)|HLA-B62(15)
C0482867|T201|COMP|4779-5|LNC|HLA-B62(15)|HLA-B62(15)
C0482868|T201|COMP|4780-3|LNC|HLA-B63(15)|HLA-B63(15)
C0482869|T201|COMP|4781-1|LNC|HLA-B63(15)|HLA-B63(15)
C0482870|T201|COMP|4782-9|LNC|HLA-B64(14)|HLA-B64(14)
C0482871|T201|COMP|4783-7|LNC|HLA-B64(14)|HLA-B64(14)
C0482872|T201|COMP|4784-5|LNC|HLA-B65(14)|HLA-B65(14)
C0482873|T201|COMP|4785-2|LNC|HLA-B65(14)|HLA-B65(14)
C0482874|T201|COMP|4786-0|LNC|HLA-B67|HLA-B67
C0482875|T201|COMP|4787-8|LNC|HLA-B67|HLA-B67
C0482876|T201|COMP|4788-6|LNC|HLA-B w6|HLA-B w6
C0482877|T201|COMP|4789-4|LNC|HLA-B w6|HLA-B w6
C0482878|T201|COMP|4790-2|LNC|HLA-B70|HLA-B70
C0482879|T201|COMP|4791-0|LNC|HLA-B70|HLA-B70
C0482880|T201|COMP|4792-8|LNC|HLA-B71(70)|HLA-B71(70)
C0482881|T201|COMP|4793-6|LNC|HLA-B71(70)|HLA-B71(70)
C0482882|T201|COMP|4794-4|LNC|HLA-B72(70)|HLA-B72(70)
C0482883|T201|COMP|4795-1|LNC|HLA-B72(70)|HLA-B72(70)
C0482884|T201|COMP|4796-9|LNC|HLA-B73|HLA-B73
C0482885|T201|COMP|4797-7|LNC|HLA-B73|HLA-B73
C0482886|T201|COMP|4798-5|LNC|HLA-B75(15)|HLA-B75(15)
C0482887|T201|COMP|4799-3|LNC|HLA-B75(15)|HLA-B75(15)
C0482888|T201|COMP|4800-9|LNC|HLA-B76(15)|HLA-B76(15)
C0482889|T201|COMP|4801-7|LNC|HLA-B76(15)|HLA-B76(15)
C0482890|T201|COMP|4802-5|LNC|HLA-B77(15)|HLA-B77(15)
C0482891|T201|COMP|4803-3|LNC|HLA-B77(15)|HLA-B77(15)
C0482892|T201|COMP|4804-1|LNC|HLA-B12|HLA-B12
C0482893|T201|COMP|4805-8|LNC|HLA-B12|HLA-B12
C0482894|T201|COMP|4806-6|LNC|HLA-B13|HLA-B13
C0482895|T201|COMP|4807-4|LNC|HLA-B13|HLA-B13
C0482896|T201|COMP|4808-2|LNC|HLA-B14|HLA-B14
C0482897|T201|COMP|4809-0|LNC|HLA-B14|HLA-B14
C0482898|T201|COMP|4810-8|LNC|HLA-B15|HLA-B15
C0482899|T201|COMP|4811-6|LNC|HLA-B15|HLA-B15
C0482900|T201|COMP|4812-4|LNC|HLA-B16|HLA-B16
C0482901|T201|COMP|4813-2|LNC|HLA-B16|HLA-B16
C0482902|T201|COMP|4814-0|LNC|HLA-B17|HLA-B17
C0482903|T201|COMP|4815-7|LNC|HLA-B17|HLA-B17
C0482904|T201|COMP|4816-5|LNC|HLA-B18|HLA-B18
C0482905|T201|COMP|4817-3|LNC|HLA-B18|HLA-B18
C0482906|T201|COMP|4818-1|LNC|HLA-B21|HLA-B21
C0482907|T201|COMP|4819-9|LNC|HLA-B21|HLA-B21
C0482908|T201|COMP|4820-7|LNC|HLA-B27|HLA-B27
C0482909|T201|COMP|4821-5|LNC|HLA-B27|HLA-B27
C0482910|T201|COMP|4822-3|LNC|HLA-B35|HLA-B35
C0482911|T201|COMP|4823-1|LNC|HLA-B35|HLA-B35
C0482912|T201|COMP|4824-9|LNC|HLA-B37|HLA-B37
C0482913|T201|COMP|4825-6|LNC|HLA-B37|HLA-B37
C0482914|T201|COMP|4826-4|LNC|HLA-B38(16)|HLA-B38(16)
C0482915|T201|COMP|4827-2|LNC|HLA-B38(16)|HLA-B38(16)
C0482916|T201|COMP|4828-0|LNC|HLA-B39(16)|HLA-B39(16)
C0482917|T201|COMP|4829-8|LNC|HLA-B39(16)|HLA-B39(16)
C0482918|T201|COMP|4830-6|LNC|HLA-B40|HLA-B40
C0482919|T201|COMP|4831-4|LNC|HLA-B40|HLA-B40
C0482920|T201|COMP|4832-2|LNC|HLA-B44(12)|HLA-B44(12)
C0482921|T201|COMP|4833-0|LNC|HLA-B44(12)|HLA-B44(12)
C0482922|T201|COMP|4834-8|LNC|HLA-B45(12)|HLA-B45(12)
C0482923|T201|COMP|4835-5|LNC|HLA-B45(12)|HLA-B45(12)
C0482924|T201|COMP|4836-3|LNC|HLA-B49(21)|HLA-B49(21)
C0482925|T201|COMP|4837-1|LNC|HLA-B49(21)|HLA-B49(21)
C0482926|T201|COMP|4838-9|LNC|HLA-B51(5)|HLA-B51(5)
C0482927|T201|COMP|4839-7|LNC|HLA-B51(5)|HLA-B51(5)
C0482928|T201|COMP|4840-5|LNC|HLA-B5|HLA-B5
C0482929|T201|COMP|4841-3|LNC|HLA-B5|HLA-B5
C0482930|T201|COMP|4842-1|LNC|HLA-B7|HLA-B7
C0482931|T201|COMP|4843-9|LNC|HLA-B7|HLA-B7
C0482932|T201|COMP|4844-7|LNC|HLA-B8|HLA-B8
C0482933|T201|COMP|4845-4|LNC|HLA-B8|HLA-B8
C0482934|T201|COMP|4846-2|LNC|HLA-Cw10(w3)|HLA-Cw10(w3)
C0482935|T201|COMP|4847-0|LNC|HLA-Cw10(w3)|HLA-Cw10(w3)
C0482936|T201|COMP|4848-8|LNC|HLA-Cw11|HLA-Cw11
C0482937|T201|COMP|4849-6|LNC|HLA-Cw11|HLA-Cw11
C0482938|T201|COMP|4850-4|LNC|HLA-Cw1|HLA-Cw1
C0482939|T201|COMP|4851-2|LNC|HLA-Cw1|HLA-Cw1
C0482940|T201|COMP|4852-0|LNC|HLA-Cw2|HLA-Cw2
C0482941|T201|COMP|4853-8|LNC|HLA-Cw2|HLA-Cw2
C0482942|T201|COMP|4854-6|LNC|HLA-Cw3|HLA-Cw3
C0482943|T201|COMP|4855-3|LNC|HLA-Cw3|HLA-Cw3
C0482944|T201|COMP|4856-1|LNC|HLA-Cw4|HLA-Cw4
C0482945|T201|COMP|4857-9|LNC|HLA-Cw4|HLA-Cw4
C0482946|T201|COMP|4858-7|LNC|HLA-Cw5|HLA-Cw5
C0482947|T201|COMP|4859-5|LNC|HLA-Cw5|HLA-Cw5
C0482948|T201|COMP|4860-3|LNC|HLA-Cw6|HLA-Cw6
C0482949|T201|COMP|4861-1|LNC|HLA-Cw6|HLA-Cw6
C0482950|T201|COMP|4862-9|LNC|HLA-Cw7|HLA-Cw7
C0482951|T201|COMP|4863-7|LNC|HLA-Cw7|HLA-Cw7
C0482952|T201|COMP|4864-5|LNC|HLA-Cw8|HLA-Cw8
C0482953|T201|COMP|4865-2|LNC|HLA-Cw8|HLA-Cw8
C0482954|T201|COMP|4866-0|LNC|HLA-Cw9(w3)|HLA-Cw9(w3)
C0482955|T201|COMP|4867-8|LNC|HLA-Cw9(w3)|HLA-Cw9(w3)
C0482956|T201|COMP|4868-6|LNC|HLA-Dw10|HLA-Dw10
C0482957|T201|COMP|4869-4|LNC|HLA-Dw10|HLA-Dw10
C0482958|T201|COMP|4870-2|LNC|HLA-Dw11(w7)|HLA-Dw11(w7)
C0482959|T201|COMP|4871-0|LNC|HLA-Dw11(w7)|HLA-Dw11(w7)
C0482960|T201|COMP|4872-8|LNC|HLA-Dw12|HLA-Dw12
C0482961|T201|COMP|4873-6|LNC|HLA-Dw12|HLA-Dw12
C0482962|T201|COMP|4874-4|LNC|HLA-Dw13|HLA-Dw13
C0482963|T201|COMP|4875-1|LNC|HLA-Dw13|HLA-Dw13
C0482964|T201|COMP|4876-9|LNC|HLA-Dw14|HLA-Dw14
C0482965|T201|COMP|4877-7|LNC|HLA-Dw14|HLA-Dw14
C0482966|T201|COMP|4878-5|LNC|HLA-Dw15|HLA-Dw15
C0482967|T201|COMP|4879-3|LNC|HLA-Dw15|HLA-Dw15
C0482968|T201|COMP|4880-1|LNC|HLA-Dw16|HLA-Dw16
C0482969|T201|COMP|4881-9|LNC|HLA-Dw16|HLA-Dw16
C0482970|T201|COMP|4882-7|LNC|HLA-Dw17(w7)|HLA-Dw17(w7)
C0482971|T201|COMP|4883-5|LNC|HLA-Dw17(w7)|HLA-Dw17(w7)
C0482972|T201|COMP|4884-3|LNC|HLA-Dw18(w6)|HLA-Dw18(w6)
C0482973|T201|COMP|4885-0|LNC|HLA-Dw18(w6)|HLA-Dw18(w6)
C0482974|T201|COMP|4886-8|LNC|HLA-Dw19(w6)|HLA-Dw19(w6)
C0482975|T201|COMP|4887-6|LNC|HLA-Dw19(w6)|HLA-Dw19(w6)
C0482976|T201|COMP|4888-4|LNC|HLA-Dw1|HLA-Dw1
C0482977|T201|COMP|4889-2|LNC|HLA-Dw1|HLA-Dw1
C0482978|T201|COMP|4890-0|LNC|HLA-Dw20|HLA-Dw20
C0482979|T201|COMP|4891-8|LNC|HLA-Dw20|HLA-Dw20
C0482980|T201|COMP|4892-6|LNC|HLA-Dw21|HLA-Dw21
C0482981|T201|COMP|4893-4|LNC|HLA-Dw21|HLA-Dw21
C0482982|T201|COMP|4894-2|LNC|HLA-Dw22|HLA-Dw22
C0482983|T201|COMP|4895-9|LNC|HLA-Dw22|HLA-Dw22
C0482984|T201|COMP|4896-7|LNC|HLA-Dw23|HLA-Dw23
C0482985|T201|COMP|4897-5|LNC|HLA-Dw23|HLA-Dw23
C0482986|T201|COMP|4898-3|LNC|HLA-Dw24|HLA-Dw24
C0482987|T201|COMP|4899-1|LNC|HLA-Dw24|HLA-Dw24
C0482988|T201|COMP|4900-7|LNC|HLA-Dw25|HLA-Dw25
C0482989|T201|COMP|4901-5|LNC|HLA-Dw25|HLA-Dw25
C0482990|T201|COMP|4902-3|LNC|HLA-Dw26|HLA-Dw26
C0482991|T201|COMP|4903-1|LNC|HLA-Dw26|HLA-Dw26
C0482992|T201|COMP|4904-9|LNC|HLA-Dw2|HLA-Dw2
C0482993|T201|COMP|4905-6|LNC|HLA-Dw2|HLA-Dw2
C0482994|T201|COMP|4906-4|LNC|HLA-Dw3|HLA-Dw3
C0482995|T201|COMP|4907-2|LNC|HLA-Dw3|HLA-Dw3
C0482996|T201|COMP|4908-0|LNC|HLA-Dw4|HLA-Dw4
C0482997|T201|COMP|4909-8|LNC|HLA-Dw4|HLA-Dw4
C0482998|T201|COMP|4910-6|LNC|HLA-Dw5|HLA-Dw5
C0482999|T201|COMP|4911-4|LNC|HLA-Dw5|HLA-Dw5
C0483000|T201|COMP|4912-2|LNC|HLA-Dw6|HLA-Dw6
C0483001|T201|COMP|4913-0|LNC|HLA-Dw6|HLA-Dw6
C0483002|T201|COMP|4914-8|LNC|HLA-Dw7|HLA-Dw7
C0483003|T201|COMP|4915-5|LNC|HLA-Dw7|HLA-Dw7
C0483004|T201|COMP|4916-3|LNC|HLA-Dw8|HLA-Dw8
C0483005|T201|COMP|4917-1|LNC|HLA-Dw8|HLA-Dw8
C0483006|T201|COMP|4918-9|LNC|HLA-Dw9|HLA-Dw9
C0483007|T201|COMP|4919-7|LNC|HLA-Dw9|HLA-Dw9
C0483008|T201|COMP|4920-5|LNC|HLA-DPw1|HLA-DPw1
C0483009|T201|COMP|4921-3|LNC|HLA-DPw1|HLA-DPw1
C0483010|T201|COMP|4922-1|LNC|HLA-DPw2|HLA-DPw2
C0483011|T201|COMP|4923-9|LNC|HLA-DPw2|HLA-DPw2
C0483012|T201|COMP|4924-7|LNC|HLA-DPw3|HLA-DPw3
C0483013|T201|COMP|4925-4|LNC|HLA-DPw3|HLA-DPw3
C0483014|T201|COMP|4926-2|LNC|HLA-DPw4|HLA-DPw4
C0483015|T201|COMP|4927-0|LNC|HLA-DPw4|HLA-DPw4
C0483016|T201|COMP|4928-8|LNC|HLA-DPw5|HLA-DPw5
C0483017|T201|COMP|4929-6|LNC|HLA-DPw5|HLA-DPw5
C0483018|T201|COMP|4930-4|LNC|HLA-DPw6|HLA-DPw6
C0483019|T201|COMP|4931-2|LNC|HLA-DPw6|HLA-DPw6
C0483020|T201|COMP|4932-0|LNC|HLA-DQ1|HLA-DQ1
C0483021|T201|COMP|4933-8|LNC|HLA-DQ1|HLA-DQ1
C0483022|T201|COMP|4934-6|LNC|HLA-DQ2|HLA-DQ2
C0483023|T201|COMP|4935-3|LNC|HLA-DQ2|HLA-DQ2
C0483024|T201|COMP|4936-1|LNC|HLA-DQ3|HLA-DQ3
C0483025|T201|COMP|4937-9|LNC|HLA-DQ3|HLA-DQ3
C0483026|T201|COMP|4938-7|LNC|HLA-DQ4|HLA-DQ4
C0483027|T201|COMP|4939-5|LNC|HLA-DQ4|HLA-DQ4
C0483028|T201|COMP|4940-3|LNC|HLA-DQ5(1)|HLA-DQ5(1)
C0483029|T201|COMP|4941-1|LNC|HLA-DQ5(1)|HLA-DQ5(1)
C0483030|T201|COMP|4942-9|LNC|HLA-DQ6(1)|HLA-DQ6(1)
C0483031|T201|COMP|4943-7|LNC|HLA-DQ6(1)|HLA-DQ6(1)
C0483032|T201|COMP|4944-5|LNC|HLA-DQ7(3)|HLA-DQ7(3)
C0483033|T201|COMP|4945-2|LNC|HLA-DQ7(3)|HLA-DQ7(3)
C0483034|T201|COMP|4946-0|LNC|HLA-DQ8(3)|HLA-DQ8(3)
C0483035|T201|COMP|4947-8|LNC|HLA-DQ8(3)|HLA-DQ8(3)
C0483036|T201|COMP|4948-6|LNC|HLA-DQ9(3)|HLA-DQ9(3)
C0483037|T201|COMP|4949-4|LNC|HLA-DQ9(3)|HLA-DQ9(3)
C0483038|T201|COMP|4950-2|LNC|HLA-DR10|HLA-DR10
C0483039|T201|COMP|4951-0|LNC|HLA-DR10|HLA-DR10
C0483040|T201|COMP|4952-8|LNC|HLA-DR11(5)|HLA-DR11(5)
C0483041|T201|COMP|4953-6|LNC|HLA-DR11(5)|HLA-DR11(5)
C0483042|T201|COMP|4954-4|LNC|HLA-DR12(5)|HLA-DR12(5)
C0483043|T201|COMP|4955-1|LNC|HLA-DR12(5)|HLA-DR12(5)
C0483044|T201|COMP|4956-9|LNC|HLA-DR13(6)|HLA-DR13(6)
C0483045|T201|COMP|4957-7|LNC|HLA-DR13(6)|HLA-DR13(6)
C0483046|T201|COMP|4958-5|LNC|HLA-DR14(6)|HLA-DR14(6)
C0483047|T201|COMP|4959-3|LNC|HLA-DR14(6)|HLA-DR14(6)
C0483048|T201|COMP|4960-1|LNC|HLA-DR15(2)|HLA-DR15(2)
C0483049|T201|COMP|4961-9|LNC|HLA-DR15(2)|HLA-DR15(2)
C0483050|T201|COMP|4962-7|LNC|HLA-DR16(2)|HLA-DR16(2)
C0483051|T201|COMP|4963-5|LNC|HLA-DR16(2)|HLA-DR16(2)
C0483052|T201|COMP|4964-3|LNC|HLA-DR17(3)|HLA-DR17(3)
C0483053|T201|COMP|4965-0|LNC|HLA-DR17(3)|HLA-DR17(3)
C0483054|T201|COMP|4966-8|LNC|HLA-DR18(3)|HLA-DR18(3)
C0483055|T201|COMP|4967-6|LNC|HLA-DR18(3)|HLA-DR18(3)
C0483056|T201|COMP|4968-4|LNC|HLA-DR52|HLA-DR52
C0483057|T201|COMP|4969-2|LNC|HLA-DR52|HLA-DR52
C0483058|T201|COMP|4970-0|LNC|HLA-DR53|HLA-DR53
C0483059|T201|COMP|4971-8|LNC|HLA-DR53|HLA-DR53
C0483060|T201|COMP|4972-6|LNC|HLA-DR6|HLA-DR6
C0483061|T201|COMP|4973-4|LNC|HLA-DR6|HLA-DR6
C0483062|T201|COMP|4974-2|LNC|HLA-DR8|HLA-DR8
C0483063|T201|COMP|4975-9|LNC|HLA-DR8|HLA-DR8
C0483064|T201|COMP|4976-7|LNC|HLA-DR1|HLA-DR1
C0483065|T201|COMP|4977-5|LNC|HLA-DR1|HLA-DR1
C0483066|T201|COMP|4978-3|LNC|HLA-DR2|HLA-DR2
C0483067|T201|COMP|4979-1|LNC|HLA-DR2|HLA-DR2
C0483068|T201|COMP|4980-9|LNC|HLA-DR3|HLA-DR3
C0483069|T201|COMP|4981-7|LNC|HLA-DR3|HLA-DR3
C0483070|T201|COMP|4982-5|LNC|HLA-DR4|HLA-DR4
C0483071|T201|COMP|4983-3|LNC|HLA-DR4|HLA-DR4
C0483072|T201|COMP|4984-1|LNC|HLA-DR5|HLA-DR5
C0483073|T201|COMP|4985-8|LNC|HLA-DR5|HLA-DR5
C0483074|T201|COMP|4986-6|LNC|HLA-DR7|HLA-DR7
C0483075|T201|COMP|4987-4|LNC|HLA-DR7|HLA-DR7
C0483076|T201|COMP|4988-2|LNC|HLA-DR9|HLA-DR9
C0483077|T201|COMP|4989-0|LNC|HLA-DR9|HLA-DR9
C0483078|T201|COMP|6575-5|LNC|Escherichia coli verotoxin 1 Ab|Escherichia coli verotoxin 1 Ab
C0483079|T201|COMP|6577-1|LNC|Escherichia coli verotoxin 2 Ab|Escherichia coli verotoxin 2 Ab
C0483082|T201|COMP|5097-1|LNC|Cold agglutinin|Cold agglutinin
C0483083|T201|COMP|5098-9|LNC|Cold agglutinin|Cold agglutinin
C0483084|T201|COMP|5234-0|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C0483085|T201|COMP|5235-7|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C0483086|T201|COMP|5276-1|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C0483087|T201|COMP|5275-3|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C0483088|T201|COMP|5301-7|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0483089|T201|COMP|5302-5|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0483090|T201|COMP|5348-8|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C0483091|T201|COMP|5349-6|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C0483092|T201|COMP|5351-2|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C0483093|T201|COMP|5352-0|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C0483094|T201|COMP|5353-8|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C0483095|T201|COMP|5354-6|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C0483096|T201|COMP|5355-3|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0483097|T201|COMP|5356-1|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0483098|T201|COMP|5357-9|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0483099|T201|COMP|5361-1|LNC|Spermatozoa Ab|Spermatozoa Ab
C0483100|T201|COMP|5379-3|LNC|Platelet Ab|Platelet Ab
C0483101|T201|COMP|5380-1|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C0483102|T201|COMP|5381-9|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C0483103|T201|COMP|5415-5|LNC|CD10+CD20+|CD10+CD20+
C0483104|T201|COMP|5438-7|LNC|CD16+CD56+CD3-|CD16+CD56+CD3-
C0483105|T201|COMP|6707-4|LNC|CD16-CD57+|CD16-CD57+
C0483106|T201|COMP|5440-3|LNC|CD16+CD57-|CD16+CD57-
C0483107|T201|COMP|5445-2|LNC|CD19+SmIg kappa+|CD19+SmIg kappa+
C0483108|T201|COMP|5446-0|LNC|CD19+SmIg lambda+|CD19+SmIg lambda+
C0483109|T201|COMP|5451-0|LNC|CD22+CD19+|CD22+CD19+
C0483110|T201|COMP|694-0|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0483111|T201|COMP|5460-1|LNC|CD3+DR+|CD3+DR+
C0483112|T201|COMP|5466-8|LNC|CD34+DR+|CD34+DR+
C0483113|T201|COMP|5473-4|LNC|CD4+CD8+|CD4+CD8+
C0483114|T201|COMP|5498-1|LNC|CD5+CD2-|CD5+CD2-
C0483115|T201|COMP|5524-4|LNC|CD7+CD3-|CD7+CD3-
C0483116|T201|COMP|5566-5|LNC|Acetone|Acetone
C0483117|T201|COMP|5641-6|LNC|Ethanol|Ethanol
C0483118|T201|COMP|5690-3|LNC|Methanol|Methanol
C0483119|T201|COMP|5691-1|LNC|Methanol|Methanol
C0483120|T201|COMP|5693-7|LNC|Methanol|Methanol
C0483121|T201|COMP|5309-0|LNC|Rickettsia spotted fever group Ab|Rickettsia spotted fever group Ab
C0483122|T201|COMP|5310-8|LNC|Rickettsia spotted fever group Ab|Rickettsia spotted fever group Ab
C0483123|T201|COMP|5311-6|LNC|Rickettsia spotted fever group Ab|Rickettsia spotted fever group Ab
C0483124|T201|COMP|5312-4|LNC|Rickettsia spotted fever group Ab.IgG|Rickettsia spotted fever group Ab.IgG
C0483125|T201|COMP|5313-2|LNC|Rickettsia spotted fever group Ab.IgG|Rickettsia spotted fever group Ab.IgG
C0483126|T201|COMP|5314-0|LNC|Rickettsia spotted fever group Ab.IgM|Rickettsia spotted fever group Ab.IgM
C0483127|T201|COMP|5702-6|LNC|Nickel|Nickel
C0483128|T201|COMP|5315-7|LNC|Rickettsia spotted fever group Ab.IgM|Rickettsia spotted fever group Ab.IgM
C0483129|T201|COMP|5316-5|LNC|Rickettsia typhus group Ab|Rickettsia typhus group Ab
C0483130|T201|COMP|5317-3|LNC|Rickettsia typhus group Ab|Rickettsia typhus group Ab
C0483131|T201|COMP|5318-1|LNC|Rickettsia typhus group Ab|Rickettsia typhus group Ab
C0483132|T201|COMP|5319-9|LNC|Rickettsia typhus group Ab.IgG|Rickettsia typhus group Ab.IgG
C0483133|T201|COMP|5320-7|LNC|Rickettsia typhus group Ab.IgG|Rickettsia typhus group Ab.IgG
C0483134|T201|COMP|5321-5|LNC|Rickettsia typhus group Ab.IgM|Rickettsia typhus group Ab.IgM
C0483135|T201|COMP|5322-3|LNC|Rickettsia typhus group Ab.IgM|Rickettsia typhus group Ab.IgM
C0483136|T201|COMP|5326-4|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C0483137|T201|COMP|5327-2|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C0483138|T201|COMP|5336-3|LNC|Saccharomonospora viridis Ab|Saccharomonospora viridis Ab
C0483139|T201|COMP|5040-1|LNC|Actinomyces sp Ab|Actinomyces sp Ab
C0483140|T201|COMP|5058-3|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0483141|T201|COMP|6313-1|LNC|Blastomyces dermatitidis Ag|Blastomyces dermatitidis Ag
C0483142|T201|COMP|6314-9|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C0483143|T201|COMP|5059-1|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C0483144|T201|COMP|5073-2|LNC|La Crosse virus Ab|La Crosse virus Ab
C0483145|T201|COMP|5100-3|LNC|Coxiella burnetii Ab|Coxiella burnetii Ab
C0483146|T201|COMP|5115-1|LNC|Corynebacterium diphtheriae Ab|Corynebacterium diphtheriae Ab
C0483147|T201|COMP|5116-9|LNC|Corynebacterium diphtheriae Ab|Corynebacterium diphtheriae Ab
C0483148|T201|COMP|566-0|LNC|Cryptosporidium sp Ag|Cryptosporidium sp Ag
C0483149|T201|COMP|6382-6|LNC|Dengue virus Ab|Dengue virus Ab
C0483150|T201|COMP|6383-4|LNC|Dengue virus Ab|Dengue virus Ab
C0483151|T201|COMP|5153-2|LNC|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C0483152|T201|COMP|5154-0|LNC|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C0483153|T201|COMP|5155-7|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0483154|T201|COMP|5156-5|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0483155|T201|COMP|5157-3|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0483156|T201|COMP|5158-1|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0483157|T201|COMP|5159-9|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0483158|T201|COMP|5160-7|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0483159|T201|COMP|6400-6|LNC|Ehrlichia canis Ab|Ehrlichia canis Ab
C0483160|T201|COMP|6401-4|LNC|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C0483161|T201|COMP|6402-2|LNC|Ehrlichia chaffeensis Ab.IgM|Ehrlichia chaffeensis Ab.IgM
C0483162|T201|COMP|6403-0|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C0483163|T201|COMP|6404-8|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C0483164|T201|COMP|6405-5|LNC|Ehrlichia sp Ab|Ehrlichia sp Ab
C0483165|T201|COMP|6414-7|LNC|Haemophilus influenzae A Ag|Haemophilus influenzae A Ag
C0483166|T201|COMP|6416-2|LNC|Haemophilus influenzae D Ag|Haemophilus influenzae D Ag
C0483167|T201|COMP|6417-0|LNC|Haemophilus influenzae E Ag|Haemophilus influenzae E Ag
C0483168|T201|COMP|6418-8|LNC|Haemophilus influenzae F Ag|Haemophilus influenzae F Ag
C0483169|T201|COMP|5189-6|LNC|Hepatitis B virus little e Ab|Hepatitis B virus little e Ab
C0483170|T201|COMP|5190-4|LNC|Hepatitis B virus little e Ab|Hepatitis B virus little e Ab
C0483171|T201|COMP|5191-2|LNC|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C0483172|T201|COMP|5192-0|LNC|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C0483173|T201|COMP|6457-6|LNC|DNA double strand Ab|DNA double strand Ab
C0483174|T201|COMP|623-9|LNC|Bacteria identified|Bacteria identified
C0483526|T201|COMP|6975-7|LNC|Amikacin|Amikacin
C0483527|T201|COMP|6976-5|LNC|Amoxicillin|Amoxicillin
C0483528|T201|COMP|6977-3|LNC|Amoxicillin+Clavulanate|Amoxicillin+Clavulanate
C0483529|T201|COMP|6978-1|LNC|Amphotericin B|Amphotericin B
C0483530|T201|COMP|6979-9|LNC|Ampicillin|Ampicillin
C0483531|T201|COMP|6980-7|LNC|Ampicillin+Sulbactam|Ampicillin+Sulbactam
C0483532|T201|COMP|6981-5|LNC|Azithromycin|Azithromycin
C0483533|T201|COMP|6982-3|LNC|Aztreonam|Aztreonam
C0483534|T201|COMP|6827-0|LNC|Bacitracin|Bacitracin
C0483535|T201|COMP|6983-1|LNC|Bacitracin|Bacitracin
C0483536|T201|COMP|6984-9|LNC|Beta lactamase.extended spectrum|Beta lactamase.extended spectrum
C0483537|T201|COMP|6985-6|LNC|Beta lactamase.usual|Beta lactamase.usual
C0483538|T201|COMP|6986-4|LNC|Cefaclor|Cefaclor
C0483539|T201|COMP|6643-1|LNC|Cefepime|Cefepime
C0483540|T201|COMP|6644-9|LNC|Cefepime|Cefepime
C0483541|T201|COMP|8272-7|LNC|Cefepime|Cefepime
C0483542|T201|COMP|6987-2|LNC|Cefepime|Cefepime
C0483543|T201|COMP|8273-5|LNC|Cefepime|Cefepime
C0483544|T201|COMP|6988-0|LNC|Cefodizime|Cefodizime
C0483545|T201|COMP|6989-8|LNC|Cefotaxime|Cefotaxime
C0483546|T201|COMP|6990-6|LNC|cefoTEtan|cefoTEtan
C0483547|T201|COMP|6991-4|LNC|cefOXitin|cefOXitin
C0483548|T201|COMP|8274-3|LNC|Cefpirome|Cefpirome
C0483549|T201|COMP|8275-0|LNC|Cefpirome|Cefpirome
C0483550|T201|COMP|8276-8|LNC|Cefpirome|Cefpirome
C0483551|T201|COMP|6992-2|LNC|Cefpirome|Cefpirome
C0483552|T201|COMP|6650-6|LNC|Cefpirome|Cefpirome
C0483553|T201|COMP|6993-0|LNC|Cefpodoxime|Cefpodoxime
C0483554|T201|COMP|6994-8|LNC|Cefprozil|Cefprozil
C0483555|T201|COMP|6995-5|LNC|cefTAZidime|cefTAZidime
C0483556|T201|COMP|6996-3|LNC|Ceftibuten|Ceftibuten
C0483557|T201|COMP|6997-1|LNC|Ceftizoxime|Ceftizoxime
C0483558|T201|COMP|6998-9|LNC|cefTRIAXone|cefTRIAXone
C0483559|T201|COMP|6999-7|LNC|Cefuroxime.parenteral|Cefuroxime.parenteral
C0483560|T201|COMP|7000-3|LNC|Cephalothin|Cephalothin
C0483561|T201|COMP|7001-1|LNC|Chloramphenicol|Chloramphenicol
C0483562|T201|COMP|7002-9|LNC|Ciprofloxacin|Ciprofloxacin
C0483563|T201|COMP|7003-7|LNC|Clarithromycin|Clarithromycin
C0483564|T201|COMP|7004-5|LNC|Clinafloxacin|Clinafloxacin
C0483565|T201|COMP|7005-2|LNC|Clindamycin|Clindamycin
C0483566|T201|COMP|7006-0|LNC|Demeclocycline|Demeclocycline
C0483567|T201|COMP|7007-8|LNC|Dirithromycin|Dirithromycin
C0483568|T201|COMP|7008-6|LNC|Doxycycline|Doxycycline
C0483569|T201|COMP|7009-4|LNC|Erythromycin|Erythromycin
C0483570|T201|COMP|7010-2|LNC|Ethambutol|Ethambutol
C0483571|T201|COMP|7011-0|LNC|Ethionamide|Ethionamide
C0483572|T201|COMP|7012-8|LNC|Fleroxacin|Fleroxacin
C0483573|T201|COMP|7013-6|LNC|Fluconazole|Fluconazole
C0483574|T201|COMP|7014-4|LNC|5-Fluorocytosine|5-Fluorocytosine
C0483575|T201|COMP|7015-1|LNC|Fusidate|Fusidate
C0483576|T201|COMP|7016-9|LNC|Gentamicin|Gentamicin
C0483577|T201|COMP|7017-7|LNC|Gentamicin.high potency|Gentamicin.high potency
C0483578|T201|COMP|7018-5|LNC|Gentamicin.high potency|Gentamicin.high potency
C0483579|T201|COMP|7019-3|LNC|Imipenem|Imipenem
C0483580|T201|COMP|7020-1|LNC|Isoniazid|Isoniazid
C0483581|T201|COMP|7021-9|LNC|Itraconazole|Itraconazole
C0483582|T201|COMP|7022-7|LNC|Kanamycin|Kanamycin
C0483583|T201|COMP|7023-5|LNC|Kanamycin.high potency|Kanamycin.high potency
C0483584|T201|COMP|7024-3|LNC|Kanamycin.high potency|Kanamycin.high potency
C0483585|T201|COMP|7025-0|LNC|Ketoconazole|Ketoconazole
C0483586|T201|COMP|7026-8|LNC|levoFLOXacin|levoFLOXacin
C0483587|T201|COMP|7027-6|LNC|Loracarbef|Loracarbef
C0483588|T201|COMP|7028-4|LNC|Amdinocillin|Amdinocillin
C0483589|T201|COMP|6651-4|LNC|Meropenem|Meropenem
C0483590|T201|COMP|6652-2|LNC|Meropenem|Meropenem
C0483591|T201|COMP|6653-0|LNC|Meropenem|Meropenem
C0483592|T201|COMP|7029-2|LNC|Meropenem|Meropenem
C0483593|T201|COMP|6654-8|LNC|Meropenem|Meropenem
C0483594|T201|COMP|7030-0|LNC|Methicillin|Methicillin
C0483595|T201|COMP|7031-8|LNC|metroNIDAZOLE|metroNIDAZOLE
C0483596|T201|COMP|7032-6|LNC|Minocycline|Minocycline
C0483597|T201|COMP|7033-4|LNC|Mupirocin|Mupirocin
C0483598|T201|COMP|7034-2|LNC|Nalidixate|Nalidixate
C0483599|T201|COMP|7035-9|LNC|Netilmicin|Netilmicin
C0483600|T201|COMP|7036-7|LNC|Nitrofurantoin|Nitrofurantoin
C0483601|T201|COMP|7037-5|LNC|Norfloxacin|Norfloxacin
C0483602|T201|COMP|7038-3|LNC|Ofloxacin|Ofloxacin
C0483603|T201|COMP|7039-1|LNC|Oxacillin|Oxacillin
C0483604|T201|COMP|7040-9|LNC|Pefloxacin|Pefloxacin
C0483605|T201|COMP|6932-8|LNC|Penicillin|Penicillin
C0483606|T201|COMP|7041-7|LNC|Penicillin G|Penicillin G
C0483607|T201|COMP|7042-5|LNC|Penicillin V|Penicillin V
C0483608|T201|COMP|7043-3|LNC|Piperacillin|Piperacillin
C0483609|T201|COMP|7044-1|LNC|Piperacillin+Tazobactam|Piperacillin+Tazobactam
C0483610|T201|COMP|7045-8|LNC|rifAMPin|rifAMPin
C0483611|T201|COMP|7046-6|LNC|Roxithromycin|Roxithromycin
C0483612|T201|COMP|7047-4|LNC|Sparfloxacin|Sparfloxacin
C0483613|T201|COMP|7048-2|LNC|Streptomycin|Streptomycin
C0483614|T201|COMP|6933-6|LNC|Streptomycin.high potency|Streptomycin.high potency
C0483615|T201|COMP|7049-0|LNC|Streptomycin.high potency|Streptomycin.high potency
C0483616|T201|COMP|7050-8|LNC|sulfADIAZINE|sulfADIAZINE
C0483617|T201|COMP|7051-6|LNC|Teicoplanin|Teicoplanin
C0483618|T201|COMP|7052-4|LNC|Tetracycline|Tetracycline
C0483619|T201|COMP|7053-2|LNC|Ticarcillin|Ticarcillin
C0483620|T201|COMP|7054-0|LNC|Ticarcillin+Clavulanate|Ticarcillin+Clavulanate
C0483621|T201|COMP|7055-7|LNC|Tobramycin|Tobramycin
C0483622|T201|COMP|7056-5|LNC|Trimethoprim|Trimethoprim
C0483623|T201|COMP|7057-3|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0483624|T201|COMP|7058-1|LNC|Trovafloxacin|Trovafloxacin
C0483625|T201|COMP|7059-9|LNC|Vancomycin|Vancomycin
C0483626|T201|COMP|7060-7|LNC|Haliotis spp Ab.IgE|Haliotis spp Ab.IgE
C0483627|T201|COMP|6711-6|LNC|Acetaminophen Ab.IgE|Acetaminophen Ab.IgE
C0483628|T201|COMP|7108-4|LNC|Acetylsalicylate Ab.IgE|Acetylsalicylate Ab.IgE
C0483629|T201|COMP|7061-5|LNC|Alder Ab.IgG|Alder Ab.IgG
C0483630|T201|COMP|7062-3|LNC|Alnus rubra Ab.IgE|Alnus rubra Ab.IgE
C0483631|T201|COMP|7063-1|LNC|Alnus rugosa Ab.IgE|Alnus rugosa Ab.IgE
C0483632|T201|COMP|7064-9|LNC|Alnus rhombifolia Ab.IgE|Alnus rhombifolia Ab.IgE
C0483633|T201|COMP|7065-6|LNC|Medicago sativa Ab.IgE|Medicago sativa Ab.IgE
C0483634|T201|COMP|7066-4|LNC|Medicago sativa Ab.IgG|Medicago sativa Ab.IgG
C0483635|T201|COMP|7067-2|LNC|Medicago sativa pollen Ab.IgE|Medicago sativa pollen Ab.IgE
C0483636|T201|COMP|7068-0|LNC|Algae Ab.IgE|Algae Ab.IgE
C0483637|T201|COMP|7069-8|LNC|Pimenta dioica Ab.IgE|Pimenta dioica Ab.IgE
C0483638|T201|COMP|7070-6|LNC|Prunus dulcis Ab.IgG|Prunus dulcis Ab.IgG
C0483639|T201|COMP|7071-4|LNC|Prunus dulcis basophil bound Ab|Prunus dulcis basophil bound Ab
C0483640|T201|COMP|7072-2|LNC|Prunus dulcis tree Ab.IgE|Prunus dulcis tree Ab.IgE
C0483641|T201|COMP|7073-0|LNC|Amylase Ab.IgE|Amylase Ab.IgE
C0483642|T201|COMP|6020-2|LNC|Alternaria alternata Ab.IgE|Alternaria alternata Ab.IgE
C0483643|T201|COMP|7074-8|LNC|Alternaria sp Ab.IgE|Alternaria sp Ab.IgE
C0483644|T201|COMP|7075-5|LNC|Alternaria sp Ab.IgG|Alternaria sp Ab.IgG
C0483646|T201|COMP|7077-1|LNC|Alternaria alternata basophil bound Ab|Alternaria alternata basophil bound Ab
C0483647|T201|COMP|6829-6|LNC|Amoxicillin Ab.IgE|Amoxicillin Ab.IgE
C0483648|T201|COMP|6712-4|LNC|Ampicillin Ab.IgE|Ampicillin Ab.IgE
C0483649|T201|COMP|7078-9|LNC|Ampicillin Ab.IgM|Ampicillin Ab.IgM
C0483650|T201|COMP|7079-7|LNC|Engraulis encrasicolus Ab.IgE|Engraulis encrasicolus Ab.IgE
C0483651|T201|COMP|7080-5|LNC|Engraulis encrasicolus Ab.IgG|Engraulis encrasicolus Ab.IgG
C0483652|T201|COMP|7081-3|LNC|Pimpinella anisum Ab.IgE|Pimpinella anisum Ab.IgE
C0483653|T201|COMP|7082-1|LNC|Monomorium minimum Ab.IgG|Monomorium minimum Ab.IgG
C0483654|T201|COMP|7083-9|LNC|Monomorium minimum basophil bound Ab|Monomorium minimum basophil bound Ab
C0483655|T201|COMP|7084-7|LNC|Solenopsis geminata Ab.IgG|Solenopsis geminata Ab.IgG
C0483656|T201|COMP|6117-6|LNC|Solenopsis invicta Ab.IgE|Solenopsis invicta Ab.IgE
C0483657|T201|COMP|7086-2|LNC|Solenopsis richteri Ab.IgE|Solenopsis richteri Ab.IgE
C0483658|T201|COMP|7087-0|LNC|Pogonomyrmex barbatus Ab.IgE|Pogonomyrmex barbatus Ab.IgE
C0483659|T201|COMP|7088-8|LNC|Malus sylvestris Ab.IgG|Malus sylvestris Ab.IgG
C0483660|T201|COMP|7089-6|LNC|Malus sylvestris basophil bound Ab|Malus sylvestris basophil bound Ab
C0483661|T201|COMP|7090-4|LNC|Malus sylvestris tree Ab.IgE|Malus sylvestris tree Ab.IgE
C0483662|T201|COMP|7091-2|LNC|Prunus armeniaca Ab.IgE|Prunus armeniaca Ab.IgE
C0483663|T201|COMP|7092-0|LNC|Prunus armeniaca Ab.IgG|Prunus armeniaca Ab.IgG
C0483664|T201|COMP|7093-8|LNC|Maranta arundinacea Ab.IgE|Maranta arundinacea Ab.IgE
C0483665|T201|COMP|7094-6|LNC|Cynara scolymus Ab.IgE|Cynara scolymus Ab.IgE
C0483666|T201|COMP|7095-3|LNC|Fraxinus velutina Ab.IgE|Fraxinus velutina Ab.IgE
C0483667|T201|COMP|6832-0|LNC|Fraxinus latifolia Ab.IgE|Fraxinus latifolia Ab.IgE
C0483668|T201|COMP|7097-9|LNC|Ash Ab.IgG|Ash Ab.IgG
C0483669|T201|COMP|7098-7|LNC|Fraxinus americana basophil bound Ab|Fraxinus americana basophil bound Ab
C0483670|T201|COMP|7099-5|LNC|Asparagus officinalis Ab.IgE|Asparagus officinalis Ab.IgE
C0483671|T201|COMP|7100-1|LNC|Asparagus officinalis Ab.IgG|Asparagus officinalis Ab.IgG
C0483672|T201|COMP|7101-9|LNC|Populus tremula Ab.IgE|Populus tremula Ab.IgE
C0483673|T201|COMP|7102-7|LNC|Populus tremula Ab.IgG|Populus tremula Ab.IgG
C0483674|T201|COMP|7103-5|LNC|Aspergillus fumigatus Ab.IgG|Aspergillus fumigatus Ab.IgG
C0483675|T201|COMP|7104-3|LNC|Aspergillus fumigatus basophil bound Ab|Aspergillus fumigatus basophil bound Ab
C0483676|T201|COMP|7105-0|LNC|Aspergillus nidulans Ab.IgE|Aspergillus nidulans Ab.IgE
C0483677|T201|COMP|6830-4|LNC|Aspergillus niger Ab.IgE|Aspergillus niger Ab.IgE
C0483678|T201|COMP|7106-8|LNC|Aspergillus sp Ab.IgE|Aspergillus sp Ab.IgE
C0483679|T201|COMP|7107-6|LNC|Aspergillus sp Ab.IgG|Aspergillus sp Ab.IgG
C0483680|T201|COMP|7109-2|LNC|Persea americana Ab.IgG|Persea americana Ab.IgG
C0483681|T201|COMP|7110-0|LNC|Baccharis spp Ab.IgE|Baccharis spp Ab.IgE
C0483682|T201|COMP|7112-6|LNC|Musa spp Ab.IgG|Musa spp Ab.IgG
C0483683|T201|COMP|7113-4|LNC|Musa spp basophil bound Ab|Musa spp basophil bound Ab
C0483684|T201|COMP|7114-2|LNC|Hordeum vulgare Ab.IgG|Hordeum vulgare Ab.IgG
C0483685|T201|COMP|7115-9|LNC|Hordeum vulgare basophil bound Ab|Hordeum vulgare basophil bound Ab
C0483686|T201|COMP|7116-7|LNC|Hordeum vulgare pollen Ab.IgE|Hordeum vulgare pollen Ab.IgE
C0483687|T201|COMP|7117-5|LNC|(Avena sativa+Hordeum vulgare) Ab.IgE|(Avena sativa+Hordeum vulgare) Ab.IgE
C0483688|T201|COMP|7118-3|LNC|Ocimum basilicum Ab.IgE|Ocimum basilicum Ab.IgE
C0483689|T201|COMP|7119-1|LNC|Ocimum basilicum Ab.IgG|Ocimum basilicum Ab.IgG
C0483690|T201|COMP|7120-9|LNC|Micropterus salmoides Ab.IgE|Micropterus salmoides Ab.IgE
C0483691|T201|COMP|7121-7|LNC|Bassiai Ab.IgE|Bassiai Ab.IgE
C0483692|T201|COMP|7122-5|LNC|Tilia americana Ab.IgE|Tilia americana Ab.IgE
C0483693|T201|COMP|7123-3|LNC|Myrica spp Ab.IgE|Myrica spp Ab.IgE
C0483694|T201|COMP|7124-1|LNC|Myrica spp pollen Ab.IgE|Myrica spp pollen Ab.IgE
C0483695|T201|COMP|7125-8|LNC|Laurus nobilis Ab.IgE|Laurus nobilis Ab.IgE
C0483696|T201|COMP|7126-6|LNC|Laurus nobilis Ab.IgG|Laurus nobilis Ab.IgG
C0483697|T201|COMP|6831-2|LNC|Bean green Ab.IgE|Bean green Ab.IgE
C0483698|T201|COMP|7127-4|LNC|Bean green Ab.IgG|Bean green Ab.IgG
C0483699|T201|COMP|7128-2|LNC|Bean green basophil bound Ab|Bean green basophil bound Ab
C0483700|T201|COMP|7129-0|LNC|Bean kidney red Ab.IgE|Bean kidney red Ab.IgE
C0483701|T201|COMP|7130-8|LNC|Bean kidney red Ab.IgG|Bean kidney red Ab.IgG
C0483702|T201|COMP|7131-6|LNC|Phaseolus limensis Ab.IgE|Phaseolus limensis Ab.IgE
C0483703|T201|COMP|7132-4|LNC|Phaseolus limensis Ab.IgG|Phaseolus limensis Ab.IgG
C0483704|T201|COMP|7133-2|LNC|Vigna radiata Ab.IgE|Vigna radiata Ab.IgE
C0483705|T201|COMP|7134-0|LNC|Vigna radiata Ab.IgG|Vigna radiata Ab.IgG
C0483706|T201|COMP|7135-7|LNC|Bean pinto Ab.IgE|Bean pinto Ab.IgE
C0483707|T201|COMP|7136-5|LNC|Bean pinto Ab.IgG|Bean pinto Ab.IgG
C0483708|T201|COMP|6735-5|LNC|Glycine max Ab.IgG|Glycine max Ab.IgG
C0483709|T201|COMP|7137-3|LNC|Glycine max basophil bound Ab|Glycine max basophil bound Ab
C0483710|T201|COMP|7138-1|LNC|Glycine max dust Ab.IgE|Glycine max dust Ab.IgE
C0483711|T201|COMP|7139-9|LNC|Bean string Ab.IgG|Bean string Ab.IgG
C0483712|T201|COMP|7140-7|LNC|Bean wax Ab.IgE|Bean wax Ab.IgE
C0483713|T201|COMP|7141-5|LNC|Bean white Ab.IgG|Bean white Ab.IgG
C0483714|T201|COMP|7142-3|LNC|Bean yellow Ab.IgG|Bean yellow Ab.IgG
C0483715|T201|COMP|6844-5|LNC|Apis mellifera Ab.IgE|Apis mellifera Ab.IgE
C0483716|T201|COMP|6727-2|LNC|Apis mellifera Ab.IgG|Apis mellifera Ab.IgG
C0483717|T201|COMP|6714-0|LNC|Beef Ab.IgG|Beef Ab.IgG
C0483718|T201|COMP|7143-1|LNC|Beef basophil bound Ab|Beef basophil bound Ab
C0483719|T201|COMP|7144-9|LNC|Liver beef basophil bound Ab|Liver beef basophil bound Ab
C0483720|T201|COMP|7145-6|LNC|Beet Ab.IgG|Beet Ab.IgG
C0483721|T201|COMP|7146-4|LNC|Beet red Ab.IgE|Beet red Ab.IgE
C0483722|T201|COMP|7147-2|LNC|Beta vulgaris Ab.IgE|Beta vulgaris Ab.IgE
C0483723|T201|COMP|7148-0|LNC|Berry Ab.IgE|Berry Ab.IgE
C0483724|T201|COMP|7149-8|LNC|Bipolanis curvularia Ab.IgE|Bipolanis curvularia Ab.IgE
C0483725|T201|COMP|7150-6|LNC|Birch White Ab.IgE|Birch White Ab.IgE
C0483726|T201|COMP|7151-4|LNC|Rubus fruticosus Ab.IgE|Rubus fruticosus Ab.IgE
C0483727|T201|COMP|7152-2|LNC|Vaccinium myrtillus Ab.IgE|Vaccinium myrtillus Ab.IgE
C0483728|T201|COMP|7153-0|LNC|Vaccinium myrtillus Ab.IgG|Vaccinium myrtillus Ab.IgG
C0483729|T201|COMP|7154-8|LNC|Vaccinium myrtillus basophil bound Ab|Vaccinium myrtillus basophil bound Ab
C0483730|T201|COMP|7155-5|LNC|Acer negundo Ab.IgE|Acer negundo Ab.IgE
C0483731|T201|COMP|7156-3|LNC|Acer negundo Ab.IgG|Acer negundo Ab.IgG
C0483732|T201|COMP|7157-1|LNC|Bertholletia excelsa Ab.IgG|Bertholletia excelsa Ab.IgG
C0483733|T201|COMP|7158-9|LNC|Bertholletia excelsa basophil bound Ab|Bertholletia excelsa basophil bound Ab
C0483734|T201|COMP|7159-7|LNC|Brassica oleracea var italica Ab.IgG|Brassica oleracea var italica Ab.IgG
C0483735|T201|COMP|7160-5|LNC|Brassica oleracea var gemmifera Ab.IgE|Brassica oleracea var gemmifera Ab.IgE
C0483736|T201|COMP|7161-3|LNC|Brassica oleracea var gemmifera Ab.IgG|Brassica oleracea var gemmifera Ab.IgG
C0483737|T201|COMP|7162-1|LNC|Fagopyrum esculentum Ab.IgG|Fagopyrum esculentum Ab.IgG
C0483740|T201|COMP|7164-7|LNC|Hymenoclea salsola Ab.IgE|Hymenoclea salsola Ab.IgE
C0483741|T201|COMP|7166-2|LNC|Burweed Ab.IgE|Burweed Ab.IgE
C0483742|T201|COMP|7167-0|LNC|Butterfly Ab.IgE|Butterfly Ab.IgE
C0483743|T201|COMP|7168-8|LNC|Buttermilk basophil bound Ab|Buttermilk basophil bound Ab
C0483744|T201|COMP|7169-6|LNC|Brassica oleracea var capitata Ab.IgE|Brassica oleracea var capitata Ab.IgE
C0483745|T201|COMP|7170-4|LNC|Brassica oleracea var capitata Ab.IgG|Brassica oleracea var capitata Ab.IgG
C0483746|T201|COMP|7171-2|LNC|Canary feather Ab.IgE|Canary feather Ab.IgE
C0483747|T201|COMP|9729-5|LNC|Canary serum proteins Ab.IgE|Canary serum proteins Ab.IgE
C0483748|T201|COMP|7172-0|LNC|Candida albicans Ab.IgG|Candida albicans Ab.IgG
C0483749|T201|COMP|7173-8|LNC|Candida albicans basophil bound Ab|Candida albicans basophil bound Ab
C0483750|T201|COMP|7174-6|LNC|Candida sp Ab.IgG|Candida sp Ab.IgG
C0483753|T201|COMP|7177-9|LNC|Cucumis melo spp basophil bound Ab|Cucumis melo spp basophil bound Ab
C0483754|T201|COMP|7178-7|LNC|Carum carvi Ab.IgE|Carum carvi Ab.IgE
C0483755|T201|COMP|7179-5|LNC|Ceratonia siliqua Ab.IgE|Ceratonia siliqua Ab.IgE
C0483756|T201|COMP|7180-3|LNC|Daucus carota Ab.IgG|Daucus carota Ab.IgG
C0483757|T201|COMP|7181-1|LNC|Daucus carota basophil bound Ab|Daucus carota basophil bound Ab
C0483758|T201|COMP|7182-9|LNC|Casein Ab.IgG|Casein Ab.IgG
C0483759|T201|COMP|6718-1|LNC|Anacardium occidentale Ab.IgE|Anacardium occidentale Ab.IgE
C0483760|T201|COMP|7183-7|LNC|Anacardium occidentale Ab.IgG|Anacardium occidentale Ab.IgG
C0483761|T201|COMP|6833-8|LNC|Cat dander Ab.IgE|Cat dander Ab.IgE
C0483762|T201|COMP|7184-5|LNC|Cat dander Ab.IgG|Cat dander Ab.IgG
C0483763|T201|COMP|7185-2|LNC|Cat dander basophil bound Ab|Cat dander basophil bound Ab
C0483764|T201|COMP|7186-0|LNC|Cat hair Ab.IgE|Cat hair Ab.IgE
C0483765|T201|COMP|6834-6|LNC|Cat hair+Cat epithelium Ab.IgE|Cat hair+Cat epithelium Ab.IgE
C0483766|T201|COMP|7187-8|LNC|Ictalurus punctatus Ab.IgE|Ictalurus punctatus Ab.IgE
C0483767|T201|COMP|7188-6|LNC|Ictalurus punctatus basophil bound Ab|Ictalurus punctatus basophil bound Ab
C0483768|T201|COMP|7189-4|LNC|Typhaceae sp Ab.IgE|Typhaceae sp Ab.IgE
C0483769|T201|COMP|6835-3|LNC|Brassica oleracea var botrytis Ab.IgE|Brassica oleracea var botrytis Ab.IgE
C0483770|T201|COMP|7190-2|LNC|Brassica oleracea var botrytis Ab.IgG|Brassica oleracea var botrytis Ab.IgG
C0483771|T201|COMP|7191-0|LNC|Brassica oleracea var botrytis basophil bound Ab|Brassica oleracea var botrytis basophil bound Ab
C0483772|T201|COMP|7192-8|LNC|Cedar dust Ab.IgE|Cedar dust Ab.IgE
C0483773|T201|COMP|7193-6|LNC|Juniperus sabinoides Ab.IgG|Juniperus sabinoides Ab.IgG
C0483774|T201|COMP|7194-4|LNC|Juniperus sabinoides basophil bound Ab|Juniperus sabinoides basophil bound Ab
C0483775|T201|COMP|7195-1|LNC|Juniperus virginiana Ab.IgE|Juniperus virginiana Ab.IgE
C0483776|T201|COMP|7196-9|LNC|Tamarix spp Ab.IgE|Tamarix spp Ab.IgE
C0483777|T201|COMP|7197-7|LNC|Apium graveolens Ab.IgG|Apium graveolens Ab.IgG
C0483778|T201|COMP|7198-5|LNC|Apium graveolens basophil bound Ab|Apium graveolens basophil bound Ab
C0483779|T201|COMP|7199-3|LNC|Cephalosporine mold Ab.IgE|Cephalosporine mold Ab.IgE
C0483780|T201|COMP|7200-9|LNC|Chaetomium globosum Ab.IgE|Chaetomium globosum Ab.IgE
C0483781|T201|COMP|7201-7|LNC|Cheese American Ab.IgE|Cheese American Ab.IgE
C0483782|T201|COMP|7202-5|LNC|Cheese American Ab.IgG|Cheese American Ab.IgG
C0483783|T201|COMP|7203-3|LNC|Cheese blue Ab.IgE|Cheese blue Ab.IgE
C0483784|T201|COMP|7204-1|LNC|Cheese cheddar type Ab.IgG|Cheese cheddar type Ab.IgG
C0483785|T201|COMP|7205-8|LNC|Cheese cheddar type basophil bound Ab|Cheese cheddar type basophil bound Ab
C0483786|T201|COMP|7206-6|LNC|Cheese cottage Ab.IgE|Cheese cottage Ab.IgE
C0483787|T201|COMP|7207-4|LNC|Cheese cottage Ab.IgG|Cheese cottage Ab.IgG
C0483788|T201|COMP|7208-2|LNC|Cheese cream basophil bound Ab|Cheese cream basophil bound Ab
C0483789|T201|COMP|7209-0|LNC|Cheese mozzarella Ab.IgE|Cheese mozzarella Ab.IgE
C0483790|T201|COMP|7210-8|LNC|Cheese mozzarella Ab.IgG|Cheese mozzarella Ab.IgG
C0483791|T201|COMP|7211-6|LNC|Cheese mozzarella basophil bound Ab|Cheese mozzarella basophil bound Ab
C0483792|T201|COMP|7212-4|LNC|Cheese parmesan Ab.IgE|Cheese parmesan Ab.IgE
C0483793|T201|COMP|7213-2|LNC|Cheese parmesan basophil bound Ab|Cheese parmesan basophil bound Ab
C0483794|T201|COMP|7214-0|LNC|Cheese roquefort Ab.IgE|Cheese roquefort Ab.IgE
C0483795|T201|COMP|7215-7|LNC|Cheese swiss Ab.IgE|Cheese swiss Ab.IgE
C0483796|T201|COMP|7216-5|LNC|Cheese swiss Ab.IgG|Cheese swiss Ab.IgG
C0483797|T201|COMP|6719-9|LNC|Prunus avium Ab.IgE|Prunus avium Ab.IgE
C0483798|T201|COMP|7217-3|LNC|Prunus avium Ab.IgG|Prunus avium Ab.IgG
C0483799|T201|COMP|7218-1|LNC|Prunus avium basophil bound Ab|Prunus avium basophil bound Ab
C0483800|T201|COMP|6259-6|LNC|Castanea sativa Ab.IgE|Castanea sativa Ab.IgE
C0483801|T201|COMP|7220-7|LNC|Aesculus hippocastanum Ab.IgE|Aesculus hippocastanum Ab.IgE
C0483802|T201|COMP|7221-5|LNC|Chewing gum Ab.IgE|Chewing gum Ab.IgE
C0483803|T201|COMP|7222-3|LNC|Chicken Ab.IgG|Chicken Ab.IgG
C0483804|T201|COMP|7223-1|LNC|Chicken basophil bound Ab|Chicken basophil bound Ab
C0483805|T201|COMP|7224-9|LNC|Chicken feather Ab.IgG|Chicken feather Ab.IgG
C0483806|T201|COMP|6836-1|LNC|Chicken serum proteins Ab.IgE|Chicken serum proteins Ab.IgE
C0483807|T201|COMP|7225-6|LNC|Cichorium intybus Ab.IgE|Cichorium intybus Ab.IgE
C0483808|T201|COMP|7226-4|LNC|Sapium sebiferum Ab.IgE|Sapium sebiferum Ab.IgE
C0483809|T201|COMP|6720-7|LNC|Chocolate Ab.IgG|Chocolate Ab.IgG
C0483810|T201|COMP|7227-2|LNC|Chocolate basophil bound Ab|Chocolate basophil bound Ab
C0483811|T201|COMP|7228-0|LNC|Chymodiactin Ab.IgE|Chymodiactin Ab.IgE
C0483812|T201|COMP|6837-9|LNC|Cinnamomum spp Ab.IgE|Cinnamomum spp Ab.IgE
C0483813|T201|COMP|7229-8|LNC|Cinnamomum spp Ab.IgG|Cinnamomum spp Ab.IgG
C0483814|T201|COMP|7230-6|LNC|Cladosporium herbarum Ab.IgG|Cladosporium herbarum Ab.IgG
C0483815|T201|COMP|7231-4|LNC|Cladosporium herbarum basophil bound Ab|Cladosporium herbarum basophil bound Ab
C0483816|T201|COMP|7232-2|LNC|Ruditapes spp Ab.IgG|Ruditapes spp Ab.IgG
C0483817|T201|COMP|7233-0|LNC|Ruditapes spp basophil bound Ab|Ruditapes spp basophil bound Ab
C0483818|T201|COMP|7234-8|LNC|Syzygium aromaticum Ab.IgE|Syzygium aromaticum Ab.IgE
C0483819|T201|COMP|7235-5|LNC|Syzygium aromaticum Ab.IgG|Syzygium aromaticum Ab.IgG
C0483820|T201|COMP|7236-3|LNC|Clover Ab.IgE|Clover Ab.IgE
C0483821|T201|COMP|6838-7|LNC|Cockatiel droppings Ab.IgE|Cockatiel droppings Ab.IgE
C0483822|T201|COMP|7237-1|LNC|Cockatoo Ab.IgE|Cockatoo Ab.IgE
C0483823|T201|COMP|7238-9|LNC|Xanthium commune Ab.IgG|Xanthium commune Ab.IgG
C0483824|T201|COMP|7239-7|LNC|Xanthium commune basophil bound Ab|Xanthium commune basophil bound Ab
C0483825|T201|COMP|7240-5|LNC|Cocos nucifera Ab.IgG|Cocos nucifera Ab.IgG
C0483826|T201|COMP|7241-3|LNC|Cocos nucifera basophil bound Ab|Cocos nucifera basophil bound Ab
C0483827|T201|COMP|6721-5|LNC|Gadus morhua Ab.IgG|Gadus morhua Ab.IgG
C0483828|T201|COMP|7242-1|LNC|Gadus morhua basophil bound Ab|Gadus morhua basophil bound Ab
C0483829|T201|COMP|6722-3|LNC|Coffea spp Ab.IgG|Coffea spp Ab.IgG
C0483830|T201|COMP|7243-9|LNC|Coffee bean Ab.IgE|Coffee bean Ab.IgE
C0483831|T201|COMP|7244-7|LNC|Cola Ab.IgE|Cola Ab.IgE
C0483832|T201|COMP|7245-4|LNC|Cola Ab.IgG|Cola Ab.IgG
C0483833|T201|COMP|7246-2|LNC|Cola nut basophil bound Ab|Cola nut basophil bound Ab
C0483834|T201|COMP|6723-1|LNC|Zea mays Ab.IgG|Zea mays Ab.IgG
C0483835|T201|COMP|7247-0|LNC|Zea mays basophil bound Ab|Zea mays basophil bound Ab
C0483836|T201|COMP|7248-8|LNC|Zea mays pollen Ab.IgE|Zea mays pollen Ab.IgE
C0483837|T201|COMP|7249-6|LNC|Cornish hen basophil bound Ab|Cornish hen basophil bound Ab
C0483838|T201|COMP|7250-4|LNC|Cotton gin dust Ab.IgE|Cotton gin dust Ab.IgE
C0483839|T201|COMP|7251-2|LNC|Cotton linters Ab.IgE|Cotton linters Ab.IgE
C0483840|T201|COMP|7252-0|LNC|Cotton linters basophil bound Ab|Cotton linters basophil bound Ab
C0483841|T201|COMP|7253-8|LNC|Cottonseed Ab.IgG|Cottonseed Ab.IgG
C0483844|T201|COMP|7255-3|LNC|Populus fremontii Ab.IgE|Populus fremontii Ab.IgE
C0483845|T201|COMP|7257-9|LNC|Cow epithelium Ab.IgE|Cow epithelium Ab.IgE
C0483846|T201|COMP|7258-7|LNC|Cow milk Ab.IgE|Cow milk Ab.IgE
C0483847|T201|COMP|6729-8|LNC|Cow milk Ab.IgG|Cow milk Ab.IgG
C0483848|T201|COMP|7259-5|LNC|Cow milk basophil bound Ab|Cow milk basophil bound Ab
C0483849|T201|COMP|7260-3|LNC|Cancer pagurus Ab.IgG|Cancer pagurus Ab.IgG
C0483850|T201|COMP|7261-1|LNC|Cancer pagurus basophil bound Ab|Cancer pagurus basophil bound Ab
C0483851|T201|COMP|7262-9|LNC|Vaccinium oxycoccos Ab.IgE|Vaccinium oxycoccos Ab.IgE
C0483852|T201|COMP|7263-7|LNC|Vaccinium oxycoccos Ab.IgG|Vaccinium oxycoccos Ab.IgG
C0483853|T201|COMP|7264-5|LNC|Vaccinium oxycoccos basophil bound Ab|Vaccinium oxycoccos basophil bound Ab
C0483854|T201|COMP|7265-2|LNC|Astacus astacus Ab.IgE|Astacus astacus Ab.IgE
C0483855|T201|COMP|7266-0|LNC|Cricket Ab.IgE|Cricket Ab.IgE
C0483856|T201|COMP|7267-8|LNC|Cryptococcus terreus Ab.IgE|Cryptococcus terreus Ab.IgE
C0483857|T201|COMP|6839-5|LNC|Cryptostroma corticale Ab.IgE|Cryptostroma corticale Ab.IgE
C0483858|T201|COMP|6724-9|LNC|Cucumis sativus Ab.IgE|Cucumis sativus Ab.IgE
C0483859|T201|COMP|7268-6|LNC|Cucumis sativus Ab.IgG|Cucumis sativus Ab.IgG
C0483860|T201|COMP|7269-4|LNC|Cucumis sativus basophil bound Ab|Cucumis sativus basophil bound Ab
C0483861|T201|COMP|7270-2|LNC|Curry Ab.IgE|Curry Ab.IgE
C0483862|T201|COMP|7271-0|LNC|Curvularia sp Ab.IgE|Curvularia sp Ab.IgE
C0483863|T201|COMP|7272-8|LNC|Taxodium distichum Ab.IgE|Taxodium distichum Ab.IgE
C0483864|T201|COMP|7273-6|LNC|Dahlia sp Ab.IgE|Dahlia sp Ab.IgE
C0483865|T201|COMP|7274-4|LNC|Bellis perennis Ab.IgE|Bellis perennis Ab.IgE
C0483866|T201|COMP|7275-1|LNC|Phoenix canariensis pollen Ab.IgE|Phoenix canariensis pollen Ab.IgE
C0483867|T201|COMP|7276-9|LNC|Dermatophagoides farinae Ab.IgG|Dermatophagoides farinae Ab.IgG
C0483868|T201|COMP|7277-7|LNC|Dermatophagoides farinae basophil bound Ab|Dermatophagoides farinae basophil bound Ab
C0483869|T201|COMP|7278-5|LNC|Dermatophagoides pteronyssinus Ab.IgG|Dermatophagoides pteronyssinus Ab.IgG
C0483870|T201|COMP|7279-3|LNC|Dermatophagoides pteronyssinus basophil bound Ab|Dermatophagoides pteronyssinus basophil bound Ab
C0483871|T201|COMP|7280-1|LNC|Anethum graveolens Ab.IgE|Anethum graveolens Ab.IgE
C0483872|T201|COMP|7281-9|LNC|Anethum graveolens Ab.IgG|Anethum graveolens Ab.IgG
C0483873|T201|COMP|7282-7|LNC|Discase Ab.IgE|Discase Ab.IgE
C0483874|T201|COMP|6738-9|LNC|Rumex crispus Ab.IgE|Rumex crispus Ab.IgE
C0483875|T201|COMP|7283-5|LNC|Rumex crispus basophil bound Ab|Rumex crispus basophil bound Ab
C0483876|T201|COMP|7284-3|LNC|Dog dander Ab.IgG|Dog dander Ab.IgG
C0483877|T201|COMP|7285-0|LNC|Dog epithelium Ab.IgG|Dog epithelium Ab.IgG
C0483878|T201|COMP|7286-8|LNC|Dog epithelium basophil bound Ab|Dog epithelium basophil bound Ab
C0483879|T201|COMP|7287-6|LNC|Anthemis cotula Ab.IgE|Anthemis cotula Ab.IgE
C0483880|T201|COMP|7288-4|LNC|Dogwood pollen Ab.IgE|Dogwood pollen Ab.IgE
C0483881|T201|COMP|7289-2|LNC|Duck feather Ab.IgG|Duck feather Ab.IgG
C0483882|T201|COMP|6725-6|LNC|Egg white Ab.IgG|Egg white Ab.IgG
C0483883|T201|COMP|7290-0|LNC|Egg white basophil bound Ab|Egg white basophil bound Ab
C0483884|T201|COMP|7291-8|LNC|Egg whole Ab.IgE|Egg whole Ab.IgE
C0483885|T201|COMP|7292-6|LNC|Egg whole Ab.IgG|Egg whole Ab.IgG
C0483886|T201|COMP|7293-4|LNC|Egg whole basophil bound Ab|Egg whole basophil bound Ab
C0483887|T201|COMP|7294-2|LNC|Egg yolk Ab.IgG|Egg yolk Ab.IgG
C0483888|T201|COMP|7295-9|LNC|Egg yolk basophil bound Ab|Egg yolk basophil bound Ab
C0483889|T201|COMP|7296-7|LNC|Solanum melongena Ab.IgE|Solanum melongena Ab.IgE
C0483890|T201|COMP|7297-5|LNC|Solanum melongena Ab.IgG|Solanum melongena Ab.IgG
C0483891|T201|COMP|7484-9|LNC|Iva xanthifolia Ab.IgE|Iva xanthifolia Ab.IgE
C0483892|T201|COMP|7485-6|LNC|Iva xanthifolia Ab.IgG|Iva xanthifolia Ab.IgG
C0483893|T201|COMP|7298-3|LNC|Sambucus nigra Ab.IgG|Sambucus nigra Ab.IgG
C0483894|T201|COMP|6108-5|LNC|Sambucus nigra Ab.IgE|Sambucus nigra Ab.IgE
C0483895|T201|COMP|6109-3|LNC|Ulmus americana Ab.IgE|Ulmus americana Ab.IgE
C0483896|T201|COMP|7301-5|LNC|Ulmus americana basophil bound Ab|Ulmus americana basophil bound Ab
C0483898|T201|COMP|7302-3|LNC|Ulmus pumila Ab.IgE|Ulmus pumila Ab.IgE
C0483899|T201|COMP|7304-9|LNC|Cichorium endivia Ab.IgE|Cichorium endivia Ab.IgE
C0483900|T201|COMP|7305-6|LNC|Cichorium endivia Ab.IgG|Cichorium endivia Ab.IgG
C0483901|T201|COMP|6111-9|LNC|Epicoccum purpurascens Ab.IgE|Epicoccum purpurascens Ab.IgE
C0483902|T201|COMP|7307-2|LNC|Epidermophyton floccosum Ab.IgE|Epidermophyton floccosum Ab.IgE
C0483903|T201|COMP|7308-0|LNC|Esterase Ab.IgE|Esterase Ab.IgE
C0483904|T201|COMP|7309-8|LNC|Ficus benjamina Ab.IgE|Ficus benjamina Ab.IgE
C0483905|T201|COMP|7310-6|LNC|Pseudotsuga taxifolia Ab.IgE|Pseudotsuga taxifolia Ab.IgE
C0483906|T201|COMP|7491-4|LNC|Firebush mexican Ab.IgE|Firebush mexican Ab.IgE
C0483907|T201|COMP|7311-4|LNC|Fish Ab.IgE|Fish Ab.IgE
C0483908|T201|COMP|7312-2|LNC|Linum usitatissimum Ab.IgE|Linum usitatissimum Ab.IgE
C0483909|T201|COMP|7313-0|LNC|Ctenocephalides sp Ab.IgE|Ctenocephalides sp Ab.IgE
C0483910|T201|COMP|7314-8|LNC|Ctenocephalides sp Ab.IgG|Ctenocephalides sp Ab.IgG
C0483911|T201|COMP|7315-5|LNC|Ctenocephalides sp basophil bound Ab|Ctenocephalides sp basophil bound Ab
C0483912|T201|COMP|7316-3|LNC|Flounder Ab.IgE|Flounder Ab.IgE
C0483913|T201|COMP|7317-1|LNC|Flounder Ab.IgG|Flounder Ab.IgG
C0483914|T201|COMP|7318-9|LNC|Flounder basophil bound Ab|Flounder basophil bound Ab
C0483915|T201|COMP|7319-7|LNC|Chrysops flavidus (whole body) Ab.IgE|Chrysops flavidus (whole body) Ab.IgE
C0483916|T201|COMP|7320-5|LNC|Tabanus spp Ab.IgG|Tabanus spp Ab.IgG
C0483917|T201|COMP|7321-3|LNC|Musca domestica basophil bound Ab|Musca domestica basophil bound Ab
C0483918|T201|COMP|7322-1|LNC|Formaldehyde basophil bound Ab|Formaldehyde basophil bound Ab
C0483919|T201|COMP|7323-9|LNC|Fruit Ab.IgE|Fruit Ab.IgE
C0483920|T201|COMP|7324-7|LNC|Fusarium culmorum Ab.IgG|Fusarium culmorum Ab.IgG
C0483921|T201|COMP|7325-4|LNC|Fusarium moniliforme Ab.IgG|Fusarium moniliforme Ab.IgG
C0483923|T201|COMP|7327-0|LNC|Fusarium solani Ab.IgE|Fusarium solani Ab.IgE
C0483924|T201|COMP|7328-8|LNC|Fusarium solani Ab.IgG|Fusarium solani Ab.IgG
C0483925|T201|COMP|7326-2|LNC|Fusarium oxysporum Ab.IgE|Fusarium oxysporum Ab.IgE
C0483926|T201|COMP|7330-4|LNC|Allium sativum Ab.IgG|Allium sativum Ab.IgG
C0483927|T201|COMP|7331-2|LNC|Allium sativum basophil bound Ab|Allium sativum basophil bound Ab
C0483928|T201|COMP|7332-0|LNC|Gelatin Ab.IgE|Gelatin Ab.IgE
C0483929|T201|COMP|7333-8|LNC|Geotrichum candidum Ab.IgE|Geotrichum candidum Ab.IgE
C0483930|T201|COMP|6840-3|LNC|Gerbil Ab.IgE|Gerbil Ab.IgE
C0483931|T201|COMP|7334-6|LNC|Gerbil epithelium Ab.IgE|Gerbil epithelium Ab.IgE
C0483932|T201|COMP|7335-3|LNC|Zingiber officinale Ab.IgE|Zingiber officinale Ab.IgE
C0483933|T201|COMP|7336-1|LNC|Zingiber officinale Ab.IgG|Zingiber officinale Ab.IgG
C0483934|T201|COMP|7337-9|LNC|Gladiolus sp Ab.IgE|Gladiolus sp Ab.IgE
C0483935|T201|COMP|7338-7|LNC|Gluten Ab.IgG|Gluten Ab.IgG
C0483936|T201|COMP|7339-5|LNC|Gnat whole body Ab.IgE|Gnat whole body Ab.IgE
C0483937|T201|COMP|7340-3|LNC|Goat milk Ab.IgE|Goat milk Ab.IgE
C0483938|T201|COMP|7341-1|LNC|Goat milk Ab.IgG|Goat milk Ab.IgG
C0483939|T201|COMP|7342-9|LNC|Solidago virgaurea Ab.IgG|Solidago virgaurea Ab.IgG
C0483940|T201|COMP|7343-7|LNC|Solidago virgaurea basophil bound Ab|Solidago virgaurea basophil bound Ab
C0483941|T201|COMP|7344-5|LNC|Goose feather Ab.IgG|Goose feather Ab.IgG
C0483942|T201|COMP|7345-2|LNC|Grain Ab.IgE|Grain Ab.IgE
C0483943|T201|COMP|7346-0|LNC|Grain dust Ab.IgE|Grain dust Ab.IgE
C0483944|T201|COMP|7347-8|LNC|Grain mill dust Ab.IgE|Grain mill dust Ab.IgE
C0483945|T201|COMP|6841-1|LNC|Vitis vinifera Ab.IgE|Vitis vinifera Ab.IgE
C0483946|T201|COMP|7348-6|LNC|Vitis vinifera Ab.IgG|Vitis vinifera Ab.IgG
C0483947|T201|COMP|7349-4|LNC|Grape raisin basophil bound Ab|Grape raisin basophil bound Ab
C0483948|T201|COMP|7350-2|LNC|Citrus paradisis Ab.IgG|Citrus paradisis Ab.IgG
C0483949|T201|COMP|7351-0|LNC|Citrus paradisis basophil bound Ab|Citrus paradisis basophil bound Ab
C0483950|T201|COMP|7111-8|LNC|Paspalum notatum basophil bound Ab|Paspalum notatum basophil bound Ab
C0483951|T201|COMP|6228-1|LNC|Agrostis stolonifera Ab.IgE|Agrostis stolonifera Ab.IgE
C0483952|T201|COMP|7353-6|LNC|Cynodon dactylon Ab.IgG|Cynodon dactylon Ab.IgG
C0483953|T201|COMP|7354-4|LNC|Cynodon dactylon basophil bound Ab|Cynodon dactylon basophil bound Ab
C0483954|T201|COMP|7355-1|LNC|Poa annua Ab.IgE|Poa annua Ab.IgE
C0483955|T201|COMP|7356-9|LNC|Poa compressa Ab.IgE|Poa compressa Ab.IgE
C0483957|T201|COMP|7358-5|LNC|Poa pratensis basophil bound Ab|Poa pratensis basophil bound Ab
C0483958|T201|COMP|6726-4|LNC|Arrhenatherum elatius Ab.IgE|Arrhenatherum elatius Ab.IgE
C0483959|T201|COMP|7359-3|LNC|Festuca elatior basophil bound Ab|Festuca elatior basophil bound Ab
C0483960|T201|COMP|7360-1|LNC|Bouteloua gracilis Ab.IgE|Bouteloua gracilis Ab.IgE
C0483961|T201|COMP|7361-9|LNC|Sorghum halepense basophil bound Ab|Sorghum halepense basophil bound Ab
C0483962|T201|COMP|7362-7|LNC|Grass koehlers Ab.IgE|Grass koehlers Ab.IgE
C0483963|T201|COMP|6169-7|LNC|Festuca elatior Ab.IgE|Festuca elatior Ab.IgE
C0483964|T201|COMP|7364-3|LNC|Festuca elatior Ab.IgG|Festuca elatior Ab.IgG
C0483965|T201|COMP|7365-0|LNC|Dactylis glomerata Ab.IgG|Dactylis glomerata Ab.IgG
C0483966|T201|COMP|7366-8|LNC|Dactylis glomerata basophil bound Ab|Dactylis glomerata basophil bound Ab
C0483967|T201|COMP|7367-6|LNC|Agropyron repens Ab.IgE|Agropyron repens Ab.IgE
C0483968|T201|COMP|7368-4|LNC|Agrostis stolonifera basophil bound Ab|Agrostis stolonifera basophil bound Ab
C0483969|T201|COMP|7369-2|LNC|Lolium perenne Ab.IgE|Lolium perenne Ab.IgE
C0483972|T201|COMP|7370-0|LNC|Lolium perenne Ab.IgG|Lolium perenne Ab.IgG
C0483973|T201|COMP|7374-2|LNC|Lolium perenne basophil bound Ab|Lolium perenne basophil bound Ab
C0483974|T201|COMP|7375-9|LNC|Grass sorghum Ab.IgE|Grass sorghum Ab.IgE
C0483975|T201|COMP|7376-7|LNC|Sorghum sudanense Ab.IgE|Sorghum sudanense Ab.IgE
C0483976|T201|COMP|7377-5|LNC|Anthoxanthum odoratum basophil bound Ab|Anthoxanthum odoratum basophil bound Ab
C0483977|T201|COMP|7378-3|LNC|Grass tall oat Ab.IgE|Grass tall oat Ab.IgE
C0483978|T201|COMP|7379-1|LNC|Grass wheat Ab.IgG|Grass wheat Ab.IgG
C0483979|T201|COMP|7380-9|LNC|Grayfish Ab.IgE|Grayfish Ab.IgE
C0483980|T201|COMP|7381-7|LNC|Sarcobatus vermiculatus Ab.IgE|Sarcobatus vermiculatus Ab.IgE
C0483981|T201|COMP|7382-5|LNC|Gum arabic Ab.IgE|Gum arabic Ab.IgE
C0483982|T201|COMP|7383-3|LNC|Celtis occidentalis Ab.IgE|Celtis occidentalis Ab.IgE
C0483983|T201|COMP|7384-1|LNC|Melanogrammus aeglefinus Ab.IgE|Melanogrammus aeglefinus Ab.IgE
C0483984|T201|COMP|7385-8|LNC|Melanogrammus aeglefinus Ab.IgG|Melanogrammus aeglefinus Ab.IgG
C0483985|T201|COMP|6842-9|LNC|Hippoglossus hippoglossus Ab.IgE|Hippoglossus hippoglossus Ab.IgE
C0483986|T201|COMP|7386-6|LNC|Hippoglossus hippoglossus Ab.IgG|Hippoglossus hippoglossus Ab.IgG
C0483987|T201|COMP|7387-4|LNC|Hippoglossus hippoglossus basophil bound Ab|Hippoglossus hippoglossus basophil bound Ab
C0483988|T201|COMP|7388-2|LNC|Ham basophil bound Ab|Ham basophil bound Ab
C0483989|T201|COMP|7389-0|LNC|Hay Ab.IgE|Hay Ab.IgE
C0483990|T201|COMP|7391-6|LNC|Corylus avellana Ab.IgG|Corylus avellana Ab.IgG
C0483991|T201|COMP|7392-4|LNC|Corylus avellana basophil bound Ab|Corylus avellana basophil bound Ab
C0483992|T201|COMP|7393-2|LNC|Helminthosporium interseminatum Ab.IgE|Helminthosporium interseminatum Ab.IgE
C0483993|T201|COMP|7394-0|LNC|Helminthosporium maydis Ab.IgE|Helminthosporium maydis Ab.IgE
C0483994|T201|COMP|7395-7|LNC|Helminthosporium sp Ab.IgE|Helminthosporium sp Ab.IgE
C0483995|T201|COMP|7396-5|LNC|Helminthosporium sp Ab.IgG|Helminthosporium sp Ab.IgG
C0483996|T201|COMP|7397-3|LNC|Tsuga canadensis Ab.IgE|Tsuga canadensis Ab.IgE
C0483997|T201|COMP|7398-1|LNC|Hemp Ab.IgE|Hemp Ab.IgE
C0483998|T201|COMP|7399-9|LNC|Hemp fiber Ab.IgE|Hemp fiber Ab.IgE
C0483999|T201|COMP|7400-5|LNC|Amaranthus tuberculatus Ab.IgE|Amaranthus tuberculatus Ab.IgE
C0484000|T201|COMP|7401-3|LNC|Clupea harengus Ab.IgG|Clupea harengus Ab.IgG
C0484002|T201|COMP|7403-9|LNC|Hickory basophil bound Ab|Hickory basophil bound Ab
C0484003|T201|COMP|7404-7|LNC|Carya ovata Ab.IgE|Carya ovata Ab.IgE
C0484004|T201|COMP|7405-4|LNC|Carya laciniosa Ab.IgE|Carya laciniosa Ab.IgE
C0484005|T201|COMP|6209-1|LNC|Carya illinoinensis tree Ab.IgE|Carya illinoinensis tree Ab.IgE
C0484006|T201|COMP|7407-0|LNC|Carya tomentosa Ab.IgE|Carya tomentosa Ab.IgE
C0484007|T201|COMP|7408-8|LNC|Histamine extract basophil bound Ab|Histamine extract basophil bound Ab
C0484008|T201|COMP|7412-0|LNC|Honey Ab.IgE|Honey Ab.IgE
C0484009|T201|COMP|7411-2|LNC|Honey Ab.IgG|Honey Ab.IgG
C0484010|T201|COMP|7413-8|LNC|Honeysuckle Ab.IgE|Honeysuckle Ab.IgE
C0484011|T201|COMP|7414-6|LNC|Humulus lupus Ab.IgG|Humulus lupus Ab.IgG
C0484012|T201|COMP|7415-3|LNC|Cladosporium sphaerospermum Ab.IgE|Cladosporium sphaerospermum Ab.IgE
C0484013|T201|COMP|7416-1|LNC|Carpinus betulus Ab.IgE|Carpinus betulus Ab.IgE
C0484014|T201|COMP|7417-9|LNC|Dolichovespula maculata Ab.IgG|Dolichovespula maculata Ab.IgG
C0484015|T201|COMP|6739-7|LNC|Dolichovespula arenaria Ab.IgG|Dolichovespula arenaria Ab.IgG
C0484016|T201|COMP|7418-7|LNC|Horse dander basophil bound Ab|Horse dander basophil bound Ab
C0484017|T201|COMP|7419-5|LNC|Horse epithelium Ab.IgE|Horse epithelium Ab.IgE
C0484018|T201|COMP|7420-3|LNC|Armoracia rusticana Ab.IgE|Armoracia rusticana Ab.IgE
C0484019|T201|COMP|7421-1|LNC|House dust AP Ab.IgE|House dust AP Ab.IgE
C0484020|T201|COMP|7422-9|LNC|House dust AP Ab.IgG|House dust AP Ab.IgG
C0484021|T201|COMP|7423-7|LNC|House dust basophil bound Ab|House dust basophil bound Ab
C0484022|T201|COMP|7424-5|LNC|House dust Greer Ab.IgG|House dust Greer Ab.IgG
C0484023|T201|COMP|9444-1|LNC|House dust Hausstaub Ab.IgE|House dust Hausstaub Ab.IgE
C0484024|T201|COMP|7425-2|LNC|House dust Hollister Stier Ab.IgE|House dust Hollister Stier Ab.IgE
C0484025|T201|COMP|7426-0|LNC|House dust Hollister Stier Ab.IgG|House dust Hollister Stier Ab.IgG
C0484026|T201|COMP|9828-5|LNC|House dust Greer Ab.IgE|House dust Greer Ab.IgE
C0484027|T201|COMP|7427-8|LNC|Hymenopterase Ab.IgE|Hymenopterase Ab.IgE
C0484028|T201|COMP|7428-6|LNC|Allenrolfea occidentalis Ab.IgE|Allenrolfea occidentalis Ab.IgE
C0484029|T201|COMP|7429-4|LNC|Hexamethylene diisocyanate (HDI) Ab.IgE|Hexamethylene diisocyanate (HDI) Ab.IgE
C0484030|T201|COMP|7430-2|LNC|Diphenylmethane diisocyanate (MDI) Ab.IgE|Diphenylmethane diisocyanate (MDI) Ab.IgE
C0484031|T201|COMP|7431-0|LNC|Toluene diisocyanate (TDI) Ab.IgE|Toluene diisocyanate (TDI) Ab.IgE
C0484032|T201|COMP|7432-8|LNC|Juniper Ab.IgE|Juniper Ab.IgE
C0484033|T201|COMP|7433-6|LNC|Juniper basophil bound Ab|Juniper basophil bound Ab
C0484034|T201|COMP|7434-4|LNC|Juniperus pinchotii Ab.IgE|Juniperus pinchotii Ab.IgE
C0484035|T201|COMP|7435-1|LNC|Juniperus occidentalis Ab.IgE|Juniperus occidentalis Ab.IgE
C0484036|T201|COMP|7436-9|LNC|Chorchorus capsularis Ab.IgE|Chorchorus capsularis Ab.IgE
C0484037|T201|COMP|7437-7|LNC|Kapok Ab.IgE|Kapok Ab.IgE
C0484038|T201|COMP|7438-5|LNC|Kapok basophil bound Ab|Kapok basophil bound Ab
C0484039|T201|COMP|7439-3|LNC|Karaya gum Ab.IgE|Karaya gum Ab.IgE
C0484040|T201|COMP|7440-1|LNC|Actinidia chinensis Ab.IgG|Actinidia chinensis Ab.IgG
C0484041|T201|COMP|7441-9|LNC|Actinidia chinensis basophil bound Ab|Actinidia chinensis basophil bound Ab
C0484042|T201|COMP|7442-7|LNC|Kochia scoparia Ab.IgA|Kochia scoparia Ab.IgA
C0484043|T201|COMP|7443-5|LNC|Kochia scoparia Ab.IgE|Kochia scoparia Ab.IgE
C0484043|T201|COMP|7163-9|LNC|Kochia scoparia Ab.IgE|Kochia scoparia Ab.IgE
C0484043|T201|COMP|6118-4|LNC|Kochia scoparia Ab.IgE|Kochia scoparia Ab.IgE
C0484044|T201|COMP|7444-3|LNC|Lactalbumin Ab.IgG|Lactalbumin Ab.IgG
C0484045|T201|COMP|7445-0|LNC|Lactalbumin alpha Ab.IgE|Lactalbumin alpha Ab.IgE
C0484046|T201|COMP|7446-8|LNC|Lactalbumin basophil bound Ab|Lactalbumin basophil bound Ab
C0484047|T201|COMP|7447-6|LNC|Lactoglobulin Ab.IgG|Lactoglobulin Ab.IgG
C0484048|T201|COMP|7448-4|LNC|Lamb Ab.IgG|Lamb Ab.IgG
C0484049|T201|COMP|7449-2|LNC|Lamb basophil bound Ab|Lamb basophil bound Ab
C0484050|T201|COMP|7450-0|LNC|Chenopodium album basophil bound Ab|Chenopodium album basophil bound Ab
C0484051|T201|COMP|7451-8|LNC|Latex ALK basophil bound Ab|Latex ALK basophil bound Ab
C0484052|T201|COMP|7452-6|LNC|Latex Bencard basophil bound Ab|Latex Bencard basophil bound Ab
C0484053|T201|COMP|6728-0|LNC|Latex glove extract Ab.IgE|Latex glove extract Ab.IgE
C0484054|T201|COMP|6845-2|LNC|Latex glove extract ammoniated Ab.IgE|Latex glove extract ammoniated Ab.IgE
C0484055|T201|COMP|6846-0|LNC|Latex glove extract buffered Ab.IgE|Latex glove extract buffered Ab.IgE
C0484056|T201|COMP|7453-4|LNC|Latex Greer basophil bound Ab|Latex Greer basophil bound Ab
C0484057|T201|COMP|7454-2|LNC|Latex Stallerg basophil bound Ab|Latex Stallerg basophil bound Ab
C0484058|T201|COMP|7455-9|LNC|Citrus limon Ab.IgG|Citrus limon Ab.IgG
C0484059|T201|COMP|7456-7|LNC|Citrus limon basophil bound Ab|Citrus limon basophil bound Ab
C0484060|T201|COMP|6239-8|LNC|Atriplex lentiformis Ab.IgE|Atriplex lentiformis Ab.IgE
C0484061|T201|COMP|7458-3|LNC|Lens esculenta Ab.IgE|Lens esculenta Ab.IgE
C0484062|T201|COMP|7459-1|LNC|Lens esculenta Ab.IgG|Lens esculenta Ab.IgG
C0484063|T201|COMP|7460-9|LNC|Lactuca sativa Ab.IgG|Lactuca sativa Ab.IgG
C0484064|T201|COMP|7461-7|LNC|Lactuca sativa basophil bound Ab|Lactuca sativa basophil bound Ab
C0484065|T201|COMP|7462-5|LNC|Glycyrrhiza lepidota Ab.IgE|Glycyrrhiza lepidota Ab.IgE
C0484066|T201|COMP|7463-3|LNC|Lilium longiflorum Ab.IgE|Lilium longiflorum Ab.IgE
C0484067|T201|COMP|7464-1|LNC|Citrus aurantifolia Ab.IgE|Citrus aurantifolia Ab.IgE
C0484068|T201|COMP|7465-8|LNC|Citrus aurantifolia Ab.IgG|Citrus aurantifolia Ab.IgG
C0484069|T201|COMP|7466-6|LNC|Linen Ab.IgE|Linen Ab.IgE
C0484070|T201|COMP|7467-4|LNC|Lipolase Ab.IgE|Lipolase Ab.IgE
C0484071|T201|COMP|7468-2|LNC|Liver Ab.IgE|Liver Ab.IgE
C0484072|T201|COMP|7469-0|LNC|Liver calf Ab.IgE|Liver calf Ab.IgE
C0484073|T201|COMP|7470-8|LNC|Llama fur Ab.IgE|Llama fur Ab.IgE
C0484074|T201|COMP|7471-6|LNC|Homarus gammarus Ab.IgG|Homarus gammarus Ab.IgG
C0484075|T201|COMP|7472-4|LNC|Locust tree Ab.IgE|Locust tree Ab.IgE
C0484076|T201|COMP|7473-2|LNC|Robinia pseudoacacia Ab.IgE|Robinia pseudoacacia Ab.IgE
C0484077|T201|COMP|7474-0|LNC|Scomber scombrus Ab.IgE|Scomber scombrus Ab.IgE
C0484078|T201|COMP|7475-7|LNC|Scomber scombrus basophil bound Ab|Scomber scombrus basophil bound Ab
C0484079|T201|COMP|7476-5|LNC|Malt Ab.IgG|Malt Ab.IgG
C0484080|T201|COMP|7477-3|LNC|Mangifera indica pollen Ab.IgE|Mangifera indica pollen Ab.IgE
C0484081|T201|COMP|7478-1|LNC|Acer macrophyllum Ab.IgE|Acer macrophyllum Ab.IgE
C0484082|T201|COMP|7479-9|LNC|Acer rubrum Ab.IgE|Acer rubrum Ab.IgE
C0484083|T201|COMP|7480-7|LNC|Acer rubrum basophil bound Ab|Acer rubrum basophil bound Ab
C0484084|T201|COMP|7481-5|LNC|Maple red+Silver Ab.IgE|Maple red+Silver Ab.IgE
C0484085|T201|COMP|7482-3|LNC|Maple sugar Ab.IgE|Maple sugar Ab.IgE
C0484086|T201|COMP|7483-1|LNC|Maple syrup Ab.IgE|Maple syrup Ab.IgE
C0484087|T201|COMP|7486-4|LNC|Mattress dust Ab.IgE|Mattress dust Ab.IgE
C0484088|T201|COMP|7487-2|LNC|Mayfly Ab.IgE|Mayfly Ab.IgE
C0484089|T201|COMP|7488-0|LNC|Mayfly basophil bound Ab|Mayfly basophil bound Ab
C0484090|T201|COMP|7489-8|LNC|Melaleuca leucadendron basophil bound Ab|Melaleuca leucadendron basophil bound Ab
C0484091|T201|COMP|57880-7|LNC|Cucumis melo spp Ab.IgG|Cucumis melo spp Ab.IgG
C0484092|T201|COMP|6847-8|LNC|Chenopodium ambrosioides Ab.IgE|Chenopodium ambrosioides Ab.IgE
C0484093|T201|COMP|7492-2|LNC|Multiple inhalant allergen Ab.IgE|Multiple inhalant allergen Ab.IgE
C0484094|T201|COMP|7493-0|LNC|Milk evaporated Ab.IgE|Milk evaporated Ab.IgE
C0484095|T201|COMP|7494-8|LNC|Panicum milliaceum Ab.IgG|Panicum milliaceum Ab.IgG
C0484096|T201|COMP|7495-5|LNC|Mite dust Ab.IgE|Mite dust Ab.IgE
C0484097|T201|COMP|7496-3|LNC|Cheese mold type Ab.IgG|Cheese mold type Ab.IgG
C0484098|T201|COMP|7497-1|LNC|Cheese mold type basophil bound Ab|Cheese mold type basophil bound Ab
C0484099|T201|COMP|7498-9|LNC|Chrysonilia sitophila Ab.IgE|Chrysonilia sitophila Ab.IgE
C0484100|T201|COMP|7499-7|LNC|Monkey epithelium Ab.IgE|Monkey epithelium Ab.IgE
C0484101|T201|COMP|7500-2|LNC|Aedes communis basophil bound Ab|Aedes communis basophil bound Ab
C0484102|T201|COMP|7501-0|LNC|Tillandsia usneoides Ab.IgE|Tillandsia usneoides Ab.IgE
C0484103|T201|COMP|7502-8|LNC|Moth Ab.IgE|Moth Ab.IgE
C0484104|T201|COMP|7503-6|LNC|Moth basophil bound Ab|Moth basophil bound Ab
C0484105|T201|COMP|7504-4|LNC|Mouse hair Ab.IgE|Mouse hair Ab.IgE
C0484106|T201|COMP|7505-1|LNC|Mouse multi Ab.IgE|Mouse multi Ab.IgE
C0484107|T201|COMP|7506-9|LNC|Mucor plumbeus Ab.IgE|Mucor plumbeus Ab.IgE
C0484108|T201|COMP|7507-7|LNC|Mucor racemosus Ab.IgG|Mucor racemosus Ab.IgG
C0484109|T201|COMP|7508-5|LNC|Mucor racemosus basophil bound Ab|Mucor racemosus basophil bound Ab
C0484110|T201|COMP|7509-3|LNC|Mucor sp Ab.IgG|Mucor sp Ab.IgG
C0484111|T201|COMP|7510-1|LNC|Artemisia vulgaris basophil bound Ab|Artemisia vulgaris basophil bound Ab
C0484112|T201|COMP|7511-9|LNC|Artemisia douglasiana Ab.IgE|Artemisia douglasiana Ab.IgE
C0484113|T201|COMP|7512-7|LNC|Morus alba Ab.IgE|Morus alba Ab.IgE
C0484113|T201|COMP|6281-0|LNC|Morus alba Ab.IgE|Morus alba Ab.IgE
C0484113|T201|COMP|17291-6|LNC|Morus alba Ab.IgE|Morus alba Ab.IgE
C0484114|T201|COMP|7513-5|LNC|Morus alba Ab.IgG|Morus alba Ab.IgG
C0484115|T201|COMP|7514-3|LNC|Morus rubra Ab.IgE|Morus rubra Ab.IgE
C0484116|T201|COMP|6848-6|LNC|Agaricus hortensis Ab.IgE|Agaricus hortensis Ab.IgE
C0484117|T201|COMP|7515-0|LNC|Agaricus hortensis Ab.IgG|Agaricus hortensis Ab.IgG
C0484118|T201|COMP|7516-8|LNC|Agaricus hortensis basophil bound Ab|Agaricus hortensis basophil bound Ab
C0484119|T201|COMP|7517-6|LNC|Pleurotus ostreatus Ab.IgE|Pleurotus ostreatus Ab.IgE
C0484120|T201|COMP|57884-9|LNC|Cucumis melo spp Ab.IgE|Cucumis melo spp Ab.IgE
C0484121|T201|COMP|7519-2|LNC|Mytilus edulis Ab.IgG|Mytilus edulis Ab.IgG
C0484122|T201|COMP|7520-0|LNC|Mytilus edulis basophil bound Ab|Mytilus edulis basophil bound Ab
C0484123|T201|COMP|7521-8|LNC|Mustard Ab.IgG|Mustard Ab.IgG
C0484124|T201|COMP|7522-6|LNC|Mycogone sp Ab.IgE|Mycogone sp Ab.IgE
C0484125|T201|COMP|7523-4|LNC|Prunus persica var nucipersica Ab.IgE|Prunus persica var nucipersica Ab.IgE
C0484126|T201|COMP|7524-2|LNC|Prunus persica var nucipersica Ab.IgG|Prunus persica var nucipersica Ab.IgG
C0484127|T201|COMP|7525-9|LNC|Nigrospora oryzae Ab.IgE|Nigrospora oryzae Ab.IgE
C0484128|T201|COMP|7526-7|LNC|Nigrospora sphaerica Ab.IgE|Nigrospora sphaerica Ab.IgE
C0484129|T201|COMP|7527-5|LNC|Nutmeg Ab.IgG|Nutmeg Ab.IgG
C0484130|T201|COMP|7528-3|LNC|Quercus velutina Ab.IgE|Quercus velutina Ab.IgE
C0484131|T201|COMP|7529-1|LNC|Quercus kelloggii Ab.IgE|Quercus kelloggii Ab.IgE
C0484132|T201|COMP|7530-9|LNC|Quercus gambelii Ab.IgE|Quercus gambelii Ab.IgE
C0484133|T201|COMP|7531-7|LNC|Chenopodium botrys Ab.IgE|Chenopodium botrys Ab.IgE
C0484134|T201|COMP|7532-5|LNC|Quercus agrifolia Ab.IgE|Quercus agrifolia Ab.IgE
C0484135|T201|COMP|7533-3|LNC|Quercus wislizeni Ab.IgE|Quercus wislizeni Ab.IgE
C0484136|T201|COMP|7534-1|LNC|Quercus rubra Ab.IgE|Quercus rubra Ab.IgE
C0484137|T201|COMP|7535-8|LNC|Quercus lobata Ab.IgE|Quercus lobata Ab.IgE
C0484138|T201|COMP|6189-5|LNC|Quercus alba Ab.IgE|Quercus alba Ab.IgE
C0484139|T201|COMP|7536-6|LNC|Quercus alba Ab.IgG|Quercus alba Ab.IgG
C0484140|T201|COMP|7537-4|LNC|Quercus alba basophil bound Ab|Quercus alba basophil bound Ab
C0484141|T201|COMP|7538-2|LNC|Avena sativa Ab.IgG|Avena sativa Ab.IgG
C0484142|T201|COMP|7539-0|LNC|Avena sativa basophil bound Ab|Avena sativa basophil bound Ab
C0484144|T201|COMP|6190-3|LNC|Avena sativa Ab.IgE|Avena sativa Ab.IgE
C0484145|T201|COMP|7542-4|LNC|Trisetum paniceum Ab.IgE|Trisetum paniceum Ab.IgE
C0484146|T201|COMP|7543-2|LNC|Oidiodendrum spp Ab.IgE|Oidiodendrum spp Ab.IgE
C0484147|T201|COMP|7544-0|LNC|Abelmoschus esculentus Ab.IgE|Abelmoschus esculentus Ab.IgE
C0484148|T201|COMP|7545-7|LNC|Olive Ab.IgE|Olive Ab.IgE
C0484149|T201|COMP|7546-5|LNC|Olea europaea Ab.IgG|Olea europaea Ab.IgG
C0484150|T201|COMP|7547-3|LNC|Olive green Ab.IgE|Olive green Ab.IgE
C0484151|T201|COMP|7548-1|LNC|Allium cepa Ab.IgG|Allium cepa Ab.IgG
C0484152|T201|COMP|7549-9|LNC|Allium cepa basophil bound Ab|Allium cepa basophil bound Ab
C0484153|T201|COMP|6730-6|LNC|Citrus sinensis Ab.IgG|Citrus sinensis Ab.IgG
C0484154|T201|COMP|7550-7|LNC|Citrus sinensis basophil bound Ab|Citrus sinensis basophil bound Ab
C0484155|T201|COMP|7551-5|LNC|Citrus sinensis tree Ab.IgE|Citrus sinensis tree Ab.IgE
C0484156|T201|COMP|7552-3|LNC|Origanum vulgare Ab.IgE|Origanum vulgare Ab.IgE
C0484157|T201|COMP|7553-1|LNC|Origanum vulgare Ab.IgG|Origanum vulgare Ab.IgG
C0484158|T201|COMP|7554-9|LNC|Origanum vulgare basophil bound Ab|Origanum vulgare basophil bound Ab
C0484159|T201|COMP|7555-6|LNC|Iris germanica var florentina Ab.IgE|Iris germanica var florentina Ab.IgE
C0484160|T201|COMP|7556-4|LNC|Ovalbumin Ab.IgE|Ovalbumin Ab.IgE
C0484161|T201|COMP|7557-2|LNC|Ovomucoid Ab.IgE|Ovomucoid Ab.IgE
C0484162|T201|COMP|7558-0|LNC|Ostrea edulis Ab.IgE|Ostrea edulis Ab.IgE
C0484163|T201|COMP|7559-8|LNC|Ostrea edulis Ab.IgG|Ostrea edulis Ab.IgG
C0484164|T201|COMP|7560-6|LNC|Ostrea edulis basophil bound Ab|Ostrea edulis basophil bound Ab
C0484165|T201|COMP|6060-8|LNC|Amaranthus palmeri Ab.IgE|Amaranthus palmeri Ab.IgE
C0484166|T201|COMP|6850-2|LNC|Carica papaya Ab.IgE|Carica papaya Ab.IgE
C0484167|T201|COMP|7562-2|LNC|Paper Ab.IgE|Paper Ab.IgE
C0484168|T201|COMP|7563-0|LNC|Capsicum annuum Ab.IgE|Capsicum annuum Ab.IgE
C0484169|T201|COMP|7564-8|LNC|Parakeet droppings Ab.IgE|Parakeet droppings Ab.IgE
C0484170|T201|COMP|7565-5|LNC|Parakeet feather Ab.IgE|Parakeet feather Ab.IgE
C0484171|T201|COMP|7566-3|LNC|Parakeet serum Ab.IgE|Parakeet serum Ab.IgE
C0484172|T201|COMP|7567-1|LNC|Parrot serum Ab.IgE|Parrot serum Ab.IgE
C0484173|T201|COMP|7568-9|LNC|Petroselinum crispum Ab.IgG|Petroselinum crispum Ab.IgG
C0484174|T201|COMP|7569-7|LNC|Pastinaca sativa Ab.IgE|Pastinaca sativa Ab.IgE
C0484175|T201|COMP|7570-5|LNC|Pisum sativum Ab.IgG|Pisum sativum Ab.IgG
C0484176|T201|COMP|7571-3|LNC|Vigna sinensis Ab.IgE|Vigna sinensis Ab.IgE
C0484177|T201|COMP|7572-1|LNC|Vigna sinensis Ab.IgG|Vigna sinensis Ab.IgG
C0484178|T201|COMP|7573-9|LNC|Cicer arietinus Ab.IgE|Cicer arietinus Ab.IgE
C0484179|T201|COMP|7574-7|LNC|Pisum sativum basophil bound Ab|Pisum sativum basophil bound Ab
C0484180|T201|COMP|7575-4|LNC|Prunus persica Ab.IgG|Prunus persica Ab.IgG
C0484181|T201|COMP|7576-2|LNC|Prunus persica basophil bound Ab|Prunus persica basophil bound Ab
C0484182|T201|COMP|6732-2|LNC|Arachis hypogaea Ab.IgG|Arachis hypogaea Ab.IgG
C0484183|T201|COMP|7577-0|LNC|Arachis hypogaea basophil bound Ab|Arachis hypogaea basophil bound Ab
C0484184|T201|COMP|7578-8|LNC|Pyrus communis Ab.IgG|Pyrus communis Ab.IgG
C0484185|T201|COMP|7579-6|LNC|Pyrus communis pollen Ab.IgE|Pyrus communis pollen Ab.IgE
C0484186|T201|COMP|7580-4|LNC|Carya illinoinensis nut Ab.IgG|Carya illinoinensis nut Ab.IgG
C0484187|T201|COMP|7402-1|LNC|Carya illinoinensis nut basophil bound Ab|Carya illinoinensis nut basophil bound Ab
C0484188|T201|COMP|6851-0|LNC|Penicillin G Ab.IgE|Penicillin G Ab.IgE
C0484189|T201|COMP|7583-8|LNC|Penicillium sp Ab.IgG|Penicillium sp Ab.IgG
C0484190|T201|COMP|7584-6|LNC|Penicillium notatum Ab.IgG|Penicillium notatum Ab.IgG
C0484191|T201|COMP|7585-3|LNC|Penicillium notatum basophil bound Ab|Penicillium notatum basophil bound Ab
C0484192|T201|COMP|7586-1|LNC|Pepper bell Ab.IgE|Pepper bell Ab.IgE
C0484193|T201|COMP|7587-9|LNC|Pepper bell Ab.IgG|Pepper bell Ab.IgG
C0484194|T201|COMP|7588-7|LNC|Piper nigrum Ab.IgG|Piper nigrum Ab.IgG
C0484195|T201|COMP|7589-5|LNC|Piper nigrum basophil bound Ab|Piper nigrum basophil bound Ab
C0484196|T201|COMP|7590-3|LNC|Pepper cayenne Ab.IgG|Pepper cayenne Ab.IgG
C0484197|T201|COMP|7591-1|LNC|Capsicum frutescens Ab.IgE|Capsicum frutescens Ab.IgE
C0484198|T201|COMP|7592-9|LNC|Capsicum frutescens Ab.IgG|Capsicum frutescens Ab.IgG
C0484199|T201|COMP|7593-7|LNC|Capsicum frutescens basophil bound Ab|Capsicum frutescens basophil bound Ab
C0484200|T201|COMP|6852-8|LNC|Pepper green Ab.IgE|Pepper green Ab.IgE
C0484201|T201|COMP|7594-5|LNC|Pepper green Ab.IgG|Pepper green Ab.IgG
C0484202|T201|COMP|7595-2|LNC|Pepper red basophil bound Ab|Pepper red basophil bound Ab
C0484203|T201|COMP|7596-0|LNC|Pepper white Ab.IgE|Pepper white Ab.IgE
C0484204|T201|COMP|7597-8|LNC|Pepper white Ab.IgG|Pepper white Ab.IgG
C0484205|T201|COMP|7598-6|LNC|Perca spp Ab.IgG|Perca spp Ab.IgG
C0484206|T201|COMP|7599-4|LNC|Phadiatop Ab.IgE|Phadiatop Ab.IgE
C0484207|T201|COMP|7600-0|LNC|Phospholipase Ab.IgE|Phospholipase Ab.IgE
C0484208|T201|COMP|7601-8|LNC|Phthalic anhydride Ab.IgE|Phthalic anhydride Ab.IgE
C0484209|T201|COMP|7602-6|LNC|Salicornia spp Ab.IgE|Salicornia spp Ab.IgE
C0484210|T201|COMP|7603-4|LNC|Pigeon droppings Ab.IgG|Pigeon droppings Ab.IgG
C0484211|T201|COMP|6733-0|LNC|Pigeon serum Ab|Pigeon serum Ab
C0484212|T201|COMP|7604-2|LNC|Pigweed common Ab.IgE|Pigweed common Ab.IgE
C0484213|T201|COMP|7605-9|LNC|Pigweed Ab.IgG|Pigweed Ab.IgG
C0484214|T201|COMP|7606-7|LNC|Pigweed basophil bound Ab|Pigweed basophil bound Ab
C0484215|T201|COMP|7761-0|LNC|Stizostedion vitreum Ab.IgE|Stizostedion vitreum Ab.IgE
C0484216|T201|COMP|6282-8|LNC|Pinus strobus Ab.IgE|Pinus strobus Ab.IgE
C0484217|T201|COMP|7608-3|LNC|Pinus taeda Ab.IgE|Pinus taeda Ab.IgE
C0484219|T201|COMP|7610-9|LNC|Pinus ponderosa Ab.IgE|Pinus ponderosa Ab.IgE
C0484220|T201|COMP|7611-7|LNC|Pinus monticola Ab.IgE|Pinus monticola Ab.IgE
C0484221|T201|COMP|7612-5|LNC|Ananas comosus Ab.IgG|Ananas comosus Ab.IgG
C0484222|T201|COMP|7613-3|LNC|Pistacia vera Ab.IgE|Pistacia vera Ab.IgE
C0484223|T201|COMP|7614-1|LNC|Pitosporium basophil bound Ab|Pitosporium basophil bound Ab
C0484224|T201|COMP|7615-8|LNC|Plantain Ab.IgE|Plantain Ab.IgE
C0484225|T201|COMP|7616-6|LNC|Plantago lanceolata basophil bound Ab|Plantago lanceolata basophil bound Ab
C0484226|T201|COMP|6853-6|LNC|Prunus domestica Ab.IgE|Prunus domestica Ab.IgE
C0484227|T201|COMP|7617-4|LNC|Prunus domestica Ab.IgG|Prunus domestica Ab.IgG
C0484228|T201|COMP|7618-2|LNC|Prunus domestica pollen Ab.IgE|Prunus domestica pollen Ab.IgE
C0484229|T201|COMP|7619-0|LNC|Poison ivy Ab.IgE|Poison ivy Ab.IgE
C0484230|T201|COMP|7254-6|LNC|Populus nigra Ab.IgE|Populus nigra Ab.IgE
C0484231|T201|COMP|7621-6|LNC|Poplar sp Ab.IgE|Poplar sp Ab.IgE
C0484232|T201|COMP|7622-4|LNC|Populus alba basophil bound Ab|Populus alba basophil bound Ab
C0484233|T201|COMP|7623-2|LNC|Papaver somniferum Ab.IgE|Papaver somniferum Ab.IgE
C0484234|T201|COMP|6734-8|LNC|Pork Ab.IgG|Pork Ab.IgG
C0484235|T201|COMP|7624-0|LNC|Pork basophil bound Ab|Pork basophil bound Ab
C0484237|T201|COMP|7626-5|LNC|Solanum tuberosum basophil bound Ab|Solanum tuberosum basophil bound Ab
C0484238|T201|COMP|7627-3|LNC|Ipomoea batatas Ab.IgE|Ipomoea batatas Ab.IgE
C0484239|T201|COMP|7628-1|LNC|Ipomoea batatas Ab.IgG|Ipomoea batatas Ab.IgG
C0484240|T201|COMP|7629-9|LNC|Ipomoea batatas basophil bound Ab|Ipomoea batatas basophil bound Ab
C0484241|T201|COMP|7625-7|LNC|Solanum tuberosum Ab.IgG|Solanum tuberosum Ab.IgG
C0484242|T201|COMP|7631-5|LNC|Iva axillaris Ab.IgE|Iva axillaris Ab.IgE
C0484243|T201|COMP|7632-3|LNC|Ligustrum vulgare Ab.IgE|Ligustrum vulgare Ab.IgE
C0484244|T201|COMP|7633-1|LNC|Ligustrum vulgare Ab.IgG|Ligustrum vulgare Ab.IgG
C0484245|T201|COMP|7634-9|LNC|Prune Ab.IgE|Prune Ab.IgE
C0484246|T201|COMP|7635-6|LNC|Psyllium seed Ab.IgE|Psyllium seed Ab.IgE
C0484247|T201|COMP|7636-4|LNC|Pullularia pullulans Ab.IgE|Pullularia pullulans Ab.IgE
C0484248|T201|COMP|7637-2|LNC|Pullularia sp Ab.IgE|Pullularia sp Ab.IgE
C0484249|T201|COMP|7638-0|LNC|Pullularia sp Ab.IgG|Pullularia sp Ab.IgG
C0484250|T201|COMP|6854-4|LNC|Cucurbita pepo Ab.IgE|Cucurbita pepo Ab.IgE
C0484251|T201|COMP|7639-8|LNC|Chrysanthemum cinerariifolium Ab.IgE|Chrysanthemum cinerariifolium Ab.IgE
C0484252|T201|COMP|7640-6|LNC|Chrysanthemum cinerariifolium basophil bound Ab|Chrysanthemum cinerariifolium basophil bound Ab
C0484253|T201|COMP|7641-4|LNC|Chrysothamnus nauseosus Ab.IgE|Chrysothamnus nauseosus Ab.IgE
C0484254|T201|COMP|7642-2|LNC|Rabbit meat Ab.IgE|Rabbit meat Ab.IgE
C0484255|T201|COMP|7643-0|LNC|Raphanus sativus Ab.IgE|Raphanus sativus Ab.IgE
C0484256|T201|COMP|7644-8|LNC|Raphanus sativus Ab.IgG|Raphanus sativus Ab.IgG
C0484257|T201|COMP|7645-5|LNC|Ambrosia ambrosioides Ab.IgE|Ambrosia ambrosioides Ab.IgE
C0484258|T201|COMP|7646-3|LNC|Ambrosia elatior Ab.IgG|Ambrosia elatior Ab.IgG
C0484259|T201|COMP|7647-1|LNC|Ambrosia dumosa Ab.IgE|Ambrosia dumosa Ab.IgE
C0484260|T201|COMP|7648-9|LNC|Franseria acanthicarpa basophil bound Ab|Franseria acanthicarpa basophil bound Ab
C0484261|T201|COMP|7649-7|LNC|Ambrosia trifida basophil bound Ab|Ambrosia trifida basophil bound Ab
C0484262|T201|COMP|7650-5|LNC|Ambrosia elatior Ab.IgE|Ambrosia elatior Ab.IgE
C0484262|T201|COMP|6086-3|LNC|Ambrosia elatior Ab.IgE|Ambrosia elatior Ab.IgE
C0484263|T201|COMP|7651-3|LNC|Ambrosia elatior Ab.IgG|Ambrosia elatior Ab.IgG
C0484264|T201|COMP|7652-1|LNC|Ambrosia elatior basophil bound Ab|Ambrosia elatior basophil bound Ab
C0484265|T201|COMP|7653-9|LNC|Ambrosia elatior+Ambrosia trifida Ab.IgG|Ambrosia elatior+Ambrosia trifida Ab.IgG
C0484266|T201|COMP|7654-7|LNC|Ambrosia confertiflora Ab.IgE|Ambrosia confertiflora Ab.IgE
C0484267|T201|COMP|7655-4|LNC|Ambrosia bidentata Ab.IgE|Ambrosia bidentata Ab.IgE
C0484268|T201|COMP|7656-2|LNC|Rubus idaeus Ab.IgE|Rubus idaeus Ab.IgE
C0484269|T201|COMP|7657-0|LNC|Rubus idaeus Ab.IgG|Rubus idaeus Ab.IgG
C0484270|T201|COMP|7658-8|LNC|Rubus idaeus basophil bound Ab|Rubus idaeus basophil bound Ab
C0484271|T201|COMP|6934-4|LNC|RAST class|RAST class
C0484272|T201|COMP|7659-6|LNC|Rat hair Ab.IgE|Rat hair Ab.IgE
C0484273|T201|COMP|7660-4|LNC|Rat muliialgro Ab.IgE|Rat muliialgro Ab.IgE
C0484274|T201|COMP|7661-2|LNC|Snapper red Ab.IgE|Snapper red Ab.IgE
C0484275|T201|COMP|7662-0|LNC|Snapper red Ab.IgG|Snapper red Ab.IgG
C0484276|T201|COMP|7663-8|LNC|Sequoia spp dust Ab.IgE|Sequoia spp dust Ab.IgE
C0484277|T201|COMP|7664-6|LNC|Sequoia spp Ab.IgE|Sequoia spp Ab.IgE
C0484278|T201|COMP|6855-1|LNC|Phragmites communis Ab.IgE|Phragmites communis Ab.IgE
C0484279|T201|COMP|7665-3|LNC|Rhodotorula spp Ab.IgE|Rhodotorula spp Ab.IgE
C0484280|T201|COMP|7667-9|LNC|Rheum spp Ab.IgE|Rheum spp Ab.IgE
C0484281|T201|COMP|7668-7|LNC|Oryza sativa Ab.IgG|Oryza sativa Ab.IgG
C0484282|T201|COMP|7669-5|LNC|Oryza sativa basophil bound Ab|Oryza sativa basophil bound Ab
C0484283|T201|COMP|7777-6|LNC|Zizania spp Ab.IgE|Zizania spp Ab.IgE
C0484284|T201|COMP|7670-3|LNC|Rubber tree brazilian Ab.IgE|Rubber tree brazilian Ab.IgE
C0484285|T201|COMP|7672-9|LNC|Puccinia graminis triticu Ab.IgE|Puccinia graminis triticu Ab.IgE
C0484286|T201|COMP|7673-7|LNC|Secale cereale basophil bound Ab|Secale cereale basophil bound Ab
C0484288|T201|COMP|7675-2|LNC|Secale cereale Ab.IgG|Secale cereale Ab.IgG
C0484289|T201|COMP|7676-0|LNC|Carthamus tinctorius Ab.IgE|Carthamus tinctorius Ab.IgE
C0484290|T201|COMP|7677-8|LNC|Carthamus tinctorius Ab.IgG|Carthamus tinctorius Ab.IgG
C0484291|T201|COMP|7678-6|LNC|Salvia officinalis Ab.IgE|Salvia officinalis Ab.IgE
C0484292|T201|COMP|7680-2|LNC|Salvia officinalis Ab.IgG|Salvia officinalis Ab.IgG
C0484294|T201|COMP|7682-8|LNC|Artemisia tridentata Ab.IgG|Artemisia tridentata Ab.IgG
C0484295|T201|COMP|7683-6|LNC|Artemisia californica Ab.IgE|Artemisia californica Ab.IgE
C0484296|T201|COMP|7681-0|LNC|Artemisia tridentata Ab.IgE|Artemisia tridentata Ab.IgE
C0484297|T201|COMP|7685-1|LNC|Salmo salar Ab.IgG|Salmo salar Ab.IgG
C0484298|T201|COMP|7686-9|LNC|Saltbush Ab.IgE|Saltbush Ab.IgE
C0484299|T201|COMP|7687-7|LNC|Saltbush annual Ab.IgE|Saltbush annual Ab.IgE
C0484300|T201|COMP|7688-5|LNC|Sardine Ab.IgG|Sardine Ab.IgG
C0484301|T201|COMP|7689-3|LNC|Savinase Ab.IgE|Savinase Ab.IgE
C0484302|T201|COMP|7690-1|LNC|Atriplex polycarpa Ab.IgE|Atriplex polycarpa Ab.IgE
C0484303|T201|COMP|7691-9|LNC|Pecten spp Ab.IgE|Pecten spp Ab.IgE
C0484304|T201|COMP|7692-7|LNC|Pecten spp Ab.IgG|Pecten spp Ab.IgG
C0484305|T201|COMP|7693-5|LNC|Schistosoma sp Ab.IgE|Schistosoma sp Ab.IgE
C0484306|T201|COMP|7694-3|LNC|Scorpion Ab.IgE|Scorpion Ab.IgE
C0484307|T201|COMP|7695-0|LNC|Cytisus scoparius Ab.IgE|Cytisus scoparius Ab.IgE
C0484308|T201|COMP|7696-8|LNC|Sesamum indicum Ab.IgG|Sesamum indicum Ab.IgG
C0484309|T201|COMP|7697-6|LNC|Sesamum indicum basophil bound Ab|Sesamum indicum basophil bound Ab
C0484310|T201|COMP|7698-4|LNC|Sheep epithelium basophil bound Ab|Sheep epithelium basophil bound Ab
C0484311|T201|COMP|7699-2|LNC|Rumex acetosella basophil bound Ab|Rumex acetosella basophil bound Ab
C0484312|T201|COMP|7700-8|LNC|Pandalus borealis Ab.IgG|Pandalus borealis Ab.IgG
C0484313|T201|COMP|7701-6|LNC|Pandalus borealis basophil bound Ab|Pandalus borealis basophil bound Ab
C0484314|T201|COMP|9676-8|LNC|Silicone Ab.IgE|Silicone Ab.IgE
C0484315|T201|COMP|7702-4|LNC|Smelt Ab.IgE|Smelt Ab.IgE
C0484316|T201|COMP|7704-0|LNC|Ustilago cynodontis Ab.IgE|Ustilago cynodontis Ab.IgE
C0484317|T201|COMP|7703-2|LNC|Ustilago maydis Ab.IgE|Ustilago maydis Ab.IgE
C0484318|T201|COMP|7705-7|LNC|Sphacelotheca cruenta Ab.IgE|Sphacelotheca cruenta Ab.IgE
C0484319|T201|COMP|7706-5|LNC|Sphacelotheca cruenta Ab.IgG|Sphacelotheca cruenta Ab.IgG
C0484320|T201|COMP|7707-3|LNC|Ustilago avenae Ab.IgE|Ustilago avenae Ab.IgE
C0484321|T201|COMP|7708-1|LNC|Ustilago tritici Ab.IgE|Ustilago tritici Ab.IgE
C0484322|T201|COMP|7709-9|LNC|Solea solea Ab.IgE|Solea solea Ab.IgE
C0484323|T201|COMP|7710-7|LNC|Solea solea Ab.IgG|Solea solea Ab.IgG
C0484324|T201|COMP|6856-9|LNC|Spinacia oleracea Ab.IgE|Spinacia oleracea Ab.IgE
C0484325|T201|COMP|7711-5|LNC|Spinacia oleracea Ab.IgG|Spinacia oleracea Ab.IgG
C0484326|T201|COMP|7712-3|LNC|Spondylocladium atrovirens Ab.IgE|Spondylocladium atrovirens Ab.IgE
C0484327|T201|COMP|6857-7|LNC|Picea excelsa Ab.IgE|Picea excelsa Ab.IgE
C0484328|T201|COMP|7713-1|LNC|Squash Ab.IgE|Squash Ab.IgE
C0484329|T201|COMP|7714-9|LNC|Squash summer Ab.IgE|Squash summer Ab.IgE
C0484330|T201|COMP|7715-6|LNC|Squash summer Ab.IgG|Squash summer Ab.IgG
C0484331|T201|COMP|7716-4|LNC|Squash yellow Ab.IgE|Squash yellow Ab.IgE
C0484332|T201|COMP|7717-2|LNC|Squash yellow Ab.IgG|Squash yellow Ab.IgG
C0484333|T201|COMP|7718-0|LNC|Squash zucchini Ab.IgE|Squash zucchini Ab.IgE
C0484334|T201|COMP|6858-5|LNC|Loligo sp Ab.IgE|Loligo sp Ab.IgE
C0484335|T201|COMP|7719-8|LNC|Staphylococcus aureus Ab.IgE|Staphylococcus aureus Ab.IgE
C0484336|T201|COMP|7720-6|LNC|Stemphylium solani Ab.IgE|Stemphylium solani Ab.IgE
C0484337|T201|COMP|7721-4|LNC|Fragaria vesca Ab.IgG|Fragaria vesca Ab.IgG
C0484338|T201|COMP|7722-2|LNC|Fragaria vesca basophil bound Ab|Fragaria vesca basophil bound Ab
C0484339|T201|COMP|7723-0|LNC|Saccharum officinarum Ab.IgE|Saccharum officinarum Ab.IgE
C0484340|T201|COMP|7724-8|LNC|Saccharum officinarum Ab.IgG|Saccharum officinarum Ab.IgG
C0484341|T201|COMP|7725-5|LNC|Helianthus annuus Ab.IgG|Helianthus annuus Ab.IgG
C0484342|T201|COMP|7726-3|LNC|Helianthus annuus pollen Ab.IgE|Helianthus annuus pollen Ab.IgE
C0484343|T201|COMP|7727-1|LNC|Helianthus annuus seed basophil bound Ab|Helianthus annuus seed basophil bound Ab
C0484344|T201|COMP|7409-6|LNC|Swine basophil bound Ab|Swine basophil bound Ab
C0484345|T201|COMP|7410-4|LNC|Swine epithelium Ab.IgG|Swine epithelium Ab.IgG
C0484346|T201|COMP|7728-9|LNC|Xiphias gladius Ab.IgE|Xiphias gladius Ab.IgE
C0484347|T201|COMP|7729-7|LNC|Xiphias gladius Ab.IgG|Xiphias gladius Ab.IgG
C0484348|T201|COMP|6263-8|LNC|Platanus occidentalis Ab.IgE|Platanus occidentalis Ab.IgE
C0484349|T201|COMP|7731-3|LNC|Citrus reticulata Ab.IgE|Citrus reticulata Ab.IgE
C0484350|T201|COMP|7732-1|LNC|Citrus reticulata Ab.IgG|Citrus reticulata Ab.IgG
C0484351|T201|COMP|7733-9|LNC|Manihot esculenta crantz Ab.IgE|Manihot esculenta crantz Ab.IgE
C0484352|T201|COMP|7734-7|LNC|Manihot esculenta crantz Ab.IgG|Manihot esculenta crantz Ab.IgG
C0484353|T201|COMP|7735-4|LNC|Camellia sinensis Ab.IgG|Camellia sinensis Ab.IgG
C0484354|T201|COMP|7736-2|LNC|Termamyl Ab.IgE|Termamyl Ab.IgE
C0484355|T201|COMP|7671-1|LNC|Salsola kali Ab.IgG|Salsola kali Ab.IgG
C0484356|T201|COMP|7737-0|LNC|Thymus vulgaris Ab.IgE|Thymus vulgaris Ab.IgE
C0484357|T201|COMP|7738-8|LNC|Phleum pratense basophil bound Ab|Phleum pratense basophil bound Ab
C0484358|T201|COMP|7739-6|LNC|Nicotiana tabacum Ab.IgG|Nicotiana tabacum Ab.IgG
C0484359|T201|COMP|7740-4|LNC|Nicotiana tabacum basophil bound Ab|Nicotiana tabacum basophil bound Ab
C0484360|T201|COMP|7741-2|LNC|Nicotiana tabacum cigarette Ab.IgE|Nicotiana tabacum cigarette Ab.IgE
C0484361|T201|COMP|6859-3|LNC|Nicotiana tabacum Ab.IgE|Nicotiana tabacum Ab.IgE
C0484362|T201|COMP|6736-3|LNC|Lycopersicon lycopersicum Ab.IgG|Lycopersicon lycopersicum Ab.IgG
C0484363|T201|COMP|7742-0|LNC|Lycopersicon lycopersicum basophil bound Ab|Lycopersicon lycopersicum basophil bound Ab
C0484364|T201|COMP|7743-8|LNC|Astragalus spp Ab.IgE|Astragalus spp Ab.IgE
C0484365|T201|COMP|7744-6|LNC|Ailanthus altissima Ab.IgE|Ailanthus altissima Ab.IgE
C0484366|T201|COMP|7745-3|LNC|Trichophyton Ab.IgE|Trichophyton Ab.IgE
C0484367|T201|COMP|6860-1|LNC|Trichophyton rubrum Ab.IgE|Trichophyton rubrum Ab.IgE
C0484368|T201|COMP|7746-1|LNC|Trimellitic anhydride Ab.IgE|Trimellitic anhydride Ab.IgE
C0484369|T201|COMP|7747-9|LNC|Oncorhynchus mykiss Ab.IgG|Oncorhynchus mykiss Ab.IgG
C0484370|T201|COMP|7748-7|LNC|Tryptase Ab.IgE|Tryptase Ab.IgE
C0484371|T201|COMP|7749-5|LNC|Thunnus albacares Ab.IgG|Thunnus albacares Ab.IgG
C0484372|T201|COMP|7750-3|LNC|Thunnus albacares basophil bound Ab|Thunnus albacares basophil bound Ab
C0484373|T201|COMP|7751-1|LNC|Turkey Ab.IgG|Turkey Ab.IgG
C0484374|T201|COMP|7752-9|LNC|Turkey basophil bound Ab|Turkey basophil bound Ab
C0484375|T201|COMP|7753-7|LNC|Turkey feather Ab.IgE|Turkey feather Ab.IgE
C0484376|T201|COMP|7754-5|LNC|Turnip Ab.IgE|Turnip Ab.IgE
C0484377|T201|COMP|7755-2|LNC|Upholstery dust Ab.IgE|Upholstery dust Ab.IgE
C0484378|T201|COMP|7756-0|LNC|Vanilla planifolia Ab.IgE|Vanilla planifolia Ab.IgE
C0484379|T201|COMP|6861-9|LNC|Vanilla planifolia Ab.IgG|Vanilla planifolia Ab.IgG
C0484380|T201|COMP|7757-8|LNC|Veal Ab.IgE|Veal Ab.IgE
C0484381|T201|COMP|7758-6|LNC|Veal basophil bound Ab|Veal basophil bound Ab
C0484382|T201|COMP|7759-4|LNC|Venison Ab.IgE|Venison Ab.IgE
C0484383|T201|COMP|7760-2|LNC|Wall pellitory Ab.IgE|Wall pellitory Ab.IgE
C0484384|T201|COMP|7762-8|LNC|Juglans spp basophil bound Ab|Juglans spp basophil bound Ab
C0484385|T201|COMP|7763-6|LNC|Juglans nigra Ab.IgE|Juglans nigra Ab.IgE
C0484386|T201|COMP|7764-4|LNC|Walnut black western Ab.IgE|Walnut black western Ab.IgE
C0484387|T201|COMP|7765-1|LNC|Juglans regia Ab.IgE|Juglans regia Ab.IgE
C0484388|T201|COMP|7766-9|LNC|Juglans regia pollen Ab.IgE|Juglans regia pollen Ab.IgE
C0484389|T201|COMP|7767-7|LNC|Juglans spp Ab.IgG|Juglans spp Ab.IgG
C0484390|T201|COMP|6731-4|LNC|Polistes spp Ab.IgG|Polistes spp Ab.IgG
C0484391|T201|COMP|6740-5|LNC|Vespula spp Ab.IgE|Vespula spp Ab.IgE
C0484392|T201|COMP|7768-5|LNC|Vespula spp Ab.IgG|Vespula spp Ab.IgG
C0484393|T201|COMP|7769-3|LNC|Trapa natans Ab.IgE|Trapa natans Ab.IgE
C0484394|T201|COMP|7770-1|LNC|Citrullus lanatus Ab.IgE|Citrullus lanatus Ab.IgE
C0484395|T201|COMP|7771-9|LNC|Citrullus lanatus Ab.IgG|Citrullus lanatus Ab.IgG
C0484396|T201|COMP|6737-1|LNC|Triticum aestivum Ab.IgG|Triticum aestivum Ab.IgG
C0484397|T201|COMP|7772-7|LNC|Triticum aestivum basophil bound Ab|Triticum aestivum basophil bound Ab
C0484398|T201|COMP|6277-8|LNC|Triticum aestivum pollen Ab.IgE|Triticum aestivum pollen Ab.IgE
C0484399|T201|COMP|7774-3|LNC|Cow whey Ab.IgE|Cow whey Ab.IgE
C0484400|T201|COMP|7775-0|LNC|Whitefish Ab.IgE|Whitefish Ab.IgE
C0484401|T201|COMP|7776-8|LNC|Whitefish Ab.IgG|Whitefish Ab.IgG
C0484402|T201|COMP|6862-7|LNC|Salix nigra Ab.IgE|Salix nigra Ab.IgE
C0484403|T201|COMP|7778-4|LNC|Salix discolor Ab.IgE|Salix discolor Ab.IgE
C0484404|T201|COMP|7779-2|LNC|Atriplex canescens Ab.IgE|Atriplex canescens Ab.IgE
C0484405|T201|COMP|7780-0|LNC|Ceratoides arborescens Ab.IgE|Ceratoides arborescens Ab.IgE
C0484406|T201|COMP|7781-8|LNC|Artemisia absinthium Ab.IgG|Artemisia absinthium Ab.IgG
C0484407|T201|COMP|7782-6|LNC|Dioscorea batatas Ab.IgE|Dioscorea batatas Ab.IgE
C0484408|T201|COMP|7783-4|LNC|Yeast bakers Ab.IgE|Yeast bakers Ab.IgE
C0484409|T201|COMP|6713-2|LNC|Saccharomyces cerevisiae Ab.IgG|Saccharomyces cerevisiae Ab.IgG
C0484410|T201|COMP|7784-2|LNC|Saccharomyces cerevisiae basophil bound Ab|Saccharomyces cerevisiae basophil bound Ab
C0484411|T201|COMP|6715-7|LNC|Yeast brewer's Ab.IgG|Yeast brewer's Ab.IgG
C0484412|T201|COMP|7785-9|LNC|Yeast brewer's basophil bound Ab|Yeast brewer's basophil bound Ab
C0484413|T201|COMP|7786-7|LNC|Taxus spp Ab.IgE|Taxus spp Ab.IgE
C0484414|T201|COMP|7787-5|LNC|Yogurt Ab.IgE|Yogurt Ab.IgE
C0484415|T201|COMP|7788-3|LNC|Yogurt Ab.IgG|Yogurt Ab.IgG
C0484416|T201|COMP|7789-1|LNC|Acanthocytes|Acanthocytes
C0484417|T201|COMP|10371-3|LNC|Bite cells|Bite cells
C0484418|T201|COMP|10372-1|LNC|Blister cells|Blister cells
C0484419|T201|COMP|7790-9|LNC|Burr cells|Burr cells
C0484421|T201|COMP|7792-5|LNC|Dohle body|Dohle body
C0484422|T201|COMP|9727-9|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0484423|T201|COMP|10327-5|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0484424|T201|COMP|6742-1|LNC|Erythrocyte morphology finding|Erythrocyte morphology finding
C0484425|T201|COMP|6741-3|LNC|Erythrocytes|Erythrocytes
C0484426|T201|COMP|10373-9|LNC|Fragments|Fragments
C0484427|T201|COMP|10374-7|LNC|Helmet cells|Helmet cells
C0484428|T201|COMP|7793-3|LNC|Howell-Jolly bodies|Howell-Jolly bodies
C0484429|T201|COMP|10375-4|LNC|Irregularly contracted cells|Irregularly contracted cells
C0484430|T201|COMP|6690-2|LNC|Leukocytes|Leukocytes
C0484431|T201|COMP|6743-9|LNC|Leukocytes|Leukocytes
C0484432|T201|COMP|6744-7|LNC|Lymphocytes|Lymphocytes
C0484433|T201|COMP|9440-9|LNC|Lymphocytes.IgA/100 lymphocytes|Lymphocytes.IgA/100 lymphocytes
C0484434|T201|COMP|9441-7|LNC|Lymphocytes.IgD/100 lymphocytes|Lymphocytes.IgD/100 lymphocytes
C0484435|T201|COMP|9442-5|LNC|Lymphocytes.IgG/100 lymphocytes|Lymphocytes.IgG/100 lymphocytes
C0484436|T201|COMP|9443-3|LNC|Lymphocytes.IgM/100 lymphocytes|Lymphocytes.IgM/100 lymphocytes
C0484437|T201|COMP|10328-3|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0484438|T201|COMP|10376-2|LNC|Macrocytes.oval|Macrocytes.oval
C0484439|T201|COMP|33252-8|LNC|Monocytes|Monocytes
C0484440|T201|COMP|33251-0|LNC|Monocytes|Monocytes
C0484441|T201|COMP|9305-4|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0484442|T201|COMP|6745-4|LNC|Neutrophils.segmented|Neutrophils.segmented
C0484443|T201|COMP|7794-1|LNC|Normocytic/Normochromic polychromasia|Normocytic/Normochromic polychromasia
C0484444|T201|COMP|7795-8|LNC|Pappenheimer bodies|Pappenheimer bodies
C0484445|T201|COMP|10377-0|LNC|Pencil cells|Pencil cells
C0484446|T201|COMP|7796-6|LNC|Platelet clump|Platelet clump
C0484447|T201|COMP|9317-9|LNC|Platelets|Platelets
C0484448|T201|COMP|10378-8|LNC|Polychromasia|Polychromasia
C0484449|T201|COMP|9306-2|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0484450|T201|COMP|6863-5|LNC|Prolymphocytes|Prolymphocytes
C0484451|T201|COMP|6746-2|LNC|Prolymphocytes/100 leukocytes|Prolymphocytes/100 leukocytes
C0484452|T201|COMP|10379-6|LNC|Erythrocytes.dual population|Erythrocytes.dual population
C0484453|T201|COMP|7797-4|LNC|Rouleaux|Rouleaux
C0484454|T201|COMP|7798-2|LNC|Smudge cells|Smudge cells
C0484455|T201|COMP|10380-4|LNC|Stomatocytes|Stomatocytes
C0484456|T201|COMP|10381-2|LNC|Target cells|Target cells
C0484457|T201|COMP|10382-0|LNC|A,B variant NOS Ag|A,B variant NOS Ag
C0484458|T201|COMP|10383-8|LNC|A,B variant NOS Ag|A,B variant NOS Ag
C0484459|T201|COMP|10384-6|LNC|A,B variant NOS Ag|A,B variant NOS Ag
C0484460|T201|COMP|10385-3|LNC|Albumin concentration given|Albumin concentration given
C0484461|T201|COMP|10386-1|LNC|Albumin given|Albumin given
C0484462|T201|COMP|10387-9|LNC|Autologous erythrocytes given|Autologous erythrocytes given
C0484463|T201|COMP|10388-7|LNC|Autologous whole blood given|Autologous whole blood given
C0484464|T201|COMP|10389-5|LNC|Blood product.other|Blood product.other
C0484465|T201|COMP|10390-3|LNC|Blood product special preparation|Blood product special preparation
C0484466|T201|COMP|10391-1|LNC|Cytomegalovirus immune globulin given|Cytomegalovirus immune globulin given
C0484467|T201|COMP|10392-9|LNC|Cryoprecipitate given|Cryoprecipitate given
C0484468|T201|COMP|967-0|LNC|D little u Ab|D little u Ab
C0484469|T201|COMP|968-8|LNC|D little u Ab|D little u Ab
C0484470|T201|COMP|969-6|LNC|D little u Ab|D little u Ab
C0484471|T201|COMP|10393-7|LNC|Factor IX given|Factor IX given
C0484472|T201|COMP|10394-5|LNC|Factor IX given|Factor IX given
C0484473|T201|COMP|10395-2|LNC|Factor VIII given|Factor VIII given
C0484474|T201|COMP|10396-0|LNC|Factor VIII given|Factor VIII given
C0484475|T201|COMP|10397-8|LNC|Hepatitis B virus immune globulin given|Hepatitis B virus immune globulin given
C0484476|T201|COMP|10401-8|LNC|Immune serum globulin given|Immune serum globulin given
C0484477|T201|COMP|10402-6|LNC|Immune serum globulin given|Immune serum globulin given
C0484478|T201|COMP|10403-4|LNC|Inject immune serum globulin|Inject immune serum globulin
C0484479|T201|COMP|10404-2|LNC|Inject Rh immune globulin|Inject Rh immune globulin
C0484480|T201|COMP|10405-9|LNC|Inject varicella zoster virus immune globulin|Inject varicella zoster virus immune globulin
C0484481|T201|COMP|10409-1|LNC|Pentaspan given|Pentaspan given
C0484482|T201|COMP|10410-9|LNC|Plasma given|Plasma given
C0484483|T201|COMP|10411-7|LNC|Plasma given|Plasma given
C0484484|T201|COMP|10412-5|LNC|Platelets given|Platelets given
C0484485|T201|COMP|10331-7|LNC|Rh|Rh
C0484486|T201|COMP|10413-3|LNC|Rh immune globulin given|Rh immune globulin given
C0484487|T201|COMP|10414-1|LNC|Transfuse albumin|Transfuse albumin
C0484488|T201|COMP|10415-8|LNC|Transfuse blood exchange transfusion|Transfuse blood exchange transfusion
C0484489|T201|COMP|10416-6|LNC|Transfuse blood product.other|Transfuse blood product.other
C0484490|T201|COMP|10417-4|LNC|Transfuse cryoprecipitate|Transfuse cryoprecipitate
C0484491|T201|COMP|10418-2|LNC|Transfuse factor IX|Transfuse factor IX
C0484492|T201|COMP|10419-0|LNC|Transfuse factor VIII|Transfuse factor VIII
C0484493|T201|COMP|10420-8|LNC|Transfuse immune serum globulin|Transfuse immune serum globulin
C0484494|T201|COMP|10421-6|LNC|Transfuse Pentaspan|Transfuse Pentaspan
C0484495|T201|COMP|10422-4|LNC|Transfuse plasma|Transfuse plasma
C0484496|T201|COMP|10423-2|LNC|Transfuse platelets|Transfuse platelets
C0484497|T201|COMP|10424-0|LNC|Transfuse erythrocytes|Transfuse erythrocytes
C0484498|T201|COMP|10425-7|LNC|Transfuse Rh immune globulin|Transfuse Rh immune globulin
C0484499|T201|COMP|10426-5|LNC|Transfuse whole blood|Transfuse whole blood
C0484500|T201|COMP|10427-3|LNC|Transfuse whole blood autologous|Transfuse whole blood autologous
C0484501|T201|COMP|10428-1|LNC|Varicella zoster virus immune globulin given|Varicella zoster virus immune globulin given
C0484502|T201|COMP|10429-9|LNC|AE 1 Ag|AE 1 Ag
C0484503|T201|COMP|10430-7|LNC|AE 3 Ag|AE 3 Ag
C0484504|T201|COMP|10431-5|LNC|B-cell Ag|B-cell Ag
C0484506|T201|COMP|10433-1|LNC|BR-2 Ag|BR-2 Ag
C0484507|T201|COMP|10434-9|LNC|Complement C3 Ag|Complement C3 Ag
C0484508|T201|COMP|10435-6|LNC|C5B-9 Ag|C5B-9 Ag
C0484509|T201|COMP|10436-4|LNC|CD15 Ag|CD15 Ag
C0484510|T201|COMP|10437-2|LNC|CD16 Ag|CD16 Ag
C0484511|T201|COMP|10438-0|LNC|CD20 Ag|CD20 Ag
C0484512|T201|COMP|10439-8|LNC|CD3 Ag|CD3 Ag
C0484513|T201|COMP|10432-3|LNC|CD30 Ag|CD30 Ag
C0484514|T201|COMP|10441-4|LNC|CD34 Ag|CD34 Ag
C0484515|T201|COMP|10442-2|LNC|CD56 Ag|CD56 Ag
C0484516|T201|COMP|10443-0|LNC|CD43.T-Cell monocyte+Myeloid cell Ag|CD43.T-Cell monocyte+Myeloid cell Ag
C0484517|T201|COMP|10444-8|LNC|CD57 Ag|CD57 Ag
C0484518|T201|COMP|10445-5|LNC|CD11c Ag|CD11c Ag
C0484519|T201|COMP|10446-3|LNC|Leukocyte common Ag|Leukocyte common Ag
C0484520|T201|COMP|9680-0|LNC|Cells.CD16+CD57+/100 cells|Cells.CD16+CD57+/100 cells
C0484521|T201|COMP|8101-8|LNC|Cells.CD3+CD8+/100 cells|Cells.CD3+CD8+/100 cells
C0484522|T201|COMP|8102-6|LNC|Cells.CD33/100 cells|Cells.CD33/100 cells
C0484523|T201|COMP|8103-4|LNC|Cells.CD45+CD14+/100 cells|Cells.CD45+CD14+/100 cells
C0484524|T201|COMP|33595-0|LNC|Cells.CD5+CD20+|Cells.CD5+CD20+
C0484525|T201|COMP|8105-9|LNC|Cells.CD5+CD8+/100 cells|Cells.CD5+CD8+/100 cells
C0484526|T201|COMP|8106-7|LNC|Cells.CD1/100 cells|Cells.CD1/100 cells
C0484527|T201|COMP|9554-7|LNC|Cells.CD10|Cells.CD10
C0484528|T201|COMP|8107-5|LNC|Cells.CD10/100 cells|Cells.CD10/100 cells
C0484529|T201|COMP|9840-0|LNC|Cells.CD11+CD20+|Cells.CD11+CD20+
C0484530|T201|COMP|9555-4|LNC|Cells.CD11c|Cells.CD11c
C0484531|T201|COMP|9556-2|LNC|Cells.CD11c+20c+|Cells.CD11c+20c+
C0484532|T201|COMP|8108-3|LNC|Cells.CD11c+CD20+/100 cells|Cells.CD11c+CD20+/100 cells
C0484533|T201|COMP|8109-1|LNC|Cells.CD11c/100 cells|Cells.CD11c/100 cells
C0484534|T201|COMP|8110-9|LNC|Cells.CD13/100 cells|Cells.CD13/100 cells
C0484535|T201|COMP|8111-7|LNC|Cells.CD14/100 cells|Cells.CD14/100 cells
C0484536|T201|COMP|8112-5|LNC|Cells.CD3-CD16+CD56+/100 cells|Cells.CD3-CD16+CD56+/100 cells
C0484537|T201|COMP|8113-3|LNC|Cells.CD16+CD57-/100 cells|Cells.CD16+CD57-/100 cells
C0484538|T201|COMP|8115-8|LNC|Cells.CD16/100 cells|Cells.CD16/100 cells
C0484539|T201|COMP|8116-6|LNC|Cells.CD19|Cells.CD19
C0484540|T201|COMP|8117-4|LNC|Cells.CD19/100 cells|Cells.CD19/100 cells
C0484541|T201|COMP|9557-0|LNC|Cells.CD2|Cells.CD2
C0484542|T201|COMP|8118-2|LNC|Cells.CD2/100 cells|Cells.CD2/100 cells
C0484543|T201|COMP|9558-8|LNC|Cells.CD20|Cells.CD20
C0484544|T201|COMP|8119-0|LNC|Cells.CD20/100 cells|Cells.CD20/100 cells
C0484545|T201|COMP|8120-8|LNC|Cells.CD21/100 cells|Cells.CD21/100 cells
C0484546|T201|COMP|8121-6|LNC|Cells.CD25/100 cells|Cells.CD25/100 cells
C0484547|T201|COMP|8122-4|LNC|Cells.CD3|Cells.CD3
C0484548|T201|COMP|8123-2|LNC|Cells.CD3+CD4+/100 cells|Cells.CD3+CD4+/100 cells
C0484549|T201|COMP|9728-7|LNC|Cells.CD3-CD16+CD56+|Cells.CD3-CD16+CD56+
C0484550|T201|COMP|8124-0|LNC|Cells.CD3/100 cells|Cells.CD3/100 cells
C0484551|T201|COMP|8125-7|LNC|Cells.CD34/100 cells|Cells.CD34/100 cells
C0484552|T201|COMP|8126-5|LNC|Cells.CD38/100 cells|Cells.CD38/100 cells
C0484553|T201|COMP|8127-3|LNC|Cells.CD4|Cells.CD4
C0484554|T201|COMP|8128-1|LNC|Cells.CD4/100 cells|Cells.CD4/100 cells
C0484555|T201|COMP|8129-9|LNC|Cells.CD4/Cells.CD8|Cells.CD4/Cells.CD8
C0484556|T201|COMP|8130-7|LNC|Cells.CD45/100 cells|Cells.CD45/100 cells
C0484557|T201|COMP|9559-6|LNC|Cells.CD5|Cells.CD5
C0484558|T201|COMP|9561-2|LNC|Cells.CD5+CD19+|Cells.CD5+CD19+
C0484559|T201|COMP|8131-5|LNC|Cells.CD5+CD19+/100 cells|Cells.CD5+CD19+/100 cells
C0484560|T201|COMP|9771-7|LNC|Cells.CD5+CD20+|Cells.CD5+CD20+
C0484561|T201|COMP|8132-3|LNC|Cells.CD5/100 cells|Cells.CD5/100 cells
C0484562|T201|COMP|8133-1|LNC|Cells.CD56/100 cells|Cells.CD56/100 cells
C0484563|T201|COMP|8134-9|LNC|Cells.CD57/100 cells|Cells.CD57/100 cells
C0484564|T201|COMP|9563-8|LNC|Cells.CD7|Cells.CD7
C0484565|T201|COMP|8135-6|LNC|Cells.CD7/100 cells|Cells.CD7/100 cells
C0484566|T201|COMP|8136-4|LNC|Cells.CD71/100 cells|Cells.CD71/100 cells
C0484567|T201|COMP|8137-2|LNC|Cells.CD8|Cells.CD8
C0484568|T201|COMP|8138-0|LNC|Cells.CD8/100 cells|Cells.CD8/100 cells
C0484569|T201|COMP|10447-1|LNC|M-5 Ag|M-5 Ag
C0484570|T201|COMP|10448-9|LNC|T-cell Ag|T-cell Ag
C0484571|T201|COMP|9612-3|LNC|Cortisol^15M post 250 ug corticotropin IM|Cortisol^15M post 250 ug corticotropin IM
C0484572|T201|COMP|9613-1|LNC|Cortisol^2H post 250 ug corticotropin IM|Cortisol^2H post 250 ug corticotropin IM
C0484573|T201|COMP|9614-9|LNC|Cortisol^45M post 250 ug corticotropin IM|Cortisol^45M post 250 ug corticotropin IM
C0484574|T201|COMP|9615-6|LNC|Cortisol^1.5H post 250 ug corticotropin IM|Cortisol^1.5H post 250 ug corticotropin IM
C0484575|T201|COMP|10332-5|LNC|Cortisol^pre 250 ug corticotropin IM|Cortisol^pre 250 ug corticotropin IM
C0484576|T201|COMP|6762-9|LNC|Glucose^1.5H post 50 g lactose PO|Glucose^1.5H post 50 g lactose PO
C0484577|T201|COMP|6761-1|LNC|Glucose^1.5H post 50 g lactose PO|Glucose^1.5H post 50 g lactose PO
C0484578|T201|COMP|6763-7|LNC|Glucose^1.5H post 75 g glucose PO|Glucose^1.5H post 75 g glucose PO
C0484579|T201|COMP|6747-0|LNC|Glucose^1H post 50 g lactose PO|Glucose^1H post 50 g lactose PO
C0484580|T201|COMP|6748-8|LNC|Glucose^1H post 75 g glucose PO|Glucose^1H post 75 g glucose PO
C0484581|T201|COMP|10449-7|LNC|Glucose^1H post meal|Glucose^1H post meal
C0484582|T201|COMP|9375-7|LNC|Glucose^2.5H post 100 g glucose PO|Glucose^2.5H post 100 g glucose PO
C0484583|T201|COMP|6749-6|LNC|Glucose^2.5H post 75 g glucose PO|Glucose^2.5H post 75 g glucose PO
C0484584|T201|COMP|6750-4|LNC|Glucose^2H post 50 g lactose PO|Glucose^2H post 50 g lactose PO
C0484585|T201|COMP|6751-2|LNC|Glucose^2H post 75 g glucose PO|Glucose^2H post 75 g glucose PO
C0484586|T201|COMP|6689-4|LNC|Glucose^2H post meal|Glucose^2H post meal
C0484587|T201|COMP|9376-5|LNC|Glucose^3.5H post 100 g glucose PO|Glucose^3.5H post 100 g glucose PO
C0484588|T201|COMP|6752-0|LNC|Glucose^3.5H post 75 g glucose PO|Glucose^3.5H post 75 g glucose PO
C0484589|T201|COMP|6753-8|LNC|Glucose^30M post 50 g lactose PO|Glucose^30M post 50 g lactose PO
C0484590|T201|COMP|6754-6|LNC|Glucose^30M post 75 g glucose PO|Glucose^30M post 75 g glucose PO
C0484591|T201|COMP|6755-3|LNC|Glucose^3H post 75 g glucose PO|Glucose^3H post 75 g glucose PO
C0484592|T201|COMP|9377-3|LNC|Glucose^4.5H post 100 g glucose PO|Glucose^4.5H post 100 g glucose PO
C0484593|T201|COMP|6756-1|LNC|Glucose^4.5H post 75 g glucose PO|Glucose^4.5H post 75 g glucose PO
C0484594|T201|COMP|6757-9|LNC|Glucose^4H post 75 g glucose PO|Glucose^4H post 75 g glucose PO
C0484595|T201|COMP|9378-1|LNC|Glucose^5.5H post 100 g glucose PO|Glucose^5.5H post 100 g glucose PO
C0484596|T201|COMP|6758-7|LNC|Glucose^5H post 75 g glucose PO|Glucose^5H post 75 g glucose PO
C0484597|T201|COMP|6760-3|LNC|Glucose^6H post 75 g glucose PO|Glucose^6H post 75 g glucose PO
C0484598|T201|COMP|6759-5|LNC|Glucose^6H post 75 g glucose PO|Glucose^6H post 75 g glucose PO
C0484599|T201|COMP|10450-5|LNC|Glucose^post 10H CFst|Glucose^post 10H CFst
C0484600|T201|COMP|6764-5|LNC|Glucose^post CFst|Glucose^post CFst
C0484601|T201|COMP|9307-0|LNC|Insulin^30M post 75 g glucose PO|Insulin^30M post 75 g glucose PO
C0484602|T201|COMP|9339-3|LNC|Insulin^6H post 75 g glucose PO|Insulin^6H post 75 g glucose PO
C0484603|T201|COMP|9570-3|LNC|Para aminobenzoate^6H post 500 mg bentiromide PO|Para aminobenzoate^6H post 500 mg bentiromide PO
C0484604|T201|COMP|10451-3|LNC|Proinsulin^post 12H CFst|Proinsulin^post 12H CFst
C0484605|T201|COMP|9772-5|LNC|Xylose^1H post 25 g xylose PO|Xylose^1H post 25 g xylose PO
C0484606|T201|COMP|10452-1|LNC|Xylose^1H post 25 g xylose PO|Xylose^1H post 25 g xylose PO
C0484607|T201|COMP|10453-9|LNC|Xylose^1H post dose xylose PO|Xylose^1H post dose xylose PO
C0484608|T201|COMP|10454-7|LNC|Xylose^2H post 25 g xylose PO|Xylose^2H post 25 g xylose PO
C0484609|T201|COMP|10455-4|LNC|Xylose^30M post 25 g xylose PO|Xylose^30M post 25 g xylose PO
C0484610|T201|COMP|10456-2|LNC|Xylose^post 6H CFst|Xylose^post 6H CFst
C0484611|T201|COMP|6865-0|LNC|1-Methylhistidine|1-Methylhistidine
C0484612|T201|COMP|6701-7|LNC|11-Hydroxyandrosterone|11-Hydroxyandrosterone
C0484613|T201|COMP|6700-9|LNC|11-Hydroxyetiocholanolone|11-Hydroxyetiocholanolone
C0484614|T201|COMP|6702-5|LNC|11-Ketoandrosterone|11-Ketoandrosterone
C0484615|T201|COMP|6703-3|LNC|11-Ketoetiocholanolone|11-Ketoetiocholanolone
C0484616|T201|COMP|6704-1|LNC|11-Ketopregnanetriol|11-Ketopregnanetriol
C0484617|T201|COMP|9445-8|LNC|11-Oxopregnanetriol|11-Oxopregnanetriol
C0484618|T201|COMP|6866-8|LNC|17-Hydroxycorticosteroids|17-Hydroxycorticosteroids
C0484619|T201|COMP|6765-2|LNC|17-Hydroxypregnenolone|17-Hydroxypregnenolone
C0484620|T201|COMP|9616-4|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C0484621|T201|COMP|6766-0|LNC|17-Ketosteroids|17-Ketosteroids
C0484622|T201|COMP|6767-8|LNC|18-Hydroxycorticosteroids|18-Hydroxycorticosteroids
C0484623|T201|COMP|9639-6|LNC|18-Hydroxycorticosterone|18-Hydroxycorticosterone
C0484624|T201|COMP|9308-8|LNC|2,4-Dinitrophenylhydrazine reacting substances|2,4-Dinitrophenylhydrazine reacting substances
C0484625|T201|COMP|9695-8|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C0484626|T201|COMP|6867-6|LNC|3-Methylhistidine|3-Methylhistidine
C0484627|T201|COMP|10457-0|LNC|Actin Ag|Actin Ag
C0484628|T201|COMP|9402-9|LNC|Acyl carnitine|Acyl carnitine
C0484629|T201|COMP|9403-7|LNC|Acylcarnitine|Acylcarnitine
C0484630|T201|COMP|9404-5|LNC|Adenosine deaminase|Adenosine deaminase
C0484631|T201|COMP|6868-4|LNC|Adenosine monophosphate.cyclic|Adenosine monophosphate.cyclic
C0484632|T201|COMP|9318-7|LNC|Albumin/Creatinine|Albumin/Creatinine
C0484633|T201|COMP|9406-0|LNC|Albumin/Globulin|Albumin/Globulin
C0484634|T201|COMP|9405-2|LNC|Albumin/Globulin|Albumin/Globulin
C0484637|T201|COMP|10458-8|LNC|Alkaline phosphatase.placental Ag|Alkaline phosphatase.placental Ag
C0484638|T201|COMP|6768-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0484639|T201|COMP|6869-2|LNC|Allo-tetrahydrocortisol|Allo-tetrahydrocortisol
C0484640|T201|COMP|9734-5|LNC|Alpha 1 globulin|Alpha 1 globulin
C0484641|T201|COMP|6870-0|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0484642|T201|COMP|6935-1|LNC|Alpha aminoadipate|Alpha aminoadipate
C0484643|T201|COMP|10459-6|LNC|Alpha-1-Fetoprotein Ag|Alpha-1-Fetoprotein Ag
C0484644|T201|COMP|10460-4|LNC|Lactalbumin alpha Ag|Lactalbumin alpha Ag
C0484645|T201|COMP|10461-2|LNC|Alpha-1-Antichymotrypsin Ag|Alpha-1-Antichymotrypsin Ag
C0484646|T201|COMP|10462-0|LNC|Alpha 1 antitrypsin Ag|Alpha 1 antitrypsin Ag
C0484647|T201|COMP|6770-2|LNC|Alpha 1 antitrypsin phenotyping|Alpha 1 antitrypsin phenotyping
C0484648|T201|COMP|6771-0|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C0484649|T201|COMP|9407-8|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C0484650|T201|COMP|9408-6|LNC|Aminobenzoate|Aminobenzoate
C0484651|T201|COMP|9309-6|LNC|Ammonia|Ammonia
C0484652|T201|COMP|1798-8|LNC|Amylase|Amylase
C0484653|T201|COMP|10463-8|LNC|Amyloid A component Ag|Amyloid A component Ag
C0484654|T201|COMP|10464-6|LNC|Amyloid P component Ag|Amyloid P component Ag
C0484655|T201|COMP|10465-3|LNC|Amyloid.prealbumin Ag|Amyloid.prealbumin Ag
C0484656|T201|COMP|9409-4|LNC|Anabolic steroids|Anabolic steroids
C0484657|T201|COMP|9640-4|LNC|Androstanediol|Androstanediol
C0484658|T201|COMP|9310-4|LNC|Androstenedione|Androstenedione
C0484659|T201|COMP|6705-8|LNC|Androsterone|Androsterone
C0484660|T201|COMP|10466-1|LNC|Anion gap 3|Anion gap 3
C0484661|T201|COMP|6871-8|LNC|Anserine|Anserine
C0484662|T201|COMP|1874-7|LNC|Apolipoprotein B/Apolipoprotein A-I|Apolipoprotein B/Apolipoprotein A-I
C0484663|T201|COMP|9340-1|LNC|Apolipoprotein B/Apolipoprotein A-I|Apolipoprotein B/Apolipoprotein A-I
C0484664|T201|COMP|10333-3|LNC|Appearance|Appearance
C0484665|T201|COMP|1903-4|LNC|Ascorbate|Ascorbate
C0484666|T201|COMP|6872-6|LNC|Beta alanine|Beta alanine
C0484667|T201|COMP|9320-3|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0484668|T201|COMP|9744-4|LNC|Beta globulin|Beta globulin
C0484669|T201|COMP|9829-3|LNC|Beta globulin|Beta globulin
C0484670|T201|COMP|6873-4|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C0484671|T201|COMP|10467-9|LNC|Beta-2-Microglobulin amyloid Ag|Beta-2-Microglobulin amyloid Ag
C0484672|T201|COMP|10468-7|LNC|Calcitonin Ag|Calcitonin Ag
C0484673|T201|COMP|6874-2|LNC|Calcium|Calcium
C0484674|T201|COMP|9321-1|LNC|Calcium/Creatinine|Calcium/Creatinine
C0484675|T201|COMP|10334-1|LNC|Cancer Ag 125|Cancer Ag 125
C0484676|T201|COMP|6875-9|LNC|Cancer Ag 15-3|Cancer Ag 15-3
C0484677|T201|COMP|10469-5|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0484678|T201|COMP|9641-2|LNC|Catecholamines/Creatinine|Catecholamines/Creatinine
C0484679|T201|COMP|9794-9|LNC|Cathepsin D|Cathepsin D
C0484680|T201|COMP|9341-9|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C0484681|T201|COMP|9742-8|LNC|Chloride|Chloride
C0484682|T201|COMP|9342-7|LNC|Cholesterol|Cholesterol
C0484683|T201|COMP|9830-1|LNC|Cholesterol.total/Cholesterol.in HDL|Cholesterol.total/Cholesterol.in HDL
C0484684|T201|COMP|9322-9|LNC|Cholesterol.total/Cholesterol.in HDL|Cholesterol.total/Cholesterol.in HDL
C0484685|T201|COMP|9509-1|LNC|Cholinesterase|Cholinesterase
C0484686|T201|COMP|10470-3|LNC|Choriogonadotropin Ag|Choriogonadotropin Ag
C0484687|T201|COMP|9811-1|LNC|Chromogranin A|Chromogranin A
C0484688|T201|COMP|10471-1|LNC|Chromogranin A Ag|Chromogranin A Ag
C0484689|T201|COMP|10472-9|LNC|Chromogranin Ag|Chromogranin Ag
C0484690|T201|COMP|9617-2|LNC|Chylomicrons|Chylomicrons
C0484691|T201|COMP|10473-7|LNC|Chymotrypsin Ag|Chymotrypsin Ag
C0484692|T201|COMP|6687-8|LNC|Citrate|Citrate
C0484693|T201|COMP|9511-7|LNC|Citrulline|Citrulline
C0484694|T201|COMP|6876-7|LNC|Citrulline|Citrulline
C0484695|T201|COMP|10474-5|LNC|Collagen type 4 Ag|Collagen type 4 Ag
C0484696|T201|COMP|10335-8|LNC|Color|Color
C0484697|T201|COMP|9343-5|LNC|Coproporphyrin 1|Coproporphyrin 1
C0484698|T201|COMP|6877-5|LNC|Coproporphyrin 1|Coproporphyrin 1
C0484699|T201|COMP|9344-3|LNC|Coproporphyrin 1/Coproporphyrin.total|Coproporphyrin 1/Coproporphyrin.total
C0484700|T201|COMP|9345-0|LNC|Coproporphyrin 3|Coproporphyrin 3
C0484701|T201|COMP|6878-3|LNC|Coproporphyrin 3|Coproporphyrin 3
C0484702|T201|COMP|6879-1|LNC|Corticotropin|Corticotropin
C0484703|T201|COMP|10475-2|LNC|Corticotropin Ag|Corticotropin Ag
C0484704|T201|COMP|9812-9|LNC|Cortisol^PM trough specimen|Cortisol^PM trough specimen
C0484705|T201|COMP|9813-7|LNC|Cortisol^AM peak specimen|Cortisol^AM peak specimen
C0484706|T201|COMP|9642-0|LNC|Creatine kinase.BB/Creatine kinase.total|Creatine kinase.BB/Creatine kinase.total
C0484707|T201|COMP|6773-6|LNC|Creatine kinase.MB|Creatine kinase.MB
C0484708|T201|COMP|9643-8|LNC|Creatine kinase.MM/Creatine kinase.total|Creatine kinase.MM/Creatine kinase.total
C0484709|T201|COMP|6880-9|LNC|Cystathionine|Cystathionine
C0484710|T201|COMP|9644-6|LNC|Cystine|Cystine
C0484711|T201|COMP|6699-3|LNC|Delta 5-Pregnanetriol|Delta 5-Pregnanetriol
C0484712|T201|COMP|6937-7|LNC|Deoxypyridinoline|Deoxypyridinoline
C0484713|T201|COMP|6936-9|LNC|Deoxypyridinoline|Deoxypyridinoline
C0484715|T201|COMP|10476-0|LNC|Desmin Ag|Desmin Ag
C0484716|T201|COMP|6775-1|LNC|Androstanolone|Androstanolone
C0484717|T201|COMP|10477-8|LNC|Enolase.neuron specific Ag|Enolase.neuron specific Ag
C0484718|T201|COMP|10478-6|LNC|Eosinophil major basic protein Ag|Eosinophil major basic protein Ag
C0484719|T201|COMP|10479-4|LNC|CD227 Ag|CD227 Ag
C0484720|T201|COMP|10480-2|LNC|Estrogen+Progesterone receptor Ag|Estrogen+Progesterone receptor Ag
C0484721|T201|COMP|6776-9|LNC|Estrone|Estrone
C0484722|T201|COMP|6881-7|LNC|Ethanolamine|Ethanolamine
C0484723|T201|COMP|10481-0|LNC|Follitropin.alpha subunit Ag|Follitropin.alpha subunit Ag
C0484724|T201|COMP|10482-8|LNC|Follitropin.beta subunit Ag|Follitropin.beta subunit Ag
C0484725|T201|COMP|6882-5|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0484726|T201|COMP|9745-1|LNC|Gamma globulin|Gamma globulin
C0484727|T201|COMP|9831-9|LNC|Gamma globulin|Gamma globulin
C0484728|T201|COMP|10483-6|LNC|Gastrin Ag|Gastrin Ag
C0484729|T201|COMP|10484-4|LNC|Glial fibrillary acidic protein Ag|Glial fibrillary acidic protein Ag
C0484730|T201|COMP|10485-1|LNC|Glucagon Ag|Glucagon Ag
C0484731|T201|COMP|2345-7|LNC|Glucose|Glucose
C0484732|T201|COMP|6883-3|LNC|Glucose.protein bound|Glucose.protein bound
C0484733|T201|COMP|9379-9|LNC|Glutathione reductase|Glutathione reductase
C0484734|T201|COMP|10336-6|LNC|Gonadotropin peptide|Gonadotropin peptide
C0484735|T201|COMP|9832-7|LNC|Cholesterol.in HDL 2|Cholesterol.in HDL 2
C0484736|T201|COMP|9833-5|LNC|Cholesterol.in HDL 3|Cholesterol.in HDL 3
C0484737|T201|COMP|10486-9|LNC|Hemoglobin Ag|Hemoglobin Ag
C0484738|T201|COMP|9447-4|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C0484739|T201|COMP|9446-6|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C0484740|T201|COMP|9380-7|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C0484741|T201|COMP|9448-2|LNC|Heptaporphyrin|Heptaporphyrin
C0484742|T201|COMP|9449-0|LNC|Heptaporphyrin|Heptaporphyrin
C0484743|T201|COMP|9451-6|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C0484744|T201|COMP|9450-8|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C0484745|T201|COMP|9527-3|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C0484746|T201|COMP|9452-4|LNC|Hexaporphyrin|Hexaporphyrin
C0484747|T201|COMP|6709-0|LNC|Hippurate|Hippurate
C0484748|T201|COMP|9410-2|LNC|Histamine|Histamine
C0484749|T201|COMP|9453-2|LNC|Histidine|Histidine
C0484750|T201|COMP|10487-7|LNC|HMB-45 Ag|HMB-45 Ag
C0484751|T201|COMP|6884-1|LNC|Homocystine|Homocystine
C0484752|T201|COMP|9411-0|LNC|Hydrocorticosterone|Hydrocorticosterone
C0484753|T201|COMP|6885-8|LNC|Hydroxylysine|Hydroxylysine
C0484754|T201|COMP|2447-1|LNC|Hydroxyproline|Hydroxyproline
C0484755|T201|COMP|6938-5|LNC|IgA|IgA
C0484756|T201|COMP|6778-5|LNC|IgA|IgA
C0484757|T201|COMP|6779-3|LNC|IgA|IgA
C0484758|T201|COMP|10488-5|LNC|IgA Ag|IgA Ag
C0484759|T201|COMP|6886-6|LNC|IgA subclass 1|IgA subclass 1
C0484761|T201|COMP|6939-3|LNC|IgA subclass 2|IgA subclass 2
C0484762|T201|COMP|10489-3|LNC|IgA.heavy chain Ag|IgA.heavy chain Ag
C0484763|T201|COMP|10490-1|LNC|IgE Ag|IgE Ag
C0484764|T201|COMP|6780-1|LNC|IgG|IgG
C0484765|T201|COMP|6781-9|LNC|IgG|IgG
C0484766|T201|COMP|10491-9|LNC|IgG Ag|IgG Ag
C0484767|T201|COMP|10492-7|LNC|IgG.heavy chain Ag|IgG.heavy chain Ag
C0484768|T201|COMP|6782-7|LNC|IgG/Albumin|IgG/Albumin
C0484769|T201|COMP|6783-5|LNC|IgM|IgM
C0484770|T201|COMP|6784-3|LNC|IgM|IgM
C0484771|T201|COMP|10493-5|LNC|IgM Ag|IgM Ag
C0484772|T201|COMP|10494-3|LNC|IgM.heavy chain Ag|IgM.heavy chain Ag
C0484773|T201|COMP|6785-0|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C0484774|T201|COMP|6787-6|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C0484775|T201|COMP|6786-8|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C0484777|T201|COMP|6789-2|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C0484778|T201|COMP|6791-8|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C0484779|T201|COMP|6790-0|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C0484780|T201|COMP|6887-4|LNC|Indicans|Indicans
C0484781|T201|COMP|10495-0|LNC|Insulin Ag|Insulin Ag
C0484782|T201|COMP|9537-2|LNC|Intrinsic factor blocking Ab|Intrinsic factor blocking Ab
C0484783|T201|COMP|9743-6|LNC|Isoleucine|Isoleucine
C0484784|T201|COMP|10496-8|LNC|Immunoglobulin light chains.kappa Ag|Immunoglobulin light chains.kappa Ag
C0484785|T201|COMP|10497-6|LNC|Immunoglobulin light chains.kappa amyloid Ag|Immunoglobulin light chains.kappa amyloid Ag
C0484786|T201|COMP|10498-4|LNC|Keratin Ag|Keratin Ag
C0484787|T201|COMP|10499-2|LNC|Immunoglobulin light chains.lambda Ag|Immunoglobulin light chains.lambda Ag
C0484788|T201|COMP|10500-7|LNC|Immunoglobulin light chains.lambda amyloid Ag|Immunoglobulin light chains.lambda amyloid Ag
C0484789|T201|COMP|9412-8|LNC|Leucine|Leucine
C0484790|T201|COMP|9618-0|LNC|Cholesterol|Cholesterol
C0484791|T201|COMP|9413-6|LNC|Lipids|Lipids
C0484792|T201|COMP|9619-8|LNC|Triglyceride|Triglyceride
C0484793|T201|COMP|9620-6|LNC|Lipoprotein.beta|Lipoprotein.beta
C0484794|T201|COMP|9346-8|LNC|Lipoprotein.beta|Lipoprotein.beta
C0484795|T201|COMP|9621-4|LNC|Lipoprotein.pre-beta|Lipoprotein.pre-beta
C0484796|T201|COMP|10501-5|LNC|Lutropin|Lutropin
C0484797|T201|COMP|6692-8|LNC|Lutropin|Lutropin
C0484798|T201|COMP|10502-3|LNC|Lutropin Ag|Lutropin Ag
C0484799|T201|COMP|10503-1|LNC|Lysozyme Ag|Lysozyme Ag
C0484800|T201|COMP|9645-3|LNC|Metanephrine/Creatinine|Metanephrine/Creatinine
C0484801|T201|COMP|10504-9|LNC|Myelin basic protein Ag|Myelin basic protein Ag
C0484802|T201|COMP|10505-6|LNC|Myoglobin Ag|Myoglobin Ag
C0484803|T201|COMP|10506-4|LNC|Peanut agglutinin Ag|Peanut agglutinin Ag
C0484804|T201|COMP|9730-3|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C0484806|T201|COMP|9347-6|LNC|pH.combined acid|pH.combined acid
C0484807|T201|COMP|9348-4|LNC|pH.free acid|pH.free acid
C0484808|T201|COMP|9349-2|LNC|pH.total acid|pH.total acid
C0484809|T201|COMP|9731-1|LNC|Phosphoethanolamine|Phosphoethanolamine
C0484810|T201|COMP|9414-4|LNC|Phosphoserine|Phosphoserine
C0484811|T201|COMP|9732-9|LNC|Phosphoserine|Phosphoserine
C0484812|T201|COMP|9622-2|LNC|Phytonadione|Phytonadione
C0484813|T201|COMP|9733-7|LNC|Porphyrins|Porphyrins
C0484814|T201|COMP|6792-6|LNC|Potassium|Potassium
C0484815|T201|COMP|6940-1|LNC|Potassium|Potassium
C0484816|T201|COMP|9482-1|LNC|Potassium|Potassium
C0484817|T201|COMP|10337-4|LNC|Procollagen type I|Procollagen type I
C0484818|T201|COMP|10507-2|LNC|Prolactin Ag|Prolactin Ag
C0484819|T201|COMP|10508-0|LNC|Prostate specific Ag|Prostate specific Ag
C0484820|T201|COMP|10509-8|LNC|Acid phosphatase.prostatic Ag|Acid phosphatase.prostatic Ag
C0484821|T201|COMP|6888-2|LNC|Alpha 2 globulin|Alpha 2 globulin
C0484822|T201|COMP|6889-0|LNC|Beta globulin|Beta globulin
C0484823|T201|COMP|6890-8|LNC|Gamma globulin|Gamma globulin
C0484824|T201|COMP|6793-4|LNC|Prealbumin|Prealbumin
C0484825|T201|COMP|6942-7|LNC|Albumin|Albumin
C0484826|T201|COMP|6941-9|LNC|Albumin|Albumin
C0484827|T201|COMP|6794-2|LNC|Alpha 1 globulin|Alpha 1 globulin
C0484828|T201|COMP|6795-9|LNC|Alpha 2 globulin|Alpha 2 globulin
C0484829|T201|COMP|9381-5|LNC|Pyridinoline|Pyridinoline
C0484830|T201|COMP|6695-1|LNC|Riboflavin|Riboflavin
C0484831|T201|COMP|10510-6|LNC|S-100 Ag|S-100 Ag
C0484832|T201|COMP|9323-7|LNC|Sarcosine|Sarcosine
C0484833|T201|COMP|10511-4|LNC|Serotonin Ag|Serotonin Ag
C0484834|T201|COMP|9485-4|LNC|Sodium|Sodium
C0484835|T201|COMP|10512-2|LNC|Somatostatin Ag|Somatostatin Ag
C0484836|T201|COMP|10513-0|LNC|Somatotropin Ag|Somatotropin Ag
C0484837|T201|COMP|9486-2|LNC|Sulfate|Sulfate
C0484838|T201|COMP|9350-0|LNC|Sulfhydryls|Sulfhydryls
C0484839|T201|COMP|9646-1|LNC|Sulfide|Sulfide
C0484840|T201|COMP|10514-8|LNC|Synaptophysin Ag|Synaptophysin Ag
C0484841|T201|COMP|9324-5|LNC|Taurine|Taurine
C0484842|T201|COMP|6891-6|LNC|Testosterone.free+weakly bound/Testosterone.total|Testosterone.free+weakly bound/Testosterone.total
C0484843|T201|COMP|9382-3|LNC|Coproporphyrin|Coproporphyrin
C0484844|T201|COMP|9579-4|LNC|Tetrahydrocorticosterone|Tetrahydrocorticosterone
C0484845|T201|COMP|9647-9|LNC|Thiosulfate|Thiosulfate
C0484846|T201|COMP|10515-5|LNC|Thyroglobulin Ag|Thyroglobulin Ag
C0484847|T201|COMP|10516-3|LNC|Thyrotropin Ag|Thyrotropin Ag
C0484848|T201|COMP|6892-4|LNC|Thyroxine.free|Thyroxine.free
C0484849|T201|COMP|6796-7|LNC|Transferrin saturation|Transferrin saturation
C0484850|T201|COMP|6597-9|LNC|Troponin T.cardiac|Troponin T.cardiac
C0484851|T201|COMP|6598-7|LNC|Troponin T.cardiac|Troponin T.cardiac
C0484852|T201|COMP|10517-1|LNC|Trypsin Ag|Trypsin Ag
C0484853|T201|COMP|9325-2|LNC|Tryptophan|Tryptophan
C0484854|T201|COMP|10518-9|LNC|Ulex europaeus I lectin Ag|Ulex europaeus I lectin Ag
C0484855|T201|COMP|6893-2|LNC|Urobilinogen|Urobilinogen
C0484856|T201|COMP|9735-2|LNC|Uroporphyrin/Porphyrins.total|Uroporphyrin/Porphyrins.total
C0484857|T201|COMP|9623-0|LNC|Valine|Valine
C0484858|T201|COMP|9624-8|LNC|Vanillylmandelate|Vanillylmandelate
C0484859|T201|COMP|10519-7|LNC|Vimentin Ag|Vimentin Ag
C0484862|T201|COMP|10520-5|LNC|Coagulation factor VI Ag|Coagulation factor VI Ag
C0484863|T201|COMP|10521-3|LNC|Coagulation factor VIII Ag|Coagulation factor VIII Ag
C0484864|T201|COMP|10522-1|LNC|Coagulation factor XIII Ag|Coagulation factor XIII Ag
C0484865|T201|COMP|6683-7|LNC|Coagulation reptilase induced|Coagulation reptilase induced
C0484866|T201|COMP|6684-5|LNC|Coagulation reptilase induced|Coagulation reptilase induced
C0484867|T201|COMP|7799-0|LNC|Fibrin D-dimer|Fibrin D-dimer
C0484868|T201|COMP|10523-9|LNC|Fibrinogen Ag|Fibrinogen Ag
C0484869|T201|COMP|7800-6|LNC|Phospholipid Ab|Phospholipid Ab
C0484870|T201|COMP|7801-4|LNC|Phospholipid Ab.IgG|Phospholipid Ab.IgG
C0484871|T201|COMP|7802-2|LNC|Phospholipid Ab.IgM|Phospholipid Ab.IgM
C0484877|T201|COMP|9696-6|LNC|8-Hydroxyloxapine|8-Hydroxyloxapine
C0484878|T201|COMP|9383-1|LNC|9-Hydroxyrisperidone|9-Hydroxyrisperidone
C0484879|T201|COMP|6943-5|LNC|acetoHEXAMIDE|acetoHEXAMIDE
C0484880|T201|COMP|10528-8|LNC|Acetophenazine|Acetophenazine
C0484881|T201|COMP|9416-9|LNC|Acyclovir|Acyclovir
C0484882|T201|COMP|9311-2|LNC|Albuterol|Albuterol
C0484883|T201|COMP|9736-0|LNC|Allopurinol|Allopurinol
C0484884|T201|COMP|9351-8|LNC|ALPRAZolam|ALPRAZolam
C0484885|T201|COMP|9312-0|LNC|Aminocaproate|Aminocaproate
C0484886|T201|COMP|10529-6|LNC|Amoxapine metabolite|Amoxapine metabolite
C0484887|T201|COMP|9625-5|LNC|Amoxapine+8-Hydroxyamoxapine|Amoxapine+8-Hydroxyamoxapine
C0484888|T201|COMP|9352-6|LNC|Amphetamines|Amphetamines
C0484889|T201|COMP|9417-7|LNC|Anthraquinone|Anthraquinone
C0484890|T201|COMP|10530-4|LNC|Aprobarbital|Aprobarbital
C0484891|T201|COMP|6894-0|LNC|Zidovudine|Zidovudine
C0484892|T201|COMP|9353-4|LNC|Baclofen|Baclofen
C0484893|T201|COMP|10338-2|LNC|Barbiturates|Barbiturates
C0484894|T201|COMP|9384-9|LNC|Benztropine|Benztropine
C0484895|T201|COMP|9354-2|LNC|Benztropine|Benztropine
C0484896|T201|COMP|10531-2|LNC|Bretylium|Bretylium
C0484897|T201|COMP|9355-9|LNC|Bumetanide|Bumetanide
C0484898|T201|COMP|6706-6|LNC|buPROPion|buPROPion
C0484899|T201|COMP|9356-7|LNC|busPIRone|busPIRone
C0484900|T201|COMP|6895-7|LNC|Butalbital|Butalbital
C0484901|T201|COMP|9313-8|LNC|Butorphanol|Butorphanol
C0484902|T201|COMP|9415-1|LNC|carBAMazepine 10,11-Epoxide|carBAMazepine 10,11-Epoxide
C0484903|T201|COMP|9328-6|LNC|Carbidopa|Carbidopa
C0484904|T201|COMP|3042-9|LNC|Chloral hydrate|Chloral hydrate
C0484905|T201|COMP|17738-6|LNC|Chloral hydrate|Chloral hydrate
C0484906|T201|COMP|9508-3|LNC|Chlorothiazide|Chlorothiazide
C0484907|T201|COMP|9648-7|LNC|Chlorothiazide|Chlorothiazide
C0484908|T201|COMP|6896-5|LNC|cloZAPine|cloZAPine
C0484909|T201|COMP|6797-5|LNC|Cyclobenzaprine|Cyclobenzaprine
C0484910|T201|COMP|9746-9|LNC|Dantrolene|Dantrolene
C0484911|T201|COMP|9747-7|LNC|Dapsone|Dapsone
C0484912|T201|COMP|6774-4|LNC|Desethylamiodarone|Desethylamiodarone
C0484914|T201|COMP|9814-5|LNC|Dextroamphetamine|Dextroamphetamine
C0484915|T201|COMP|9737-8|LNC|Propoxyphene|Propoxyphene
C0484916|T201|COMP|10533-8|LNC|Propoxyphene+Acetaminophen|Propoxyphene+Acetaminophen
C0484917|T201|COMP|9626-3|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C0484918|T201|COMP|10534-6|LNC|Diazoxide|Diazoxide
C0484919|T201|COMP|9515-8|LNC|Diclofenac|Diclofenac
C0484920|T201|COMP|10535-3|LNC|Digoxin|Digoxin
C0484921|T201|COMP|6898-1|LNC|dilTIAZem|dilTIAZem
C0484922|T201|COMP|10536-1|LNC|Dipyridamole|Dipyridamole
C0484923|T201|COMP|9748-5|LNC|Dipyridamole|Dipyridamole
C0484924|T201|COMP|9357-5|LNC|Disulfiram|Disulfiram
C0484926|T201|COMP|9773-3|LNC|Ergotamine|Ergotamine
C0484927|T201|COMP|6899-9|LNC|Felbamate|Felbamate
C0484928|T201|COMP|10339-0|LNC|Fluoxetine+Norfluoxetine|Fluoxetine+Norfluoxetine
C0484930|T201|COMP|9738-6|LNC|Gabapentin|Gabapentin
C0484931|T201|COMP|10539-5|LNC|glipiZIDE|glipiZIDE
C0484932|T201|COMP|6944-3|LNC|glipiZIDE|glipiZIDE
C0484933|T201|COMP|6900-5|LNC|Glutethimide|Glutethimide
C0484934|T201|COMP|10540-3|LNC|glyBURIDE|glyBURIDE
C0484935|T201|COMP|6945-0|LNC|glyBURIDE|glyBURIDE
C0484936|T201|COMP|9649-5|LNC|Hydroflumethiazide|Hydroflumethiazide
C0484937|T201|COMP|9834-3|LNC|HYDROmorphone|HYDROmorphone
C0484938|T201|COMP|9835-0|LNC|HYDROmorphone|HYDROmorphone
C0484939|T201|COMP|9418-5|LNC|Hydroxybupropion|Hydroxybupropion
C0484940|T201|COMP|6946-8|LNC|Imipramine|Imipramine
C0484941|T201|COMP|9627-1|LNC|Imipramine+Desipramine|Imipramine+Desipramine
C0484942|T201|COMP|6901-3|LNC|Insulin.free|Insulin.free
C0484943|T201|COMP|6947-6|LNC|ISOtretinoin|ISOtretinoin
C0484944|T201|COMP|6948-4|LNC|lamoTRIgine|lamoTRIgine
C0484945|T201|COMP|9385-6|LNC|Levodopa|Levodopa
C0484946|T201|COMP|9815-2|LNC|Lithium|Lithium
C0484947|T201|COMP|9358-3|LNC|Lithium|Lithium
C0484948|T201|COMP|6691-0|LNC|Loxapine+8-Hydroxyamoxapine|Loxapine+8-Hydroxyamoxapine
C0484949|T201|COMP|10541-1|LNC|Mepivacaine|Mepivacaine
C0484950|T201|COMP|2609-6|LNC|Metanephrines|Metanephrines
C0484951|T201|COMP|6949-2|LNC|Metaproterenol|Metaproterenol
C0484952|T201|COMP|6902-1|LNC|Methadone|Methadone
C0484953|T201|COMP|10542-9|LNC|Metharbital|Metharbital
C0484955|T201|COMP|9650-3|LNC|Methyclothiazide|Methyclothiazide
C0484956|T201|COMP|9774-1|LNC|Metoclopramide|Metoclopramide
C0484957|T201|COMP|9651-1|LNC|metOLazone|metOLazone
C0484958|T201|COMP|10340-8|LNC|Molindone|Molindone
C0484959|T201|COMP|9775-8|LNC|Moricizine|Moricizine
C0484960|T201|COMP|9438-3|LNC|Morphine|Morphine
C0484961|T201|COMP|9652-9|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0484963|T201|COMP|9777-4|LNC|Nalbuphine|Nalbuphine
C0484964|T201|COMP|9740-2|LNC|Neopterin|Neopterin
C0484965|T201|COMP|9386-4|LNC|NIFEdipine|NIFEdipine
C0484966|T201|COMP|3536-0|LNC|Norclomipramine|Norclomipramine
C0484967|T201|COMP|10544-5|LNC|Normeperidine|Normeperidine
C0484968|T201|COMP|10545-2|LNC|Normephenytoin|Normephenytoin
C0484969|T201|COMP|10546-0|LNC|Normethsuximide|Normethsuximide
C0484970|T201|COMP|10341-6|LNC|Norpropoxyphene|Norpropoxyphene
C0484971|T201|COMP|6903-9|LNC|Norverapamil|Norverapamil
C0484972|T201|COMP|9628-9|LNC|Norvenlafaxine|Norvenlafaxine
C0484973|T201|COMP|9699-0|LNC|PARoxetine|PARoxetine
C0484974|T201|COMP|9778-2|LNC|Phenelzine|Phenelzine
C0484975|T201|COMP|10547-8|LNC|Primidone+PHENobarbital|Primidone+PHENobarbital
C0484976|T201|COMP|6904-7|LNC|Phenothiazine|Phenothiazine
C0484977|T201|COMP|10548-6|LNC|Phenytoin.free/Phenytoin.total|Phenytoin.free/Phenytoin.total
C0484978|T201|COMP|10549-4|LNC|Pirmenol|Pirmenol
C0484979|T201|COMP|9700-6|LNC|Procaine|Procaine
C0484980|T201|COMP|9387-2|LNC|Procyclidine|Procyclidine
C0484981|T201|COMP|6905-4|LNC|Propafenone|Propafenone
C0484982|T201|COMP|9388-0|LNC|Propylthiouracil|Propylthiouracil
C0484983|T201|COMP|9389-8|LNC|Pseudoephedrine|Pseudoephedrine
C0484984|T201|COMP|9390-6|LNC|Pyridostigmine|Pyridostigmine
C0484985|T201|COMP|9391-4|LNC|Quazepam|Quazepam
C0484986|T201|COMP|9392-2|LNC|Quinethazone|Quinethazone
C0484987|T201|COMP|6694-4|LNC|quiNIDine|quiNIDine
C0484988|T201|COMP|9779-0|LNC|quiNIDine.free|quiNIDine.free
C0484989|T201|COMP|6950-0|LNC|raNITIdine|raNITIdine
C0484990|T201|COMP|9393-0|LNC|risperiDONE|risperiDONE
C0484991|T201|COMP|9394-8|LNC|Risperidone+9-Hydroxyrisperidone|Risperidone+9-Hydroxyrisperidone
C0484992|T201|COMP|6906-2|LNC|Sertraline|Sertraline
C0484993|T201|COMP|9395-5|LNC|SUFentanil|SUFentanil
C0484994|T201|COMP|9396-3|LNC|SUFentanil|SUFentanil
C0484995|T201|COMP|6907-0|LNC|sulfADIAZINE|sulfADIAZINE
C0484996|T201|COMP|10342-4|LNC|Sulfamethoxazole|Sulfamethoxazole
C0484997|T201|COMP|9701-4|LNC|sulfiSOXAZOLE|sulfiSOXAZOLE
C0484998|T201|COMP|9359-1|LNC|Tacrine|Tacrine
C0485000|T201|COMP|10343-2|LNC|Temazepam|Temazepam
C0485001|T201|COMP|9702-2|LNC|Terbutaline|Terbutaline
C0485002|T201|COMP|6696-9|LNC|Thiothixene|Thiothixene
C0485003|T201|COMP|9629-7|LNC|TOLAZamide|TOLAZamide
C0485004|T201|COMP|6951-8|LNC|TOLAZamide|TOLAZamide
C0485005|T201|COMP|6952-6|LNC|TOLBUTamide|TOLBUTamide
C0485006|T201|COMP|10344-0|LNC|Tranylcypromine|Tranylcypromine
C0485007|T201|COMP|10551-0|LNC|Triamterene|Triamterene
C0485008|T201|COMP|9653-7|LNC|Trichlormethiazide|Trichlormethiazide
C0485009|T201|COMP|6799-1|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0485010|T201|COMP|10552-8|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0485011|T201|COMP|9703-0|LNC|Trihexyphenidyl|Trihexyphenidyl
C0485012|T201|COMP|10345-7|LNC|Trihexyphenidyl|Trihexyphenidyl
C0485013|T201|COMP|9630-5|LNC|Venlafaxine|Venlafaxine
C0485014|T201|COMP|6953-4|LNC|Zolpidem|Zolpidem
C0485015|T201|COMP|10553-6|LNC|Acid phosphatase.prostatic|Acid phosphatase.prostatic
C0485016|T201|COMP|10554-4|LNC|Acid phosphatase.prostatic|Acid phosphatase.prostatic
C0485017|T201|COMP|10555-1|LNC|Acrosin|Acrosin
C0485018|T201|COMP|10556-9|LNC|Adenosine triphosphatase|Adenosine triphosphatase
C0485019|T201|COMP|10557-7|LNC|Adenosine triphosphate|Adenosine triphosphate
C0485020|T201|COMP|10558-5|LNC|Albumin|Albumin
C0485021|T201|COMP|10559-3|LNC|Calcium|Calcium
C0485022|T201|COMP|10560-1|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0485023|T201|COMP|10561-9|LNC|Carnitine|Carnitine
C0485024|T201|COMP|10562-7|LNC|Cells|Cells
C0485025|T201|COMP|10563-5|LNC|Cells other than spermatozoa|Cells other than spermatozoa
C0485026|T201|COMP|10564-3|LNC|Cervical mucus|Cervical mucus
C0485027|T201|COMP|10565-0|LNC|Choriogonadotropin|Choriogonadotropin
C0485028|T201|COMP|10566-8|LNC|Choriogonadotropin|Choriogonadotropin
C0485029|T201|COMP|10567-6|LNC|Citrate|Citrate
C0485030|T201|COMP|10568-4|LNC|Clarity|Clarity
C0485031|T201|COMP|10569-2|LNC|Color|Color
C0485032|T201|COMP|10570-0|LNC|Consistency|Consistency
C0485033|T201|COMP|10571-8|LNC|Consistency|Consistency
C0485034|T201|COMP|10572-6|LNC|Duration^post ejaculation|Duration^post ejaculation
C0485036|T201|COMP|10574-2|LNC|Fructose|Fructose
C0485037|T201|COMP|10575-9|LNC|Gamma glutamyl transferase|Gamma glutamyl transferase
C0485038|T201|COMP|10576-7|LNC|Germ cells.immature|Germ cells.immature
C0485039|T201|COMP|10577-5|LNC|Glucosidase|Glucosidase
C0485040|T201|COMP|10578-3|LNC|Glycerophosphocholine|Glycerophosphocholine
C0485041|T201|COMP|10579-1|LNC|Leukocytes|Leukocytes
C0485042|T201|COMP|10580-9|LNC|Liquefaction|Liquefaction
C0485043|T201|COMP|10581-7|LNC|Number of entities|Number of entities
C0485045|T201|COMP|10583-3|LNC|Prostaglandin F1 alpha|Prostaglandin F1 alpha
C0485046|T201|COMP|10584-1|LNC|Protein|Protein
C0485047|T201|COMP|10585-8|LNC|Round cells|Round cells
C0485048|T201|COMP|10586-6|LNC|Semen|Semen
C0485049|T201|COMP|10587-4|LNC|Sexual abstinence duration|Sexual abstinence duration
C0485050|T201|COMP|6800-7|LNC|Spermatozoa.motile/100 spermatozoa|Spermatozoa.motile/100 spermatozoa
C0485051|T201|COMP|10588-2|LNC|Spermatogonia|Spermatogonia
C0485052|T201|COMP|10589-0|LNC|Spermatids|Spermatids
C0485053|T201|COMP|10590-8|LNC|Spermatids|Spermatids
C0485054|T201|COMP|10591-6|LNC|Spermatocytes.primary|Spermatocytes.primary
C0485055|T201|COMP|10592-4|LNC|Spermatocytes.secondary|Spermatocytes.secondary
C0485056|T201|COMP|9704-8|LNC|Spermatozoa|Spermatozoa
C0485057|T201|COMP|9780-8|LNC|Spermatozoa|Spermatozoa
C0485058|T201|COMP|10596-5|LNC|Spermatozoa Ab|Spermatozoa Ab
C0485059|T201|COMP|10598-1|LNC|Spermatozoa Ab|Spermatozoa Ab
C0485060|T201|COMP|10597-3|LNC|Spermatozoa Ab|Spermatozoa Ab
C0485062|T201|COMP|10599-9|LNC|Spermatozoa penetration|Spermatozoa penetration
C0485063|T201|COMP|10600-5|LNC|Spermatozoa penetration|Spermatozoa penetration
C0485064|T201|COMP|10601-3|LNC|Spermatozoa penetration^post coitus|Spermatozoa penetration^post coitus
C0485065|T201|COMP|10602-1|LNC|Spermatozoa.abnormal head/100 spermatozoa|Spermatozoa.abnormal head/100 spermatozoa
C0485066|T201|COMP|10603-9|LNC|Spermatozoa.abnormal midpiece/100 spermatozoa|Spermatozoa.abnormal midpiece/100 spermatozoa
C0485067|T201|COMP|10604-7|LNC|Spermatozoa.abnormal tail/100 spermatozoa|Spermatozoa.abnormal tail/100 spermatozoa
C0485068|T201|COMP|10605-4|LNC|Spermatozoa.agglutinated/100 spermatozoa|Spermatozoa.agglutinated/100 spermatozoa
C0485069|T201|COMP|10606-2|LNC|Spermatozoa.amorphous head/100 spermatozoa|Spermatozoa.amorphous head/100 spermatozoa
C0485070|T201|COMP|10607-0|LNC|Spermatozoa.coiled tail/100 spermatozoa|Spermatozoa.coiled tail/100 spermatozoa
C0485071|T201|COMP|10608-8|LNC|Spermatozoa.cytoplasmic droplet/100 spermatozoa|Spermatozoa.cytoplasmic droplet/100 spermatozoa
C0485072|T201|COMP|10609-6|LNC|Spermatozoa.duplicate head/100 spermatozoa|Spermatozoa.duplicate head/100 spermatozoa
C0485073|T201|COMP|10610-4|LNC|Spermatozoa.duplicate tail/100 spermatozoa|Spermatozoa.duplicate tail/100 spermatozoa
C0485074|T201|COMP|10611-2|LNC|Spermatozoa.immotile/100 spermatozoa|Spermatozoa.immotile/100 spermatozoa
C0485075|T201|COMP|10612-0|LNC|Spermatozoa.large oval head/100 spermatozoa|Spermatozoa.large oval head/100 spermatozoa
C0485076|T201|COMP|10613-8|LNC|Spermatozoa.viable/100 spermatozoa|Spermatozoa.viable/100 spermatozoa
C0485077|T201|COMP|10614-6|LNC|Spermatozoa.motile with IgA/100 spermatozoa|Spermatozoa.motile with IgA/100 spermatozoa
C0485078|T201|COMP|10615-3|LNC|Spermatozoa.motile with IgA/100 spermatozoa|Spermatozoa.motile with IgA/100 spermatozoa
C0485079|T201|COMP|10616-1|LNC|Spermatozoa.motile with IgG/100 spermatozoa|Spermatozoa.motile with IgG/100 spermatozoa
C0485080|T201|COMP|10617-9|LNC|Spermatozoa.motile with IgG/100 spermatozoa|Spermatozoa.motile with IgG/100 spermatozoa
C0485081|T201|COMP|10618-7|LNC|Spermatozoa.motile with IgM/100 spermatozoa|Spermatozoa.motile with IgM/100 spermatozoa
C0485082|T201|COMP|10619-5|LNC|Spermatozoa.motile with IgM/100 spermatozoa|Spermatozoa.motile with IgM/100 spermatozoa
C0485083|T201|COMP|10620-3|LNC|Spermatozoa.nonprogressive/100 spermatozoa|Spermatozoa.nonprogressive/100 spermatozoa
C0485084|T201|COMP|10621-1|LNC|Spermatozoa.normal head/100 spermatozoa|Spermatozoa.normal head/100 spermatozoa
C0485085|T201|COMP|10622-9|LNC|Spermatozoa.normal/100 spermatozoa|Spermatozoa.normal/100 spermatozoa
C0485086|T201|COMP|10623-7|LNC|Spermatozoa.pin head/100 spermatozoa|Spermatozoa.pin head/100 spermatozoa
C0485087|T201|COMP|10593-2|LNC|Spermatozoa.pyriform head/100 spermatozoa|Spermatozoa.pyriform head/100 spermatozoa
C0485088|T201|COMP|10624-5|LNC|Spermatozoa.rapid/100 spermatozoa|Spermatozoa.rapid/100 spermatozoa
C0485089|T201|COMP|10625-2|LNC|Spermatozoa.round head/100 spermatozoa|Spermatozoa.round head/100 spermatozoa
C0485090|T201|COMP|10626-0|LNC|Spermatozoa.slow/100 spermatozoa|Spermatozoa.slow/100 spermatozoa
C0485091|T201|COMP|10627-8|LNC|Spermatozoa.small oval head/100 spermatozoa|Spermatozoa.small oval head/100 spermatozoa
C0485092|T201|COMP|10628-6|LNC|Spermatozoa.tail swelling/100 spermatozoa|Spermatozoa.tail swelling/100 spermatozoa
C0485093|T201|COMP|10594-0|LNC|Spermatozoa.tapering head/100 spermatozoa|Spermatozoa.tapering head/100 spermatozoa
C0485094|T201|COMP|10629-4|LNC|Spermatozoa.vacuolated head/100 spermatozoa|Spermatozoa.vacuolated head/100 spermatozoa
C0485095|T201|COMP|10630-2|LNC|Spinnbarkeit|Spinnbarkeit
C0485096|T201|COMP|10631-0|LNC|Testosterone|Testosterone
C0485097|T201|COMP|10632-8|LNC|Time until next menstrual period|Time until next menstrual period
C0485098|T201|COMP|9631-3|LNC|Viscosity|Viscosity
C0485099|T201|COMP|10633-6|LNC|Zinc|Zinc
C0485101|T201|COMP|6801-5|LNC|Complement C3|Complement C3
C0485102|T201|COMP|6908-8|LNC|Complement C4|Complement C4
C0485103|T201|COMP|10346-5|LNC|Hemoglobin A|Hemoglobin A
C0485104|T201|COMP|9749-3|LNC|Hemoglobin F|Hemoglobin F
C0485105|T201|COMP|9654-5|LNC|Interleukin 2 receptor.soluble|Interleukin 2 receptor.soluble
C0485106|T201|COMP|6909-6|LNC|Mucin clot|Mucin clot
C0485107|T201|COMP|6864-3|LNC|Hemoglobin S|Hemoglobin S
C0485108|T201|COMP|9419-3|LNC|HLA-DQ6|HLA-DQ6
C0485109|T201|COMP|6802-3|LNC|HLA-DR10|HLA-DR10
C0485110|T201|COMP|6803-1|LNC|HLA-DR15|HLA-DR15
C0485111|T201|COMP|6804-9|LNC|HLA-DR52|HLA-DR52
C0485112|T201|COMP|6805-6|LNC|HLA-DR53|HLA-DR53
C0485113|T201|COMP|6806-4|LNC|HLA-DR6|HLA-DR6
C0485114|T201|COMP|6807-2|LNC|HLA-DR8|HLA-DR8
C0485115|T201|COMP|6618-3|LNC|Acanthamoeba sp Ab|Acanthamoeba sp Ab
C0485116|T201|COMP|6619-1|LNC|Acanthamoeba sp Ab|Acanthamoeba sp Ab
C0485117|T201|COMP|6620-9|LNC|Acanthamoeba sp Ab|Acanthamoeba sp Ab
C0485118|T201|COMP|7803-0|LNC|Acanthamoeba sp Ab|Acanthamoeba sp Ab
C0485119|T201|COMP|10635-1|LNC|Acanthamoeba sp identified|Acanthamoeba sp identified
C0485120|T201|COMP|10636-9|LNC|Acanthamoeba sp identified|Acanthamoeba sp identified
C0485121|T201|COMP|9781-6|LNC|Acanthamoeba sp identified|Acanthamoeba sp identified
C0485123|T201|COMP|7804-8|LNC|Actinomyces sp Ab|Actinomyces sp Ab
C0485124|T201|COMP|9816-0|LNC|Actinomyces sp identified|Actinomyces sp identified
C0485125|T201|COMP|10638-5|LNC|Actinomycetes.thermophilic colony count|Actinomycetes.thermophilic colony count
C0485126|T201|COMP|10639-3|LNC|Actinomycetes.thermophilic identified|Actinomycetes.thermophilic identified
C0485127|T201|COMP|10640-1|LNC|Adenovirus 40+41|Adenovirus 40+41
C0485128|T201|COMP|7805-5|LNC|Adenovirus Ab|Adenovirus Ab
C0485129|T201|COMP|9782-4|LNC|Adenovirus sp identified|Adenovirus sp identified
C0485130|T201|COMP|9582-8|LNC|Afipia felis Ab.IgG|Afipia felis Ab.IgG
C0485131|T201|COMP|9583-6|LNC|Afipia felis Ab.IgM|Afipia felis Ab.IgM
C0485132|T201|COMP|10641-9|LNC|Amoeba identified|Amoeba identified
C0485133|T201|COMP|10642-7|LNC|Amoeba identified|Amoeba identified
C0485134|T201|COMP|10643-5|LNC|Amoeba identified|Amoeba identified
C0485135|T201|COMP|6594-6|LNC|Amoeba identified|Amoeba identified
C0485136|T201|COMP|10644-3|LNC|Arthropod identified|Arthropod identified
C0485137|T201|COMP|7806-3|LNC|Ascaris lumbricoides Ab|Ascaris lumbricoides Ab
C0485138|T201|COMP|9490-4|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C0485139|T201|COMP|9492-0|LNC|Aspergillus sp Ab.IgM|Aspergillus sp Ab.IgM
C0485140|T201|COMP|10645-0|LNC|Aspergillus fumigatus Ag|Aspergillus fumigatus Ag
C0485141|T201|COMP|6808-0|LNC|Aspergillus fumigatus 1 Ab|Aspergillus fumigatus 1 Ab
C0485142|T201|COMP|6809-8|LNC|Aspergillus fumigatus 6 Ab|Aspergillus fumigatus 6 Ab
C0485143|T201|COMP|9632-1|LNC|Aspergillus fumigatus Ab|Aspergillus fumigatus Ab
C0485144|T201|COMP|7807-1|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C0485145|T201|COMP|7808-9|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C0485146|T201|COMP|9491-2|LNC|Aspergillus sp Ab.IgA|Aspergillus sp Ab.IgA
C0485147|T201|COMP|7809-7|LNC|Astrovirus|Astrovirus
C0485148|T201|COMP|10646-8|LNC|Astrovirus|Astrovirus
C0485149|T201|COMP|7810-5|LNC|Astrovirus Ag|Astrovirus Ag
C0485150|T201|COMP|7811-3|LNC|Astrovirus RNA|Astrovirus RNA
C0485151|T201|COMP|6810-6|LNC|Aureobasidium pullulans Ab|Aureobasidium pullulans Ab
C0485152|T201|COMP|9584-4|LNC|Babesia sp Ab.IgG|Babesia sp Ab.IgG
C0485153|T201|COMP|9585-1|LNC|Babesia sp Ab.IgM|Babesia sp Ab.IgM
C0485154|T201|COMP|7812-1|LNC|Babesia microti Ab|Babesia microti Ab
C0485155|T201|COMP|10347-3|LNC|Babesia microti identified|Babesia microti identified
C0485156|T201|COMP|7813-9|LNC|Babesia sp Ab|Babesia sp Ab
C0485157|T201|COMP|10647-6|LNC|Babesia sp identified|Babesia sp identified
C0485158|T201|COMP|10648-4|LNC|Babesia sp identified|Babesia sp identified
C0485159|T201|COMP|7814-7|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0485160|T201|COMP|7815-4|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C0485161|T201|COMP|6954-2|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C0485162|T201|COMP|6955-9|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C0485163|T201|COMP|8009-3|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C0485164|T201|COMP|9360-9|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C0485165|T201|COMP|8010-1|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C0485166|T201|COMP|9361-7|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C0485167|T201|COMP|7816-2|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0485168|T201|COMP|9494-6|LNC|Blastomyces dermatitidis Ab.IgG|Blastomyces dermatitidis Ab.IgG
C0485169|T201|COMP|10348-1|LNC|Bordetella parapertussis Ab|Bordetella parapertussis Ab
C0485170|T201|COMP|9362-5|LNC|Bordetella pertussis Ab.IgA|Bordetella pertussis Ab.IgA
C0485171|T201|COMP|9363-3|LNC|Bordetella pertussis Ab.IgG|Bordetella pertussis Ab.IgG
C0485172|T201|COMP|9364-1|LNC|Bordetella pertussis Ab.IgM|Bordetella pertussis Ab.IgM
C0485173|T201|COMP|9588-5|LNC|Borrelia burgdorferi 18kD Ab.IgG|Borrelia burgdorferi 18kD Ab.IgG
C0485174|T201|COMP|9589-3|LNC|Borrelia burgdorferi 23kD Ab.IgG|Borrelia burgdorferi 23kD Ab.IgG
C0485175|T201|COMP|9598-4|LNC|Borrelia burgdorferi 23kD Ab.IgM|Borrelia burgdorferi 23kD Ab.IgM
C0485176|T201|COMP|9590-1|LNC|Borrelia burgdorferi 28kD Ab.IgG|Borrelia burgdorferi 28kD Ab.IgG
C0485177|T201|COMP|9591-9|LNC|Borrelia burgdorferi 30kD Ab.IgG|Borrelia burgdorferi 30kD Ab.IgG
C0485178|T201|COMP|9592-7|LNC|Borrelia burgdorferi 39kD Ab.IgG|Borrelia burgdorferi 39kD Ab.IgG
C0485179|T201|COMP|9599-2|LNC|Borrelia burgdorferi 39kD Ab.IgM|Borrelia burgdorferi 39kD Ab.IgM
C0485180|T201|COMP|9593-5|LNC|Borrelia burgdorferi 41kD Ab.IgG|Borrelia burgdorferi 41kD Ab.IgG
C0485181|T201|COMP|9587-7|LNC|Borrelia burgdorferi 41kD Ab.IgM|Borrelia burgdorferi 41kD Ab.IgM
C0485182|T201|COMP|9594-3|LNC|Borrelia burgdorferi 45kD Ab.IgG|Borrelia burgdorferi 45kD Ab.IgG
C0485183|T201|COMP|9595-0|LNC|Borrelia burgdorferi 58kD Ab.IgG|Borrelia burgdorferi 58kD Ab.IgG
C0485184|T201|COMP|9596-8|LNC|Borrelia burgdorferi 66kD Ab.IgG|Borrelia burgdorferi 66kD Ab.IgG
C0485185|T201|COMP|9597-6|LNC|Borrelia burgdorferi 93kD Ab.IgG|Borrelia burgdorferi 93kD Ab.IgG
C0485186|T201|COMP|9586-9|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0485187|T201|COMP|7817-0|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0485188|T201|COMP|7818-8|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0485189|T201|COMP|6910-4|LNC|Brucella abortus Ab.IgA|Brucella abortus Ab.IgA
C0485190|T201|COMP|6911-2|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C0485191|T201|COMP|9495-3|LNC|Brucella canis Ab.IgG|Brucella canis Ab.IgG
C0485192|T201|COMP|9496-1|LNC|Brucella canis Ab.IgM|Brucella canis Ab.IgM
C0485193|T201|COMP|10349-9|LNC|Brucella sp Ab|Brucella sp Ab
C0485194|T201|COMP|6606-8|LNC|Brugia malayi Ab|Brugia malayi Ab
C0485195|T201|COMP|7819-6|LNC|Brugia malayi Ab|Brugia malayi Ab
C0485196|T201|COMP|10649-2|LNC|Calicivirus|Calicivirus
C0485197|T201|COMP|6595-3|LNC|Klebsiella granulomatis|Klebsiella granulomatis
C0485198|T201|COMP|9655-2|LNC|Campylobacter jejuni Ab|Campylobacter jejuni Ab
C0485199|T201|COMP|7820-4|LNC|Candida albicans Ab|Candida albicans Ab
C0485200|T201|COMP|9498-7|LNC|Candida sp Ab.IgA|Candida sp Ab.IgA
C0485201|T201|COMP|9500-0|LNC|Candida sp Ab.IgM|Candida sp Ab.IgM
C0485202|T201|COMP|9501-8|LNC|Candida sp Ag|Candida sp Ag
C0485203|T201|COMP|10650-0|LNC|Candida sp DNA|Candida sp DNA
C0485204|T201|COMP|6912-0|LNC|Chlamydophila pneumoniae Ab.IgA|Chlamydophila pneumoniae Ab.IgA
C0485205|T201|COMP|6913-8|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C0485206|T201|COMP|6914-6|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C0485207|T201|COMP|10651-8|LNC|Chlamydophila pneumoniae Ag|Chlamydophila pneumoniae Ag
C0485208|T201|COMP|10652-6|LNC|Chlamydophila pneumoniae DNA|Chlamydophila pneumoniae DNA
C0485209|T201|COMP|7821-2|LNC|Chlamydophila pneumoniae rRNA|Chlamydophila pneumoniae rRNA
C0485210|T201|COMP|7822-0|LNC|Chlamydophila psittaci Ab|Chlamydophila psittaci Ab
C0485211|T201|COMP|6915-3|LNC|Chlamydophila psittaci Ab.IgA|Chlamydophila psittaci Ab.IgA
C0485212|T201|COMP|6916-1|LNC|Chlamydophila psittaci Ab.IgG|Chlamydophila psittaci Ab.IgG
C0485213|T201|COMP|6917-9|LNC|Chlamydophila psittaci Ab.IgM|Chlamydophila psittaci Ab.IgM
C0485214|T201|COMP|7823-8|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0485215|T201|COMP|7824-6|LNC|Chlamydia trachomatis Ab|Chlamydia trachomatis Ab
C0485216|T201|COMP|6918-7|LNC|Chlamydia trachomatis Ab.IgA|Chlamydia trachomatis Ab.IgA
C0485217|T201|COMP|6919-5|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C0485218|T201|COMP|6920-3|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C0485219|T201|COMP|9365-8|LNC|Clostridioides difficile Ab|Clostridioides difficile Ab
C0485220|T201|COMP|10653-4|LNC|Clotrimazole|Clotrimazole
C0485221|T201|COMP|10654-2|LNC|Clotrimazole|Clotrimazole
C0485222|T201|COMP|10655-9|LNC|Coccidia identified|Coccidia identified
C0485223|T201|COMP|10656-7|LNC|Coccidia identified|Coccidia identified
C0485224|T201|COMP|7825-3|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0485225|T201|COMP|9705-5|LNC|Coccidioides immitis Ab.IgA|Coccidioides immitis Ab.IgA
C0485226|T201|COMP|7826-1|LNC|Coccidioides immitis Ab.IgG|Coccidioides immitis Ab.IgG
C0485227|T201|COMP|7827-9|LNC|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C0485228|T201|COMP|9764-2|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C0485229|T201|COMP|7828-7|LNC|Coxiella burnetii Ab|Coxiella burnetii Ab
C0485230|T201|COMP|7829-5|LNC|Coxiella burnetii phase 1 Ab.IgG|Coxiella burnetii phase 1 Ab.IgG
C0485231|T201|COMP|7830-3|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C0485232|T201|COMP|7831-1|LNC|Coxiella burnetii phase 1 Ab.IgM|Coxiella burnetii phase 1 Ab.IgM
C0485233|T201|COMP|7832-9|LNC|Coxiella burnetii phase 2 Ab.IgM|Coxiella burnetii phase 2 Ab.IgM
C0485234|T201|COMP|9706-3|LNC|Coxiella burnetii phase 1 Ab.IgA|Coxiella burnetii phase 1 Ab.IgA
C0485235|T201|COMP|9708-9|LNC|Coxiella burnetii phase 1 Ab.IgG|Coxiella burnetii phase 1 Ab.IgG
C0485236|T201|COMP|9710-5|LNC|Coxiella burnetii phase 1 Ab.IgM|Coxiella burnetii phase 1 Ab.IgM
C0485237|T201|COMP|9707-1|LNC|Coxiella burnetii phase 2 Ab.IgA|Coxiella burnetii phase 2 Ab.IgA
C0485238|T201|COMP|9709-7|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C0485239|T201|COMP|9711-3|LNC|Coxiella burnetii phase 2 Ab.IgM|Coxiella burnetii phase 2 Ab.IgM
C0485240|T201|COMP|9751-9|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C0485241|T201|COMP|9750-1|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C0485242|T201|COMP|9752-7|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C0485243|T201|COMP|7833-7|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C0485244|T201|COMP|6688-6|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C0485245|T201|COMP|9753-5|LNC|Coxsackievirus A2 Ab|Coxsackievirus A2 Ab
C0485246|T201|COMP|6956-7|LNC|Coxsackievirus A21 Ab|Coxsackievirus A21 Ab
C0485247|T201|COMP|9754-3|LNC|Coxsackievirus A4 Ab|Coxsackievirus A4 Ab
C0485248|T201|COMP|9756-8|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C0485249|T201|COMP|7834-5|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C0485250|T201|COMP|9755-0|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C0485251|T201|COMP|9758-4|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C0485252|T201|COMP|7835-2|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C0485253|T201|COMP|9757-6|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C0485254|T201|COMP|9759-2|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C0485255|T201|COMP|7836-0|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C0485256|T201|COMP|9760-0|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C0485257|T201|COMP|7837-8|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C0485258|T201|COMP|9761-8|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C0485259|T201|COMP|7838-6|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C0485260|T201|COMP|9762-6|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C0485261|T201|COMP|7839-4|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C0485262|T201|COMP|9763-4|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C0485263|T201|COMP|7840-2|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C0485264|T201|COMP|7841-0|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C0485265|T201|COMP|7842-8|LNC|Cryptococcus neoformans Ab|Cryptococcus neoformans Ab
C0485266|T201|COMP|10657-5|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C0485267|T201|COMP|7843-6|LNC|Cryptococcus sp Ab|Cryptococcus sp Ab
C0485268|T201|COMP|9817-8|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C0485269|T201|COMP|9819-4|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C0485270|T201|COMP|9818-6|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C0485271|T201|COMP|9820-2|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C0485272|T201|COMP|10658-3|LNC|Cyanobacterium identified|Cyanobacterium identified
C0485273|T201|COMP|10659-1|LNC|Cyclospora sp identified|Cyclospora sp identified
C0485274|T201|COMP|9601-6|LNC|Taenia solium larva 13kD Ab|Taenia solium larva 13kD Ab
C0485275|T201|COMP|9602-4|LNC|Taenia solium larva 14kD Ab|Taenia solium larva 14kD Ab
C0485276|T201|COMP|9603-2|LNC|Taenia solium larva 18kD Ab|Taenia solium larva 18kD Ab
C0485277|T201|COMP|9604-0|LNC|Taenia solium larva 21kD Ab|Taenia solium larva 21kD Ab
C0485278|T201|COMP|9605-7|LNC|Taenia solium larva 24kD Ab|Taenia solium larva 24kD Ab
C0485279|T201|COMP|9606-5|LNC|Taenia solium larva 39-42kD Ab|Taenia solium larva 39-42kD Ab
C0485280|T201|COMP|9607-3|LNC|Taenia solium larva 50kD Ab|Taenia solium larva 50kD Ab
C0485281|T201|COMP|9600-8|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C0485282|T201|COMP|7844-4|LNC|Taenia solium larva Ab.IgA|Taenia solium larva Ab.IgA
C0485283|T201|COMP|7845-1|LNC|Taenia solium larva Ab.IgA|Taenia solium larva Ab.IgA
C0485284|T201|COMP|7846-9|LNC|Taenia solium larva Ab.IgG|Taenia solium larva Ab.IgG
C0485285|T201|COMP|7847-7|LNC|Taenia solium larva Ab.IgG|Taenia solium larva Ab.IgG
C0485286|T201|COMP|7848-5|LNC|Taenia solium larva Ab.IgM|Taenia solium larva Ab.IgM
C0485287|T201|COMP|7849-3|LNC|Taenia solium larva Ab.IgM|Taenia solium larva Ab.IgM
C0485288|T201|COMP|7850-1|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C0485289|T201|COMP|9514-1|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0485290|T201|COMP|7851-9|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0485291|T201|COMP|9513-3|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0485292|T201|COMP|6921-1|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0485293|T201|COMP|7852-7|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0485294|T201|COMP|7853-5|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0485295|T201|COMP|10660-9|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0485296|T201|COMP|7854-3|LNC|Dengue virus 1 Ab|Dengue virus 1 Ab
C0485297|T201|COMP|7855-0|LNC|Dengue virus 1+2+3+4 RNA|Dengue virus 1+2+3+4 RNA
C0485298|T201|COMP|7856-8|LNC|Dengue virus 2 Ab|Dengue virus 2 Ab
C0485299|T201|COMP|7857-6|LNC|Dengue virus 3 Ab|Dengue virus 3 Ab
C0485300|T201|COMP|7858-4|LNC|Dengue virus 4 Ab|Dengue virus 4 Ab
C0485301|T201|COMP|7859-2|LNC|Dengue virus Ab|Dengue virus Ab
C0485302|T201|COMP|6811-4|LNC|Dengue virus Ab.IgG|Dengue virus Ab.IgG
C0485303|T201|COMP|6812-2|LNC|Dengue virus Ab.IgM|Dengue virus Ab.IgM
C0485304|T201|COMP|10661-7|LNC|Dinoflagellate identified|Dinoflagellate identified
C0485305|T201|COMP|6596-1|LNC|Diphtheria sp identified|Diphtheria sp identified
C0485306|T201|COMP|7860-0|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C0485307|T201|COMP|7861-8|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C0485308|T201|COMP|7862-6|LNC|Ebola virus Ab|Ebola virus Ab
C0485309|T201|COMP|7863-4|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0485310|T201|COMP|9656-0|LNC|Echinococcus sp Ab.IgG|Echinococcus sp Ab.IgG
C0485311|T201|COMP|9657-8|LNC|Echinococcus sp Ab.IgM|Echinococcus sp Ab.IgM
C0485312|T201|COMP|7864-2|LNC|Echovirus 1 Ab|Echovirus 1 Ab
C0485313|T201|COMP|9516-6|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C0485314|T201|COMP|7865-9|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C0485315|T201|COMP|6708-2|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C0485316|T201|COMP|6813-0|LNC|Echovirus 16 Ab|Echovirus 16 Ab
C0485317|T201|COMP|9517-4|LNC|Echovirus 18 Ab|Echovirus 18 Ab
C0485318|T201|COMP|7866-7|LNC|Echovirus 19 Ab|Echovirus 19 Ab
C0485319|T201|COMP|7867-5|LNC|Echovirus 3 Ab|Echovirus 3 Ab
C0485320|T201|COMP|9518-2|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C0485321|T201|COMP|7868-3|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C0485322|T201|COMP|9519-0|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C0485323|T201|COMP|7869-1|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C0485324|T201|COMP|7870-9|LNC|Echovirus 40 Ab|Echovirus 40 Ab
C0485325|T201|COMP|7871-7|LNC|Echovirus 6 Ab|Echovirus 6 Ab
C0485326|T201|COMP|6922-9|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C0485327|T201|COMP|9520-8|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C0485328|T201|COMP|7872-5|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C0485329|T201|COMP|16795-7|LNC|Echovirus Ab|Echovirus Ab
C0485330|T201|COMP|7874-1|LNC|Ehrlichia canis Ab|Ehrlichia canis Ab
C0485331|T201|COMP|7875-8|LNC|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C0485332|T201|COMP|9783-2|LNC|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C0485333|T201|COMP|7876-6|LNC|Ehrlichia chaffeensis Ab.IgM|Ehrlichia chaffeensis Ab.IgM
C0485334|T201|COMP|9784-0|LNC|Ehrlichia chaffeensis Ab.IgM|Ehrlichia chaffeensis Ab.IgM
C0485335|T201|COMP|7877-4|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C0485335|T201|COMP|7878-2|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C0485335|T201|COMP|20810-8|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C0485337|T201|COMP|7879-0|LNC|Ehrlichia sp Ab|Ehrlichia sp Ab
C0485339|T201|COMP|7880-8|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0485340|T201|COMP|9421-9|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0485341|T201|COMP|9420-1|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0485342|T201|COMP|9521-6|LNC|Entamoeba histolytica Ab.IgA|Entamoeba histolytica Ab.IgA
C0485343|T201|COMP|9522-4|LNC|Entamoeba histolytica Ab.IgG|Entamoeba histolytica Ab.IgG
C0485344|T201|COMP|9523-2|LNC|Entamoeba histolytica Ab.IgM|Entamoeba histolytica Ab.IgM
C0485345|T201|COMP|7881-6|LNC|Enterovirus RNA|Enterovirus RNA
C0485346|T201|COMP|6814-8|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C0485347|T201|COMP|6815-5|LNC|Epstein Barr virus nuclear Ab.IgM|Epstein Barr virus nuclear Ab.IgM
C0485348|T201|COMP|7882-4|LNC|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C0485349|T201|COMP|7883-2|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0485350|T201|COMP|7884-0|LNC|Epstein Barr virus nuclear Ab.IgM|Epstein Barr virus nuclear Ab.IgM
C0485351|T201|COMP|9633-9|LNC|Epstein Barr virus capsid Ab.IgA|Epstein Barr virus capsid Ab.IgA
C0485352|T201|COMP|7885-7|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0485353|T201|COMP|7886-5|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0485354|T201|COMP|7887-3|LNC|Filaria Ab|Filaria Ab
C0485355|T201|COMP|10662-5|LNC|Filaria identified|Filaria identified
C0485356|T201|COMP|10663-3|LNC|Filaria identified|Filaria identified
C0485357|T201|COMP|10664-1|LNC|Filaria identified|Filaria identified
C0485358|T201|COMP|7888-1|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C0485359|T201|COMP|7889-9|LNC|Francisella tularensis Ab.IgG|Francisella tularensis Ab.IgG
C0485360|T201|COMP|7890-7|LNC|Francisella tularensis Ab.IgM|Francisella tularensis Ab.IgM
C0485361|T201|COMP|10665-8|LNC|Fungus colony count|Fungus colony count
C0485362|T201|COMP|10666-6|LNC|Fungus identified|Fungus identified
C0485363|T201|COMP|10667-4|LNC|Fungus identified|Fungus identified
C0485364|T201|COMP|10668-2|LNC|Fungus identified|Fungus identified
C0485365|T201|COMP|10669-0|LNC|Fungus identified|Fungus identified
C0485366|T201|COMP|9524-0|LNC|Giardia lamblia Ab|Giardia lamblia Ab
C0485367|T201|COMP|9658-6|LNC|Giardia lamblia Ab.IgA|Giardia lamblia Ab.IgA
C0485368|T201|COMP|7891-5|LNC|Giardia lamblia Ab.IgG|Giardia lamblia Ab.IgG
C0485369|T201|COMP|7892-3|LNC|Giardia lamblia Ab.IgM|Giardia lamblia Ab.IgM
C0485370|T201|COMP|10670-8|LNC|Giardia lamblia|Giardia lamblia
C0485371|T201|COMP|7893-1|LNC|Gliadin Ab|Gliadin Ab
C0485372|T201|COMP|7894-9|LNC|Haemophilus influenzae Ab|Haemophilus influenzae Ab
C0485373|T201|COMP|6610-0|LNC|Haemophilus influenzae A Ag|Haemophilus influenzae A Ag
C0485374|T201|COMP|6611-8|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C0485375|T201|COMP|6599-5|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C0485376|T201|COMP|6612-6|LNC|Haemophilus influenzae C Ag|Haemophilus influenzae C Ag
C0485377|T201|COMP|8271-9|LNC|Haemophilus influenzae C Ag|Haemophilus influenzae C Ag
C0485378|T201|COMP|6613-4|LNC|Haemophilus influenzae D Ag|Haemophilus influenzae D Ag
C0485379|T201|COMP|6614-2|LNC|Haemophilus influenzae E Ag|Haemophilus influenzae E Ag
C0485380|T201|COMP|6615-9|LNC|Haemophilus influenzae F Ag|Haemophilus influenzae F Ag
C0485381|T201|COMP|6600-1|LNC|Haemophilus sp identified|Haemophilus sp identified
C0485382|T201|COMP|7895-6|LNC|Hantavirus hantaan Ab.IgG|Hantavirus hantaan Ab.IgG
C0485383|T201|COMP|7896-4|LNC|Hantavirus hantaan Ab.IgM|Hantavirus hantaan Ab.IgM
C0485384|T201|COMP|7897-2|LNC|Hantavirus puumala Ab.IgG|Hantavirus puumala Ab.IgG
C0485385|T201|COMP|7898-0|LNC|Hantavirus puumala Ab.IgM|Hantavirus puumala Ab.IgM
C0485386|T201|COMP|7899-8|LNC|Hantavirus RNA|Hantavirus RNA
C0485387|T201|COMP|7900-4|LNC|Helicobacter pylori Ab|Helicobacter pylori Ab
C0485388|T201|COMP|7901-2|LNC|Helicobacter pylori Ab.IgA|Helicobacter pylori Ab.IgA
C0485389|T201|COMP|7902-0|LNC|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C0485390|T201|COMP|7903-8|LNC|Helicobacter pylori Ab.IgM|Helicobacter pylori Ab.IgM
C0485391|T201|COMP|10671-6|LNC|Helminth identified|Helminth identified
C0485392|T201|COMP|10672-4|LNC|Helminth+Arthropod identified|Helminth+Arthropod identified
C0485393|T201|COMP|7904-6|LNC|Hepatitis A virus RNA|Hepatitis A virus RNA
C0485394|T201|COMP|10673-2|LNC|Hepatitis B virus core Ag|Hepatitis B virus core Ag
C0485395|T201|COMP|10674-0|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C0485396|T201|COMP|10675-7|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C0485397|T201|COMP|7905-3|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C0485398|T201|COMP|10676-5|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C0485399|T201|COMP|9608-1|LNC|Hepatitis C virus 100-3 Ab|Hepatitis C virus 100-3 Ab
C0485400|T201|COMP|9609-9|LNC|Hepatitis C virus 22-3 Ab|Hepatitis C virus 22-3 Ab
C0485401|T201|COMP|9610-7|LNC|Hepatitis C virus c33c Ab|Hepatitis C virus c33c Ab
C0485402|T201|COMP|9526-5|LNC|Hepatitis D virus Ag|Hepatitis D virus Ag
C0485403|T201|COMP|9525-7|LNC|Hepatitis D virus Ab.IgM|Hepatitis D virus Ab.IgM
C0485404|T201|COMP|7906-1|LNC|Hepatitis D virus RNA|Hepatitis D virus RNA
C0485405|T201|COMP|10677-3|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C0485406|T201|COMP|10678-1|LNC|Herpes simplex virus 1+2 Ag|Herpes simplex virus 1+2 Ag
C0485407|T201|COMP|10679-9|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C0485408|T201|COMP|10680-7|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C0485409|T201|COMP|10681-5|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C0485410|T201|COMP|9454-0|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C0485411|T201|COMP|7907-9|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C0485412|T201|COMP|9659-4|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C0485413|T201|COMP|9422-7|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C0485414|T201|COMP|10350-7|LNC|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C0485415|T201|COMP|7908-7|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C0485416|T201|COMP|7909-5|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C0485417|T201|COMP|7910-3|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C0485418|T201|COMP|7911-1|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C0485419|T201|COMP|7912-9|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0485420|T201|COMP|7913-7|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C0485421|T201|COMP|7914-5|LNC|Heterophile Ab after beef cell absorption|Heterophile Ab after beef cell absorption
C0485422|T201|COMP|7915-2|LNC|Heterophile Ab after guinea pig cell absorption|Heterophile Ab after guinea pig cell absorption
C0485423|T201|COMP|7916-0|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0485424|T201|COMP|9528-1|LNC|Histoplasma capsulatum Ab.IgA|Histoplasma capsulatum Ab.IgA
C0485425|T201|COMP|9529-9|LNC|Histoplasma capsulatum Ab.IgG|Histoplasma capsulatum Ab.IgG
C0485426|T201|COMP|9530-7|LNC|Histoplasma capsulatum Ab.IgM|Histoplasma capsulatum Ab.IgM
C0485427|T201|COMP|6816-3|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C0485428|T201|COMP|6817-1|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C0485429|T201|COMP|7917-8|LNC|HIV 1 Ab|HIV 1 Ab
C0485430|T201|COMP|9837-6|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C0485431|T201|COMP|9661-0|LNC|HIV 1 gp120 Ab|HIV 1 gp120 Ab
C0485432|T201|COMP|9660-2|LNC|HIV 1 gp160 Ab|HIV 1 gp160 Ab
C0485433|T201|COMP|9662-8|LNC|HIV 1 gp41 Ab|HIV 1 gp41 Ab
C0485434|T201|COMP|9663-6|LNC|HIV 1 p17 Ab|HIV 1 p17 Ab
C0485435|T201|COMP|9664-4|LNC|HIV 1 p24 Ab|HIV 1 p24 Ab
C0485436|T201|COMP|9665-1|LNC|HIV 1 p24 Ag|HIV 1 p24 Ag
C0485437|T201|COMP|9821-0|LNC|HIV 1 p24 Ag|HIV 1 p24 Ag
C0485438|T201|COMP|9666-9|LNC|HIV 1 p31 Ab|HIV 1 p31 Ab
C0485439|T201|COMP|9667-7|LNC|HIV 1 p51 Ab|HIV 1 p51 Ab
C0485440|T201|COMP|9668-5|LNC|HIV 1 p55 Ab|HIV 1 p55 Ab
C0485441|T201|COMP|9669-3|LNC|HIV 1 p66 Ab|HIV 1 p66 Ab
C0485443|T201|COMP|10351-5|LNC|HIV 1 RNA|HIV 1 RNA
C0485444|T201|COMP|7918-6|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C0485445|T201|COMP|7919-4|LNC|HIV 2 Ab|HIV 2 Ab
C0485446|T201|COMP|9836-8|LNC|HIV proviral DNA|HIV proviral DNA
C0485447|T201|COMP|10683-1|LNC|Hydatid cyst identified|Hydatid cyst identified
C0485448|T201|COMP|10684-9|LNC|Hydatid cyst identified|Hydatid cyst identified
C0485449|T201|COMP|10685-6|LNC|Hydatid cyst identified|Hydatid cyst identified
C0485450|T201|COMP|9531-5|LNC|Influenza virus A Ab|Influenza virus A Ab
C0485451|T201|COMP|7920-2|LNC|Influenza virus A Ab|Influenza virus A Ab
C0485452|T201|COMP|9532-3|LNC|Influenza virus A Ab.IgG|Influenza virus A Ab.IgG
C0485453|T201|COMP|9533-1|LNC|Influenza virus A Ab.IgM|Influenza virus A Ab.IgM
C0485454|T201|COMP|6639-9|LNC|Influenza virus A Bangkok Ab|Influenza virus A Bangkok Ab
C0485455|T201|COMP|7921-0|LNC|Influenza virus A Bangkok Ab|Influenza virus A Bangkok Ab
C0485456|T201|COMP|6635-7|LNC|Influenza virus A England Ab|Influenza virus A England Ab
C0485457|T201|COMP|7922-8|LNC|Influenza virus A England Ab|Influenza virus A England Ab
C0485458|T201|COMP|6634-0|LNC|Influenza virus A Hong Kong Ab|Influenza virus A Hong Kong Ab
C0485459|T201|COMP|7923-6|LNC|Influenza virus A Hong Kong Ab|Influenza virus A Hong Kong Ab
C0485460|T201|COMP|6642-3|LNC|Influenza virus A Leningrad Ab|Influenza virus A Leningrad Ab
C0485461|T201|COMP|7924-4|LNC|Influenza virus A Leningrad Ab|Influenza virus A Leningrad Ab
C0485462|T201|COMP|6641-5|LNC|Influenza virus A Mississippi Ab|Influenza virus A Mississippi Ab
C0485463|T201|COMP|7925-1|LNC|Influenza virus A Mississippi Ab|Influenza virus A Mississippi Ab
C0485464|T201|COMP|6640-7|LNC|Influenza virus A Phillipines Ab|Influenza virus A Phillipines Ab
C0485465|T201|COMP|7926-9|LNC|Influenza virus A Phillipines Ab|Influenza virus A Phillipines Ab
C0485466|T201|COMP|6636-5|LNC|Influenza virus A Port Chalmers Ab|Influenza virus A Port Chalmers Ab
C0485467|T201|COMP|7927-7|LNC|Influenza virus A Port Chalmers Ab|Influenza virus A Port Chalmers Ab
C0485468|T201|COMP|6638-1|LNC|Influenza virus A Texas Ab|Influenza virus A Texas Ab
C0485469|T201|COMP|7928-5|LNC|Influenza virus A Texas Ab|Influenza virus A Texas Ab
C0485470|T201|COMP|6637-3|LNC|Influenza virus A Victoria Ab|Influenza virus A Victoria Ab
C0485471|T201|COMP|7929-3|LNC|Influenza virus A Victoria Ab|Influenza virus A Victoria Ab
C0485472|T201|COMP|7930-1|LNC|Influenza virus A+B Ab|Influenza virus A+B Ab
C0485473|T201|COMP|9534-9|LNC|Influenza virus B Ab|Influenza virus B Ab
C0485474|T201|COMP|7931-9|LNC|Influenza virus B Ab|Influenza virus B Ab
C0485475|T201|COMP|9535-6|LNC|Influenza virus B Ab.IgG|Influenza virus B Ab.IgG
C0485476|T201|COMP|9536-4|LNC|Influenza virus B Ab.IgM|Influenza virus B Ab.IgM
C0485477|T201|COMP|7932-7|LNC|Influenza virus C Ab|Influenza virus C Ab
C0485478|T201|COMP|6601-9|LNC|Influenza virus identified|Influenza virus identified
C0485479|T201|COMP|6602-7|LNC|Influenza virus identified|Influenza virus identified
C0485480|T201|COMP|6603-5|LNC|Influenza virus identified|Influenza virus identified
C0485481|T201|COMP|6604-3|LNC|Influenza virus identified|Influenza virus identified
C0485482|T201|COMP|7933-5|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0485483|T201|COMP|7935-0|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0485484|T201|COMP|7934-3|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0485485|T201|COMP|7936-8|LNC|Japanese encephalitis virus RNA|Japanese encephalitis virus RNA
C0485486|T201|COMP|7937-6|LNC|Junin virus Ab|Junin virus Ab
C0485487|T201|COMP|9538-0|LNC|La Crosse virus Ab|La Crosse virus Ab
C0485488|T201|COMP|7938-4|LNC|La Crosse virus Ab|La Crosse virus Ab
C0485489|T201|COMP|7939-2|LNC|La Crosse virus Ab|La Crosse virus Ab
C0485490|T201|COMP|9539-8|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C0485491|T201|COMP|7940-0|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C0485492|T201|COMP|9540-6|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C0485493|T201|COMP|7941-8|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C0485494|T201|COMP|7942-6|LNC|Lassa virus Ab.IgG|Lassa virus Ab.IgG
C0485495|T201|COMP|7943-4|LNC|Lassa virus Ab.IgG|Lassa virus Ab.IgG
C0485496|T201|COMP|7944-2|LNC|Lassa virus Ab.IgM|Lassa virus Ab.IgM
C0485497|T201|COMP|7945-9|LNC|Lassa virus Ab.IgM|Lassa virus Ab.IgM
C0485498|T201|COMP|7946-7|LNC|Lassa virus Ag|Lassa virus Ag
C0485499|T201|COMP|7947-5|LNC|Legionella pneumophila Ab|Legionella pneumophila Ab
C0485500|T201|COMP|7948-3|LNC|Legionella pneumophila 1 Ab|Legionella pneumophila 1 Ab
C0485501|T201|COMP|9541-4|LNC|Legionella pneumophila 1 Ab.IgG|Legionella pneumophila 1 Ab.IgG
C0485502|T201|COMP|9542-2|LNC|Legionella pneumophila 1 Ab.IgM|Legionella pneumophila 1 Ab.IgM
C0485503|T201|COMP|9543-0|LNC|Legionella pneumophila 1 Ag|Legionella pneumophila 1 Ag
C0485504|T201|COMP|7949-1|LNC|Legionella pneumophila 2 Ab|Legionella pneumophila 2 Ab
C0485505|T201|COMP|9544-8|LNC|Legionella pneumophila 2 Ab.IgG|Legionella pneumophila 2 Ab.IgG
C0485506|T201|COMP|9545-5|LNC|Legionella pneumophila 2 Ab.IgM|Legionella pneumophila 2 Ab.IgM
C0485507|T201|COMP|7950-9|LNC|Legionella pneumophila 3 Ab|Legionella pneumophila 3 Ab
C0485508|T201|COMP|9546-3|LNC|Legionella pneumophila 3 Ab.IgG|Legionella pneumophila 3 Ab.IgG
C0485509|T201|COMP|9547-1|LNC|Legionella pneumophila 3 Ab.IgM|Legionella pneumophila 3 Ab.IgM
C0485510|T201|COMP|7951-7|LNC|Legionella pneumophila 4 Ab|Legionella pneumophila 4 Ab
C0485511|T201|COMP|9548-9|LNC|Legionella pneumophila 4 Ab.IgG|Legionella pneumophila 4 Ab.IgG
C0485512|T201|COMP|9549-7|LNC|Legionella pneumophila 4 Ab.IgM|Legionella pneumophila 4 Ab.IgM
C0485513|T201|COMP|7952-5|LNC|Legionella pneumophila 5 Ab|Legionella pneumophila 5 Ab
C0485514|T201|COMP|9550-5|LNC|Legionella pneumophila 5 Ab.IgG|Legionella pneumophila 5 Ab.IgG
C0485515|T201|COMP|9551-3|LNC|Legionella pneumophila 5 Ab.IgM|Legionella pneumophila 5 Ab.IgM
C0485516|T201|COMP|7953-3|LNC|Legionella pneumophila 6 Ab|Legionella pneumophila 6 Ab
C0485517|T201|COMP|9552-1|LNC|Legionella pneumophila 6 Ab.IgG|Legionella pneumophila 6 Ab.IgG
C0485518|T201|COMP|9553-9|LNC|Legionella pneumophila 6 Ab.IgM|Legionella pneumophila 6 Ab.IgM
C0485519|T201|COMP|7954-1|LNC|Legionella pneumophila 7 Ab|Legionella pneumophila 7 Ab
C0485520|T201|COMP|7955-8|LNC|Legionella pneumophila 8 Ab|Legionella pneumophila 8 Ab
C0485521|T201|COMP|7956-6|LNC|Legionella pneumophila 9 Ab|Legionella pneumophila 9 Ab
C0485522|T201|COMP|7957-4|LNC|Legionella sp Ab|Legionella sp Ab
C0485523|T201|COMP|10686-4|LNC|Leishmania sp identified|Leishmania sp identified
C0485524|T201|COMP|10687-2|LNC|Leishmania sp identified|Leishmania sp identified
C0485525|T201|COMP|6621-7|LNC|Leishmania sp Ab|Leishmania sp Ab
C0485526|T201|COMP|6622-5|LNC|Leishmania sp Ab|Leishmania sp Ab
C0485527|T201|COMP|6623-3|LNC|Leishmania sp Ab|Leishmania sp Ab
C0485528|T201|COMP|7958-2|LNC|Leishmania sp Ab|Leishmania sp Ab
C0485529|T201|COMP|7959-0|LNC|Leptospira sp Ab|Leptospira sp Ab
C0485530|T201|COMP|7960-8|LNC|Leptospira interrogans Ab|Leptospira interrogans Ab
C0485531|T201|COMP|6605-0|LNC|Leptospira interrogans Ag|Leptospira interrogans Ag
C0485532|T201|COMP|6609-2|LNC|Listeria sp identified|Listeria sp identified
C0485533|T201|COMP|9564-6|LNC|Lymphocytic choriomeningitis virus Ab|Lymphocytic choriomeningitis virus Ab
C0485534|T201|COMP|9766-7|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C0485535|T201|COMP|9765-9|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C0485536|T201|COMP|9768-3|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C0485537|T201|COMP|9767-5|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C0485538|T201|COMP|9565-3|LNC|Measles virus Ab|Measles virus Ab
C0485539|T201|COMP|7961-6|LNC|Measles virus Ab|Measles virus Ab
C0485540|T201|COMP|9566-1|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0485541|T201|COMP|7962-4|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0485542|T201|COMP|7963-2|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C0485543|T201|COMP|7964-0|LNC|Measles virus RNA|Measles virus RNA
C0485544|T201|COMP|9822-8|LNC|Bacteria identified|Bacteria identified
C0485545|T201|COMP|17887-1|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0485546|T201|COMP|17892-1|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0485547|T201|COMP|10354-9|LNC|Bacteria identified|Bacteria identified
C0485548|T201|COMP|6818-9|LNC|Saccharopolyspora rectivirgula Ab|Saccharopolyspora rectivirgula Ab
C0485573|T201|COMP|6674-6|LNC|Ova & parasites identified|Ova & parasites identified
C0485575|T201|COMP|6676-1|LNC|Enterobius vermicularis|Enterobius vermicularis
C0485581|T201|COMP|10690-6|LNC|Microsporidia identified|Microsporidia identified
C0485582|T201|COMP|9567-9|LNC|Mumps virus Ab|Mumps virus Ab
C0485583|T201|COMP|7965-7|LNC|Mumps virus Ab|Mumps virus Ab
C0485584|T201|COMP|7966-5|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0485585|T201|COMP|7967-3|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C0485586|T201|COMP|7968-1|LNC|Mumps virus RNA|Mumps virus RNA
C0485587|T201|COMP|10692-2|LNC|Mushroom.toxic identified|Mushroom.toxic identified
C0485588|T201|COMP|10693-0|LNC|Mushroom.toxic identified|Mushroom.toxic identified
C0485589|T201|COMP|10691-4|LNC|Mushroom.toxic identified|Mushroom.toxic identified
C0485590|T201|COMP|9823-6|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0485591|T201|COMP|9824-4|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0485592|T201|COMP|9825-1|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C0485593|T201|COMP|7969-9|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C0485594|T201|COMP|7970-7|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C0485595|T201|COMP|6624-1|LNC|Naegleria fowleri Ab|Naegleria fowleri Ab
C0485596|T201|COMP|6625-8|LNC|Naegleria fowleri Ab|Naegleria fowleri Ab
C0485597|T201|COMP|7971-5|LNC|Naegleria fowleri Ab|Naegleria fowleri Ab
C0485598|T201|COMP|10694-8|LNC|Naegleria sp identified|Naegleria sp identified
C0485599|T201|COMP|10695-5|LNC|Naegleria sp identified|Naegleria sp identified
C0485600|T201|COMP|9568-7|LNC|Neisseria gonorrhoeae Ab|Neisseria gonorrhoeae Ab
C0485601|T201|COMP|7972-3|LNC|Neisseria meningitidis serogroup Y Ab|Neisseria meningitidis serogroup Y Ab
C0485602|T201|COMP|9569-5|LNC|Nocardia sp Ab.IgG|Nocardia sp Ab.IgG
C0485603|T201|COMP|7973-1|LNC|Norovirus|Norovirus
C0485604|T201|COMP|10696-3|LNC|Norovirus|Norovirus
C0485605|T201|COMP|7974-9|LNC|Norovirus RNA|Norovirus RNA
C0485606|T201|COMP|10697-1|LNC|Nystatin|Nystatin
C0485607|T201|COMP|10698-9|LNC|Nystatin|Nystatin
C0485608|T201|COMP|10699-7|LNC|Onchocerca sp identified|Onchocerca sp identified
C0485609|T201|COMP|10700-3|LNC|Orthopoxvirus|Orthopoxvirus
C0485610|T201|COMP|10701-1|LNC|Ova & parasites identified|Ova & parasites identified
C0485611|T201|COMP|10702-9|LNC|Ova & parasites identified|Ova & parasites identified
C0485612|T201|COMP|10703-7|LNC|Ova & parasites identified|Ova & parasites identified
C0485613|T201|COMP|10704-5|LNC|Ova & parasites identified|Ova & parasites identified
C0485614|T201|COMP|7975-6|LNC|Human papilloma virus Ab|Human papilloma virus Ab
C0485615|T201|COMP|10705-2|LNC|Human papilloma virus Ag|Human papilloma virus Ag
C0485616|T201|COMP|7976-4|LNC|Paracoccidioides brasiliensis Ab|Paracoccidioides brasiliensis Ab
C0485617|T201|COMP|7977-2|LNC|Paragonimus sp Ab|Paragonimus sp Ab
C0485618|T201|COMP|7978-0|LNC|Parainfluenza virus 1 Ab|Parainfluenza virus 1 Ab
C0485619|T201|COMP|7979-8|LNC|Parainfluenza virus 2 Ab|Parainfluenza virus 2 Ab
C0485620|T201|COMP|7980-6|LNC|Parainfluenza virus 3 Ab|Parainfluenza virus 3 Ab
C0485621|T201|COMP|7981-4|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0485622|T201|COMP|7982-2|LNC|Parvovirus B19 Ab|Parvovirus B19 Ab
C0485623|T201|COMP|7983-0|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0485624|T201|COMP|7984-8|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0485625|T201|COMP|9572-9|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C0485626|T201|COMP|9571-1|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C0485627|T201|COMP|10706-0|LNC|Picornavirus|Picornavirus
C0485628|T201|COMP|10708-6|LNC|Plant.toxic identified|Plant.toxic identified
C0485629|T201|COMP|10707-8|LNC|Plant.toxic identified|Plant.toxic identified
C0485630|T201|COMP|10709-4|LNC|Plasmodium falciparum Ag|Plasmodium falciparum Ag
C0485631|T201|COMP|9670-1|LNC|Plasmodium malariae Ab.IgG|Plasmodium malariae Ab.IgG
C0485632|T201|COMP|9671-9|LNC|Plasmodium malariae Ab.IgM|Plasmodium malariae Ab.IgM
C0485633|T201|COMP|10710-2|LNC|Plasmodium sp identified|Plasmodium sp identified
C0485634|T201|COMP|10711-0|LNC|Plasmodium vivax Ag|Plasmodium vivax Ag
C0485635|T201|COMP|10712-8|LNC|Pneumocystis sp identified|Pneumocystis sp identified
C0485636|T201|COMP|7985-5|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C0485637|T201|COMP|7986-3|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C0485638|T201|COMP|7987-1|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C0485639|T201|COMP|10713-6|LNC|Prototheca identified|Prototheca identified
C0485640|T201|COMP|7988-9|LNC|Burkholderia pseudomallei Ab.IgG|Burkholderia pseudomallei Ab.IgG
C0485641|T201|COMP|7989-7|LNC|Burkholderia pseudomallei Ab.IgM|Burkholderia pseudomallei Ab.IgM
C0485642|T201|COMP|7990-5|LNC|Respiratory syncytial virus Ab|Respiratory syncytial virus Ab
C0485643|T201|COMP|7991-3|LNC|Respiratory syncytial virus Ab.IgG|Respiratory syncytial virus Ab.IgG
C0485644|T201|COMP|9573-7|LNC|Respiratory syncytial virus Ab.IgG|Respiratory syncytial virus Ab.IgG
C0485645|T201|COMP|7992-1|LNC|Respiratory syncytial virus Ab.IgM|Respiratory syncytial virus Ab.IgM
C0485646|T201|COMP|9574-5|LNC|Respiratory syncytial virus Ab.IgM|Respiratory syncytial virus Ab.IgM
C0485647|T201|COMP|7993-9|LNC|Rhinovirus RNA|Rhinovirus RNA
C0485648|T201|COMP|7994-7|LNC|Rickettsia sp Ab|Rickettsia sp Ab
C0485649|T201|COMP|7995-4|LNC|Rickettsia prowazekii Ab|Rickettsia prowazekii Ab
C0485650|T201|COMP|7996-2|LNC|Rickettsia prowazekii RNA|Rickettsia prowazekii RNA
C0485651|T201|COMP|7997-0|LNC|Rickettsia spotted fever group Ab|Rickettsia spotted fever group Ab
C0485652|T201|COMP|7998-8|LNC|Rickettsia spotted fever group Ab.IgG|Rickettsia spotted fever group Ab.IgG
C0485653|T201|COMP|7999-6|LNC|Rickettsia spotted fever group Ab.IgM|Rickettsia spotted fever group Ab.IgM
C0485654|T201|COMP|8000-2|LNC|Rickettsia typhus group Ab|Rickettsia typhus group Ab
C0485655|T201|COMP|8001-0|LNC|Rickettsia typhus group Ab.IgG|Rickettsia typhus group Ab.IgG
C0485656|T201|COMP|8002-8|LNC|Rickettsia typhus group Ab.IgM|Rickettsia typhus group Ab.IgM
C0485657|T201|COMP|8003-6|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C0485658|T201|COMP|8004-4|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C0485659|T201|COMP|8005-1|LNC|Rickettsia rickettsii RNA|Rickettsia rickettsii RNA
C0485660|T201|COMP|8006-9|LNC|Orientia tsutsugamushi Ab|Orientia tsutsugamushi Ab
C0485661|T201|COMP|8007-7|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C0485662|T201|COMP|8008-5|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C0485663|T201|COMP|8011-9|LNC|Rotavirus|Rotavirus
C0485664|T201|COMP|10714-4|LNC|Rotavirus|Rotavirus
C0485665|T201|COMP|9575-2|LNC|Rotavirus Ab|Rotavirus Ab
C0485666|T201|COMP|8012-7|LNC|Rotavirus dsRNA|Rotavirus dsRNA
C0485667|T201|COMP|9576-0|LNC|Rubella virus Ab|Rubella virus Ab
C0485668|T201|COMP|8013-5|LNC|Rubella virus Ab|Rubella virus Ab
C0485669|T201|COMP|8014-3|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0485670|T201|COMP|8015-0|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C0485671|T201|COMP|8021-8|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0485672|T201|COMP|9577-8|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0485673|T201|COMP|8022-6|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0485674|T201|COMP|8023-4|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0485675|T201|COMP|8024-2|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0485676|T201|COMP|9578-6|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0485677|T201|COMP|8016-8|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C0485678|T201|COMP|9634-7|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C0485679|T201|COMP|8017-6|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C0485680|T201|COMP|9635-4|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C0485681|T201|COMP|8025-9|LNC|Saint Louis encephalitis virus RNA|Saint Louis encephalitis virus RNA
C0485682|T201|COMP|9672-7|LNC|Salmonella sp Ab.IgA|Salmonella sp Ab.IgA
C0485683|T201|COMP|9673-5|LNC|Salmonella sp Ab.IgG|Salmonella sp Ab.IgG
C0485684|T201|COMP|9674-3|LNC|Salmonella sp Ab.IgM|Salmonella sp Ab.IgM
C0485685|T201|COMP|9787-3|LNC|Sarcoptes scabiei identified|Sarcoptes scabiei identified
C0485686|T201|COMP|8018-4|LNC|Schistosoma japonicum Ab|Schistosoma japonicum Ab
C0485687|T201|COMP|6626-6|LNC|Schistosoma japonicum Ab|Schistosoma japonicum Ab
C0485688|T201|COMP|8019-2|LNC|Schistosoma mansoni Ab|Schistosoma mansoni Ab
C0485689|T201|COMP|6627-4|LNC|Schistosoma mansoni Ab|Schistosoma mansoni Ab
C0485690|T201|COMP|6628-2|LNC|Schistosoma sp Ab|Schistosoma sp Ab
C0485691|T201|COMP|6629-0|LNC|Schistosoma sp Ab|Schistosoma sp Ab
C0485692|T201|COMP|6630-8|LNC|Schistosoma sp Ab|Schistosoma sp Ab
C0485693|T201|COMP|6631-6|LNC|Schistosoma sp Ab|Schistosoma sp Ab
C0485694|T201|COMP|8020-0|LNC|Schistosoma sp Ab|Schistosoma sp Ab
C0485695|T201|COMP|10715-1|LNC|Schistosoma sp identified|Schistosoma sp identified
C0485696|T201|COMP|10716-9|LNC|Schistosoma sp identified|Schistosoma sp identified
C0485697|T201|COMP|9712-1|LNC|Shigella boydii Ab|Shigella boydii Ab
C0485698|T201|COMP|9713-9|LNC|Shigella dysenteriae Ab|Shigella dysenteriae Ab
C0485699|T201|COMP|9714-7|LNC|Shigella flexneri Ab|Shigella flexneri Ab
C0485700|T201|COMP|9715-4|LNC|Shigella sonnei Ab|Shigella sonnei Ab
C0485701|T201|COMP|8026-7|LNC|Stain method|Stain method
C0485702|T201|COMP|9716-2|LNC|Streptococcal hyaluronidase Ab|Streptococcal hyaluronidase Ab
C0485703|T201|COMP|6819-7|LNC|Streptococcus sp Ab|Streptococcus sp Ab
C0485704|T201|COMP|6820-5|LNC|Streptococcus sp Ab|Streptococcus sp Ab
C0485705|T201|COMP|9455-7|LNC|Streptococcus pneumoniae 1 Ab.IgG|Streptococcus pneumoniae 1 Ab.IgG
C0485706|T201|COMP|9456-5|LNC|Streptococcus pneumoniae 12 Ab.IgG|Streptococcus pneumoniae 12 Ab.IgG
C0485707|T201|COMP|8027-5|LNC|Streptococcus pneumoniae 14 Ab.IgG|Streptococcus pneumoniae 14 Ab.IgG
C0485708|T201|COMP|9457-3|LNC|Streptococcus pneumoniae 19 Ab.IgG|Streptococcus pneumoniae 19 Ab.IgG
C0485709|T201|COMP|9458-1|LNC|Streptococcus pneumoniae 23 Ab.IgG|Streptococcus pneumoniae 23 Ab.IgG
C0485710|T201|COMP|8033-3|LNC|Streptococcus pneumoniae 3 Ab.IgG|Streptococcus pneumoniae 3 Ab.IgG
C0485711|T201|COMP|9459-9|LNC|Streptococcus pneumoniae 4 Ab.IgG|Streptococcus pneumoniae 4 Ab.IgG
C0485713|T201|COMP|9460-7|LNC|Streptococcus pneumoniae 6+26 Ab.IgG|Streptococcus pneumoniae 6+26 Ab.IgG
C0485715|T201|COMP|9461-5|LNC|Streptococcus pneumoniae 8 Ab.IgG|Streptococcus pneumoniae 8 Ab.IgG
C0485716|T201|COMP|8029-1|LNC|Streptococcus pneumoniae 9 Ab.IgG|Streptococcus pneumoniae 9 Ab.IgG
C0485717|T201|COMP|10717-7|LNC|Streptococcus pneumoniae Ab|Streptococcus pneumoniae Ab
C0485718|T201|COMP|8030-9|LNC|Streptococcus pneumoniae Ab|Streptococcus pneumoniae Ab
C0485719|T201|COMP|8031-7|LNC|Streptococcus pneumoniae Ab.IgG|Streptococcus pneumoniae Ab.IgG
C0485720|T201|COMP|8032-5|LNC|Streptococcus pneumoniae Ab.IgM|Streptococcus pneumoniae Ab.IgM
C0485721|T201|COMP|9788-1|LNC|Streptolysin O Ab|Streptolysin O Ab
C0485722|T201|COMP|8034-1|LNC|Strongyloides sp Ab|Strongyloides sp Ab
C0485723|T201|COMP|10718-5|LNC|Strongyloides sp Ab|Strongyloides sp Ab
C0485724|T201|COMP|6632-4|LNC|Strongyloides stercoralis Ab.IgG|Strongyloides stercoralis Ab.IgG
C0485725|T201|COMP|8035-8|LNC|Strongyloides stercoralis Ab.IgG|Strongyloides stercoralis Ab.IgG
C0485726|T201|COMP|8036-6|LNC|Taenia saginata Ab|Taenia saginata Ab
C0485727|T201|COMP|8037-4|LNC|Taenia solium adult Ab|Taenia solium adult Ab
C0485728|T201|COMP|10719-3|LNC|Taenia solium adult Ab|Taenia solium adult Ab
C0485729|T201|COMP|10358-0|LNC|Teichoate Ab|Teichoate Ab
C0485730|T201|COMP|10720-1|LNC|Terbinafine|Terbinafine
C0485731|T201|COMP|10721-9|LNC|Terbinafine|Terbinafine
C0485732|T201|COMP|9769-1|LNC|Thermoactinomyces candidus Ab|Thermoactinomyces candidus Ab
C0485733|T201|COMP|9770-9|LNC|Thermoactinomyces sacchari Ab|Thermoactinomyces sacchari Ab
C0485734|T201|COMP|6821-3|LNC|Thermoactinomyces vulgaris Ab|Thermoactinomyces vulgaris Ab
C0485735|T201|COMP|10722-7|LNC|Torovirus|Torovirus
C0485736|T201|COMP|8038-2|LNC|Toxocara canis Ab|Toxocara canis Ab
C0485737|T201|COMP|9717-0|LNC|Toxocara canis Ab.IgA|Toxocara canis Ab.IgA
C0485738|T201|COMP|9718-8|LNC|Toxocara canis Ab.IgG|Toxocara canis Ab.IgG
C0485739|T201|COMP|9719-6|LNC|Toxocara canis Ab.IgM|Toxocara canis Ab.IgM
C0485740|T201|COMP|10723-5|LNC|Toxoplasma gondii Ab.IgA|Toxoplasma gondii Ab.IgA
C0485741|T201|COMP|10724-3|LNC|Toxoplasma gondii Ab.IgE|Toxoplasma gondii Ab.IgE
C0485742|T201|COMP|8039-0|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0485743|T201|COMP|8040-8|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0485744|T201|COMP|10725-0|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C0485745|T201|COMP|9741-0|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0485746|T201|COMP|10726-8|LNC|Toxoplasma gondii|Toxoplasma gondii
C0485747|T201|COMP|10727-6|LNC|Toxoplasma gondii identified|Toxoplasma gondii identified
C0485748|T201|COMP|9826-9|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0485749|T201|COMP|8041-6|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0485750|T201|COMP|8042-4|LNC|Trichinella spiralis Ab|Trichinella spiralis Ab
C0485751|T201|COMP|8043-2|LNC|Trichinella spiralis Ab.IgG|Trichinella spiralis Ab.IgG
C0485752|T201|COMP|10728-4|LNC|Trichomonas sp identified|Trichomonas sp identified
C0485753|T201|COMP|8045-7|LNC|Trypanosoma cruzi Ab|Trypanosoma cruzi Ab
C0485754|T201|COMP|10729-2|LNC|Trypanosoma sp identified|Trypanosoma sp identified
C0485755|T201|COMP|10730-0|LNC|Trypanosoma sp identified|Trypanosoma sp identified
C0485756|T201|COMP|10731-8|LNC|Trypanosoma sp identified|Trypanosoma sp identified
C0485757|T201|COMP|10732-6|LNC|Trypanosoma sp identified|Trypanosoma sp identified
C0485758|T201|COMP|10733-4|LNC|Trypanosoma sp identified|Trypanosoma sp identified
C0485759|T201|COMP|9636-2|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C0485760|T201|COMP|8046-5|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C0485761|T201|COMP|8047-3|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0485762|T201|COMP|8048-1|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0485763|T201|COMP|8049-9|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C0485764|T201|COMP|10734-2|LNC|Varicella zoster virus identified|Varicella zoster virus identified
C0485765|T201|COMP|8050-7|LNC|Venezuelan equine encephalitis virus Ab.IgG|Venezuelan equine encephalitis virus Ab.IgG
C0485766|T201|COMP|8051-5|LNC|Venezuelan equine encephalitis virus Ab.IgM|Venezuelan equine encephalitis virus Ab.IgM
C0485767|T201|COMP|10735-9|LNC|Viral sequencing|Viral sequencing
C0485768|T201|COMP|10736-7|LNC|Virus identified|Virus identified
C0485769|T201|COMP|6608-4|LNC|Virus identified|Virus identified
C0485770|T201|COMP|10737-5|LNC|Virus identified|Virus identified
C0485771|T201|COMP|10738-3|LNC|Virus identified|Virus identified
C0485772|T201|COMP|10739-1|LNC|Virus identified|Virus identified
C0485773|T201|COMP|9314-6|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0485774|T201|COMP|9581-0|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0485775|T201|COMP|9315-3|LNC|Western equine encephalitis virus Ab.IgG|Western equine encephalitis virus Ab.IgG
C0485776|T201|COMP|8052-3|LNC|Western equine encephalitis virus Ab.IgG|Western equine encephalitis virus Ab.IgG
C0485777|T201|COMP|6957-5|LNC|Western equine encephalitis virus Ab.IgG|Western equine encephalitis virus Ab.IgG
C0485778|T201|COMP|9316-1|LNC|Western equine encephalitis virus Ab.IgM|Western equine encephalitis virus Ab.IgM
C0485779|T201|COMP|8053-1|LNC|Western equine encephalitis virus Ab.IgM|Western equine encephalitis virus Ab.IgM
C0485780|T201|COMP|6958-3|LNC|Western equine encephalitis virus Ab.IgM|Western equine encephalitis virus Ab.IgM
C0485781|T201|COMP|6633-2|LNC|Wuchereria bancrofti Ab|Wuchereria bancrofti Ab
C0485782|T201|COMP|8054-9|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C0485783|T201|COMP|8055-6|LNC|Yellow fever virus Ab.IgG|Yellow fever virus Ab.IgG
C0485784|T201|COMP|8056-4|LNC|Yellow fever virus Ab.IgM|Yellow fever virus Ab.IgM
C0485785|T201|COMP|8057-2|LNC|Yellow fever virus RNA|Yellow fever virus RNA
C0485786|T201|COMP|6959-1|LNC|Yersinia enterocolitica O:3 Ab|Yersinia enterocolitica O:3 Ab
C0485787|T201|COMP|6960-9|LNC|Yersinia enterocolitica O:5 Ab|Yersinia enterocolitica O:5 Ab
C0485788|T201|COMP|6961-7|LNC|Yersinia enterocolitica O:8 Ab|Yersinia enterocolitica O:8 Ab
C0485789|T201|COMP|6962-5|LNC|Yersinia enterocolitica O:9 Ab|Yersinia enterocolitica O:9 Ab
C0485790|T201|COMP|6963-3|LNC|Yersinia enterocolitica Ab|Yersinia enterocolitica Ab
C0485791|T201|COMP|6964-1|LNC|Yersinia enterocolitica Ab.IgA|Yersinia enterocolitica Ab.IgA
C0485792|T201|COMP|6965-8|LNC|Yersinia enterocolitica Ab.IgG|Yersinia enterocolitica Ab.IgG
C0485793|T201|COMP|6966-6|LNC|Yersinia enterocolitica Ab.IgM|Yersinia enterocolitica Ab.IgM
C0485794|T201|COMP|6967-4|LNC|Yersinia pseudotuberculosis Ab|Yersinia pseudotuberculosis Ab
C0485795|T201|COMP|8251-1|LNC|Service comment|Service comment
C0485796|T201|COMP|8252-9|LNC|Service comment 10|Service comment 10
C0485797|T201|COMP|8253-7|LNC|Service comment 11|Service comment 11
C0485798|T201|COMP|8254-5|LNC|Service comment 12|Service comment 12
C0485799|T201|COMP|8255-2|LNC|Service comment 13|Service comment 13
C0485800|T201|COMP|8256-0|LNC|Service comment 14|Service comment 14
C0485801|T201|COMP|8257-8|LNC|Service comment 15|Service comment 15
C0485802|T201|COMP|8258-6|LNC|Service comment 16|Service comment 16
C0485803|T201|COMP|8259-4|LNC|Service comment 17|Service comment 17
C0485804|T201|COMP|8260-2|LNC|Service comment 18|Service comment 18
C0485805|T201|COMP|8261-0|LNC|Service comment 19|Service comment 19
C0485806|T201|COMP|8262-8|LNC|Service comment 02|Service comment 02
C0485807|T201|COMP|8263-6|LNC|Service comment 20|Service comment 20
C0485808|T201|COMP|8264-4|LNC|Service comment 03|Service comment 03
C0485809|T201|COMP|8265-1|LNC|Service comment 04|Service comment 04
C0485810|T201|COMP|8266-9|LNC|Service comment 05|Service comment 05
C0485811|T201|COMP|8267-7|LNC|Service comment 06|Service comment 06
C0485812|T201|COMP|8268-5|LNC|Service comment 07|Service comment 07
C0485813|T201|COMP|8269-3|LNC|Service comment 08|Service comment 08
C0485814|T201|COMP|8270-1|LNC|Service comment 09|Service comment 09
C0485815|T201|COMP|9796-4|LNC|Color|Color
C0485816|T201|COMP|9795-6|LNC|Composition|Composition
C0485817|T201|COMP|9797-2|LNC|Consistency|Consistency
C0485818|T201|COMP|9798-0|LNC|Depth|Depth
C0485819|T201|COMP|9799-8|LNC|Length|Length
C0485820|T201|COMP|9800-4|LNC|Number|Number
C0485821|T201|COMP|9801-2|LNC|Shape|Shape
C0485822|T201|COMP|9802-0|LNC|Size|Size
C0485823|T201|COMP|9803-8|LNC|Texture|Texture
C0485824|T201|COMP|9804-6|LNC|Weight|Weight
C0485825|T201|COMP|9805-3|LNC|Width|Width
C0485826|T201|COMP|9326-0|LNC|Phosphatidylserine Ab.IgG|Phosphatidylserine Ab.IgG
C0485827|T201|COMP|9327-8|LNC|Phosphatidylserine Ab.IgM|Phosphatidylserine Ab.IgM
C0485828|T201|COMP|8058-0|LNC|Acetylcholine receptor Ab|Acetylcholine receptor Ab
C0485829|T201|COMP|8059-8|LNC|Adrenal Ab|Adrenal Ab
C0485830|T201|COMP|6923-7|LNC|Adrenal cortex Ab|Adrenal cortex Ab
C0485831|T201|COMP|8060-6|LNC|Adrenal cortex Ab|Adrenal cortex Ab
C0485832|T201|COMP|8061-4|LNC|Nuclear Ab|Nuclear Ab
C0485833|T201|COMP|6822-1|LNC|Nuclear Ab|Nuclear Ab
C0485834|T201|COMP|10359-8|LNC|Asialoganglioside GM1 Ab.IgM|Asialoganglioside GM1 Ab.IgM
C0485835|T201|COMP|9329-4|LNC|Basement membrane Ab|Basement membrane Ab
C0485836|T201|COMP|8062-2|LNC|Cardiolipin Ab|Cardiolipin Ab
C0485837|T201|COMP|8063-0|LNC|Cardiolipin Ab.IgA|Cardiolipin Ab.IgA
C0485838|T201|COMP|8065-5|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C0485839|T201|COMP|8067-1|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C0485840|T201|COMP|8068-9|LNC|Centromere Ab|Centromere Ab
C0485841|T201|COMP|10360-6|LNC|DNA single strand Ab.IgG|DNA single strand Ab.IgG
C0485842|T201|COMP|10361-4|LNC|DNA single strand Ab.IgM|DNA single strand Ab.IgM
C0485843|T201|COMP|10362-2|LNC|Endomysium Ab.IgA|Endomysium Ab.IgA
C0485844|T201|COMP|8069-7|LNC|Epidermis Ab|Epidermis Ab
C0485845|T201|COMP|6924-5|LNC|Gliadin Ab.IgA|Gliadin Ab.IgA
C0485846|T201|COMP|8070-5|LNC|Gliadin Ab.IgM|Gliadin Ab.IgM
C0485847|T201|COMP|8071-3|LNC|Histone Ab|Histone Ab
C0485848|T201|COMP|8072-1|LNC|Insulin Ab|Insulin Ab
C0485849|T201|COMP|8073-9|LNC|Insulin bovine Ab|Insulin bovine Ab
C0485850|T201|COMP|8074-7|LNC|Insulin human Ab|Insulin human Ab
C0485851|T201|COMP|8075-4|LNC|Insulin porcine Ab|Insulin porcine Ab
C0485852|T201|COMP|9424-3|LNC|Intercellular substance Ab|Intercellular substance Ab
C0485853|T201|COMP|8076-2|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C0485854|T201|COMP|9838-4|LNC|Liver kidney microsomal Ab|Liver kidney microsomal Ab
C0485855|T201|COMP|8077-0|LNC|Mitochondria Ab|Mitochondria Ab
C0485856|T201|COMP|6925-2|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C0485857|T201|COMP|6926-0|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C0485858|T201|COMP|8078-8|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C0485859|T201|COMP|8079-6|LNC|Myelin Ab.IgA|Myelin Ab.IgA
C0485860|T201|COMP|8080-4|LNC|Myelin Ab.IgG|Myelin Ab.IgG
C0485861|T201|COMP|8081-2|LNC|Myelin Ab.IgM|Myelin Ab.IgM
C0485862|T201|COMP|8082-0|LNC|Myelin basic protein Ab|Myelin basic protein Ab
C0485863|T201|COMP|6969-0|LNC|Myeloperoxidase Ab|Myeloperoxidase Ab
C0485864|T201|COMP|8083-8|LNC|Myocardium Ab|Myocardium Ab
C0485865|T201|COMP|8084-6|LNC|Neutrophil cytoplasmic Ab.classic|Neutrophil cytoplasmic Ab.classic
C0485866|T201|COMP|8085-3|LNC|Neutrophil cytoplasmic Ab.perinuclear|Neutrophil cytoplasmic Ab.perinuclear
C0485867|T201|COMP|9423-5|LNC|Nuclear Ab|Nuclear Ab
C0485868|T201|COMP|8086-1|LNC|Pancreatic islet cell Ab|Pancreatic islet cell Ab
C0485869|T201|COMP|8087-9|LNC|Parietal cell Ab|Parietal cell Ab
C0485870|T201|COMP|8088-7|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C0485871|T201|COMP|6927-8|LNC|Platelet Ab.IgG|Platelet Ab.IgG
C0485872|T201|COMP|8089-5|LNC|Platelet associated Ab.IgG|Platelet associated Ab.IgG
C0485873|T201|COMP|8090-3|LNC|Platelet associated Ab.IgM|Platelet associated Ab.IgM
C0485874|T201|COMP|6968-2|LNC|Proteinase 3 Ab|Proteinase 3 Ab
C0485875|T201|COMP|6970-8|LNC|Purkinje cells Ab|Purkinje cells Ab
C0485876|T201|COMP|9398-9|LNC|Reticulin Ab|Reticulin Ab
C0485877|T201|COMP|9720-4|LNC|Reticulin Ab.IgA|Reticulin Ab.IgA
C0485878|T201|COMP|9839-2|LNC|Rheumatoid arthritis nuclear Ab|Rheumatoid arthritis nuclear Ab
C0485879|T201|COMP|6928-6|LNC|Rheumatoid factor|Rheumatoid factor
C0485880|T201|COMP|6823-9|LNC|Rheumatoid factor|Rheumatoid factor
C0485881|T201|COMP|9338-5|LNC|Rheumatoid factor.IgM|Rheumatoid factor.IgM
C0485882|T201|COMP|8091-1|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0485883|T201|COMP|9399-7|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0485884|T201|COMP|9721-2|LNC|Salivary gland Ab|Salivary gland Ab
C0485885|T201|COMP|8092-9|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C0485886|T201|COMP|9675-0|LNC|Silicone Ab.IgA|Silicone Ab.IgA
C0485887|T201|COMP|9677-6|LNC|Silicone Ab.IgG|Silicone Ab.IgG
C0485888|T201|COMP|9678-4|LNC|Silicone Ab.IgM|Silicone Ab.IgM
C0485889|T201|COMP|8093-7|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C0485890|T201|COMP|8094-5|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C0485891|T201|COMP|9722-0|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0485892|T201|COMP|8095-2|LNC|Smooth muscle Ab|Smooth muscle Ab
C0485893|T201|COMP|8096-0|LNC|Somatotropin Ab|Somatotropin Ab
C0485894|T201|COMP|9723-8|LNC|Spermatozoa Ab.IgA|Spermatozoa Ab.IgA
C0485895|T201|COMP|9724-6|LNC|Spermatozoa Ab.IgG|Spermatozoa Ab.IgG
C0485896|T201|COMP|9725-3|LNC|Spermatozoa Ab.IgM|Spermatozoa Ab.IgM
C0485897|T201|COMP|9679-2|LNC|Squamous cell carcinoma Ag|Squamous cell carcinoma Ag
C0485898|T201|COMP|8097-8|LNC|Striated muscle Ab|Striated muscle Ab
C0485899|T201|COMP|8098-6|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C0485901|T201|COMP|9580-2|LNC|Thyroxine Ab|Thyroxine Ab
C0485902|T201|COMP|10740-9|LNC|Aluminum.microscopic observation|Aluminum.microscopic observation
C0485903|T201|COMP|10741-7|LNC|Amyloid.microscopic observation|Amyloid.microscopic observation
C0485904|T201|COMP|10742-5|LNC|Amyloid.microscopic observation|Amyloid.microscopic observation
C0485905|T201|COMP|10743-3|LNC|Amyloid.microscopic observation|Amyloid.microscopic observation
C0485906|T201|COMP|10744-1|LNC|Amyloid.microscopic observation|Amyloid.microscopic observation
C0485907|T201|COMP|10745-8|LNC|Bile.microscopic observation|Bile.microscopic observation
C0485908|T201|COMP|10746-6|LNC|Calcium.microscopic observation|Calcium.microscopic observation
C0485911|T201|COMP|10749-0|LNC|Collagen fibers.microscopic observation|Collagen fibers.microscopic observation
C0485912|T201|COMP|10750-8|LNC|Connective tissue.microscopic observation|Connective tissue.microscopic observation
C0485913|T201|COMP|10751-6|LNC|Copper.microscopic observation|Copper.microscopic observation
C0485914|T201|COMP|10752-4|LNC|Fat.microscopic observation|Fat.microscopic observation
C0485915|T201|COMP|10753-2|LNC|Fat.microscopic observation|Fat.microscopic observation
C0485916|T201|COMP|10754-0|LNC|Fat.microscopic observation|Fat.microscopic observation
C0485917|T201|COMP|10755-7|LNC|Fungus.microscopic observation|Fungus.microscopic observation
C0485918|T201|COMP|10756-5|LNC|Glial fibers.microscopic observation|Glial fibers.microscopic observation
C0485920|T201|COMP|10758-1|LNC|Iron.microscopic observation|Iron.microscopic observation
C0485921|T201|COMP|10759-9|LNC|Iron.microscopic observation|Iron.microscopic observation
C0485922|T201|COMP|10760-7|LNC|Iron.microscopic observation|Iron.microscopic observation
C0485923|T201|COMP|10761-5|LNC|Iron.microscopic observation|Iron.microscopic observation
C0485983|T201|COMP|10822-5|LNC|Mucin.microscopic observation|Mucin.microscopic observation
C0485984|T201|COMP|10823-3|LNC|Mucopolysaccharides.microscopic observation|Mucopolysaccharides.microscopic observation
C0485986|T201|COMP|10825-8|LNC|Myelin+Nerve cells.microscopic observation|Myelin+Nerve cells.microscopic observation
C0485987|T201|COMP|10826-6|LNC|Nissel.microscopic observation|Nissel.microscopic observation
C0485988|T201|COMP|10827-4|LNC|Reticulum.microscopic observation|Reticulum.microscopic observation
C0485989|T201|COMP|8100-0|LNC|Specimen preparation|Specimen preparation
C0485990|T201|COMP|10828-2|LNC|Urate crystals.microscopic observation|Urate crystals.microscopic observation
C0485991|T201|COMP|9681-8|LNC|1-Naphthol|1-Naphthol
C0485992|T201|COMP|6971-6|LNC|2,4 toluenediamine|2,4 toluenediamine
C0485993|T201|COMP|9806-1|LNC|2,4-Dichlorophenoxyacetate|2,4-Dichlorophenoxyacetate
C0485994|T201|COMP|6972-4|LNC|2,6 toluenediamine|2,6 toluenediamine
C0485995|T201|COMP|9682-6|LNC|2-Butanol|2-Butanol
C0485996|T201|COMP|9683-4|LNC|2-Methyl-2-Propanol|2-Methyl-2-Propanol
C0485997|T201|COMP|9432-6|LNC|Isobutyl acetate|Isobutyl acetate
C0485998|T201|COMP|9425-0|LNC|Acetone|Acetone
C0485999|T201|COMP|9430-0|LNC|Isobutylcarbinol|Isobutylcarbinol
C0486000|T201|COMP|6929-4|LNC|Aluminum|Aluminum
C0486001|T201|COMP|9462-3|LNC|Aluminum|Aluminum
C0486002|T201|COMP|8140-6|LNC|Amphetamines|Amphetamines
C0486003|T201|COMP|8141-4|LNC|Amphetamines|Amphetamines
C0486004|T201|COMP|8142-2|LNC|Amphetamines|Amphetamines
C0486005|T201|COMP|8139-8|LNC|Amphetamines|Amphetamines
C0486006|T201|COMP|8144-8|LNC|Amphetamines|Amphetamines
C0486007|T201|COMP|8145-5|LNC|Amphetamines|Amphetamines
C0486008|T201|COMP|8146-3|LNC|Amphetamines|Amphetamines
C0486009|T201|COMP|8143-0|LNC|Amphetamines|Amphetamines
C0486010|T201|COMP|8148-9|LNC|Amphetamines|Amphetamines
C0486011|T201|COMP|8149-7|LNC|Amphetamines|Amphetamines
C0486012|T201|COMP|8147-1|LNC|Amphetamines|Amphetamines
C0486013|T201|COMP|8151-3|LNC|Amphetamines|Amphetamines
C0486014|T201|COMP|8152-1|LNC|Amphetamines|Amphetamines
C0486015|T201|COMP|8150-5|LNC|Amphetamines|Amphetamines
C0486016|T201|COMP|8154-7|LNC|Amphetamines|Amphetamines
C0486017|T201|COMP|8155-4|LNC|Amphetamines|Amphetamines
C0486018|T201|COMP|8156-2|LNC|Amphetamines|Amphetamines
C0486019|T201|COMP|8153-9|LNC|Amphetamines|Amphetamines
C0486020|T201|COMP|9489-6|LNC|Arsenic|Arsenic
C0486021|T201|COMP|8157-0|LNC|Arsenic|Arsenic
C0486022|T201|COMP|8158-8|LNC|Arsenic|Arsenic
C0486023|T201|COMP|9463-1|LNC|Arsenic|Arsenic
C0486024|T201|COMP|9366-6|LNC|Arsenic|Arsenic
C0486025|T201|COMP|9427-6|LNC|Barbiturates|Barbiturates
C0486026|T201|COMP|9426-8|LNC|Barbiturates|Barbiturates
C0486027|T201|COMP|10363-0|LNC|Barbiturates|Barbiturates
C0486028|T201|COMP|9464-9|LNC|Barium|Barium
C0486029|T201|COMP|9684-2|LNC|Bendiocarb|Bendiocarb
C0486030|T201|COMP|9330-2|LNC|Benzene|Benzene
C0486031|T201|COMP|9465-6|LNC|Benzene|Benzene
C0486032|T201|COMP|9428-4|LNC|Benzodiazepines|Benzodiazepines
C0486033|T201|COMP|8159-6|LNC|Beryllium|Beryllium
C0486034|T201|COMP|8160-4|LNC|Beryllium|Beryllium
C0486035|T201|COMP|8161-2|LNC|Bismuth|Bismuth
C0486036|T201|COMP|9493-8|LNC|Bismuth|Bismuth
C0486037|T201|COMP|9367-4|LNC|Borate|Borate
C0486038|T201|COMP|9331-0|LNC|Boron|Boron
C0486039|T201|COMP|9368-2|LNC|Boron|Boron
C0486040|T201|COMP|9497-9|LNC|Butane|Butane
C0486041|T201|COMP|9685-9|LNC|Butanol|Butanol
C0486042|T201|COMP|9686-7|LNC|Cadmium|Cadmium
C0486043|T201|COMP|9466-4|LNC|Cadmium|Cadmium
C0486044|T201|COMP|9687-5|LNC|Cadmium|Cadmium
C0486045|T201|COMP|9467-2|LNC|Calcium|Calcium
C0486046|T201|COMP|9369-0|LNC|Camphor|Camphor
C0486047|T201|COMP|8163-8|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486048|T201|COMP|8164-6|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486049|T201|COMP|8165-3|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486050|T201|COMP|8162-0|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486051|T201|COMP|8167-9|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486052|T201|COMP|8168-7|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486053|T201|COMP|8169-5|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486054|T201|COMP|8166-1|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486055|T201|COMP|8171-1|LNC|Cannabinoids|Cannabinoids
C0486056|T201|COMP|8172-9|LNC|Cannabinoids|Cannabinoids
C0486057|T201|COMP|8170-3|LNC|Cannabinoids|Cannabinoids
C0486058|T201|COMP|8174-5|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486059|T201|COMP|8175-2|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486060|T201|COMP|8173-7|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486061|T201|COMP|8177-8|LNC|Cannabinoids|Cannabinoids
C0486062|T201|COMP|8178-6|LNC|Cannabinoids|Cannabinoids
C0486063|T201|COMP|8179-4|LNC|Cannabinoids|Cannabinoids
C0486064|T201|COMP|8176-0|LNC|Cannabinoids|Cannabinoids
C0486065|T201|COMP|9789-9|LNC|Carbamate pesticides|Carbamate pesticides
C0486066|T201|COMP|9688-3|LNC|Carbaryl|Carbaryl
C0486067|T201|COMP|9689-1|LNC|Carbofuran|Carbofuran
C0486068|T201|COMP|9332-8|LNC|Carbon tetrachloride|Carbon tetrachloride
C0486069|T201|COMP|9502-6|LNC|Carbophenothion|Carbophenothion
C0486070|T201|COMP|9468-0|LNC|Chloramines|Chloramines
C0486071|T201|COMP|9807-9|LNC|Chlordane|Chlordane
C0486072|T201|COMP|8180-2|LNC|Chlorobenzene|Chlorobenzene
C0486073|T201|COMP|9505-9|LNC|Chlorobenzene|Chlorobenzene
C0486074|T201|COMP|9506-7|LNC|Chloroethane|Chloroethane
C0486075|T201|COMP|9333-6|LNC|Chloroform|Chloroform
C0486076|T201|COMP|9507-5|LNC|Chloromethane|Chloromethane
C0486077|T201|COMP|9371-6|LNC|Chlorpyrifos|Chlorpyrifos
C0486078|T201|COMP|9510-9|LNC|Chromium|Chromium
C0486079|T201|COMP|8181-0|LNC|Chromium|Chromium
C0486080|T201|COMP|9469-8|LNC|Chromium|Chromium
C0486081|T201|COMP|9690-9|LNC|Chromium|Chromium
C0486082|T201|COMP|9691-7|LNC|Cobalt|Cobalt
C0486083|T201|COMP|8183-6|LNC|Benzoylecgonine|Benzoylecgonine
C0486084|T201|COMP|8184-4|LNC|Benzoylecgonine|Benzoylecgonine
C0486085|T201|COMP|8185-1|LNC|Benzoylecgonine|Benzoylecgonine
C0486086|T201|COMP|8182-8|LNC|Benzoylecgonine|Benzoylecgonine
C0486087|T201|COMP|8187-7|LNC|Benzoylecgonine|Benzoylecgonine
C0486088|T201|COMP|8188-5|LNC|Benzoylecgonine|Benzoylecgonine
C0486089|T201|COMP|8189-3|LNC|Benzoylecgonine|Benzoylecgonine
C0486090|T201|COMP|8186-9|LNC|Benzoylecgonine|Benzoylecgonine
C0486091|T201|COMP|8190-1|LNC|Cocaine|Cocaine
C0486092|T201|COMP|8191-9|LNC|Cocaine|Cocaine
C0486093|T201|COMP|8192-7|LNC|Benzoylecgonine|Benzoylecgonine
C0486094|T201|COMP|8193-5|LNC|Benzoylecgonine|Benzoylecgonine
C0486095|T201|COMP|8195-0|LNC|Cocaine|Cocaine
C0486096|T201|COMP|8196-8|LNC|Cocaine|Cocaine
C0486097|T201|COMP|8197-6|LNC|Cocaine|Cocaine
C0486098|T201|COMP|8194-3|LNC|Cocaine|Cocaine
C0486099|T201|COMP|8198-4|LNC|Copper|Copper
C0486100|T201|COMP|9470-6|LNC|Copper|Copper
C0486101|T201|COMP|10364-8|LNC|Cotinine|Cotinine
C0486102|T201|COMP|10365-5|LNC|Cotinine|Cotinine
C0486103|T201|COMP|10366-3|LNC|Cotinine|Cotinine
C0486104|T201|COMP|9372-4|LNC|Cotinine|Cotinine
C0486105|T201|COMP|9512-5|LNC|Creosol|Creosol
C0486106|T201|COMP|10367-1|LNC|Ethanol|Ethanol
C0486107|T201|COMP|8199-2|LNC|Ethyl benzene|Ethyl benzene
C0486108|T201|COMP|9471-4|LNC|Fluoride|Fluoride
C0486109|T201|COMP|8200-8|LNC|Gadolinium|Gadolinium
C0486110|T201|COMP|8201-6|LNC|Gadolinium|Gadolinium
C0486111|T201|COMP|9472-2|LNC|Heptachlor|Heptachlor
C0486112|T201|COMP|9473-0|LNC|Heptachlorepoxide|Heptachlorepoxide
C0486113|T201|COMP|9474-8|LNC|Hexachlorobenzene|Hexachlorobenzene
C0486115|T201|COMP|9476-3|LNC|Hexanoylglycine|Hexanoylglycine
C0486116|T201|COMP|9429-2|LNC|Indium|Indium
C0486117|T201|COMP|9431-8|LNC|Isobutanol|Isobutanol
C0486118|T201|COMP|9692-5|LNC|Isobutanol|Isobutanol
C0486119|T201|COMP|9433-4|LNC|Isoflurane|Isoflurane
C0486120|T201|COMP|9435-9|LNC|Isopropanol|Isopropanol
C0486121|T201|COMP|9434-2|LNC|Isopropanol|Isopropanol
C0486122|T201|COMP|10368-9|LNC|Lead|Lead
C0486123|T201|COMP|9436-7|LNC|Lead|Lead
C0486124|T201|COMP|8202-4|LNC|Lead|Lead
C0486125|T201|COMP|9477-1|LNC|Lead|Lead
C0486126|T201|COMP|9478-9|LNC|Magnesium|Magnesium
C0486127|T201|COMP|8203-2|LNC|Manganese|Manganese
C0486128|T201|COMP|9693-3|LNC|Mercury|Mercury
C0486129|T201|COMP|8204-0|LNC|Mercury|Mercury
C0486130|T201|COMP|8205-7|LNC|Mercury|Mercury
C0486131|T201|COMP|6693-6|LNC|Mercury|Mercury
C0486132|T201|COMP|9479-7|LNC|Mercury|Mercury
C0486133|T201|COMP|9726-1|LNC|Mescaline|Mescaline
C0486134|T201|COMP|9334-4|LNC|Methanol|Methanol
C0486135|T201|COMP|9790-7|LNC|Methyl bromide|Methyl bromide
C0486136|T201|COMP|9437-5|LNC|Methylhippurate|Methylhippurate
C0486138|T201|COMP|8207-3|LNC|Nickel|Nickel
C0486139|T201|COMP|8208-1|LNC|Nickel|Nickel
C0486140|T201|COMP|9480-5|LNC|Nitrate|Nitrate
C0486141|T201|COMP|8210-7|LNC|Opiates|Opiates
C0486142|T201|COMP|8211-5|LNC|Opiates|Opiates
C0486143|T201|COMP|8212-3|LNC|Opiates|Opiates
C0486144|T201|COMP|8209-9|LNC|Opiates|Opiates
C0486145|T201|COMP|10369-7|LNC|Opiates|Opiates
C0486146|T201|COMP|8214-9|LNC|Opiates|Opiates
C0486147|T201|COMP|8215-6|LNC|Opiates|Opiates
C0486148|T201|COMP|8216-4|LNC|Opiates|Opiates
C0486149|T201|COMP|8213-1|LNC|Opiates|Opiates
C0486150|T201|COMP|8218-0|LNC|Opiates|Opiates
C0486151|T201|COMP|8219-8|LNC|Opiates|Opiates
C0486152|T201|COMP|8217-2|LNC|Opiates|Opiates
C0486153|T201|COMP|8221-4|LNC|Opiates|Opiates
C0486154|T201|COMP|8222-2|LNC|Opiates|Opiates
C0486155|T201|COMP|8220-6|LNC|Opiates|Opiates
C0486156|T201|COMP|8224-8|LNC|Opiates|Opiates
C0486157|T201|COMP|8225-5|LNC|Opiates|Opiates
C0486158|T201|COMP|8226-3|LNC|Opiates|Opiates
C0486159|T201|COMP|8223-0|LNC|Opiates|Opiates
C0486160|T201|COMP|9791-5|LNC|Organochlorine pesticides|Organochlorine pesticides
C0486161|T201|COMP|9792-3|LNC|Organophosphate pesticides|Organophosphate pesticides
C0486162|T201|COMP|9827-7|LNC|Paraquat|Paraquat
C0486163|T201|COMP|8228-9|LNC|Phencyclidine|Phencyclidine
C0486164|T201|COMP|8229-7|LNC|Phencyclidine|Phencyclidine
C0486165|T201|COMP|8230-5|LNC|Phencyclidine|Phencyclidine
C0486166|T201|COMP|8227-1|LNC|Phencyclidine|Phencyclidine
C0486167|T201|COMP|10370-5|LNC|Phencyclidine|Phencyclidine
C0486168|T201|COMP|8232-1|LNC|Phencyclidine|Phencyclidine
C0486169|T201|COMP|8233-9|LNC|Phencyclidine|Phencyclidine
C0486170|T201|COMP|8234-7|LNC|Phencyclidine|Phencyclidine
C0486171|T201|COMP|8231-3|LNC|Phencyclidine|Phencyclidine
C0486172|T201|COMP|8235-4|LNC|Phencyclidine|Phencyclidine
C0486173|T201|COMP|8236-2|LNC|Phencyclidine|Phencyclidine
C0486174|T201|COMP|8237-0|LNC|Phencyclidine|Phencyclidine
C0486175|T201|COMP|8238-8|LNC|Phencyclidine|Phencyclidine
C0486176|T201|COMP|8240-4|LNC|Phencyclidine|Phencyclidine
C0486177|T201|COMP|8241-2|LNC|Phencyclidine|Phencyclidine
C0486178|T201|COMP|8242-0|LNC|Phencyclidine|Phencyclidine
C0486179|T201|COMP|8239-6|LNC|Phencyclidine|Phencyclidine
C0486180|T201|COMP|9808-7|LNC|Phenothiazines|Phenothiazines
C0486181|T201|COMP|9400-3|LNC|Platinum|Platinum
C0486182|T201|COMP|9694-1|LNC|Propoxur|Propoxur
C0486183|T201|COMP|9809-5|LNC|Propoxyphene|Propoxyphene
C0486185|T201|COMP|9810-3|LNC|quiNINE|quiNINE
C0486186|T201|COMP|9483-9|LNC|Selenium|Selenium
C0486187|T201|COMP|10829-0|LNC|Silicon|Silicon
C0486188|T201|COMP|9401-1|LNC|Silicon|Silicon
C0486189|T201|COMP|6931-0|LNC|Silver|Silver
C0486190|T201|COMP|9484-7|LNC|Silver|Silver
C0486191|T201|COMP|8243-8|LNC|Styrene|Styrene
C0486192|T201|COMP|8244-6|LNC|Titanium|Titanium
C0486193|T201|COMP|9637-0|LNC|Toluene|Toluene
C0486194|T201|COMP|9638-8|LNC|Toluene|Toluene
C0486195|T201|COMP|9793-1|LNC|Trichloroethylene|Trichloroethylene
C0486196|T201|COMP|8245-3|LNC|Zinc|Zinc
C0486197|T201|COMP|6973-2|LNC|Zinc|Zinc
C0486198|T201|COMP|9487-0|LNC|Zinc|Zinc
C0486199|T201|COMP|6974-0|LNC|Zirconium|Zirconium
C0486200|T201|COMP|8246-1|LNC|Amorphous sediment|Amorphous sediment
C0486201|T201|COMP|9335-1|LNC|Appearance|Appearance
C0486203|T201|COMP|9439-1|LNC|Casts|Casts
C0486204|T201|COMP|9842-6|LNC|Casts|Casts
C0486205|T201|COMP|9374-0|LNC|Character|Character
C0486206|T201|COMP|6824-7|LNC|Color|Color
C0486207|T201|COMP|9397-1|LNC|Color|Color
C0486208|T201|COMP|6825-4|LNC|Crystals|Crystals
C0486209|T201|COMP|6826-2|LNC|Crystals|Crystals
C0486210|T201|COMP|8247-9|LNC|Mucus|Mucus
C0486211|T201|COMP|8248-7|LNC|Spermatozoa|Spermatozoa
C0486212|T201|COMP|8249-5|LNC|Transitional cells|Transitional cells
C0486213|T201|COMP|1016-5|LNC|E Ab|E Ab
C0486214|T201|COMP|1017-3|LNC|E Ab|E Ab
C0486215|T201|COMP|1018-1|LNC|E Ab|E Ab
C0486216|T201|COMP|1019-9|LNC|E Ag|E Ag
C0486217|T201|COMP|1020-7|LNC|E Ag|E Ag
C0486218|T201|COMP|1021-5|LNC|E Ag|E Ag
C0486219|T201|COMP|1058-7|LNC|I Ab|I Ab
C0486220|T201|COMP|1059-5|LNC|I Ab|I Ab
C0486221|T201|COMP|1060-3|LNC|I Ab|I Ab
C0486222|T201|COMP|1064-5|LNC|I NOS Ag|I NOS Ag
C0486223|T201|COMP|1065-2|LNC|I NOS Ag|I NOS Ag
C0486224|T201|COMP|10400-0|LNC|I Ag|I Ag
C0486225|T201|COMP|1091-8|LNC|K Ab|K Ab
C0486226|T201|COMP|1092-6|LNC|K Ab|K Ab
C0486227|T201|COMP|1093-4|LNC|K Ab|K Ab
C0486228|T201|COMP|1094-2|LNC|K Ag|K Ag
C0486229|T201|COMP|1095-9|LNC|K Ag|K Ag
C0486230|T201|COMP|1096-7|LNC|K Ag|K Ag
C0486231|T201|COMP|1160-1|LNC|little e Ab|little e Ab
C0486232|T201|COMP|1161-9|LNC|little e Ab|little e Ab
C0486233|T201|COMP|1162-7|LNC|little e Ab|little e Ab
C0486234|T201|COMP|1163-5|LNC|little e Ag|little e Ag
C0486235|T201|COMP|1164-3|LNC|little e Ag|little e Ag
C0486236|T201|COMP|1165-0|LNC|little e Ag|little e Ag
C0486237|T201|COMP|1184-1|LNC|little i Ab|little i Ab
C0486238|T201|COMP|1185-8|LNC|little i Ab|little i Ab
C0486239|T201|COMP|1186-6|LNC|little i Ab|little i Ab
C0486240|T201|COMP|10406-7|LNC|little i Ag|little i Ag
C0486241|T201|COMP|1188-2|LNC|little i NOS Ag|little i NOS Ag
C0486242|T201|COMP|1189-0|LNC|little i NOS Ag|little i NOS Ag
C0486243|T201|COMP|1190-8|LNC|little k Ab|little k Ab
C0486244|T201|COMP|1191-6|LNC|little k Ab|little k Ab
C0486245|T201|COMP|1192-4|LNC|little k Ab|little k Ab
C0486246|T201|COMP|1193-2|LNC|little k Ag|little k Ag
C0486247|T201|COMP|1194-0|LNC|little k Ag|little k Ag
C0486248|T201|COMP|1195-7|LNC|little k Ag|little k Ag
C0486249|T201|COMP|1208-8|LNC|little s Ab|little s Ab
C0486250|T201|COMP|1209-6|LNC|little s Ab|little s Ab
C0486251|T201|COMP|1210-4|LNC|little s Ab|little s Ab
C0486252|T201|COMP|1211-2|LNC|little s Ag|little s Ag
C0486253|T201|COMP|1212-0|LNC|little s Ag|little s Ag
C0486254|T201|COMP|1213-8|LNC|little s Ag|little s Ag
C0486255|T201|COMP|1315-1|LNC|S Ab|S Ab
C0486256|T201|COMP|1316-9|LNC|S Ab|S Ab
C0486257|T201|COMP|8114-1|LNC|Cells.CD16-CD57+/100 cells|Cells.CD16-CD57+/100 cells
C0486258|T201|COMP|9336-9|LNC|IgA subclass 1/IgA.total|IgA subclass 1/IgA.total
C0486259|T201|COMP|5895-7|LNC|Coagulation tissue factor induced.INR|Coagulation tissue factor induced.INR
C0486260|T201|COMP|5896-5|LNC|Coagulation tissue factor induced.normal/Actual|Coagulation tissue factor induced.normal/Actual
C0486262|T201|COMP|4467-7|LNC|Spinnbarkeit test|Spinnbarkeit test
C0488650|T201|COMP|10226-9|LNC|Oxygen content|Oxygen content
C0488752|T201|COMP|10232-7|LNC|Oxygen content|Oxygen content
C0488753|T201|COMP|10233-5|LNC|Oxygen content|Oxygen content
C0488754|T201|COMP|10234-3|LNC|Oxygen content|Oxygen content
C0488755|T201|COMP|10235-0|LNC|Oxygen content|Oxygen content
C0488756|T201|COMP|10236-8|LNC|Oxygen content|Oxygen content
C0488757|T201|COMP|10237-6|LNC|Oxygen content|Oxygen content
C0488758|T201|COMP|10238-4|LNC|Oxygen content|Oxygen content
C0488759|T201|COMP|10239-2|LNC|Oxygen content|Oxygen content
C0488760|T201|COMP|10240-0|LNC|Oxygen content|Oxygen content
C0488761|T201|COMP|10241-8|LNC|Oxygen content|Oxygen content
C0488762|T201|COMP|10242-6|LNC|Oxygen content|Oxygen content
C0488763|T201|COMP|10243-4|LNC|Oxygen content|Oxygen content
C0488764|T201|COMP|10244-2|LNC|Oxygen content|Oxygen content
C0488765|T201|COMP|10245-9|LNC|Oxygen content|Oxygen content
C0488766|T201|COMP|10246-7|LNC|Oxygen content|Oxygen content
C0488767|T201|COMP|10247-5|LNC|Oxygen content|Oxygen content
C0488768|T201|COMP|10248-3|LNC|Oxygen content|Oxygen content
C0549668|T201|COMP|13450-2|LNC|Creatinine renal clearance/1.73 sq M|Creatinine renal clearance/1.73 sq M
C0549671|T201|COMP|13094-8|LNC|Monosialoganglioside GM1 Ab.IgA|Monosialoganglioside GM1 Ab.IgA
C0549673|T201|COMP|10868-8|LNC|Bacitracin|Bacitracin
C0549674|T201|COMP|11575-8|LNC|Cefmetazole|Cefmetazole
C0549675|T201|COMP|11576-6|LNC|Erythromycin+sulfiSOXAZOLE|Erythromycin+sulfiSOXAZOLE
C0549676|T201|COMP|11577-4|LNC|Sulfamethoxazole|Sulfamethoxazole
C0549677|T201|COMP|11578-2|LNC|sulfiSOXAZOLE|sulfiSOXAZOLE
C0549678|T201|COMP|11159-1|LNC|Alkalase Ab.IgE|Alkalase Ab.IgE
C0549679|T201|COMP|10919-9|LNC|Anisakis Ab.IgE|Anisakis Ab.IgE
C0549680|T201|COMP|10930-6|LNC|Artemia salina Ab.IgE|Artemia salina Ab.IgE
C0549681|T201|COMP|11030-4|LNC|(Aspergillus fumigatus+Aspergillus niger) Ab.IgE|(Aspergillus fumigatus+Aspergillus niger) Ab.IgE
C0549682|T201|COMP|10920-7|LNC|Phyllostachys pubescens Ab.IgE|Phyllostachys pubescens Ab.IgE
C0549683|T201|COMP|11160-9|LNC|Beta lactoglobulin Ab.IgG|Beta lactoglobulin Ab.IgG
C0549684|T201|COMP|10921-5|LNC|Blomia tropicalis Ab.IgE|Blomia tropicalis Ab.IgE
C0549685|T201|COMP|11161-7|LNC|Bran wheat Ab.IgE|Bran wheat Ab.IgE
C0549686|T201|COMP|10923-1|LNC|Bromelin Ab.IgE|Bromelin Ab.IgE
C0549688|T201|COMP|13216-7|LNC|Candida albicans immune complex|Candida albicans immune complex
C0549689|T201|COMP|11163-3|LNC|Carageenan Ab.IgE|Carageenan Ab.IgE
C0549690|T201|COMP|10924-9|LNC|Averrhoa carambola Ab.IgE|Averrhoa carambola Ab.IgE
C0549691|T201|COMP|11164-1|LNC|Cheese cream Ab.IgE|Cheese cream Ab.IgE
C0549692|T201|COMP|11165-8|LNC|Chinchilla Ab.IgE|Chinchilla Ab.IgE
C0549693|T201|COMP|11166-6|LNC|Chortoglyphus arcuatus Ab.IgE|Chortoglyphus arcuatus Ab.IgE
C0549694|T201|COMP|11167-4|LNC|Cockatiel feather Ab.IgE|Cockatiel feather Ab.IgE
C0549695|T201|COMP|13184-7|LNC|Populus deltoides Ab.IgG|Populus deltoides Ab.IgG
C0549696|T201|COMP|11168-2|LNC|Cupressus arizonica Ab.IgE|Cupressus arizonica Ab.IgE
C0549697|T201|COMP|10931-4|LNC|Daphnia Ab.IgE|Daphnia Ab.IgE
C0549698|T201|COMP|10926-4|LNC|Deer epithelium Ab.IgE|Deer epithelium Ab.IgE
C0549699|T201|COMP|11169-0|LNC|Deer hair Ab.IgE|Deer hair Ab.IgE
C0549700|T201|COMP|11170-8|LNC|Dematiaceae Ab.IgE|Dematiaceae Ab.IgE
C0549701|T201|COMP|13186-2|LNC|Rumex crispus Ab.IgG|Rumex crispus Ab.IgG
C0549702|T201|COMP|10927-2|LNC|Elk meat Ab.IgE|Elk meat Ab.IgE
C0549703|T201|COMP|13183-9|LNC|Ulmus americana Ab.IgG|Ulmus americana Ab.IgG
C0549704|T201|COMP|11171-6|LNC|Erythromycin Ab.IgE|Erythromycin Ab.IgE
C0549705|T201|COMP|10928-0|LNC|Foeniculum vulgare fresh Ab.IgE|Foeniculum vulgare fresh Ab.IgE
C0549706|T201|COMP|10929-8|LNC|Foeniculum vulgare seed Ab.IgE|Foeniculum vulgare seed Ab.IgE
C0549707|T201|COMP|11172-4|LNC|Ferret epithelium Ab.IgE|Ferret epithelium Ab.IgE
C0549708|T201|COMP|11173-2|LNC|Ficus carica Ab.IgE|Ficus carica Ab.IgE
C0549709|T201|COMP|13180-5|LNC|Formaldehyde Ab.IgG|Formaldehyde Ab.IgG
C0549710|T201|COMP|13190-4|LNC|Formaldehyde Ab.IgM|Formaldehyde Ab.IgM
C0549711|T201|COMP|13181-3|LNC|Paspalum notatum Ab.IgG|Paspalum notatum Ab.IgG
C0549712|T201|COMP|10933-0|LNC|Cyamopsis tetragonoloba Ab.IgE|Cyamopsis tetragonoloba Ab.IgE
C0549713|T201|COMP|10934-8|LNC|Psidium guajava Ab.IgE|Psidium guajava Ab.IgE
C0549714|T201|COMP|11175-7|LNC|Helminthosporium sativum Ab.IgE|Helminthosporium sativum Ab.IgE
C0549715|T201|COMP|10935-5|LNC|Horse serum proteins Ab.IgE|Horse serum proteins Ab.IgE
C0549716|T201|COMP|11176-5|LNC|Lactalbumin alpha Ab.IgG|Lactalbumin alpha Ab.IgG
C0549717|T201|COMP|11177-3|LNC|Lactalbumin beta Ab.IgE|Lactalbumin beta Ab.IgE
C0549718|T201|COMP|11178-1|LNC|Beta galactosidase Ab.IgE|Beta galactosidase Ab.IgE
C0549719|T201|COMP|11179-9|LNC|Tilia cordata Ab.IgE|Tilia cordata Ab.IgE
C0549720|T201|COMP|11180-7|LNC|Lupinus spp Ab.IgE|Lupinus spp Ab.IgE
C0549721|T201|COMP|11181-5|LNC|Lycopodium spp Ab.IgE|Lycopodium spp Ab.IgE
C0549722|T201|COMP|11182-3|LNC|Lysozyme Ab.IgE|Lysozyme Ab.IgE
C0549723|T201|COMP|11183-1|LNC|Macadamia spp Ab.IgE|Macadamia spp Ab.IgE
C0549724|T201|COMP|10925-6|LNC|Scomber japonicus Ab.IgE|Scomber japonicus Ab.IgE
C0549725|T201|COMP|11184-9|LNC|Trachurus japonicus Ab.IgE|Trachurus japonicus Ab.IgE
C0549726|T201|COMP|10936-3|LNC|Mare milk Ab.IgE|Mare milk Ab.IgE
C0549727|T201|COMP|10937-1|LNC|Origanum majorana Ab.IgE|Origanum majorana Ab.IgE
C0549728|T201|COMP|11185-6|LNC|Maxatase Ab.IgE|Maxatase Ab.IgE
C0549729|T201|COMP|10939-7|LNC|Lepidorhombus whiffiagonis Ab.IgE|Lepidorhombus whiffiagonis Ab.IgE
C0549730|T201|COMP|13182-1|LNC|Prosopis juliflora Ab.IgG|Prosopis juliflora Ab.IgG
C0549731|T201|COMP|10940-5|LNC|Cow milk boiled Ab.IgE|Cow milk boiled Ab.IgE
C0549732|T201|COMP|10941-3|LNC|Milk powder Ab.IgE|Milk powder Ab.IgE
C0549733|T201|COMP|11186-4|LNC|Setaria italica Ab.IgE|Setaria italica Ab.IgE
C0549734|T201|COMP|10942-1|LNC|Echinochloa crus-galli Ab.IgE|Echinochloa crus-galli Ab.IgE
C0549735|T201|COMP|10943-9|LNC|Mink epithelium Ab.IgE|Mink epithelium Ab.IgE
C0549736|T201|COMP|10938-9|LNC|Ephestia kuehniella Ab.IgE|Ephestia kuehniella Ab.IgE
C0549737|T201|COMP|13188-8|LNC|Artemisia vulgaris Ab.IgG|Artemisia vulgaris Ab.IgG
C0549738|T201|COMP|13185-4|LNC|Urtica dioica Ab.IgG|Urtica dioica Ab.IgG
C0549739|T201|COMP|10944-7|LNC|Octopus vulgaris Ab.IgE|Octopus vulgaris Ab.IgE
C0549740|T201|COMP|13177-1|LNC|Elaeagnus angustifolia Ab.IgE|Elaeagnus angustifolia Ab.IgE
C0549741|T201|COMP|10945-4|LNC|Papain Ab.IgE|Papain Ab.IgE
C0549742|T201|COMP|10946-2|LNC|Passiflora edulis Ab.IgE|Passiflora edulis Ab.IgE
C0549743|T201|COMP|11187-2|LNC|Penicillium frequentans Ab.IgE|Penicillium frequentans Ab.IgE
C0549744|T201|COMP|11188-0|LNC|Pepper cayenne Ab.IgE|Pepper cayenne Ab.IgE
C0549745|T201|COMP|11189-8|LNC|Pepper jalapeno Ab.IgE|Pepper jalapeno Ab.IgE
C0549746|T201|COMP|11190-6|LNC|Mentha piperita Ab.IgE|Mentha piperita Ab.IgE
C0549747|T201|COMP|10947-0|LNC|Diospyros kaki Ab.IgE|Diospyros kaki Ab.IgE
C0549748|T201|COMP|13240-7|LNC|Phoma herbarum Ab.IgE|Phoma herbarum Ab.IgE
C0549749|T201|COMP|10948-8|LNC|Pigeon feather Ab.IgE|Pigeon feather Ab.IgE
C0549750|T201|COMP|10955-3|LNC|Pinus palustris Ab.IgE|Pinus palustris Ab.IgE
C0549751|T201|COMP|10954-6|LNC|Pinus edulis Ab.IgE|Pinus edulis Ab.IgE
C0549752|T201|COMP|10956-1|LNC|Pinus echinata Ab.IgE|Pinus echinata Ab.IgE
C0549753|T201|COMP|10957-9|LNC|Pinus elliottii Ab.IgE|Pinus elliottii Ab.IgE
C0549754|T201|COMP|10958-7|LNC|Pinus virginiana Ab.IgE|Pinus virginiana Ab.IgE
C0549755|T201|COMP|10949-6|LNC|Malassezia furfur Ab.IgE|Malassezia furfur Ab.IgE
C0549756|T201|COMP|13189-6|LNC|Plantago lanceolata Ab.IgG|Plantago lanceolata Ab.IgG
C0549757|T201|COMP|10959-5|LNC|Pleuronectes platessa Ab.IgE|Pleuronectes platessa Ab.IgE
C0549758|T201|COMP|11191-4|LNC|Pollachius virens Ab.IgE|Pollachius virens Ab.IgE
C0549759|T201|COMP|11192-2|LNC|Protamine Ab.IgE|Protamine Ab.IgE
C0549760|T201|COMP|11193-0|LNC|Cucurbita pepo seed Ab.IgE|Cucurbita pepo seed Ab.IgE
C0549761|T201|COMP|10960-3|LNC|Rabbit serum proteins Ab.IgE|Rabbit serum proteins Ab.IgE
C0549762|T201|COMP|10961-1|LNC|Rabbit urine proteins Ab.IgE|Rabbit urine proteins Ab.IgE
C0549763|T201|COMP|13187-0|LNC|Franseria acanthicarpa Ab.IgG|Franseria acanthicarpa Ab.IgG
C0549764|T201|COMP|11194-8|LNC|Brassica napus pollen Ab.IgE|Brassica napus pollen Ab.IgE
C0549765|T201|COMP|11195-5|LNC|Brassica rapa Ab.IgE|Brassica rapa Ab.IgE
C0549766|T201|COMP|10950-4|LNC|Reindeer epithelium Ab.IgE|Reindeer epithelium Ab.IgE
C0549767|T201|COMP|11196-3|LNC|Hoplostethus atlanticus Ab.IgE|Hoplostethus atlanticus Ab.IgE
C0549769|T201|COMP|11197-1|LNC|Sardina pilchardus Ab.IgE|Sardina pilchardus Ab.IgE
C0549770|T201|COMP|10951-2|LNC|Sericin Ab.IgE|Sericin Ab.IgE
C0549771|T201|COMP|10922-3|LNC|Bovine serum albumin Ab.IgE|Bovine serum albumin Ab.IgE
C0549772|T201|COMP|11198-9|LNC|Shark Ab.IgE|Shark Ab.IgE
C0549773|T201|COMP|11199-7|LNC|Silver Ab.IgE|Silver Ab.IgE
C0549774|T201|COMP|11200-3|LNC|Helix aspersa Ab.IgE|Helix aspersa Ab.IgE
C0549775|T201|COMP|10963-7|LNC|Spondylocladium citrovirens Ab.IgE|Spondylocladium citrovirens Ab.IgE
C0549776|T201|COMP|11201-1|LNC|Succinylcholine Ab.IgE|Succinylcholine Ab.IgE
C0549777|T201|COMP|10952-0|LNC|Swine urine proteins Ab.IgE|Swine urine proteins Ab.IgE
C0549778|T201|COMP|11202-9|LNC|Artemisia dracunculus Ab.IgE|Artemisia dracunculus Ab.IgE
C0549779|T201|COMP|10932-2|LNC|Tetramin Ab.IgE|Tetramin Ab.IgE
C0549780|T201|COMP|10953-8|LNC|Phleum pratense Ab.IgG|Phleum pratense Ab.IgG
C0549781|T201|COMP|11203-7|LNC|Trichosporon pullulans Ab.IgE|Trichosporon pullulans Ab.IgE
C0549782|T201|COMP|11204-5|LNC|Ulocladium chartarum Ab.IgE|Ulocladium chartarum Ab.IgE
C0549783|T201|COMP|13179-7|LNC|Juglans regia Ab.IgG|Juglans regia Ab.IgG
C0549784|T201|COMP|6198-6|LNC|Polistes spp Ab.IgE|Polistes spp Ab.IgE
C0549785|T201|COMP|13176-3|LNC|Wasp venom Ab.IgE|Wasp venom Ab.IgE
C0549786|T201|COMP|13178-9|LNC|Wasp venom Ab.IgG|Wasp venom Ab.IgG
C0549787|T201|COMP|11174-0|LNC|Sitophilus granarius Ab.IgE|Sitophilus granarius Ab.IgE
C0549788|T201|COMP|11281-3|LNC|Auer rods|Auer rods
C0549789|T201|COMP|13330-6|LNC|Barr bodies|Barr bodies
C0549790|T201|COMP|12179-8|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0549791|T201|COMP|11105-4|LNC|Basophils/100 cells|Basophils/100 cells
C0549792|T201|COMP|11150-0|LNC|Blasts/100 cells|Blasts/100 cells
C0549793|T201|COMP|11280-5|LNC|Cabot rings|Cabot rings
C0549794|T201|COMP|12182-2|LNC|Cells|Cells
C0549795|T201|COMP|11282-1|LNC|Cells counted.total|Cells counted.total
C0549796|T201|COMP|11274-8|LNC|Elliptocytes|Elliptocytes
C0549797|T201|COMP|12209-3|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0549798|T201|COMP|11152-6|LNC|Eosinophils/100 cells|Eosinophils/100 cells
C0549799|T201|COMP|11106-2|LNC|Eosinophils/100 cells|Eosinophils/100 cells
C0549800|T201|COMP|12211-9|LNC|Epithelial cells|Epithelial cells
C0549801|T201|COMP|11131-0|LNC|Erythroblasts early/100 cells|Erythroblasts early/100 cells
C0549802|T201|COMP|11136-9|LNC|Erythroblasts late/100 erythrocytes|Erythroblasts late/100 erythrocytes
C0549803|T201|COMP|11137-7|LNC|Erythroblasts mid/100 erythrocytes|Erythroblasts mid/100 erythrocytes
C0549804|T201|COMP|11273-0|LNC|Erythrocytes|Erythrocytes
C0549805|T201|COMP|11127-8|LNC|Erythrocytes|Erythrocytes
C0549806|T201|COMP|11156-7|LNC|Leukocyte morphology finding|Leukocyte morphology finding
C0549807|T201|COMP|12226-7|LNC|Leukocytes|Leukocytes
C0549808|T201|COMP|11157-5|LNC|Leukocytes|Leukocytes
C0549809|T201|COMP|12224-2|LNC|Leukocytes|Leukocytes
C0549810|T201|COMP|12225-9|LNC|Leukocytes|Leukocytes
C0549811|T201|COMP|13349-6|LNC|Leukocytes|Leukocytes
C0549812|T201|COMP|13351-2|LNC|Leukocytes other|Leukocytes other
C0549813|T201|COMP|13046-8|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C0549814|T201|COMP|11107-0|LNC|Lymphocytes.variant/100 cells|Lymphocytes.variant/100 cells
C0549815|T201|COMP|11275-5|LNC|Lymphocytes.large granular/100 leukocytes|Lymphocytes.large granular/100 leukocytes
C0549816|T201|COMP|11031-2|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0549817|T201|COMP|11108-8|LNC|Lymphocytes/100 cells|Lymphocytes/100 cells
C0549818|T201|COMP|12229-1|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C0549819|T201|COMP|12230-9|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C0549820|T201|COMP|11109-6|LNC|Mast cells/100 cells|Mast cells/100 cells
C0549821|T201|COMP|11110-4|LNC|Megakaryocytes/100 cells|Megakaryocytes/100 cells
C0549822|T201|COMP|12233-3|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C0549823|T201|COMP|12234-1|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C0549824|T201|COMP|11111-2|LNC|Metamyelocytes/100 cells|Metamyelocytes/100 cells
C0549825|T201|COMP|11112-0|LNC|Monocytes/100 cells|Monocytes/100 cells
C0549826|T201|COMP|12236-6|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0549827|T201|COMP|11113-8|LNC|Myeloblasts/100 cells|Myeloblasts/100 cells
C0549828|T201|COMP|11114-6|LNC|Myelocytes/100 cells|Myelocytes/100 cells
C0549829|T201|COMP|11138-5|LNC|Myeloid cells/Erythroid cells|Myeloid cells/Erythroid cells
C0549830|T201|COMP|11128-6|LNC|Neutrophils.segmented/100 cells|Neutrophils.segmented/100 cells
C0549831|T201|COMP|12278-8|LNC|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0549832|T201|COMP|13354-6|LNC|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0549833|T201|COMP|11103-9|LNC|Neutrophils.band form/100 cells|Neutrophils.band form/100 cells
C0549834|T201|COMP|11115-3|LNC|Neutrophils/100 cells|Neutrophils/100 cells
C0549835|T201|COMP|11104-7|LNC|Normoblasts.basophilic/100 cells|Normoblasts.basophilic/100 cells
C0549836|T201|COMP|11116-1|LNC|Normoblasts.orthochromic/100 cells|Normoblasts.orthochromic/100 cells
C0549837|T201|COMP|11119-5|LNC|Normoblasts.polychromatophilic/100 cells|Normoblasts.polychromatophilic/100 cells
C0549838|T201|COMP|12241-6|LNC|Osmotic fragility|Osmotic fragility
C0549839|T201|COMP|11117-9|LNC|Plasma cells.immature/100 cells|Plasma cells.immature/100 cells
C0549840|T201|COMP|13047-6|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C0549841|T201|COMP|11118-7|LNC|Plasma cells/100 cells|Plasma cells/100 cells
C0549842|T201|COMP|11125-2|LNC|Platelet morphology finding|Platelet morphology finding
C0549843|T201|COMP|13057-5|LNC|Platelets|Platelets
C0549844|T201|COMP|11126-0|LNC|Platelets|Platelets
C0549845|T201|COMP|13056-7|LNC|Platelets|Platelets
C0549846|T201|COMP|12244-0|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0549847|T201|COMP|11129-4|LNC|Pronormoblasts|Pronormoblasts
C0549848|T201|COMP|11120-3|LNC|Promyelocytes/100 cells|Promyelocytes/100 cells
C0549849|T201|COMP|11121-1|LNC|Prolymphocytes/100 cells|Prolymphocytes/100 cells
C0549850|T201|COMP|11122-9|LNC|Promonocytes/100 cells|Promonocytes/100 cells
C0549851|T201|COMP|11123-7|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C0549852|T201|COMP|11124-5|LNC|Pronormoblasts/100 cells|Pronormoblasts/100 cells
C0549853|T201|COMP|12248-1|LNC|Epithelial cells.renal|Epithelial cells.renal
C0549855|T201|COMP|13048-4|LNC|Sezary cells|Sezary cells
C0549856|T201|COMP|12258-0|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C0549857|T201|COMP|11276-3|LNC|Tubular cells|Tubular cells
C0549858|T201|COMP|13355-3|LNC|Unspecified cells/100 leukocytes|Unspecified cells/100 leukocytes
C0549859|T201|COMP|12273-9|LNC|Xanthochromia|Xanthochromia
C0549860|T201|COMP|13310-8|LNC|Kell group Ag|Kell group Ag
C0549861|T201|COMP|13309-0|LNC|Duffy group Ag|Duffy group Ag
C0549862|T201|COMP|11130-2|LNC|Lymphocytes B|Lymphocytes B
C0549863|T201|COMP|13331-4|LNC|Cells.CD2+CD26+/100 cells|Cells.CD2+CD26+/100 cells
C0549864|T201|COMP|13333-0|LNC|Cells.CD3+CD25+/100 cells|Cells.CD3+CD25+/100 cells
C0549865|T201|COMP|13341-3|LNC|Cells.CD3+CD25+/100 cells|Cells.CD3+CD25+/100 cells
C0549866|T201|COMP|13342-1|LNC|Cells.CD3+CD26+/100 cells|Cells.CD3+CD26+/100 cells
C0549867|T201|COMP|13340-5|LNC|Cells.CD3+CD38+/100 cells|Cells.CD3+CD38+/100 cells
C0549868|T201|COMP|13346-2|LNC|Cells.CD35/100 cells|Cells.CD35/100 cells
C0549869|T201|COMP|13491-6|LNC|Cells.CD4+CD25+|Cells.CD4+CD25+
C0549870|T201|COMP|13332-2|LNC|Cells.CD4+CD25+/100 cells|Cells.CD4+CD25+/100 cells
C0549871|T201|COMP|13335-5|LNC|Cells.CD4+CD29+/100 cells|Cells.CD4+CD29+/100 cells
C0549872|T201|COMP|13336-3|LNC|Cells.CD4+CD45RA+/100 cells|Cells.CD4+CD45RA+/100 cells
C0549873|T201|COMP|13492-4|LNC|Cells.CD4+HLA-DR+|Cells.CD4+HLA-DR+
C0549874|T201|COMP|13343-9|LNC|Cells.CD4+HLA-DR+/100 cells|Cells.CD4+HLA-DR+/100 cells
C0549875|T201|COMP|13345-4|LNC|Cells.CD8+CD11b+/100 cells|Cells.CD8+CD11b+/100 cells
C0549876|T201|COMP|13493-2|LNC|Cells.CD8+CD25+|Cells.CD8+CD25+
C0549877|T201|COMP|13334-8|LNC|Cells.CD8+CD25+/100 cells|Cells.CD8+CD25+/100 cells
C0549878|T201|COMP|13344-7|LNC|Cells.CD8+CD38+/100 cells|Cells.CD8+CD38+/100 cells
C0549879|T201|COMP|13339-7|LNC|Cells.CD8+CD56+/100 cells|Cells.CD8+CD56+/100 cells
C0549880|T201|COMP|13338-9|LNC|Cells.CD8+CD57+/100 cells|Cells.CD8+CD57+/100 cells
C0549881|T201|COMP|13337-1|LNC|Cells.CD8+HLA-DR+/100 cells|Cells.CD8+HLA-DR+/100 cells
C0549888|T201|COMP|13040-1|LNC|C peptide^1.5H post XXX challenge|C peptide^1.5H post XXX challenge
C0549889|T201|COMP|13039-3|LNC|C peptide^1H post XXX challenge|C peptide^1H post XXX challenge
C0549890|T201|COMP|13042-7|LNC|C peptide^2.5H post XXX challenge|C peptide^2.5H post XXX challenge
C0549891|T201|COMP|13041-9|LNC|C peptide^2H post XXX challenge|C peptide^2H post XXX challenge
C0549892|T201|COMP|13032-8|LNC|C peptide^2nd specimen post XXX challenge|C peptide^2nd specimen post XXX challenge
C0549893|T201|COMP|13038-5|LNC|C peptide^30M post XXX challenge|C peptide^30M post XXX challenge
C0549894|T201|COMP|13043-5|LNC|C peptide^3H post XXX challenge|C peptide^3H post XXX challenge
C0549895|T201|COMP|13033-6|LNC|C peptide^3rd specimen post XXX challenge|C peptide^3rd specimen post XXX challenge
C0549896|T201|COMP|13034-4|LNC|C peptide^4th specimen post XXX challenge|C peptide^4th specimen post XXX challenge
C0549897|T201|COMP|13044-3|LNC|C peptide^5H post XXX challenge|C peptide^5H post XXX challenge
C0549898|T201|COMP|13035-1|LNC|C peptide^5th specimen post XXX challenge|C peptide^5th specimen post XXX challenge
C0549899|T201|COMP|13045-0|LNC|C peptide^6H post XXX challenge|C peptide^6H post XXX challenge
C0549900|T201|COMP|13036-9|LNC|C peptide^6th specimen post XXX challenge|C peptide^6th specimen post XXX challenge
C0549901|T201|COMP|13037-7|LNC|C peptide^post CFst|C peptide^post CFst
C0549902|T201|COMP|12506-2|LNC|Calcitonin^2nd specimen post XXX challenge|Calcitonin^2nd specimen post XXX challenge
C0549903|T201|COMP|12507-0|LNC|Calcitonin^3rd specimen post XXX challenge|Calcitonin^3rd specimen post XXX challenge
C0549904|T201|COMP|12508-8|LNC|Calcitonin^4th specimen post XXX challenge|Calcitonin^4th specimen post XXX challenge
C0549905|T201|COMP|12509-6|LNC|Calcitonin^5th specimen post XXX challenge|Calcitonin^5th specimen post XXX challenge
C0549906|T201|COMP|12510-4|LNC|Calcitonin^6th specimen post XXX challenge|Calcitonin^6th specimen post XXX challenge
C0549907|T201|COMP|12516-1|LNC|Catecholamines^2nd specimen post XXX challenge|Catecholamines^2nd specimen post XXX challenge
C0549908|T201|COMP|12522-9|LNC|Catecholamines^2nd specimen post XXX challenge|Catecholamines^2nd specimen post XXX challenge
C0549909|T201|COMP|12523-7|LNC|Catecholamines^3rd specimen post XXX challenge|Catecholamines^3rd specimen post XXX challenge
C0549910|T201|COMP|12517-9|LNC|Catecholamines^3rd specimen post XXX challenge|Catecholamines^3rd specimen post XXX challenge
C0549911|T201|COMP|12524-5|LNC|Catecholamines^4th specimen post XXX challenge|Catecholamines^4th specimen post XXX challenge
C0549912|T201|COMP|12518-7|LNC|Catecholamines^4th specimen post XXX challenge|Catecholamines^4th specimen post XXX challenge
C0549913|T201|COMP|12519-5|LNC|Catecholamines^5th specimen post XXX challenge|Catecholamines^5th specimen post XXX challenge
C0549914|T201|COMP|12520-3|LNC|Catecholamines^6th specimen post XXX challenge|Catecholamines^6th specimen post XXX challenge
C0549915|T201|COMP|12521-1|LNC|Catecholamines^7th specimen post XXX challenge|Catecholamines^7th specimen post XXX challenge
C0549916|T201|COMP|12458-6|LNC|Corticotropin^2nd specimen post XXX challenge|Corticotropin^2nd specimen post XXX challenge
C0549917|T201|COMP|12459-4|LNC|Corticotropin^3rd specimen post XXX challenge|Corticotropin^3rd specimen post XXX challenge
C0549918|T201|COMP|12460-2|LNC|Corticotropin^4th specimen post XXX challenge|Corticotropin^4th specimen post XXX challenge
C0549919|T201|COMP|12461-0|LNC|Corticotropin^5th specimen post XXX challenge|Corticotropin^5th specimen post XXX challenge
C0549920|T201|COMP|12462-8|LNC|Corticotropin^6th specimen post XXX challenge|Corticotropin^6th specimen post XXX challenge
C0549921|T201|COMP|12463-6|LNC|Corticotropin^7th specimen post XXX challenge|Corticotropin^7th specimen post XXX challenge
C0549922|T201|COMP|12464-4|LNC|Corticotropin^8th specimen post XXX challenge|Corticotropin^8th specimen post XXX challenge
C0549923|T201|COMP|12565-8|LNC|Cortisol^10th specimen post XXX challenge|Cortisol^10th specimen post XXX challenge
C0549924|T201|COMP|12567-4|LNC|Cortisol^1H post XXX challenge|Cortisol^1H post XXX challenge
C0549925|T201|COMP|12569-0|LNC|Cortisol^2.5H post XXX challenge|Cortisol^2.5H post XXX challenge
C0549926|T201|COMP|12568-2|LNC|Cortisol^20M post XXX challenge|Cortisol^20M post XXX challenge
C0549927|T201|COMP|12557-5|LNC|Cortisol^2nd specimen post XXX challenge|Cortisol^2nd specimen post XXX challenge
C0549928|T201|COMP|12566-6|LNC|Cortisol^30M post XXX challenge|Cortisol^30M post XXX challenge
C0549929|T201|COMP|12558-3|LNC|Cortisol^3rd specimen post XXX challenge|Cortisol^3rd specimen post XXX challenge
C0549930|T201|COMP|12559-1|LNC|Cortisol^4th specimen post XXX challenge|Cortisol^4th specimen post XXX challenge
C0549931|T201|COMP|12560-9|LNC|Cortisol^5th specimen post XXX challenge|Cortisol^5th specimen post XXX challenge
C0549932|T201|COMP|12561-7|LNC|Cortisol^6th specimen post XXX challenge|Cortisol^6th specimen post XXX challenge
C0549933|T201|COMP|12562-5|LNC|Cortisol^7th specimen post XXX challenge|Cortisol^7th specimen post XXX challenge
C0549934|T201|COMP|12563-3|LNC|Cortisol^8th specimen post XXX challenge|Cortisol^8th specimen post XXX challenge
C0549935|T201|COMP|12564-1|LNC|Cortisol^9th specimen post XXX challenge|Cortisol^9th specimen post XXX challenge
C0549936|T201|COMP|12570-8|LNC|Cortisol^post XXX challenge|Cortisol^post XXX challenge
C0549937|T201|COMP|13432-0|LNC|DOPamine^2nd specimen post XXX challenge|DOPamine^2nd specimen post XXX challenge
C0549938|T201|COMP|13433-8|LNC|DOPamine^3rd specimen post XXX challenge|DOPamine^3rd specimen post XXX challenge
C0549939|T201|COMP|13434-6|LNC|DOPamine^4th specimen post XXX challenge|DOPamine^4th specimen post XXX challenge
C0549940|T201|COMP|13435-3|LNC|DOPamine^5th specimen post XXX challenge|DOPamine^5th specimen post XXX challenge
C0549941|T201|COMP|13436-1|LNC|DOPamine^6th specimen post XXX challenge|DOPamine^6th specimen post XXX challenge
C0549942|T201|COMP|13437-9|LNC|DOPamine^7th specimen post XXX challenge|DOPamine^7th specimen post XXX challenge
C0549943|T201|COMP|12529-4|LNC|EPINEPHrine^2H post XXX challenge|EPINEPHrine^2H post XXX challenge
C0549944|T201|COMP|13420-5|LNC|EPINEPHrine^2nd specimen post XXX challenge|EPINEPHrine^2nd specimen post XXX challenge
C0549945|T201|COMP|13421-3|LNC|EPINEPHrine^3rd specimen post XXX challenge|EPINEPHrine^3rd specimen post XXX challenge
C0549946|T201|COMP|13422-1|LNC|EPINEPHrine^4th specimen post XXX challenge|EPINEPHrine^4th specimen post XXX challenge
C0549947|T201|COMP|13423-9|LNC|EPINEPHrine^5th specimen post XXX challenge|EPINEPHrine^5th specimen post XXX challenge
C0549948|T201|COMP|13424-7|LNC|EPINEPHrine^6th specimen post XXX challenge|EPINEPHrine^6th specimen post XXX challenge
C0549949|T201|COMP|13425-4|LNC|EPINEPHrine^7th specimen post XXX challenge|EPINEPHrine^7th specimen post XXX challenge
C0549950|T201|COMP|12596-3|LNC|Estradiol^3H post XXX challenge|Estradiol^3H post XXX challenge
C0549951|T201|COMP|12597-1|LNC|Estrogen^2nd specimen post XXX challenge|Estrogen^2nd specimen post XXX challenge
C0549952|T201|COMP|12667-2|LNC|Follitropin^5th specimen post XXX challenge|Follitropin^5th specimen post XXX challenge
C0549953|T201|COMP|12661-5|LNC|Follitropin^10M post XXX challenge|Follitropin^10M post XXX challenge
C0549954|T201|COMP|12662-3|LNC|Follitropin^20M post XXX challenge|Follitropin^20M post XXX challenge
C0549955|T201|COMP|12664-9|LNC|Follitropin^2nd specimen post XXX challenge|Follitropin^2nd specimen post XXX challenge
C0549956|T201|COMP|12660-7|LNC|Follitropin^3H post XXX challenge|Follitropin^3H post XXX challenge
C0549957|T201|COMP|12665-6|LNC|Follitropin^3rd specimen post XXX challenge|Follitropin^3rd specimen post XXX challenge
C0549958|T201|COMP|12663-1|LNC|Follitropin^40M post XXX challenge|Follitropin^40M post XXX challenge
C0549959|T201|COMP|12666-4|LNC|Follitropin^4th specimen post XXX challenge|Follitropin^4th specimen post XXX challenge
C0549960|T201|COMP|12668-0|LNC|Follitropin^6th specimen post XXX challenge|Follitropin^6th specimen post XXX challenge
C0549961|T201|COMP|12669-8|LNC|Follitropin^7th specimen post XXX challenge|Follitropin^7th specimen post XXX challenge
C0549962|T201|COMP|12670-6|LNC|Follitropin^8th specimen post XXX challenge|Follitropin^8th specimen post XXX challenge
C0549963|T201|COMP|12671-4|LNC|Follitropin^9th specimen post XXX challenge|Follitropin^9th specimen post XXX challenge
C0549964|T201|COMP|12645-8|LNC|Glucose^10H post XXX challenge|Glucose^10H post XXX challenge
C0549965|T201|COMP|12654-0|LNC|Glucose^10M post XXX challenge|Glucose^10M post XXX challenge
C0549966|T201|COMP|12651-6|LNC|Glucose^10M pre XXX challenge|Glucose^10M pre XXX challenge
C0549967|T201|COMP|12622-7|LNC|Glucose^10th specimen post XXX challenge|Glucose^10th specimen post XXX challenge
C0549968|T201|COMP|12623-5|LNC|Glucose^11th specimen post XXX challenge|Glucose^11th specimen post XXX challenge
C0549969|T201|COMP|12647-4|LNC|Glucose^12H post XXX challenge|Glucose^12H post XXX challenge
C0549970|T201|COMP|12624-3|LNC|Glucose^12th specimen post XXX challenge|Glucose^12th specimen post XXX challenge
C0549971|T201|COMP|12625-0|LNC|Glucose^13th specimen post XXX challenge|Glucose^13th specimen post XXX challenge
C0549972|T201|COMP|12626-8|LNC|Glucose^14th specimen post XXX challenge|Glucose^14th specimen post XXX challenge
C0549973|T201|COMP|10832-4|LNC|Glucose^15M post 50 g lactose PO|Glucose^15M post 50 g lactose PO
C0549974|T201|COMP|12639-1|LNC|Glucose^15M post XXX challenge|Glucose^15M post XXX challenge
C0549975|T201|COMP|12648-2|LNC|Glucose^15M post dose lactose PO|Glucose^15M post dose lactose PO
C0549976|T201|COMP|12627-6|LNC|Glucose^15th specimen post XXX challenge|Glucose^15th specimen post XXX challenge
C0549977|T201|COMP|12646-6|LNC|Glucose^1H post XXX challenge|Glucose^1H post XXX challenge
C0549978|T201|COMP|12615-1|LNC|Glucose^1st specimen post XXX challenge|Glucose^1st specimen post XXX challenge
C0549979|T201|COMP|10966-0|LNC|Glucose^2.5H post 75 g glucose PO|Glucose^2.5H post 75 g glucose PO
C0549980|T201|COMP|12655-7|LNC|Glucose^20M post XXX challenge|Glucose^20M post XXX challenge
C0549981|T201|COMP|12610-2|LNC|Glucose^2H post XXX challenge|Glucose^2H post XXX challenge
C0549982|T201|COMP|12652-4|LNC|Glucose^2M post XXX challenge|Glucose^2M post XXX challenge
C0549983|T201|COMP|12616-9|LNC|Glucose^2nd specimen post XXX challenge|Glucose^2nd specimen post XXX challenge
C0549984|T201|COMP|10967-8|LNC|Glucose^3.5H post 75 g glucose PO|Glucose^3.5H post 75 g glucose PO
C0549985|T201|COMP|12650-8|LNC|Glucose^3.5H post dose lactose PO|Glucose^3.5H post dose lactose PO
C0549986|T201|COMP|12617-7|LNC|Glucose^3rd specimen post XXX challenge|Glucose^3rd specimen post XXX challenge
C0549987|T201|COMP|10968-6|LNC|Glucose^4.5H post 75 g glucose PO|Glucose^4.5H post 75 g glucose PO
C0549988|T201|COMP|12657-3|LNC|Glucose^40M post XXX challenge|Glucose^40M post XXX challenge
C0549989|T201|COMP|11032-0|LNC|Glucose^45M post 50 g lactose PO|Glucose^45M post 50 g lactose PO
C0549990|T201|COMP|12656-5|LNC|Glucose^4M post XXX challenge|Glucose^4M post XXX challenge
C0549991|T201|COMP|12618-5|LNC|Glucose^4th specimen post XXX challenge|Glucose^4th specimen post XXX challenge
C0549992|T201|COMP|12658-1|LNC|Glucose^50M post XXX challenge|Glucose^50M post XXX challenge
C0549993|T201|COMP|12619-3|LNC|Glucose^5th specimen post XXX challenge|Glucose^5th specimen post XXX challenge
C0549994|T201|COMP|12640-9|LNC|Glucose^6.5H post XXX challenge|Glucose^6.5H post XXX challenge
C0549995|T201|COMP|12620-1|LNC|Glucose^6th specimen post XXX challenge|Glucose^6th specimen post XXX challenge
C0549996|T201|COMP|12649-0|LNC|Glucose^6th specimen post dose lactose|Glucose^6th specimen post dose lactose
C0549997|T201|COMP|12642-5|LNC|Glucose^7.5H post XXX challenge|Glucose^7.5H post XXX challenge
C0549998|T201|COMP|12659-9|LNC|Glucose^70M post XXX challenge|Glucose^70M post XXX challenge
C0549999|T201|COMP|12641-7|LNC|Glucose^7H post XXX challenge|Glucose^7H post XXX challenge
C0550000|T201|COMP|12614-4|LNC|Glucose^7H post meal|Glucose^7H post meal
C0550001|T201|COMP|12643-3|LNC|Glucose^8H post XXX challenge|Glucose^8H post XXX challenge
C0550002|T201|COMP|12653-2|LNC|Glucose^8M post XXX challenge|Glucose^8M post XXX challenge
C0550003|T201|COMP|12637-5|LNC|Glucose^8th specimen post XXX challenge|Glucose^8th specimen post XXX challenge
C0550004|T201|COMP|12644-1|LNC|Glucose^9H post XXX challenge|Glucose^9H post XXX challenge
C0550005|T201|COMP|12621-9|LNC|Glucose^9th specimen post XXX challenge|Glucose^9th specimen post XXX challenge
C0550006|T201|COMP|12638-3|LNC|Glucose^pre dose lactose PO|Glucose^pre dose lactose PO
C0550010|T201|COMP|12747-2|LNC|Insulin^3.5H post XXX challenge|Insulin^3.5H post XXX challenge
C0550011|T201|COMP|12754-8|LNC|Insulin^10H post XXX challenge|Insulin^10H post XXX challenge
C0550012|T201|COMP|12755-5|LNC|Insulin^11H post XXX challenge|Insulin^11H post XXX challenge
C0550013|T201|COMP|12756-3|LNC|Insulin^12H post XXX challenge|Insulin^12H post XXX challenge
C0550014|T201|COMP|12762-1|LNC|Insulin^15M post XXX challenge|Insulin^15M post XXX challenge
C0550015|T201|COMP|12763-9|LNC|Insulin^19M post XXX challenge|Insulin^19M post XXX challenge
C0550016|T201|COMP|12764-7|LNC|Insulin^22M post XXX challenge|Insulin^22M post XXX challenge
C0550017|T201|COMP|12759-7|LNC|Insulin^2M post XXX challenge|Insulin^2M post XXX challenge
C0550018|T201|COMP|12739-9|LNC|Insulin^2nd specimen post XXX challenge|Insulin^2nd specimen post XXX challenge
C0550019|T201|COMP|12740-7|LNC|Insulin^3rd specimen post XXX challenge|Insulin^3rd specimen post XXX challenge
C0550020|T201|COMP|12748-0|LNC|Insulin^4.5H post XXX challenge|Insulin^4.5H post XXX challenge
C0550021|T201|COMP|12765-4|LNC|Insulin^40M post XXX challenge|Insulin^40M post XXX challenge
C0550022|T201|COMP|12766-2|LNC|Insulin^45M post XXX challenge|Insulin^45M post XXX challenge
C0550023|T201|COMP|12760-5|LNC|Insulin^4M post XXX challenge|Insulin^4M post XXX challenge
C0550024|T201|COMP|12741-5|LNC|Insulin^4th specimen post XXX challenge|Insulin^4th specimen post XXX challenge
C0550025|T201|COMP|12749-8|LNC|Insulin^5.5H post XXX challenge|Insulin^5.5H post XXX challenge
C0550026|T201|COMP|12767-0|LNC|Insulin^50M post XXX challenge|Insulin^50M post XXX challenge
C0550027|T201|COMP|12742-3|LNC|Insulin^5th specimen post XXX challenge|Insulin^5th specimen post XXX challenge
C0550028|T201|COMP|12743-1|LNC|Insulin^6th specimen post XXX challenge|Insulin^6th specimen post XXX challenge
C0550029|T201|COMP|12751-4|LNC|Insulin^7.5H post XXX challenge|Insulin^7.5H post XXX challenge
C0550030|T201|COMP|12768-8|LNC|Insulin^70M post XXX challenge|Insulin^70M post XXX challenge
C0550031|T201|COMP|12750-6|LNC|Insulin^7H post XXX challenge|Insulin^7H post XXX challenge
C0550032|T201|COMP|12744-9|LNC|Insulin^7th specimen post XXX challenge|Insulin^7th specimen post XXX challenge
C0550033|T201|COMP|12752-2|LNC|Insulin^8H post XXX challenge|Insulin^8H post XXX challenge
C0550034|T201|COMP|12761-3|LNC|Insulin^8M post XXX challenge|Insulin^8M post XXX challenge
C0550035|T201|COMP|12745-6|LNC|Insulin^8th specimen post XXX challenge|Insulin^8th specimen post XXX challenge
C0550036|T201|COMP|12753-0|LNC|Insulin^9H post XXX challenge|Insulin^9H post XXX challenge
C0550037|T201|COMP|12746-4|LNC|Insulin^9th specimen post XXX challenge|Insulin^9th specimen post XXX challenge
C0550038|T201|COMP|12758-9|LNC|Insulin^15M pre XXX challenge|Insulin^15M pre XXX challenge
C0550039|T201|COMP|12757-1|LNC|Insulin^30M pre XXX challenge|Insulin^30M pre XXX challenge
C0550040|T201|COMP|12738-1|LNC|Insulin^pre XXX challenge|Insulin^pre XXX challenge
C0550041|T201|COMP|10833-2|LNC|Insulin^7H post 75 g glucose PO|Insulin^7H post 75 g glucose PO
C0550042|T201|COMP|12448-7|LNC|Ketones^post CFst|Ketones^post CFst
C0550043|T201|COMP|12449-5|LNC|Ketones^1H post XXX challenge|Ketones^1H post XXX challenge
C0550044|T201|COMP|12450-3|LNC|Ketones^2H post XXX challenge|Ketones^2H post XXX challenge
C0550045|T201|COMP|12451-1|LNC|Ketones^3H post XXX challenge|Ketones^3H post XXX challenge
C0550046|T201|COMP|12672-2|LNC|Lutropin^10M post XXX challenge|Lutropin^10M post XXX challenge
C0550047|T201|COMP|12674-8|LNC|Lutropin^15M pre XXX challenge|Lutropin^15M pre XXX challenge
C0550048|T201|COMP|12675-5|LNC|Lutropin^20M post XXX challenge|Lutropin^20M post XXX challenge
C0550049|T201|COMP|12677-1|LNC|Lutropin^2nd specimen post XXX challenge|Lutropin^2nd specimen post XXX challenge
C0550050|T201|COMP|12673-0|LNC|Lutropin^3H post XXX challenge|Lutropin^3H post XXX challenge
C0550051|T201|COMP|12678-9|LNC|Lutropin^3rd specimen post XXX challenge|Lutropin^3rd specimen post XXX challenge
C0550052|T201|COMP|12676-3|LNC|Lutropin^40M post XXX challenge|Lutropin^40M post XXX challenge
C0550053|T201|COMP|12679-7|LNC|Lutropin^4th specimen post XXX challenge|Lutropin^4th specimen post XXX challenge
C0550054|T201|COMP|12680-5|LNC|Lutropin^5th specimen post XXX challenge|Lutropin^5th specimen post XXX challenge
C0550055|T201|COMP|12681-3|LNC|Lutropin^6th specimen post XXX challenge|Lutropin^6th specimen post XXX challenge
C0550056|T201|COMP|12682-1|LNC|Lutropin^7th specimen post XXX challenge|Lutropin^7th specimen post XXX challenge
C0550057|T201|COMP|12683-9|LNC|Lutropin^8th specimen post XXX challenge|Lutropin^8th specimen post XXX challenge
C0550058|T201|COMP|12684-7|LNC|Lutropin^9th specimen post XXX challenge|Lutropin^9th specimen post XXX challenge
C0550059|T201|COMP|12832-2|LNC|Prolactin^10M post XXX challenge|Prolactin^10M post XXX challenge
C0550060|T201|COMP|12831-4|LNC|Prolactin^10th specimen post XXX challenge|Prolactin^10th specimen post XXX challenge
C0550061|T201|COMP|12834-8|LNC|Prolactin^15M post XXX challenge|Prolactin^15M post XXX challenge
C0550062|T201|COMP|12833-0|LNC|Prolactin^20M post XXX challenge|Prolactin^20M post XXX challenge
C0550063|T201|COMP|12823-1|LNC|Prolactin^2nd specimen post XXX challenge|Prolactin^2nd specimen post XXX challenge
C0550064|T201|COMP|12824-9|LNC|Prolactin^3rd specimen post XXX challenge|Prolactin^3rd specimen post XXX challenge
C0550065|T201|COMP|12835-5|LNC|Prolactin^45M post XXX challenge|Prolactin^45M post XXX challenge
C0550066|T201|COMP|12825-6|LNC|Prolactin^4th specimen post XXX challenge|Prolactin^4th specimen post XXX challenge
C0550067|T201|COMP|12826-4|LNC|Prolactin^5th specimen post XXX challenge|Prolactin^5th specimen post XXX challenge
C0550068|T201|COMP|12827-2|LNC|Prolactin^6th specimen post XXX challenge|Prolactin^6th specimen post XXX challenge
C0550069|T201|COMP|12828-0|LNC|Prolactin^7th specimen post XXX challenge|Prolactin^7th specimen post XXX challenge
C0550070|T201|COMP|12829-8|LNC|Prolactin^8th specimen post XXX challenge|Prolactin^8th specimen post XXX challenge
C0550071|T201|COMP|12830-6|LNC|Prolactin^9th specimen post XXX challenge|Prolactin^9th specimen post XXX challenge
C0550072|T201|COMP|12525-2|LNC|Norepinephrine^1H post XXX challenge|Norepinephrine^1H post XXX challenge
C0550073|T201|COMP|12526-0|LNC|Norepinephrine^2H post XXX challenge|Norepinephrine^2H post XXX challenge
C0550074|T201|COMP|13426-2|LNC|Norepinephrine^2nd specimen post XXX challenge|Norepinephrine^2nd specimen post XXX challenge
C0550075|T201|COMP|12527-8|LNC|Norepinephrine^3H post XXX challenge|Norepinephrine^3H post XXX challenge
C0550076|T201|COMP|13427-0|LNC|Norepinephrine^3rd specimen post XXX challenge|Norepinephrine^3rd specimen post XXX challenge
C0550077|T201|COMP|12528-6|LNC|Norepinephrine^4H post XXX challenge|Norepinephrine^4H post XXX challenge
C0550078|T201|COMP|13428-8|LNC|Norepinephrine^4th specimen post XXX challenge|Norepinephrine^4th specimen post XXX challenge
C0550079|T201|COMP|13429-6|LNC|Norepinephrine^5th specimen post XXX challenge|Norepinephrine^5th specimen post XXX challenge
C0550080|T201|COMP|13430-4|LNC|Norepinephrine^6th specimen post XXX challenge|Norepinephrine^6th specimen post XXX challenge
C0550081|T201|COMP|13431-2|LNC|Norepinephrine^7th specimen post XXX challenge|Norepinephrine^7th specimen post XXX challenge
C0550082|T201|COMP|12798-5|LNC|Oxalate^10th specimen post XXX challenge|Oxalate^10th specimen post XXX challenge
C0550083|T201|COMP|12790-2|LNC|Oxalate^2nd specimen post XXX challenge|Oxalate^2nd specimen post XXX challenge
C0550084|T201|COMP|12791-0|LNC|Oxalate^3rd specimen post XXX challenge|Oxalate^3rd specimen post XXX challenge
C0550085|T201|COMP|12792-8|LNC|Oxalate^4th specimen post XXX challenge|Oxalate^4th specimen post XXX challenge
C0550086|T201|COMP|12793-6|LNC|Oxalate^5th specimen post XXX challenge|Oxalate^5th specimen post XXX challenge
C0550087|T201|COMP|12794-4|LNC|Oxalate^6th specimen post XXX challenge|Oxalate^6th specimen post XXX challenge
C0550088|T201|COMP|12795-1|LNC|Oxalate^7th specimen post XXX challenge|Oxalate^7th specimen post XXX challenge
C0550089|T201|COMP|12796-9|LNC|Oxalate^8th specimen post XXX challenge|Oxalate^8th specimen post XXX challenge
C0550090|T201|COMP|12797-7|LNC|Oxalate^9th specimen post XXX challenge|Oxalate^9th specimen post XXX challenge
C0550091|T201|COMP|12822-3|LNC|Progesterone^1H post XXX challenge|Progesterone^1H post XXX challenge
C0550092|T201|COMP|12815-7|LNC|Progesterone^2nd specimen post XXX challenge|Progesterone^2nd specimen post XXX challenge
C0550093|T201|COMP|12821-5|LNC|Progesterone^30M post XXX challenge|Progesterone^30M post XXX challenge
C0550094|T201|COMP|12816-5|LNC|Progesterone^3rd specimen post XXX challenge|Progesterone^3rd specimen post XXX challenge
C0550095|T201|COMP|12817-3|LNC|Progesterone^4th specimen post XXX challenge|Progesterone^4th specimen post XXX challenge
C0550096|T201|COMP|12818-1|LNC|Progesterone^5th specimen post XXX challenge|Progesterone^5th specimen post XXX challenge
C0550097|T201|COMP|12819-9|LNC|Progesterone^6th specimen post XXX challenge|Progesterone^6th specimen post XXX challenge
C0550098|T201|COMP|12900-7|LNC|Renin^2nd specimen post XXX challenge|Renin^2nd specimen post XXX challenge
C0550099|T201|COMP|12901-5|LNC|Renin^3rd specimen post XXX challenge|Renin^3rd specimen post XXX challenge
C0550100|T201|COMP|12902-3|LNC|Renin^4th specimen post XXX challenge|Renin^4th specimen post XXX challenge
C0550101|T201|COMP|12903-1|LNC|Renin^5th specimen post XXX challenge|Renin^5th specimen post XXX challenge
C0550102|T201|COMP|12904-9|LNC|Renin^6th specimen post XXX challenge|Renin^6th specimen post XXX challenge
C0550103|T201|COMP|12905-6|LNC|Renin^7th specimen post XXX challenge|Renin^7th specimen post XXX challenge
C0550104|T201|COMP|12906-4|LNC|Renin^8th specimen post XXX challenge|Renin^8th specimen post XXX challenge
C0550105|T201|COMP|12697-9|LNC|Somatotropin^10M post XXX challenge|Somatotropin^10M post XXX challenge
C0550106|T201|COMP|12693-8|LNC|Somatotropin^10th specimen post XXX challenge|Somatotropin^10th specimen post XXX challenge
C0550107|T201|COMP|12698-7|LNC|Somatotropin^15M post XXX challenge|Somatotropin^15M post XXX challenge
C0550108|T201|COMP|12701-9|LNC|Somatotropin^2.5H post XXX challenge|Somatotropin^2.5H post XXX challenge
C0550109|T201|COMP|12699-5|LNC|Somatotropin^20M post XXX challenge|Somatotropin^20M post XXX challenge
C0550110|T201|COMP|12685-4|LNC|Somatotropin^2nd specimen post XXX challenge|Somatotropin^2nd specimen post XXX challenge
C0550111|T201|COMP|12686-2|LNC|Somatotropin^3rd specimen post XXX challenge|Somatotropin^3rd specimen post XXX challenge
C0550112|T201|COMP|12700-1|LNC|Somatotropin^45M post XXX challenge|Somatotropin^45M post XXX challenge
C0550113|T201|COMP|12687-0|LNC|Somatotropin^4th specimen post XXX challenge|Somatotropin^4th specimen post XXX challenge
C0550114|T201|COMP|12688-8|LNC|Somatotropin^5th specimen post XXX challenge|Somatotropin^5th specimen post XXX challenge
C0550115|T201|COMP|12689-6|LNC|Somatotropin^6th specimen post XXX challenge|Somatotropin^6th specimen post XXX challenge
C0550116|T201|COMP|12690-4|LNC|Somatotropin^7th specimen post XXX challenge|Somatotropin^7th specimen post XXX challenge
C0550117|T201|COMP|12691-2|LNC|Somatotropin^8th specimen post XXX challenge|Somatotropin^8th specimen post XXX challenge
C0550118|T201|COMP|12692-0|LNC|Somatotropin^9th specimen post XXX challenge|Somatotropin^9th specimen post XXX challenge
C0550119|T201|COMP|12695-3|LNC|Somatotropin^15M pre XXX challenge|Somatotropin^15M pre XXX challenge
C0550120|T201|COMP|12696-1|LNC|Somatotropin^pre XXX challenge|Somatotropin^pre XXX challenge
C0550121|T201|COMP|12694-6|LNC|Somatotropin^post XXX challenge|Somatotropin^post XXX challenge
C0550122|T201|COMP|12922-1|LNC|Testosterone^1H post XXX challenge|Testosterone^1H post XXX challenge
C0550123|T201|COMP|12921-3|LNC|Testosterone^3H post XXX challenge|Testosterone^3H post XXX challenge
C0550124|T201|COMP|12938-7|LNC|Thyrotropin^1.5H post XXX challenge|Thyrotropin^1.5H post XXX challenge
C0550125|T201|COMP|12933-8|LNC|Thyrotropin^10M post XXX challenge|Thyrotropin^10M post XXX challenge
C0550126|T201|COMP|12934-6|LNC|Thyrotropin^15M post XXX challenge|Thyrotropin^15M post XXX challenge
C0550127|T201|COMP|12935-3|LNC|Thyrotropin^20M post XXX challenge|Thyrotropin^20M post XXX challenge
C0550128|T201|COMP|12939-5|LNC|Thyrotropin^2H post XXX challenge|Thyrotropin^2H post XXX challenge
C0550129|T201|COMP|12941-1|LNC|Thyrotropin^2nd specimen post XXX challenge|Thyrotropin^2nd specimen post XXX challenge
C0550130|T201|COMP|12942-9|LNC|Thyrotropin^3rd specimen post XXX challenge|Thyrotropin^3rd specimen post XXX challenge
C0550131|T201|COMP|12936-1|LNC|Thyrotropin^40M post XXX challenge|Thyrotropin^40M post XXX challenge
C0550132|T201|COMP|12937-9|LNC|Thyrotropin^45M post XXX challenge|Thyrotropin^45M post XXX challenge
C0550133|T201|COMP|11033-8|LNC|Thyrotropin^45M post dose TRH IV|Thyrotropin^45M post dose TRH IV
C0550134|T201|COMP|12943-7|LNC|Thyrotropin^4th specimen post XXX challenge|Thyrotropin^4th specimen post XXX challenge
C0550135|T201|COMP|12944-5|LNC|Thyrotropin^5th specimen post XXX challenge|Thyrotropin^5th specimen post XXX challenge
C0550136|T201|COMP|12945-2|LNC|Thyrotropin^6th specimen post XXX challenge|Thyrotropin^6th specimen post XXX challenge
C0550137|T201|COMP|12946-0|LNC|Thyrotropin^7th specimen post XXX challenge|Thyrotropin^7th specimen post XXX challenge
C0550138|T201|COMP|12947-8|LNC|Thyrotropin^8th specimen post XXX challenge|Thyrotropin^8th specimen post XXX challenge
C0550139|T201|COMP|12948-6|LNC|Thyrotropin^9th specimen post XXX challenge|Thyrotropin^9th specimen post XXX challenge
C0550140|T201|COMP|12940-3|LNC|Thyrotropin^30M pre XXX challenge|Thyrotropin^30M pre XXX challenge
C0550141|T201|COMP|12932-0|LNC|Thyrotropin^post XXX challenge|Thyrotropin^post XXX challenge
C0550142|T201|COMP|12952-8|LNC|Thyroxine uptake^1H post XXX challenge|Thyroxine uptake^1H post XXX challenge
C0550143|T201|COMP|12931-2|LNC|Thyroxine^1H post XXX challenge|Thyroxine^1H post XXX challenge
C0550144|T201|COMP|12923-9|LNC|Thyroxine^2nd specimen post XXX challenge|Thyroxine^2nd specimen post XXX challenge
C0550145|T201|COMP|12924-7|LNC|Thyroxine^3rd specimen post XXX challenge|Thyroxine^3rd specimen post XXX challenge
C0550146|T201|COMP|12925-4|LNC|Thyroxine^4th specimen post XXX challenge|Thyroxine^4th specimen post XXX challenge
C0550147|T201|COMP|12926-2|LNC|Thyroxine^5th specimen post XXX challenge|Thyroxine^5th specimen post XXX challenge
C0550148|T201|COMP|12927-0|LNC|Thyroxine^6th specimen post XXX challenge|Thyroxine^6th specimen post XXX challenge
C0550149|T201|COMP|12928-8|LNC|Thyroxine^7th specimen post XXX challenge|Thyroxine^7th specimen post XXX challenge
C0550150|T201|COMP|12929-6|LNC|Thyroxine^8th specimen post XXX challenge|Thyroxine^8th specimen post XXX challenge
C0550151|T201|COMP|12930-4|LNC|Thyroxine^9th specimen post XXX challenge|Thyroxine^9th specimen post XXX challenge
C0550152|T201|COMP|12982-5|LNC|Vasopressin^2nd specimen post XXX challenge|Vasopressin^2nd specimen post XXX challenge
C0550153|T201|COMP|13028-6|LNC|Xylose^1.5H post XXX challenge|Xylose^1.5H post XXX challenge
C0550154|T201|COMP|10869-6|LNC|Xylose^3H post 25 g xylose PO|Xylose^3H post 25 g xylose PO
C0550155|T201|COMP|13029-4|LNC|Xylose^3H post XXX challenge|Xylose^3H post XXX challenge
C0550156|T201|COMP|10870-4|LNC|Xylose^4H post 25 g xylose PO|Xylose^4H post 25 g xylose PO
C0550157|T201|COMP|13030-2|LNC|Xylose^4H post XXX challenge|Xylose^4H post XXX challenge
C0550158|T201|COMP|10871-2|LNC|Xylose^5H post 25 g xylose PO|Xylose^5H post 25 g xylose PO
C0550159|T201|COMP|13031-0|LNC|Xylose^5H post XXX challenge|Xylose^5H post XXX challenge
C0550160|T201|COMP|10872-0|LNC|Xylose^baseline|Xylose^baseline
C0550161|T201|COMP|12997-3|LNC|1,4-Dioxane|1,4-Dioxane
C0550162|T201|COMP|13406-4|LNC|1-Methylhistidine|1-Methylhistidine
C0550163|T201|COMP|13377-7|LNC|1-Methylhistidine|1-Methylhistidine
C0550164|T201|COMP|12769-6|LNC|17-Ketosteroids.total neutral|17-Ketosteroids.total neutral
C0550165|T201|COMP|11206-0|LNC|18-Hydroxydeoxycorticosterone|18-Hydroxydeoxycorticosterone
C0550166|T201|COMP|13480-9|LNC|18-Hydroxydeoxycortisol/Creatinine|18-Hydroxydeoxycortisol/Creatinine
C0550167|T201|COMP|12986-6|LNC|2,5-Hexanedione|2,5-Hexanedione
C0550168|T201|COMP|12540-1|LNC|2-Methylcitrate|2-Methylcitrate
C0550169|T201|COMP|12539-3|LNC|2-Methylcitrate|2-Methylcitrate
C0550170|T201|COMP|12533-6|LNC|Thiazolidine-2-Thione-4-Carboxylic acid|Thiazolidine-2-Thione-4-Carboxylic acid
C0550172|T201|COMP|12541-9|LNC|Meta methylhippurate+Para methylhippurate|Meta methylhippurate+Para methylhippurate
C0550173|T201|COMP|13407-2|LNC|3-Methylhistidine|3-Methylhistidine
C0550174|T201|COMP|13378-5|LNC|3-Methylhistidine|3-Methylhistidine
C0550175|T201|COMP|12172-3|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C0550176|T201|COMP|11145-0|LNC|5-Hydroxyindoleacetate/Creatinine|5-Hydroxyindoleacetate/Creatinine
C0550177|T201|COMP|12987-4|LNC|Acetonitrile|Acetonitrile
C0550178|T201|COMP|11034-6|LNC|Acetylcholine receptor binding Ab|Acetylcholine receptor binding Ab
C0550179|T201|COMP|12899-1|LNC|Acetylene|Acetylene
C0550180|T201|COMP|12804-1|LNC|Acid phosphatase|Acid phosphatase
C0550181|T201|COMP|12173-1|LNC|Acid phosphatase.non-prostatic|Acid phosphatase.non-prostatic
C0550182|T201|COMP|12988-2|LNC|Acrylamide|Acrylamide
C0550183|T201|COMP|11035-3|LNC|Adenylate kinase|Adenylate kinase
C0550184|T201|COMP|12280-4|LNC|Alanine|Alanine
C0550185|T201|COMP|12174-9|LNC|Albumin/Globulin|Albumin/Globulin
C0550186|T201|COMP|12175-6|LNC|Albumin/Globulin|Albumin/Globulin
C0550187|T201|COMP|2299-6|LNC|Aldolase|Aldolase
C0550188|T201|COMP|13482-5|LNC|Aldosterone/Creatinine|Aldosterone/Creatinine
C0550189|T201|COMP|12805-8|LNC|Alkaline phosphatase isoenzyme|Alkaline phosphatase isoenzyme
C0550190|T201|COMP|12806-6|LNC|Alkaline phosphatase.lung|Alkaline phosphatase.lung
C0550191|T201|COMP|13383-5|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0550192|T201|COMP|13384-3|LNC|Alpha aminoadipate|Alpha aminoadipate
C0550193|T201|COMP|13366-0|LNC|Alpha aminoadipate|Alpha aminoadipate
C0550194|T201|COMP|11037-9|LNC|Alpha-N-acetylgalactosaminidase|Alpha-N-acetylgalactosaminidase
C0550195|T201|COMP|12728-2|LNC|Alpha subunit|Alpha subunit
C0550196|T201|COMP|12960-1|LNC|Alpha 1 antitrypsin fecal clearance|Alpha 1 antitrypsin fecal clearance
C0550197|T201|COMP|12466-9|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C0550198|T201|COMP|11207-8|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0550199|T201|COMP|13500-4|LNC|Amino acid pattern|Amino acid pattern
C0550200|T201|COMP|12176-4|LNC|Amino acids|Amino acids
C0550201|T201|COMP|12468-5|LNC|Amino acids|Amino acids
C0550202|T201|COMP|12467-7|LNC|Amino acids|Amino acids
C0550203|T201|COMP|12177-2|LNC|Amino acids/Creatinine|Amino acids/Creatinine
C0550204|T201|COMP|12472-7|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0550209|T201|COMP|12479-2|LNC|Androsterone|Androsterone
C0550210|T201|COMP|12480-0|LNC|Angiotensin converting enzyme|Angiotensin converting enzyme
C0550211|T201|COMP|13386-8|LNC|Anserine|Anserine
C0550212|T201|COMP|13462-7|LNC|Apolipoprotein A-I/Apolipoprotein B|Apolipoprotein A-I/Apolipoprotein B
C0550213|T201|COMP|11135-1|LNC|Appearance|Appearance
C0550214|T201|COMP|11134-4|LNC|Appearance|Appearance
C0550215|T201|COMP|11158-3|LNC|Appearance|Appearance
C0550216|T201|COMP|13387-6|LNC|Arginine|Arginine
C0550217|T201|COMP|12482-6|LNC|Ascorbate|Ascorbate
C0550218|T201|COMP|13388-4|LNC|Asparagine|Asparagine
C0550219|T201|COMP|13389-2|LNC|Aspartate|Aspartate
C0550220|T201|COMP|11208-6|LNC|Atrial natriuretic factor|Atrial natriuretic factor
C0550221|T201|COMP|11555-0|LNC|Base excess|Base excess
C0550222|T201|COMP|13390-0|LNC|Beta alanine|Beta alanine
C0550223|T201|COMP|13368-6|LNC|Beta alanine|Beta alanine
C0550224|T201|COMP|13385-0|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0550225|T201|COMP|13367-8|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0550226|T201|COMP|12915-5|LNC|Beta galactosidase|Beta galactosidase
C0550227|T201|COMP|11038-7|LNC|Beta+gamma tocopherol|Beta+gamma tocopherol
C0550228|T201|COMP|11209-4|LNC|Beta glucuronidase|Beta glucuronidase
C0550229|T201|COMP|10873-8|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C0550230|T201|COMP|13485-8|LNC|Beta-2-Microglobulin/Creatinine|Beta-2-Microglobulin/Creatinine
C0550231|T201|COMP|12913-0|LNC|Beta-N-acetylhexosaminidase|Beta-N-acetylhexosaminidase
C0550232|T201|COMP|12514-6|LNC|Bicarbonate|Bicarbonate
C0550233|T201|COMP|12513-8|LNC|Bicarbonate|Bicarbonate
C0550235|T201|COMP|12476-8|LNC|Bilirubin|Bilirubin
C0550236|T201|COMP|10874-6|LNC|Bombesin|Bombesin
C0550237|T201|COMP|11039-5|LNC|C reactive protein|C reactive protein
C0550238|T201|COMP|13454-4|LNC|Calcium-phosphorus product|Calcium-phosphorus product
C0550239|T201|COMP|12180-6|LNC|Calcium.ionized|Calcium.ionized
C0550240|T201|COMP|12181-4|LNC|Calcium|Calcium
C0550241|T201|COMP|12511-2|LNC|Calcium|Calcium
C0550242|T201|COMP|13444-5|LNC|Calcium/Albumin|Calcium/Albumin
C0550243|T201|COMP|13448-6|LNC|Calcium/Osmolality|Calcium/Osmolality
C0550244|T201|COMP|11210-2|LNC|Cancer Ag 125|Cancer Ag 125
C0550245|T201|COMP|13127-6|LNC|Cancer Ag DM-70K|Cancer Ag DM-70K
C0550246|T201|COMP|11557-6|LNC|Carbon dioxide|Carbon dioxide
C0550247|T201|COMP|11211-0|LNC|Carbon dioxide|Carbon dioxide
C0550248|T201|COMP|12515-3|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0550249|T201|COMP|10876-1|LNC|Carnitine esters|Carnitine esters
C0550250|T201|COMP|10875-3|LNC|Carnitine esters|Carnitine esters
C0550251|T201|COMP|10877-9|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C0550252|T201|COMP|13391-8|LNC|Carnosine|Carnosine
C0550253|T201|COMP|13369-4|LNC|Carnosine|Carnosine
C0550254|T201|COMP|12474-3|LNC|Carnosine|Carnosine
C0550255|T201|COMP|11133-6|LNC|Catecholamines.free|Catecholamines.free
C0550256|T201|COMP|12898-3|LNC|Chloride|Chloride
C0550257|T201|COMP|12530-2|LNC|Chloride|Chloride
C0550258|T201|COMP|11054-4|LNC|Cholesterol.in LDL/Cholesterol.in HDL|Cholesterol.in LDL/Cholesterol.in HDL
C0550259|T201|COMP|12772-0|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C0550260|T201|COMP|12771-2|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C0550261|T201|COMP|12773-8|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C0550262|T201|COMP|13459-3|LNC|Cholesterol.in LDL/Cholesterol.total|Cholesterol.in LDL/Cholesterol.total
C0550264|T201|COMP|13457-7|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C0550265|T201|COMP|13458-5|LNC|Cholesterol.in VLDL|Cholesterol.in VLDL
C0550266|T201|COMP|12183-0|LNC|Cholesterol|Cholesterol
C0550267|T201|COMP|11154-2|LNC|Cholinesterase|Cholinesterase
C0550268|T201|COMP|12184-8|LNC|Choriogonadotropin|Choriogonadotropin
C0550269|T201|COMP|13392-6|LNC|Citrulline|Citrulline
C0550270|T201|COMP|12186-3|LNC|Colloid oncotic pressure|Colloid oncotic pressure
C0550271|T201|COMP|11212-8|LNC|Coproporphyrin|Coproporphyrin
C0550272|T201|COMP|12809-0|LNC|Coproporphyrin|Coproporphyrin
C0550273|T201|COMP|11213-6|LNC|Corticotropin releasing hormone|Corticotropin releasing hormone
C0550274|T201|COMP|12283-8|LNC|Corticotropin releasing hormone|Corticotropin releasing hormone
C0550275|T201|COMP|11040-3|LNC|Cortisol.free|Cortisol.free
C0550276|T201|COMP|11155-9|LNC|Cortisol/Creatinine|Cortisol/Creatinine
C0550277|T201|COMP|12189-7|LNC|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C0550278|T201|COMP|12188-9|LNC|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C0550279|T201|COMP|12187-1|LNC|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C0550280|T201|COMP|13484-1|LNC|Creatine/Creatinine|Creatine/Creatinine
C0550281|T201|COMP|12190-5|LNC|Creatinine|Creatinine
C0550282|T201|COMP|12192-1|LNC|Creatinine^2H post peritoneal dialysis|Creatinine^2H post peritoneal dialysis
C0550283|T201|COMP|12193-9|LNC|Creatinine^4H post peritoneal dialysis|Creatinine^4H post peritoneal dialysis
C0550284|T201|COMP|12191-3|LNC|Creatinine|Creatinine
C0550285|T201|COMP|12589-8|LNC|Creatinine|Creatinine
C0550286|T201|COMP|12585-6|LNC|Creatinine|Creatinine
C0550287|T201|COMP|12586-4|LNC|Creatinine|Creatinine
C0550288|T201|COMP|12587-2|LNC|Creatinine|Creatinine
C0550289|T201|COMP|12588-0|LNC|Creatinine|Creatinine
C0550290|T201|COMP|11214-4|LNC|Creatinine|Creatinine
C0550291|T201|COMP|12584-9|LNC|Creatinine|Creatinine
C0550292|T201|COMP|13451-0|LNC|Creatinine dialysis fluid clearance|Creatinine dialysis fluid clearance
C0550293|T201|COMP|13441-1|LNC|Creatinine renal clearance|Creatinine renal clearance
C0550294|T201|COMP|13442-9|LNC|Creatinine renal clearance|Creatinine renal clearance
C0550295|T201|COMP|13443-7|LNC|Creatinine renal clearance|Creatinine renal clearance
C0550296|T201|COMP|12194-7|LNC|Creatinine^12H post peritoneal dialysis|Creatinine^12H post peritoneal dialysis
C0550297|T201|COMP|12576-5|LNC|Creatinine^1st specimen|Creatinine^1st specimen
C0550298|T201|COMP|12574-0|LNC|Creatinine^24H specimen|Creatinine^24H specimen
C0550299|T201|COMP|12572-4|LNC|Creatinine^2H dwell specimen|Creatinine^2H dwell specimen
C0550300|T201|COMP|12577-3|LNC|Creatinine^2nd specimen|Creatinine^2nd specimen
C0550301|T201|COMP|12578-1|LNC|Creatinine^3rd specimen|Creatinine^3rd specimen
C0550302|T201|COMP|12573-2|LNC|Creatinine^4H dwell specimen|Creatinine^4H dwell specimen
C0550303|T201|COMP|12579-9|LNC|Creatinine^4th specimen|Creatinine^4th specimen
C0550304|T201|COMP|12580-7|LNC|Creatinine^5th specimen|Creatinine^5th specimen
C0550305|T201|COMP|12581-5|LNC|Creatinine^6th specimen|Creatinine^6th specimen
C0550306|T201|COMP|12582-3|LNC|Creatinine^7th specimen|Creatinine^7th specimen
C0550307|T201|COMP|12583-1|LNC|Creatinine^8th specimen|Creatinine^8th specimen
C0550308|T201|COMP|12575-7|LNC|Creatinine^baseline|Creatinine^baseline
C0550309|T201|COMP|11041-1|LNC|Creatinine^post dialysis|Creatinine^post dialysis
C0550310|T201|COMP|11042-9|LNC|Creatinine^pre dialysis|Creatinine^pre dialysis
C0550311|T201|COMP|11043-7|LNC|Cryofibrinogen|Cryofibrinogen
C0550312|T201|COMP|12197-0|LNC|Cryofibrinogen|Cryofibrinogen
C0550313|T201|COMP|12198-8|LNC|Cryofibrinogen|Cryofibrinogen
C0550314|T201|COMP|12199-6|LNC|Cryofibrinogen|Cryofibrinogen
C0550315|T201|COMP|12196-2|LNC|Cryofibrinogen|Cryofibrinogen
C0550316|T201|COMP|12207-7|LNC|Cryoglobulin|Cryoglobulin
C0550317|T201|COMP|12201-0|LNC|Cryoglobulin|Cryoglobulin
C0550318|T201|COMP|12202-8|LNC|Cryoglobulin|Cryoglobulin
C0550319|T201|COMP|12203-6|LNC|Cryoglobulin|Cryoglobulin
C0550320|T201|COMP|12204-4|LNC|Cryoglobulin|Cryoglobulin
C0550321|T201|COMP|12200-2|LNC|Cryoglobulin|Cryoglobulin
C0550322|T201|COMP|12205-1|LNC|Cryoglobulin|Cryoglobulin
C0550323|T201|COMP|12206-9|LNC|Cryoglobulin|Cryoglobulin
C0550324|T201|COMP|13393-4|LNC|Cystathionine|Cystathionine
C0550325|T201|COMP|13370-2|LNC|Cystathionine|Cystathionine
C0550326|T201|COMP|13394-2|LNC|Cystine|Cystine
C0550327|T201|COMP|13371-0|LNC|Cystine|Cystine
C0550328|T201|COMP|10969-4|LNC|Cystine+Homocysteine|Cystine+Homocysteine
C0550334|T201|COMP|11215-1|LNC|Delta aminolevulinate|Delta aminolevulinate
C0550335|T201|COMP|12475-0|LNC|Delta aminolevulinate|Delta aminolevulinate
C0550336|T201|COMP|11216-9|LNC|Deoxypyridinoline|Deoxypyridinoline
C0550337|T201|COMP|11044-5|LNC|Diphosphoglycerate mutase|Diphosphoglycerate mutase
C0550338|T201|COMP|11045-2|LNC|Enolase|Enolase
C0550339|T201|COMP|11046-0|LNC|EPINEPHrine|EPINEPHrine
C0550340|T201|COMP|12214-3|LNC|Estradiol|Estradiol
C0550341|T201|COMP|12213-5|LNC|Estradiol|Estradiol
C0550342|T201|COMP|12595-5|LNC|Estradiol|Estradiol
C0550344|T201|COMP|12598-9|LNC|Fat.neutral|Fat.neutral
C0550345|T201|COMP|12215-0|LNC|Fatty acids.very long chain|Fatty acids.very long chain
C0550346|T201|COMP|13489-0|LNC|Follitropin/Creatinine|Follitropin/Creatinine
C0550347|T201|COMP|10970-2|LNC|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C0550348|T201|COMP|12217-6|LNC|Globulin|Globulin
C0550349|T201|COMP|10834-0|LNC|Globulin|Globulin
C0550350|T201|COMP|12629-2|LNC|Glucose|Glucose
C0550351|T201|COMP|12628-4|LNC|Glucose|Glucose
C0550352|T201|COMP|12220-0|LNC|Glucose^12H post peritoneal dialysis|Glucose^12H post peritoneal dialysis
C0550353|T201|COMP|12218-4|LNC|Glucose^2H post peritoneal dialysis|Glucose^2H post peritoneal dialysis
C0550354|T201|COMP|12219-2|LNC|Glucose^4H post peritoneal dialysis|Glucose^4H post peritoneal dialysis
C0550355|T201|COMP|13453-6|LNC|Glucose mean value|Glucose mean value
C0550356|T201|COMP|11047-8|LNC|Glucose phosphate isomerase|Glucose phosphate isomerase
C0550357|T201|COMP|11142-7|LNC|Glucose^15M post 100 g glucose PO|Glucose^15M post 100 g glucose PO
C0550358|T201|COMP|12630-0|LNC|Glucose^1st specimen|Glucose^1st specimen
C0550359|T201|COMP|12612-8|LNC|Glucose^2H specimen|Glucose^2H specimen
C0550360|T201|COMP|12608-6|LNC|Glucose^2H dwell specimen|Glucose^2H dwell specimen
C0550361|T201|COMP|12631-8|LNC|Glucose^2nd specimen|Glucose^2nd specimen
C0550362|T201|COMP|12632-6|LNC|Glucose^3rd specimen|Glucose^3rd specimen
C0550363|T201|COMP|11143-5|LNC|Glucose^45M post 100 g glucose PO|Glucose^45M post 100 g glucose PO
C0550364|T201|COMP|12613-6|LNC|Glucose^4H specimen|Glucose^4H specimen
C0550365|T201|COMP|12609-4|LNC|Glucose^4H dwell specimen|Glucose^4H dwell specimen
C0550366|T201|COMP|12611-0|LNC|Glucose^4H specimen|Glucose^4H specimen
C0550367|T201|COMP|12633-4|LNC|Glucose^4th specimen|Glucose^4th specimen
C0550368|T201|COMP|12634-2|LNC|Glucose^5th specimen|Glucose^5th specimen
C0550369|T201|COMP|12635-9|LNC|Glucose^6th specimen|Glucose^6th specimen
C0550370|T201|COMP|12636-7|LNC|Glucose^7th specimen|Glucose^7th specimen
C0550371|T201|COMP|12607-8|LNC|Glucose^pre dialysis|Glucose^pre dialysis
C0550372|T201|COMP|13395-9|LNC|Glutamate|Glutamate
C0550373|T201|COMP|13396-7|LNC|Glutamine|Glutamine
C0550374|T201|COMP|11048-6|LNC|Glyceraldehyde 3 phosphate dehydrogenase|Glyceraldehyde 3 phosphate dehydrogenase
C0550375|T201|COMP|13397-5|LNC|Glycine|Glycine
C0550376|T201|COMP|13481-7|LNC|Gonadotropin peptide/Creatinine|Gonadotropin peptide/Creatinine
C0550377|T201|COMP|12503-9|LNC|Hemoglobin.gastrointestinal^4th specimen|Hemoglobin.gastrointestinal^4th specimen
C0550378|T201|COMP|12504-7|LNC|Hemoglobin.gastrointestinal^5th specimen|Hemoglobin.gastrointestinal^5th specimen
C0550379|T201|COMP|11217-7|LNC|Hexaporphyrin|Hexaporphyrin
C0550380|T201|COMP|13398-3|LNC|Histidine|Histidine
C0550381|T201|COMP|12470-1|LNC|Homocysteine|Homocysteine
C0550382|T201|COMP|13399-1|LNC|Homocystine|Homocystine
C0550383|T201|COMP|13372-8|LNC|Homocystine|Homocystine
C0550384|T201|COMP|11144-3|LNC|Homovanillate|Homovanillate
C0550385|T201|COMP|12715-9|LNC|Homovanillate|Homovanillate
C0550386|T201|COMP|11146-8|LNC|Homovanillate/Creatinine|Homovanillate/Creatinine
C0550387|T201|COMP|13400-7|LNC|Hydroxylysine|Hydroxylysine
C0550388|T201|COMP|13373-6|LNC|Hydroxylysine|Hydroxylysine
C0550389|T201|COMP|13401-5|LNC|Hydroxyproline|Hydroxyproline
C0550390|T201|COMP|13374-4|LNC|Hydroxyproline|Hydroxyproline
C0550392|T201|COMP|12720-9|LNC|Hydroxyproline|Hydroxyproline
C0550393|T201|COMP|13312-4|LNC|IgA Ab.IgG|IgA Ab.IgG
C0550394|T201|COMP|12725-8|LNC|IgA.secretory|IgA.secretory
C0550395|T201|COMP|13456-9|LNC|IgG synthesis rate|IgG synthesis rate
C0550396|T201|COMP|13313-2|LNC|IgM Ab.IgM|IgM Ab.IgM
C0550397|T201|COMP|11219-3|LNC|Immunoglobulin light chains|Immunoglobulin light chains
C0550398|T201|COMP|11050-2|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C0550399|T201|COMP|11051-0|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C0550400|T201|COMP|12722-5|LNC|Insulin-like growth factor binding protein 1|Insulin-like growth factor binding protein 1
C0550401|T201|COMP|12723-3|LNC|Insulin-like growth factor binding protein 2|Insulin-like growth factor binding protein 2
C0550402|T201|COMP|11220-1|LNC|Iodine.free|Iodine.free
C0550403|T201|COMP|13452-8|LNC|Iron/Transferrin|Iron/Transferrin
C0550404|T201|COMP|13402-3|LNC|Isoleucine|Isoleucine
C0550405|T201|COMP|10879-5|LNC|Isovalerylglycine|Isovalerylglycine
C0550406|T201|COMP|12777-9|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C0550407|T201|COMP|11053-6|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0550408|T201|COMP|12778-7|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C0550409|T201|COMP|13403-1|LNC|Leucine|Leucine
C0550410|T201|COMP|12726-6|LNC|Leucine-enkephalin|Leucine-enkephalin
C0550411|T201|COMP|12912-2|LNC|Lipids|Lipids
C0550413|T201|COMP|10835-7|LNC|Lipoprotein (little a)|Lipoprotein (little a)
C0550414|T201|COMP|13490-8|LNC|Lutropin/Creatinine|Lutropin/Creatinine
C0550415|T201|COMP|13404-9|LNC|Lysine|Lysine
C0550416|T201|COMP|13375-1|LNC|Lysine|Lysine
C0550417|T201|COMP|10971-0|LNC|Lysozyme|Lysozyme
C0550419|T201|COMP|10880-3|LNC|Magnesium|Magnesium
C0550420|T201|COMP|13474-2|LNC|Magnesium/Creatinine|Magnesium/Creatinine
C0550421|T201|COMP|12231-7|LNC|Prolactin^baseline|Prolactin^baseline
C0550422|T201|COMP|13000-5|LNC|Mandelate|Mandelate
C0550423|T201|COMP|13001-3|LNC|Mandelate/Creatinine|Mandelate/Creatinine
C0550424|T201|COMP|11055-1|LNC|Melatonin|Melatonin
C0550425|T201|COMP|12721-7|LNC|Melatonin|Melatonin
C0550426|T201|COMP|11056-9|LNC|Melatonin|Melatonin
C0550427|T201|COMP|11140-1|LNC|Metanephrine|Metanephrine
C0550428|T201|COMP|13405-6|LNC|Methionine|Methionine
C0550429|T201|COMP|13376-9|LNC|Methionine|Methionine
C0550430|T201|COMP|11057-7|LNC|Monophosphoglyceromutase|Monophosphoglyceromutase
C0550431|T201|COMP|11147-6|LNC|Myoglobin/Creatinine|Myoglobin/Creatinine
C0550432|T201|COMP|10836-5|LNC|Niacin|Niacin
C0550433|T201|COMP|12239-0|LNC|Oligosaccharides|Oligosaccharides
C0550434|T201|COMP|10837-3|LNC|Organic acids|Organic acids
C0550435|T201|COMP|10972-8|LNC|Organic acids|Organic acids
C0550436|T201|COMP|13408-0|LNC|Ornithine|Ornithine
C0550437|T201|COMP|13379-3|LNC|Ornithine|Ornithine
C0550438|T201|COMP|12240-8|LNC|Orotidine|Orotidine
C0550439|T201|COMP|13483-3|LNC|Oxalate/Creatinine|Oxalate/Creatinine
C0550440|T201|COMP|11556-8|LNC|Oxygen|Oxygen
C0550441|T201|COMP|11559-2|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C0550442|T201|COMP|12334-9|LNC|Para aminophenol|Para aminophenol
C0550443|T201|COMP|10882-9|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C0550444|T201|COMP|10881-1|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C0550445|T201|COMP|11221-9|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C0550446|T201|COMP|11222-7|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C0550448|T201|COMP|13487-4|LNC|Phenol/Creatinine|Phenol/Creatinine
C0550449|T201|COMP|10883-7|LNC|Phenolphthalein|Phenolphthalein
C0550450|T201|COMP|12317-4|LNC|Phenolphthalein|Phenolphthalein
C0550451|T201|COMP|11223-5|LNC|Phenolphthalein|Phenolphthalein
C0550452|T201|COMP|13409-8|LNC|Phenylalanine|Phenylalanine
C0550453|T201|COMP|12803-3|LNC|Phenylalanine|Phenylalanine
C0550454|T201|COMP|12537-7|LNC|Phenylglyoxylate|Phenylglyoxylate
C0550455|T201|COMP|12242-4|LNC|Phosphate|Phosphate
C0550456|T201|COMP|10884-5|LNC|Phosphate|Phosphate
C0550457|T201|COMP|11141-9|LNC|Phosphate/Creatinine|Phosphate/Creatinine
C0550458|T201|COMP|13410-6|LNC|Phosphoethanolamine|Phosphoethanolamine
C0550459|T201|COMP|11224-3|LNC|Phosphoethanolamine|Phosphoethanolamine
C0550460|T201|COMP|12473-5|LNC|Phosphoethanolamine|Phosphoethanolamine
C0550461|T201|COMP|11058-5|LNC|Phosphofructokinase|Phosphofructokinase
C0550462|T201|COMP|11059-3|LNC|Phosphoglycerate kinase|Phosphoglycerate kinase
C0550463|T201|COMP|13411-4|LNC|Phosphoserine|Phosphoserine
C0550464|T201|COMP|12807-4|LNC|Phosphoserine|Phosphoserine
C0550465|T201|COMP|10838-1|LNC|Phosphoserine|Phosphoserine
C0550466|T201|COMP|12245-7|LNC|Porphobilinogen|Porphobilinogen
C0550467|T201|COMP|12916-3|LNC|Porphobilinogen synthase|Porphobilinogen synthase
C0550468|T201|COMP|12917-1|LNC|Porphobilinogen synthase|Porphobilinogen synthase
C0550469|T201|COMP|11225-0|LNC|Porphyrins|Porphyrins
C0550470|T201|COMP|12246-5|LNC|Porphyrins|Porphyrins
C0550471|T201|COMP|10885-2|LNC|Porphyrins|Porphyrins
C0550472|T201|COMP|12814-0|LNC|Potassium|Potassium
C0550473|T201|COMP|11148-4|LNC|Potassium/Creatinine|Potassium/Creatinine
C0550474|T201|COMP|12812-4|LNC|Potassium^2nd specimen|Potassium^2nd specimen
C0550475|T201|COMP|12813-2|LNC|Potassium^3rd specimen|Potassium^3rd specimen
C0550476|T201|COMP|12599-7|LNC|Pristanate|Pristanate
C0550477|T201|COMP|12600-3|LNC|Pristanate/Phytanate|Pristanate/Phytanate
C0550478|T201|COMP|12820-7|LNC|Progesterone|Progesterone
C0550479|T201|COMP|13412-2|LNC|Proline|Proline
C0550480|T201|COMP|11226-8|LNC|Prorenin|Prorenin
C0550481|T201|COMP|12839-7|LNC|Prostaglandin D2|Prostaglandin D2
C0550482|T201|COMP|12838-9|LNC|Prostaglandin D2|Prostaglandin D2
C0550483|T201|COMP|12837-1|LNC|Prostaglandin E1|Prostaglandin E1
C0550484|T201|COMP|12836-3|LNC|Prostaglandin E2|Prostaglandin E2
C0550485|T201|COMP|12840-5|LNC|Prostaglandin F2 alpha|Prostaglandin F2 alpha
C0550486|T201|COMP|10886-0|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C0550488|T201|COMP|13439-5|LNC|Protein pattern|Protein pattern
C0550489|T201|COMP|12851-2|LNC|Protein pattern|Protein pattern
C0550490|T201|COMP|13438-7|LNC|Protein pattern|Protein pattern
C0550491|T201|COMP|12782-9|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C0550492|T201|COMP|12783-7|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C0550493|T201|COMP|13128-4|LNC|Immunosuppressive acidic protein|Immunosuppressive acidic protein
C0550494|T201|COMP|12843-9|LNC|Protein|Protein
C0550495|T201|COMP|12842-1|LNC|Protein|Protein
C0550496|T201|COMP|12844-7|LNC|Protein^2nd specimen|Protein^2nd specimen
C0550497|T201|COMP|12845-4|LNC|Protein^3rd specimen|Protein^3rd specimen
C0550498|T201|COMP|12846-2|LNC|Protein^4th specimen|Protein^4th specimen
C0550499|T201|COMP|12847-0|LNC|Protein^5th specimen|Protein^5th specimen
C0550500|T201|COMP|12848-8|LNC|Protein^6th specimen|Protein^6th specimen
C0550501|T201|COMP|12849-6|LNC|Protein^7th specimen|Protein^7th specimen
C0550502|T201|COMP|12850-4|LNC|Protein^8th specimen|Protein^8th specimen
C0550503|T201|COMP|10887-8|LNC|Pyridinoline|Pyridinoline
C0550504|T201|COMP|12247-3|LNC|Pyruvate|Pyruvate
C0550505|T201|COMP|11227-6|LNC|Pyruvate kinase|Pyruvate kinase
C0550506|T201|COMP|11060-1|LNC|Reducing substances|Reducing substances
C0550507|T201|COMP|12249-9|LNC|Renin|Renin
C0550508|T201|COMP|13413-0|LNC|Sarcosine|Sarcosine
C0550509|T201|COMP|13380-1|LNC|Sarcosine|Sarcosine
C0550510|T201|COMP|13414-8|LNC|Serine|Serine
C0550511|T201|COMP|12907-2|LNC|Sodium|Sodium
C0550512|T201|COMP|12908-0|LNC|Sodium|Sodium
C0550513|T201|COMP|11149-2|LNC|Sodium/Creatinine|Sodium/Creatinine
C0550514|T201|COMP|12252-3|LNC|Somatomedin C|Somatomedin C
C0550515|T201|COMP|12284-6|LNC|Growth hormone-releasing hormone|Growth hormone-releasing hormone
C0550516|T201|COMP|12253-1|LNC|Somatotropin^baseline|Somatotropin^baseline
C0550517|T201|COMP|12260-6|LNC|Sucrose hemolysis|Sucrose hemolysis
C0550518|T201|COMP|12920-5|LNC|Sulfate|Sulfate
C0550519|T201|COMP|13123-5|LNC|Sulfate-3-Glucuronyl paragloboside Ab|Sulfate-3-Glucuronyl paragloboside Ab
C0550520|T201|COMP|13101-1|LNC|Sulfate-3-Glucuronyl paragloboside Ab.IgM|Sulfate-3-Glucuronyl paragloboside Ab.IgM
C0550521|T201|COMP|13100-3|LNC|Sulfate-3-Glucuronyl paragloboside Ab.IgM|Sulfate-3-Glucuronyl paragloboside Ab.IgM
C0550522|T201|COMP|13415-5|LNC|Taurine|Taurine
C0550523|T201|COMP|13486-6|LNC|Testosterone/Creatinine|Testosterone/Creatinine
C0550524|T201|COMP|12420-6|LNC|Thiosulfate|Thiosulfate
C0550525|T201|COMP|12421-4|LNC|Thiosulfate/Creatinine|Thiosulfate/Creatinine
C0550526|T201|COMP|13416-3|LNC|Threonine|Threonine
C0550527|T201|COMP|11061-9|LNC|11-Dehydro thromboxane beta 2|11-Dehydro thromboxane beta 2
C0550528|T201|COMP|11580-8|LNC|Thyrotropin|Thyrotropin
C0550529|T201|COMP|11579-0|LNC|Thyrotropin|Thyrotropin
C0550530|T201|COMP|11062-7|LNC|Thyroxine.albumin bound|Thyroxine.albumin bound
C0550531|T201|COMP|12949-4|LNC|Transferrin.carbohydrate deficient|Transferrin.carbohydrate deficient
C0550532|T201|COMP|10888-6|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C0550533|T201|COMP|12228-3|LNC|Triglyceride|Triglyceride
C0550533|T201|COMP|12950-2|LNC|Triglyceride|Triglyceride
C0550533|T201|COMP|13899-0|LNC|Triglyceride|Triglyceride
C0550534|T201|COMP|12951-0|LNC|Triglyceride|Triglyceride
C0550535|T201|COMP|12953-6|LNC|Triiodothyronine^2nd specimen post XXX challenge|Triiodothyronine^2nd specimen post XXX challenge
C0550536|T201|COMP|12954-4|LNC|Triiodothyronine^3rd specimen post XXX challenge|Triiodothyronine^3rd specimen post XXX challenge
C0550537|T201|COMP|12955-1|LNC|Triiodothyronine^4th specimen post XXX challenge|Triiodothyronine^4th specimen post XXX challenge
C0550538|T201|COMP|12956-9|LNC|Triiodothyronine^5th specimen post XXX challenge|Triiodothyronine^5th specimen post XXX challenge
C0550539|T201|COMP|12957-7|LNC|Triiodothyronine^6th specimen post XXX challenge|Triiodothyronine^6th specimen post XXX challenge
C0550540|T201|COMP|12958-5|LNC|Triiodothyronine^7th specimen post XXX challenge|Triiodothyronine^7th specimen post XXX challenge
C0550541|T201|COMP|12959-3|LNC|Triiodothyronine^8th specimen post XXX challenge|Triiodothyronine^8th specimen post XXX challenge
C0550542|T201|COMP|11063-5|LNC|Triosephosphate isomerase|Triosephosphate isomerase
C0550543|T201|COMP|10839-9|LNC|Troponin I.cardiac|Troponin I.cardiac
C0550544|T201|COMP|12733-2|LNC|Tryptase|Tryptase
C0550545|T201|COMP|13418-9|LNC|Tryptophan|Tryptophan
C0550546|T201|COMP|13417-1|LNC|Tyrosine|Tyrosine
C0550547|T201|COMP|13381-9|LNC|Tyrosine|Tyrosine
C0550548|T201|COMP|12264-8|LNC|Epstein Barr virus early restricted Ab|Epstein Barr virus early restricted Ab
C0550549|T201|COMP|12961-9|LNC|Urea nitrogen|Urea nitrogen
C0550550|T201|COMP|12963-5|LNC|Urea nitrogen|Urea nitrogen
C0550551|T201|COMP|12962-7|LNC|Urea nitrogen|Urea nitrogen
C0550552|T201|COMP|12268-9|LNC|Urea nitrogen^12H post peritoneal dialysis|Urea nitrogen^12H post peritoneal dialysis
C0550553|T201|COMP|12266-3|LNC|Urea nitrogen^2H post peritoneal dialysis|Urea nitrogen^2H post peritoneal dialysis
C0550554|T201|COMP|12267-1|LNC|Urea nitrogen^4H post peritoneal dialysis|Urea nitrogen^4H post peritoneal dialysis
C0550555|T201|COMP|12265-5|LNC|Urea nitrogen|Urea nitrogen
C0550556|T201|COMP|13506-1|LNC|Urea nitrogen renal clearance|Urea nitrogen renal clearance
C0550557|T201|COMP|12981-7|LNC|Urea nitrogen^post dialysis/pre dialysis|Urea nitrogen^post dialysis/pre dialysis
C0550558|T201|COMP|12967-6|LNC|Urea nitrogen|Urea nitrogen
C0550559|T201|COMP|12972-6|LNC|Urea nitrogen^1st specimen|Urea nitrogen^1st specimen
C0550560|T201|COMP|12979-1|LNC|Urea nitrogen^24H specimen|Urea nitrogen^24H specimen
C0550561|T201|COMP|12970-0|LNC|Urea nitrogen^2H dwell specimen|Urea nitrogen^2H dwell specimen
C0550562|T201|COMP|12966-8|LNC|Urea nitrogen^2H specimen|Urea nitrogen^2H specimen
C0550563|T201|COMP|12974-2|LNC|Urea nitrogen^3rd specimen|Urea nitrogen^3rd specimen
C0550564|T201|COMP|12968-4|LNC|Urea nitrogen^4H specimen|Urea nitrogen^4H specimen
C0550565|T201|COMP|12971-8|LNC|Urea nitrogen^4H dwell specimen|Urea nitrogen^4H dwell specimen
C0550566|T201|COMP|12973-4|LNC|Urea nitrogen^4th specimen|Urea nitrogen^4th specimen
C0550567|T201|COMP|12975-9|LNC|Urea nitrogen^5th specimen|Urea nitrogen^5th specimen
C0550568|T201|COMP|12976-7|LNC|Urea nitrogen^6th specimen|Urea nitrogen^6th specimen
C0550569|T201|COMP|12965-0|LNC|Urea nitrogen^70M specimen|Urea nitrogen^70M specimen
C0550570|T201|COMP|12978-3|LNC|Urea nitrogen^7th specimen|Urea nitrogen^7th specimen
C0550571|T201|COMP|12977-5|LNC|Urea nitrogen^8th specimen|Urea nitrogen^8th specimen
C0550572|T201|COMP|12964-3|LNC|Urea nitrogen^baseline|Urea nitrogen^baseline
C0550573|T201|COMP|12969-2|LNC|Urea nitrogen^baseline|Urea nitrogen^baseline
C0550574|T201|COMP|11064-3|LNC|Urea nitrogen^post dialysis|Urea nitrogen^post dialysis
C0550575|T201|COMP|11065-0|LNC|Urea nitrogen^pre dialysis|Urea nitrogen^pre dialysis
C0550576|T201|COMP|12269-7|LNC|Urobilinogen|Urobilinogen
C0550577|T201|COMP|12270-5|LNC|Uroporphyrin|Uroporphyrin
C0550578|T201|COMP|11228-4|LNC|Uroporphyrin|Uroporphyrin
C0550579|T201|COMP|12808-2|LNC|Uroporphyrin|Uroporphyrin
C0550580|T201|COMP|12810-8|LNC|Porphobilinogen deaminase|Porphobilinogen deaminase
C0550581|T201|COMP|12811-6|LNC|Uroporphyrinogen III synthase|Uroporphyrinogen III synthase
C0550582|T201|COMP|11066-8|LNC|Uroporphyrinogen III synthase|Uroporphyrinogen III synthase
C0550583|T201|COMP|13419-7|LNC|Valine|Valine
C0550584|T201|COMP|12274-7|LNC|Xylose|Xylose
C0550585|T201|COMP|11067-6|LNC|Bleeding time|Bleeding time
C0550587|T201|COMP|13488-2|LNC|Coagulation surface induced|Coagulation surface induced
C0550588|T201|COMP|13058-3|LNC|Coagulation surface induced^2nd specimen|Coagulation surface induced^2nd specimen
C0550589|T201|COMP|13059-1|LNC|Coagulation surface induced^3rd specimen|Coagulation surface induced^3rd specimen
C0550590|T201|COMP|13060-9|LNC|Coagulation surface induced^4th specimen|Coagulation surface induced^4th specimen
C0550591|T201|COMP|13053-4|LNC|Coagulation kaolin induced|Coagulation kaolin induced
C0550592|T201|COMP|13054-2|LNC|Fibrin+Fibrinogen fragments|Fibrin+Fibrinogen fragments
C0550593|T201|COMP|13050-0|LNC|Protein C/Coagulation factor IX|Protein C/Coagulation factor IX
C0550594|T201|COMP|13051-8|LNC|Protein S|Protein S
C0550595|T201|COMP|13052-6|LNC|Protein S/Coagulation factor IX|Protein S/Coagulation factor IX
C0550597|T201|COMP|12551-8|LNC|Isocarboxazid|Isocarboxazid
C0550601|T201|COMP|10973-6|LNC|3 methoxy O desmethylencainide|3 methoxy O desmethylencainide
C0550602|T201|COMP|11229-2|LNC|3-O-Methyldopa|3-O-Methyldopa
C0550603|T201|COMP|10974-4|LNC|5-Fluorocytosine|5-Fluorocytosine
C0550604|T201|COMP|10975-1|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0550605|T201|COMP|10976-9|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0550606|T201|COMP|12407-3|LNC|6-Beta naltrexone|6-Beta naltrexone
C0550607|T201|COMP|12788-6|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0550608|T201|COMP|12442-0|LNC|Acetaminophen|Acetaminophen
C0550609|T201|COMP|12502-1|LNC|Allobarbital|Allobarbital
C0550610|T201|COMP|10977-7|LNC|ALPRAZolam|ALPRAZolam
C0550611|T201|COMP|10978-5|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C0550612|T201|COMP|12485-9|LNC|Amobarbital|Amobarbital
C0550613|T201|COMP|12494-1|LNC|Amobarbital|Amobarbital
C0550614|T201|COMP|11230-0|LNC|Amobarbital|Amobarbital
C0550615|T201|COMP|12350-5|LNC|Amphetamines|Amphetamines
C0550616|T201|COMP|12332-3|LNC|Antihistamines|Antihistamines
C0550617|T201|COMP|12344-8|LNC|Antipsychotics|Antipsychotics
C0550618|T201|COMP|12313-3|LNC|Aprobarbital|Aprobarbital
C0550619|T201|COMP|11231-8|LNC|Astemizole|Astemizole
C0550620|T201|COMP|10840-7|LNC|Atropine|Atropine
C0550621|T201|COMP|12495-8|LNC|Barbital|Barbital
C0550622|T201|COMP|12360-4|LNC|Barbital|Barbital
C0550623|T201|COMP|12352-1|LNC|Benzoylecgonine|Benzoylecgonine
C0550624|T201|COMP|13479-1|LNC|Benzoylecgonine/Creatinine|Benzoylecgonine/Creatinine
C0550625|T201|COMP|12328-1|LNC|Beta blockers|Beta blockers
C0550626|T201|COMP|10889-4|LNC|Bisacodyl|Bisacodyl
C0550627|T201|COMP|11232-6|LNC|Bromocriptine|Bromocriptine
C0550628|T201|COMP|11233-4|LNC|Brompheniramine|Brompheniramine
C0550629|T201|COMP|12486-7|LNC|Butabarbital|Butabarbital
C0550630|T201|COMP|12496-6|LNC|Butabarbital|Butabarbital
C0550631|T201|COMP|12487-5|LNC|Butalbital|Butalbital
C0550632|T201|COMP|12497-4|LNC|Butalbital|Butalbital
C0550633|T201|COMP|11071-8|LNC|Butalbital|Butalbital
C0550634|T201|COMP|12394-3|LNC|Butorphanol|Butorphanol
C0550635|T201|COMP|12395-0|LNC|Butorphanol|Butorphanol
C0550636|T201|COMP|12333-1|LNC|Butorphanol|Butorphanol
C0550637|T201|COMP|12363-8|LNC|carBAMazepine|carBAMazepine
C0550638|T201|COMP|10979-3|LNC|Carisoprodol|Carisoprodol
C0550639|T201|COMP|10980-1|LNC|Cephapirin|Cephapirin
C0550640|T201|COMP|12305-9|LNC|Chlordecone|Chlordecone
C0550641|T201|COMP|12427-1|LNC|Chlormezanone|Chlormezanone
C0550642|T201|COMP|12396-8|LNC|chlorproPAMIDE|chlorproPAMIDE
C0550643|T201|COMP|12329-9|LNC|chlorproPAMIDE|chlorproPAMIDE
C0550644|T201|COMP|12425-5|LNC|Chlorzoxazone|Chlorzoxazone
C0550645|T201|COMP|12374-5|LNC|cloBAZam|cloBAZam
C0550646|T201|COMP|10981-9|LNC|cloNIDine|cloNIDine
C0550647|T201|COMP|12314-1|LNC|Clorazepate|Clorazepate
C0550648|T201|COMP|12375-2|LNC|Clozapine+Norclozapine|Clozapine+Norclozapine
C0550649|T201|COMP|12784-5|LNC|Codeine.free|Codeine.free
C0550650|T201|COMP|12345-5|LNC|Cyclothiazide|Cyclothiazide
C0550651|T201|COMP|10982-7|LNC|Demeclocycline|Demeclocycline
C0550652|T201|COMP|12377-8|LNC|Demoxepam|Demoxepam
C0550653|T201|COMP|12709-2|LNC|Norastemizole|Norastemizole
C0550654|T201|COMP|12385-1|LNC|Desmethyldoxepin|Desmethyldoxepin
C0550655|T201|COMP|10983-5|LNC|Norparamethadione|Norparamethadione
C0550656|T201|COMP|12444-6|LNC|Nortrimipramine|Nortrimipramine
C0550657|T201|COMP|11072-6|LNC|Despropionylfentanyl|Despropionylfentanyl
C0550658|T201|COMP|11073-4|LNC|Despropionylfentanyl|Despropionylfentanyl
C0550659|T201|COMP|11234-2|LNC|Propoxyphene|Propoxyphene
C0550660|T201|COMP|12357-0|LNC|Propoxyphene|Propoxyphene
C0550661|T201|COMP|12326-5|LNC|Diamorphine|Diamorphine
C0550662|T201|COMP|12378-6|LNC|diazePAM|diazePAM
C0550663|T201|COMP|10984-3|LNC|Dicloxacillin|Dicloxacillin
C0550664|T201|COMP|12785-2|LNC|Dihydrocodeine.free|Dihydrocodeine.free
C0550665|T201|COMP|12391-9|LNC|dimenhyDRINATE|dimenhyDRINATE
C0550666|T201|COMP|12365-3|LNC|dimenhyDRINATE|dimenhyDRINATE
C0550667|T201|COMP|12372-9|LNC|Dimethylacetamide|Dimethylacetamide
C0550668|T201|COMP|12337-2|LNC|Dimethylsulfoxide|Dimethylsulfoxide
C0550669|T201|COMP|12292-9|LNC|Dimethyltryptamine|Dimethyltryptamine
C0550670|T201|COMP|12398-4|LNC|Diphenoxylate|Diphenoxylate
C0550671|T201|COMP|12366-1|LNC|Disopyramide|Disopyramide
C0550672|T201|COMP|12288-7|LNC|Diuretics|Diuretics
C0550673|T201|COMP|10985-0|LNC|Doxapram|Doxapram
C0550674|T201|COMP|10986-8|LNC|Doxycycline|Doxycycline
C0550675|T201|COMP|12399-2|LNC|Emetine|Emetine
C0550676|T201|COMP|12400-8|LNC|Emetine|Emetine
C0550677|T201|COMP|12298-6|LNC|Erythromycin|Erythromycin
C0550678|T201|COMP|11235-9|LNC|fentaNYL|fentaNYL
C0550679|T201|COMP|10987-6|LNC|Fluconazole|Fluconazole
C0550680|T201|COMP|12439-6|LNC|FLUoxetine|FLUoxetine
C0550681|T201|COMP|12605-2|LNC|Flurazepam|Flurazepam
C0550682|T201|COMP|12428-9|LNC|Flurbiprofen|Flurbiprofen
C0550683|T201|COMP|10988-4|LNC|fluvoxaMINE|fluvoxaMINE
C0550684|T201|COMP|11236-7|LNC|Gemfibrozil|Gemfibrozil
C0550685|T201|COMP|12402-4|LNC|Griseofulvin|Griseofulvin
C0550686|T201|COMP|12379-4|LNC|Halazepam|Halazepam
C0550687|T201|COMP|12493-3|LNC|Hexobarbital|Hexobarbital
C0550688|T201|COMP|11237-5|LNC|hydrALAZINE|hydrALAZINE
C0550689|T201|COMP|12336-4|LNC|hydrALAZINE|hydrALAZINE
C0550690|T201|COMP|12308-3|LNC|HYDROcodone|HYDROcodone
C0550691|T201|COMP|12786-0|LNC|HYDROcodone.free|HYDROcodone.free
C0550692|T201|COMP|12787-8|LNC|HYDROmorphone.free|HYDROmorphone.free
C0550693|T201|COMP|11238-3|LNC|Hydroxyalprazolam|Hydroxyalprazolam
C0550694|T201|COMP|12604-5|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C0550695|T201|COMP|12602-9|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C0550696|T201|COMP|12383-6|LNC|Hydroxytriazolam|Hydroxytriazolam
C0550697|T201|COMP|12432-1|LNC|Hydroxytriazolam|Hydroxytriazolam
C0550698|T201|COMP|11240-9|LNC|hydrOXYzine|hydrOXYzine
C0550699|T201|COMP|12324-0|LNC|hydrOXYzine|hydrOXYzine
C0550700|T201|COMP|11239-1|LNC|hydrOXYzine|hydrOXYzine
C0550701|T201|COMP|11241-7|LNC|Hyoscyamine|Hyoscyamine
C0550702|T201|COMP|12330-7|LNC|Hypoglycemics.oral|Hypoglycemics.oral
C0550704|T201|COMP|10989-2|LNC|Itraconazole|Itraconazole
C0550705|T201|COMP|11052-8|LNC|Ketamine|Ketamine
C0550706|T201|COMP|12327-3|LNC|Ketamine|Ketamine
C0550707|T201|COMP|10990-0|LNC|Ketoconazole|Ketoconazole
C0550709|T201|COMP|13455-1|LNC|Lithium.plasma/Lithium.RBC|Lithium.plasma/Lithium.RBC
C0550710|T201|COMP|12380-2|LNC|LORazepam|LORazepam
C0550711|T201|COMP|12341-4|LNC|Mazindol|Mazindol
C0550712|T201|COMP|12532-8|LNC|Meclizine|Meclizine
C0550713|T201|COMP|12403-2|LNC|Mephentermine|Mephentermine
C0550714|T201|COMP|12291-1|LNC|Mephentermine|Mephentermine
C0550715|T201|COMP|12315-8|LNC|Mephobarbital|Mephobarbital
C0550716|T201|COMP|11242-5|LNC|Mercaptopurine|Mercaptopurine
C0550717|T201|COMP|12367-9|LNC|Mesoridazine|Mesoridazine
C0550718|T201|COMP|12498-2|LNC|Metharbital|Metharbital
C0550719|T201|COMP|11243-3|LNC|Methadone|Methadone
C0550720|T201|COMP|12356-2|LNC|Methadone|Methadone
C0550721|T201|COMP|12353-9|LNC|Methaqualone|Methaqualone
C0550722|T201|COMP|10841-5|LNC|methazolAMIDE|methazolAMIDE
C0550723|T201|COMP|12346-3|LNC|Methyclothiazide|Methyclothiazide
C0550724|T201|COMP|12347-1|LNC|metOLazone|metOLazone
C0550725|T201|COMP|10991-8|LNC|metroNIDAZOLE|metroNIDAZOLE
C0550726|T201|COMP|12440-4|LNC|Midazolam|Midazolam
C0550727|T201|COMP|11244-1|LNC|Morphine.free|Morphine.free
C0550728|T201|COMP|12603-7|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0550730|T201|COMP|12406-5|LNC|Nadolol|Nadolol
C0550731|T201|COMP|10993-4|LNC|Nafcillin|Nafcillin
C0550732|T201|COMP|10994-2|LNC|Naltrexone|Naltrexone
C0550733|T201|COMP|12309-1|LNC|Naltrexone|Naltrexone
C0550734|T201|COMP|12544-3|LNC|Nefazodone|Nefazodone
C0550735|T201|COMP|10995-9|LNC|Neomycin|Neomycin
C0550736|T201|COMP|12294-5|LNC|Nicotine|Nicotine
C0550737|T201|COMP|12404-0|LNC|Nitroglycerin|Nitroglycerin
C0550738|T201|COMP|9776-6|LNC|Norchlordiazepoxide|Norchlordiazepoxide
C0550739|T201|COMP|10992-6|LNC|Norclozapine|Norclozapine
C0550740|T201|COMP|12386-9|LNC|Nordoxepin|Nordoxepin
C0550741|T201|COMP|12431-3|LNC|Norfenfluramine|Norfenfluramine
C0550742|T201|COMP|11074-2|LNC|Norfentanyl|Norfentanyl
C0550743|T201|COMP|11075-9|LNC|Norfentanyl|Norfentanyl
C0550744|T201|COMP|12445-3|LNC|Norfluoxetine|Norfluoxetine
C0550745|T201|COMP|10996-7|LNC|Normeperidine|Normeperidine
C0550746|T201|COMP|10890-2|LNC|Normethsuximide|Normethsuximide
C0550747|T201|COMP|10997-5|LNC|O-desmethylencainide|O-desmethylencainide
C0550748|T201|COMP|12438-8|LNC|Nortramadol|Nortramadol
C0550749|T201|COMP|12389-3|LNC|OLANZapine|OLANZapine
C0550750|T201|COMP|11245-8|LNC|Orphenadrine|Orphenadrine
C0550751|T201|COMP|12362-0|LNC|Oxazepam|Oxazepam
C0550752|T201|COMP|12381-0|LNC|Oxazepam|Oxazepam
C0550753|T201|COMP|12361-2|LNC|Oxazepam|Oxazepam
C0550754|T201|COMP|11246-6|LNC|oxyCODONE|oxyCODONE
C0550755|T201|COMP|10998-3|LNC|oxyCODONE|oxyCODONE
C0550756|T201|COMP|12789-4|LNC|oxyCODONE.free|oxyCODONE.free
C0550757|T201|COMP|12342-2|LNC|oxyMORphone|oxyMORphone
C0550758|T201|COMP|11247-4|LNC|oxyMORphone|oxyMORphone
C0550759|T201|COMP|10891-0|LNC|Oxyphenisatin|Oxyphenisatin
C0550760|T201|COMP|12550-0|LNC|Papaverine|Papaverine
C0550761|T201|COMP|10999-1|LNC|Paramethadione|Paramethadione
C0550762|T201|COMP|12488-3|LNC|PENTobarbital|PENTobarbital
C0550763|T201|COMP|12499-0|LNC|PENTobarbital|PENTobarbital
C0550765|T201|COMP|10892-8|LNC|Pentoxifylline|Pentoxifylline
C0550766|T201|COMP|11248-2|LNC|Pergolide|Pergolide
C0550767|T201|COMP|11249-0|LNC|Phenacemide|Phenacemide
C0550768|T201|COMP|12368-7|LNC|Phenacetin|Phenacetin
C0550769|T201|COMP|12484-2|LNC|PHENobarbital|PHENobarbital
C0550770|T201|COMP|12501-3|LNC|PHENobarbital|PHENobarbital
C0550771|T201|COMP|12388-5|LNC|Phenylethylmalonamide|Phenylethylmalonamide
C0550772|T201|COMP|12447-9|LNC|Phenylethylmalonamide|Phenylethylmalonamide
C0550773|T201|COMP|11250-8|LNC|Phenylethylmalonate|Phenylethylmalonate
C0550774|T201|COMP|12310-9|LNC|Phenytoin|Phenytoin
C0550775|T201|COMP|12410-7|LNC|Pimozide|Pimozide
C0550776|T201|COMP|11251-6|LNC|Piroxicam|Piroxicam
C0550777|T201|COMP|12300-0|LNC|Polythiazide|Polythiazide
C0550778|T201|COMP|12311-7|LNC|Prazepam|Prazepam
C0550779|T201|COMP|12727-4|LNC|prednisoLONE|prednisoLONE
C0550780|T201|COMP|12434-7|LNC|predniSONE|predniSONE
C0550781|T201|COMP|12387-7|LNC|Primidone|Primidone
C0550782|T201|COMP|12301-8|LNC|Procaine|Procaine
C0550783|T201|COMP|12290-3|LNC|Procyclidine|Procyclidine
C0550784|T201|COMP|12411-5|LNC|Promazine|Promazine
C0550785|T201|COMP|11000-7|LNC|Promethazine|Promethazine
C0550786|T201|COMP|11001-5|LNC|Pyrazinamide|Pyrazinamide
C0550787|T201|COMP|12546-8|LNC|Quinethazone|Quinethazone
C0550788|T201|COMP|12348-9|LNC|Quinethazone|Quinethazone
C0550789|T201|COMP|11252-4|LNC|Scopolamine|Scopolamine
C0550790|T201|COMP|11002-3|LNC|Scopolamine|Scopolamine
C0550791|T201|COMP|12489-1|LNC|Secobarbital|Secobarbital
C0550792|T201|COMP|12500-5|LNC|Secobarbital|Secobarbital
C0550793|T201|COMP|12416-4|LNC|Sotalol|Sotalol
C0550794|T201|COMP|12318-2|LNC|Spironolactone|Spironolactone
C0550795|T201|COMP|11253-2|LNC|Tacrolimus|Tacrolimus
C0550796|T201|COMP|12382-8|LNC|Temazepam|Temazepam
C0550797|T201|COMP|12418-0|LNC|Terfenadine|Terfenadine
C0550798|T201|COMP|12419-8|LNC|Terfenadine|Terfenadine
C0550799|T201|COMP|12325-7|LNC|Tetrahydrocortisone|Tetrahydrocortisone
C0550800|T201|COMP|12302-6|LNC|Theobromine|Theobromine
C0550801|T201|COMP|12303-4|LNC|Theobromine|Theobromine
C0550802|T201|COMP|12370-3|LNC|Thiopental|Thiopental
C0550803|T201|COMP|12319-0|LNC|Thioridazine|Thioridazine
C0550804|T201|COMP|12320-8|LNC|Thiothixene|Thiothixene
C0550805|T201|COMP|11003-1|LNC|Ticlopidine|Ticlopidine
C0550806|T201|COMP|12437-0|LNC|traMADol|traMADol
C0550807|T201|COMP|10893-6|LNC|Trenbolone|Trenbolone
C0550808|T201|COMP|12384-4|LNC|Triazolam|Triazolam
C0550809|T201|COMP|12349-7|LNC|Trichlormethiazide|Trichlormethiazide
C0550810|T201|COMP|11004-9|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0550811|T201|COMP|12321-6|LNC|Trifluoperazine|Trifluoperazine
C0550812|T201|COMP|12422-2|LNC|Triflupromazine|Triflupromazine
C0550813|T201|COMP|12322-4|LNC|Triflupromazine|Triflupromazine
C0550814|T201|COMP|12423-0|LNC|Trimeprazine|Trimeprazine
C0550815|T201|COMP|12800-9|LNC|Trimeprazine|Trimeprazine
C0550816|T201|COMP|12323-2|LNC|Trimeprazine|Trimeprazine
C0550817|T201|COMP|11005-6|LNC|Trimethoprim|Trimethoprim
C0550818|T201|COMP|12443-8|LNC|Trimipramine|Trimipramine
C0550819|T201|COMP|12548-4|LNC|Tybamate|Tybamate
C0550820|T201|COMP|12282-0|LNC|Warfarin|Warfarin
C0550821|T201|COMP|12545-0|LNC|Zomepirac|Zomepirac
C0550822|T201|COMP|13359-5|LNC|Character|Character
C0550823|T201|COMP|13360-3|LNC|Color|Color
C0550824|T201|COMP|12452-9|LNC|Epithelial cells|Epithelial cells
C0550825|T201|COMP|13361-1|LNC|Semen analysis panel|Semen analysis panel
C0550826|T201|COMP|12257-2|LNC|Spermatozoa.motile/100 spermatozoa^post vasectomy|Spermatozoa.motile/100 spermatozoa^post vasectomy
C0550827|T201|COMP|12256-4|LNC|Spermatozoa^post vasectomy|Spermatozoa^post vasectomy
C0550828|T201|COMP|13172-2|LNC|Complement C1q Ag|Complement C1q Ag
C0550829|T201|COMP|13086-4|LNC|C3 nephritic factor|C3 nephritic factor
C0550830|T201|COMP|13085-6|LNC|C4 nephritic factor|C4 nephritic factor
C0550831|T201|COMP|13117-7|LNC|Complement Sc5b-9 Ab|Complement Sc5b-9 Ab
C0550832|T201|COMP|13087-2|LNC|Complement alternate pathway AH50|Complement alternate pathway AH50
C0550833|T201|COMP|13088-0|LNC|Complement total hemolytic CH100|Complement total hemolytic CH100
C0550834|T201|COMP|11151-8|LNC|Hematocrit|Hematocrit
C0550835|T201|COMP|11271-4|LNC|Hematocrit|Hematocrit
C0550836|T201|COMP|11153-4|LNC|Hematocrit|Hematocrit
C0550837|T201|COMP|12711-8|LNC|Hemoglobin A region|Hemoglobin A region
C0550838|T201|COMP|12713-4|LNC|Hemoglobin C+E+O+A2 region|Hemoglobin C+E+O+A2 region
C0550839|T201|COMP|12710-0|LNC|Hemoglobin pattern|Hemoglobin pattern
C0550840|T201|COMP|12712-6|LNC|Hemoglobin S+D+G region|Hemoglobin S+D+G region
C0550841|T201|COMP|13055-9|LNC|Heparin|Heparin
C0550842|T201|COMP|12731-6|LNC|Interferon.alpha|Interferon.alpha
C0550843|T201|COMP|12730-8|LNC|Interferon.beta|Interferon.beta
C0550844|T201|COMP|12729-0|LNC|Interferon.gamma|Interferon.gamma
C0550845|T201|COMP|12732-4|LNC|Interleukin 12|Interleukin 12
C0550846|T201|COMP|12227-5|LNC|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C0550847|T201|COMP|11272-2|LNC|Erythrocyte mean corpuscular volume|Erythrocyte mean corpuscular volume
C0550848|T201|COMP|12243-2|LNC|Platelets|Platelets
C0550849|T201|COMP|13298-5|LNC|HLA-A|HLA-A
C0550850|T201|COMP|13300-9|LNC|HLA-A+B|HLA-A+B
C0550851|T201|COMP|13301-7|LNC|HLA-A+B+Bw|HLA-A+B+Bw
C0550852|T201|COMP|13303-3|LNC|HLA-A+B+C|HLA-A+B+C
C0550853|T201|COMP|13299-3|LNC|HLA-B|HLA-B
C0550854|T201|COMP|13302-5|LNC|HLA-C|HLA-C
C0550855|T201|COMP|12285-3|LNC|HLA-DP|HLA-DP
C0550856|T201|COMP|13305-8|LNC|HLA-DQ|HLA-DQ
C0550857|T201|COMP|13307-4|LNC|HLA-DQ alpha|HLA-DQ alpha
C0550858|T201|COMP|10842-3|LNC|HLA-DQ1|HLA-DQ1
C0550859|T201|COMP|10843-1|LNC|HLA-DQ2|HLA-DQ2
C0550860|T201|COMP|10844-9|LNC|HLA-DQ3|HLA-DQ3
C0550861|T201|COMP|10845-6|LNC|HLA-DQ4|HLA-DQ4
C0550862|T201|COMP|13304-1|LNC|HLA-DR|HLA-DR
C0550863|T201|COMP|13306-6|LNC|HLA-DR beta|HLA-DR beta
C0550864|T201|COMP|13192-0|LNC|Adenovirus Ab|Adenovirus Ab
C0550865|T201|COMP|13193-8|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C0550866|T201|COMP|11583-2|LNC|Aspergillus fumigatus 1 Ab|Aspergillus fumigatus 1 Ab
C0550867|T201|COMP|11592-3|LNC|Aspergillus fumigatus 6 Ab|Aspergillus fumigatus 6 Ab
C0550868|T201|COMP|13194-6|LNC|Aspergillus glaucus Ab|Aspergillus glaucus Ab
C0550869|T201|COMP|10894-4|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C0550870|T201|COMP|11584-0|LNC|Aureobasidium pullulans Ab|Aureobasidium pullulans Ab
C0550871|T201|COMP|11467-8|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0550872|T201|COMP|11468-6|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0550873|T201|COMP|11469-4|LNC|Bacillus anthracis|Bacillus anthracis
C0550874|T201|COMP|12178-0|LNC|Bacteria|Bacteria
C0550875|T201|COMP|13201-9|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0550876|T201|COMP|11585-7|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C0550877|T201|COMP|11550-1|LNC|Borrelia burgdorferi|Borrelia burgdorferi
C0550878|T201|COMP|12866-0|LNC|Borrelia burgdorferi 18kD Ab|Borrelia burgdorferi 18kD Ab
C0550879|T201|COMP|12883-5|LNC|Borrelia burgdorferi 18kD Ab|Borrelia burgdorferi 18kD Ab
C0550880|T201|COMP|12864-5|LNC|Borrelia burgdorferi 25kD Ab|Borrelia burgdorferi 25kD Ab
C0550881|T201|COMP|12888-4|LNC|Borrelia burgdorferi 25kD Ab|Borrelia burgdorferi 25kD Ab
C0550882|T201|COMP|12879-3|LNC|Borrelia burgdorferi 25kD Ab|Borrelia burgdorferi 25kD Ab
C0550883|T201|COMP|12865-2|LNC|Borrelia burgdorferi 29kD Ab|Borrelia burgdorferi 29kD Ab
C0550884|T201|COMP|12882-7|LNC|Borrelia burgdorferi 29kD Ab|Borrelia burgdorferi 29kD Ab
C0550885|T201|COMP|12878-5|LNC|Borrelia burgdorferi 29kD Ab|Borrelia burgdorferi 29kD Ab
C0550886|T201|COMP|12869-4|LNC|Borrelia burgdorferi 30kD Ab|Borrelia burgdorferi 30kD Ab
C0550887|T201|COMP|12889-2|LNC|Borrelia burgdorferi 30kD Ab|Borrelia burgdorferi 30kD Ab
C0550888|T201|COMP|12892-6|LNC|Borrelia burgdorferi 30kD Ab|Borrelia burgdorferi 30kD Ab
C0550889|T201|COMP|12860-3|LNC|Borrelia burgdorferi 39kD Ab|Borrelia burgdorferi 39kD Ab
C0550890|T201|COMP|12884-3|LNC|Borrelia burgdorferi 39kD Ab|Borrelia burgdorferi 39kD Ab
C0550891|T201|COMP|12863-7|LNC|Borrelia burgdorferi 41kD Ab|Borrelia burgdorferi 41kD Ab
C0550892|T201|COMP|12887-6|LNC|Borrelia burgdorferi 41kD Ab|Borrelia burgdorferi 41kD Ab
C0550893|T201|COMP|12891-8|LNC|Borrelia burgdorferi 41kD Ab|Borrelia burgdorferi 41kD Ab
C0550894|T201|COMP|12890-0|LNC|Borrelia burgdorferi 45kD Ab|Borrelia burgdorferi 45kD Ab
C0550895|T201|COMP|12868-6|LNC|Borrelia burgdorferi 47kD Ab|Borrelia burgdorferi 47kD Ab
C0550896|T201|COMP|12881-9|LNC|Borrelia burgdorferi 47kD Ab|Borrelia burgdorferi 47kD Ab
C0550897|T201|COMP|12877-7|LNC|Borrelia burgdorferi 47kD Ab|Borrelia burgdorferi 47kD Ab
C0550898|T201|COMP|12867-8|LNC|Borrelia burgdorferi 58kD Ab|Borrelia burgdorferi 58kD Ab
C0550899|T201|COMP|12880-1|LNC|Borrelia burgdorferi 58kD Ab|Borrelia burgdorferi 58kD Ab
C0550900|T201|COMP|12896-7|LNC|Borrelia burgdorferi 58kD Ab|Borrelia burgdorferi 58kD Ab
C0550901|T201|COMP|12862-9|LNC|Borrelia burgdorferi 66kD Ab|Borrelia burgdorferi 66kD Ab
C0550902|T201|COMP|12886-8|LNC|Borrelia burgdorferi 66kD Ab|Borrelia burgdorferi 66kD Ab
C0550903|T201|COMP|12861-1|LNC|Borrelia burgdorferi 88kD Ab|Borrelia burgdorferi 88kD Ab
C0550904|T201|COMP|12885-0|LNC|Borrelia burgdorferi 88kD Ab|Borrelia burgdorferi 88kD Ab
C0550905|T201|COMP|12873-6|LNC|Borrelia burgdorferi 88kD Ab|Borrelia burgdorferi 88kD Ab
C0550906|T201|COMP|12874-4|LNC|Borrelia burgdorferi 93kD Ab|Borrelia burgdorferi 93kD Ab
C0550907|T201|COMP|11006-4|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0550909|T201|COMP|12781-1|LNC|Borrelia burgdorferi Ab band pattern|Borrelia burgdorferi Ab band pattern
C0550910|T201|COMP|13204-3|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0550911|T201|COMP|13202-7|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0550912|T201|COMP|13206-8|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0550913|T201|COMP|13502-0|LNC|Borrelia burgdorferi Ab.IgG band pattern|Borrelia burgdorferi Ab.IgG band pattern
C0550914|T201|COMP|13205-0|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0550915|T201|COMP|13203-5|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0550916|T201|COMP|13207-6|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0550917|T201|COMP|13503-8|LNC|Borrelia burgdorferi Ab.IgM band pattern|Borrelia burgdorferi Ab.IgM band pattern
C0550918|T201|COMP|11007-2|LNC|Borrelia burgdorferi Ag|Borrelia burgdorferi Ag
C0550919|T201|COMP|10846-4|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C0550920|T201|COMP|11551-9|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C0550921|T201|COMP|10847-2|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C0550922|T201|COMP|13208-4|LNC|Borrelia hermsii Ab.IgG|Borrelia hermsii Ab.IgG
C0550923|T201|COMP|13209-2|LNC|Borrelia hermsii Ab.IgM|Borrelia hermsii Ab.IgM
C0550924|T201|COMP|11586-5|LNC|Brucella abortus Ab|Brucella abortus Ab
C0550925|T201|COMP|13212-6|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C0550926|T201|COMP|13213-4|LNC|Brucella abortus Ab.IgM|Brucella abortus Ab.IgM
C0550927|T201|COMP|11587-3|LNC|Brucella canis Ab|Brucella canis Ab
C0550928|T201|COMP|13214-2|LNC|Brucella canis Ab.IgG|Brucella canis Ab.IgG
C0550929|T201|COMP|13215-9|LNC|Brucella canis Ab.IgM|Brucella canis Ab.IgM
C0550930|T201|COMP|11588-1|LNC|Brucella melitensis Ab|Brucella melitensis Ab
C0550931|T201|COMP|13211-8|LNC|Brucella sp Ab.IgA|Brucella sp Ab.IgA
C0550932|T201|COMP|13210-0|LNC|Brucella sp Ab.IgG|Brucella sp Ab.IgG
C0550933|T201|COMP|11589-9|LNC|Brucella suis Ab|Brucella suis Ab
C0550934|T201|COMP|11102-1|LNC|Charcot-leyden crystals|Charcot-leyden crystals
C0550935|T201|COMP|11254-0|LNC|Chlamydophila pneumoniae Ab|Chlamydophila pneumoniae Ab
C0550936|T201|COMP|10848-0|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C0550937|T201|COMP|10849-8|LNC|Chlamydia sp Ab.IgM|Chlamydia sp Ab.IgM
C0550939|T201|COMP|13217-5|LNC|Chlamydia trachomatis B Ab|Chlamydia trachomatis B Ab
C0550941|T201|COMP|13220-9|LNC|Chlamydia trachomatis C Ab.IgM|Chlamydia trachomatis C Ab.IgM
C0550942|T201|COMP|13218-3|LNC|Chlamydia trachomatis C Ab|Chlamydia trachomatis C Ab
C0550944|T201|COMP|13221-7|LNC|Chlamydia trachomatis G+F+K Ab.IgM|Chlamydia trachomatis G+F+K Ab.IgM
C0550945|T201|COMP|13219-1|LNC|Chlamydia trachomatis G+F+K Ab|Chlamydia trachomatis G+F+K Ab
C0550946|T201|COMP|11470-2|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C0550947|T201|COMP|10895-1|LNC|Clostridioides difficile toxin B|Clostridioides difficile toxin B
C0550948|T201|COMP|13292-8|LNC|Colorado tick fever virus Ab.IgG|Colorado tick fever virus Ab.IgG
C0550949|T201|COMP|13293-6|LNC|Colorado tick fever virus Ab.IgM|Colorado tick fever virus Ab.IgM
C0550950|T201|COMP|13227-4|LNC|Corynebacterium diphtheriae Ab.IgG|Corynebacterium diphtheriae Ab.IgG
C0550951|T201|COMP|13232-4|LNC|Coxsackievirus A Ab|Coxsackievirus A Ab
C0550952|T201|COMP|13297-7|LNC|Coxsackievirus A1 Ab|Coxsackievirus A1 Ab
C0550953|T201|COMP|13295-1|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C0550954|T201|COMP|11590-7|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C0550955|T201|COMP|13296-9|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C0550956|T201|COMP|13235-7|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C0550957|T201|COMP|13233-2|LNC|Coxsackievirus A2 Ab|Coxsackievirus A2 Ab
C0550958|T201|COMP|11591-5|LNC|Coxsackievirus A2 Ab|Coxsackievirus A2 Ab
C0550959|T201|COMP|11599-8|LNC|Coxsackievirus A21 Ab|Coxsackievirus A21 Ab
C0550960|T201|COMP|13234-0|LNC|Coxsackievirus A4 Ab|Coxsackievirus A4 Ab
C0550961|T201|COMP|11593-1|LNC|Coxsackievirus A4 Ab|Coxsackievirus A4 Ab
C0550962|T201|COMP|11472-8|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C0550963|T201|COMP|11471-0|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C0550964|T201|COMP|11473-6|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C0550965|T201|COMP|10850-6|LNC|Cyclospora cayetanensis|Cyclospora cayetanensis
C0550966|T201|COMP|11008-0|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0550967|T201|COMP|13225-8|LNC|Cytomegalovirus Ab.IgG^1st specimen|Cytomegalovirus Ab.IgG^1st specimen
C0550968|T201|COMP|13226-6|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0550969|T201|COMP|13228-2|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C0550970|T201|COMP|10897-7|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C0550971|T201|COMP|10896-9|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C0550972|T201|COMP|13229-0|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C0550973|T201|COMP|10899-3|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C0550974|T201|COMP|10898-5|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C0550975|T201|COMP|11581-6|LNC|Ebola virus Ab|Ebola virus Ab
C0550976|T201|COMP|11594-9|LNC|Echovirus 16 Ab|Echovirus 16 Ab
C0550977|T201|COMP|11595-6|LNC|Echovirus 18 Ab|Echovirus 18 Ab
C0550978|T201|COMP|11601-2|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C0550979|T201|COMP|13195-3|LNC|Ehrlichia chaffeensis Ab|Ehrlichia chaffeensis Ab
C0550980|T201|COMP|13196-1|LNC|Ehrlichia sp Ab.IgG|Ehrlichia sp Ab.IgG
C0550981|T201|COMP|13197-9|LNC|Ehrlichia sp Ab.IgM|Ehrlichia sp Ab.IgM
C0550982|T201|COMP|13316-5|LNC|Enterococcus species.vancomycin resistant|Enterococcus species.vancomycin resistant
C0550983|T201|COMP|13238-1|LNC|Epstein Barr virus Ab|Epstein Barr virus Ab
C0550984|T201|COMP|13239-9|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0550985|T201|COMP|13236-5|LNC|Epstein Barr virus early diffuse Ab|Epstein Barr virus early diffuse Ab
C0550986|T201|COMP|13237-3|LNC|Epstein Barr virus early restricted Ab|Epstein Barr virus early restricted Ab
C0550987|T201|COMP|12212-7|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0550988|T201|COMP|11009-8|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0550989|T201|COMP|11010-6|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0550990|T201|COMP|13318-1|LNC|Escherichia coli enteroinvasive identified|Escherichia coli enteroinvasive identified
C0550991|T201|COMP|13329-8|LNC|Escherichia coli labile toxin|Escherichia coli labile toxin
C0550992|T201|COMP|12276-2|LNC|Escherichia coli O157:H7|Escherichia coli O157:H7
C0550993|T201|COMP|10851-4|LNC|Escherichia coli O157:H7|Escherichia coli O157:H7
C0550994|T201|COMP|13244-9|LNC|Filaria Ab.IgG|Filaria Ab.IgG
C0550995|T201|COMP|13245-6|LNC|Filaria Ab.IgM|Filaria Ab.IgM
C0550997|T201|COMP|11255-7|LNC|Haemophilus ducreyi|Haemophilus ducreyi
C0550998|T201|COMP|11256-5|LNC|Haemophilus influenzae B Ab.IgG|Haemophilus influenzae B Ab.IgG
C0550999|T201|COMP|13246-4|LNC|Haemophilus influenzae B Ab|Haemophilus influenzae B Ab
C0551000|T201|COMP|11257-3|LNC|Haemophilus influenzae B Ab.IgG|Haemophilus influenzae B Ab.IgG
C0551001|T201|COMP|13289-4|LNC|Hantavirus hantaan Ab|Hantavirus hantaan Ab
C0551002|T201|COMP|13126-8|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C0551003|T201|COMP|11258-1|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C0551004|T201|COMP|10900-9|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0551005|T201|COMP|11076-7|LNC|Hepatitis C virus 5-1-1 Ab|Hepatitis C virus 5-1-1 Ab
C0551006|T201|COMP|11077-5|LNC|Hepatitis C virus superoxide dismutase Ab|Hepatitis C virus superoxide dismutase Ab
C0551008|T201|COMP|11011-4|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C0551009|T201|COMP|11259-9|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C0551010|T201|COMP|13248-0|LNC|Hepatitis D virus Ab|Hepatitis D virus Ab
C0551011|T201|COMP|13294-4|LNC|Hepatitis E virus Ab|Hepatitis E virus Ab
C0551012|T201|COMP|13505-3|LNC|Herpes simplex virus 1+2 Ab pattern|Herpes simplex virus 1+2 Ab pattern
C0551013|T201|COMP|13249-8|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C0551014|T201|COMP|13501-2|LNC|Herpes simplex virus 2 Ab pattern|Herpes simplex virus 2 Ab pattern
C0551015|T201|COMP|13324-9|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C0551016|T201|COMP|13251-4|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C0551017|T201|COMP|13323-1|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C0551018|T201|COMP|13252-2|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C0551019|T201|COMP|13250-6|LNC|Herpes virus 6 Ab.IgG+IgM|Herpes virus 6 Ab.IgG+IgM
C0551020|T201|COMP|11610-3|LNC|Heterophile Ab|Heterophile Ab
C0551021|T201|COMP|12456-0|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C0551022|T201|COMP|12455-2|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C0551023|T201|COMP|13499-9|LNC|HIV 1 Ab band pattern|HIV 1 Ab band pattern
C0551024|T201|COMP|12893-4|LNC|HIV 1 gp105 Ab|HIV 1 gp105 Ab
C0551025|T201|COMP|12870-2|LNC|HIV 1 gp34 Ab|HIV 1 gp34 Ab
C0551026|T201|COMP|12872-8|LNC|HIV 1 p15 Ab|HIV 1 p15 Ab
C0551027|T201|COMP|12859-5|LNC|HIV 1 p18 Ab|HIV 1 p18 Ab
C0551028|T201|COMP|12855-3|LNC|HIV 1 p23 Ab|HIV 1 p23 Ab
C0551029|T201|COMP|12871-0|LNC|HIV 1 p26 Ab|HIV 1 p26 Ab
C0551030|T201|COMP|12857-9|LNC|HIV 1 p28 Ab|HIV 1 p28 Ab
C0551031|T201|COMP|12858-7|LNC|HIV 1 p32 Ab|HIV 1 p32 Ab
C0551032|T201|COMP|12876-9|LNC|HIV 1 p53 Ab|HIV 1 p53 Ab
C0551033|T201|COMP|12895-9|LNC|HIV 1 p58 Ab|HIV 1 p58 Ab
C0551034|T201|COMP|12875-1|LNC|HIV 1 p64 Ab|HIV 1 p64 Ab
C0551035|T201|COMP|12856-1|LNC|HIV 1 p65 Ab|HIV 1 p65 Ab
C0551036|T201|COMP|12894-2|LNC|HIV 1 p68 Ab|HIV 1 p68 Ab
C0551037|T201|COMP|10901-7|LNC|HIV 2 gp125 Ab|HIV 2 gp125 Ab
C0551038|T201|COMP|10902-5|LNC|HIV 2 gp36 Ab|HIV 2 gp36 Ab
C0551039|T201|COMP|11078-3|LNC|HIV 2 gp80 Ab|HIV 2 gp80 Ab
C0551040|T201|COMP|11079-1|LNC|HIV 2 p26 Ab|HIV 2 p26 Ab
C0551041|T201|COMP|11080-9|LNC|HIV 2 p53 Ab|HIV 2 p53 Ab
C0551042|T201|COMP|11081-7|LNC|HIV 2 p56 Ab|HIV 2 p56 Ab
C0551043|T201|COMP|11082-5|LNC|HIV 2 p68 Ab|HIV 2 p68 Ab
C0551044|T201|COMP|11609-5|LNC|HTLV I Ab|HTLV I Ab
C0551045|T201|COMP|11260-7|LNC|HTLV I Ab|HTLV I Ab
C0551046|T201|COMP|13247-2|LNC|HTLV I+II Ab|HTLV I+II Ab
C0551047|T201|COMP|10903-3|LNC|Hyaluronidase Ab|Hyaluronidase Ab
C0551048|T201|COMP|11474-4|LNC|Hydatid cyst identified|Hydatid cyst identified
C0551049|T201|COMP|10853-0|LNC|Isospora belli|Isospora belli
C0551050|T201|COMP|11608-7|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0551051|T201|COMP|11607-9|LNC|Junin virus Ab|Junin virus Ab
C0551052|T201|COMP|10904-1|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C0551053|T201|COMP|10905-8|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C0551054|T201|COMP|13255-5|LNC|Legionella longbeachae 1+2 Ab|Legionella longbeachae 1+2 Ab
C0551055|T201|COMP|13253-0|LNC|Legionella non pneumophila sp Ab|Legionella non pneumophila sp Ab
C0551056|T201|COMP|13254-8|LNC|Legionella pneumophila atypical Ab|Legionella pneumophila atypical Ab
C0551057|T201|COMP|13258-9|LNC|Leishmania braziliensis Ab.IgG|Leishmania braziliensis Ab.IgG
C0551058|T201|COMP|13259-7|LNC|Leishmania braziliensis Ab.IgM|Leishmania braziliensis Ab.IgM
C0551059|T201|COMP|13256-3|LNC|Leishmania donovani Ab.IgG|Leishmania donovani Ab.IgG
C0551060|T201|COMP|13257-1|LNC|Leishmania donovani Ab.IgM|Leishmania donovani Ab.IgM
C0551061|T201|COMP|13260-5|LNC|Leishmania mexicana Ab.IgG|Leishmania mexicana Ab.IgG
C0551062|T201|COMP|13261-3|LNC|Leishmania mexicana Ab.IgM|Leishmania mexicana Ab.IgM
C0551063|T201|COMP|13262-1|LNC|Leishmania tropica Ab.IgG|Leishmania tropica Ab.IgG
C0551064|T201|COMP|13263-9|LNC|Leishmania tropica Ab.IgM|Leishmania tropica Ab.IgM
C0551065|T201|COMP|13264-7|LNC|Leptospira sp Ab.IgG|Leptospira sp Ab.IgG
C0551066|T201|COMP|13265-4|LNC|Leptospira sp Ab.IgM|Leptospira sp Ab.IgM
C0551067|T201|COMP|11606-1|LNC|Leptospira interrogans Ab|Leptospira interrogans Ab
C0551068|T201|COMP|11605-3|LNC|Lymphocytic choriomeningitis virus Ab|Lymphocytic choriomeningitis virus Ab
C0551069|T201|COMP|12232-5|LNC|Measles virus Ag|Measles virus Ag
C0551070|T201|COMP|10854-8|LNC|Microfilaria sp identified|Microfilaria sp identified
C0551071|T201|COMP|12281-2|LNC|Bacteria identified|Bacteria identified
C0551072|T201|COMP|11261-5|LNC|Bacteria identified|Bacteria identified
C0551073|T201|COMP|13314-0|LNC|Bacteria identified|Bacteria identified
C0551074|T201|COMP|13315-7|LNC|Bacteria identified|Bacteria identified
C0551075|T201|COMP|11475-1|LNC|Microorganism identified|Microorganism identified
C0551077|T201|COMP|11552-7|LNC|Microscopic exam|Microscopic exam
C0551078|T201|COMP|10855-5|LNC|Ova & parasites identified|Ova & parasites identified
C0551088|T201|COMP|13319-9|LNC|Ova & parasites identified^2nd specimen|Ova & parasites identified^2nd specimen
C0551089|T201|COMP|13320-7|LNC|Ova & parasites identified^3rd specimen|Ova & parasites identified^3rd specimen
C0551090|T201|COMP|10857-1|LNC|Microsporidia identified|Microsporidia identified
C0551091|T201|COMP|13266-2|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0551092|T201|COMP|13267-0|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C0551093|T201|COMP|12237-4|LNC|Mumps virus Ag|Mumps virus Ag
C0551094|T201|COMP|13270-4|LNC|Mycoplasma pneumoniae Ab.IgA|Mycoplasma pneumoniae Ab.IgA
C0551095|T201|COMP|13268-8|LNC|Mycoplasma pneumoniae Ab^1st specimen|Mycoplasma pneumoniae Ab^1st specimen
C0551096|T201|COMP|13269-6|LNC|Mycoplasma pneumoniae Ab^2nd specimen|Mycoplasma pneumoniae Ab^2nd specimen
C0551097|T201|COMP|13271-2|LNC|Neisseria meningitidis serogroup A Ab|Neisseria meningitidis serogroup A Ab
C0551098|T201|COMP|13272-0|LNC|Neisseria meningitidis serogroup C Ab|Neisseria meningitidis serogroup C Ab
C0551099|T201|COMP|13321-5|LNC|Human papilloma virus Ab.IgG|Human papilloma virus Ab.IgG
C0551100|T201|COMP|13322-3|LNC|Human papilloma virus Ab.IgM|Human papilloma virus Ab.IgM
C0551101|T201|COMP|12222-6|LNC|Human papilloma virus Ag|Human papilloma virus Ag
C0551102|T201|COMP|12223-4|LNC|Human papilloma virus 16+18 Ag|Human papilloma virus 16+18 Ag
C0551103|T201|COMP|11083-3|LNC|Human papilloma virus identified|Human papilloma virus identified
C0551104|T201|COMP|11481-9|LNC|Human papilloma virus identified|Human papilloma virus identified
C0551105|T201|COMP|13327-2|LNC|Parainfluenza virus Ag|Parainfluenza virus Ag
C0551106|T201|COMP|11262-3|LNC|Parainfluenza virus 3 Ab.IgG|Parainfluenza virus 3 Ab.IgG
C0551107|T201|COMP|11263-1|LNC|Parainfluenza virus 3 Ab.IgM|Parainfluenza virus 3 Ab.IgM
C0551108|T201|COMP|13326-4|LNC|Pneumocystis sp identified|Pneumocystis sp identified
C0551109|T201|COMP|11604-6|LNC|Burkholderia pseudomallei Ab|Burkholderia pseudomallei Ab
C0551110|T201|COMP|11084-1|LNC|Reagin Ab|Reagin Ab
C0551111|T201|COMP|11012-2|LNC|Reovirus Ab|Reovirus Ab
C0551112|T201|COMP|13199-5|LNC|Rickettsia conorii Ab.IgG|Rickettsia conorii Ab.IgG
C0551113|T201|COMP|13200-1|LNC|Rickettsia conorii Ab.IgM|Rickettsia conorii Ab.IgM
C0551114|T201|COMP|11482-7|LNC|Rickettsia rickettsii RNA|Rickettsia rickettsii RNA
C0551115|T201|COMP|13325-6|LNC|Bartonella sp identified|Bartonella sp identified
C0551116|T201|COMP|13281-1|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0551117|T201|COMP|13279-5|LNC|Rubella virus Ab.IgG^1st specimen|Rubella virus Ab.IgG^1st specimen
C0551118|T201|COMP|13280-3|LNC|Rubella virus Ab.IgG^2nd specimen|Rubella virus Ab.IgG^2nd specimen
C0551119|T201|COMP|13282-9|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C0551120|T201|COMP|12251-5|LNC|Rubella virus Ag|Rubella virus Ag
C0551121|T201|COMP|13283-7|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C0551122|T201|COMP|13328-0|LNC|Measles virus Ag|Measles virus Ag
C0551123|T201|COMP|13230-8|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C0551124|T201|COMP|10906-6|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C0551125|T201|COMP|13231-6|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C0551126|T201|COMP|10907-4|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C0551127|T201|COMP|11264-9|LNC|Salmonella paratyphi A Ab|Salmonella paratyphi A Ab
C0551128|T201|COMP|11265-6|LNC|Salmonella paratyphi B Ab|Salmonella paratyphi B Ab
C0551129|T201|COMP|11603-8|LNC|Salmonella sp Ab|Salmonella sp Ab
C0551130|T201|COMP|13284-5|LNC|Salmonella typhi H D Ab|Salmonella typhi H D Ab
C0551131|T201|COMP|13285-2|LNC|Salmonella typhi O D Ab|Salmonella typhi O D Ab
C0551132|T201|COMP|13277-9|LNC|Schistosoma sp Ab.IgG|Schistosoma sp Ab.IgG
C0551133|T201|COMP|13278-7|LNC|Schistosoma sp Ab.IgM|Schistosoma sp Ab.IgM
C0551134|T201|COMP|11085-8|LNC|Schistosoma sp identified|Schistosoma sp identified
C0551135|T201|COMP|11602-0|LNC|Shigella boydii Ab|Shigella boydii Ab
C0551136|T201|COMP|11596-4|LNC|Shigella dysenteriae Ab|Shigella dysenteriae Ab
C0551137|T201|COMP|11600-4|LNC|Shigella flexneri Ab|Shigella flexneri Ab
C0551138|T201|COMP|11611-1|LNC|Shigella sonnei Ab|Shigella sonnei Ab
C0551139|T201|COMP|13243-1|LNC|Sporothrix schenckii Ab.IgA|Sporothrix schenckii Ab.IgA
C0551140|T201|COMP|13241-5|LNC|Sporothrix schenckii Ab.IgG|Sporothrix schenckii Ab.IgG
C0551141|T201|COMP|13242-3|LNC|Sporothrix schenckii Ab.IgM|Sporothrix schenckii Ab.IgM
C0551142|T201|COMP|13273-8|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C0551144|T201|COMP|11266-4|LNC|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C0551145|T201|COMP|11267-2|LNC|Streptococcus.beta-hemolytic|Streptococcus.beta-hemolytic
C0551146|T201|COMP|13131-8|LNC|Streptococcus pneumoniae 1 Ab|Streptococcus pneumoniae 1 Ab
C0551149|T201|COMP|13135-9|LNC|Streptococcus pneumoniae 12 Ab|Streptococcus pneumoniae 12 Ab
C0551155|T201|COMP|13136-7|LNC|Streptococcus pneumoniae Danish serotype 18C Ab|Streptococcus pneumoniae Danish serotype 18C Ab
C0551158|T201|COMP|13137-5|LNC|Streptococcus pneumoniae 19 Ab|Streptococcus pneumoniae 19 Ab
C0551160|T201|COMP|13159-9|LNC|Streptococcus pneumoniae 19 Ab^1st specimen|Streptococcus pneumoniae 19 Ab^1st specimen
C0551162|T201|COMP|13138-3|LNC|Streptococcus pneumoniae 23 Ab|Streptococcus pneumoniae 23 Ab
C0551168|T201|COMP|13132-6|LNC|Streptococcus pneumoniae 4 Ab|Streptococcus pneumoniae 4 Ab
C0551171|T201|COMP|13167-2|LNC|Streptococcus pneumoniae Danish serotype 7F Ab|Streptococcus pneumoniae Danish serotype 7F Ab
C0551172|T201|COMP|13168-0|LNC|Streptococcus pneumoniae 6+26 Ab|Streptococcus pneumoniae 6+26 Ab
C0551173|T201|COMP|13133-4|LNC|Streptococcus pneumoniae Danish serotype 6B Ab|Streptococcus pneumoniae Danish serotype 6B Ab
C0551176|T201|COMP|10908-2|LNC|Streptococcus pneumoniae 7 Ab.IgG|Streptococcus pneumoniae 7 Ab.IgG
C0551179|T201|COMP|13134-2|LNC|Streptococcus pneumoniae 8 Ab|Streptococcus pneumoniae 8 Ab
C0551180|T201|COMP|13149-0|LNC|Streptococcus pneumoniae 8 Ab^1st specimen|Streptococcus pneumoniae 8 Ab^1st specimen
C0551181|T201|COMP|13150-8|LNC|Streptococcus pneumoniae 8 Ab^2nd specimen|Streptococcus pneumoniae 8 Ab^2nd specimen
C0551184|T201|COMP|11086-6|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C0551185|T201|COMP|11268-0|LNC|Streptococcus pyogenes|Streptococcus pyogenes
C0551186|T201|COMP|11269-8|LNC|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C0551187|T201|COMP|12259-8|LNC|Streptococcus pyogenes enzyme Ab|Streptococcus pyogenes enzyme Ab
C0551188|T201|COMP|10858-9|LNC|Teichoate Ab|Teichoate Ab
C0551189|T201|COMP|13198-7|LNC|Thermoactinomyces sp Ab|Thermoactinomyces sp Ab
C0551190|T201|COMP|13274-6|LNC|Toxocara canis Ab|Toxocara canis Ab
C0551193|T201|COMP|11598-0|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C0551194|T201|COMP|12261-4|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0551195|T201|COMP|13286-0|LNC|Toxoplasma gondii Ab.IgG^2nd specimen|Toxoplasma gondii Ab.IgG^2nd specimen
C0551196|T201|COMP|12262-2|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0551197|T201|COMP|13287-8|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C0551198|T201|COMP|12263-0|LNC|Epstein Barr virus early diffuse Ab|Epstein Barr virus early diffuse Ab
C0551199|T201|COMP|13288-6|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0551200|T201|COMP|11597-2|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0551201|T201|COMP|13291-0|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C0551202|T201|COMP|13290-2|LNC|Trypanosoma cruzi Ab.IgM|Trypanosoma cruzi Ab.IgM
C0551203|T201|COMP|10859-7|LNC|Trypanosoma sp|Trypanosoma sp
C0551204|T201|COMP|12271-3|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C0551205|T201|COMP|10860-5|LNC|Varicella zoster virus|Varicella zoster virus
C0551206|T201|COMP|11483-5|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C0551207|T201|COMP|11270-6|LNC|Viral inclusion bodies|Viral inclusion bodies
C0551208|T201|COMP|11484-3|LNC|Virus identified|Virus identified
C0551209|T201|COMP|12272-1|LNC|Virus identified|Virus identified
C0551210|T201|COMP|11582-4|LNC|Wuchereria bancrofti Ab|Wuchereria bancrofti Ab
C0551211|T201|COMP|12275-4|LNC|Yeast|Yeast
C0551212|T201|COMP|13363-7|LNC|Collection duration|Collection duration
C0551214|T201|COMP|13358-7|LNC|Collection time|Collection time
C0551215|T201|COMP|12426-3|LNC|Brodifacoum|Brodifacoum
C0551216|T201|COMP|12397-6|LNC|Colchicine|Colchicine
C0551217|T201|COMP|12430-5|LNC|Cumene|Cumene
C0551218|T201|COMP|12306-7|LNC|Cyclohexane|Cyclohexane
C0551219|T201|COMP|12995-7|LNC|Cyclohexanone|Cyclohexanone
C0551220|T201|COMP|12312-5|LNC|Cyclopropane|Cyclopropane
C0551221|T201|COMP|12339-8|LNC|Diquat|Diquat
C0551222|T201|COMP|12606-0|LNC|Dolichol|Dolichol
C0551223|T201|COMP|12737-3|LNC|Endothelin|Endothelin
C0551224|T201|COMP|12999-9|LNC|Epichlorohydrin|Epichlorohydrin
C0551225|T201|COMP|12401-6|LNC|Ethinamate|Ethinamate
C0551226|T201|COMP|12299-4|LNC|Ethinamate|Ethinamate
C0551227|T201|COMP|12335-6|LNC|Halothane|Halothane
C0551229|T201|COMP|12736-5|LNC|Hyaluronate|Hyaluronate
C0551230|T201|COMP|13174-8|LNC|Interpretation|Interpretation
C0551231|T201|COMP|13169-8|LNC|Interpretation|Interpretation
C0551232|T201|COMP|13440-3|LNC|Interpretation|Interpretation
C0551233|T201|COMP|12801-7|LNC|Methdilazine|Methdilazine
C0551234|T201|COMP|12491-7|LNC|Methohexital|Methohexital
C0551235|T201|COMP|12316-6|LNC|Methopyrilene|Methopyrilene
C0551236|T201|COMP|12714-2|LNC|N-methylhistamine|N-methylhistamine
C0551237|T201|COMP|13311-6|LNC|MNSs group Ag|MNSs group Ag
C0551238|T201|COMP|13461-9|LNC|Monoacetyldapsone/Dapsone|Monoacetyldapsone/Dapsone
C0551239|T201|COMP|12919-7|LNC|Monoamine oxidase|Monoamine oxidase
C0551240|T201|COMP|12918-9|LNC|Monoamine oxidase|Monoamine oxidase
C0551241|T201|COMP|13348-8|LNC|Monoclonal band observed|Monoclonal band observed
C0551242|T201|COMP|13130-0|LNC|Motilin|Motilin
C0551243|T201|COMP|12542-7|LNC|N-methylacetamide|N-methylacetamide
C0551244|T201|COMP|12543-5|LNC|Methyl formamide|Methyl formamide
C0551245|T201|COMP|12405-7|LNC|Nabumetone|Nabumetone
C0551246|T201|COMP|12435-4|LNC|Naphthalene|Naphthalene
C0551247|T201|COMP|12436-2|LNC|Naphthol|Naphthol
C0551248|T201|COMP|13016-1|LNC|Nitrophenol|Nitrophenol
C0551249|T201|COMP|13026-0|LNC|Orthocresol|Orthocresol
C0551250|T201|COMP|13477-5|LNC|Orthocresol/Creatinine|Orthocresol/Creatinine
C0551251|T201|COMP|12408-1|LNC|Oxybutynin|Oxybutynin
C0551252|T201|COMP|12994-0|LNC|Oxychlordane|Oxychlordane
C0551253|T201|COMP|13006-2|LNC|1,4-Dichlorobenzene|1,4-Dichlorobenzene
C0551254|T201|COMP|11100-5|LNC|Tetrachloroethylene|Tetrachloroethylene
C0551255|T201|COMP|12331-5|LNC|Phenethylamine|Phenethylamine
C0551256|T201|COMP|12802-5|LNC|Propiomazine|Propiomazine
C0551257|T201|COMP|12412-3|LNC|Pyridine|Pyridine
C0551258|T201|COMP|12413-1|LNC|Resperine|Resperine
C0551259|T201|COMP|12414-9|LNC|Resperine|Resperine
C0551260|T201|COMP|12415-6|LNC|Selegiline|Selegiline
C0551261|T201|COMP|12429-7|LNC|Succinylcholine|Succinylcholine
C0551262|T201|COMP|12390-1|LNC|sulfaSALAzine|sulfaSALAzine
C0551263|T201|COMP|12417-2|LNC|Sulindac|Sulindac
C0551264|T201|COMP|12369-5|LNC|Sympathomimetics|Sympathomimetics
C0551265|T201|COMP|13357-9|LNC|Synovial cells|Synovial cells
C0551266|T201|COMP|12490-9|LNC|Allyl-sec-butyl-barbiturate|Allyl-sec-butyl-barbiturate
C0551267|T201|COMP|12492-5|LNC|Thiamylal|Thiamylal
C0551268|T201|COMP|12547-6|LNC|Phorate|Phorate
C0551269|T201|COMP|12441-2|LNC|Tolmetin|Tolmetin
C0551270|T201|COMP|12424-8|LNC|Triprolidine|Triprolidine
C0551271|T201|COMP|10861-3|LNC|Progesterone receptor|Progesterone receptor
C0551272|T201|COMP|13496-5|LNC|Triple phosphate crystals|Triple phosphate crystals
C0551273|T201|COMP|11560-0|LNC|Acetylcholine receptor binding Ab|Acetylcholine receptor binding Ab
C0551274|T201|COMP|11561-8|LNC|Acetylcholine receptor blocking Ab|Acetylcholine receptor blocking Ab
C0551275|T201|COMP|11562-6|LNC|Acetylcholine receptor modulation Ab|Acetylcholine receptor modulation Ab
C0551276|T201|COMP|10862-1|LNC|Basement membrane Ab|Basement membrane Ab
C0551277|T201|COMP|13110-2|LNC|Beta tubulin Ab.IgM|Beta tubulin Ab.IgM
C0551278|T201|COMP|12852-0|LNC|Bovine inner ear Ag|Bovine inner ear Ag
C0551279|T201|COMP|12724-1|LNC|Voltage-gated calcium channel Ab.IgG|Voltage-gated calcium channel Ab.IgG
C0551280|T201|COMP|12735-7|LNC|Collagen Ab|Collagen Ab
C0551281|T201|COMP|12734-0|LNC|Soluble liver Ab|Soluble liver Ab
C0551282|T201|COMP|13091-4|LNC|Deoxyribonucleoprotein Ab|Deoxyribonucleoprotein Ab
C0551283|T201|COMP|13107-8|LNC|Disialylganglioside GD1a Ab|Disialylganglioside GD1a Ab
C0551284|T201|COMP|13102-9|LNC|Disialylganglioside GD1b Ab|Disialylganglioside GD1b Ab
C0551285|T201|COMP|13103-7|LNC|Disialylganglioside GD1b Ab.IgG|Disialylganglioside GD1b Ab.IgG
C0551286|T201|COMP|13104-5|LNC|Disialylganglioside GD1b Ab.IgM|Disialylganglioside GD1b Ab.IgM
C0551287|T201|COMP|13308-2|LNC|DNA|DNA
C0551288|T201|COMP|11013-0|LNC|DNA double strand Ab|DNA double strand Ab
C0551290|T201|COMP|12277-0|LNC|DNA double strand Ab|DNA double strand Ab
C0551291|T201|COMP|13092-2|LNC|Endomysium Ab|Endomysium Ab
C0551292|T201|COMP|10863-9|LNC|Endomysium Ab.IgA|Endomysium Ab.IgA
C0551293|T201|COMP|13173-0|LNC|Fibronectin aggregate Ab.IgA|Fibronectin aggregate Ab.IgA
C0551294|T201|COMP|13089-8|LNC|Asialoganglioside GM1 Ab|Asialoganglioside GM1 Ab
C0551295|T201|COMP|13090-6|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C0551296|T201|COMP|12221-8|LNC|Heterophile Ab|Heterophile Ab
C0551297|T201|COMP|10864-7|LNC|Immune complex|Immune complex
C0551299|T201|COMP|13171-4|LNC|Immune complex|Immune complex
C0551300|T201|COMP|11087-4|LNC|Insulin Ab|Insulin Ab
C0551301|T201|COMP|10865-4|LNC|Intercellular substance Ab|Intercellular substance Ab
C0551302|T201|COMP|11564-2|LNC|Intrinsic factor Ab|Intrinsic factor Ab
C0551303|T201|COMP|11565-9|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C0551304|T201|COMP|13175-5|LNC|Liver cytosol Ab|Liver cytosol Ab
C0551305|T201|COMP|11566-7|LNC|Liver kidney microsomal Ab|Liver kidney microsomal Ab
C0551306|T201|COMP|13093-0|LNC|Monosialoganglioside GM1 Ab.IgM|Monosialoganglioside GM1 Ab.IgM
C0551307|T201|COMP|12776-1|LNC|Mucin-like carcinoma associated Ag|Mucin-like carcinoma associated Ag
C0551308|T201|COMP|13164-9|LNC|Human antimouse Ab|Human antimouse Ab
C0551309|T201|COMP|12897-5|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C0551310|T201|COMP|13119-3|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C0551311|T201|COMP|13118-5|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C0551312|T201|COMP|13096-3|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C0551313|T201|COMP|11089-0|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C0551314|T201|COMP|11088-2|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C0551315|T201|COMP|12854-6|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C0551316|T201|COMP|13115-1|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C0551317|T201|COMP|13114-4|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C0551318|T201|COMP|5128-4|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C0551319|T201|COMP|13066-6|LNC|Nuclear Ab|Nuclear Ab
C0551320|T201|COMP|13111-0|LNC|Nuclear Ab|Nuclear Ab
C0551321|T201|COMP|13112-8|LNC|Nuclear Ab|Nuclear Ab
C0551322|T201|COMP|13067-4|LNC|Nuclear Ab pattern|Nuclear Ab pattern
C0551323|T201|COMP|13068-2|LNC|Nuclear Ab pattern|Nuclear Ab pattern
C0551324|T201|COMP|13120-1|LNC|Ovary Ab|Ovary Ab
C0551325|T201|COMP|13129-2|LNC|Pancreatic oncofetal Ag|Pancreatic oncofetal Ag
C0551326|T201|COMP|12799-3|LNC|Parathyrin Ab|Parathyrin Ab
C0551327|T201|COMP|13072-4|LNC|Phosphatidate Ab.IgA|Phosphatidate Ab.IgA
C0551328|T201|COMP|13070-8|LNC|Phosphatidate Ab.IgG|Phosphatidate Ab.IgG
C0551329|T201|COMP|13071-6|LNC|Phosphatidate Ab.IgM|Phosphatidate Ab.IgM
C0551330|T201|COMP|13075-7|LNC|Phosphatidylcholine Ab.IgA|Phosphatidylcholine Ab.IgA
C0551331|T201|COMP|13073-2|LNC|Phosphatidylcholine Ab.IgG|Phosphatidylcholine Ab.IgG
C0551332|T201|COMP|13074-0|LNC|Phosphatidylcholine Ab.IgM|Phosphatidylcholine Ab.IgM
C0551333|T201|COMP|13078-1|LNC|Phosphatidylethanolamine Ab.IgA|Phosphatidylethanolamine Ab.IgA
C0551334|T201|COMP|13076-5|LNC|Phosphatidylethanolamine Ab.IgG|Phosphatidylethanolamine Ab.IgG
C0551335|T201|COMP|13077-3|LNC|Phosphatidylethanolamine Ab.IgM|Phosphatidylethanolamine Ab.IgM
C0551336|T201|COMP|13081-5|LNC|Phosphatidylglycerol Ab.IgA|Phosphatidylglycerol Ab.IgA
C0551337|T201|COMP|13079-9|LNC|Phosphatidylglycerol Ab.IgG|Phosphatidylglycerol Ab.IgG
C0551338|T201|COMP|13080-7|LNC|Phosphatidylglycerol Ab.IgM|Phosphatidylglycerol Ab.IgM
C0551339|T201|COMP|13084-9|LNC|Phosphatidylinositol Ab.IgA|Phosphatidylinositol Ab.IgA
C0551340|T201|COMP|13082-3|LNC|Phosphatidylinositol Ab.IgG|Phosphatidylinositol Ab.IgG
C0551341|T201|COMP|13083-1|LNC|Phosphatidylinositol Ab.IgM|Phosphatidylinositol Ab.IgM
C0551342|T201|COMP|13069-0|LNC|Phosphatidylserine Ab.IgA|Phosphatidylserine Ab.IgA
C0551343|T201|COMP|11568-3|LNC|Phosphatidylserine Ab.IgG|Phosphatidylserine Ab.IgG
C0551344|T201|COMP|11569-1|LNC|Phosphatidylserine Ab.IgM|Phosphatidylserine Ab.IgM
C0551345|T201|COMP|13065-8|LNC|Platelet Ab.circulating|Platelet Ab.circulating
C0551346|T201|COMP|13063-3|LNC|Drug induced platelet Ab|Drug induced platelet Ab
C0551347|T201|COMP|13062-5|LNC|Platelet Ab.IgA|Platelet Ab.IgA
C0551348|T201|COMP|11570-9|LNC|Platelet Ab.IgG|Platelet Ab.IgG
C0551349|T201|COMP|13061-7|LNC|Platelet Ab.IgM|Platelet Ab.IgM
C0551350|T201|COMP|13064-1|LNC|Platelet associated Ab.IgA|Platelet associated Ab.IgA
C0551351|T201|COMP|13097-1|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C0551352|T201|COMP|12853-8|LNC|Purkinje cells Ab|Purkinje cells Ab
C0551353|T201|COMP|13116-9|LNC|Reticulin Ab.IgG|Reticulin Ab.IgG
C0551354|T201|COMP|11571-7|LNC|Rheumatoid arthritis nuclear Ab|Rheumatoid arthritis nuclear Ab
C0551356|T201|COMP|11572-5|LNC|Rheumatoid factor|Rheumatoid factor
C0551357|T201|COMP|11573-3|LNC|Rheumatoid factor.IgM|Rheumatoid factor.IgM
C0551358|T201|COMP|13121-9|LNC|Ribosomal P protein Ab|Ribosomal P protein Ab
C0551359|T201|COMP|13347-0|LNC|RNA polymerase I+II+III Ab|RNA polymerase I+II+III Ab
C0551360|T201|COMP|11090-8|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0551361|T201|COMP|11014-8|LNC|Somatotropin Ab|Somatotropin Ab
C0551362|T201|COMP|11015-5|LNC|Somatotropin binding protein|Somatotropin binding protein
C0551363|T201|COMP|10866-2|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C0551364|T201|COMP|13098-9|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C0551365|T201|COMP|10867-0|LNC|Sulfatide Ab.IgM|Sulfatide Ab.IgM
C0551366|T201|COMP|13106-0|LNC|Tetrasialylganglioside GQ1b Ab|Tetrasialylganglioside GQ1b Ab
C0551367|T201|COMP|13105-2|LNC|Tetrasialylganglioside GQ1b Ab.IgG|Tetrasialylganglioside GQ1b Ab.IgG
C0551368|T201|COMP|8099-4|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C0551375|T201|COMP|12984-1|LNC|2,4 toluenediamine|2,4 toluenediamine
C0551376|T201|COMP|12985-8|LNC|2,6 toluenediamine|2,6 toluenediamine
C0551377|T201|COMP|12989-0|LNC|Allyl alcohol|Allyl alcohol
C0551378|T201|COMP|11091-6|LNC|Alpha chlordane|Alpha chlordane
C0551379|T201|COMP|13470-0|LNC|Aluminum/Creatinine|Aluminum/Creatinine
C0551380|T201|COMP|12535-1|LNC|Amyl nitrite|Amyl nitrite
C0551381|T201|COMP|12702-7|LNC|Antimony|Antimony
C0551382|T201|COMP|12481-8|LNC|Arsenic.inorganic|Arsenic.inorganic
C0551383|T201|COMP|13463-5|LNC|Arsenic/Creatinine|Arsenic/Creatinine
C0551384|T201|COMP|11092-4|LNC|Barbiturates|Barbiturates
C0551385|T201|COMP|11022-1|LNC|Barbiturates|Barbiturates
C0551386|T201|COMP|12358-8|LNC|Barbiturates|Barbiturates
C0551387|T201|COMP|10909-0|LNC|Benzidine|Benzidine
C0551388|T201|COMP|12364-6|LNC|Benzodiazepines|Benzodiazepines
C0551389|T201|COMP|11023-9|LNC|Benzodiazepines|Benzodiazepines
C0551390|T201|COMP|11024-7|LNC|Benzodiazepines|Benzodiazepines
C0551391|T201|COMP|12359-6|LNC|Benzodiazepines|Benzodiazepines
C0551392|T201|COMP|12304-2|LNC|Benzyl alcohol|Benzyl alcohol
C0551393|T201|COMP|10910-8|LNC|Borate|Borate
C0551394|T201|COMP|12433-9|LNC|Bufotenine|Bufotenine
C0551395|T201|COMP|12536-9|LNC|Butyl nitrate|Butyl nitrate
C0551396|T201|COMP|12505-4|LNC|Cadmium|Cadmium
C0551397|T201|COMP|13471-8|LNC|Cadmium/Creatinine|Cadmium/Creatinine
C0551398|T201|COMP|13478-3|LNC|Tetrahydrocannabinol/Creatinine|Tetrahydrocannabinol/Creatinine
C0551399|T201|COMP|12351-3|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0551400|T201|COMP|12297-8|LNC|Chlorate|Chlorate
C0551401|T201|COMP|12993-2|LNC|Hydrocarbons.chlorinated|Hydrocarbons.chlorinated
C0551402|T201|COMP|13464-3|LNC|Chromium/Creatinine|Chromium/Creatinine
C0551403|T201|COMP|13468-4|LNC|Cobalt/Creatinine|Cobalt/Creatinine
C0551404|T201|COMP|12556-7|LNC|Copper|Copper
C0551405|T201|COMP|12293-7|LNC|Cotinine|Cotinine
C0551406|T201|COMP|13497-3|LNC|Dextroamphetamine/Levoamphetamine|Dextroamphetamine/Levoamphetamine
C0551408|T201|COMP|13498-1|LNC|Dextromethamphetamine/Levomethamphetamine|Dextromethamphetamine/Levomethamphetamine
C0551409|T201|COMP|10911-6|LNC|Dichlorobenzidine|Dichlorobenzidine
C0551410|T201|COMP|12996-5|LNC|Dichlorodifluoroethane|Dichlorodifluoroethane
C0551411|T201|COMP|11093-2|LNC|Dichlorodiphenyldichloroethylene|Dichlorodiphenyldichloroethylene
C0551412|T201|COMP|11094-0|LNC|Dichlorodiphenyltrichloroethane|Dichlorodiphenyltrichloroethane
C0551413|T201|COMP|12307-5|LNC|Dichloroethane|Dichloroethane
C0551414|T201|COMP|12998-1|LNC|Methylene chloride|Methylene chloride
C0551415|T201|COMP|11095-7|LNC|Dieldrin|Dieldrin
C0551416|T201|COMP|13015-3|LNC|Diisobutylketone|Diisobutylketone
C0551417|T201|COMP|12287-9|LNC|Drugs identified|Drugs identified
C0551418|T201|COMP|12289-5|LNC|Drugs identified|Drugs identified
C0551419|T201|COMP|13007-0|LNC|Ethane|Ethane
C0551420|T201|COMP|12465-1|LNC|Ethanol|Ethanol
C0551421|T201|COMP|13027-8|LNC|Ethyl acetate|Ethyl acetate
C0551422|T201|COMP|12340-6|LNC|Ethylene|Ethylene
C0551423|T201|COMP|12601-1|LNC|Fluoride|Fluoride
C0551424|T201|COMP|13475-9|LNC|Fluoride/Creatinine|Fluoride/Creatinine
C0551425|T201|COMP|12703-5|LNC|Gallium|Gallium
C0551426|T201|COMP|11096-5|LNC|Gamma chlordane|Gamma chlordane
C0551427|T201|COMP|12295-2|LNC|Hallucinogens|Hallucinogens
C0551428|T201|COMP|13005-4|LNC|2,4,5-Trichlorophenoxyacetate|2,4,5-Trichlorophenoxyacetate
C0551429|T201|COMP|13003-9|LNC|Hydrocarbons.halogenated|Hydrocarbons.halogenated
C0551430|T201|COMP|12446-1|LNC|Hydrocarbons.halogenated|Hydrocarbons.halogenated
C0551431|T201|COMP|13004-7|LNC|Hydrocarbons.halogenated.volatile|Hydrocarbons.halogenated.volatile
C0551432|T201|COMP|12992-4|LNC|Isobutane|Isobutane
C0551433|T201|COMP|12371-1|LNC|Isopropyl ether|Isopropyl ether
C0551434|T201|COMP|12478-4|LNC|Levomethamphetamine|Levomethamphetamine
C0551435|T201|COMP|10912-4|LNC|Lead|Lead
C0551436|T201|COMP|12770-4|LNC|Lead|Lead
C0551437|T201|COMP|13466-8|LNC|Lead/Creatinine|Lead/Creatinine
C0551438|T201|COMP|12704-3|LNC|Length|Length
C0551439|T201|COMP|11097-3|LNC|Lindane|Lindane
C0551440|T201|COMP|11098-1|LNC|Malaoxon|Malaoxon
C0551441|T201|COMP|12775-3|LNC|Mercury|Mercury
C0551442|T201|COMP|12774-6|LNC|Mercury|Mercury
C0551443|T201|COMP|13465-0|LNC|Mercury/Creatinine|Mercury/Creatinine
C0551444|T201|COMP|12296-0|LNC|Mescaline|Mescaline
C0551445|T201|COMP|13002-1|LNC|Mesityl oxide|Mesityl oxide
C0551446|T201|COMP|11025-4|LNC|Methadone|Methadone
C0551447|T201|COMP|11026-2|LNC|Methaqualone|Methaqualone
C0551448|T201|COMP|11099-9|LNC|Methoxychlor|Methoxychlor
C0551449|T201|COMP|13011-2|LNC|Methyl ethyl ketone|Methyl ethyl ketone
C0551450|T201|COMP|13009-6|LNC|Methyl ethyl ketone|Methyl ethyl ketone
C0551451|T201|COMP|13012-0|LNC|Methyl isoamyl ketone|Methyl isoamyl ketone
C0551452|T201|COMP|13013-8|LNC|Methyl isobutyl ketone|Methyl isobutyl ketone
C0551453|T201|COMP|13010-4|LNC|Methyl amyl ketone|Methyl amyl ketone
C0551454|T201|COMP|13014-6|LNC|Methyl butyl ketone|Methyl butyl ketone
C0551455|T201|COMP|13008-8|LNC|Methyl propyl ketone|Methyl propyl ketone
C0551456|T201|COMP|10913-2|LNC|4,4'-Methylene bis(2-Chloroaniline)|4,4'-Methylene bis(2-Chloroaniline)
C0551457|T201|COMP|10914-0|LNC|Methylenediamine|Methylenediamine
C0551458|T201|COMP|12554-2|LNC|Narcotics|Narcotics
C0551459|T201|COMP|12780-3|LNC|Nickel|Nickel
C0551460|T201|COMP|12779-5|LNC|Nickel|Nickel
C0551461|T201|COMP|13472-6|LNC|Nickel/Creatinine|Nickel/Creatinine
C0551462|T201|COMP|12538-5|LNC|Nitrate|Nitrate
C0551463|T201|COMP|12354-7|LNC|Opiates|Opiates
C0551464|T201|COMP|12338-0|LNC|Pentachlorophenol|Pentachlorophenol
C0551465|T201|COMP|13020-3|LNC|Pesticides|Pesticides
C0551466|T201|COMP|13021-1|LNC|Pesticides|Pesticides
C0551467|T201|COMP|13019-5|LNC|Pesticides|Pesticides
C0551468|T201|COMP|13018-7|LNC|Pesticides|Pesticides
C0551469|T201|COMP|12355-4|LNC|Phencyclidine|Phencyclidine
C0551470|T201|COMP|10915-7|LNC|Phencyclidine|Phencyclidine
C0551471|T201|COMP|10916-5|LNC|Platinum|Platinum
C0551472|T201|COMP|12991-6|LNC|Polychlorinated biphenyl.Aroclor 1254|Polychlorinated biphenyl.Aroclor 1254
C0551473|T201|COMP|12990-8|LNC|Polychlorinated biphenyl.Aroclor 1260|Polychlorinated biphenyl.Aroclor 1260
C0551474|T201|COMP|13022-9|LNC|Propane|Propane
C0551475|T201|COMP|11027-0|LNC|Propoxyphene|Propoxyphene
C0551476|T201|COMP|12552-6|LNC|Propylene glycol|Propylene glycol
C0551477|T201|COMP|13467-6|LNC|Selenium/Creatinine|Selenium/Creatinine
C0551478|T201|COMP|13476-7|LNC|Silver/Creatinine|Silver/Creatinine
C0551479|T201|COMP|12553-4|LNC|Stimulants|Stimulants
C0551480|T201|COMP|12705-0|LNC|Strontium|Strontium
C0551481|T201|COMP|12706-8|LNC|Tellurium|Tellurium
C0551482|T201|COMP|13469-2|LNC|Thallium/Creatinine|Thallium/Creatinine
C0551483|T201|COMP|12343-0|LNC|Thiazides|Thiazides
C0551484|T201|COMP|12707-6|LNC|Thorium|Thorium
C0551485|T201|COMP|12708-4|LNC|Tin|Tin
C0551486|T201|COMP|13024-5|LNC|Trichlorofluoroethane|Trichlorofluoroethane
C0551487|T201|COMP|13023-7|LNC|Trichlorofluoromethane|Trichlorofluoromethane
C0551488|T201|COMP|13025-2|LNC|Trichlorotrifluoroethane|Trichlorotrifluoroethane
C0551489|T201|COMP|12483-4|LNC|Tungsten|Tungsten
C0551490|T201|COMP|12549-2|LNC|Turpentine|Turpentine
C0551491|T201|COMP|12555-9|LNC|Turpentine|Turpentine
C0551492|T201|COMP|12983-3|LNC|Volatiles|Volatiles
C0551493|T201|COMP|11028-8|LNC|Zinc|Zinc
C0551494|T201|COMP|10917-3|LNC|Zinc|Zinc
C0551495|T201|COMP|10918-1|LNC|Zinc|Zinc
C0551496|T201|COMP|13473-4|LNC|Zinc/Creatinine|Zinc/Creatinine
C0551497|T201|COMP|11218-5|LNC|Albumin|Albumin
C0551498|T201|COMP|12453-7|LNC|Phosphate crystals.amorphous|Phosphate crystals.amorphous
C0551499|T201|COMP|12454-5|LNC|Urate crystals.amorphous|Urate crystals.amorphous
C0551500|T201|COMP|11101-3|LNC|Bacteria|Bacteria
C0551501|T201|COMP|11278-9|LNC|Bladder cells|Bladder cells
C0551502|T201|COMP|12512-0|LNC|Calcium hydrogen phosphate dihydrate crystals|Calcium hydrogen phosphate dihydrate crystals
C0551503|T201|COMP|11029-6|LNC|Consistency|Consistency
C0551504|T201|COMP|12469-3|LNC|Cystine crystals|Cystine crystals
C0551505|T201|COMP|12210-1|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0551506|T201|COMP|11277-1|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C0551507|T201|COMP|11279-7|LNC|Urine sediment comments|Urine sediment comments
C0552286|T201|COMP|13495-7|LNC|Specimen volume|Specimen volume
C0552287|T201|COMP|13494-0|LNC|Specimen volume|Specimen volume
C0552288|T201|COMP|12457-8|LNC|Specimen volume|Specimen volume
C0552289|T201|COMP|12254-9|LNC|Specimen volume|Specimen volume
C0552290|T201|COMP|12255-6|LNC|Specimen volume|Specimen volume
C0678220|T201|COMP|13099-7|LNC|Sulfatide Ab.IgM|Sulfatide Ab.IgM
C0699860|T201|COMP|10878-7|LNC|Iodine.protein bound|Iodine.protein bound
C0700435|T201|COMP|1196-5|LNC|Little NOS Ab|Little NOS Ab
C0700436|T201|COMP|1544-6|LNC|Glucose^6H post 100 g glucose PO|Glucose^6H post 100 g glucose PO
C0796701|T201|COMP|13507-9|LNC|Lupus erythematosus cells|Lupus erythematosus cells
C0796702|T201|COMP|13508-7|LNC|Hematocrit|Hematocrit
C0796705|T201|COMP|13511-1|LNC|Cyanide ascorbate screen|Cyanide ascorbate screen
C0796707|T201|COMP|13513-7|LNC|Iron.microscopic observation|Iron.microscopic observation
C0796708|T201|COMP|13514-5|LNC|Hemoglobin pattern|Hemoglobin pattern
C0796709|T201|COMP|13515-2|LNC|Hemoglobin pattern|Hemoglobin pattern
C0796710|T201|COMP|13516-0|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0796711|T201|COMP|13517-8|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C0796712|T201|COMP|13518-6|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C0796713|T201|COMP|13519-4|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0796714|T201|COMP|13521-0|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C0796715|T201|COMP|13522-8|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C0796716|T201|COMP|13523-6|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0796717|T201|COMP|13524-4|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0796718|T201|COMP|13525-1|LNC|Nonhematic cells/100 leukocytes|Nonhematic cells/100 leukocytes
C0796719|T201|COMP|13526-9|LNC|Nonhematic cells/100 leukocytes|Nonhematic cells/100 leukocytes
C0796720|T201|COMP|13527-7|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C0796721|T201|COMP|13528-5|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C0796722|T201|COMP|13529-3|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C0796723|T201|COMP|13530-1|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C0796724|T201|COMP|13531-9|LNC|Fat.microscopic observation|Fat.microscopic observation
C0796725|T201|COMP|13532-7|LNC|Xanthochromia|Xanthochromia
C0796726|T201|COMP|13533-5|LNC|Acid hemolysis|Acid hemolysis
C0796727|T201|COMP|13534-3|LNC|Sucrose hemolysis|Sucrose hemolysis
C0796728|T201|COMP|13535-0|LNC|Sucrose hemolysis|Sucrose hemolysis
C0796729|T201|COMP|13536-8|LNC|Globulin|Globulin
C0796730|T201|COMP|13537-6|LNC|Protein|Protein
C0796730|T201|COMP|14897-3|LNC|Protein|Protein
C0796731|T201|COMP|13538-4|LNC|Carbon dioxide|Carbon dioxide
C0796732|T201|COMP|13539-2|LNC|Phosphate|Phosphate
C0796733|T201|COMP|13540-0|LNC|Carbon dioxide|Carbon dioxide
C0796734|T201|COMP|13542-6|LNC|Phosphate|Phosphate
C0796735|T201|COMP|13544-2|LNC|4-Hydroxyglutethimide|4-Hydroxyglutethimide
C0796736|T201|COMP|13545-9|LNC|ALPRAZolam|ALPRAZolam
C0796737|T201|COMP|13546-7|LNC|Amikacin|Amikacin
C0796738|T201|COMP|13547-5|LNC|Butriptyline|Butriptyline
C0796739|T201|COMP|13548-3|LNC|chlorproMAZINE|chlorproMAZINE
C0796740|T201|COMP|13549-1|LNC|clomiPRAMINE|clomiPRAMINE
C0796741|T201|COMP|13550-9|LNC|clonazePAM|clonazePAM
C0796742|T201|COMP|13551-7|LNC|Clorazepate|Clorazepate
C0796743|T201|COMP|13552-5|LNC|cloZAPine|cloZAPine
C0796744|T201|COMP|13553-3|LNC|Cocaethylene|Cocaethylene
C0796745|T201|COMP|13554-1|LNC|Cyclobenzaprine|Cyclobenzaprine
C0796746|T201|COMP|13555-8|LNC|D-pseudoephedrine|D-pseudoephedrine
C0796747|T201|COMP|13556-6|LNC|Demoxepam|Demoxepam
C0796748|T201|COMP|13557-4|LNC|Norsertraline|Norsertraline
C0796749|T201|COMP|13558-2|LNC|Disopyramide|Disopyramide
C0796750|T201|COMP|13559-0|LNC|Flecainide|Flecainide
C0796751|T201|COMP|13560-8|LNC|fluvoxaMINE|fluvoxaMINE
C0796752|T201|COMP|13561-6|LNC|Gentamicin|Gentamicin
C0796753|T201|COMP|13562-4|LNC|Gentamicin|Gentamicin
C0796754|T201|COMP|13563-2|LNC|Glutethimide|Glutethimide
C0796755|T201|COMP|13564-0|LNC|Ibuprofen|Ibuprofen
C0796756|T201|COMP|13565-7|LNC|LORazepam|LORazepam
C0796757|T201|COMP|13566-5|LNC|Mesoridazine|Mesoridazine
C0796758|T201|COMP|13567-3|LNC|Mexiletine|Mexiletine
C0796759|T201|COMP|13568-1|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0796760|T201|COMP|13569-9|LNC|Norchlordiazepoxide|Norchlordiazepoxide
C0796761|T201|COMP|13570-7|LNC|Norclomipramine|Norclomipramine
C0796762|T201|COMP|13571-5|LNC|Norclozapine|Norclozapine
C0796763|T201|COMP|13572-3|LNC|Nordiazepam|Nordiazepam
C0796764|T201|COMP|13573-1|LNC|Nordoxepin|Nordoxepin
C0796765|T201|COMP|13574-9|LNC|Norfluoxetine|Norfluoxetine
C0796766|T201|COMP|13575-6|LNC|Normaprotiline|Normaprotiline
C0796767|T201|COMP|13576-4|LNC|oxyCODONE|oxyCODONE
C0796768|T201|COMP|13577-2|LNC|PARoxetine|PARoxetine
C0796769|T201|COMP|13578-0|LNC|Promazine|Promazine
C0796770|T201|COMP|13579-8|LNC|Sertraline|Sertraline
C0796771|T201|COMP|13580-6|LNC|Temazepam|Temazepam
C0796772|T201|COMP|13581-4|LNC|Theophylline|Theophylline
C0796773|T201|COMP|13582-2|LNC|Theophylline|Theophylline
C0796774|T201|COMP|13583-0|LNC|Thioridazine|Thioridazine
C0796775|T201|COMP|13584-8|LNC|Tobramycin|Tobramycin
C0796776|T201|COMP|13585-5|LNC|Trifluoperazine|Trifluoperazine
C0796777|T201|COMP|13586-3|LNC|Vancomycin|Vancomycin
C0796778|T201|COMP|13587-1|LNC|Vancomycin|Vancomycin
C0796779|T201|COMP|13588-9|LNC|Venlafaxine|Venlafaxine
C0796780|T201|COMP|13589-7|LNC|Activated protein C resistance|Activated protein C resistance
C0796781|T201|COMP|13590-5|LNC|Activated protein C resistance|Activated protein C resistance
C0796782|T201|COMP|13591-3|LNC|Factor inhibitor XXX|Factor inhibitor XXX
C0796783|T201|COMP|13592-1|LNC|Platelet aggregation.XXX induced|Platelet aggregation.XXX induced
C0796784|T201|COMP|13593-9|LNC|Platelet aggregation.prostaglandin induced|Platelet aggregation.prostaglandin induced
C0796785|T201|COMP|13594-7|LNC|Prekallikrein|Prekallikrein
C0796786|T201|COMP|13595-4|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0796787|T201|COMP|13596-2|LNC|Histiocytes|Histiocytes
C0796788|T201|COMP|13597-0|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0796789|T201|COMP|783-1|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C0796790|T201|COMP|33855-8|LNC|Promonocytes|Promonocytes
C0796791|T201|COMP|13600-2|LNC|11-Deoxycortisol^15M post 250 ug corticotropin|11-Deoxycortisol^15M post 250 ug corticotropin
C0796792|T201|COMP|13601-0|LNC|11-Deoxycortisol^1H post 250 ug corticotropin|11-Deoxycortisol^1H post 250 ug corticotropin
C0796793|T201|COMP|13602-8|LNC|11-Deoxycortisol^30M post 250 ug corticotropin|11-Deoxycortisol^30M post 250 ug corticotropin
C0796797|T201|COMP|13606-9|LNC|Glucose^3H post 50 g lactose PO|Glucose^3H post 50 g lactose PO
C0796798|T201|COMP|13607-7|LNC|Glucose^4H post 50 g lactose PO|Glucose^4H post 50 g lactose PO
C0796799|T201|COMP|13608-5|LNC|Insulin^1.5H post 75 g glucose PO|Insulin^1.5H post 75 g glucose PO
C0796800|T201|COMP|13609-3|LNC|Insulin^2.5H post 75 g glucose PO|Insulin^2.5H post 75 g glucose PO
C0796801|T201|COMP|13610-1|LNC|3-Beta-Androstanediol|3-Beta-Androstanediol
C0796802|T201|COMP|13611-9|LNC|6-Beta-Hydroxycortisol|6-Beta-Hydroxycortisol
C0796803|T201|COMP|13612-7|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C0796804|T201|COMP|13613-5|LNC|Ethanolamine|Ethanolamine
C0796805|T201|COMP|13614-3|LNC|Etiocholanolone|Etiocholanolone
C0796806|T201|COMP|13615-0|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0796807|T201|COMP|13616-8|LNC|Nitrite|Nitrite
C0796808|T201|COMP|13617-6|LNC|Prostaglandin D2|Prostaglandin D2
C0796809|T201|COMP|13618-4|LNC|Tetrahydroaldosterone|Tetrahydroaldosterone
C0796810|T201|COMP|13619-2|LNC|Specimen volume|Specimen volume
C0796811|T201|COMP|13620-0|LNC|Specimen volume|Specimen volume
C0796812|T201|COMP|13621-8|LNC|Coagulation thrombin induced|Coagulation thrombin induced
C0796813|T201|COMP|13622-6|LNC|Acetaminophen|Acetaminophen
C0796814|T201|COMP|13623-4|LNC|Dextromethorphan|Dextromethorphan
C0796815|T201|COMP|13624-2|LNC|DOXOrubicin|DOXOrubicin
C0796816|T201|COMP|13625-9|LNC|Methoxsalen|Methoxsalen
C0796817|T201|COMP|13626-7|LNC|Mitotane|Mitotane
C0796818|T201|COMP|13627-5|LNC|Erythrocytes|Erythrocytes
C0796820|T201|COMP|13629-1|LNC|Interleukin 1 beta|Interleukin 1 beta
C0796821|T201|COMP|13170-6|LNC|Immune complex|Immune complex
C0796822|T201|COMP|13631-7|LNC|Immune complex|Immune complex
C0796823|T201|COMP|13632-5|LNC|Insulin receptor Ab|Insulin receptor Ab
C0796824|T201|COMP|13633-3|LNC|Insulin receptor Ab|Insulin receptor Ab
C0796825|T201|COMP|13634-1|LNC|Rheumatoid factor|Rheumatoid factor
C0796826|T201|COMP|13635-8|LNC|Ribosomal Ab|Ribosomal Ab
C0796827|T201|COMP|13636-6|LNC|Ribosomal P Ab|Ribosomal P Ab
C0796828|T201|COMP|13637-4|LNC|Trichloroethane|Trichloroethane
C0796829|T201|COMP|13638-2|LNC|Chlordecone|Chlordecone
C0796830|T201|COMP|13639-0|LNC|Chlordecone|Chlordecone
C0796831|T201|COMP|13640-8|LNC|Vinyl chloride|Vinyl chloride
C0796832|T201|COMP|13641-6|LNC|Codeine|Codeine
C0796833|T201|COMP|13642-4|LNC|Ethylene glycol|Ethylene glycol
C0796834|T201|COMP|13643-2|LNC|Lindane|Lindane
C0796835|T201|COMP|13644-0|LNC|1,3-Dimethylbenzene|1,3-Dimethylbenzene
C0796836|T201|COMP|13645-7|LNC|Manganese|Manganese
C0796837|T201|COMP|13646-5|LNC|Methaqualone|Methaqualone
C0796839|T201|COMP|13648-1|LNC|Morphine|Morphine
C0796840|T201|COMP|13649-9|LNC|Nickel|Nickel
C0796841|T201|COMP|13650-7|LNC|1,2-Dimethylbenzene|1,2-Dimethylbenzene
C0796842|T201|COMP|13651-5|LNC|1,4-Dimethylbenzene|1,4-Dimethylbenzene
C0796843|T201|COMP|13652-3|LNC|Zinc|Zinc
C0796844|T201|COMP|13653-1|LNC|Epithelial cells.renal|Epithelial cells.renal
C0796845|T201|COMP|13654-9|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C0796846|T201|COMP|13655-6|LNC|Leukocytes|Leukocytes
C0796847|T201|COMP|13656-4|LNC|Phosphate crystals.amorphous|Phosphate crystals.amorphous
C0796848|T201|COMP|13657-2|LNC|Urate crystals.amorphous|Urate crystals.amorphous
C0796849|T201|COMP|13658-0|LNC|Urobilinogen|Urobilinogen
C0796850|T201|COMP|13659-8|LNC|Epidermal growth factor receptor|Epidermal growth factor receptor
C0796851|T201|COMP|13660-6|LNC|Gonadotropin releasing hormone|Gonadotropin releasing hormone
C0796852|T201|COMP|13661-4|LNC|Ganglioside GD1b Ab.IgM|Ganglioside GD1b Ab.IgM
C0796853|T201|COMP|13662-2|LNC|Ganglioside GD1b Ab.IgG|Ganglioside GD1b Ab.IgG
C0796854|T201|COMP|13663-0|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C0796856|T201|COMP|13665-5|LNC|1-Methylhistidine/Creatinine|1-Methylhistidine/Creatinine
C0796857|T201|COMP|13666-3|LNC|Alpha aminoadipate/Creatinine|Alpha aminoadipate/Creatinine
C0796858|T201|COMP|13667-1|LNC|Alpha aminobutyrate/Creatinine|Alpha aminobutyrate/Creatinine
C0796859|T201|COMP|13668-9|LNC|2-Ethyl-3-Hydroxypropionate/Creatinine|2-Ethyl-3-Hydroxypropionate/Creatinine
C0796860|T201|COMP|13669-7|LNC|2-Hydroxy-3-Methylvalerate/Creatinine|2-Hydroxy-3-Methylvalerate/Creatinine
C0796861|T201|COMP|13670-5|LNC|2-Hydroxyadipate/Creatinine|2-Hydroxyadipate/Creatinine
C0796862|T201|COMP|13671-3|LNC|Alpha hydroxybutyrate/Creatinine|Alpha hydroxybutyrate/Creatinine
C0796863|T201|COMP|13672-1|LNC|2-Hydroxyglutarate/Creatinine|2-Hydroxyglutarate/Creatinine
C0796864|T201|COMP|13673-9|LNC|2-Hydroxyisocaproate/Creatinine|2-Hydroxyisocaproate/Creatinine
C0796865|T201|COMP|13674-7|LNC|2-Hydroxyisovalerate/Creatinine|2-Hydroxyisovalerate/Creatinine
C0796866|T201|COMP|13675-4|LNC|2-Methyl-3-Hydroxybutyrate/Creatinine|2-Methyl-3-Hydroxybutyrate/Creatinine
C0796867|T201|COMP|13676-2|LNC|2-Oxo,3-Methylvalerate/Creatinine|2-Oxo,3-Methylvalerate/Creatinine
C0796868|T201|COMP|13677-0|LNC|2-Oxoadipate/Creatinine|2-Oxoadipate/Creatinine
C0796869|T201|COMP|13678-8|LNC|Alpha ketoglutarate/Creatinine|Alpha ketoglutarate/Creatinine
C0796870|T201|COMP|13679-6|LNC|2-Oxoisocaproate/Creatinine|2-Oxoisocaproate/Creatinine
C0796871|T201|COMP|13680-4|LNC|2-Oxoisovalerate/Creatinine|2-Oxoisovalerate/Creatinine
C0796872|T201|COMP|13681-2|LNC|Beta aminoisobutyrate/Creatinine|Beta aminoisobutyrate/Creatinine
C0796873|T201|COMP|13682-0|LNC|3-Hydroxy,3-Methylglutarate/Creatinine|3-Hydroxy,3-Methylglutarate/Creatinine
C0796874|T201|COMP|13683-8|LNC|3-Hydroxyadipate/Creatinine|3-Hydroxyadipate/Creatinine
C0796875|T201|COMP|13684-6|LNC|Beta hydroxybutyrate/Creatinine|Beta hydroxybutyrate/Creatinine
C0796876|T201|COMP|13685-3|LNC|3-Hydroxyglutarate/Creatinine|3-Hydroxyglutarate/Creatinine
C0796877|T201|COMP|13686-1|LNC|3-Hydroxyisobutyrate/Creatinine|3-Hydroxyisobutyrate/Creatinine
C0796878|T201|COMP|13687-9|LNC|3-Hydroxyisovalerate/Creatinine|3-Hydroxyisovalerate/Creatinine
C0796879|T201|COMP|13688-7|LNC|3-Hydroxypropionate/Creatinine|3-Hydroxypropionate/Creatinine
C0796880|T201|COMP|13689-5|LNC|3-Hydroxyvalerate/Creatinine|3-Hydroxyvalerate/Creatinine
C0796881|T201|COMP|13690-3|LNC|Vanillylmandelate/Creatinine|Vanillylmandelate/Creatinine
C0796882|T201|COMP|13691-1|LNC|3-Methylcrotonylglycine/Creatinine|3-Methylcrotonylglycine/Creatinine
C0796883|T201|COMP|13692-9|LNC|3-Methylglutaconate/Creatinine|3-Methylglutaconate/Creatinine
C0796884|T201|COMP|13693-7|LNC|3-Methylglutarate/Creatinine|3-Methylglutarate/Creatinine
C0796885|T201|COMP|13694-5|LNC|3-Methylhistidine/Creatinine|3-Methylhistidine/Creatinine
C0796886|T201|COMP|13695-2|LNC|Gamma aminobutyrate/Creatinine|Gamma aminobutyrate/Creatinine
C0796887|T201|COMP|13696-0|LNC|4-Hydroxyphenylacetate/Creatinine|4-Hydroxyphenylacetate/Creatinine
C0796888|T201|COMP|13697-8|LNC|4-Hydroxyphenyllactate/Creatinine|4-Hydroxyphenyllactate/Creatinine
C0796889|T201|COMP|13698-6|LNC|4-Hydroxyphenylpyruvate/Creatinine|4-Hydroxyphenylpyruvate/Creatinine
C0796890|T201|COMP|13699-4|LNC|5-Hydroxyhexanoate/Creatinine|5-Hydroxyhexanoate/Creatinine
C0796891|T201|COMP|13700-0|LNC|5-Oxoproline/Creatinine|5-Oxoproline/Creatinine
C0796892|T201|COMP|13701-8|LNC|Acetoacetate/Creatinine|Acetoacetate/Creatinine
C0796893|T201|COMP|13702-6|LNC|Aconitate/Creatinine|Aconitate/Creatinine
C0796894|T201|COMP|13703-4|LNC|Adipate/Creatinine|Adipate/Creatinine
C0796895|T201|COMP|13704-2|LNC|Alanine/Creatinine|Alanine/Creatinine
C0796896|T201|COMP|13705-9|LNC|Albumin/Creatinine|Albumin/Creatinine
C0796897|T201|COMP|13706-7|LNC|Amylase/Creatinine|Amylase/Creatinine
C0796898|T201|COMP|13707-5|LNC|Anserine/Creatinine|Anserine/Creatinine
C0796899|T201|COMP|13708-3|LNC|Arginine/Creatinine|Arginine/Creatinine
C0796900|T201|COMP|13709-1|LNC|Argininosuccinate/Creatinine|Argininosuccinate/Creatinine
C0796901|T201|COMP|13710-9|LNC|Asparagine/Creatinine|Asparagine/Creatinine
C0796902|T201|COMP|13711-7|LNC|Aspartate/Creatinine|Aspartate/Creatinine
C0796903|T201|COMP|13712-5|LNC|Azelate/Creatinine|Azelate/Creatinine
C0796904|T201|COMP|13713-3|LNC|Benzoate/Creatinine|Benzoate/Creatinine
C0796905|T201|COMP|13714-1|LNC|Beta alanine/Creatinine|Beta alanine/Creatinine
C0796906|T201|COMP|13715-8|LNC|C peptide/Creatinine|C peptide/Creatinine
C0796907|T201|COMP|13716-6|LNC|C peptide/Creatinine|C peptide/Creatinine
C0796908|T201|COMP|13717-4|LNC|Calcium/Creatinine|Calcium/Creatinine
C0796909|T201|COMP|13718-2|LNC|Carnitine.free (C0)/Creatinine|Carnitine.free (C0)/Creatinine
C0796910|T201|COMP|13719-0|LNC|Carnitine/Creatinine|Carnitine/Creatinine
C0796911|T201|COMP|13720-8|LNC|Carnosine/Creatinine|Carnosine/Creatinine
C0796912|T201|COMP|13721-6|LNC|Chloride/Creatinine|Chloride/Creatinine
C0796913|T201|COMP|13722-4|LNC|Citrate/Creatinine|Citrate/Creatinine
C0796914|T201|COMP|13723-2|LNC|Citrulline/Creatinine|Citrulline/Creatinine
C0796915|T201|COMP|13724-0|LNC|Cystathionine/Creatinine|Cystathionine/Creatinine
C0796916|T201|COMP|13725-7|LNC|Cystine/Creatinine|Cystine/Creatinine
C0796917|T201|COMP|13726-5|LNC|Decadienediate/Creatinine|Decadienediate/Creatinine
C0796918|T201|COMP|13727-3|LNC|Decenedioate/Creatinine|Decenedioate/Creatinine
C0796919|T201|COMP|13728-1|LNC|Delta aminolevulinate/Creatinine|Delta aminolevulinate/Creatinine
C0796920|T201|COMP|13729-9|LNC|Deoxypyridinoline/Creatinine|Deoxypyridinoline/Creatinine
C0796921|T201|COMP|13730-7|LNC|Deoxypyridinoline/Creatinine|Deoxypyridinoline/Creatinine
C0796922|T201|COMP|13731-5|LNC|Deoxypyridinoline/Creatinine|Deoxypyridinoline/Creatinine
C0796923|T201|COMP|13732-3|LNC|Dodecanedioate/Creatinine|Dodecanedioate/Creatinine
C0796924|T201|COMP|13733-1|LNC|DOPamine/Creatinine|DOPamine/Creatinine
C0796925|T201|COMP|13734-9|LNC|EPINEPHrine/Creatinine|EPINEPHrine/Creatinine
C0796926|T201|COMP|13735-6|LNC|Epinephrine+Norepinephrine/Creatinine|Epinephrine+Norepinephrine/Creatinine
C0796927|T201|COMP|13736-4|LNC|Estradiol/Creatinine|Estradiol/Creatinine
C0796928|T201|COMP|13737-2|LNC|Estriol/Creatinine|Estriol/Creatinine
C0796929|T201|COMP|13739-8|LNC|Estrone/Creatinine|Estrone/Creatinine
C0796930|T201|COMP|13740-6|LNC|Ethanolamine/Creatinine|Ethanolamine/Creatinine
C0796931|T201|COMP|13741-4|LNC|Ethylmalonate/Creatinine|Ethylmalonate/Creatinine
C0796932|T201|COMP|13742-2|LNC|Formate/Creatinine|Formate/Creatinine
C0796933|T201|COMP|13743-0|LNC|Fumarate/Creatinine|Fumarate/Creatinine
C0796934|T201|COMP|13744-8|LNC|Galactose/Creatinine|Galactose/Creatinine
C0796935|T201|COMP|13745-5|LNC|Glutaconate/Creatinine|Glutaconate/Creatinine
C0796936|T201|COMP|13746-3|LNC|Glutamate/Creatinine|Glutamate/Creatinine
C0796937|T201|COMP|13747-1|LNC|Glutamine/Creatinine|Glutamine/Creatinine
C0796938|T201|COMP|13748-9|LNC|Glutarate/Creatinine|Glutarate/Creatinine
C0796939|T201|COMP|13749-7|LNC|Glycerate/Creatinine|Glycerate/Creatinine
C0796940|T201|COMP|13750-5|LNC|Glycine/Creatinine|Glycine/Creatinine
C0796941|T201|COMP|13751-3|LNC|Glycolate/Creatinine|Glycolate/Creatinine
C0796942|T201|COMP|13752-1|LNC|Glyoxylate/Creatinine|Glyoxylate/Creatinine
C0796943|T201|COMP|13753-9|LNC|Hexanoylglycine/Creatinine|Hexanoylglycine/Creatinine
C0796944|T201|COMP|13754-7|LNC|Hippurate/Creatinine|Hippurate/Creatinine
C0796945|T201|COMP|13755-4|LNC|Histamine/Creatinine|Histamine/Creatinine
C0796946|T201|COMP|13756-2|LNC|Histamine/Creatinine|Histamine/Creatinine
C0796947|T201|COMP|13757-0|LNC|Histidine/Creatinine|Histidine/Creatinine
C0796948|T201|COMP|13758-8|LNC|Homocysteine/Creatinine|Homocysteine/Creatinine
C0796949|T201|COMP|13759-6|LNC|Homocystine/Creatinine|Homocystine/Creatinine
C0796950|T201|COMP|13760-4|LNC|Homovanillate/Creatinine|Homovanillate/Creatinine
C0796951|T201|COMP|13761-2|LNC|Hydroxydecanedioate/Creatinine|Hydroxydecanedioate/Creatinine
C0796952|T201|COMP|13762-0|LNC|Hydroxylysine/Creatinine|Hydroxylysine/Creatinine
C0796953|T201|COMP|13763-8|LNC|Hydroxyproline/Creatinine|Hydroxyproline/Creatinine
C0796954|T201|COMP|13764-6|LNC|Isocitrate/Creatinine|Isocitrate/Creatinine
C0796955|T201|COMP|13765-3|LNC|Isoleucine/Creatinine|Isoleucine/Creatinine
C0796956|T201|COMP|13766-1|LNC|Isovalerylglycine/Creatinine|Isovalerylglycine/Creatinine
C0796957|T201|COMP|13767-9|LNC|Lactate/Creatinine|Lactate/Creatinine
C0796958|T201|COMP|13768-7|LNC|Leucine/Creatinine|Leucine/Creatinine
C0796959|T201|COMP|13769-5|LNC|Lysine/Creatinine|Lysine/Creatinine
C0796960|T201|COMP|13770-3|LNC|Malate/Creatinine|Malate/Creatinine
C0796961|T201|COMP|13771-1|LNC|Metanephrines/Creatinine|Metanephrines/Creatinine
C0796962|T201|COMP|13772-9|LNC|Methionine/Creatinine|Methionine/Creatinine
C0796963|T201|COMP|13773-7|LNC|2-Methylcitrate/Creatinine|2-Methylcitrate/Creatinine
C0796964|T201|COMP|13774-5|LNC|Methylhippurate/Creatinine|Methylhippurate/Creatinine
C0796965|T201|COMP|13775-2|LNC|Methylmalonate/Creatinine|Methylmalonate/Creatinine
C0796966|T201|COMP|13776-0|LNC|Methylmalonate/Creatinine|Methylmalonate/Creatinine
C0796967|T201|COMP|13777-8|LNC|Methylsuccinate/Creatinine|Methylsuccinate/Creatinine
C0796968|T201|COMP|13778-6|LNC|Mevalonate/Creatinine|Mevalonate/Creatinine
C0796969|T201|COMP|13779-4|LNC|N-acetyl-L-aspartate/Creatinine|N-acetyl-L-aspartate/Creatinine
C0796970|T201|COMP|13780-2|LNC|N-acetyltyrosine/Creatinine|N-acetyltyrosine/Creatinine
C0796971|T201|COMP|13781-0|LNC|N-methylhistamine/Creatinine|N-methylhistamine/Creatinine
C0796972|T201|COMP|13782-8|LNC|Norepinephrine/Creatinine|Norepinephrine/Creatinine
C0796973|T201|COMP|13783-6|LNC|Normetanephrine/Creatinine|Normetanephrine/Creatinine
C0796974|T201|COMP|13784-4|LNC|Octanoate/Creatinine|Octanoate/Creatinine
C0796975|T201|COMP|13785-1|LNC|Octenedioate/Creatinine|Octenedioate/Creatinine
C0796976|T201|COMP|13786-9|LNC|Ornithine/Creatinine|Ornithine/Creatinine
C0796977|T201|COMP|13787-7|LNC|Orotate/Creatinine|Orotate/Creatinine
C0796978|T201|COMP|13788-5|LNC|Oxalate/Creatinine|Oxalate/Creatinine
C0796979|T201|COMP|13789-3|LNC|Phosphoethanolamine/Creatinine|Phosphoethanolamine/Creatinine
C0796980|T201|COMP|13790-1|LNC|Para nitrophenol/Creatinine|Para nitrophenol/Creatinine
C0796981|T201|COMP|13791-9|LNC|Phenylacetate/Creatinine|Phenylacetate/Creatinine
C0796982|T201|COMP|13792-7|LNC|Phenyllactate/Creatinine|Phenyllactate/Creatinine
C0796983|T201|COMP|13793-5|LNC|Phenylpropionylglycine/Creatinine|Phenylpropionylglycine/Creatinine
C0796984|T201|COMP|13794-3|LNC|Phenylpyruvate/Creatinine|Phenylpyruvate/Creatinine
C0796985|T201|COMP|13795-0|LNC|Phosphate/Creatinine|Phosphate/Creatinine
C0796986|T201|COMP|13796-8|LNC|Phosphoserine/Creatinine|Phosphoserine/Creatinine
C0796987|T201|COMP|13797-6|LNC|Porphobilinogen/Creatinine|Porphobilinogen/Creatinine
C0796988|T201|COMP|13798-4|LNC|Potassium/Creatinine|Potassium/Creatinine
C0796989|T201|COMP|13799-2|LNC|Proline/Creatinine|Proline/Creatinine
C0796990|T201|COMP|13800-8|LNC|Propionylglycine/Creatinine|Propionylglycine/Creatinine
C0796991|T201|COMP|13801-6|LNC|Protein/Creatinine|Protein/Creatinine
C0796992|T201|COMP|13802-4|LNC|Pyridinoline/Creatinine|Pyridinoline/Creatinine
C0796993|T201|COMP|13803-2|LNC|Pyridinoline/Creatinine|Pyridinoline/Creatinine
C0796994|T201|COMP|13804-0|LNC|Pyridinoline/Creatinine|Pyridinoline/Creatinine
C0796995|T201|COMP|13805-7|LNC|Pyruvate/Creatinine|Pyruvate/Creatinine
C0796996|T201|COMP|13806-5|LNC|Sarcosine/Creatinine|Sarcosine/Creatinine
C0796997|T201|COMP|13807-3|LNC|Sebacate/Creatinine|Sebacate/Creatinine
C0796998|T201|COMP|13808-1|LNC|Serine/Creatinine|Serine/Creatinine
C0796999|T201|COMP|13809-9|LNC|Sodium/Creatinine|Sodium/Creatinine
C0797000|T201|COMP|13810-7|LNC|Suberate/Creatinine|Suberate/Creatinine
C0797001|T201|COMP|13811-5|LNC|Suberylglycine/Creatinine|Suberylglycine/Creatinine
C0797002|T201|COMP|13812-3|LNC|Succinate/Creatinine|Succinate/Creatinine
C0797003|T201|COMP|13813-1|LNC|Succinylacetone/Creatinine|Succinylacetone/Creatinine
C0797004|T201|COMP|13814-9|LNC|Taurine/Creatinine|Taurine/Creatinine
C0797005|T201|COMP|13815-6|LNC|Threonine/Creatinine|Threonine/Creatinine
C0797006|T201|COMP|13816-4|LNC|Tiglylglycine/Creatinine|Tiglylglycine/Creatinine
C0797007|T201|COMP|13817-2|LNC|Tryptophan/Creatinine|Tryptophan/Creatinine
C0797008|T201|COMP|13818-0|LNC|Tyrosine/Creatinine|Tyrosine/Creatinine
C0797009|T201|COMP|13819-8|LNC|Uracil/Creatinine|Uracil/Creatinine
C0797010|T201|COMP|13820-6|LNC|Urate/Creatinine|Urate/Creatinine
C0797011|T201|COMP|13821-4|LNC|Urea nitrogen/Creatinine|Urea nitrogen/Creatinine
C0797012|T201|COMP|13822-2|LNC|Valine/Creatinine|Valine/Creatinine
C0797013|T201|COMP|13823-0|LNC|Antimony/Creatinine|Antimony/Creatinine
C0797014|T201|COMP|13824-8|LNC|Arsenic/Creatinine|Arsenic/Creatinine
C0797015|T201|COMP|13825-5|LNC|Arsenic.inorganic/Creatinine|Arsenic.inorganic/Creatinine
C0797016|T201|COMP|13826-3|LNC|Barium/Creatinine|Barium/Creatinine
C0797017|T201|COMP|13827-1|LNC|Beryllium/Creatinine|Beryllium/Creatinine
C0797018|T201|COMP|13828-9|LNC|Cadmium/Creatinine|Cadmium/Creatinine
C0797019|T201|COMP|13829-7|LNC|Copper/Creatinine|Copper/Creatinine
C0797020|T201|COMP|13830-5|LNC|Phenylglyoxylate/Creatinine|Phenylglyoxylate/Creatinine
C0797021|T201|COMP|13831-3|LNC|Vanadium/Creatinine|Vanadium/Creatinine
C0797022|T201|COMP|13832-1|LNC|Dimethylbenzene/Creatinine|Dimethylbenzene/Creatinine
C0797023|T201|COMP|13833-9|LNC|Finch feather Ab.IgE|Finch feather Ab.IgE
C0797024|T201|COMP|13834-7|LNC|IgE.total|IgE.total
C0797025|T201|COMP|13835-4|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0797026|T201|COMP|13836-2|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0797027|T201|COMP|13837-0|LNC|Blasts.CD10/100 blasts|Blasts.CD10/100 blasts
C0797028|T201|COMP|13838-8|LNC|Blasts.CD13/100 blasts|Blasts.CD13/100 blasts
C0797029|T201|COMP|13839-6|LNC|Blasts.CD14/100 blasts|Blasts.CD14/100 blasts
C0797030|T201|COMP|13840-4|LNC|Blasts.CD19/100 blasts|Blasts.CD19/100 blasts
C0797031|T201|COMP|13841-2|LNC|Blasts.CD2/100 blasts|Blasts.CD2/100 blasts
C0797032|T201|COMP|13842-0|LNC|Blasts.CD20/100 blasts|Blasts.CD20/100 blasts
C0797033|T201|COMP|13843-8|LNC|Blasts.CD33/100 blasts|Blasts.CD33/100 blasts
C0797034|T201|COMP|13844-6|LNC|Blasts.CD34/100 blasts|Blasts.CD34/100 blasts
C0797035|T201|COMP|13845-3|LNC|Blasts.CD5/100 blasts|Blasts.CD5/100 blasts
C0797036|T201|COMP|13846-1|LNC|Blasts.CD7/100 blasts|Blasts.CD7/100 blasts
C0797038|T201|COMP|13848-7|LNC|Cells.CD3+CD26+|Cells.CD3+CD26+
C0797039|T201|COMP|13850-3|LNC|Cells.CD5+CD25+|Cells.CD5+CD25+
C0797040|T201|COMP|13851-1|LNC|Cells.CD5+CD25+/100 cells|Cells.CD5+CD25+/100 cells
C0797041|T201|COMP|13852-9|LNC|Aldosterone^1H post 250 ug corticotropin IM|Aldosterone^1H post 250 ug corticotropin IM
C0797042|T201|COMP|13853-7|LNC|Aldosterone^1H post 25 mg captopril PO|Aldosterone^1H post 25 mg captopril PO
C0797043|T201|COMP|13854-5|LNC|Aldosterone^2H post 25 mg captopril PO|Aldosterone^2H post 25 mg captopril PO
C0797044|T201|COMP|13855-2|LNC|Aldosterone^30M post 250 ug corticotropin IM|Aldosterone^30M post 250 ug corticotropin IM
C0797045|T201|COMP|13856-0|LNC|Androstenedione^15M post 250 ug corticotropin IM|Androstenedione^15M post 250 ug corticotropin IM
C0797046|T201|COMP|13857-8|LNC|Androstenedione^1H post 250 ug corticotropin IM|Androstenedione^1H post 250 ug corticotropin IM
C0797047|T201|COMP|13858-6|LNC|Androstenedione^30M post 250 ug corticotropin IM|Androstenedione^30M post 250 ug corticotropin IM
C0797048|T201|COMP|13859-4|LNC|C peptide^10M post 1 mg glucagon IV|C peptide^10M post 1 mg glucagon IV
C0797049|T201|COMP|13860-2|LNC|C peptide^15M post 1 mg glucagon IV|C peptide^15M post 1 mg glucagon IV
C0797050|T201|COMP|13861-0|LNC|C peptide^5M post 1 mg glucagon IV|C peptide^5M post 1 mg glucagon IV
C0797054|T201|COMP|13865-1|LNC|Glucose^2.5H post 50 g lactose PO|Glucose^2.5H post 50 g lactose PO
C0797055|T201|COMP|13866-9|LNC|Glucose^5H post 50 g lactose PO|Glucose^5H post 50 g lactose PO
C0797056|T201|COMP|13867-7|LNC|Renin^1H post 25 mg captopril PO|Renin^1H post 25 mg captopril PO
C0797057|T201|COMP|13868-5|LNC|Renin^2H post 25 mg captopril PO|Renin^2H post 25 mg captopril PO
C0797058|T201|COMP|13869-3|LNC|Thyrotropin^1.5H post dose TRH IV|Thyrotropin^1.5H post dose TRH IV
C0797059|T201|COMP|13870-1|LNC|Thyrotropin^15M post dose TRH IV|Thyrotropin^15M post dose TRH IV
C0797060|T201|COMP|13871-9|LNC|Thyrotropin^2H post dose TRH IV|Thyrotropin^2H post dose TRH IV
C0797061|T201|COMP|13872-7|LNC|11-Deoxycortisol|11-Deoxycortisol
C0797062|T201|COMP|13873-5|LNC|Albumin.glycated/Albumin.total|Albumin.glycated/Albumin.total
C0797063|T201|COMP|13874-3|LNC|Alkaline phosphatase.liver 1|Alkaline phosphatase.liver 1
C0797064|T201|COMP|13875-0|LNC|Alkaline phosphatase.liver 2|Alkaline phosphatase.liver 2
C0797065|T201|COMP|13876-8|LNC|Beta-2 transferrin|Beta-2 transferrin
C0797066|T201|COMP|13877-6|LNC|Bilirubin|Bilirubin
C0797067|T201|COMP|13878-4|LNC|Collagen type 1 Ab.IgG|Collagen type 1 Ab.IgG
C0797068|T201|COMP|13879-2|LNC|Collagen type 2 Ab.IgG|Collagen type 2 Ab.IgG
C0797069|T201|COMP|13880-0|LNC|Collagen type 4 Ab.IgG|Collagen type 4 Ab.IgG
C0797070|T201|COMP|13881-8|LNC|Deoxypyridinoline.free/Creatinine|Deoxypyridinoline.free/Creatinine
C0797071|T201|COMP|13882-6|LNC|Androstanolone.free/Androstanolone.total|Androstanolone.free/Androstanolone.total
C0797072|T201|COMP|13883-4|LNC|Estradiol.bioavailable/Estradiol.total|Estradiol.bioavailable/Estradiol.total
C0797073|T201|COMP|13884-2|LNC|Estradiol.bioavailable|Estradiol.bioavailable
C0797074|T201|COMP|13738-0|LNC|Estrogen/Creatinine|Estrogen/Creatinine
C0797080|T201|COMP|13891-7|LNC|Motilin|Motilin
C0797081|T201|COMP|13892-5|LNC|Nitrosonaphthol|Nitrosonaphthol
C0797082|T201|COMP|13893-3|LNC|Phenylalanine|Phenylalanine
C0797083|T201|COMP|13894-1|LNC|Pregnenolone|Pregnenolone
C0797084|T201|COMP|13895-8|LNC|Sodium|Sodium
C0797085|T201|COMP|13896-6|LNC|Insulin-like growth factor-I|Insulin-like growth factor-I
C0797086|T201|COMP|13897-4|LNC|Thyrotropin.beta subunit|Thyrotropin.beta subunit
C0797087|T201|COMP|13898-2|LNC|Trichloroacetate|Trichloroacetate
C0797088|T201|COMP|13900-6|LNC|Tumor necrosis factor.alpha|Tumor necrosis factor.alpha
C0797089|T201|COMP|13901-4|LNC|Tyrosine|Tyrosine
C0797090|T201|COMP|13902-2|LNC|Urate|Urate
C0797091|T201|COMP|13903-0|LNC|Vasopressin|Vasopressin
C0797093|T201|COMP|13905-5|LNC|Meclofenamate|Meclofenamate
C0797094|T201|COMP|13906-3|LNC|Mesoridazine|Mesoridazine
C0797095|T201|COMP|13907-1|LNC|Norethindrone|Norethindrone
C0797096|T201|COMP|13908-9|LNC|Oxipurinol|Oxipurinol
C0797097|T201|COMP|13909-7|LNC|Tamoxifen|Tamoxifen
C0797098|T201|COMP|13910-5|LNC|HLA-B22|HLA-B22
C0797099|T201|COMP|13911-3|LNC|HLA-B27 related Ag|HLA-B27 related Ag
C0797100|T201|COMP|13912-1|LNC|HLA-B42|HLA-B42
C0797101|T201|COMP|13913-9|LNC|Adenovirus Ab|Adenovirus Ab
C0797102|T201|COMP|13914-7|LNC|Adenovirus Ab.IgG|Adenovirus Ab.IgG
C0797103|T201|COMP|13915-4|LNC|Adenovirus Ab.IgM|Adenovirus Ab.IgM
C0797104|T201|COMP|13916-2|LNC|Bordetella parapertussis Ag|Bordetella parapertussis Ag
C0797105|T201|COMP|13917-0|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0797106|T201|COMP|13918-8|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0797107|T201|COMP|13919-6|LNC|Hepatitis B virus core Ab.IgG|Hepatitis B virus core Ab.IgG
C0797108|T201|COMP|13920-4|LNC|HIV 2 p41 Ab|HIV 2 p41 Ab
C0797109|T201|COMP|13921-2|LNC|Mumps virus|Mumps virus
C0797110|T201|COMP|13922-0|LNC|Trichinella spiralis Ab.IgA|Trichinella spiralis Ab.IgA
C0797111|T201|COMP|13923-8|LNC|Trichinella spiralis Ab.IgM|Trichinella spiralis Ab.IgM
C0797112|T201|COMP|13924-6|LNC|Calcitonin Ab|Calcitonin Ab
C0797113|T201|COMP|13925-3|LNC|Soluble liver Ab|Soluble liver Ab
C0797114|T201|COMP|13926-1|LNC|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C0797115|T201|COMP|13927-9|LNC|Pancreatic islet cell Ab|Pancreatic islet cell Ab
C0797116|T201|COMP|13928-7|LNC|Parathyrin Ab|Parathyrin Ab
C0797117|T201|COMP|13929-5|LNC|Rheumatoid factor|Rheumatoid factor
C0797118|T201|COMP|13930-3|LNC|Rheumatoid factor|Rheumatoid factor
C0797119|T201|COMP|13931-1|LNC|Striated muscle Ab|Striated muscle Ab
C0797120|T201|COMP|13932-9|LNC|Testes Ab.IgG|Testes Ab.IgG
C0797121|T201|COMP|13933-7|LNC|Benzodiazepines|Benzodiazepines
C0797122|T201|COMP|13934-5|LNC|Butanol|Butanol
C0797123|T201|COMP|13935-2|LNC|Dichlorodifluoromethane|Dichlorodifluoromethane
C0797124|T201|COMP|13936-0|LNC|Diethyl ether|Diethyl ether
C0797125|T201|COMP|13937-8|LNC|Ethyl acetate|Ethyl acetate
C0797126|T201|COMP|13938-6|LNC|Trichloroethane|Trichloroethane
C0797127|T201|COMP|13939-4|LNC|Trichlorotrifluoroethane|Trichlorotrifluoroethane
C0797128|T201|COMP|13940-2|LNC|Dimethylbenzene|Dimethylbenzene
C0797129|T201|COMP|13941-0|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0797130|T201|COMP|13942-8|LNC|Spermatozoa.motile|Spermatozoa.motile
C0797131|T201|COMP|13943-6|LNC|Fructose|Fructose
C0797132|T201|COMP|13944-4|LNC|Phosphatase.leukocyte|Phosphatase.leukocyte
C0797133|T201|COMP|13945-1|LNC|Erythrocytes|Erythrocytes
C0797134|T201|COMP|13946-9|LNC|Complement+Immunoglobulin|Complement+Immunoglobulin
C0797135|T201|COMP|13947-7|LNC|Coccidioides immitis Ab.IgG|Coccidioides immitis Ab.IgG
C0797136|T201|COMP|13948-5|LNC|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C0797137|T201|COMP|13949-3|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0797138|T201|COMP|13950-1|LNC|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C0797139|T201|COMP|13951-9|LNC|Hepatitis A virus Ab|Hepatitis A virus Ab
C0797140|T201|COMP|13952-7|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C0797141|T201|COMP|13953-5|LNC|Hepatitis B virus little e Ab|Hepatitis B virus little e Ab
C0797142|T201|COMP|13954-3|LNC|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C0797143|T201|COMP|13955-0|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C0797144|T201|COMP|13956-8|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C0797145|T201|COMP|13957-6|LNC|Clostridioides difficile toxin A|Clostridioides difficile toxin A
C0797146|T201|COMP|13958-4|LNC|Arsenic|Arsenic
C0797147|T201|COMP|13959-2|LNC|Calcium.ionized|Calcium.ionized
C0797148|T201|COMP|13960-0|LNC|Coproporphyrin|Coproporphyrin
C0797149|T201|COMP|13961-8|LNC|Mercury|Mercury
C0797150|T201|COMP|13962-6|LNC|Beta glucuronidase|Beta glucuronidase
C0797151|T201|COMP|13963-4|LNC|Orotate|Orotate
C0797152|T201|COMP|13964-2|LNC|Methylmalonate|Methylmalonate
C0797153|T201|COMP|13965-9|LNC|Homocysteine|Homocysteine
C0797154|T201|COMP|13966-7|LNC|Cystine|Cystine
C0797155|T201|COMP|13967-5|LNC|Sex hormone binding globulin|Sex hormone binding globulin
C0797156|T201|COMP|13968-3|LNC|Penicillin|Penicillin
C0797157|T201|COMP|13969-1|LNC|Creatine kinase.MB|Creatine kinase.MB
C0797158|T201|COMP|13970-9|LNC|Delta tocopherol|Delta tocopherol
C0797159|T201|COMP|13971-7|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C0797160|T201|COMP|13972-5|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0797161|T201|COMP|13973-3|LNC|Prealbumin/Protein.total|Prealbumin/Protein.total
C0797162|T201|COMP|13974-1|LNC|Albumin/Protein.total|Albumin/Protein.total
C0797163|T201|COMP|13975-8|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0797164|T201|COMP|13976-6|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C0797165|T201|COMP|13977-4|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0797166|T201|COMP|13978-2|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0797167|T201|COMP|13979-0|LNC|Prealbumin/Protein.total|Prealbumin/Protein.total
C0797168|T201|COMP|13980-8|LNC|Albumin/Protein.total|Albumin/Protein.total
C0797169|T201|COMP|13981-6|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0797170|T201|COMP|13982-4|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C0797171|T201|COMP|13983-2|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0797172|T201|COMP|13984-0|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0797173|T201|COMP|13985-7|LNC|Prealbumin/Protein.total|Prealbumin/Protein.total
C0797174|T201|COMP|13986-5|LNC|Albumin/Protein.total|Albumin/Protein.total
C0797175|T201|COMP|13987-3|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0797176|T201|COMP|13988-1|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C0797177|T201|COMP|13989-9|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0797178|T201|COMP|13990-7|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0797179|T201|COMP|13991-5|LNC|Prealbumin/Protein.total|Prealbumin/Protein.total
C0797180|T201|COMP|13992-3|LNC|Albumin/Protein.total|Albumin/Protein.total
C0797181|T201|COMP|13993-1|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0797182|T201|COMP|13994-9|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C0797183|T201|COMP|13995-6|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0797184|T201|COMP|13996-4|LNC|Hydroxyproline/Creatinine|Hydroxyproline/Creatinine
C0797185|T201|COMP|13997-2|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C0797186|T201|COMP|13998-0|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C0797187|T201|COMP|13999-8|LNC|Transferrin.carbohydrate deficient|Transferrin.carbohydrate deficient
C0797188|T201|COMP|14000-4|LNC|Urea nitrogen|Urea nitrogen
C0797189|T201|COMP|14001-2|LNC|IgE|IgE
C0797190|T201|COMP|14002-0|LNC|IgM|IgM
C0797191|T201|COMP|14003-8|LNC|Carbon dioxide|Carbon dioxide
C0797192|T201|COMP|14004-6|LNC|Prostaglandin A|Prostaglandin A
C0797193|T201|COMP|14005-3|LNC|Prostaglandin E1|Prostaglandin E1
C0797194|T201|COMP|14006-1|LNC|Prostaglandin E2|Prostaglandin E2
C0797195|T201|COMP|14007-9|LNC|Prostaglandin F2 alpha|Prostaglandin F2 alpha
C0797196|T201|COMP|14008-7|LNC|Phosphatidylcholine Ab.IgG|Phosphatidylcholine Ab.IgG
C0797197|T201|COMP|14009-5|LNC|Phosphatidylcholine Ab.IgM|Phosphatidylcholine Ab.IgM
C0797198|T201|COMP|14010-3|LNC|Phosphatidylcholine Ab.IgA|Phosphatidylcholine Ab.IgA
C0797199|T201|COMP|14011-1|LNC|Platelet associated Ab.IgA|Platelet associated Ab.IgA
C0797200|T201|COMP|14012-9|LNC|Platelet associated Ab.IgG|Platelet associated Ab.IgG
C0797201|T201|COMP|14013-7|LNC|Platelet associated Ab.IgM|Platelet associated Ab.IgM
C0797202|T201|COMP|14014-5|LNC|Thyroxine.prealbumin bound|Thyroxine.prealbumin bound
C0797203|T201|COMP|14015-2|LNC|Thyroxine.prealbumin bound/Prealbumin|Thyroxine.prealbumin bound/Prealbumin
C0797204|T201|COMP|14016-0|LNC|Thyroxine.thyroxine binding globulin bound|Thyroxine.thyroxine binding globulin bound
C0797205|T201|COMP|14017-8|LNC|Cells.CD22/100 cells|Cells.CD22/100 cells
C0797206|T201|COMP|14018-6|LNC|Cells.CD23/100 cells|Cells.CD23/100 cells
C0797207|T201|COMP|14019-4|LNC|HTLV I+II gp46 Ab|HTLV I+II gp46 Ab
C0797208|T201|COMP|14020-2|LNC|HTLV I+II p19 Ab|HTLV I+II p19 Ab
C0797209|T201|COMP|14021-0|LNC|HTLV I+II p24 Ab|HTLV I+II p24 Ab
C0797210|T201|COMP|14022-8|LNC|HTLV I+II p26 Ab|HTLV I+II p26 Ab
C0797211|T201|COMP|14023-6|LNC|HTLV I+II p28 Ab|HTLV I+II p28 Ab
C0797212|T201|COMP|14024-4|LNC|HTLV I+II p32 Ab|HTLV I+II p32 Ab
C0797213|T201|COMP|14025-1|LNC|HTLV I+II p36 Ab|HTLV I+II p36 Ab
C0797214|T201|COMP|14026-9|LNC|HTLV I+II p53 Ab|HTLV I+II p53 Ab
C0797215|T201|COMP|14027-7|LNC|HTLV I+II rgp21 Ab|HTLV I+II rgp21 Ab
C0797216|T201|COMP|14028-5|LNC|HTLV I+II rgp46-I Ab|HTLV I+II rgp46-I Ab
C0797217|T201|COMP|14029-3|LNC|HTLV I+II rgp46-II Ab|HTLV I+II rgp46-II Ab
C0797219|T201|COMP|14031-9|LNC|Ciprofloxacin^peak|Ciprofloxacin^peak
C0797220|T201|COMP|14032-7|LNC|Ciprofloxacin^trough|Ciprofloxacin^trough
C0797221|T201|COMP|14033-5|LNC|1,4-Dioxane|1,4-Dioxane
C0797222|T201|COMP|14034-3|LNC|Rheumatoid factor|Rheumatoid factor
C0797223|T201|COMP|14035-0|LNC|Cryptomeria japonica Ab.IgE|Cryptomeria japonica Ab.IgE
C0797224|T201|COMP|14036-8|LNC|Dermatophagoides microceras Ab.IgE|Dermatophagoides microceras Ab.IgE
C0797225|T201|COMP|14037-6|LNC|Fox Ab.IgE|Fox Ab.IgE
C0797226|T201|COMP|14038-4|LNC|Todarodes pacificus Ab.IgE|Todarodes pacificus Ab.IgE
C0797227|T201|COMP|14039-2|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0797228|T201|COMP|14040-0|LNC|Carbon dioxide|Carbon dioxide
C0797229|T201|COMP|14041-8|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0797230|T201|COMP|14042-6|LNC|Corticosterone|Corticosterone
C0797231|T201|COMP|14043-4|LNC|Cortisol.free|Cortisol.free
C0797232|T201|COMP|14044-2|LNC|Cortisone|Cortisone
C0797233|T201|COMP|14045-9|LNC|D-lactate|D-lactate
C0797234|T201|COMP|14046-7|LNC|D-lactate|D-lactate
C0797235|T201|COMP|14047-5|LNC|Androstanolone.free|Androstanolone.free
C0797236|T201|COMP|14048-3|LNC|Elastase.pancreatic|Elastase.pancreatic
C0797237|T201|COMP|14049-1|LNC|Epidermal growth factor|Epidermal growth factor
C0797238|T201|COMP|14050-9|LNC|Epidermal growth factor receptor|Epidermal growth factor receptor
C0797239|T201|COMP|14051-7|LNC|Estrogen binding protein|Estrogen binding protein
C0797240|T201|COMP|14052-5|LNC|Formate|Formate
C0797241|T201|COMP|14053-3|LNC|Homocystine|Homocystine
C0797242|T201|COMP|14054-1|LNC|Prostaglandin D2|Prostaglandin D2
C0797243|T201|COMP|14055-8|LNC|Sodium|Sodium
C0797244|T201|COMP|14056-6|LNC|carBAMazepine 10,11-Epoxide.free|carBAMazepine 10,11-Epoxide.free
C0797245|T201|COMP|14057-4|LNC|carBAMazepine.free|carBAMazepine.free
C0797246|T201|COMP|14058-2|LNC|Ciprofloxacin^peak|Ciprofloxacin^peak
C0797247|T201|COMP|14059-0|LNC|Ciprofloxacin^trough|Ciprofloxacin^trough
C0797248|T201|COMP|14060-8|LNC|Cyclobenzaprine|Cyclobenzaprine
C0797249|T201|COMP|14061-6|LNC|Cyclobenzaprine|Cyclobenzaprine
C0797250|T201|COMP|14062-4|LNC|Dexamethasone|Dexamethasone
C0797251|T201|COMP|14063-2|LNC|Dezocine|Dezocine
C0797252|T201|COMP|14064-0|LNC|Diethylstilbestrol|Diethylstilbestrol
C0797253|T201|COMP|14065-7|LNC|Diflunisal|Diflunisal
C0797254|T201|COMP|14066-5|LNC|Dihydrocodeine|Dihydrocodeine
C0797255|T201|COMP|14067-3|LNC|Dihydrocodeine|Dihydrocodeine
C0797256|T201|COMP|14068-1|LNC|Triamterene+hydroCHLOROthiazide|Triamterene+hydroCHLOROthiazide
C0797257|T201|COMP|14069-9|LNC|Estazolam|Estazolam
C0797258|T201|COMP|14070-7|LNC|fluPHENAZine|fluPHENAZine
C0797259|T201|COMP|14071-5|LNC|Ibuprofen|Ibuprofen
C0797260|T201|COMP|14072-3|LNC|Monoacetyldapsone|Monoacetyldapsone
C0797261|T201|COMP|14073-1|LNC|Phenytoin|Phenytoin
C0797262|T201|COMP|14074-9|LNC|Spironolactone|Spironolactone
C0797263|T201|COMP|14075-6|LNC|Sulfapyridine|Sulfapyridine
C0797264|T201|COMP|14076-4|LNC|Complement total hemolytic CH100|Complement total hemolytic CH100
C0797265|T201|COMP|14077-2|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0797266|T201|COMP|14078-0|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0797267|T201|COMP|14079-8|LNC|Brucella canis Ab.IgG|Brucella canis Ab.IgG
C0797268|T201|COMP|14080-6|LNC|Brucella canis Ab.IgM|Brucella canis Ab.IgM
C0797269|T201|COMP|14081-4|LNC|Coliform bacteria|Coliform bacteria
C0797270|T201|COMP|14082-2|LNC|Echinococcus sp Ab.IgG|Echinococcus sp Ab.IgG
C0797271|T201|COMP|14083-0|LNC|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C0797272|T201|COMP|14084-8|LNC|Herpes simplex virus 1|Herpes simplex virus 1
C0797273|T201|COMP|14085-5|LNC|Herpes simplex virus 2|Herpes simplex virus 2
C0797274|T201|COMP|14086-3|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C0797275|T201|COMP|14087-1|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C0797276|T201|COMP|14088-9|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C0797277|T201|COMP|14089-7|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0797278|T201|COMP|14090-5|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C0797279|T201|COMP|14091-3|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C0797280|T201|COMP|14092-1|LNC|HIV 1 Ab|HIV 1 Ab
C0797281|T201|COMP|14093-9|LNC|Bacteria identified|Bacteria identified
C0797282|T201|COMP|14094-7|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C0797283|T201|COMP|14095-4|LNC|Fibronectin aggregate Ab.IgG|Fibronectin aggregate Ab.IgG
C0797284|T201|COMP|14096-2|LNC|Intercalated disk Ab|Intercalated disk Ab
C0797285|T201|COMP|14097-0|LNC|Antimony|Antimony
C0797286|T201|COMP|14098-8|LNC|Dimethylsulfoxide|Dimethylsulfoxide
C0797287|T201|COMP|14099-6|LNC|Nickel|Nickel
C0797288|T201|COMP|14100-2|LNC|Strontium|Strontium
C0797289|T201|COMP|14101-0|LNC|Strychnine|Strychnine
C0797290|T201|COMP|14102-8|LNC|Strychnine|Strychnine
C0797291|T201|COMP|14103-6|LNC|Epithelial cells|Epithelial cells
C0797292|T201|COMP|14104-4|LNC|Ustilago nuda+Ustilago tritici Ab.IgE|Ustilago nuda+Ustilago tritici Ab.IgE
C0797293|T201|COMP|14105-1|LNC|Leukocytes|Leukocytes
C0797294|T201|COMP|14106-9|LNC|Lymphocytes|Lymphocytes
C0797295|T201|COMP|14107-7|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C0797296|T201|COMP|14108-5|LNC|Cells.CD16c+CD56+|Cells.CD16c+CD56+
C0797297|T201|COMP|14109-3|LNC|Cells.CD16c+CD56+/100 cells|Cells.CD16c+CD56+/100 cells
C0797298|T201|COMP|14112-7|LNC|Cells.CD25+CD19+/100 cells|Cells.CD25+CD19+/100 cells
C0797299|T201|COMP|14113-5|LNC|Cells.CD56|Cells.CD56
C0797301|T201|COMP|14115-0|LNC|Collagen crosslinked N-telopeptide/Creatinine|Collagen crosslinked N-telopeptide/Creatinine
C0797302|T201|COMP|14116-8|LNC|IgG synthesis rate|IgG synthesis rate
C0797303|T201|COMP|14117-6|LNC|IgG clearance/Albumin clearance|IgG clearance/Albumin clearance
C0797304|T201|COMP|14118-4|LNC|Lactate|Lactate
C0797305|T201|COMP|14119-2|LNC|Lactate dehydrogenase 1/Lactate dehydrogenase 2|Lactate dehydrogenase 1/Lactate dehydrogenase 2
C0797307|T201|COMP|14121-8|LNC|Pyruvate|Pyruvate
C0797308|T201|COMP|14122-6|LNC|Pyruvate|Pyruvate
C0797309|T201|COMP|14123-4|LNC|Thyroxine.albumin bound/Albumin|Thyroxine.albumin bound/Albumin
C0797310|T201|COMP|14124-2|LNC|Bacteria|Bacteria
C0797311|T201|COMP|14125-9|LNC|Entamoeba histolytica|Entamoeba histolytica
C0797312|T201|COMP|14126-7|LNC|HIV 1 gp120+gp160 Ab|HIV 1 gp120+gp160 Ab
C0797313|T201|COMP|14127-5|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0797314|T201|COMP|14128-3|LNC|Rabies virus Ab|Rabies virus Ab
C0797315|T201|COMP|14129-1|LNC|Respiratory syncytial virus|Respiratory syncytial virus
C0797316|T201|COMP|14130-9|LNC|Estrogen receptor|Estrogen receptor
C0797317|T201|COMP|14131-7|LNC|PM-1 Ab|PM-1 Ab
C0797318|T201|COMP|14132-5|LNC|Color|Color
C0797319|T201|COMP|14133-3|LNC|Maple silver Ab.IgE|Maple silver Ab.IgE
C0797320|T201|COMP|14134-1|LNC|Hemoglobin.free|Hemoglobin.free
C0797321|T201|COMP|14135-8|LNC|Cells.CD3+CD8+|Cells.CD3+CD8+
C0797322|T201|COMP|14136-6|LNC|Cells.CD34|Cells.CD34
C0797323|T201|COMP|14137-4|LNC|Glucose^5.5H post 75 g glucose PO|Glucose^5.5H post 75 g glucose PO
C0797324|T201|COMP|14138-2|LNC|Ketones^30M post XXX challenge|Ketones^30M post XXX challenge
C0797325|T201|COMP|14139-0|LNC|Ketones^4H post XXX challenge|Ketones^4H post XXX challenge
C0797326|T201|COMP|14140-8|LNC|Ketones^5H post XXX challenge|Ketones^5H post XXX challenge
C0797327|T201|COMP|14141-6|LNC|Ketones^6H post XXX challenge|Ketones^6H post XXX challenge
C0797328|T201|COMP|14142-4|LNC|Somatotropin^15M post XXX challenge|Somatotropin^15M post XXX challenge
C0797329|T201|COMP|14143-2|LNC|Somatotropin^20M post XXX challenge|Somatotropin^20M post XXX challenge
C0797330|T201|COMP|14144-0|LNC|Somatotropin^2H post XXX challenge|Somatotropin^2H post XXX challenge
C0797331|T201|COMP|14145-7|LNC|Somatotropin^40M post XXX challenge|Somatotropin^40M post XXX challenge
C0797332|T201|COMP|14146-5|LNC|Somatotropin^1H post XXX challenge|Somatotropin^1H post XXX challenge
C0797333|T201|COMP|14147-3|LNC|Somatotropin^1.5H post XXX challenge|Somatotropin^1.5H post XXX challenge
C0797334|T201|COMP|14148-1|LNC|18-Hydroxycortisol|18-Hydroxycortisol
C0797335|T201|COMP|14149-9|LNC|Corticotropin.big fragment|Corticotropin.big fragment
C0797336|T201|COMP|14151-5|LNC|Bicarbonate|Bicarbonate
C0797337|T201|COMP|14152-3|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C0797338|T201|COMP|14153-1|LNC|Carnitine esters/Creatinine|Carnitine esters/Creatinine
C0797339|T201|COMP|14154-9|LNC|Cholesterol sulfate|Cholesterol sulfate
C0797340|T201|COMP|14155-6|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C0797341|T201|COMP|14156-4|LNC|Coproporphyrin|Coproporphyrin
C0797342|T201|COMP|14157-2|LNC|Coproporphyrin|Coproporphyrin
C0797343|T201|COMP|14158-0|LNC|Cortisol|Cortisol
C0797344|T201|COMP|14159-8|LNC|Cortisone|Cortisone
C0797345|T201|COMP|14160-6|LNC|Estrone.unconjugated/Estrone.total|Estrone.unconjugated/Estrone.total
C0797346|T201|COMP|14161-4|LNC|Formaldehyde|Formaldehyde
C0797347|T201|COMP|14162-2|LNC|Gamma melanocyte stimulating hormone|Gamma melanocyte stimulating hormone
C0797348|T201|COMP|14163-0|LNC|IgA.secretory|IgA.secretory
C0797349|T201|COMP|14164-8|LNC|Immunosuppressive acidic protein|Immunosuppressive acidic protein
C0797350|T201|COMP|14165-5|LNC|Lactate|Lactate
C0797351|T201|COMP|14166-3|LNC|Methane|Methane
C0797352|T201|COMP|14167-1|LNC|N-methylimidazoleacetate|N-methylimidazoleacetate
C0797353|T201|COMP|14168-9|LNC|Palatinase|Palatinase
C0797354|T201|COMP|14169-7|LNC|Peptide histidine isoleucine|Peptide histidine isoleucine
C0797355|T201|COMP|14170-5|LNC|Pituitary glycoprotein hormone.alpha subunit|Pituitary glycoprotein hormone.alpha subunit
C0797356|T201|COMP|14171-3|LNC|Porphyrins|Porphyrins
C0797357|T201|COMP|14172-1|LNC|Potassium|Potassium
C0797358|T201|COMP|14173-9|LNC|Progesterone.free|Progesterone.free
C0797359|T201|COMP|14174-7|LNC|Prostaglandin F2 alpha|Prostaglandin F2 alpha
C0797360|T201|COMP|14175-4|LNC|Protoporphyrin|Protoporphyrin
C0797361|T201|COMP|14176-2|LNC|Pyrroles|Pyrroles
C0797362|T201|COMP|14177-0|LNC|Growth hormone-releasing hormone|Growth hormone-releasing hormone
C0797363|T201|COMP|14178-8|LNC|Sucrase|Sucrase
C0797364|T201|COMP|14179-6|LNC|Tissue polypeptide Ag|Tissue polypeptide Ag
C0797365|T201|COMP|14180-4|LNC|Uroporphyrin|Uroporphyrin
C0797366|T201|COMP|14181-2|LNC|Uroporphyrin|Uroporphyrin
C0797367|T201|COMP|14182-0|LNC|Thrombin antithrombin complex Ag|Thrombin antithrombin complex Ag
C0797368|T201|COMP|14183-8|LNC|Aprobarbital|Aprobarbital
C0797369|T201|COMP|14184-6|LNC|Atropine|Atropine
C0797370|T201|COMP|14185-3|LNC|methIMAzole|methIMAzole
C0797371|T201|COMP|14186-1|LNC|Methylprednisolone|Methylprednisolone
C0797372|T201|COMP|14187-9|LNC|OKT3|OKT3
C0797373|T201|COMP|14188-7|LNC|Omeprazole|Omeprazole
C0797374|T201|COMP|14189-5|LNC|Phenyltoloxamine|Phenyltoloxamine
C0797375|T201|COMP|14190-3|LNC|Phenytoin.free|Phenytoin.free
C0797376|T201|COMP|14191-1|LNC|Prazosin|Prazosin
C0797377|T201|COMP|14192-9|LNC|Triazolam|Triazolam
C0797378|T201|COMP|14193-7|LNC|Tripelennamine|Tripelennamine
C0797379|T201|COMP|14194-5|LNC|Spermatozoa.progressive/100 spermatozoa|Spermatozoa.progressive/100 spermatozoa
C0797380|T201|COMP|14195-2|LNC|Complement C3b.inactive|Complement C3b.inactive
C0797381|T201|COMP|14196-0|LNC|Reticulocytes|Reticulocytes
C0797383|T201|COMP|14198-6|LNC|Chlamydophila psittaci Ab|Chlamydophila psittaci Ab
C0797384|T201|COMP|14199-4|LNC|Chlamydia trachomatis B Ab.IgA|Chlamydia trachomatis B Ab.IgA
C0797385|T201|COMP|14200-0|LNC|Chlamydia trachomatis B Ab.IgG|Chlamydia trachomatis B Ab.IgG
C0797386|T201|COMP|14201-8|LNC|Chlamydia trachomatis B Ab.IgM|Chlamydia trachomatis B Ab.IgM
C0797387|T201|COMP|14202-6|LNC|Chlamydia trachomatis C Ab.IgA|Chlamydia trachomatis C Ab.IgA
C0797388|T201|COMP|14203-4|LNC|Chlamydia trachomatis C Ab.IgG|Chlamydia trachomatis C Ab.IgG
C0797389|T201|COMP|14204-2|LNC|Chlamydia trachomatis C Ab.IgM|Chlamydia trachomatis C Ab.IgM
C0797390|T201|COMP|14205-9|LNC|Coccidioides immitis Ag|Coccidioides immitis Ag
C0797391|T201|COMP|14206-7|LNC|Coccidioides immitis exoantigen identification|Coccidioides immitis exoantigen identification
C0797392|T201|COMP|14207-5|LNC|DNAse B Ab.Streptococcal|DNAse B Ab.Streptococcal
C0797393|T201|COMP|14208-3|LNC|Filaria Ab.IgG4|Filaria Ab.IgG4
C0797394|T201|COMP|14209-1|LNC|Francisella tularensis Ab.IgA|Francisella tularensis Ab.IgA
C0797395|T201|COMP|14210-9|LNC|Giardia lamblia Ag|Giardia lamblia Ag
C0797396|T201|COMP|14211-7|LNC|Hepatitis E virus Ab.IgG|Hepatitis E virus Ab.IgG
C0797397|T201|COMP|14212-5|LNC|Hepatitis E virus Ab.IgM|Hepatitis E virus Ab.IgM
C0797398|T201|COMP|14213-3|LNC|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C0797399|T201|COMP|14214-1|LNC|Histoplasma capsulatum exoantigen identification|Histoplasma capsulatum exoantigen identification
C0797400|T201|COMP|14215-8|LNC|HTLV I g46 Ab|HTLV I g46 Ab
C0797401|T201|COMP|14216-6|LNC|HTLV I gp46 Ab|HTLV I gp46 Ab
C0797402|T201|COMP|14217-4|LNC|HTLV I p19 Ab|HTLV I p19 Ab
C0797403|T201|COMP|14218-2|LNC|HTLV I p24 Ab|HTLV I p24 Ab
C0797404|T201|COMP|14219-0|LNC|HTLV I p26 Ab|HTLV I p26 Ab
C0797405|T201|COMP|14220-8|LNC|HTLV I p28 Ab|HTLV I p28 Ab
C0797406|T201|COMP|14221-6|LNC|HTLV I p32 Ab|HTLV I p32 Ab
C0797407|T201|COMP|14222-4|LNC|HTLV I p36 Ab|HTLV I p36 Ab
C0797408|T201|COMP|14223-2|LNC|HTLV I p53 Ab|HTLV I p53 Ab
C0797409|T201|COMP|14224-0|LNC|HTLV I rgp21 Ab|HTLV I rgp21 Ab
C0797410|T201|COMP|14225-7|LNC|HTLV II g46 Ab|HTLV II g46 Ab
C0797411|T201|COMP|14226-5|LNC|Nocardia sp identified|Nocardia sp identified
C0797412|T201|COMP|14227-3|LNC|Salmonella typhi H D Ab|Salmonella typhi H D Ab
C0797413|T201|COMP|14228-1|LNC|Cells.estrogen receptor/100 cells|Cells.estrogen receptor/100 cells
C0797414|T201|COMP|14229-9|LNC|P53 protein Ag|P53 protein Ag
C0797415|T201|COMP|14230-7|LNC|Cells.progesterone receptor/100 cells|Cells.progesterone receptor/100 cells
C0797416|T201|COMP|14231-5|LNC|H2a-H2b DNA Ab.IgG|H2a-H2b DNA Ab.IgG
C0797417|T201|COMP|14232-3|LNC|Adrenal Ab|Adrenal Ab
C0797418|T201|COMP|14233-1|LNC|Beta tubulin Ab.IgG|Beta tubulin Ab.IgG
C0797419|T201|COMP|14234-9|LNC|Beta tubulin Ab.IgM|Beta tubulin Ab.IgM
C0797420|T201|COMP|14235-6|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C0797421|T201|COMP|14236-4|LNC|Mitochondria Ab|Mitochondria Ab
C0797422|T201|COMP|14237-2|LNC|Myelin basic protein Ab.IgA|Myelin basic protein Ab.IgA
C0797423|T201|COMP|14238-0|LNC|Myelin basic protein Ab.IgG|Myelin basic protein Ab.IgG
C0797424|T201|COMP|14239-8|LNC|Myelin basic protein Ab.IgM|Myelin basic protein Ab.IgM
C0797425|T201|COMP|14240-6|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C0797426|T201|COMP|14241-4|LNC|Parietal cell Ab|Parietal cell Ab
C0797427|T201|COMP|14242-2|LNC|Phosphatidylcholine Ab.IgA|Phosphatidylcholine Ab.IgA
C0797428|T201|COMP|14243-0|LNC|Phosphatidylcholine Ab.IgG|Phosphatidylcholine Ab.IgG
C0797429|T201|COMP|14244-8|LNC|Phosphatidylcholine Ab.IgM|Phosphatidylcholine Ab.IgM
C0797430|T201|COMP|14245-5|LNC|Phosphatidylserine Ab.IgG|Phosphatidylserine Ab.IgG
C0797431|T201|COMP|14246-3|LNC|Phosphatidylserine Ab.IgM|Phosphatidylserine Ab.IgM
C0797432|T201|COMP|14247-1|LNC|Purkinje cells Ab|Purkinje cells Ab
C0797433|T201|COMP|14248-9|LNC|Purkinje cells Ab|Purkinje cells Ab
C0797434|T201|COMP|14249-7|LNC|Purkinje cells Ab|Purkinje cells Ab
C0797435|T201|COMP|14250-5|LNC|Purkinje cells Ab.IgG|Purkinje cells Ab.IgG
C0797437|T201|COMP|14252-1|LNC|Smooth muscle Ab|Smooth muscle Ab
C0797438|T201|COMP|14253-9|LNC|Somatotropin Ab|Somatotropin Ab
C0797439|T201|COMP|14254-7|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C0797440|T201|COMP|14255-4|LNC|Thyrotropin blocking Ab|Thyrotropin blocking Ab
C0797441|T201|COMP|14256-2|LNC|Tetrachlorodiphenylethane|Tetrachlorodiphenylethane
C0797442|T201|COMP|14257-0|LNC|Tetrachlorodiphenylethane|Tetrachlorodiphenylethane
C0797443|T201|COMP|14258-8|LNC|1,4-Dioxane|1,4-Dioxane
C0797444|T201|COMP|14259-6|LNC|1-Pentanol|1-Pentanol
C0797445|T201|COMP|14260-4|LNC|Bromoform|Bromoform
C0797446|T201|COMP|14261-2|LNC|Codeine|Codeine
C0797447|T201|COMP|14262-0|LNC|Dichlorodiphenyldichloroethylene|Dichlorodiphenyldichloroethylene
C0797448|T201|COMP|14263-8|LNC|Dichlorodiphenyltrichloroethane|Dichlorodiphenyltrichloroethane
C0797449|T201|COMP|14264-6|LNC|Enflurane|Enflurane
C0797450|T201|COMP|14265-3|LNC|Isobutyl acetate|Isobutyl acetate
C0797451|T201|COMP|14266-1|LNC|Methoxyflurane|Methoxyflurane
C0797452|T201|COMP|14267-9|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0797453|T201|COMP|14268-7|LNC|Butyl acetate|Butyl acetate
C0797454|T201|COMP|14269-5|LNC|Sec-butyl acetate|Sec-butyl acetate
C0797455|T201|COMP|14270-3|LNC|Tert-butyl acetate|Tert-butyl acetate
C0797456|T201|COMP|14271-1|LNC|Character|Character
C0797457|T201|COMP|14272-9|LNC|Liver kidney microsomal Ab|Liver kidney microsomal Ab
C0797458|T201|COMP|14273-7|LNC|Reticulin Ab.IgA|Reticulin Ab.IgA
C0797459|T201|COMP|14274-5|LNC|Uroporphyrin|Uroporphyrin
C0797460|T201|COMP|14275-2|LNC|Immune complex|Immune complex
C0797461|T201|COMP|14276-0|LNC|Hemoglobin F distribution|Hemoglobin F distribution
C0797462|T201|COMP|14277-8|LNC|Neutrophil cytoplasmic Ab.classic|Neutrophil cytoplasmic Ab.classic
C0797463|T201|COMP|14278-6|LNC|Neutrophil cytoplasmic Ab.perinuclear|Neutrophil cytoplasmic Ab.perinuclear
C0797464|T201|COMP|14282-8|LNC|Acylcarnitine|Acylcarnitine
C0797465|T201|COMP|14283-6|LNC|Acylcarnitine|Acylcarnitine
C0797466|T201|COMP|14284-4|LNC|Beta glucuronidase|Beta glucuronidase
C0797467|T201|COMP|14285-1|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C0797468|T201|COMP|14286-9|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C0797469|T201|COMP|14287-7|LNC|Carnitine|Carnitine
C0797470|T201|COMP|14288-5|LNC|Carnitine|Carnitine
C0797471|T201|COMP|14290-1|LNC|Erythrocytes|Erythrocytes
C0797472|T201|COMP|14291-9|LNC|Follitropin^baseline|Follitropin^baseline
C0797473|T201|COMP|14292-7|LNC|IgE|IgE
C0797474|T201|COMP|14293-5|LNC|Insulin^baseline|Insulin^baseline
C0797475|T201|COMP|14294-3|LNC|Lysosomal enzymes screen|Lysosomal enzymes screen
C0797476|T201|COMP|14295-0|LNC|Organic acids/Creatinine|Organic acids/Creatinine
C0797477|T201|COMP|14296-8|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C0797478|T201|COMP|14297-6|LNC|Thyrotropin|Thyrotropin
C0797479|T201|COMP|14298-4|LNC|Plasma units available|Plasma units available
C0797480|T201|COMP|14299-2|LNC|Cryoprecipitate units available|Cryoprecipitate units available
C0797481|T201|COMP|14300-8|LNC|Plateletpheresis units available|Plateletpheresis units available
C0797482|T201|COMP|14301-6|LNC|Platelet concentrate units available|Platelet concentrate units available
C0797483|T201|COMP|14302-4|LNC|Packed erythrocytes units available|Packed erythrocytes units available
C0797484|T201|COMP|14303-2|LNC|Transfuse plateletpheresis|Transfuse plateletpheresis
C0797485|T201|COMP|14304-0|LNC|Measles virus Ab.IgG^1st specimen|Measles virus Ab.IgG^1st specimen
C0797486|T201|COMP|14305-7|LNC|Measles virus Ab.IgG^2nd specimen|Measles virus Ab.IgG^2nd specimen
C0797487|T201|COMP|14306-5|LNC|Varicella zoster virus Ab.IgG^1st specimen|Varicella zoster virus Ab.IgG^1st specimen
C0797488|T201|COMP|14307-3|LNC|Varicella zoster virus Ab.IgG^2nd specimen|Varicella zoster virus Ab.IgG^2nd specimen
C0797489|T201|COMP|14308-1|LNC|Amphetamines|Amphetamines
C0797490|T201|COMP|14309-9|LNC|Amphetamines|Amphetamines
C0797491|T201|COMP|14310-7|LNC|Phencyclidine|Phencyclidine
C0797492|T201|COMP|14311-5|LNC|Phencyclidine|Phencyclidine
C0797493|T201|COMP|14312-3|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0797494|T201|COMP|14313-1|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0797495|T201|COMP|14314-9|LNC|Benzoylecgonine|Benzoylecgonine
C0797496|T201|COMP|14315-6|LNC|Benzoylecgonine|Benzoylecgonine
C0797497|T201|COMP|14316-4|LNC|Benzodiazepines|Benzodiazepines
C0797501|T201|COMP|14320-6|LNC|Bacteria identified|Bacteria identified
C0797502|T201|COMP|14321-4|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C0797503|T201|COMP|14322-2|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C0797504|T201|COMP|14323-0|LNC|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C0797505|T201|COMP|14324-8|LNC|Escherichia coli K1 Ag|Escherichia coli K1 Ag
C0797506|T201|COMP|14325-5|LNC|Bacteria identified|Bacteria identified
C0797507|T201|COMP|14326-3|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0797508|T201|COMP|14327-1|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C0797509|T201|COMP|14328-9|LNC|Leukocytes|Leukocytes
C0797510|T201|COMP|14329-7|LNC|Mucus|Mucus
C0797511|T201|COMP|14330-5|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0797512|T201|COMP|14331-3|LNC|Erythrocytes|Erythrocytes
C0797513|T201|COMP|14332-1|LNC|Para aminosalicylate|Para aminosalicylate
C0797514|T201|COMP|14333-9|LNC|Lead|Lead
C0797515|T201|COMP|14334-7|LNC|Lithium|Lithium
C0797516|T201|COMP|14335-4|LNC|Optical density|Optical density
C0797517|T201|COMP|14336-2|LNC|Ethanol|Ethanol
C0797518|T201|COMP|34540-5|LNC|Phenytoin free & total panel|Phenytoin free & total panel
C0797519|T201|COMP|14338-8|LNC|Prealbumin|Prealbumin
C0797520|T201|COMP|14339-6|LNC|IgG/Protein.total|IgG/Protein.total
C0797521|T201|COMP|14340-4|LNC|Gammopathy|Gammopathy
C0797522|T201|COMP|14341-2|LNC|Globulin/Protein.total|Globulin/Protein.total
C0797523|T201|COMP|14343-8|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0797524|T201|COMP|14344-6|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0797525|T201|COMP|14345-3|LNC|Specific gravity|Specific gravity
C0797526|T201|COMP|14346-1|LNC|Specific gravity|Specific gravity
C0797527|T201|COMP|14347-9|LNC|Specific gravity|Specific gravity
C0797528|T201|COMP|14348-7|LNC|Specific gravity|Specific gravity
C0797529|T201|COMP|14349-5|LNC|Specific gravity|Specific gravity
C0797530|T201|COMP|14350-3|LNC|Specific gravity|Specific gravity
C0797531|T201|COMP|14351-1|LNC|Specific gravity|Specific gravity
C0797532|T201|COMP|14352-9|LNC|Specific gravity|Specific gravity
C0797546|T201|COMP|14366-9|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C0797547|T201|COMP|14367-7|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C0797548|T201|COMP|14368-5|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C0797549|T201|COMP|14369-3|LNC|Yeast|Yeast
C0797550|T201|COMP|14370-1|LNC|Yeast|Yeast
C0797551|T201|COMP|14371-9|LNC|Yeast|Yeast
C0797552|T201|COMP|14372-7|LNC|Erythrocytes|Erythrocytes
C0797553|T201|COMP|14373-5|LNC|Leukocytes|Leukocytes
C0797554|T201|COMP|14374-3|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0797555|T201|COMP|14375-0|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0797556|T201|COMP|14376-8|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0797557|T201|COMP|14377-6|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0797558|T201|COMP|14378-4|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0797559|T201|COMP|14379-2|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0797560|T201|COMP|14380-0|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0797561|T201|COMP|14381-8|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0797562|T201|COMP|14382-6|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0797563|T201|COMP|14383-4|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0797564|T201|COMP|14384-2|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0797565|T201|COMP|14385-9|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0797566|T201|COMP|14386-7|LNC|Glucose|Glucose
C0797567|T201|COMP|14387-5|LNC|Protein|Protein
C0797568|T201|COMP|14388-3|LNC|Amylase|Amylase
C0797569|T201|COMP|14389-1|LNC|Amylase|Amylase
C0797570|T201|COMP|14390-9|LNC|Amylase|Amylase
C0797571|T201|COMP|14391-7|LNC|Amylase|Amylase
C0797572|T201|COMP|14392-5|LNC|Amylase|Amylase
C0797573|T201|COMP|14393-3|LNC|Urea nitrogen|Urea nitrogen
C0797574|T201|COMP|14394-1|LNC|Urea nitrogen|Urea nitrogen
C0797575|T201|COMP|14396-6|LNC|Urea nitrogen|Urea nitrogen
C0797576|T201|COMP|14397-4|LNC|Urea nitrogen|Urea nitrogen
C0797577|T201|COMP|14398-2|LNC|Creatinine|Creatinine
C0797578|T201|COMP|14399-0|LNC|Creatinine|Creatinine
C0797579|T201|COMP|14401-4|LNC|Creatinine|Creatinine
C0797580|T201|COMP|14402-2|LNC|Creatinine|Creatinine
C0797581|T201|COMP|14403-0|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0797582|T201|COMP|14404-8|LNC|Phosphate|Phosphate
C0797583|T201|COMP|14405-5|LNC|Phosphate|Phosphate
C0797584|T201|COMP|14406-3|LNC|Phosphate|Phosphate
C0797585|T201|COMP|14407-1|LNC|Phosphate|Phosphate
C0797586|T201|COMP|14408-9|LNC|Phosphate|Phosphate
C0797587|T201|COMP|14409-7|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0797588|T201|COMP|14410-5|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0797589|T201|COMP|14411-3|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0797590|T201|COMP|14412-1|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0797591|T201|COMP|14413-9|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0797592|T201|COMP|14414-7|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0797593|T201|COMP|14415-4|LNC|Calcium|Calcium
C0797594|T201|COMP|14416-2|LNC|Calcium|Calcium
C0797595|T201|COMP|14417-0|LNC|Calcium|Calcium
C0797596|T201|COMP|14418-8|LNC|Calcium|Calcium
C0797597|T201|COMP|14419-6|LNC|Calcium|Calcium
C0797598|T201|COMP|14420-4|LNC|Bilirubin|Bilirubin
C0797599|T201|COMP|14421-2|LNC|Bilirubin|Bilirubin
C0797600|T201|COMP|14422-0|LNC|Bilirubin|Bilirubin
C0797601|T201|COMP|14423-8|LNC|Bilirubin|Bilirubin
C0797602|T201|COMP|14424-6|LNC|Bilirubin|Bilirubin
C0797603|T201|COMP|14425-3|LNC|Globulin|Globulin
C0797604|T201|COMP|14426-1|LNC|Globulin|Globulin
C0797605|T201|COMP|14427-9|LNC|Globulin|Globulin
C0797606|T201|COMP|14428-7|LNC|Globulin|Globulin
C0797607|T201|COMP|14429-5|LNC|Globulin|Globulin
C0797608|T201|COMP|14430-3|LNC|Globulin|Globulin
C0797609|T201|COMP|14431-1|LNC|Globulin|Globulin
C0797610|T201|COMP|14432-9|LNC|Albumin/Globulin|Albumin/Globulin
C0797611|T201|COMP|14433-7|LNC|Albumin/Globulin|Albumin/Globulin
C0797612|T201|COMP|14434-5|LNC|Albumin/Globulin|Albumin/Globulin
C0797613|T201|COMP|14435-2|LNC|Albumin/Globulin|Albumin/Globulin
C0797614|T201|COMP|14436-0|LNC|Albumin/Globulin|Albumin/Globulin
C0797615|T201|COMP|14437-8|LNC|Albumin/Globulin|Albumin/Globulin
C0797616|T201|COMP|14438-6|LNC|Cholesterol|Cholesterol
C0797617|T201|COMP|14439-4|LNC|Cholesterol|Cholesterol
C0797618|T201|COMP|14441-0|LNC|Cholesterol|Cholesterol
C0797619|T201|COMP|14442-8|LNC|Cholesterol|Cholesterol
C0797620|T201|COMP|14443-6|LNC|Cholesterol|Cholesterol
C0797621|T201|COMP|14444-4|LNC|Cholesterol|Cholesterol
C0797622|T201|COMP|14445-1|LNC|Triglyceride|Triglyceride
C0797623|T201|COMP|14446-9|LNC|Triglyceride|Triglyceride
C0797624|T201|COMP|14447-7|LNC|Triglyceride|Triglyceride
C0797625|T201|COMP|14448-5|LNC|Triglyceride|Triglyceride
C0797626|T201|COMP|14449-3|LNC|Triglyceride|Triglyceride
C0797627|T201|COMP|14450-1|LNC|Triglyceride|Triglyceride
C0797628|T201|COMP|14451-9|LNC|Virus identified|Virus identified
C0797629|T201|COMP|14452-7|LNC|Virus identified|Virus identified
C0797630|T201|COMP|14453-5|LNC|Virus identified|Virus identified
C0797631|T201|COMP|14454-3|LNC|Virus identified|Virus identified
C0797632|T201|COMP|14455-0|LNC|Virus identified|Virus identified
C0797633|T201|COMP|14456-8|LNC|Virus identified|Virus identified
C0797634|T201|COMP|14457-6|LNC|Virus identified|Virus identified
C0797635|T201|COMP|14458-4|LNC|Virus identified|Virus identified
C0797636|T201|COMP|14459-2|LNC|Virus identified|Virus identified
C0797637|T201|COMP|14460-0|LNC|Virus identified|Virus identified
C0797638|T201|COMP|14461-8|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C0797639|T201|COMP|14462-6|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C0797640|T201|COMP|14463-4|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C0797641|T201|COMP|14464-2|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C0797642|T201|COMP|14465-9|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C0797643|T201|COMP|14466-7|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C0797644|T201|COMP|14467-5|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C0797645|T201|COMP|14468-3|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797646|T201|COMP|14469-1|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797647|T201|COMP|14470-9|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797648|T201|COMP|14471-7|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797649|T201|COMP|14472-5|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797650|T201|COMP|14473-3|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797651|T201|COMP|14474-1|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797652|T201|COMP|14475-8|LNC|Bacteria identified|Bacteria identified
C0797653|T201|COMP|14477-4|LNC|Bacteria identified|Bacteria identified
C0797654|T201|COMP|14478-2|LNC|Bacteria identified|Bacteria identified
C0797655|T201|COMP|14479-0|LNC|Diphtheria sp identified|Diphtheria sp identified
C0797656|T201|COMP|14480-8|LNC|Diphtheria sp identified|Diphtheria sp identified
C0797657|T201|COMP|14481-6|LNC|Diphtheria sp identified|Diphtheria sp identified
C0797658|T201|COMP|14482-4|LNC|Diphtheria sp identified|Diphtheria sp identified
C0797659|T201|COMP|14483-2|LNC|Diphtheria sp identified|Diphtheria sp identified
C0797660|T201|COMP|14484-0|LNC|Mycoplasma sp & Ureaplasma sp|Mycoplasma sp & Ureaplasma sp
C0797661|T201|COMP|14485-7|LNC|Mycoplasma sp & Ureaplasma sp|Mycoplasma sp & Ureaplasma sp
C0797662|T201|COMP|14486-5|LNC|Mycoplasma sp & Ureaplasma sp|Mycoplasma sp & Ureaplasma sp
C0797663|T201|COMP|14487-3|LNC|Mycoplasma sp & Ureaplasma sp|Mycoplasma sp & Ureaplasma sp
C0797664|T201|COMP|14488-1|LNC|Virus identified|Virus identified
C0797665|T201|COMP|14489-9|LNC|Virus identified|Virus identified
C0797666|T201|COMP|14490-7|LNC|Virus identified|Virus identified
C0797667|T201|COMP|14491-5|LNC|Virus identified|Virus identified
C0797668|T201|COMP|14492-3|LNC|Virus identified|Virus identified
C0797669|T201|COMP|14493-1|LNC|Virus identified|Virus identified
C0797670|T201|COMP|14494-9|LNC|Virus identified|Virus identified
C0797671|T201|COMP|14495-6|LNC|Virus identified|Virus identified
C0797672|T201|COMP|14496-4|LNC|Virus identified|Virus identified
C0797673|T201|COMP|14497-2|LNC|Virus identified|Virus identified
C0797674|T201|COMP|14498-0|LNC|Virus identified|Virus identified
C0797675|T201|COMP|14499-8|LNC|Human papilloma virus Ag|Human papilloma virus Ag
C0797676|T201|COMP|14500-3|LNC|Human papilloma virus Ag|Human papilloma virus Ag
C0797677|T201|COMP|14501-1|LNC|Human papilloma virus Ag|Human papilloma virus Ag
C0797678|T201|COMP|14502-9|LNC|Human papilloma virus Ag|Human papilloma virus Ag
C0797679|T201|COMP|14503-7|LNC|Human papilloma virus 16+18 Ag|Human papilloma virus 16+18 Ag
C0797680|T201|COMP|14504-5|LNC|Human papilloma virus 16+18 Ag|Human papilloma virus 16+18 Ag
C0797681|T201|COMP|14505-2|LNC|Human papilloma virus 16+18 Ag|Human papilloma virus 16+18 Ag
C0797682|T201|COMP|14506-0|LNC|Human papilloma virus 16+18 Ag|Human papilloma virus 16+18 Ag
C0797683|T201|COMP|14507-8|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797684|T201|COMP|14508-6|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797685|T201|COMP|14509-4|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797686|T201|COMP|14510-2|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797687|T201|COMP|14511-0|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797688|T201|COMP|14512-8|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797689|T201|COMP|14513-6|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C0797690|T201|COMP|14514-4|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0797691|T201|COMP|14515-1|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0797692|T201|COMP|14516-9|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0797693|T201|COMP|14517-7|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0797694|T201|COMP|14518-5|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0797695|T201|COMP|14519-3|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0797696|T201|COMP|14520-1|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0797697|T201|COMP|14521-9|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0797698|T201|COMP|14522-7|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C0797699|T201|COMP|14523-5|LNC|Rubella virus Ag|Rubella virus Ag
C0797700|T201|COMP|14524-3|LNC|Rubella virus Ag|Rubella virus Ag
C0797701|T201|COMP|14525-0|LNC|Rubella virus Ag|Rubella virus Ag
C0797702|T201|COMP|14526-8|LNC|Rubella virus Ag|Rubella virus Ag
C0797703|T201|COMP|14527-6|LNC|Rubella virus Ag|Rubella virus Ag
C0797704|T201|COMP|14528-4|LNC|Rubella virus Ag|Rubella virus Ag
C0797705|T201|COMP|14529-2|LNC|Rubella virus Ag|Rubella virus Ag
C0797706|T201|COMP|14530-0|LNC|Rubella virus Ag|Rubella virus Ag
C0797707|T201|COMP|14531-8|LNC|Rubella virus Ag|Rubella virus Ag
C0797708|T201|COMP|14532-6|LNC|Rubella virus Ag|Rubella virus Ag
C0797709|T201|COMP|14533-4|LNC|Rubella virus Ag|Rubella virus Ag
C0797710|T201|COMP|14534-2|LNC|Measles virus Ag|Measles virus Ag
C0797711|T201|COMP|14535-9|LNC|Measles virus Ag|Measles virus Ag
C0797712|T201|COMP|14536-7|LNC|Measles virus Ag|Measles virus Ag
C0797713|T201|COMP|14537-5|LNC|Measles virus Ag|Measles virus Ag
C0797714|T201|COMP|14538-3|LNC|Measles virus Ag|Measles virus Ag
C0797715|T201|COMP|14539-1|LNC|Measles virus Ag|Measles virus Ag
C0797716|T201|COMP|14540-9|LNC|Measles virus Ag|Measles virus Ag
C0797717|T201|COMP|14541-7|LNC|Measles virus Ag|Measles virus Ag
C0797718|T201|COMP|14542-5|LNC|Measles virus Ag|Measles virus Ag
C0797719|T201|COMP|14543-3|LNC|Measles virus Ag|Measles virus Ag
C0797720|T201|COMP|14544-1|LNC|Measles virus Ag|Measles virus Ag
C0797721|T201|COMP|14545-8|LNC|Mumps virus Ag|Mumps virus Ag
C0797722|T201|COMP|14546-6|LNC|Mumps virus Ag|Mumps virus Ag
C0797723|T201|COMP|14547-4|LNC|Mumps virus Ag|Mumps virus Ag
C0797724|T201|COMP|14548-2|LNC|Mumps virus Ag|Mumps virus Ag
C0797725|T201|COMP|14549-0|LNC|Mumps virus Ag|Mumps virus Ag
C0797726|T201|COMP|14550-8|LNC|Mumps virus Ag|Mumps virus Ag
C0797727|T201|COMP|14551-6|LNC|Mumps virus Ag|Mumps virus Ag
C0797728|T201|COMP|14552-4|LNC|Mumps virus Ag|Mumps virus Ag
C0797729|T201|COMP|14553-2|LNC|Mumps virus Ag|Mumps virus Ag
C0797730|T201|COMP|14554-0|LNC|Mumps virus Ag|Mumps virus Ag
C0797731|T201|COMP|14555-7|LNC|Mumps virus Ag|Mumps virus Ag
C0797732|T201|COMP|14556-5|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C0797733|T201|COMP|14557-3|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C0797734|T201|COMP|14558-1|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C0797735|T201|COMP|14559-9|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C0797736|T201|COMP|14560-7|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C0797737|T201|COMP|14561-5|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C0797738|T201|COMP|14562-3|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C0797739|T201|COMP|14563-1|LNC|Hemoglobin.gastrointestinal^1st specimen|Hemoglobin.gastrointestinal^1st specimen
C0797740|T201|COMP|14564-9|LNC|Hemoglobin.gastrointestinal^2nd specimen|Hemoglobin.gastrointestinal^2nd specimen
C0797741|T201|COMP|14565-6|LNC|Hemoglobin.gastrointestinal^3rd specimen|Hemoglobin.gastrointestinal^3rd specimen
C0797742|T201|COMP|14566-4|LNC|Calcitriol|Calcitriol
C0797743|T201|COMP|14567-2|LNC|11-Deoxycortisol|11-Deoxycortisol
C0797744|T201|COMP|14568-0|LNC|17-Hydroxycorticosteroids|17-Hydroxycorticosteroids
C0797745|T201|COMP|14569-8|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C0797746|T201|COMP|14570-6|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C0797747|T201|COMP|14571-4|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C0797748|T201|COMP|14572-2|LNC|17-Ketosteroids|17-Ketosteroids
C0797749|T201|COMP|14573-0|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C0797750|T201|COMP|14574-8|LNC|8-Hydroxyamoxapine|8-Hydroxyamoxapine
C0797751|T201|COMP|14575-5|LNC|Blood group antibody investigation|Blood group antibody investigation
C0797752|T201|COMP|14576-3|LNC|Blood group antibody investigation|Blood group antibody investigation
C0797753|T201|COMP|14577-1|LNC|ABO & Rh group|ABO & Rh group
C0797754|T201|COMP|14578-9|LNC|ABO group|ABO group
C0797755|T201|COMP|14579-7|LNC|ABO group|ABO group
C0797756|T201|COMP|14580-5|LNC|ABO group|ABO group
C0797757|T201|COMP|14581-3|LNC|Acetaminophen|Acetaminophen
C0797758|T201|COMP|14582-1|LNC|Acetone|Acetone
C0797759|T201|COMP|14583-9|LNC|Acidity.titratable|Acidity.titratable
C0797760|T201|COMP|14584-7|LNC|Adenosine monophosphate.cyclic|Adenosine monophosphate.cyclic
C0797761|T201|COMP|14585-4|LNC|Albumin/Creatinine|Albumin/Creatinine
C0797762|T201|COMP|14586-2|LNC|Aldosterone|Aldosterone
C0797763|T201|COMP|14587-0|LNC|Aldosterone|Aldosterone
C0797764|T201|COMP|14588-8|LNC|Alkaline phosphatase isoenzymes|Alkaline phosphatase isoenzymes
C0797765|T201|COMP|14589-6|LNC|Amylase isoenzymes|Amylase isoenzymes
C0797766|T201|COMP|14590-4|LNC|Alpha tocopherol|Alpha tocopherol
C0797767|T201|COMP|14591-2|LNC|ALPRAZolam|ALPRAZolam
C0797768|T201|COMP|14592-0|LNC|Aluminum|Aluminum
C0797769|T201|COMP|14593-8|LNC|Aluminum|Aluminum
C0797770|T201|COMP|14594-6|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C0797771|T201|COMP|14595-3|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C0797772|T201|COMP|14596-1|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C0797773|T201|COMP|14597-9|LNC|Amitriptyline|Amitriptyline
C0797774|T201|COMP|14598-7|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C0797775|T201|COMP|14599-5|LNC|Ammonium|Ammonium
C0797776|T201|COMP|14600-1|LNC|Amoxapine|Amoxapine
C0797777|T201|COMP|14601-9|LNC|Amoxapine+8-Hydroxyamoxapine|Amoxapine+8-Hydroxyamoxapine
C0797778|T201|COMP|14603-5|LNC|Androstenedione|Androstenedione
C0797779|T201|COMP|14604-3|LNC|Blood group antibodies identified|Blood group antibodies identified
C0797780|T201|COMP|14605-0|LNC|Blood group antibodies identified|Blood group antibodies identified
C0797781|T201|COMP|14606-8|LNC|Blood group antibody screen|Blood group antibody screen
C0797782|T201|COMP|14607-6|LNC|Nuclear Ab|Nuclear Ab
C0797783|T201|COMP|14608-4|LNC|Nuclear Ab|Nuclear Ab
C0797784|T201|COMP|14609-2|LNC|Nuclear Ab|Nuclear Ab
C0797785|T201|COMP|14610-0|LNC|Nuclear Ab|Nuclear Ab
C0797786|T201|COMP|14611-8|LNC|Nuclear Ab pattern|Nuclear Ab pattern
C0797787|T201|COMP|14612-6|LNC|Nuclear Ab|Nuclear Ab
C0797788|T201|COMP|14613-4|LNC|Nuclear Ab|Nuclear Ab
C0797789|T201|COMP|14614-2|LNC|Nuclear Ab|Nuclear Ab
C0797790|T201|COMP|14615-9|LNC|Nuclear Ab|Nuclear Ab
C0797791|T201|COMP|14616-7|LNC|Nuclear Ab|Nuclear Ab
C0797792|T201|COMP|14617-5|LNC|Appearance|Appearance
C0797793|T201|COMP|14618-3|LNC|Appearance|Appearance
C0797794|T201|COMP|14619-1|LNC|Appearance|Appearance
C0797795|T201|COMP|14620-9|LNC|Appearance|Appearance
C0797796|T201|COMP|14621-7|LNC|Appearance|Appearance
C0797797|T201|COMP|14622-5|LNC|Ascorbate|Ascorbate
C0797798|T201|COMP|14623-3|LNC|Barbital|Barbital
C0797799|T201|COMP|14624-1|LNC|Barbiturates|Barbiturates
C0797800|T201|COMP|14625-8|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0797801|T201|COMP|14626-6|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C0797802|T201|COMP|14627-4|LNC|Bicarbonate|Bicarbonate
C0797803|T201|COMP|14628-2|LNC|Bile acid|Bile acid
C0797804|T201|COMP|14629-0|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C0797805|T201|COMP|14630-8|LNC|Bilirubin.non-glucuronidated|Bilirubin.non-glucuronidated
C0797806|T201|COMP|14631-6|LNC|Bilirubin|Bilirubin
C0797807|T201|COMP|14632-4|LNC|Buffy coat|Buffy coat
C0797808|T201|COMP|14633-2|LNC|C peptide|C peptide
C0797809|T201|COMP|14634-0|LNC|C reactive protein|C reactive protein
C0797810|T201|COMP|14635-7|LNC|Calcidiol|Calcidiol
C0797811|T201|COMP|14636-5|LNC|Calcium|Calcium
C0797812|T201|COMP|14637-3|LNC|Calcium|Calcium
C0797814|T201|COMP|14639-9|LNC|carBAMazepine|carBAMazepine
C0797815|T201|COMP|14640-7|LNC|Carbon dioxide|Carbon dioxide
C0797816|T201|COMP|14641-5|LNC|Carbonate|Carbonate
C0797817|T201|COMP|14642-3|LNC|Carotene|Carotene
C0797818|T201|COMP|14643-1|LNC|Catecholamines.free|Catecholamines.free
C0797819|T201|COMP|14644-9|LNC|chlorproMAZINE|chlorproMAZINE
C0797820|T201|COMP|14645-6|LNC|chlorproMAZINE|chlorproMAZINE
C0797821|T201|COMP|14646-4|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C0797822|T201|COMP|14647-2|LNC|Cholesterol|Cholesterol
C0797823|T201|COMP|14648-0|LNC|Chylomicrons|Chylomicrons
C0797824|T201|COMP|14649-8|LNC|Cimetidine|Cimetidine
C0797825|T201|COMP|14650-6|LNC|Citrate|Citrate
C0797826|T201|COMP|14651-4|LNC|cloBAZam|cloBAZam
C0797827|T201|COMP|14652-2|LNC|clomiPRAMINE|clomiPRAMINE
C0797828|T201|COMP|14653-0|LNC|clomiPRAMINE|clomiPRAMINE
C0797829|T201|COMP|14654-8|LNC|Clomipramine+Norclomipramine|Clomipramine+Norclomipramine
C0797830|T201|COMP|14655-5|LNC|clonazePAM|clonazePAM
C0797831|T201|COMP|14656-3|LNC|cloZAPine|cloZAPine
C0797832|T201|COMP|14657-1|LNC|Clozapine+Norclozapine|Clozapine+Norclozapine
C0797833|T201|COMP|14658-9|LNC|Cold agglutinin|Cold agglutinin
C0797834|T201|COMP|14660-5|LNC|Color|Color
C0797835|T201|COMP|14661-3|LNC|Color|Color
C0797836|T201|COMP|14662-1|LNC|Color|Color
C0797837|T201|COMP|14663-9|LNC|Color|Color
C0797838|T201|COMP|14664-7|LNC|Color|Color
C0797839|T201|COMP|14665-4|LNC|Copper|Copper
C0797840|T201|COMP|14666-2|LNC|Copper|Copper
C0797841|T201|COMP|14667-0|LNC|Coproporphyrin 1|Coproporphyrin 1
C0797842|T201|COMP|14668-8|LNC|Coproporphyrin 1|Coproporphyrin 1
C0797843|T201|COMP|14669-6|LNC|Coproporphyrin 1|Coproporphyrin 1
C0797844|T201|COMP|14670-4|LNC|Coproporphyrin 1/Porphyrins.total|Coproporphyrin 1/Porphyrins.total
C0797845|T201|COMP|14671-2|LNC|Coproporphyrin 3|Coproporphyrin 3
C0797846|T201|COMP|14672-0|LNC|Coproporphyrin 3|Coproporphyrin 3
C0797847|T201|COMP|14673-8|LNC|Coproporphyrin 3|Coproporphyrin 3
C0797848|T201|COMP|14674-6|LNC|Corticotropin|Corticotropin
C0797849|T201|COMP|14675-3|LNC|Cortisol|Cortisol
C0797850|T201|COMP|14676-1|LNC|Cortisol.free|Cortisol.free
C0797852|T201|COMP|14678-7|LNC|Cortisol^PM trough specimen|Cortisol^PM trough specimen
C0797853|T201|COMP|14679-5|LNC|Cortisol^AM peak specimen|Cortisol^AM peak specimen
C0797854|T201|COMP|14680-3|LNC|Creatine kinase isoenzymes|Creatine kinase isoenzymes
C0797855|T201|COMP|14681-1|LNC|Creatinine|Creatinine
C0797856|T201|COMP|14682-9|LNC|Creatinine|Creatinine
C0797857|T201|COMP|14683-7|LNC|Creatinine|Creatinine
C0797858|T201|COMP|14684-5|LNC|Creatinine|Creatinine
C0797859|T201|COMP|14685-2|LNC|Cobalamins|Cobalamins
C0797860|T201|COMP|14686-0|LNC|Cystine|Cystine
C0797861|T201|COMP|14687-8|LNC|Transfusion date|Transfusion date
C0797862|T201|COMP|14688-6|LNC|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C0797863|T201|COMP|14689-4|LNC|Delta aminolevulinate|Delta aminolevulinate
C0797864|T201|COMP|14690-2|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0797865|T201|COMP|14691-0|LNC|Desipramine|Desipramine
C0797866|T201|COMP|14692-8|LNC|Desipramine|Desipramine
C0797867|T201|COMP|14693-6|LNC|Norclobazam|Norclobazam
C0797868|T201|COMP|14694-4|LNC|Norclomipramine|Norclomipramine
C0797869|T201|COMP|14695-1|LNC|Nordoxepin|Nordoxepin
C0797870|T201|COMP|14696-9|LNC|Deuteroporphyrin|Deuteroporphyrin
C0797871|T201|COMP|14697-7|LNC|diazePAM|diazePAM
C0797872|T201|COMP|14698-5|LNC|Digoxin|Digoxin
C0797873|T201|COMP|14699-3|LNC|diphenhydrAMINE+Dimenhydrinate|diphenhydrAMINE+Dimenhydrinate
C0797874|T201|COMP|14700-9|LNC|diphenhydrAMINE+Dimenhydrinate|diphenhydrAMINE+Dimenhydrinate
C0797875|T201|COMP|14701-7|LNC|diphenhydrAMINE+Dimenhydrinate|diphenhydrAMINE+Dimenhydrinate
C0797876|T201|COMP|14702-5|LNC|Disopyramide|Disopyramide
C0797877|T201|COMP|14703-3|LNC|DOPamine|DOPamine
C0797878|T201|COMP|14704-1|LNC|Doxepin|Doxepin
C0797879|T201|COMP|14705-8|LNC|Doxepin|Doxepin
C0797880|T201|COMP|14706-6|LNC|Doxepin|Doxepin
C0797881|T201|COMP|14707-4|LNC|Doxepin+Nordoxepin|Doxepin+Nordoxepin
C0797882|T201|COMP|14708-2|LNC|Endomysium Ab|Endomysium Ab
C0797883|T201|COMP|14709-0|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0797884|T201|COMP|14710-8|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C0797885|T201|COMP|14711-6|LNC|EPINEPHrine|EPINEPHrine
C0797886|T201|COMP|14712-4|LNC|EPINEPHrine|EPINEPHrine
C0797887|T201|COMP|14713-2|LNC|Erythrocytes|Erythrocytes
C0797888|T201|COMP|14714-0|LNC|Erythropoietin|Erythropoietin
C0797889|T201|COMP|14715-7|LNC|Estradiol|Estradiol
C0797890|T201|COMP|14716-5|LNC|Estriol|Estriol
C0797891|T201|COMP|14717-3|LNC|Estriol|Estriol
C0797892|T201|COMP|14718-1|LNC|Estriol|Estriol
C0797893|T201|COMP|14719-9|LNC|Ethanol|Ethanol
C0797894|T201|COMP|14720-7|LNC|Ethosuximide|Ethosuximide
C0797895|T201|COMP|14721-5|LNC|Ethylene glycol|Ethylene glycol
C0797896|T201|COMP|14722-3|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C0797897|T201|COMP|14723-1|LNC|Ferritin|Ferritin
C0797898|T201|COMP|14724-9|LNC|Ferritin|Ferritin
C0797899|T201|COMP|14725-6|LNC|Fluid|Fluid
C0797900|T201|COMP|14726-4|LNC|Fluoride|Fluoride
C0797901|T201|COMP|14727-2|LNC|FLUoxetine|FLUoxetine
C0797902|T201|COMP|14728-0|LNC|FLUoxetine|FLUoxetine
C0797903|T201|COMP|14729-8|LNC|Flurazepam|Flurazepam
C0797904|T201|COMP|14730-6|LNC|Flurazepam+N-desalkylflurazepam|Flurazepam+N-desalkylflurazepam
C0797905|T201|COMP|14731-4|LNC|Folate|Folate
C0797906|T201|COMP|14732-2|LNC|Folate|Folate
C0797907|T201|COMP|14733-0|LNC|Folate+Cyanocobalamin|Folate+Cyanocobalamin
C0797908|T201|COMP|14734-8|LNC|Follitropin|Follitropin
C0797909|T201|COMP|14735-5|LNC|Gastrin^10M post 0.2 U/kg secretin|Gastrin^10M post 0.2 U/kg secretin
C0797910|T201|COMP|14736-3|LNC|Gastrin^15M post 0.2 U/kg secretin|Gastrin^15M post 0.2 U/kg secretin
C0797911|T201|COMP|14737-1|LNC|Gastrin^20M post 0.2 U/kg secretin|Gastrin^20M post 0.2 U/kg secretin
C0797912|T201|COMP|14738-9|LNC|Gastrin^25M post 0.2 U/kg secretin|Gastrin^25M post 0.2 U/kg secretin
C0797913|T201|COMP|14739-7|LNC|Gastrin^2M post 0.2 U/kg secretin|Gastrin^2M post 0.2 U/kg secretin
C0797914|T201|COMP|14740-5|LNC|Gastrin^30M post 0.2 U/kg secretin|Gastrin^30M post 0.2 U/kg secretin
C0797915|T201|COMP|14741-3|LNC|Gastrin^5M post 0.2 U/kg secretin|Gastrin^5M post 0.2 U/kg secretin
C0797916|T201|COMP|14742-1|LNC|Gastrin^pre 0.2 U/kg secretin|Gastrin^pre 0.2 U/kg secretin
C0797917|T201|COMP|14743-9|LNC|Glucose|Glucose
C0797918|T201|COMP|14744-7|LNC|Glucose|Glucose
C0797919|T201|COMP|14745-4|LNC|Glucose|Glucose
C0797920|T201|COMP|14746-2|LNC|Glucose|Glucose
C0797921|T201|COMP|14747-0|LNC|Glucose|Glucose
C0797922|T201|COMP|14748-8|LNC|Glucose|Glucose
C0797923|T201|COMP|14749-6|LNC|Glucose|Glucose
C0797924|T201|COMP|14750-4|LNC|Glucose|Glucose
C0797925|T201|COMP|14751-2|LNC|Glucose^1.5H post 50 g lactose PO|Glucose^1.5H post 50 g lactose PO
C0797926|T201|COMP|14752-0|LNC|Glucose^1.5H post dose glucose|Glucose^1.5H post dose glucose
C0797927|T201|COMP|14753-8|LNC|Glucose^1H post 100 g glucose PO|Glucose^1H post 100 g glucose PO
C0797928|T201|COMP|14754-6|LNC|Glucose^1H post 50 g glucose PO|Glucose^1H post 50 g glucose PO
C0797929|T201|COMP|14755-3|LNC|Glucose^1H post 50 g lactose PO|Glucose^1H post 50 g lactose PO
C0797930|T201|COMP|14756-1|LNC|Glucose^1H post dose glucose|Glucose^1H post dose glucose
C0797931|T201|COMP|14757-9|LNC|Glucose^2H post 100 g glucose PO|Glucose^2H post 100 g glucose PO
C0797932|T201|COMP|14758-7|LNC|Glucose^2H post 50 g lactose PO|Glucose^2H post 50 g lactose PO
C0797933|T201|COMP|14759-5|LNC|Glucose^2H post dose glucose|Glucose^2H post dose glucose
C0797934|T201|COMP|14760-3|LNC|Glucose^2H post meal|Glucose^2H post meal
C0797935|T201|COMP|14761-1|LNC|Glucose^2H post meal|Glucose^2H post meal
C0797936|T201|COMP|14762-9|LNC|Glucose^30M post 50 g lactose PO|Glucose^30M post 50 g lactose PO
C0797937|T201|COMP|14763-7|LNC|Glucose^30M post dose glucose|Glucose^30M post dose glucose
C0797938|T201|COMP|14764-5|LNC|Glucose^3H post 100 g glucose PO|Glucose^3H post 100 g glucose PO
C0797939|T201|COMP|14765-2|LNC|Glucose^3H post dose glucose|Glucose^3H post dose glucose
C0797940|T201|COMP|14766-0|LNC|Glucose^4H post dose glucose|Glucose^4H post dose glucose
C0797941|T201|COMP|14767-8|LNC|Glucose^5H post dose glucose|Glucose^5H post dose glucose
C0797942|T201|COMP|14768-6|LNC|Glucose^baseline|Glucose^baseline
C0797943|T201|COMP|14769-4|LNC|Glucose^pre 12H CFst|Glucose^pre 12H CFst
C0797944|T201|COMP|14770-2|LNC|Glucose^post CFst|Glucose^post CFst
C0797945|T201|COMP|14771-0|LNC|Glucose^post CFst|Glucose^post CFst
C0797946|T201|COMP|14772-8|LNC|Gold|Gold
C0797947|T201|COMP|14773-6|LNC|Granulocytes/100 leukocytes|Granulocytes/100 leukocytes
C0797948|T201|COMP|14774-4|LNC|Haloperidol|Haloperidol
C0797949|T201|COMP|14775-1|LNC|Hemoglobin|Hemoglobin
C0797950|T201|COMP|14776-9|LNC|Heptacarboxylate|Heptacarboxylate
C0797951|T201|COMP|14777-7|LNC|Heptacarboxylate|Heptacarboxylate
C0797952|T201|COMP|14778-5|LNC|Heptacarboxylate|Heptacarboxylate
C0797953|T201|COMP|14779-3|LNC|Hexacarboxylate|Hexacarboxylate
C0797954|T201|COMP|14780-1|LNC|Hexacarboxylate|Hexacarboxylate
C0797955|T201|COMP|14781-9|LNC|Hexacarboxylate|Hexacarboxylate
C0797956|T201|COMP|14782-7|LNC|Homovanillate|Homovanillate
C0797957|T201|COMP|14783-5|LNC|Homovanillate|Homovanillate
C0797958|T201|COMP|14784-3|LNC|Hydroxyproline.free|Hydroxyproline.free
C0797959|T201|COMP|14785-0|LNC|Hydroxyproline|Hydroxyproline
C0797960|T201|COMP|14786-8|LNC|Arthropod identified|Arthropod identified
C0797961|T201|COMP|14787-6|LNC|Arthropod identified|Arthropod identified
C0797962|T201|COMP|14788-4|LNC|Helminth+Arthropod identified|Helminth+Arthropod identified
C0797963|T201|COMP|14789-2|LNC|Helminth identified|Helminth identified
C0797964|T201|COMP|14790-0|LNC|Helminth identified|Helminth identified
C0797965|T201|COMP|14791-8|LNC|Imipramine+Desipramine|Imipramine+Desipramine
C0797966|T201|COMP|14792-6|LNC|Imipramine+Desipramine|Imipramine+Desipramine
C0797967|T201|COMP|14793-4|LNC|Imipramine+Desipramine|Imipramine+Desipramine
C0797968|T201|COMP|14794-2|LNC|Imipramine+Desipramine|Imipramine+Desipramine
C0797969|T201|COMP|14795-9|LNC|Immunoglobulin light chains|Immunoglobulin light chains
C0797970|T201|COMP|14796-7|LNC|Insulin|Insulin
C0797971|T201|COMP|14797-5|LNC|Iron|Iron
C0797972|T201|COMP|14798-3|LNC|Iron|Iron
C0797973|T201|COMP|14799-1|LNC|Iron|Iron
C0797974|T201|COMP|14800-7|LNC|Iron binding capacity|Iron binding capacity
C0797975|T201|COMP|14801-5|LNC|Iron saturation|Iron saturation
C0797976|T201|COMP|14802-3|LNC|Isopropanol|Isopropanol
C0797977|T201|COMP|14803-1|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0797978|T201|COMP|14804-9|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0797979|T201|COMP|14805-6|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0797980|T201|COMP|14806-4|LNC|Lactose.PO|Lactose.PO
C0797981|T201|COMP|14807-2|LNC|Lead|Lead
C0797982|T201|COMP|14808-0|LNC|Lead|Lead
C0797983|T201|COMP|14809-8|LNC|Lead|Lead
C0797984|T201|COMP|14810-6|LNC|Leukocytes|Leukocytes
C0797985|T201|COMP|14811-4|LNC|Leukocytes|Leukocytes
C0797986|T201|COMP|14812-2|LNC|Lidocaine|Lidocaine
C0797987|T201|COMP|14813-0|LNC|Lipoprotein.alpha|Lipoprotein.alpha
C0797988|T201|COMP|14814-8|LNC|Lipoprotein.beta|Lipoprotein.beta
C0797989|T201|COMP|14815-5|LNC|Lipoprotein.beta|Lipoprotein.beta
C0797990|T201|COMP|14816-3|LNC|Lipoprotein.pre-beta|Lipoprotein.pre-beta
C0797991|T201|COMP|14817-1|LNC|LORazepam|LORazepam
C0797992|T201|COMP|14818-9|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0797993|T201|COMP|14819-7|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0797994|T201|COMP|14820-5|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0797995|T201|COMP|14821-3|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0797996|T201|COMP|32697-5|LNC|Lymphocytes|Lymphocytes
C0797997|T201|COMP|14823-9|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C0797998|T201|COMP|14824-7|LNC|Magnesium|Magnesium
C0797999|T201|COMP|14825-4|LNC|Maprotiline|Maprotiline
C0798000|T201|COMP|14826-2|LNC|Meperidine|Meperidine
C0798001|T201|COMP|14827-0|LNC|Mesoporphyrin|Mesoporphyrin
C0798002|T201|COMP|14828-8|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C0798003|T201|COMP|14829-6|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C0798004|T201|COMP|14830-4|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C0798005|T201|COMP|14831-2|LNC|Metanephrine/Creatinine|Metanephrine/Creatinine
C0798006|T201|COMP|34339-2|LNC|Metanephrine|Metanephrine
C0798007|T201|COMP|14833-8|LNC|Metanephrines|Metanephrines
C0798008|T201|COMP|14834-6|LNC|Methamphetamine|Methamphetamine
C0798009|T201|COMP|14835-3|LNC|Methanol|Methanol
C0798010|T201|COMP|14836-1|LNC|Methotrexate|Methotrexate
C0798011|T201|COMP|14837-9|LNC|Methsuximide|Methsuximide
C0798012|T201|COMP|14838-7|LNC|Toxoplasma gondii|Toxoplasma gondii
C0798013|T201|COMP|14839-5|LNC|Trypanosoma sp identified|Trypanosoma sp identified
C0798014|T201|COMP|14840-3|LNC|Trypanosoma sp identified|Trypanosoma sp identified
C0798017|T201|COMP|14843-7|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0798018|T201|COMP|14844-5|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0798019|T201|COMP|27073-6|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0798020|T201|COMP|14846-0|LNC|N-acetylprocainamide|N-acetylprocainamide
C0798021|T201|COMP|14847-8|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0798022|T201|COMP|14848-6|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0798023|T201|COMP|14849-4|LNC|Nitrazepam|Nitrazepam
C0798024|T201|COMP|14850-2|LNC|Nitrazepam|Nitrazepam
C0798025|T201|COMP|14851-0|LNC|Norclozapine|Norclozapine
C0798026|T201|COMP|14852-8|LNC|Norepinephrine|Norepinephrine
C0798027|T201|COMP|14853-6|LNC|Norepinephrine|Norepinephrine
C0798028|T201|COMP|14854-4|LNC|Norepinephrine|Norepinephrine
C0798029|T201|COMP|14855-1|LNC|Norfluoxetine|Norfluoxetine
C0798030|T201|COMP|14856-9|LNC|Nortriptyline|Nortriptyline
C0798031|T201|COMP|14857-7|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0798032|T201|COMP|14858-5|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0798033|T201|COMP|14859-3|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0798034|T201|COMP|14860-1|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0798035|T201|COMP|14861-9|LNC|Oxalate|Oxalate
C0798036|T201|COMP|14862-7|LNC|Oxalate|Oxalate
C0798037|T201|COMP|14863-5|LNC|oxyCODONE|oxyCODONE
C0798038|T201|COMP|14864-3|LNC|Oxygen|Oxygen
C0798039|T201|COMP|14865-0|LNC|Parathyrin|Parathyrin
C0798040|T201|COMP|14866-8|LNC|Parathyrin.intact|Parathyrin.intact
C0798041|T201|COMP|14867-6|LNC|PARoxetine|PARoxetine
C0798042|T201|COMP|14868-4|LNC|Pathologist report|Pathologist report
C0798043|T201|COMP|14869-2|LNC|Pathologist review|Pathologist review
C0798044|T201|COMP|14870-0|LNC|Pentacarboxylate|Pentacarboxylate
C0798045|T201|COMP|14871-8|LNC|Pentacarboxylate|Pentacarboxylate
C0798046|T201|COMP|14872-6|LNC|Pentacarboxylate|Pentacarboxylate
C0798048|T201|COMP|14874-2|LNC|PHENobarbital|PHENobarbital
C0798049|T201|COMP|14875-9|LNC|Phenylalanine|Phenylalanine
C0798050|T201|COMP|14876-7|LNC|Phenylpropanolamine|Phenylpropanolamine
C0798051|T201|COMP|14877-5|LNC|Phenytoin|Phenytoin
C0798052|T201|COMP|14878-3|LNC|Phosphate|Phosphate
C0798053|T201|COMP|14879-1|LNC|Phosphate|Phosphate
C0798055|T201|COMP|14881-7|LNC|Phosphate|Phosphate
C0798056|T201|COMP|14882-5|LNC|Porphobilinogen|Porphobilinogen
C0798057|T201|COMP|14883-3|LNC|Porphyrins|Porphyrins
C0798058|T201|COMP|14884-1|LNC|Porphyrins|Porphyrins
C0798059|T201|COMP|14885-8|LNC|Pregnanediol|Pregnanediol
C0798060|T201|COMP|14886-6|LNC|Pregnanetriol|Pregnanetriol
C0798061|T201|COMP|14887-4|LNC|Primidone|Primidone
C0798062|T201|COMP|14888-2|LNC|Procainamide|Procainamide
C0798063|T201|COMP|14889-0|LNC|Procainamide+N-acetylprocainamide|Procainamide+N-acetylprocainamide
C0798064|T201|COMP|14890-8|LNC|Progesterone|Progesterone
C0798065|T201|COMP|14891-6|LNC|Propranolol|Propranolol
C0798066|T201|COMP|14892-4|LNC|Propranolol|Propranolol
C0798067|T201|COMP|14893-2|LNC|Propranolol|Propranolol
C0798068|T201|COMP|14894-0|LNC|Propylene glycol|Propylene glycol
C0798069|T201|COMP|14895-7|LNC|Protein pattern|Protein pattern
C0798070|T201|COMP|14896-5|LNC|Protein pattern|Protein pattern
C0798071|T201|COMP|14898-1|LNC|Protriptyline|Protriptyline
C0798072|T201|COMP|14899-9|LNC|quiNIDine|quiNIDine
C0798073|T201|COMP|14900-5|LNC|raNITIdine|raNITIdine
C0798074|T201|COMP|14901-3|LNC|raNITIdine|raNITIdine
C0798075|T201|COMP|14902-1|LNC|raNITIdine|raNITIdine
C0798076|T201|COMP|14903-9|LNC|Folate|Folate
C0798077|T201|COMP|14904-7|LNC|Reagin Ab|Reagin Ab
C0798078|T201|COMP|14905-4|LNC|Retinol|Retinol
C0798079|T201|COMP|14906-2|LNC|Rh|Rh
C0798080|T201|COMP|14907-0|LNC|Rh|Rh
C0798081|T201|COMP|14908-8|LNC|Rh|Rh
C0798082|T201|COMP|14909-6|LNC|Salicylates|Salicylates
C0798083|T201|COMP|14910-4|LNC|Serotonin|Serotonin
C0798084|T201|COMP|14911-2|LNC|Sertraline|Sertraline
C0798085|T201|COMP|14912-0|LNC|Smudge cells/100 leukocytes|Smudge cells/100 leukocytes
C0798086|T201|COMP|14913-8|LNC|Testosterone|Testosterone
C0798087|T201|COMP|14914-6|LNC|Testosterone.free|Testosterone.free
C0798088|T201|COMP|14915-3|LNC|Theophylline|Theophylline
C0798089|T201|COMP|14916-1|LNC|Thiocyanate|Thiocyanate
C0798090|T201|COMP|14917-9|LNC|Thioridazine|Thioridazine
C0798091|T201|COMP|14918-7|LNC|Thyroglobulin|Thyroglobulin
C0798092|T201|COMP|14919-5|LNC|Thyrotropin binding inhibitory immunoglobulins|Thyrotropin binding inhibitory immunoglobulins
C0798093|T201|COMP|14920-3|LNC|Thyroxine.free|Thyroxine.free
C0798094|T201|COMP|14921-1|LNC|Thyroxine|Thyroxine
C0798095|T201|COMP|14922-9|LNC|Toxoplasma gondii Ab.IgA+IgE|Toxoplasma gondii Ab.IgA+IgE
C0798096|T201|COMP|14923-7|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C0798097|T201|COMP|14924-5|LNC|Transfusion reaction|Transfusion reaction
C0798098|T201|COMP|14925-2|LNC|traZODone|traZODone
C0798099|T201|COMP|14926-0|LNC|Triazolam|Triazolam
C0798100|T201|COMP|14927-8|LNC|Triglyceride|Triglyceride
C0798101|T201|COMP|14928-6|LNC|Triiodothyronine.free|Triiodothyronine.free
C0798102|T201|COMP|14929-4|LNC|Triiodothyronine.reverse|Triiodothyronine.reverse
C0798103|T201|COMP|14930-2|LNC|Triiodothyronine|Triiodothyronine
C0798104|T201|COMP|14931-0|LNC|Trimipramine|Trimipramine
C0798105|T201|COMP|14932-8|LNC|Urate|Urate
C0798106|T201|COMP|14933-6|LNC|Urate|Urate
C0798107|T201|COMP|14934-4|LNC|Urate|Urate
C0798108|T201|COMP|14935-1|LNC|Urate|Urate
C0798109|T201|COMP|14936-9|LNC|Urea nitrogen|Urea nitrogen
C0798110|T201|COMP|14937-7|LNC|Urea nitrogen|Urea nitrogen
C0798111|T201|COMP|14938-5|LNC|Urea nitrogen|Urea nitrogen
C0798112|T201|COMP|14939-3|LNC|Urea nitrogen|Urea nitrogen
C0798113|T201|COMP|14940-1|LNC|Uroporphyrin 1 isomer|Uroporphyrin 1 isomer
C0798114|T201|COMP|14941-9|LNC|Uroporphyrin 1 isomer|Uroporphyrin 1 isomer
C0798115|T201|COMP|14942-7|LNC|Uroporphyrin 1 isomer|Uroporphyrin 1 isomer
C0798116|T201|COMP|14943-5|LNC|Uroporphyrin 3 isomer|Uroporphyrin 3 isomer
C0798117|T201|COMP|14944-3|LNC|Uroporphyrin 3 isomer|Uroporphyrin 3 isomer
C0798118|T201|COMP|14945-0|LNC|Uroporphyrin 3 isomer|Uroporphyrin 3 isomer
C0798119|T201|COMP|14946-8|LNC|Valproate|Valproate
C0798120|T201|COMP|14947-6|LNC|Vanillylmandelate|Vanillylmandelate
C0798121|T201|COMP|14948-4|LNC|Vanillylmandelate/Creatinine|Vanillylmandelate/Creatinine
C0798122|T201|COMP|14949-2|LNC|Vasopressin|Vasopressin
C0798123|T201|COMP|14950-0|LNC|Viscosity|Viscosity
C0798124|T201|COMP|14951-8|LNC|Volatile drugs positive|Volatile drugs positive
C0798125|T201|COMP|14952-6|LNC|Xylose^1H post 25 g xylose PO|Xylose^1H post 25 g xylose PO
C0798126|T201|COMP|14953-4|LNC|Xylose^2H post 25 g xylose PO|Xylose^2H post 25 g xylose PO
C0798127|T201|COMP|14954-2|LNC|Xylose^post dose PO|Xylose^post dose PO
C0798128|T201|COMP|14955-9|LNC|Zinc|Zinc
C0798129|T201|COMP|14956-7|LNC|Albumin|Albumin
C0798130|T201|COMP|14957-5|LNC|Albumin|Albumin
C0798131|T201|COMP|14958-3|LNC|Albumin/Creatinine|Albumin/Creatinine
C0798132|T201|COMP|14959-1|LNC|Albumin/Creatinine|Albumin/Creatinine
C0798133|T201|COMP|14960-9|LNC|Estradiol.free/Estradiol.total|Estradiol.free/Estradiol.total
C0798143|T201|COMP|14970-8|LNC|Estrone.bioavailable|Estrone.bioavailable
C0798144|T201|COMP|14971-6|LNC|Estrone.bioavailable/Estrone.total|Estrone.bioavailable/Estrone.total
C0798145|T201|COMP|14972-4|LNC|Mycobacterium sp DNA|Mycobacterium sp DNA
C0798146|T201|COMP|14973-2|LNC|Mycobacterium sp DNA|Mycobacterium sp DNA
C0798147|T201|COMP|14974-0|LNC|Mycobacterium sp DNA|Mycobacterium sp DNA
C0798148|T201|COMP|14975-7|LNC|Human antimouse Ab|Human antimouse Ab
C0798149|T201|COMP|14976-5|LNC|Lecithin/Sphingomyelin|Lecithin/Sphingomyelin
C0798150|T201|COMP|14977-3|LNC|Immunoglobulin light chains.free|Immunoglobulin light chains.free
C0798151|T201|COMP|14978-1|LNC|cycloSPORINE|cycloSPORINE
C0798152|T201|COMP|14979-9|LNC|Coagulation surface induced|Coagulation surface induced
C0798153|T201|COMP|14980-7|LNC|A variant subtype Ab|A variant subtype Ab
C0798154|T201|COMP|14981-5|LNC|A variant subtype Ab|A variant subtype Ab
C0798155|T201|COMP|14982-3|LNC|A variant subtype Ab|A variant subtype Ab
C0798156|T201|COMP|14983-1|LNC|I (int) subtype|I (int) subtype
C0798157|T201|COMP|14984-9|LNC|I (int) subtype|I (int) subtype
C0798158|T201|COMP|14985-6|LNC|I (int) subtype|I (int) subtype
C0798159|T201|COMP|14986-4|LNC|little i-1 subtype|little i-1 subtype
C0798160|T201|COMP|14987-2|LNC|little i-1 subtype|little i-1 subtype
C0798161|T201|COMP|14988-0|LNC|little i-1 subtype|little i-1 subtype
C0798162|T201|COMP|14989-8|LNC|little i-2 subtype|little i-2 subtype
C0798163|T201|COMP|14990-6|LNC|little i-2 subtype|little i-2 subtype
C0798164|T201|COMP|14991-4|LNC|little i-2 subtype|little i-2 subtype
C0798165|T201|COMP|14992-2|LNC|O group|O group
C0798166|T201|COMP|14993-0|LNC|O group|O group
C0798167|T201|COMP|14994-8|LNC|O group|O group
C0798168|T201|COMP|14995-5|LNC|Glucose^2H post 75 g glucose PO|Glucose^2H post 75 g glucose PO
C0798169|T201|COMP|14996-3|LNC|Glucose^pre 75 g glucose PO|Glucose^pre 75 g glucose PO
C0798170|T201|COMP|14997-1|LNC|Thyrotropin^30M post dose TRH IV|Thyrotropin^30M post dose TRH IV
C0798171|T201|COMP|14998-9|LNC|Thyrotropin^1H post dose TRH IV|Thyrotropin^1H post dose TRH IV
C0798172|T201|COMP|14999-7|LNC|Thyrotropin^baseline|Thyrotropin^baseline
C0798173|T201|COMP|15000-3|LNC|Thyrotropin^pre dose TRH IV|Thyrotropin^pre dose TRH IV
C0798174|T201|COMP|15001-1|LNC|Xylose^1H post 25 g xylose PO|Xylose^1H post 25 g xylose PO
C0798175|T201|COMP|15002-9|LNC|Xylose^2H post 25 g xylose PO|Xylose^2H post 25 g xylose PO
C0798176|T201|COMP|15003-7|LNC|11-Hydroxyandrosterone|11-Hydroxyandrosterone
C0798177|T201|COMP|15004-5|LNC|11-Hydroxyetiocholanolone|11-Hydroxyetiocholanolone
C0798178|T201|COMP|15005-2|LNC|11-Ketoandrosterone|11-Ketoandrosterone
C0798179|T201|COMP|15006-0|LNC|11-Ketoetiocholanolone|11-Ketoetiocholanolone
C0798180|T201|COMP|15007-8|LNC|2,3-Diphosphoglycerate|2,3-Diphosphoglycerate
C0798181|T201|COMP|15008-6|LNC|3-Alpha-Androstanediol glucuronide|3-Alpha-Androstanediol glucuronide
C0798182|T201|COMP|15009-4|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C0798183|T201|COMP|15010-2|LNC|Aldosterone|Aldosterone
C0798184|T201|COMP|15011-0|LNC|Aldosterone^supine|Aldosterone^supine
C0798185|T201|COMP|15012-8|LNC|Aldosterone^upright|Aldosterone^upright
C0798192|T201|COMP|15019-3|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0798193|T201|COMP|15020-1|LNC|Amylase.P1/Amylase.total|Amylase.P1/Amylase.total
C0798194|T201|COMP|15021-9|LNC|Amylase.P2/Amylase.total|Amylase.P2/Amylase.total
C0798195|T201|COMP|15022-7|LNC|Amylase.P3/Amylase.total|Amylase.P3/Amylase.total
C0798196|T201|COMP|15023-5|LNC|Amylase.S1/Amylase.total|Amylase.S1/Amylase.total
C0798197|T201|COMP|15024-3|LNC|Amylase.S2/Amylase.total|Amylase.S2/Amylase.total
C0798198|T201|COMP|15025-0|LNC|Amylase.S3/Amylase.total|Amylase.S3/Amylase.total
C0798199|T201|COMP|15026-8|LNC|Androstanediol|Androstanediol
C0798200|T201|COMP|15027-6|LNC|Androstenedione|Androstenedione
C0798201|T201|COMP|15028-4|LNC|Androstenedione|Androstenedione
C0798202|T201|COMP|15029-2|LNC|Androsterone|Androsterone
C0798203|T201|COMP|15030-0|LNC|Androsterone|Androsterone
C0798204|T201|COMP|15031-8|LNC|Angiotensin I|Angiotensin I
C0798205|T201|COMP|15032-6|LNC|Angiotensin II|Angiotensin II
C0798206|T201|COMP|15033-4|LNC|Ascorbate|Ascorbate
C0798207|T201|COMP|15034-2|LNC|Bromide|Bromide
C0798208|T201|COMP|15035-9|LNC|Calcitonin|Calcitonin
C0798209|T201|COMP|15036-7|LNC|Catecholamines|Catecholamines
C0798210|T201|COMP|15037-5|LNC|Chymotrypsin|Chymotrypsin
C0798211|T201|COMP|15038-3|LNC|Citrate|Citrate
C0798212|T201|COMP|15039-1|LNC|Cobalamin|Cobalamin
C0798213|T201|COMP|15040-9|LNC|Coproporphyrin|Coproporphyrin
C0798214|T201|COMP|15041-7|LNC|Coproporphyrin|Coproporphyrin
C0798215|T201|COMP|15042-5|LNC|Corticotropin|Corticotropin
C0798216|T201|COMP|15043-3|LNC|Cortisol|Cortisol
C0798217|T201|COMP|15044-1|LNC|Cortisol.free|Cortisol.free
C0798218|T201|COMP|15045-8|LNC|Creatine|Creatine
C0798219|T201|COMP|15046-6|LNC|Creatine|Creatine
C0798220|T201|COMP|15047-4|LNC|Creatine|Creatine
C0798221|T201|COMP|15048-2|LNC|Creatine kinase.BB/Creatine kinase.total|Creatine kinase.BB/Creatine kinase.total
C0798222|T201|COMP|15049-0|LNC|Creatine kinase.MM/Creatine kinase.total|Creatine kinase.MM/Creatine kinase.total
C0798223|T201|COMP|15050-8|LNC|Creatinine|Creatinine
C0798224|T201|COMP|15051-6|LNC|Creatinine|Creatinine
C0798225|T201|COMP|15052-4|LNC|Cobalamins.unsaturated binding capacity|Cobalamins.unsaturated binding capacity
C0798226|T201|COMP|15053-2|LNC|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C0798227|T201|COMP|15054-0|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C0798228|T201|COMP|15055-7|LNC|Deoxypyridinoline|Deoxypyridinoline
C0798229|T201|COMP|15057-3|LNC|Androstanolone|Androstanolone
C0798230|T201|COMP|15058-1|LNC|DOPamine|DOPamine
C0798231|T201|COMP|15059-9|LNC|DOPamine|DOPamine
C0798232|T201|COMP|15060-7|LNC|Enolase.neuron specific|Enolase.neuron specific
C0798233|T201|COMP|15061-5|LNC|Erythropoietin|Erythropoietin
C0798234|T201|COMP|15062-3|LNC|Estradiol.unconjugated|Estradiol.unconjugated
C0798235|T201|COMP|15063-1|LNC|Estriol.conjugated|Estriol.conjugated
C0798236|T201|COMP|15064-9|LNC|Estriol.unconjugated|Estriol.unconjugated
C0798237|T201|COMP|15065-6|LNC|Etiocholanolone|Etiocholanolone
C0798239|T201|COMP|15067-2|LNC|Follitropin|Follitropin
C0798240|T201|COMP|15068-0|LNC|Follitropin|Follitropin
C0798241|T201|COMP|15069-8|LNC|Fructosamine|Fructosamine
C0798242|T201|COMP|15070-6|LNC|Fructose|Fructose
C0798243|T201|COMP|15071-4|LNC|Galactose|Galactose
C0798244|T201|COMP|15072-2|LNC|Gastrin|Gastrin
C0798245|T201|COMP|15073-0|LNC|Glucagon|Glucagon
C0798246|T201|COMP|15074-8|LNC|Glucose|Glucose
C0798247|T201|COMP|15075-5|LNC|Glucose|Glucose
C0798248|T201|COMP|15076-3|LNC|Glucose|Glucose
C0798249|T201|COMP|15077-1|LNC|Glucose|Glucose
C0798250|T201|COMP|15078-9|LNC|Lactate|Lactate
C0798251|T201|COMP|15079-7|LNC|Lutropin|Lutropin
C0798252|T201|COMP|15080-5|LNC|Lutropin|Lutropin
C0798253|T201|COMP|15081-3|LNC|Prolactin|Prolactin
C0798254|T201|COMP|15082-1|LNC|Methemoglobin|Methemoglobin
C0798255|T201|COMP|15083-9|LNC|Normetanephrine|Normetanephrine
C0798256|T201|COMP|15084-7|LNC|Osteocalcin|Osteocalcin
C0798257|T201|COMP|15085-4|LNC|Oxalate|Oxalate
C0798258|T201|COMP|15086-2|LNC|Oxalate|Oxalate
C0798259|T201|COMP|15087-0|LNC|Parathyrin related protein|Parathyrin related protein
C0798260|T201|COMP|15088-8|LNC|Parathyrin.C-terminal|Parathyrin.C-terminal
C0798261|T201|COMP|15089-6|LNC|Phospholipid|Phospholipid
C0798262|T201|COMP|15090-4|LNC|Porphyrins|Porphyrins
C0798263|T201|COMP|15091-2|LNC|Pregnanediol|Pregnanediol
C0798264|T201|COMP|15092-0|LNC|Pregnanetriol|Pregnanetriol
C0798265|T201|COMP|15093-8|LNC|Protoporphyrin.free|Protoporphyrin.free
C0798266|T201|COMP|15094-6|LNC|Testosterone|Testosterone
C0798267|T201|COMP|15095-3|LNC|Testosterone|Testosterone
C0798268|T201|COMP|15096-1|LNC|Uroporphyrin|Uroporphyrin
C0798269|T201|COMP|15097-9|LNC|Vanillylmandelate|Vanillylmandelate
C0798270|T201|COMP|15098-7|LNC|Amikacin^random|Amikacin^random
C0798271|T201|COMP|15099-5|LNC|Amiodarone|Amiodarone
C0798272|T201|COMP|15100-1|LNC|Barbiturates|Barbiturates
C0798273|T201|COMP|15101-9|LNC|Chloramphenicol|Chloramphenicol
C0798274|T201|COMP|15102-7|LNC|Codeine|Codeine
C0798275|T201|COMP|15103-5|LNC|cycloSPORINE|cycloSPORINE
C0798276|T201|COMP|15104-3|LNC|Digitoxin|Digitoxin
C0798277|T201|COMP|15105-0|LNC|Flecainide|Flecainide
C0798278|T201|COMP|15106-8|LNC|Gentamicin^random|Gentamicin^random
C0798279|T201|COMP|15107-6|LNC|Imipramine|Imipramine
C0798280|T201|COMP|15108-4|LNC|Methadone|Methadone
C0798281|T201|COMP|15109-2|LNC|Midazolam|Midazolam
C0798282|T201|COMP|15110-0|LNC|Morphine|Morphine
C0798283|T201|COMP|15111-8|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0798284|T201|COMP|15112-6|LNC|Phosphatase.leukocyte|Phosphatase.leukocyte
C0798285|T201|COMP|15113-4|LNC|Aluminum|Aluminum
C0798286|T201|COMP|15114-2|LNC|Arsenic|Arsenic
C0798287|T201|COMP|15115-9|LNC|Arsenic|Arsenic
C0798288|T201|COMP|15117-5|LNC|Cadmium|Cadmium
C0798289|T201|COMP|15118-3|LNC|Chromium|Chromium
C0798290|T201|COMP|15119-1|LNC|Cobalt|Cobalt
C0798291|T201|COMP|15120-9|LNC|Ethanol|Ethanol
C0798292|T201|COMP|15121-7|LNC|Lipoprotein.alpha/Lipoprotein.total|Lipoprotein.alpha/Lipoprotein.total
C0798293|T201|COMP|15122-5|LNC|Lipoprotein.beta/Lipoprotein.total|Lipoprotein.beta/Lipoprotein.total
C0798294|T201|COMP|15123-3|LNC|Lipoprotein.pre-beta/Lipoprotein.total|Lipoprotein.pre-beta/Lipoprotein.total
C0798295|T201|COMP|15124-1|LNC|Albumin/Protein.total|Albumin/Protein.total
C0798296|T201|COMP|15125-8|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0798297|T201|COMP|15126-6|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0798298|T201|COMP|15127-4|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C0798299|T201|COMP|15128-2|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0798300|T201|COMP|15129-0|LNC|Fibrin D-dimer|Fibrin D-dimer
C0798301|T201|COMP|15130-8|LNC|Methionine+Tryptophan|Methionine+Tryptophan
C0798302|T201|COMP|15131-6|LNC|Isoleucine+Leucine|Isoleucine+Leucine
C0798303|T201|COMP|15132-4|LNC|Beta aminoisobutyrate+Proline|Beta aminoisobutyrate+Proline
C0798304|T201|COMP|15133-2|LNC|Anserine+Carnosine+Cysteine+Histidine+Ornithine|Anserine+Carnosine+Cysteine+Histidine+Ornithine
C0798305|T201|COMP|15134-0|LNC|Glutamate+Glutamine+Threonine|Glutamate+Glutamine+Threonine
C0798307|T201|COMP|15136-5|LNC|Arginine+Argininosuccinate+Lysine+Serine+Taurine|Arginine+Argininosuccinate+Lysine+Serine+Taurine
C0798308|T201|COMP|15137-3|LNC|Alanine+Ethanolamine|Alanine+Ethanolamine
C0798309|T201|COMP|15138-1|LNC|Isoleucine+Leucine|Isoleucine+Leucine
C0798310|T201|COMP|15139-9|LNC|Anserine+Carnosine+Cysteine+Histidine+Ornithine|Anserine+Carnosine+Cysteine+Histidine+Ornithine
C0798311|T201|COMP|15140-7|LNC|Arginine+Argininosuccinate+Lysine+Serine+Taurine|Arginine+Argininosuccinate+Lysine+Serine+Taurine
C0798312|T201|COMP|15141-5|LNC|Beta aminoisobutyrate+Proline|Beta aminoisobutyrate+Proline
C0798313|T201|COMP|15142-3|LNC|Alanine+Ethanolamine|Alanine+Ethanolamine
C0798315|T201|COMP|15144-9|LNC|Glutamate+Glutamine+Threonine|Glutamate+Glutamine+Threonine
C0798316|T201|COMP|15145-6|LNC|Methionine+Tryptophan|Methionine+Tryptophan
C0798317|T201|COMP|15146-4|LNC|Acetone|Acetone
C0798318|T201|COMP|15147-2|LNC|Acetone|Acetone
C0798319|T201|COMP|15148-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798320|T201|COMP|15149-8|LNC|Ammonia|Ammonia
C0798321|T201|COMP|15150-6|LNC|Anisocytosis|Anisocytosis
C0798322|T201|COMP|15151-4|LNC|Aspergillus fumigatus 3 Ab|Aspergillus fumigatus 3 Ab
C0798323|T201|COMP|15152-2|LNC|Bilirubin.glucuronidated|Bilirubin.glucuronidated
C0798324|T201|COMP|15153-0|LNC|Bilirubin.non-glucuronidated|Bilirubin.non-glucuronidated
C0798325|T201|COMP|15154-8|LNC|Blasts|Blasts
C0798326|T201|COMP|15155-5|LNC|Calcium|Calcium
C0798327|T201|COMP|15156-3|LNC|Cancer Ag 125|Cancer Ag 125
C0798328|T201|COMP|15157-1|LNC|Cancer Ag 125|Cancer Ag 125
C0798329|T201|COMP|15158-9|LNC|Chloride|Chloride
C0798330|T201|COMP|15159-7|LNC|Coagulation factor.extrinsic pathway|Coagulation factor.extrinsic pathway
C0798331|T201|COMP|15160-5|LNC|Coagulation factor.intrinsic factor|Coagulation factor.intrinsic factor
C0798332|T201|COMP|15161-3|LNC|Complement C1 esterase inhibitor.functional|Complement C1 esterase inhibitor.functional
C0798333|T201|COMP|15162-1|LNC|Complement C1q|Complement C1q
C0798334|T201|COMP|15163-9|LNC|Complement C2|Complement C2
C0798335|T201|COMP|15164-7|LNC|Complement C3|Complement C3
C0798336|T201|COMP|15165-4|LNC|Complement C4|Complement C4
C0798337|T201|COMP|15166-2|LNC|Complement C5|Complement C5
C0798338|T201|COMP|15167-0|LNC|Complement C6|Complement C6
C0798339|T201|COMP|15168-8|LNC|Complement total hemolytic C50|Complement total hemolytic C50
C0798340|T201|COMP|15169-6|LNC|Complement total hemolytic C50|Complement total hemolytic C50
C0798341|T201|COMP|15170-4|LNC|Complement total hemolytic C50|Complement total hemolytic C50
C0798342|T201|COMP|15171-2|LNC|Cryoglobulin.IgA|Cryoglobulin.IgA
C0798343|T201|COMP|15172-0|LNC|Cryoglobulin.IgG|Cryoglobulin.IgG
C0798344|T201|COMP|15173-8|LNC|Cryoglobulin.IgM|Cryoglobulin.IgM
C0798345|T201|COMP|15174-6|LNC|Cryoglobulin/Serum.total|Cryoglobulin/Serum.total
C0798346|T201|COMP|15175-3|LNC|Cryoproteins|Cryoproteins
C0798347|T201|COMP|15176-1|LNC|Cryoproteins identified|Cryoproteins identified
C0798348|T201|COMP|15177-9|LNC|DNA double strand Ab|DNA double strand Ab
C0798349|T201|COMP|15178-7|LNC|Complement factor B|Complement factor B
C0798350|T201|COMP|15179-5|LNC|Fibrin D-dimer|Fibrin D-dimer
C0798351|T201|COMP|15180-3|LNC|Hypochromia|Hypochromia
C0798352|T201|COMP|15181-1|LNC|IgA|IgA
C0798353|T201|COMP|15182-9|LNC|IgA|IgA
C0798354|T201|COMP|15183-7|LNC|IgG|IgG
C0798355|T201|COMP|15184-5|LNC|IgG|IgG
C0798356|T201|COMP|15185-2|LNC|IgM|IgM
C0798357|T201|COMP|15186-0|LNC|IgM|IgM
C0798358|T201|COMP|15187-8|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C0798359|T201|COMP|15188-6|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C0798361|T201|COMP|15190-2|LNC|Leukocytes other|Leukocytes other
C0798363|T201|COMP|15192-8|LNC|Lymphocytes.variant|Lymphocytes.variant
C0798364|T201|COMP|15193-6|LNC|Cells.CD3-CD16+|Cells.CD3-CD16+
C0798365|T201|COMP|15194-4|LNC|Cells.CD3-CD16+/100 cells|Cells.CD3-CD16+/100 cells
C0798366|T201|COMP|15195-1|LNC|Cells.CD3-CD19+|Cells.CD3-CD19+
C0798367|T201|COMP|15196-9|LNC|Cells.CD3-CD19+/100 cells|Cells.CD3-CD19+/100 cells
C0798368|T201|COMP|15197-7|LNC|Lymphocytes.clefted/100 leukocytes|Lymphocytes.clefted/100 leukocytes
C0798369|T201|COMP|15198-5|LNC|Macrocytes|Macrocytes
C0798370|T201|COMP|15199-3|LNC|Microcytes|Microcytes
C0798371|T201|COMP|15200-9|LNC|Osmolality|Osmolality
C0798372|T201|COMP|15201-7|LNC|Platelets.large fragments|Platelets.large fragments
C0798373|T201|COMP|15202-5|LNC|Potassium|Potassium
C0798374|T201|COMP|15203-3|LNC|Rheumatoid factor|Rheumatoid factor
C0798375|T201|COMP|15204-1|LNC|Rheumatoid factor|Rheumatoid factor
C0798376|T201|COMP|15205-8|LNC|Rheumatoid factor|Rheumatoid factor
C0798377|T201|COMP|15206-6|LNC|Rheumatoid factor|Rheumatoid factor
C0798378|T201|COMP|15207-4|LNC|Sodium|Sodium
C0798379|T201|COMP|15208-2|LNC|Taurine|Taurine
C0798380|T201|COMP|15209-0|LNC|Saccharomonospora viridis Ab|Saccharomonospora viridis Ab
C0798381|T201|COMP|15210-8|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C0798382|T201|COMP|15211-6|LNC|Biopsy|Biopsy
C0798383|T201|COMP|15212-4|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C0798434|T201|COMP|15263-7|LNC|(Cottonwood+Elm+Maple+Oak+Pecan tree) Ab.IgE|(Cottonwood+Elm+Maple+Oak+Pecan tree) Ab.IgE
C0798448|T201|COMP|15278-5|LNC|Levisticum officinale Ab.IgE|Levisticum officinale Ab.IgE
C0798449|T201|COMP|15279-3|LNC|Elettaria cardamomum Ab.IgE|Elettaria cardamomum Ab.IgE
C0798450|T201|COMP|15280-1|LNC|Mace Ab.IgE|Mace Ab.IgE
C0798451|T201|COMP|15281-9|LNC|Gasterophilus intestinalis Ab.IgE|Gasterophilus intestinalis Ab.IgE
C0798452|T201|COMP|6236-4|LNC|Secale cereale pollen Ab.IgE|Secale cereale pollen Ab.IgE
C0798453|T201|COMP|15283-5|LNC|Betula verrucosa Ab.IgE|Betula verrucosa Ab.IgE
C0798454|T201|COMP|15284-3|LNC|Alnus incana Ab.IgE|Alnus incana Ab.IgE
C0798455|T201|COMP|15285-0|LNC|Platanus acerifolia Ab.IgE|Platanus acerifolia Ab.IgE
C0798505|T201|COMP|15336-1|LNC|Antibiotic XXX|Antibiotic XXX
C0798506|T201|COMP|15337-9|LNC|Antibiotic XXX^peak|Antibiotic XXX^peak
C0798507|T201|COMP|15338-7|LNC|Antibiotic XXX^trough|Antibiotic XXX^trough
C0798508|T201|COMP|15339-5|LNC|Trogoderma angustum Ab.IgE|Trogoderma angustum Ab.IgE
C0798509|T201|COMP|15340-3|LNC|Cedar italian Ab.IgE|Cedar italian Ab.IgE
C0798510|T201|COMP|15341-1|LNC|Simulium venustum Ab.IgE|Simulium venustum Ab.IgE
C0798511|T201|COMP|15342-9|LNC|Vespa crabro Ab.IgE|Vespa crabro Ab.IgE
C0798512|T201|COMP|15343-7|LNC|Blood group antibody screen|Blood group antibody screen
C0798513|T201|COMP|15344-5|LNC|little i Ab|little i Ab
C0798514|T201|COMP|15345-2|LNC|Aldosterone^1H post XXX challenge|Aldosterone^1H post XXX challenge
C0798515|T201|COMP|15346-0|LNC|Aldosterone^30M post XXX challenge|Aldosterone^30M post XXX challenge
C0798516|T201|COMP|15347-8|LNC|Somatotropin^30M post XXX challenge|Somatotropin^30M post XXX challenge
C0798519|T201|COMP|15350-2|LNC|Amylase|Amylase
C0798520|T201|COMP|15351-0|LNC|Apolipoprotein E2|Apolipoprotein E2
C0798521|T201|COMP|15352-8|LNC|Apolipoprotein E3|Apolipoprotein E3
C0798522|T201|COMP|15353-6|LNC|Apolipoprotein E4|Apolipoprotein E4
C0798523|T201|COMP|15354-4|LNC|Bombesin Ag|Bombesin Ag
C0798524|T201|COMP|15355-1|LNC|Estrone sulfate|Estrone sulfate
C0798525|T201|COMP|15356-9|LNC|Globulin|Globulin
C0798526|T201|COMP|15357-7|LNC|Iron|Iron
C0798527|T201|COMP|15358-5|LNC|Macroamylase|Macroamylase
C0798531|T201|COMP|15362-7|LNC|Coagulation surface induced.inhibitor sensitive|Coagulation surface induced.inhibitor sensitive
C0798532|T201|COMP|15363-5|LNC|Busulfan|Busulfan
C0798533|T201|COMP|15364-3|LNC|Codeine|Codeine
C0798534|T201|COMP|15365-0|LNC|Codeine|Codeine
C0798535|T201|COMP|15366-8|LNC|Dextroamphetamine|Dextroamphetamine
C0798536|T201|COMP|15367-6|LNC|Ganciclovir|Ganciclovir
C0798537|T201|COMP|15368-4|LNC|Hypoglycemics.sulfonyluric|Hypoglycemics.sulfonyluric
C0798538|T201|COMP|15369-2|LNC|Lithium.saliva/Lithium.serum|Lithium.saliva/Lithium.serum
C0798539|T201|COMP|15370-0|LNC|Morphine|Morphine
C0798540|T201|COMP|15371-8|LNC|Morphine|Morphine
C0798541|T201|COMP|15372-6|LNC|Nordiazepam|Nordiazepam
C0798542|T201|COMP|15373-4|LNC|Phenyltoloxamine|Phenyltoloxamine
C0798543|T201|COMP|15374-2|LNC|Sulfonylurea|Sulfonylurea
C0798544|T201|COMP|15375-9|LNC|Valproate.free|Valproate.free
C0798545|T201|COMP|15376-7|LNC|Spermatozoa.abnormal/100 spermatozoa|Spermatozoa.abnormal/100 spermatozoa
C0798546|T201|COMP|15377-5|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0798547|T201|COMP|15378-3|LNC|Fungus identified|Fungus identified
C0798548|T201|COMP|15379-1|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C0798549|T201|COMP|15380-9|LNC|Leishmania braziliensis Ab.IgG|Leishmania braziliensis Ab.IgG
C0798550|T201|COMP|15381-7|LNC|Leishmania braziliensis Ab.IgM|Leishmania braziliensis Ab.IgM
C0798551|T201|COMP|15382-5|LNC|Leishmania donovani Ab.IgG|Leishmania donovani Ab.IgG
C0798552|T201|COMP|15383-3|LNC|Leishmania donovani Ab.IgM|Leishmania donovani Ab.IgM
C0798553|T201|COMP|15384-1|LNC|Leishmania mexicana Ab.IgG|Leishmania mexicana Ab.IgG
C0798554|T201|COMP|15385-8|LNC|Leishmania mexicana Ab.IgM|Leishmania mexicana Ab.IgM
C0798555|T201|COMP|15386-6|LNC|Leishmania tropica Ab.IgG|Leishmania tropica Ab.IgG
C0798556|T201|COMP|15387-4|LNC|Leishmania tropica Ab.IgM|Leishmania tropica Ab.IgM
C0798557|T201|COMP|15388-2|LNC|Mycoplasma hominis|Mycoplasma hominis
C0798558|T201|COMP|15389-0|LNC|Parainfluenza virus 1 Ab.IgG|Parainfluenza virus 1 Ab.IgG
C0798559|T201|COMP|15390-8|LNC|Parainfluenza virus 1 Ab.IgM|Parainfluenza virus 1 Ab.IgM
C0798560|T201|COMP|15391-6|LNC|Parainfluenza virus 1 Ab.IgM|Parainfluenza virus 1 Ab.IgM
C0798561|T201|COMP|15392-4|LNC|Parainfluenza virus 2 Ab.IgG|Parainfluenza virus 2 Ab.IgG
C0798562|T201|COMP|15393-2|LNC|Parainfluenza virus 2 Ab.IgM|Parainfluenza virus 2 Ab.IgM
C0798563|T201|COMP|15394-0|LNC|Parainfluenza virus 3 Ab.IgG|Parainfluenza virus 3 Ab.IgG
C0798564|T201|COMP|15395-7|LNC|Parainfluenza virus 3 Ab.IgM|Parainfluenza virus 3 Ab.IgM
C0798565|T201|COMP|15396-5|LNC|Toxoplasma sp Ab.IgG|Toxoplasma sp Ab.IgG
C0798566|T201|COMP|15397-3|LNC|Trypanosoma cruzi Ab.IgM|Trypanosoma cruzi Ab.IgM
C0798567|T201|COMP|15398-1|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C0798568|T201|COMP|15399-9|LNC|Neuronal nuclear Ab.IgG|Neuronal nuclear Ab.IgG
C0798569|T201|COMP|15400-5|LNC|Platelet Ab.IgG|Platelet Ab.IgG
C0798570|T201|COMP|15401-3|LNC|Drugs identified|Drugs identified
C0798571|T201|COMP|15402-1|LNC|Ethanol|Ethanol
C0798572|T201|COMP|15403-9|LNC|Isopropanol|Isopropanol
C0798573|T201|COMP|15404-7|LNC|Levomethamphetamine/Amphetamines.total|Levomethamphetamine/Amphetamines.total
C0798574|T201|COMP|15405-4|LNC|Methamphetamine|Methamphetamine
C0798575|T201|COMP|15406-2|LNC|Methamphetamine|Methamphetamine
C0798576|T201|COMP|15407-0|LNC|Methanol|Methanol
C0798577|T201|COMP|15408-8|LNC|Thallium|Thallium
C0798578|T201|COMP|15409-6|LNC|Thallium|Thallium
C0798579|T201|COMP|15410-4|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0798580|T201|COMP|15411-2|LNC|Ergosterol|Ergosterol
C0798581|T201|COMP|15412-0|LNC|Service comment 21|Service comment 21
C0798582|T201|COMP|15413-8|LNC|Service comment 22|Service comment 22
C0798583|T201|COMP|15414-6|LNC|Service comment 23|Service comment 23
C0798584|T201|COMP|15415-3|LNC|Service comment 24|Service comment 24
C0798585|T201|COMP|15416-1|LNC|Service comment 25|Service comment 25
C0798586|T201|COMP|15417-9|LNC|Service comment 26|Service comment 26
C0798587|T201|COMP|15418-7|LNC|Service comment 27|Service comment 27
C0798588|T201|COMP|15419-5|LNC|Service comment 28|Service comment 28
C0798589|T201|COMP|15420-3|LNC|Service comment 29|Service comment 29
C0798590|T201|COMP|15421-1|LNC|Service comment 30|Service comment 30
C0798591|T201|COMP|15422-9|LNC|Service comment 31|Service comment 31
C0798592|T201|COMP|15423-7|LNC|Service comment 32|Service comment 32
C0798593|T201|COMP|15424-5|LNC|Service comment 33|Service comment 33
C0798594|T201|COMP|15425-2|LNC|Service comment 34|Service comment 34
C0798595|T201|COMP|15426-0|LNC|Service comment 35|Service comment 35
C0798596|T201|COMP|15427-8|LNC|Service comment 36|Service comment 36
C0798597|T201|COMP|15428-6|LNC|Service comment 37|Service comment 37
C0798598|T201|COMP|15429-4|LNC|Service comment 38|Service comment 38
C0798599|T201|COMP|15430-2|LNC|Service comment 39|Service comment 39
C0798600|T201|COMP|15431-0|LNC|Service comment 40|Service comment 40
C0798601|T201|COMP|15432-8|LNC|Testosterone.free/Testosterone.total|Testosterone.free/Testosterone.total
C0798602|T201|COMP|15433-6|LNC|Anaplasma marginale Ab|Anaplasma marginale Ab
C0798603|T201|COMP|15434-4|LNC|Avian adenovirus Ab|Avian adenovirus Ab
C0798604|T201|COMP|15435-1|LNC|Avian adenovirus 2 Ab|Avian adenovirus 2 Ab
C0798605|T201|COMP|15436-9|LNC|Avian encephalomyelitis virus Ab|Avian encephalomyelitis virus Ab
C0798606|T201|COMP|15437-7|LNC|Avian encephalomyelitis virus Ab|Avian encephalomyelitis virus Ab
C0798607|T201|COMP|15438-5|LNC|Avian hemorrhagic enteritis virus Ab|Avian hemorrhagic enteritis virus Ab
C0798608|T201|COMP|15439-3|LNC|Infectious bronchitis virus Ark-99 Ab|Infectious bronchitis virus Ark-99 Ab
C0798609|T201|COMP|15440-1|LNC|Infectious bronchitis virus Mass-41 Ab|Infectious bronchitis virus Mass-41 Ab
C0798610|T201|COMP|15441-9|LNC|Infectious bronchitis virus Conn-42 Ab|Infectious bronchitis virus Conn-42 Ab
C0798611|T201|COMP|15442-7|LNC|Avian infectious laryngotracheitis virus Ab|Avian infectious laryngotracheitis virus Ab
C0798612|T201|COMP|15443-5|LNC|Avian infectious laryngotracheitis virus Ab|Avian infectious laryngotracheitis virus Ab
C0798613|T201|COMP|15444-3|LNC|Influenza virus A Ab|Influenza virus A Ab
C0798614|T201|COMP|15445-0|LNC|Avian leukosis virus Ag|Avian leukosis virus Ag
C0798615|T201|COMP|15446-8|LNC|Avian leukosis virus Ag|Avian leukosis virus Ag
C0798616|T201|COMP|15447-6|LNC|Avian paramyxovirus 1 Ab|Avian paramyxovirus 1 Ab
C0798617|T201|COMP|15448-4|LNC|Avian paramyxovirus 1 Ab|Avian paramyxovirus 1 Ab
C0798618|T201|COMP|15449-2|LNC|Avian paramyxovirus 2 Ab|Avian paramyxovirus 2 Ab
C0798619|T201|COMP|15450-0|LNC|Avian paramyxovirus 3 Ab|Avian paramyxovirus 3 Ab
C0798620|T201|COMP|15451-8|LNC|Avian pox virus Ab|Avian pox virus Ab
C0798621|T201|COMP|15452-6|LNC|Avian reovirus Ab|Avian reovirus Ab
C0798622|T201|COMP|15453-4|LNC|Avian reovirus Ab|Avian reovirus Ab
C0798623|T201|COMP|15454-2|LNC|Reticuloendotheliosis virus Ab|Reticuloendotheliosis virus Ab
C0798624|T201|COMP|15455-9|LNC|Bluetongue virus Ab|Bluetongue virus Ab
C0798625|T201|COMP|15456-7|LNC|Bluetongue virus Ab|Bluetongue virus Ab
C0798626|T201|COMP|15457-5|LNC|Bordetella avium Ab|Bordetella avium Ab
C0798627|T201|COMP|15458-3|LNC|Bordetella avium Ab|Bordetella avium Ab
C0798628|T201|COMP|15459-1|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C0798629|T201|COMP|15460-9|LNC|Bovine leukemia virus Ab|Bovine leukemia virus Ab
C0798630|T201|COMP|15461-7|LNC|Bovine leukemia virus Ab|Bovine leukemia virus Ab
C0798631|T201|COMP|15462-5|LNC|Bovine diarrhea virus 1 Ab|Bovine diarrhea virus 1 Ab
C0798632|T201|COMP|15463-3|LNC|Bovine diarrhea virus 2 Ab|Bovine diarrhea virus 2 Ab
C0798635|T201|COMP|15466-6|LNC|Epizootic hemorrhagic disease virus Ab|Epizootic hemorrhagic disease virus Ab
C0798636|T201|COMP|15467-4|LNC|Equine herpesvirus 1 Ab|Equine herpesvirus 1 Ab
C0798637|T201|COMP|15468-2|LNC|Equine infectious anemia virus Ab|Equine infectious anemia virus Ab
C0798638|T201|COMP|15469-0|LNC|Equine influenza virus A1 Ab|Equine influenza virus A1 Ab
C0798639|T201|COMP|15470-8|LNC|Equine influenza virus A2 Ab|Equine influenza virus A2 Ab
C0798640|T201|COMP|15471-6|LNC|Equine influenza virus A2 Ab|Equine influenza virus A2 Ab
C0798641|T201|COMP|15472-4|LNC|Equine influenza virus Ag|Equine influenza virus Ag
C0798642|T201|COMP|15473-2|LNC|Equine arteritis virus Ab|Equine arteritis virus Ab
C0798643|T201|COMP|15474-0|LNC|Infectious bursal disease virus Ab|Infectious bursal disease virus Ab
C0798644|T201|COMP|15475-7|LNC|Infectious bursal disease virus Ab|Infectious bursal disease virus Ab
C0798645|T201|COMP|15476-5|LNC|Leptospira interrogans serovar Bratislava Ab|Leptospira interrogans serovar Bratislava Ab
C0798646|T201|COMP|15477-3|LNC|Leptospira interrogans serovar Canicola Ab|Leptospira interrogans serovar Canicola Ab
C0798647|T201|COMP|15478-1|LNC|Leptospira interrogans serovar Grippotyphosa Ab|Leptospira interrogans serovar Grippotyphosa Ab
C0798648|T201|COMP|15479-9|LNC|Leptospira interrogans serovar Hardjo Ab|Leptospira interrogans serovar Hardjo Ab
C0798650|T201|COMP|15481-5|LNC|Leptospira interrogans serovar Pomona Ab|Leptospira interrogans serovar Pomona Ab
C0798653|T201|COMP|15484-9|LNC|Mycoplasma gallisepticum Ab|Mycoplasma gallisepticum Ab
C0798654|T201|COMP|15485-6|LNC|Mycoplasma gallisepticum Ab|Mycoplasma gallisepticum Ab
C0798655|T201|COMP|15486-4|LNC|Mycoplasma gallisepticum rRNA|Mycoplasma gallisepticum rRNA
C0798656|T201|COMP|15487-2|LNC|Mycoplasma meleagridis Ab|Mycoplasma meleagridis Ab
C0798657|T201|COMP|15488-0|LNC|Mycoplasma meleagridis Ab|Mycoplasma meleagridis Ab
C0798658|T201|COMP|15489-8|LNC|Mycoplasma synoviae Ab|Mycoplasma synoviae Ab
C0798659|T201|COMP|15490-6|LNC|Mycoplasma synoviae Ab|Mycoplasma synoviae Ab
C0798660|T201|COMP|15491-4|LNC|Mycoplasma synoviae rRNA|Mycoplasma synoviae rRNA
C0798661|T201|COMP|15492-2|LNC|Neospora caninum Ab|Neospora caninum Ab
C0798662|T201|COMP|15493-0|LNC|Parainfluenza virus 3 Ab|Parainfluenza virus 3 Ab
C0798663|T201|COMP|15494-8|LNC|Pasteurella multocida Ab|Pasteurella multocida Ab
C0798666|T201|COMP|15497-1|LNC|Pseudorabies virus Ab|Pseudorabies virus Ab
C0798667|T201|COMP|15498-9|LNC|Pseudorabies virus Ab|Pseudorabies virus Ab
C0798668|T201|COMP|15499-7|LNC|Pseudorabies virus Ab|Pseudorabies virus Ab
C0798669|T201|COMP|15500-2|LNC|Pseudorabies virus.ClinEase gene deletion Ab|Pseudorabies virus.ClinEase gene deletion Ab
C0798670|T201|COMP|15501-0|LNC|Pseudorabies virus.HerdCheck gene deletion Ab|Pseudorabies virus.HerdCheck gene deletion Ab
C0798671|T201|COMP|15502-8|LNC|Pseudorabies virus.OmniMark gene deletion Ab|Pseudorabies virus.OmniMark gene deletion Ab
C0798672|T201|COMP|15503-6|LNC|Pseudorabies virus.Tolvid gene deletion Ab|Pseudorabies virus.Tolvid gene deletion Ab
C0798673|T201|COMP|15504-4|LNC|Salmonella arizonae Ab|Salmonella arizonae Ab
C0798674|T201|COMP|15505-1|LNC|Salmonella pullorum Ab|Salmonella pullorum Ab
C0798675|T201|COMP|15506-9|LNC|Salmonella typhimurium Ab|Salmonella typhimurium Ab
C0798685|T201|COMP|15518-4|LNC|Haliotis spp Ab.IgE.RAST class|Haliotis spp Ab.IgE.RAST class
C0798686|T201|COMP|15519-2|LNC|Acacia longifolia Ab.IgE.RAST class|Acacia longifolia Ab.IgE.RAST class
C0798687|T201|COMP|15520-0|LNC|Corticotropin Ab.IgE.RAST class|Corticotropin Ab.IgE.RAST class
C0798688|T201|COMP|15521-8|LNC|Alnus rhombifolia Ab.IgE.RAST class|Alnus rhombifolia Ab.IgE.RAST class
C0798689|T201|COMP|15522-6|LNC|Alder Ab.IgE.RAST class|Alder Ab.IgE.RAST class
C0798690|T201|COMP|15523-4|LNC|Alnus rugosa Ab.IgE.RAST class|Alnus rugosa Ab.IgE.RAST class
C0798691|T201|COMP|15524-2|LNC|Medicago sativa Ab.IgE.RAST class|Medicago sativa Ab.IgE.RAST class
C0798692|T201|COMP|15525-9|LNC|Alkalase Ab.IgE.RAST class|Alkalase Ab.IgE.RAST class
C0798693|T201|COMP|15526-7|LNC|Pimenta dioica Ab.IgE.RAST class|Pimenta dioica Ab.IgE.RAST class
C0798694|T201|COMP|15527-5|LNC|Prunus dulcis Ab.IgE.RAST class|Prunus dulcis Ab.IgE.RAST class
C0798695|T201|COMP|15528-3|LNC|Prunus dulcis tree Ab.IgE.RAST class|Prunus dulcis tree Ab.IgE.RAST class
C0798696|T201|COMP|15529-1|LNC|Lactalbumin alpha Ab.IgE.RAST class|Lactalbumin alpha Ab.IgE.RAST class
C0798698|T201|COMP|15530-9|LNC|Alternaria alternata Ab.IgE.RAST class|Alternaria alternata Ab.IgE.RAST class
C0798699|T201|COMP|15532-5|LNC|Amoxicillin Ab.IgE.RAST class|Amoxicillin Ab.IgE.RAST class
C0798700|T201|COMP|15533-3|LNC|Ampicillin Ab.IgE.RAST class|Ampicillin Ab.IgE.RAST class
C0798701|T201|COMP|15534-1|LNC|Engraulis encrasicolus Ab.IgE.RAST class|Engraulis encrasicolus Ab.IgE.RAST class
C0798702|T201|COMP|15535-8|LNC|Anisakis Ab.IgE.RAST class|Anisakis Ab.IgE.RAST class
C0798703|T201|COMP|15536-6|LNC|Pimpinella anisum Ab.IgE.RAST class|Pimpinella anisum Ab.IgE.RAST class
C0798705|T201|COMP|15537-4|LNC|Solenopsis invicta Ab.IgE.RAST class|Solenopsis invicta Ab.IgE.RAST class
C0798706|T201|COMP|15539-0|LNC|Malus sylvestris Ab.IgE.RAST class|Malus sylvestris Ab.IgE.RAST class
C0798707|T201|COMP|15540-8|LNC|Malus sylvestris tree Ab.IgE.RAST class|Malus sylvestris tree Ab.IgE.RAST class
C0798708|T201|COMP|15541-6|LNC|Prunus armeniaca Ab.IgE.RAST class|Prunus armeniaca Ab.IgE.RAST class
C0798709|T201|COMP|15542-4|LNC|Maranta arundinacea Ab.IgE.RAST class|Maranta arundinacea Ab.IgE.RAST class
C0798710|T201|COMP|15543-2|LNC|Cynara scolymus Ab.IgE.RAST class|Cynara scolymus Ab.IgE.RAST class
C0798711|T201|COMP|15544-0|LNC|Ascaris sp Ab.IgE.RAST class|Ascaris sp Ab.IgE.RAST class
C0798712|T201|COMP|15545-7|LNC|Fraxinus velutina Ab.IgE.RAST class|Fraxinus velutina Ab.IgE.RAST class
C0798713|T201|COMP|15546-5|LNC|Fraxinus americana Ab.IgE.RAST class|Fraxinus americana Ab.IgE.RAST class
C0798714|T201|COMP|15547-3|LNC|Asparagus officinalis Ab.IgE.RAST class|Asparagus officinalis Ab.IgE.RAST class
C0798716|T201|COMP|15549-9|LNC|Aspergillus fumigatus Ab.IgE.RAST class|Aspergillus fumigatus Ab.IgE.RAST class
C0798717|T201|COMP|15550-7|LNC|Aspergillus niger Ab.IgE.RAST class|Aspergillus niger Ab.IgE.RAST class
C0798718|T201|COMP|15551-5|LNC|Persea americana Ab.IgE.RAST class|Persea americana Ab.IgE.RAST class
C0798720|T201|COMP|15553-1|LNC|Phyllostachys pubescens Ab.IgE.RAST class|Phyllostachys pubescens Ab.IgE.RAST class
C0798721|T201|COMP|15554-9|LNC|Musa spp Ab.IgE.RAST class|Musa spp Ab.IgE.RAST class
C0798722|T201|COMP|15555-6|LNC|Hordeum vulgare Ab.IgE.RAST class|Hordeum vulgare Ab.IgE.RAST class
C0798723|T201|COMP|15556-4|LNC|Hordeum vulgare pollen Ab.IgE.RAST class|Hordeum vulgare pollen Ab.IgE.RAST class
C0798724|T201|COMP|15557-2|LNC|Ocimum basilicum Ab.IgE.RAST class|Ocimum basilicum Ab.IgE.RAST class
C0798725|T201|COMP|15558-0|LNC|Micropterus salmoides Ab.IgE.RAST class|Micropterus salmoides Ab.IgE.RAST class
C0798726|T201|COMP|15559-8|LNC|Bassia hyssopifolia Ab.IgE.RAST class|Bassia hyssopifolia Ab.IgE.RAST class
C0798727|T201|COMP|15560-6|LNC|Myrica spp Ab.IgE.RAST class|Myrica spp Ab.IgE.RAST class
C0798728|T201|COMP|15561-4|LNC|Laurus nobilis Ab.IgE.RAST class|Laurus nobilis Ab.IgE.RAST class
C0798729|T201|COMP|15562-2|LNC|Ricinus communis Ab.IgE.RAST class|Ricinus communis Ab.IgE.RAST class
C0798730|T201|COMP|15563-0|LNC|Coffee bean green Ab.IgE.RAST class|Coffee bean green Ab.IgE.RAST class
C0798731|T201|COMP|15564-8|LNC|Bean green Ab.IgE.RAST class|Bean green Ab.IgE.RAST class
C0798732|T201|COMP|15565-5|LNC|Bean kidney red Ab.IgE.RAST class|Bean kidney red Ab.IgE.RAST class
C0798733|T201|COMP|15566-3|LNC|Phaseolus limensis Ab.IgE.RAST class|Phaseolus limensis Ab.IgE.RAST class
C0798734|T201|COMP|15567-1|LNC|Bean pinto Ab.IgE.RAST class|Bean pinto Ab.IgE.RAST class
C0798735|T201|COMP|15568-9|LNC|Glycine max Ab.IgE.RAST class|Glycine max Ab.IgE.RAST class
C0798736|T201|COMP|15569-7|LNC|Bean white Ab.IgE.RAST class|Bean white Ab.IgE.RAST class
C0798737|T201|COMP|15570-5|LNC|Apis mellifera Ab.IgE.RAST class|Apis mellifera Ab.IgE.RAST class
C0798738|T201|COMP|15571-3|LNC|Fagus grandifolia Ab.IgE.RAST class|Fagus grandifolia Ab.IgE.RAST class
C0798739|T201|COMP|15572-1|LNC|Beef Ab.IgE.RAST class|Beef Ab.IgE.RAST class
C0798740|T201|COMP|15573-9|LNC|Beet Ab.IgE.RAST class|Beet Ab.IgE.RAST class
C0798741|T201|COMP|15574-7|LNC|Beta vulgaris seed Ab.IgE.RAST class|Beta vulgaris seed Ab.IgE.RAST class
C0798742|T201|COMP|15575-4|LNC|Trogoderma angustum Ab.IgE.RAST class|Trogoderma angustum Ab.IgE.RAST class
C0798743|T201|COMP|15576-2|LNC|Lactalbumin beta Ab.IgE.RAST class|Lactalbumin beta Ab.IgE.RAST class
C0798744|T201|COMP|15577-0|LNC|Beta lactoglobulin Ab.IgE.RAST class|Beta lactoglobulin Ab.IgE.RAST class
C0798745|T201|COMP|15578-8|LNC|Birch Ab.IgE.RAST class|Birch Ab.IgE.RAST class
C0798746|T201|COMP|15579-6|LNC|Betula verrucosa Ab.IgE.RAST class|Betula verrucosa Ab.IgE.RAST class
C0798747|T201|COMP|15580-4|LNC|Rubus fruticosus Ab.IgE.RAST class|Rubus fruticosus Ab.IgE.RAST class
C0798748|T201|COMP|15581-2|LNC|Blomia tropicalis Ab.IgE.RAST class|Blomia tropicalis Ab.IgE.RAST class
C0798749|T201|COMP|15582-0|LNC|Chironomus thummi Ab.IgE.RAST class|Chironomus thummi Ab.IgE.RAST class
C0798750|T201|COMP|15583-8|LNC|Vaccinium myrtillus Ab.IgE.RAST class|Vaccinium myrtillus Ab.IgE.RAST class
C0798751|T201|COMP|15584-6|LNC|Botrytis cinerea Ab.IgE.RAST class|Botrytis cinerea Ab.IgE.RAST class
C0798752|T201|COMP|15585-3|LNC|Acer negundo Ab.IgE.RAST class|Acer negundo Ab.IgE.RAST class
C0798753|T201|COMP|15586-1|LNC|Bertholletia excelsa Ab.IgE.RAST class|Bertholletia excelsa Ab.IgE.RAST class
C0798754|T201|COMP|15587-9|LNC|Brassica oleracea var italica Ab.IgE.RAST class|Brassica oleracea var italica Ab.IgE.RAST class
C0798755|T201|COMP|15588-7|LNC|Bromelin Ab.IgE.RAST class|Bromelin Ab.IgE.RAST class
C0798756|T201|COMP|15589-5|LNC|Brassica oleracea var gemmifera Ab.IgE.RAST class|Brassica oleracea var gemmifera Ab.IgE.RAST class
C0798757|T201|COMP|15590-3|LNC|Bovine serum albumin Ab.IgE.RAST class|Bovine serum albumin Ab.IgE.RAST class
C0798758|T201|COMP|15591-1|LNC|Fagopyrum esculentum Ab.IgE.RAST class|Fagopyrum esculentum Ab.IgE.RAST class
C0798759|T201|COMP|15592-9|LNC|Budgerigar feather Ab.IgE.RAST class|Budgerigar feather Ab.IgE.RAST class
C0798760|T201|COMP|15593-7|LNC|Bombus terrestris Ab.IgE.RAST class|Bombus terrestris Ab.IgE.RAST class
C0798761|T201|COMP|15594-5|LNC|Hymenoclea salsola Ab.IgE.RAST class|Hymenoclea salsola Ab.IgE.RAST class
C0798762|T201|COMP|15595-2|LNC|Iva xanthifolia Ab.IgE.RAST class|Iva xanthifolia Ab.IgE.RAST class
C0798762|T201|COMP|21256-3|LNC|Iva xanthifolia Ab.IgE.RAST class|Iva xanthifolia Ab.IgE.RAST class
C0798762|T201|COMP|21257-1|LNC|Iva xanthifolia Ab.IgE.RAST class|Iva xanthifolia Ab.IgE.RAST class
C0798763|T201|COMP|15596-0|LNC|Brassica oleracea var capitata Ab.IgE.RAST class|Brassica oleracea var capitata Ab.IgE.RAST class
C0798765|T201|COMP|15598-6|LNC|Canary feather Ab.IgE.RAST class|Canary feather Ab.IgE.RAST class
C0798766|T201|COMP|15599-4|LNC|Candida albicans Ab.IgE.RAST class|Candida albicans Ab.IgE.RAST class
C0798768|T201|COMP|15601-8|LNC|Averrhoa carambola Ab.IgE.RAST class|Averrhoa carambola Ab.IgE.RAST class
C0798769|T201|COMP|15602-6|LNC|Carum carvi Ab.IgE.RAST class|Carum carvi Ab.IgE.RAST class
C0798770|T201|COMP|15603-4|LNC|Amaranthus palmeri Ab.IgE.RAST class|Amaranthus palmeri Ab.IgE.RAST class
C0798771|T201|COMP|15604-2|LNC|Ceratonia siliqua Ab.IgE.RAST class|Ceratonia siliqua Ab.IgE.RAST class
C0798772|T201|COMP|15605-9|LNC|Daucus carota Ab.IgE.RAST class|Daucus carota Ab.IgE.RAST class
C0798773|T201|COMP|15606-7|LNC|Casein Ab.IgE.RAST class|Casein Ab.IgE.RAST class
C0798774|T201|COMP|15607-5|LNC|Anacardium occidentale Ab.IgE.RAST class|Anacardium occidentale Ab.IgE.RAST class
C0798775|T201|COMP|15608-3|LNC|Cat Ab.IgE.RAST class|Cat Ab.IgE.RAST class
C0798776|T201|COMP|15609-1|LNC|Cat dander Ab.IgE.RAST class|Cat dander Ab.IgE.RAST class
C0798777|T201|COMP|15610-9|LNC|Cat epithelium Ab.IgE.RAST class|Cat epithelium Ab.IgE.RAST class
C0798778|T201|COMP|15611-7|LNC|Ictalurus punctatus Ab.IgE.RAST class|Ictalurus punctatus Ab.IgE.RAST class
C0798779|T201|COMP|15612-5|LNC|Brassica oleracea var botrytis Ab.IgE.RAST class|Brassica oleracea var botrytis Ab.IgE.RAST class
C0798780|T201|COMP|15613-3|LNC|Cedar italian Ab.IgE.RAST class|Cedar italian Ab.IgE.RAST class
C0798781|T201|COMP|15614-1|LNC|Cryptomeria japonica Ab.IgE.RAST class|Cryptomeria japonica Ab.IgE.RAST class
C0798782|T201|COMP|15615-8|LNC|Juniperus sabinoides Ab.IgE.RAST class|Juniperus sabinoides Ab.IgE.RAST class
C0798783|T201|COMP|15616-6|LNC|Juniperus virginiana Ab.IgE.RAST class|Juniperus virginiana Ab.IgE.RAST class
C0798784|T201|COMP|15617-4|LNC|Tamarix spp Ab.IgE.RAST class|Tamarix spp Ab.IgE.RAST class
C0798785|T201|COMP|15618-2|LNC|Apium graveolens Ab.IgE.RAST class|Apium graveolens Ab.IgE.RAST class
C0798786|T201|COMP|15619-0|LNC|Acremonium sp Ab.IgE.RAST class|Acremonium sp Ab.IgE.RAST class
C0798787|T201|COMP|15620-8|LNC|Chaetomium globosum Ab.IgE.RAST class|Chaetomium globosum Ab.IgE.RAST class
C0798788|T201|COMP|15621-6|LNC|Matricaria chamomilla Ab.IgE.RAST class|Matricaria chamomilla Ab.IgE.RAST class
C0798789|T201|COMP|15622-4|LNC|Cheese American Ab.IgE.RAST class|Cheese American Ab.IgE.RAST class
C0798790|T201|COMP|15623-2|LNC|Cheese cheddar type Ab.IgE.RAST class|Cheese cheddar type Ab.IgE.RAST class
C0798791|T201|COMP|15624-0|LNC|Cheese cottage Ab.IgE.RAST class|Cheese cottage Ab.IgE.RAST class
C0798792|T201|COMP|15625-7|LNC|Cheese mozzarella Ab.IgE.RAST class|Cheese mozzarella Ab.IgE.RAST class
C0798793|T201|COMP|15626-5|LNC|Cheese parmesan Ab.IgE.RAST class|Cheese parmesan Ab.IgE.RAST class
C0798794|T201|COMP|15627-3|LNC|Cheese swiss Ab.IgE.RAST class|Cheese swiss Ab.IgE.RAST class
C0798795|T201|COMP|15628-1|LNC|Prunus avium Ab.IgE.RAST class|Prunus avium Ab.IgE.RAST class
C0798797|T201|COMP|15630-7|LNC|Aesculus hippocastanum Ab.IgE.RAST class|Aesculus hippocastanum Ab.IgE.RAST class
C0798798|T201|COMP|15629-9|LNC|Castanea sativa Ab.IgE.RAST class|Castanea sativa Ab.IgE.RAST class
C0798799|T201|COMP|15632-3|LNC|Castanea sativa pollen Ab.IgE.RAST class|Castanea sativa pollen Ab.IgE.RAST class
C0798800|T201|COMP|15633-1|LNC|Chicken feather Ab.IgE.RAST class|Chicken feather Ab.IgE.RAST class
C0798801|T201|COMP|15634-9|LNC|Chicken meat Ab.IgE.RAST class|Chicken meat Ab.IgE.RAST class
C0798802|T201|COMP|15635-6|LNC|Cichorium intybus Ab.IgE.RAST class|Cichorium intybus Ab.IgE.RAST class
C0798803|T201|COMP|15636-4|LNC|Chinchilla Ab.IgE.RAST class|Chinchilla Ab.IgE.RAST class
C0798804|T201|COMP|15637-2|LNC|Chloramin T Ab.IgE.RAST class|Chloramin T Ab.IgE.RAST class
C0798805|T201|COMP|15638-0|LNC|Chortoglyphus arcuatus Ab.IgE.RAST class|Chortoglyphus arcuatus Ab.IgE.RAST class
C0798806|T201|COMP|15639-8|LNC|Chymofast Ab.IgE.RAST class|Chymofast Ab.IgE.RAST class
C0798807|T201|COMP|15640-6|LNC|Chymopapain Ab.IgE.RAST class|Chymopapain Ab.IgE.RAST class
C0798808|T201|COMP|15641-4|LNC|Cinnamomum spp Ab.IgE.RAST class|Cinnamomum spp Ab.IgE.RAST class
C0798809|T201|COMP|15642-2|LNC|Cladosporium herbarum Ab.IgE.RAST class|Cladosporium herbarum Ab.IgE.RAST class
C0798810|T201|COMP|15643-0|LNC|Ruditapes spp Ab.IgE.RAST class|Ruditapes spp Ab.IgE.RAST class
C0798811|T201|COMP|15644-8|LNC|Syzygium aromaticum Ab.IgE.RAST class|Syzygium aromaticum Ab.IgE.RAST class
C0798812|T201|COMP|15645-5|LNC|Clover Ab.IgE.RAST class|Clover Ab.IgE.RAST class
C0798813|T201|COMP|15646-3|LNC|Xanthium commune Ab.IgE.RAST class|Xanthium commune Ab.IgE.RAST class
C0798814|T201|COMP|15647-1|LNC|Blatella germanica Ab.IgE.RAST class|Blatella germanica Ab.IgE.RAST class
C0798815|T201|COMP|15597-8|LNC|Theobroma cacao Ab.IgE.RAST class|Theobroma cacao Ab.IgE.RAST class
C0798816|T201|COMP|15649-7|LNC|Cocos nucifera Ab.IgE.RAST class|Cocos nucifera Ab.IgE.RAST class
C0798817|T201|COMP|15650-5|LNC|Gadus morhua Ab.IgE.RAST class|Gadus morhua Ab.IgE.RAST class
C0798818|T201|COMP|15651-3|LNC|Coffea spp Ab.IgE.RAST class|Coffea spp Ab.IgE.RAST class
C0798819|T201|COMP|15652-1|LNC|Cola Ab.IgE.RAST class|Cola Ab.IgE.RAST class
C0798821|T201|COMP|15654-7|LNC|Zea mays pollen Ab.IgE.RAST class|Zea mays pollen Ab.IgE.RAST class
C0798822|T201|COMP|15655-4|LNC|Cotton cultivated Ab.IgE.RAST class|Cotton cultivated Ab.IgE.RAST class
C0798823|T201|COMP|15656-2|LNC|Cotton fibers Ab.IgE.RAST class|Cotton fibers Ab.IgE.RAST class
C0798824|T201|COMP|15657-0|LNC|Cotton western Ab.IgE.RAST class|Cotton western Ab.IgE.RAST class
C0798825|T201|COMP|15658-8|LNC|Cottonseed Ab.IgE.RAST class|Cottonseed Ab.IgE.RAST class
C0798826|T201|COMP|15659-6|LNC|Populus deltoides Ab.IgE.RAST class|Populus deltoides Ab.IgE.RAST class
C0798827|T201|COMP|15660-4|LNC|Populus fremontii Ab.IgE.RAST class|Populus fremontii Ab.IgE.RAST class
C0798828|T201|COMP|15661-2|LNC|Cow dander Ab.IgE.RAST class|Cow dander Ab.IgE.RAST class
C0798829|T201|COMP|15662-0|LNC|Cow epithelium Ab.IgE.RAST class|Cow epithelium Ab.IgE.RAST class
C0798830|T201|COMP|15663-8|LNC|Cancer pagurus Ab.IgE.RAST class|Cancer pagurus Ab.IgE.RAST class
C0798831|T201|COMP|15664-6|LNC|Vaccinium oxycoccos Ab.IgE.RAST class|Vaccinium oxycoccos Ab.IgE.RAST class
C0798832|T201|COMP|15665-3|LNC|Astacus astacus Ab.IgE.RAST class|Astacus astacus Ab.IgE.RAST class
C0798833|T201|COMP|15666-1|LNC|Cryptococcus terreus Ab.IgE.RAST class|Cryptococcus terreus Ab.IgE.RAST class
C0798834|T201|COMP|15667-9|LNC|Cucumis sativus Ab.IgE.RAST class|Cucumis sativus Ab.IgE.RAST class
C0798835|T201|COMP|15668-7|LNC|Curry Ab.IgE.RAST class|Curry Ab.IgE.RAST class
C0798836|T201|COMP|15669-5|LNC|Curvularia lunata Ab.IgE.RAST class|Curvularia lunata Ab.IgE.RAST class
C0798837|T201|COMP|15670-3|LNC|Curvularia specifera Ab.IgE.RAST class|Curvularia specifera Ab.IgE.RAST class
C0798838|T201|COMP|15671-1|LNC|Cupressus arizonica Ab.IgE.RAST class|Cupressus arizonica Ab.IgE.RAST class
C0798839|T201|COMP|15672-9|LNC|Taxodium distichum Ab.IgE.RAST class|Taxodium distichum Ab.IgE.RAST class
C0798840|T201|COMP|15673-7|LNC|Cupressus sempervirens Ab.IgE.RAST class|Cupressus sempervirens Ab.IgE.RAST class
C0798841|T201|COMP|15674-5|LNC|Bellis perennis Ab.IgE.RAST class|Bellis perennis Ab.IgE.RAST class
C0798842|T201|COMP|15675-2|LNC|Chrysanthemum leucanthemum Ab.IgE.RAST class|Chrysanthemum leucanthemum Ab.IgE.RAST class
C0798843|T201|COMP|15676-0|LNC|Taraxacum vulgare Ab.IgE.RAST class|Taraxacum vulgare Ab.IgE.RAST class
C0798844|T201|COMP|15677-8|LNC|Daphnia Ab.IgE.RAST class|Daphnia Ab.IgE.RAST class
C0798845|T201|COMP|15678-6|LNC|Phoenix canariensis pollen Ab.IgE.RAST class|Phoenix canariensis pollen Ab.IgE.RAST class
C0798846|T201|COMP|15679-4|LNC|Deer epithelium Ab.IgE.RAST class|Deer epithelium Ab.IgE.RAST class
C0798847|T201|COMP|15680-2|LNC|Dermatophagoides farinae Ab.IgE.RAST class|Dermatophagoides farinae Ab.IgE.RAST class
C0798848|T201|COMP|15681-0|LNC|Dermatophagoides microceras Ab.IgE.RAST class|Dermatophagoides microceras Ab.IgE.RAST class
C0798849|T201|COMP|15682-8|LNC|Dermatophagoides pteronyssinus Ab.IgE.RAST class|Dermatophagoides pteronyssinus Ab.IgE.RAST class
C0798850|T201|COMP|15683-6|LNC|Anethum graveolens Ab.IgE.RAST class|Anethum graveolens Ab.IgE.RAST class
C0798851|T201|COMP|15684-4|LNC|Rumex crispus Ab.IgE.RAST class|Rumex crispus Ab.IgE.RAST class
C0798852|T201|COMP|15685-1|LNC|Dog dander Ab.IgE.RAST class|Dog dander Ab.IgE.RAST class
C0798853|T201|COMP|15686-9|LNC|Dog epithelium Ab.IgE.RAST class|Dog epithelium Ab.IgE.RAST class
C0798854|T201|COMP|15687-7|LNC|Duck feather Ab.IgE.RAST class|Duck feather Ab.IgE.RAST class
C0798855|T201|COMP|15688-5|LNC|Echinococcus sp Ab.IgE.RAST class|Echinococcus sp Ab.IgE.RAST class
C0798856|T201|COMP|15689-3|LNC|Egg white Ab.IgE.RAST class|Egg white Ab.IgE.RAST class
C0798857|T201|COMP|15690-1|LNC|Egg whole Ab.IgE.RAST class|Egg whole Ab.IgE.RAST class
C0798858|T201|COMP|15691-9|LNC|Egg yolk Ab.IgE.RAST class|Egg yolk Ab.IgE.RAST class
C0798859|T201|COMP|15692-7|LNC|Solanum melongena Ab.IgE.RAST class|Solanum melongena Ab.IgE.RAST class
C0798860|T201|COMP|15693-5|LNC|Iva ciliata Ab.IgE.RAST class|Iva ciliata Ab.IgE.RAST class
C0798862|T201|COMP|15694-3|LNC|Sambucus nigra Ab.IgE.RAST class|Sambucus nigra Ab.IgE.RAST class
C0798863|T201|COMP|15696-8|LNC|Elk meat Ab.IgE.RAST class|Elk meat Ab.IgE.RAST class
C0798864|T201|COMP|15697-6|LNC|Ulmus americana Ab.IgE.RAST class|Ulmus americana Ab.IgE.RAST class
C0798865|T201|COMP|15698-4|LNC|Ulmus pumila Ab.IgE.RAST class|Ulmus pumila Ab.IgE.RAST class
C0798866|T201|COMP|15699-2|LNC|Cichorium endivia Ab.IgE.RAST class|Cichorium endivia Ab.IgE.RAST class
C0798867|T201|COMP|15700-8|LNC|Epicoccum purpurascens Ab.IgE.RAST class|Epicoccum purpurascens Ab.IgE.RAST class
C0798868|T201|COMP|15701-6|LNC|Epidermophyton floccosum Ab.IgE.RAST class|Epidermophyton floccosum Ab.IgE.RAST class
C0798869|T201|COMP|15702-4|LNC|Ethylene oxide Ab.IgE.RAST class|Ethylene oxide Ab.IgE.RAST class
C0798870|T201|COMP|15703-2|LNC|Eucalyptus spp Ab.IgE.RAST class|Eucalyptus spp Ab.IgE.RAST class
C0798871|T201|COMP|15704-0|LNC|Euroglyphus maynei Ab.IgE.RAST class|Euroglyphus maynei Ab.IgE.RAST class
C0798872|T201|COMP|15705-7|LNC|Anthemis cotula Ab.IgE.RAST class|Anthemis cotula Ab.IgE.RAST class
C0798873|T201|COMP|15706-5|LNC|Foeniculum vulgare fresh Ab.IgE.RAST class|Foeniculum vulgare fresh Ab.IgE.RAST class
C0798874|T201|COMP|15707-3|LNC|Foeniculum vulgare seed Ab.IgE.RAST class|Foeniculum vulgare seed Ab.IgE.RAST class
C0798875|T201|COMP|15708-1|LNC|Ferret epithelium Ab.IgE.RAST class|Ferret epithelium Ab.IgE.RAST class
C0798876|T201|COMP|15709-9|LNC|Festuca elatior Ab.IgE.RAST class|Festuca elatior Ab.IgE.RAST class
C0798877|T201|COMP|15710-7|LNC|Finch feather Ab.IgE.RAST class|Finch feather Ab.IgE.RAST class
C0798878|T201|COMP|15711-5|LNC|Pseudotsuga taxifolia Ab.IgE.RAST class|Pseudotsuga taxifolia Ab.IgE.RAST class
C0798879|T201|COMP|15712-3|LNC|Kochia scoparia Ab.IgE.RAST class|Kochia scoparia Ab.IgE.RAST class
C0798880|T201|COMP|15713-1|LNC|Fiscus sp Ab.IgE.RAST class|Fiscus sp Ab.IgE.RAST class
C0798881|T201|COMP|15714-9|LNC|Ctenocephalides sp Ab.IgE.RAST class|Ctenocephalides sp Ab.IgE.RAST class
C0798882|T201|COMP|15715-6|LNC|Flounder Ab.IgE.RAST class|Flounder Ab.IgE.RAST class
C0798883|T201|COMP|15716-4|LNC|Simulium venustum Ab.IgE.RAST class|Simulium venustum Ab.IgE.RAST class
C0798884|T201|COMP|15717-2|LNC|Tabanus spp Ab.IgE.RAST class|Tabanus spp Ab.IgE.RAST class
C0798885|T201|COMP|15718-0|LNC|Formaldehyde Ab.IgE.RAST class|Formaldehyde Ab.IgE.RAST class
C0798886|T201|COMP|15719-8|LNC|Fox Ab.IgE.RAST class|Fox Ab.IgE.RAST class
C0798887|T201|COMP|15720-6|LNC|Alopercurus pratensis Ab.IgE.RAST class|Alopercurus pratensis Ab.IgE.RAST class
C0798888|T201|COMP|15721-4|LNC|Fusarium culmorum Ab.IgE.RAST class|Fusarium culmorum Ab.IgE.RAST class
C0798889|T201|COMP|15722-2|LNC|Fusarium moniliforme Ab.IgE.RAST class|Fusarium moniliforme Ab.IgE.RAST class
C0798890|T201|COMP|15723-0|LNC|Fusarium solani Ab.IgE.RAST class|Fusarium solani Ab.IgE.RAST class
C0798891|T201|COMP|15724-8|LNC|Allium sativum Ab.IgE.RAST class|Allium sativum Ab.IgE.RAST class
C0798892|T201|COMP|15725-5|LNC|Gelatin Ab.IgE.RAST class|Gelatin Ab.IgE.RAST class
C0798893|T201|COMP|15726-3|LNC|Geotrichum candidum Ab.IgE.RAST class|Geotrichum candidum Ab.IgE.RAST class
C0798894|T201|COMP|15727-1|LNC|Gerbil Ab.IgE.RAST class|Gerbil Ab.IgE.RAST class
C0798895|T201|COMP|15728-9|LNC|Zingiber officinale Ab.IgE.RAST class|Zingiber officinale Ab.IgE.RAST class
C0798896|T201|COMP|15729-7|LNC|Gluten Ab.IgE.RAST class|Gluten Ab.IgE.RAST class
C0798897|T201|COMP|15730-5|LNC|Glycyphagus domesticus Ab.IgE.RAST class|Glycyphagus domesticus Ab.IgE.RAST class
C0798898|T201|COMP|15731-3|LNC|Goat epithelium Ab.IgE.RAST class|Goat epithelium Ab.IgE.RAST class
C0798899|T201|COMP|15732-1|LNC|Goat milk Ab.IgE.RAST class|Goat milk Ab.IgE.RAST class
C0798900|T201|COMP|15733-9|LNC|Solidago virgaurea Ab.IgE.RAST class|Solidago virgaurea Ab.IgE.RAST class
C0798901|T201|COMP|15734-7|LNC|Goose feather Ab.IgE.RAST class|Goose feather Ab.IgE.RAST class
C0798902|T201|COMP|15735-4|LNC|Vitis vinifera Ab.IgE.RAST class|Vitis vinifera Ab.IgE.RAST class
C0798903|T201|COMP|15736-2|LNC|Citrus paradisis Ab.IgE.RAST class|Citrus paradisis Ab.IgE.RAST class
C0798904|T201|COMP|15737-0|LNC|Paspalum notatum Ab.IgE.RAST class|Paspalum notatum Ab.IgE.RAST class
C0798905|T201|COMP|15738-8|LNC|Cynodon dactylon Ab.IgE.RAST class|Cynodon dactylon Ab.IgE.RAST class
C0798906|T201|COMP|15739-6|LNC|Poa compressa Ab.IgE.RAST class|Poa compressa Ab.IgE.RAST class
C0798907|T201|COMP|15740-4|LNC|Bromus inermis Ab.IgE.RAST class|Bromus inermis Ab.IgE.RAST class
C0798908|T201|COMP|15741-2|LNC|Arrhenatherum elatius Ab.IgE.RAST class|Arrhenatherum elatius Ab.IgE.RAST class
C0798909|T201|COMP|15742-0|LNC|Bouteloua gracilis Ab.IgE.RAST class|Bouteloua gracilis Ab.IgE.RAST class
C0798910|T201|COMP|15743-8|LNC|Sorghum halepense Ab.IgE.RAST class|Sorghum halepense Ab.IgE.RAST class
C0798911|T201|COMP|15744-6|LNC|Poa pratensis Ab.IgE.RAST class|Poa pratensis Ab.IgE.RAST class
C0798912|T201|COMP|15745-3|LNC|Grass koehlers Ab.IgE.RAST class|Grass koehlers Ab.IgE.RAST class
C0798913|T201|COMP|15746-1|LNC|Dactylis glomerata Ab.IgE.RAST class|Dactylis glomerata Ab.IgE.RAST class
C0798914|T201|COMP|15747-9|LNC|Agropyron repens Ab.IgE.RAST class|Agropyron repens Ab.IgE.RAST class
C0798915|T201|COMP|15748-7|LNC|Agrostis stolonifera Ab.IgE.RAST class|Agrostis stolonifera Ab.IgE.RAST class
C0798918|T201|COMP|15751-1|LNC|Elymus triticoides Ab.IgE.RAST class|Elymus triticoides Ab.IgE.RAST class
C0798919|T201|COMP|15752-9|LNC|Distichlis spicata Ab.IgE.RAST class|Distichlis spicata Ab.IgE.RAST class
C0798920|T201|COMP|15753-7|LNC|Grass sorghum Ab.IgE.RAST class|Grass sorghum Ab.IgE.RAST class
C0798921|T201|COMP|15754-5|LNC|Sorghum sudanense Ab.IgE.RAST class|Sorghum sudanense Ab.IgE.RAST class
C0798922|T201|COMP|15755-2|LNC|Anthoxanthum odoratum Ab.IgE.RAST class|Anthoxanthum odoratum Ab.IgE.RAST class
C0798923|T201|COMP|15756-0|LNC|Holcus lanatus Ab.IgE.RAST class|Holcus lanatus Ab.IgE.RAST class
C0798924|T201|COMP|15757-8|LNC|Cyamopsis tetragonoloba Ab.IgE.RAST class|Cyamopsis tetragonoloba Ab.IgE.RAST class
C0798925|T201|COMP|15758-6|LNC|Psidium guajava Ab.IgE.RAST class|Psidium guajava Ab.IgE.RAST class
C0798926|T201|COMP|15759-4|LNC|Guinea pig epithelium Ab.IgE.RAST class|Guinea pig epithelium Ab.IgE.RAST class
C0798927|T201|COMP|15760-2|LNC|Gum arabic Ab.IgE.RAST class|Gum arabic Ab.IgE.RAST class
C0798929|T201|COMP|15762-8|LNC|Celtis occidentalis Ab.IgE.RAST class|Celtis occidentalis Ab.IgE.RAST class
C0798930|T201|COMP|15763-6|LNC|Melanogrammus aeglefinus Ab.IgE.RAST class|Melanogrammus aeglefinus Ab.IgE.RAST class
C0798931|T201|COMP|15764-4|LNC|Hippoglossus hippoglossus Ab.IgE.RAST class|Hippoglossus hippoglossus Ab.IgE.RAST class
C0798932|T201|COMP|15765-1|LNC|Hamster epithelium Ab.IgE.RAST class|Hamster epithelium Ab.IgE.RAST class
C0798933|T201|COMP|15766-9|LNC|Corylus avellana Ab.IgE.RAST class|Corylus avellana Ab.IgE.RAST class
C0798934|T201|COMP|15767-7|LNC|Corylus avellana pollen Ab.IgE.RAST class|Corylus avellana pollen Ab.IgE.RAST class
C0798936|T201|COMP|15769-3|LNC|Setomelanomma rostrata Ab.IgE.RAST class|Setomelanomma rostrata Ab.IgE.RAST class
C0798937|T201|COMP|15770-1|LNC|Tsuga canadensis Ab.IgE.RAST class|Tsuga canadensis Ab.IgE.RAST class
C0798938|T201|COMP|15771-9|LNC|Amaranthus tuberculatus Ab.IgE.RAST class|Amaranthus tuberculatus Ab.IgE.RAST class
C0798939|T201|COMP|15772-7|LNC|Clupea harengus Ab.IgE.RAST class|Clupea harengus Ab.IgE.RAST class
C0798942|T201|COMP|15775-0|LNC|Carya laciniosa Ab.IgE.RAST class|Carya laciniosa Ab.IgE.RAST class
C0798943|T201|COMP|15776-8|LNC|Carya tomentosa Ab.IgE.RAST class|Carya tomentosa Ab.IgE.RAST class
C0798944|T201|COMP|15777-6|LNC|Honey Ab.IgE.RAST class|Honey Ab.IgE.RAST class
C0798945|T201|COMP|15778-4|LNC|Honeysuckle Ab.IgE.RAST class|Honeysuckle Ab.IgE.RAST class
C0798946|T201|COMP|15779-2|LNC|Humulus lupus Ab.IgE.RAST class|Humulus lupus Ab.IgE.RAST class
C0798947|T201|COMP|15780-0|LNC|Carpinus betulus Ab.IgE.RAST class|Carpinus betulus Ab.IgE.RAST class
C0798948|T201|COMP|15781-8|LNC|Hornet Ab.IgE.RAST class|Hornet Ab.IgE.RAST class
C0798949|T201|COMP|15782-6|LNC|Dolichovespula maculata Ab.IgE.RAST class|Dolichovespula maculata Ab.IgE.RAST class
C0798950|T201|COMP|15783-4|LNC|Dolichovespula arenaria Ab.IgE.RAST class|Dolichovespula arenaria Ab.IgE.RAST class
C0798951|T201|COMP|15784-2|LNC|Horse dander Ab.IgE.RAST class|Horse dander Ab.IgE.RAST class
C0798952|T201|COMP|15785-9|LNC|Horse epithelium Ab.IgE.RAST class|Horse epithelium Ab.IgE.RAST class
C0798953|T201|COMP|15786-7|LNC|Horse serum proteins Ab.IgE.RAST class|Horse serum proteins Ab.IgE.RAST class
C0798954|T201|COMP|15787-5|LNC|Armoracia rusticana Ab.IgE.RAST class|Armoracia rusticana Ab.IgE.RAST class
C0798955|T201|COMP|15788-3|LNC|House dust Ab.IgE.RAST class|House dust Ab.IgE.RAST class
C0798956|T201|COMP|15789-1|LNC|House dust Greer Ab.IgE.RAST class|House dust Greer Ab.IgE.RAST class
C0798957|T201|COMP|15790-9|LNC|House dust Hausstaub Ab.IgE.RAST class|House dust Hausstaub Ab.IgE.RAST class
C0798958|T201|COMP|15791-7|LNC|House dust Hollister Stier Ab.IgE.RAST class|House dust Hollister Stier Ab.IgE.RAST class
C0798959|T201|COMP|15792-5|LNC|Insulin bovine Ab.IgE.RAST class|Insulin bovine Ab.IgE.RAST class
C0798960|T201|COMP|15793-3|LNC|Insulin human Ab.IgE.RAST class|Insulin human Ab.IgE.RAST class
C0798961|T201|COMP|15794-1|LNC|Insulin porcine Ab.IgE.RAST class|Insulin porcine Ab.IgE.RAST class
C0798962|T201|COMP|15795-8|LNC|Allenrolfea occidentalis Ab.IgE.RAST class|Allenrolfea occidentalis Ab.IgE.RAST class
C0798965|T201|COMP|15798-2|LNC|Toluene diisocyanate (TDI) Ab.IgE.RAST class|Toluene diisocyanate (TDI) Ab.IgE.RAST class
C0798966|T201|COMP|15799-0|LNC|Ispaghula laxative Ab.IgE.RAST class|Ispaghula laxative Ab.IgE.RAST class
C0798967|T201|COMP|15800-6|LNC|Juniper Ab.IgE.RAST class|Juniper Ab.IgE.RAST class
C0798968|T201|COMP|15801-4|LNC|Kapok Ab.IgE.RAST class|Kapok Ab.IgE.RAST class
C0798969|T201|COMP|15802-2|LNC|Actinidia chinensis Ab.IgE.RAST class|Actinidia chinensis Ab.IgE.RAST class
C0798970|T201|COMP|15803-0|LNC|Lamb Ab.IgE.RAST class|Lamb Ab.IgE.RAST class
C0798971|T201|COMP|15804-8|LNC|Mutton Ab.IgE.RAST class|Mutton Ab.IgE.RAST class
C0798972|T201|COMP|15805-5|LNC|Chenopodium album Ab.IgE.RAST class|Chenopodium album Ab.IgE.RAST class
C0798973|T201|COMP|15806-3|LNC|Latex Ab.IgE.RAST class|Latex Ab.IgE.RAST class
C0798974|T201|COMP|15807-1|LNC|Latex glove extract Ab.IgE.RAST class|Latex glove extract Ab.IgE.RAST class
C0798975|T201|COMP|15808-9|LNC|Latex glove extract ammoniated Ab.IgE.RAST class|Latex glove extract ammoniated Ab.IgE.RAST class
C0798976|T201|COMP|15809-7|LNC|Latex glove extract buffered Ab.IgE.RAST class|Latex glove extract buffered Ab.IgE.RAST class
C0798977|T201|COMP|15810-5|LNC|Legume Ab.IgE.RAST class|Legume Ab.IgE.RAST class
C0798978|T201|COMP|15811-3|LNC|Citrus limon Ab.IgE.RAST class|Citrus limon Ab.IgE.RAST class
C0798980|T201|COMP|15813-9|LNC|Lens esculenta Ab.IgE.RAST class|Lens esculenta Ab.IgE.RAST class
C0798981|T201|COMP|15814-7|LNC|Lepidoglyphus destructor Ab.IgE.RAST class|Lepidoglyphus destructor Ab.IgE.RAST class
C0798982|T201|COMP|15815-4|LNC|Lactuca sativa Ab.IgE.RAST class|Lactuca sativa Ab.IgE.RAST class
C0798983|T201|COMP|15816-2|LNC|Syringa vulgaris Ab.IgE.RAST class|Syringa vulgaris Ab.IgE.RAST class
C0798984|T201|COMP|15817-0|LNC|Lilium longiflorum Ab.IgE.RAST class|Lilium longiflorum Ab.IgE.RAST class
C0798985|T201|COMP|15818-8|LNC|Citrus aurantifolia Ab.IgE.RAST class|Citrus aurantifolia Ab.IgE.RAST class
C0798986|T201|COMP|15819-6|LNC|Tilia cordata Ab.IgE.RAST class|Tilia cordata Ab.IgE.RAST class
C0798987|T201|COMP|15820-4|LNC|Liver beef Ab.IgE.RAST class|Liver beef Ab.IgE.RAST class
C0798988|T201|COMP|15821-2|LNC|Homarus gammarus Ab.IgE.RAST class|Homarus gammarus Ab.IgE.RAST class
C0798989|T201|COMP|15822-0|LNC|Palinurus spp Ab.IgE.RAST class|Palinurus spp Ab.IgE.RAST class
C0798990|T201|COMP|15823-8|LNC|Robinia pseudoacacia Ab.IgE.RAST class|Robinia pseudoacacia Ab.IgE.RAST class
C0798991|T201|COMP|15824-6|LNC|Lupinus spp Ab.IgE.RAST class|Lupinus spp Ab.IgE.RAST class
C0798992|T201|COMP|15825-3|LNC|Lycopodium spp Ab.IgE.RAST class|Lycopodium spp Ab.IgE.RAST class
C0798993|T201|COMP|15826-1|LNC|Lysozyme Ab.IgE.RAST class|Lysozyme Ab.IgE.RAST class
C0798994|T201|COMP|15827-9|LNC|Scomber scombrus Ab.IgE.RAST class|Scomber scombrus Ab.IgE.RAST class
C0798995|T201|COMP|15828-7|LNC|Scomber japonicus Ab.IgE.RAST class|Scomber japonicus Ab.IgE.RAST class
C0798996|T201|COMP|15829-5|LNC|Trachurus japonicus Ab.IgE.RAST class|Trachurus japonicus Ab.IgE.RAST class
C0798997|T201|COMP|15653-9|LNC|Zea mays Ab.IgE.RAST class|Zea mays Ab.IgE.RAST class
C0798998|T201|COMP|15831-1|LNC|Malt Ab.IgE.RAST class|Malt Ab.IgE.RAST class
C0798999|T201|COMP|15832-9|LNC|Mangifera indica Ab.IgE.RAST class|Mangifera indica Ab.IgE.RAST class
C0799000|T201|COMP|15833-7|LNC|Acer macrophyllum Ab.IgE.RAST class|Acer macrophyllum Ab.IgE.RAST class
C0799001|T201|COMP|15834-5|LNC|Acer rubrum Ab.IgE.RAST class|Acer rubrum Ab.IgE.RAST class
C0799002|T201|COMP|15835-2|LNC|Maple silver Ab.IgE.RAST class|Maple silver Ab.IgE.RAST class
C0799003|T201|COMP|15836-0|LNC|Maple sugar Ab.IgE.RAST class|Maple sugar Ab.IgE.RAST class
C0799004|T201|COMP|15837-8|LNC|Mare milk Ab.IgE.RAST class|Mare milk Ab.IgE.RAST class
C0799005|T201|COMP|15838-6|LNC|Origanum majorana Ab.IgE.RAST class|Origanum majorana Ab.IgE.RAST class
C0799006|T201|COMP|15839-4|LNC|Maxatase Ab.IgE.RAST class|Maxatase Ab.IgE.RAST class
C0799007|T201|COMP|15840-2|LNC|Lepidorhombus whiffiagonis Ab.IgE.RAST class|Lepidorhombus whiffiagonis Ab.IgE.RAST class
C0799008|T201|COMP|15841-0|LNC|Melaleuca leucadendron Ab.IgE.RAST class|Melaleuca leucadendron Ab.IgE.RAST class
C0799010|T201|COMP|15843-6|LNC|Prosopis juliflora Ab.IgE.RAST class|Prosopis juliflora Ab.IgE.RAST class
C0799011|T201|COMP|15844-4|LNC|Chenopodium ambrosioides Ab.IgE.RAST class|Chenopodium ambrosioides Ab.IgE.RAST class
C0799012|T201|COMP|15845-1|LNC|Cladotanytarsus lewisi Ab.IgE.RAST class|Cladotanytarsus lewisi Ab.IgE.RAST class
C0799013|T201|COMP|15846-9|LNC|Milk Ab.IgE.RAST class|Milk Ab.IgE.RAST class
C0799014|T201|COMP|15847-7|LNC|Cow milk boiled Ab.IgE.RAST class|Cow milk boiled Ab.IgE.RAST class
C0799015|T201|COMP|15848-5|LNC|Milk powder Ab.IgE.RAST class|Milk powder Ab.IgE.RAST class
C0799017|T201|COMP|15850-1|LNC|Setaria italica Ab.IgE.RAST class|Setaria italica Ab.IgE.RAST class
C0799018|T201|COMP|15851-9|LNC|Echinochloa crus-galli Ab.IgE.RAST class|Echinochloa crus-galli Ab.IgE.RAST class
C0799019|T201|COMP|15852-7|LNC|Mink epithelium Ab.IgE.RAST class|Mink epithelium Ab.IgE.RAST class
C0799020|T201|COMP|15853-5|LNC|Mentha piperita Ab.IgE.RAST class|Mentha piperita Ab.IgE.RAST class
C0799021|T201|COMP|15854-3|LNC|Cheese mold type Ab.IgE.RAST class|Cheese mold type Ab.IgE.RAST class
C0799022|T201|COMP|15855-0|LNC|Chrysonilia sitophila Ab.IgE.RAST class|Chrysonilia sitophila Ab.IgE.RAST class
C0799023|T201|COMP|15856-8|LNC|Aedes communis Ab.IgE.RAST class|Aedes communis Ab.IgE.RAST class
C0799024|T201|COMP|15857-6|LNC|Moth Ab.IgE.RAST class|Moth Ab.IgE.RAST class
C0799025|T201|COMP|15858-4|LNC|Ephestia kuehniella Ab.IgE.RAST class|Ephestia kuehniella Ab.IgE.RAST class
C0799026|T201|COMP|15859-2|LNC|Mouse epithelium Ab.IgE.RAST class|Mouse epithelium Ab.IgE.RAST class
C0799027|T201|COMP|15860-0|LNC|Mouse serum proteins Ab.IgE.RAST class|Mouse serum proteins Ab.IgE.RAST class
C0799028|T201|COMP|15861-8|LNC|Mouse urine proteins Ab.IgE.RAST class|Mouse urine proteins Ab.IgE.RAST class
C0799029|T201|COMP|15862-6|LNC|Mucor racemosus Ab.IgE.RAST class|Mucor racemosus Ab.IgE.RAST class
C0799030|T201|COMP|15863-4|LNC|Artemisia vulgaris Ab.IgE.RAST class|Artemisia vulgaris Ab.IgE.RAST class
C0799031|T201|COMP|15864-2|LNC|Morus alba Ab.IgE.RAST class|Morus alba Ab.IgE.RAST class
C0799032|T201|COMP|15865-9|LNC|Morus alba Ab.IgE.RAST class|Morus alba Ab.IgE.RAST class
C0799033|T201|COMP|15866-7|LNC|Agaricus hortensis Ab.IgE.RAST class|Agaricus hortensis Ab.IgE.RAST class
C0799034|T201|COMP|57882-3|LNC|Cucumis melo spp Ab.IgE.RAST class|Cucumis melo spp Ab.IgE.RAST class
C0799035|T201|COMP|15868-3|LNC|Mussel Ab.IgE.RAST class|Mussel Ab.IgE.RAST class
C0799036|T201|COMP|15869-1|LNC|Mytilus edulis Ab.IgE.RAST class|Mytilus edulis Ab.IgE.RAST class
C0799037|T201|COMP|15870-9|LNC|Mustard Ab.IgE.RAST class|Mustard Ab.IgE.RAST class
C0799038|T201|COMP|15871-7|LNC|Prunus persica var nucipersica Ab.IgE.RAST class|Prunus persica var nucipersica Ab.IgE.RAST class
C0799039|T201|COMP|15872-5|LNC|Urtica dioica Ab.IgE.RAST class|Urtica dioica Ab.IgE.RAST class
C0799040|T201|COMP|15873-3|LNC|Nigrospora sphaerica Ab.IgE.RAST class|Nigrospora sphaerica Ab.IgE.RAST class
C0799041|T201|COMP|15874-1|LNC|Nutmeg Ab.IgE.RAST class|Nutmeg Ab.IgE.RAST class
C0799043|T201|COMP|15876-6|LNC|Quercus kelloggii Ab.IgE.RAST class|Quercus kelloggii Ab.IgE.RAST class
C0799044|T201|COMP|15877-4|LNC|Quercus parvula Ab.IgE.RAST class|Quercus parvula Ab.IgE.RAST class
C0799045|T201|COMP|15878-2|LNC|Quercus gambelii Ab.IgE.RAST class|Quercus gambelii Ab.IgE.RAST class
C0799046|T201|COMP|15879-0|LNC|Chenopodium botrys Ab.IgE.RAST class|Chenopodium botrys Ab.IgE.RAST class
C0799048|T201|COMP|15881-6|LNC|Quercus rubra Ab.IgE.RAST class|Quercus rubra Ab.IgE.RAST class
C0799049|T201|COMP|15882-4|LNC|Quercus lobata Ab.IgE.RAST class|Quercus lobata Ab.IgE.RAST class
C0799050|T201|COMP|15880-8|LNC|Quercus virginiana Ab.IgE.RAST class|Quercus virginiana Ab.IgE.RAST class
C0799051|T201|COMP|15875-8|LNC|Quercus alba Ab.IgE.RAST class|Quercus alba Ab.IgE.RAST class
C0799053|T201|COMP|15886-5|LNC|Avena sativa cultivated Ab.IgE.RAST class|Avena sativa cultivated Ab.IgE.RAST class
C0799054|T201|COMP|15887-3|LNC|Avena sativa cultivated Ab.IgE.RAST class|Avena sativa cultivated Ab.IgE.RAST class
C0799055|T201|COMP|15888-1|LNC|Octopus vulgaris Ab.IgE.RAST class|Octopus vulgaris Ab.IgE.RAST class
C0799056|T201|COMP|15889-9|LNC|Oidiodendrum spp Ab.IgE.RAST class|Oidiodendrum spp Ab.IgE.RAST class
C0799057|T201|COMP|15890-7|LNC|Abelmoschus esculentus Ab.IgE.RAST class|Abelmoschus esculentus Ab.IgE.RAST class
C0799058|T201|COMP|15891-5|LNC|Olive Ab.IgE.RAST class|Olive Ab.IgE.RAST class
C0799059|T201|COMP|15892-3|LNC|Olea europaea pollen Ab.IgE.RAST class|Olea europaea pollen Ab.IgE.RAST class
C0799060|T201|COMP|15893-1|LNC|Allium cepa Ab.IgE.RAST class|Allium cepa Ab.IgE.RAST class
C0799061|T201|COMP|15894-9|LNC|Citrus sinensis Ab.IgE.RAST class|Citrus sinensis Ab.IgE.RAST class
C0799062|T201|COMP|15895-6|LNC|Origanum vulgare Ab.IgE.RAST class|Origanum vulgare Ab.IgE.RAST class
C0799063|T201|COMP|15896-4|LNC|Iris germanica var florentina Ab.IgE.RAST class|Iris germanica var florentina Ab.IgE.RAST class
C0799064|T201|COMP|15897-2|LNC|Ovalbumin Ab.IgE.RAST class|Ovalbumin Ab.IgE.RAST class
C0799065|T201|COMP|15898-0|LNC|Ovomucoid Ab.IgE.RAST class|Ovomucoid Ab.IgE.RAST class
C0799066|T201|COMP|15899-8|LNC|Ostrea edulis Ab.IgE.RAST class|Ostrea edulis Ab.IgE.RAST class
C0799067|T201|COMP|15900-4|LNC|Syagrus romanzoffianum Ab.IgE.RAST class|Syagrus romanzoffianum Ab.IgE.RAST class
C0799068|T201|COMP|15901-2|LNC|Carica papaya Ab.IgE.RAST class|Carica papaya Ab.IgE.RAST class
C0799069|T201|COMP|15902-0|LNC|Capsicum annuum Ab.IgE.RAST class|Capsicum annuum Ab.IgE.RAST class
C0799070|T201|COMP|15903-8|LNC|Parakeet feather Ab.IgE.RAST class|Parakeet feather Ab.IgE.RAST class
C0799071|T201|COMP|15904-6|LNC|Budgerigar droppings Ab.IgE.RAST class|Budgerigar droppings Ab.IgE.RAST class
C0799072|T201|COMP|15905-3|LNC|Budgerigar feather Ab.IgE.RAST class|Budgerigar feather Ab.IgE.RAST class
C0799073|T201|COMP|15906-1|LNC|Budgerigar serum proteins Ab.IgE.RAST class|Budgerigar serum proteins Ab.IgE.RAST class
C0799074|T201|COMP|15907-9|LNC|Parrot droppings Ab.IgE.RAST class|Parrot droppings Ab.IgE.RAST class
C0799075|T201|COMP|15908-7|LNC|Parrot feather Ab.IgE.RAST class|Parrot feather Ab.IgE.RAST class
C0799076|T201|COMP|15909-5|LNC|Parrot serum proteins Ab.IgE.RAST class|Parrot serum proteins Ab.IgE.RAST class
C0799077|T201|COMP|15910-3|LNC|Petroselinum crispum Ab.IgE.RAST class|Petroselinum crispum Ab.IgE.RAST class
C0799078|T201|COMP|15911-1|LNC|Pastinaca sativa Ab.IgE.RAST class|Pastinaca sativa Ab.IgE.RAST class
C0799079|T201|COMP|15912-9|LNC|Passiflora edulis Ab.IgE.RAST class|Passiflora edulis Ab.IgE.RAST class
C0799080|T201|COMP|15913-7|LNC|Pisum sativum Ab.IgE.RAST class|Pisum sativum Ab.IgE.RAST class
C0799081|T201|COMP|15914-5|LNC|Vigna sinensis Ab.IgE.RAST class|Vigna sinensis Ab.IgE.RAST class
C0799082|T201|COMP|15915-2|LNC|Cicer arietinus Ab.IgE.RAST class|Cicer arietinus Ab.IgE.RAST class
C0799083|T201|COMP|15916-0|LNC|Prunus persica Ab.IgE.RAST class|Prunus persica Ab.IgE.RAST class
C0799084|T201|COMP|15917-8|LNC|Arachis hypogaea Ab.IgE.RAST class|Arachis hypogaea Ab.IgE.RAST class
C0799085|T201|COMP|15918-6|LNC|Pyrus communis Ab.IgE.RAST class|Pyrus communis Ab.IgE.RAST class
C0799086|T201|COMP|15773-5|LNC|Carya illinoinensis nut Ab.IgE.RAST class|Carya illinoinensis nut Ab.IgE.RAST class
C0799087|T201|COMP|15774-3|LNC|Carya illinoinensis tree Ab.IgE.RAST class|Carya illinoinensis tree Ab.IgE.RAST class
C0799088|T201|COMP|15921-0|LNC|Penicillin G Ab.IgE.RAST class|Penicillin G Ab.IgE.RAST class
C0799089|T201|COMP|15922-8|LNC|Penicillin V Ab.IgE.RAST class|Penicillin V Ab.IgE.RAST class
C0799090|T201|COMP|15923-6|LNC|Penicillium frequentans Ab.IgE.RAST class|Penicillium frequentans Ab.IgE.RAST class
C0799091|T201|COMP|15924-4|LNC|Penicillium notatum Ab.IgE.RAST class|Penicillium notatum Ab.IgE.RAST class
C0799092|T201|COMP|15925-1|LNC|Piper nigrum Ab.IgE.RAST class|Piper nigrum Ab.IgE.RAST class
C0799093|T201|COMP|15926-9|LNC|Pepper cayenne Ab.IgE.RAST class|Pepper cayenne Ab.IgE.RAST class
C0799094|T201|COMP|15927-7|LNC|Capsicum frutescens Ab.IgE.RAST class|Capsicum frutescens Ab.IgE.RAST class
C0799095|T201|COMP|15928-5|LNC|Pepper green Ab.IgE.RAST class|Pepper green Ab.IgE.RAST class
C0799096|T201|COMP|15929-3|LNC|Schinus molle Ab.IgE.RAST class|Schinus molle Ab.IgE.RAST class
C0799097|T201|COMP|15930-1|LNC|Perca spp Ab.IgE.RAST class|Perca spp Ab.IgE.RAST class
C0799098|T201|COMP|15931-9|LNC|Phoma betae Ab.IgE.RAST class|Phoma betae Ab.IgE.RAST class
C0799099|T201|COMP|15932-7|LNC|Phospholipase Ab.IgE.RAST class|Phospholipase Ab.IgE.RAST class
C0799100|T201|COMP|15933-5|LNC|Phthalic anhydride Ab.IgE.RAST class|Phthalic anhydride Ab.IgE.RAST class
C0799101|T201|COMP|15934-3|LNC|Pigeon droppings Ab.IgE.RAST class|Pigeon droppings Ab.IgE.RAST class
C0799102|T201|COMP|15935-0|LNC|Pigeon feather Ab.IgE.RAST class|Pigeon feather Ab.IgE.RAST class
C0799103|T201|COMP|15936-8|LNC|Pigweed common Ab.IgE.RAST class|Pigweed common Ab.IgE.RAST class
C0799104|T201|COMP|15937-6|LNC|Pigweed rough Ab.IgE.RAST class|Pigweed rough Ab.IgE.RAST class
C0799105|T201|COMP|15938-4|LNC|Pigweed spiny Ab.IgE.RAST class|Pigweed spiny Ab.IgE.RAST class
C0799106|T201|COMP|15939-2|LNC|Pinus nigra Ab.IgE.RAST class|Pinus nigra Ab.IgE.RAST class
C0799107|T201|COMP|15940-0|LNC|Pinus taeda Ab.IgE.RAST class|Pinus taeda Ab.IgE.RAST class
C0799108|T201|COMP|15941-8|LNC|Pinus palustris Ab.IgE.RAST class|Pinus palustris Ab.IgE.RAST class
C0799110|T201|COMP|15943-4|LNC|Pinus edulis Ab.IgE.RAST class|Pinus edulis Ab.IgE.RAST class
C0799111|T201|COMP|15944-2|LNC|Pinus echinata Ab.IgE.RAST class|Pinus echinata Ab.IgE.RAST class
C0799112|T201|COMP|15945-9|LNC|Pinus elliottii Ab.IgE.RAST class|Pinus elliottii Ab.IgE.RAST class
C0799113|T201|COMP|15946-7|LNC|Pinus virginiana Ab.IgE.RAST class|Pinus virginiana Ab.IgE.RAST class
C0799114|T201|COMP|15947-5|LNC|Pinus strobus Ab.IgE.RAST class|Pinus strobus Ab.IgE.RAST class
C0799115|T201|COMP|15948-3|LNC|Ananas comosus Ab.IgE.RAST class|Ananas comosus Ab.IgE.RAST class
C0799116|T201|COMP|15949-1|LNC|Pistacia vera Ab.IgE.RAST class|Pistacia vera Ab.IgE.RAST class
C0799117|T201|COMP|15950-9|LNC|Malassezia furfur Ab.IgE.RAST class|Malassezia furfur Ab.IgE.RAST class
C0799118|T201|COMP|15951-7|LNC|Pleuronectes platessa Ab.IgE.RAST class|Pleuronectes platessa Ab.IgE.RAST class
C0799119|T201|COMP|15952-5|LNC|Plantago lanceolata Ab.IgE.RAST class|Plantago lanceolata Ab.IgE.RAST class
C0799120|T201|COMP|15953-3|LNC|Prunus domestica Ab.IgE.RAST class|Prunus domestica Ab.IgE.RAST class
C0799121|T201|COMP|15954-1|LNC|Populus nigra Ab.IgE.RAST class|Populus nigra Ab.IgE.RAST class
C0799122|T201|COMP|15955-8|LNC|Papaver somniferum Ab.IgE.RAST class|Papaver somniferum Ab.IgE.RAST class
C0799123|T201|COMP|15956-6|LNC|Pork Ab.IgE.RAST class|Pork Ab.IgE.RAST class
C0799125|T201|COMP|15958-2|LNC|Ipomoea batatas Ab.IgE.RAST class|Ipomoea batatas Ab.IgE.RAST class
C0799126|T201|COMP|15959-0|LNC|Iva axillaris Ab.IgE.RAST class|Iva axillaris Ab.IgE.RAST class
C0799127|T201|COMP|15960-8|LNC|Ligustrum vulgare Ab.IgE.RAST class|Ligustrum vulgare Ab.IgE.RAST class
C0799128|T201|COMP|15961-6|LNC|Protamine Ab.IgE.RAST class|Protamine Ab.IgE.RAST class
C0799129|T201|COMP|15962-4|LNC|Prune Ab.IgE.RAST class|Prune Ab.IgE.RAST class
C0799130|T201|COMP|15963-2|LNC|Psyllium seed Ab.IgE.RAST class|Psyllium seed Ab.IgE.RAST class
C0799131|T201|COMP|15964-0|LNC|Aureobasidium pullulans Ab.IgE.RAST class|Aureobasidium pullulans Ab.IgE.RAST class
C0799131|T201|COMP|25329-4|LNC|Aureobasidium pullulans Ab.IgE.RAST class|Aureobasidium pullulans Ab.IgE.RAST class
C0799132|T201|COMP|15965-7|LNC|Pullularia pullulans Ab.IgE.RAST class|Pullularia pullulans Ab.IgE.RAST class
C0799133|T201|COMP|15966-5|LNC|Cucurbita pepo Ab.IgE.RAST class|Cucurbita pepo Ab.IgE.RAST class
C0799134|T201|COMP|15967-3|LNC|Cucurbita pepo seed Ab.IgE.RAST class|Cucurbita pepo seed Ab.IgE.RAST class
C0799135|T201|COMP|15968-1|LNC|Chrysanthemum cinerariifolium Ab.IgE.RAST class|Chrysanthemum cinerariifolium Ab.IgE.RAST class
C0799136|T201|COMP|15969-9|LNC|Rabbit meat Ab.IgE.RAST class|Rabbit meat Ab.IgE.RAST class
C0799137|T201|COMP|15970-7|LNC|Chrysothamnus nauseosus Ab.IgE.RAST class|Chrysothamnus nauseosus Ab.IgE.RAST class
C0799138|T201|COMP|15971-5|LNC|Rabbit epithelium Ab.IgE.RAST class|Rabbit epithelium Ab.IgE.RAST class
C0799139|T201|COMP|15972-3|LNC|Rabbit serum proteins Ab.IgE.RAST class|Rabbit serum proteins Ab.IgE.RAST class
C0799140|T201|COMP|15973-1|LNC|Rabbit urine proteins Ab.IgE.RAST class|Rabbit urine proteins Ab.IgE.RAST class
C0799141|T201|COMP|15974-9|LNC|Raphanus sativus Ab.IgE.RAST class|Raphanus sativus Ab.IgE.RAST class
C0799142|T201|COMP|15975-6|LNC|Ambrosia elatior Ab.IgE.RAST class|Ambrosia elatior Ab.IgE.RAST class
C0799143|T201|COMP|15976-4|LNC|Ambrosia dumosa Ab.IgE.RAST class|Ambrosia dumosa Ab.IgE.RAST class
C0799144|T201|COMP|15977-2|LNC|Franseria acanthicarpa Ab.IgE.RAST class|Franseria acanthicarpa Ab.IgE.RAST class
C0799145|T201|COMP|15978-0|LNC|Ambrosia trifida Ab.IgE.RAST class|Ambrosia trifida Ab.IgE.RAST class
C0799146|T201|COMP|15979-8|LNC|Ambrosia elatior Ab.IgE.RAST class|Ambrosia elatior Ab.IgE.RAST class
C0799147|T201|COMP|15980-6|LNC|Ambrosia bidentata Ab.IgE.RAST class|Ambrosia bidentata Ab.IgE.RAST class
C0799148|T201|COMP|15981-4|LNC|Ambrosia psilostachya Ab.IgE.RAST class|Ambrosia psilostachya Ab.IgE.RAST class
C0799149|T201|COMP|15982-2|LNC|Brassica rapa Ab.IgE.RAST class|Brassica rapa Ab.IgE.RAST class
C0799150|T201|COMP|15983-0|LNC|Rubus idaeus Ab.IgE.RAST class|Rubus idaeus Ab.IgE.RAST class
C0799151|T201|COMP|15984-8|LNC|Rat epithelium Ab.IgE.RAST class|Rat epithelium Ab.IgE.RAST class
C0799152|T201|COMP|15985-5|LNC|Rat serum proteins Ab.IgE.RAST class|Rat serum proteins Ab.IgE.RAST class
C0799153|T201|COMP|15986-3|LNC|Rat urine proteins Ab.IgE.RAST class|Rat urine proteins Ab.IgE.RAST class
C0799154|T201|COMP|15987-1|LNC|Sequoia spp Ab.IgE.RAST class|Sequoia spp Ab.IgE.RAST class
C0799155|T201|COMP|15988-9|LNC|Phalaris arundinacea Ab.IgE.RAST class|Phalaris arundinacea Ab.IgE.RAST class
C0799156|T201|COMP|15989-7|LNC|Phragmites communis Ab.IgE.RAST class|Phragmites communis Ab.IgE.RAST class
C0799157|T201|COMP|15990-5|LNC|Reindeer epithelium Ab.IgE.RAST class|Reindeer epithelium Ab.IgE.RAST class
C0799158|T201|COMP|15991-3|LNC|Rhizopus nigricans Ab.IgE.RAST class|Rhizopus nigricans Ab.IgE.RAST class
C0799159|T201|COMP|15992-1|LNC|Rhodotorula spp Ab.IgE.RAST class|Rhodotorula spp Ab.IgE.RAST class
C0799160|T201|COMP|15993-9|LNC|Rheum spp Ab.IgE.RAST class|Rheum spp Ab.IgE.RAST class
C0799161|T201|COMP|15994-7|LNC|Oryza sativa Ab.IgE.RAST class|Oryza sativa Ab.IgE.RAST class
C0799162|T201|COMP|15995-4|LNC|Zizania spp Ab.IgE.RAST class|Zizania spp Ab.IgE.RAST class
C0799163|T201|COMP|15996-2|LNC|Rosa spp hip Ab.IgE.RAST class|Rosa spp hip Ab.IgE.RAST class
C0799165|T201|COMP|15998-8|LNC|Secale cereale Ab.IgE.RAST class|Secale cereale Ab.IgE.RAST class
C0799166|T201|COMP|15997-0|LNC|Secale cereale pollen Ab.IgE.RAST class|Secale cereale pollen Ab.IgE.RAST class
C0799167|T201|COMP|16000-2|LNC|Lolium perenne Ab.IgE.RAST class|Lolium perenne Ab.IgE.RAST class
C0799167|T201|COMP|15749-5|LNC|Lolium perenne Ab.IgE.RAST class|Lolium perenne Ab.IgE.RAST class
C0799167|T201|COMP|15750-3|LNC|Lolium perenne Ab.IgE.RAST class|Lolium perenne Ab.IgE.RAST class
C0799168|T201|COMP|16001-0|LNC|Carthamus tinctorius Ab.IgE.RAST class|Carthamus tinctorius Ab.IgE.RAST class
C0799169|T201|COMP|16002-8|LNC|Salvia officinalis Ab.IgE.RAST class|Salvia officinalis Ab.IgE.RAST class
C0799171|T201|COMP|16003-6|LNC|Artemisia tridentata Ab.IgE.RAST class|Artemisia tridentata Ab.IgE.RAST class
C0799172|T201|COMP|16005-1|LNC|Saline fish feed Ab.IgE.RAST class|Saline fish feed Ab.IgE.RAST class
C0799173|T201|COMP|16006-9|LNC|Salmo salar Ab.IgE.RAST class|Salmo salar Ab.IgE.RAST class
C0799174|T201|COMP|16007-7|LNC|Saltbush Ab.IgE.RAST class|Saltbush Ab.IgE.RAST class
C0799175|T201|COMP|16008-5|LNC|Sardina pilchardus Ab.IgE.RAST class|Sardina pilchardus Ab.IgE.RAST class
C0799176|T201|COMP|16009-3|LNC|Savinase Ab.IgE.RAST class|Savinase Ab.IgE.RAST class
C0799177|T201|COMP|15812-1|LNC|Atriplex lentiformis Ab.IgE.RAST class|Atriplex lentiformis Ab.IgE.RAST class
C0799178|T201|COMP|16011-9|LNC|Pecten spp Ab.IgE.RAST class|Pecten spp Ab.IgE.RAST class
C0799179|T201|COMP|16012-7|LNC|Cytisus scoparius Ab.IgE.RAST class|Cytisus scoparius Ab.IgE.RAST class
C0799180|T201|COMP|16013-5|LNC|Sericin Ab.IgE.RAST class|Sericin Ab.IgE.RAST class
C0799181|T201|COMP|16014-3|LNC|Sesamum indicum Ab.IgE.RAST class|Sesamum indicum Ab.IgE.RAST class
C0799182|T201|COMP|16015-0|LNC|Sheep epithelium Ab.IgE.RAST class|Sheep epithelium Ab.IgE.RAST class
C0799183|T201|COMP|16016-8|LNC|Rumex acetosella Ab.IgE.RAST class|Rumex acetosella Ab.IgE.RAST class
C0799184|T201|COMP|16017-6|LNC|Sheep wool Ab.IgE.RAST class|Sheep wool Ab.IgE.RAST class
C0799185|T201|COMP|16018-4|LNC|Pandalus borealis Ab.IgE.RAST class|Pandalus borealis Ab.IgE.RAST class
C0799186|T201|COMP|16019-2|LNC|Silk Ab.IgE.RAST class|Silk Ab.IgE.RAST class
C0799187|T201|COMP|16020-0|LNC|Silk waste Ab.IgE.RAST class|Silk waste Ab.IgE.RAST class
C0799188|T201|COMP|16021-8|LNC|Silver Ab.IgE.RAST class|Silver Ab.IgE.RAST class
C0799189|T201|COMP|16022-6|LNC|Ustilago cynodontis Ab.IgE.RAST class|Ustilago cynodontis Ab.IgE.RAST class
C0799190|T201|COMP|16023-4|LNC|Sphacelotheca cruenta Ab.IgE.RAST class|Sphacelotheca cruenta Ab.IgE.RAST class
C0799191|T201|COMP|16024-2|LNC|Helix aspersa Ab.IgE.RAST class|Helix aspersa Ab.IgE.RAST class
C0799192|T201|COMP|16025-9|LNC|Snapper red Ab.IgE.RAST class|Snapper red Ab.IgE.RAST class
C0799193|T201|COMP|16026-7|LNC|Solea solea Ab.IgE.RAST class|Solea solea Ab.IgE.RAST class
C0799194|T201|COMP|16027-5|LNC|Spinacia oleracea Ab.IgE.RAST class|Spinacia oleracea Ab.IgE.RAST class
C0799195|T201|COMP|16028-3|LNC|Spondylocladium citrovirens Ab.IgE.RAST class|Spondylocladium citrovirens Ab.IgE.RAST class
C0799196|T201|COMP|16029-1|LNC|Picea excelsa Ab.IgE.RAST class|Picea excelsa Ab.IgE.RAST class
C0799197|T201|COMP|16030-9|LNC|Squash Ab.IgE.RAST class|Squash Ab.IgE.RAST class
C0799198|T201|COMP|16031-7|LNC|Loligo sp Ab.IgE.RAST class|Loligo sp Ab.IgE.RAST class
C0799199|T201|COMP|16032-5|LNC|Todarodes pacificus Ab.IgE.RAST class|Todarodes pacificus Ab.IgE.RAST class
C0799200|T201|COMP|16033-3|LNC|Stemphylium botryosum Ab.IgE.RAST class|Stemphylium botryosum Ab.IgE.RAST class
C0799201|T201|COMP|16034-1|LNC|Stemphylium solani Ab.IgE.RAST class|Stemphylium solani Ab.IgE.RAST class
C0799202|T201|COMP|16035-8|LNC|Acarus siro Ab.IgE.RAST class|Acarus siro Ab.IgE.RAST class
C0799203|T201|COMP|16037-4|LNC|Tyrophagus putrescentiae Ab.IgE.RAST class|Tyrophagus putrescentiae Ab.IgE.RAST class
C0799204|T201|COMP|16038-2|LNC|Fragaria vesca Ab.IgE.RAST class|Fragaria vesca Ab.IgE.RAST class
C0799205|T201|COMP|16039-0|LNC|Succinylcholine Ab.IgE.RAST class|Succinylcholine Ab.IgE.RAST class
C0799206|T201|COMP|16040-8|LNC|Saccharum officinarum Ab.IgE.RAST class|Saccharum officinarum Ab.IgE.RAST class
C0799207|T201|COMP|16041-6|LNC|Helianthus annuus pollen Ab.IgE.RAST class|Helianthus annuus pollen Ab.IgE.RAST class
C0799208|T201|COMP|16042-4|LNC|Helianthus annuus seed Ab.IgE.RAST class|Helianthus annuus seed Ab.IgE.RAST class
C0799209|T201|COMP|16043-2|LNC|Swine epithelium Ab.IgE.RAST class|Swine epithelium Ab.IgE.RAST class
C0799210|T201|COMP|16044-0|LNC|Swine urine proteins Ab.IgE.RAST class|Swine urine proteins Ab.IgE.RAST class
C0799211|T201|COMP|16045-7|LNC|Xiphias gladius Ab.IgE.RAST class|Xiphias gladius Ab.IgE.RAST class
C0799212|T201|COMP|16046-5|LNC|Platanus occidentalis Ab.IgE.RAST class|Platanus occidentalis Ab.IgE.RAST class
C0799213|T201|COMP|16047-3|LNC|Citrus reticulata Ab.IgE.RAST class|Citrus reticulata Ab.IgE.RAST class
C0799214|T201|COMP|16048-1|LNC|Manihot esculenta crantz Ab.IgE.RAST class|Manihot esculenta crantz Ab.IgE.RAST class
C0799215|T201|COMP|16049-9|LNC|Artemisia dracunculus Ab.IgE.RAST class|Artemisia dracunculus Ab.IgE.RAST class
C0799216|T201|COMP|16050-7|LNC|Camellia sinensis Ab.IgE.RAST class|Camellia sinensis Ab.IgE.RAST class
C0799217|T201|COMP|16051-5|LNC|Tetramin Ab.IgE.RAST class|Tetramin Ab.IgE.RAST class
C0799218|T201|COMP|16052-3|LNC|Salsola kali Ab.IgE.RAST class|Salsola kali Ab.IgE.RAST class
C0799219|T201|COMP|16053-1|LNC|Thymus vulgaris Ab.IgE.RAST class|Thymus vulgaris Ab.IgE.RAST class
C0799220|T201|COMP|16054-9|LNC|Phleum pratense Ab.IgE.RAST class|Phleum pratense Ab.IgE.RAST class
C0799221|T201|COMP|16055-6|LNC|Nicotiana tabacum cigarette Ab.IgE.RAST class|Nicotiana tabacum cigarette Ab.IgE.RAST class
C0799222|T201|COMP|16056-4|LNC|Nicotiana tabacum Ab.IgE.RAST class|Nicotiana tabacum Ab.IgE.RAST class
C0799223|T201|COMP|16057-2|LNC|Lycopersicon lycopersicum Ab.IgE.RAST class|Lycopersicon lycopersicum Ab.IgE.RAST class
C0799224|T201|COMP|16058-0|LNC|Astragalus spp Ab.IgE.RAST class|Astragalus spp Ab.IgE.RAST class
C0799225|T201|COMP|16059-8|LNC|Trichoderma viride Ab.IgE.RAST class|Trichoderma viride Ab.IgE.RAST class
C0799226|T201|COMP|16060-6|LNC|Trichophyton Ab.IgE.RAST class|Trichophyton Ab.IgE.RAST class
C0799227|T201|COMP|16061-4|LNC|Trichophyton rubrum Ab.IgE.RAST class|Trichophyton rubrum Ab.IgE.RAST class
C0799228|T201|COMP|16062-2|LNC|Trichosporon spp Ab.IgE.RAST class|Trichosporon spp Ab.IgE.RAST class
C0799229|T201|COMP|16063-0|LNC|Trimellitic anhydride Ab.IgE.RAST class|Trimellitic anhydride Ab.IgE.RAST class
C0799230|T201|COMP|16064-8|LNC|Oncorhynchus mykiss Ab.IgE.RAST class|Oncorhynchus mykiss Ab.IgE.RAST class
C0799231|T201|COMP|16065-5|LNC|Thunnus albacares Ab.IgE.RAST class|Thunnus albacares Ab.IgE.RAST class
C0799232|T201|COMP|16066-3|LNC|Turkey meat Ab.IgE.RAST class|Turkey meat Ab.IgE.RAST class
C0799233|T201|COMP|16067-1|LNC|Turnip Ab.IgE.RAST class|Turnip Ab.IgE.RAST class
C0799234|T201|COMP|16069-7|LNC|Ulocladium chartarum Ab.IgE.RAST class|Ulocladium chartarum Ab.IgE.RAST class
C0799235|T201|COMP|16070-5|LNC|Ustilago nuda Ab.IgE.RAST class|Ustilago nuda Ab.IgE.RAST class
C0799236|T201|COMP|16071-3|LNC|Vanilla planifolia Ab.IgE.RAST class|Vanilla planifolia Ab.IgE.RAST class
C0799237|T201|COMP|16072-1|LNC|Veal Ab.IgE.RAST class|Veal Ab.IgE.RAST class
C0799238|T201|COMP|16073-9|LNC|Wall pellitory Ab.IgE.RAST class|Wall pellitory Ab.IgE.RAST class
C0799239|T201|COMP|16074-7|LNC|Juglans spp Ab.IgE.RAST class|Juglans spp Ab.IgE.RAST class
C0799240|T201|COMP|16075-4|LNC|Juglans nigra Ab.IgE.RAST class|Juglans nigra Ab.IgE.RAST class
C0799241|T201|COMP|16076-2|LNC|Juglans nigra pollen Ab.IgE.RAST class|Juglans nigra pollen Ab.IgE.RAST class
C0799242|T201|COMP|16077-0|LNC|Juglans regia pollen Ab.IgE.RAST class|Juglans regia pollen Ab.IgE.RAST class
C0799244|T201|COMP|16078-8|LNC|Juglans california pollen Ab.IgE.RAST class|Juglans california pollen Ab.IgE.RAST class
C0799246|T201|COMP|16080-4|LNC|Polistes spp Ab.IgE.RAST class|Polistes spp Ab.IgE.RAST class
C0799247|T201|COMP|16082-0|LNC|Vespula spp Ab.IgE.RAST class|Vespula spp Ab.IgE.RAST class
C0799248|T201|COMP|16083-8|LNC|Citrullus lanatus Ab.IgE.RAST class|Citrullus lanatus Ab.IgE.RAST class
C0799249|T201|COMP|16084-6|LNC|Sitophilus granarius Ab.IgE.RAST class|Sitophilus granarius Ab.IgE.RAST class
C0799250|T201|COMP|16085-3|LNC|Triticum aestivum Ab.IgE.RAST class|Triticum aestivum Ab.IgE.RAST class
C0799251|T201|COMP|16086-1|LNC|Triticum aestivum pollen Ab.IgE.RAST class|Triticum aestivum pollen Ab.IgE.RAST class
C0799252|T201|COMP|16087-9|LNC|Triticum aestivum pollen Ab.IgE.RAST class|Triticum aestivum pollen Ab.IgE.RAST class
C0799253|T201|COMP|16088-7|LNC|Puccinia graminis triticu Ab.IgE.RAST class|Puccinia graminis triticu Ab.IgE.RAST class
C0799254|T201|COMP|16089-5|LNC|Cow whey Ab.IgE.RAST class|Cow whey Ab.IgE.RAST class
C0799255|T201|COMP|16090-3|LNC|Whitefish Ab.IgE.RAST class|Whitefish Ab.IgE.RAST class
C0799256|T201|COMP|16091-1|LNC|Salix caprea Ab.IgE.RAST class|Salix caprea Ab.IgE.RAST class
C0799257|T201|COMP|16092-9|LNC|Salix nigra Ab.IgE.RAST class|Salix nigra Ab.IgE.RAST class
C0799258|T201|COMP|16093-7|LNC|Salix discolor Ab.IgE.RAST class|Salix discolor Ab.IgE.RAST class
C0799259|T201|COMP|16094-5|LNC|Atriplex canescens Ab.IgE.RAST class|Atriplex canescens Ab.IgE.RAST class
C0799260|T201|COMP|16095-2|LNC|Artemisia absinthium Ab.IgE.RAST class|Artemisia absinthium Ab.IgE.RAST class
C0799261|T201|COMP|16096-0|LNC|Saccharomyces cerevisiae Ab.IgE.RAST class|Saccharomyces cerevisiae Ab.IgE.RAST class
C0799262|T201|COMP|16097-8|LNC|Yeast bakers Ab.IgE.RAST class|Yeast bakers Ab.IgE.RAST class
C0799263|T201|COMP|16098-6|LNC|Yeast brewer's Ab.IgE.RAST class|Yeast brewer's Ab.IgE.RAST class
C0799264|T201|COMP|16099-4|LNC|Ethionamide|Ethionamide
C0799266|T201|COMP|16101-8|LNC|Cuminum cyminum Ab.IgE|Cuminum cyminum Ab.IgE
C0799267|T201|COMP|16102-6|LNC|Gelatin bovine Ab.IgE|Gelatin bovine Ab.IgE
C0799268|T201|COMP|16103-4|LNC|Gelatin porcine Ab.IgE|Gelatin porcine Ab.IgE
C0799269|T201|COMP|16104-2|LNC|Broussonetia papyrifera Ab.IgE|Broussonetia papyrifera Ab.IgE
C0799270|T201|COMP|16105-9|LNC|Pheasant Ab.IgE|Pheasant Ab.IgE
C0799271|T201|COMP|16106-7|LNC|Cells.CD8+CD28+|Cells.CD8+CD28+
C0799272|T201|COMP|16107-5|LNC|Cells.CD8+HLA-DR+|Cells.CD8+HLA-DR+
C0799274|T201|COMP|16109-1|LNC|Prolactin^2H post XXX challenge|Prolactin^2H post XXX challenge
C0799275|T201|COMP|16110-9|LNC|11-Deoxycorticosterone|11-Deoxycorticosterone
C0799276|T201|COMP|16111-7|LNC|Epinephrine+Norepinephrine|Epinephrine+Norepinephrine
C0799277|T201|COMP|16112-5|LNC|Estrogen receptor|Estrogen receptor
C0799278|T201|COMP|16113-3|LNC|Progesterone receptor|Progesterone receptor
C0799279|T201|COMP|16114-1|LNC|Amitriptyline|Amitriptyline
C0799280|T201|COMP|16115-8|LNC|Doxepin|Doxepin
C0799281|T201|COMP|16116-6|LNC|Tetrahydrocortisone|Tetrahydrocortisone
C0799282|T201|COMP|16117-4|LNC|Babesia microti Ab.IgG|Babesia microti Ab.IgG
C0799283|T201|COMP|16118-2|LNC|Babesia microti Ab.IgM|Babesia microti Ab.IgM
C0799284|T201|COMP|16119-0|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C0799285|T201|COMP|16120-8|LNC|Brucella abortus Ab.IgM|Brucella abortus Ab.IgM
C0799286|T201|COMP|16121-6|LNC|Colorado tick fever virus Ab.IgG|Colorado tick fever virus Ab.IgG
C0799287|T201|COMP|16122-4|LNC|Colorado tick fever virus Ab.IgM|Colorado tick fever virus Ab.IgM
C0799288|T201|COMP|16123-2|LNC|Cryptococcus sp Ab|Cryptococcus sp Ab
C0799289|T201|COMP|16124-0|LNC|Cryptococcus sp Ab|Cryptococcus sp Ab
C0799290|T201|COMP|16125-7|LNC|Helicobacter pylori Ab.IgA|Helicobacter pylori Ab.IgA
C0799291|T201|COMP|16126-5|LNC|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C0799292|T201|COMP|16127-3|LNC|Helicobacter pylori Ab.IgM|Helicobacter pylori Ab.IgM
C0799293|T201|COMP|16128-1|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C0799294|T201|COMP|16129-9|LNC|Hepatitis C virus Ab.IgG|Hepatitis C virus Ab.IgG
C0799295|T201|COMP|16130-7|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C0799296|T201|COMP|16131-5|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C0799297|T201|COMP|16132-3|LNC|HIV 1 p15+p18 Ab|HIV 1 p15+p18 Ab
C0799298|T201|COMP|16133-1|LNC|Legionella pneumophila Ab.IgM|Legionella pneumophila Ab.IgM
C0799299|T201|COMP|16134-9|LNC|Neisseria meningitidis|Neisseria meningitidis
C0799300|T201|COMP|16135-6|LNC|Beta 2 glycoprotein 1 Ab.IgG|Beta 2 glycoprotein 1 Ab.IgG
C0799301|T201|COMP|16136-4|LNC|Beta 2 glycoprotein 1 Ab.IgM|Beta 2 glycoprotein 1 Ab.IgM
C0799302|T201|COMP|16137-2|LNC|Centromere Ab|Centromere Ab
C0799303|T201|COMP|16138-0|LNC|Ganglioside GM1 Ab.IgA|Ganglioside GM1 Ab.IgA
C0799304|T201|COMP|16139-8|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C0799305|T201|COMP|16140-6|LNC|Tellurium|Tellurium
C0799306|T201|COMP|16141-4|LNC|Nitrogen|Nitrogen
C0799309|T201|COMP|16144-8|LNC|Droperidol|Droperidol
C0799310|T201|COMP|16145-5|LNC|Mescaline|Mescaline
C0799311|T201|COMP|16146-3|LNC|Psilocin|Psilocin
C0799312|T201|COMP|16147-1|LNC|Aldosterone^3rd specimen post XXX challenge|Aldosterone^3rd specimen post XXX challenge
C0799313|T201|COMP|16148-9|LNC|Aldosterone^4th specimen post XXX challenge|Aldosterone^4th specimen post XXX challenge
C0799314|T201|COMP|16149-7|LNC|Aldosterone^5th specimen post XXX challenge|Aldosterone^5th specimen post XXX challenge
C0799315|T201|COMP|16150-5|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0799316|T201|COMP|16151-3|LNC|Dechlorane|Dechlorane
C0799317|T201|COMP|16152-1|LNC|Gastrin^2nd specimen post XXX challenge|Gastrin^2nd specimen post XXX challenge
C0799318|T201|COMP|16153-9|LNC|Gastrin^3rd specimen post XXX challenge|Gastrin^3rd specimen post XXX challenge
C0799319|T201|COMP|16154-7|LNC|Gastrin^4th specimen post XXX challenge|Gastrin^4th specimen post XXX challenge
C0799320|T201|COMP|16155-4|LNC|Gastrin^5th specimen post XXX challenge|Gastrin^5th specimen post XXX challenge
C0799321|T201|COMP|16156-2|LNC|Gastrin^6th specimen post XXX challenge|Gastrin^6th specimen post XXX challenge
C0799322|T201|COMP|16157-0|LNC|Gastrin^7th specimen post XXX challenge|Gastrin^7th specimen post XXX challenge
C0799323|T201|COMP|16158-8|LNC|Gastrin^8th specimen post XXX challenge|Gastrin^8th specimen post XXX challenge
C0799324|T201|COMP|16159-6|LNC|Gastrin^9th specimen post XXX challenge|Gastrin^9th specimen post XXX challenge
C0799325|T201|COMP|16160-4|LNC|Gastrin^10th specimen post XXX challenge|Gastrin^10th specimen post XXX challenge
C0799326|T201|COMP|16161-2|LNC|Gastrin^post XXX challenge|Gastrin^post XXX challenge
C0799327|T201|COMP|16162-0|LNC|Parathyrin.intact^30M post XXX challenge|Parathyrin.intact^30M post XXX challenge
C0799328|T201|COMP|16163-8|LNC|Parathyrin.intact^1H post XXX challenge|Parathyrin.intact^1H post XXX challenge
C0799329|T201|COMP|16164-6|LNC|Parathyrin.intact^2H post XXX challenge|Parathyrin.intact^2H post XXX challenge
C0799330|T201|COMP|16165-3|LNC|Glucose^10 AM specimen|Glucose^10 AM specimen
C0799331|T201|COMP|16166-1|LNC|Glucose^11 AM specimen|Glucose^11 AM specimen
C0799332|T201|COMP|16167-9|LNC|Glucose^2 PM specimen|Glucose^2 PM specimen
C0799333|T201|COMP|16168-7|LNC|Glucose^3 PM specimen|Glucose^3 PM specimen
C0799334|T201|COMP|16169-5|LNC|Glucose^4 PM specimen|Glucose^4 PM specimen
C0799335|T201|COMP|16170-3|LNC|Glucose^5 PM specimen|Glucose^5 PM specimen
C0799336|T201|COMP|16171-1|LNC|Cocaethylene|Cocaethylene
C0799337|T201|COMP|16172-9|LNC|Magnesium|Magnesium
C0799338|T201|COMP|16173-7|LNC|Amyl ether|Amyl ether
C0799339|T201|COMP|16174-5|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C0799340|T201|COMP|16175-2|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C0799341|T201|COMP|16176-0|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C0799342|T201|COMP|16177-8|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C0799343|T201|COMP|16178-6|LNC|Beryllium|Beryllium
C0799344|T201|COMP|16179-4|LNC|Polychlorinated biphenyl|Polychlorinated biphenyl
C0799345|T201|COMP|16180-2|LNC|Zinc|Zinc
C0799346|T201|COMP|16181-0|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0799347|T201|COMP|16182-8|LNC|Alkaline phosphatase isoenzymes|Alkaline phosphatase isoenzymes
C0799348|T201|COMP|16183-6|LNC|Phenolphthalein|Phenolphthalein
C0799349|T201|COMP|16184-4|LNC|Temazepam|Temazepam
C0799350|T201|COMP|16185-1|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0799351|T201|COMP|16186-9|LNC|Hydroxyalprazolam|Hydroxyalprazolam
C0799352|T201|COMP|16187-7|LNC|ALPRAZolam|ALPRAZolam
C0799353|T201|COMP|16188-5|LNC|Creatinine^2H specimen|Creatinine^2H specimen
C0799354|T201|COMP|16189-3|LNC|Creatinine^4H specimen|Creatinine^4H specimen
C0799355|T201|COMP|16190-1|LNC|Amobarbital|Amobarbital
C0799356|T201|COMP|16191-9|LNC|Butabarbital|Butabarbital
C0799357|T201|COMP|16192-7|LNC|PHENobarbital|PHENobarbital
C0799358|T201|COMP|16193-5|LNC|PENTobarbital|PENTobarbital
C0799359|T201|COMP|16194-3|LNC|Secobarbital|Secobarbital
C0799360|T201|COMP|16195-0|LNC|Benzodiazepines|Benzodiazepines
C0799361|T201|COMP|16196-8|LNC|Morphine|Morphine
C0799362|T201|COMP|16197-6|LNC|Codeine|Codeine
C0799363|T201|COMP|16198-4|LNC|Diamorphine|Diamorphine
C0799364|T201|COMP|16199-2|LNC|Methadone|Methadone
C0799365|T201|COMP|16200-8|LNC|Propoxyphene|Propoxyphene
C0799366|T201|COMP|16201-6|LNC|Oxazepam|Oxazepam
C0799367|T201|COMP|16202-4|LNC|Nordiazepam|Nordiazepam
C0799368|T201|COMP|16203-2|LNC|ALPRAZolam|ALPRAZolam
C0799369|T201|COMP|16204-0|LNC|clonazePAM|clonazePAM
C0799370|T201|COMP|16205-7|LNC|LORazepam|LORazepam
C0799371|T201|COMP|16206-5|LNC|Temazepam|Temazepam
C0799372|T201|COMP|16207-3|LNC|Meperidine|Meperidine
C0799373|T201|COMP|16208-1|LNC|Buprenorphine|Buprenorphine
C0799374|T201|COMP|16209-9|LNC|Chlorpheniramine|Chlorpheniramine
C0799375|T201|COMP|16210-7|LNC|Diethylpropion|Diethylpropion
C0799376|T201|COMP|16211-5|LNC|Dihydrocodeine|Dihydrocodeine
C0799377|T201|COMP|16212-3|LNC|Ethylamphetamine|Ethylamphetamine
C0799378|T201|COMP|16213-1|LNC|Levorphanol|Levorphanol
C0799379|T201|COMP|16214-9|LNC|Lysergate diethylamide|Lysergate diethylamide
C0799380|T201|COMP|16215-6|LNC|Mephobarbital|Mephobarbital
C0799381|T201|COMP|16216-4|LNC|MethylePHEDrine|MethylePHEDrine
C0799382|T201|COMP|16217-2|LNC|Methyprylon|Methyprylon
C0799383|T201|COMP|16218-0|LNC|Nalbuphine|Nalbuphine
C0799384|T201|COMP|16219-8|LNC|Pentazocine|Pentazocine
C0799385|T201|COMP|16220-6|LNC|Phenmetrazine|Phenmetrazine
C0799386|T201|COMP|16221-4|LNC|Phenothiazines|Phenothiazines
C0799387|T201|COMP|16222-2|LNC|Phentermine|Phentermine
C0799388|T201|COMP|16223-0|LNC|Thiopental|Thiopental
C0799389|T201|COMP|16224-8|LNC|Triazolam|Triazolam
C0799390|T201|COMP|16225-5|LNC|Amitriptyline|Amitriptyline
C0799391|T201|COMP|16226-3|LNC|Benzoylecgonine|Benzoylecgonine
C0799392|T201|COMP|16227-1|LNC|diazePAM|diazePAM
C0799393|T201|COMP|16228-9|LNC|Nordiazepam|Nordiazepam
C0799394|T201|COMP|16229-7|LNC|clonazePAM|clonazePAM
C0799395|T201|COMP|16230-5|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0799396|T201|COMP|16231-3|LNC|Flurazepam|Flurazepam
C0799397|T201|COMP|16232-1|LNC|Triazolam|Triazolam
C0799398|T201|COMP|16233-9|LNC|Midazolam|Midazolam
C0799399|T201|COMP|16234-7|LNC|Amphetamine|Amphetamine
C0799400|T201|COMP|16235-4|LNC|Methamphetamine|Methamphetamine
C0799401|T201|COMP|16236-2|LNC|Butabarbital|Butabarbital
C0799402|T201|COMP|16237-0|LNC|Butalbital|Butalbital
C0799403|T201|COMP|16238-8|LNC|Secobarbital|Secobarbital
C0799404|T201|COMP|16239-6|LNC|Amobarbital|Amobarbital
C0799405|T201|COMP|16240-4|LNC|PENTobarbital|PENTobarbital
C0799406|T201|COMP|16241-2|LNC|PHENobarbital|PHENobarbital
C0799407|T201|COMP|16242-0|LNC|Propoxyphene|Propoxyphene
C0799408|T201|COMP|16243-8|LNC|Cannabinoids|Cannabinoids
C0799409|T201|COMP|16244-6|LNC|Methaqualone|Methaqualone
C0799410|T201|COMP|16245-3|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C0799411|T201|COMP|16246-1|LNC|Methadone|Methadone
C0799412|T201|COMP|16247-9|LNC|Dextromethorphan|Dextromethorphan
C0799413|T201|COMP|16248-7|LNC|6-Monoacetylmorphine.free|6-Monoacetylmorphine.free
C0799414|T201|COMP|16249-5|LNC|oxyCODONE|oxyCODONE
C0799415|T201|COMP|16250-3|LNC|Codeine|Codeine
C0799416|T201|COMP|16251-1|LNC|Morphine|Morphine
C0799417|T201|COMP|16252-9|LNC|HYDROcodone|HYDROcodone
C0799418|T201|COMP|16253-7|LNC|Meperidine|Meperidine
C0799419|T201|COMP|16254-5|LNC|Phencyclidine|Phencyclidine
C0799420|T201|COMP|16255-2|LNC|Troponin I.cardiac|Troponin I.cardiac
C0799421|T201|COMP|16257-8|LNC|Sodium urate crystals|Sodium urate crystals
C0799422|T201|COMP|16258-6|LNC|Ammonium urate crystals|Ammonium urate crystals
C0799423|T201|COMP|16259-4|LNC|Urate dihydrate crystals|Urate dihydrate crystals
C0799424|T201|COMP|16260-2|LNC|Triamterene crystals|Triamterene crystals
C0799425|T201|COMP|16261-0|LNC|Calcium bilirubinate crystals|Calcium bilirubinate crystals
C0799426|T201|COMP|16262-8|LNC|Newberyite crystals|Newberyite crystals
C0799427|T201|COMP|16263-6|LNC|Calcium oxalate dihydrate crystals|Calcium oxalate dihydrate crystals
C0799428|T201|COMP|16264-4|LNC|Calcium oxalate monohydrate crystals|Calcium oxalate monohydrate crystals
C0799429|T201|COMP|16265-1|LNC|Triple phosphate crystals|Triple phosphate crystals
C0799430|T201|COMP|16266-9|LNC|Calcium hydrogen phosphate crystals|Calcium hydrogen phosphate crystals
C0799431|T201|COMP|16267-7|LNC|Calcium carbonate crystals|Calcium carbonate crystals
C0799432|T201|COMP|16268-5|LNC|Calcium phosphate crystals|Calcium phosphate crystals
C0799433|T201|COMP|16269-3|LNC|Urate crystals|Urate crystals
C0799434|T201|COMP|16270-1|LNC|Calcium^1H post XXX challenge|Calcium^1H post XXX challenge
C0799435|T201|COMP|16271-9|LNC|Calcium^30M post XXX challenge|Calcium^30M post XXX challenge
C0799436|T201|COMP|16272-7|LNC|Calcium^2H post XXX challenge|Calcium^2H post XXX challenge
C0799437|T201|COMP|16273-5|LNC|Calcium|Calcium
C0799438|T201|COMP|16274-3|LNC|Cells.CD4/Cells.C4|Cells.CD4/Cells.C4
C0799439|T201|COMP|16275-0|LNC|Bartonella sp DNA|Bartonella sp DNA
C0799440|T201|COMP|16276-8|LNC|Bartonella henselae DNA|Bartonella henselae DNA
C0799441|T201|COMP|16277-6|LNC|Bartonella quintana DNA|Bartonella quintana DNA
C0799442|T201|COMP|16278-4|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C0799443|T201|COMP|16279-2|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C0799444|T201|COMP|16280-0|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C0799445|T201|COMP|16281-8|LNC|traZODone|traZODone
C0799446|T201|COMP|16282-6|LNC|Acetaminophen|Acetaminophen
C0799447|T201|COMP|16283-4|LNC|Escherichia coli verotoxin|Escherichia coli verotoxin
C0799448|T201|COMP|16284-2|LNC|Polio virus Ab|Polio virus Ab
C0799449|T201|COMP|16285-9|LNC|Creatinine/Protein|Creatinine/Protein
C0799450|T201|COMP|16286-7|LNC|Testosterone.free/Testosterone.total|Testosterone.free/Testosterone.total
C0799451|T201|COMP|16287-5|LNC|Sulfatide Ab|Sulfatide Ab
C0799452|T201|COMP|16288-3|LNC|Monosialoganglioside GM1 Ab.IgG+IgM|Monosialoganglioside GM1 Ab.IgG+IgM
C0799453|T201|COMP|16289-1|LNC|Monosialoganglioside GM1 Ab|Monosialoganglioside GM1 Ab
C0799454|T201|COMP|16290-9|LNC|Neutrophils|Neutrophils
C0799455|T201|COMP|16291-7|LNC|Herpes simplex virus 1|Herpes simplex virus 1
C0799456|T201|COMP|16292-5|LNC|1,4-Dioxane|1,4-Dioxane
C0799457|T201|COMP|16293-3|LNC|11-Deoxycorticosteroids|11-Deoxycorticosteroids
C0799458|T201|COMP|16294-1|LNC|11-Deoxycorticosterone^post XXX challenge|11-Deoxycorticosterone^post XXX challenge
C0799459|T201|COMP|16295-8|LNC|11-Deoxycortisol^post XXX challenge|11-Deoxycortisol^post XXX challenge
C0799460|T201|COMP|16296-6|LNC|11-Hydroxyandrosterone|11-Hydroxyandrosterone
C0799461|T201|COMP|16297-4|LNC|17-Hydroxypregnenolone|17-Hydroxypregnenolone
C0799462|T201|COMP|16298-2|LNC|17-Hydroxypregnenolone^45M post XXX challenge|17-Hydroxypregnenolone^45M post XXX challenge
C0799463|T201|COMP|16299-0|LNC|17-Hydroxypregnenolone^6H post XXX challenge|17-Hydroxypregnenolone^6H post XXX challenge
C0799464|T201|COMP|16300-6|LNC|17-Ketogenic steroids|17-Ketogenic steroids
C0799465|T201|COMP|16301-4|LNC|17-Ketogenic steroids^baseline|17-Ketogenic steroids^baseline
C0799466|T201|COMP|16302-2|LNC|1-Methylhistidine|1-Methylhistidine
C0799467|T201|COMP|16303-0|LNC|2-Hexanol|2-Hexanol
C0799468|T201|COMP|16304-8|LNC|2-Hexanol/Creatinine|2-Hexanol/Creatinine
C0799469|T201|COMP|16305-5|LNC|2-Methoxyethanol|2-Methoxyethanol
C0799470|T201|COMP|16306-3|LNC|3-Methylhistidine|3-Methylhistidine
C0799471|T201|COMP|16307-1|LNC|Acetate|Acetate
C0799472|T201|COMP|16308-9|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C0799473|T201|COMP|16309-7|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C0799474|T201|COMP|16310-5|LNC|Acetone|Acetone
C0799475|T201|COMP|16311-3|LNC|Acetone|Acetone
C0799476|T201|COMP|16312-1|LNC|Acetonitrile|Acetonitrile
C0799477|T201|COMP|16313-9|LNC|Acetylene|Acetylene
C0799478|T201|COMP|16314-7|LNC|Acetylsalicylate|Acetylsalicylate
C0799479|T201|COMP|16315-4|LNC|Acid phosphatase|Acid phosphatase
C0799480|T201|COMP|16316-2|LNC|Acid phosphatase.tartrate resistant|Acid phosphatase.tartrate resistant
C0799481|T201|COMP|16317-0|LNC|Acid phosphatase.prostatic|Acid phosphatase.prostatic
C0799482|T201|COMP|16318-8|LNC|Acrylamide|Acrylamide
C0799483|T201|COMP|16319-6|LNC|Acrylamide|Acrylamide
C0799484|T201|COMP|16320-4|LNC|Acyclovir|Acyclovir
C0799486|T201|COMP|16322-0|LNC|Biperiden|Biperiden
C0799487|T201|COMP|16323-8|LNC|Alanine|Alanine
C0799488|T201|COMP|16324-6|LNC|Alanine aminotransferase|Alanine aminotransferase
C0799490|T201|COMP|16327-9|LNC|Allyl alcohol|Allyl alcohol
C0799491|T201|COMP|16328-7|LNC|Benzyl alcohol|Benzyl alcohol
C0799492|T201|COMP|16329-5|LNC|Aldosterone^6th specimen post XXX challenge|Aldosterone^6th specimen post XXX challenge
C0799493|T201|COMP|16330-3|LNC|Aldosterone^7th specimen post XXX challenge|Aldosterone^7th specimen post XXX challenge
C0799494|T201|COMP|16331-1|LNC|Aldosterone^8th specimen post XXX challenge|Aldosterone^8th specimen post XXX challenge
C0799495|T201|COMP|16332-9|LNC|Aldosterone^9th specimen post XXX challenge|Aldosterone^9th specimen post XXX challenge
C0799496|T201|COMP|16333-7|LNC|Aldrin|Aldrin
C0799497|T201|COMP|16334-5|LNC|Alfentanil|Alfentanil
C0799498|T201|COMP|16335-2|LNC|Hydrocarbons.aliphatic|Hydrocarbons.aliphatic
C0799500|T201|COMP|16337-8|LNC|Alkaline phosphatase|Alkaline phosphatase
C0799501|T201|COMP|16338-6|LNC|Alpha aminoadipate|Alpha aminoadipate
C0799502|T201|COMP|16339-4|LNC|Alpha aminoisobutyrate|Alpha aminoisobutyrate
C0799503|T201|COMP|16340-2|LNC|Alpha aminoisobutyrate|Alpha aminoisobutyrate
C0799504|T201|COMP|16341-0|LNC|Alpha aminoisobutyrate|Alpha aminoisobutyrate
C0799505|T201|COMP|16342-8|LNC|Alpha aminoisobutyrate|Alpha aminoisobutyrate
C0799506|T201|COMP|16343-6|LNC|Alpha aminoisobutyrate|Alpha aminoisobutyrate
C0799507|T201|COMP|16344-4|LNC|Alpha aminoisobutyrate|Alpha aminoisobutyrate
C0799508|T201|COMP|16345-1|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0799509|T201|COMP|16346-9|LNC|Alpha chlordane|Alpha chlordane
C0799510|T201|COMP|16347-7|LNC|Alpha chlordane|Alpha chlordane
C0799511|T201|COMP|16348-5|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C0799512|T201|COMP|16349-3|LNC|Aluminum|Aluminum
C0799513|T201|COMP|16350-1|LNC|Amantadine|Amantadine
C0799514|T201|COMP|16351-9|LNC|aMILoride|aMILoride
C0799515|T201|COMP|16352-7|LNC|aMILoride|aMILoride
C0799516|T201|COMP|16353-5|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0799517|T201|COMP|12471-9|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0799518|T201|COMP|16355-0|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0799519|T201|COMP|13364-5|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0799520|T201|COMP|13365-2|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0799521|T201|COMP|13382-7|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0799522|T201|COMP|16359-2|LNC|Amiodarone+Desethylamiodarone|Amiodarone+Desethylamiodarone
C0799523|T201|COMP|16360-0|LNC|Amitriptyline^peak|Amitriptyline^peak
C0799524|T201|COMP|16361-8|LNC|Amitriptyline^trough|Amitriptyline^trough
C0799525|T201|COMP|16362-6|LNC|Ammonia|Ammonia
C0799526|T201|COMP|16363-4|LNC|Ammonia|Ammonia
C0799527|T201|COMP|16364-2|LNC|Amobarbital|Amobarbital
C0799528|T201|COMP|16365-9|LNC|Amoxicillin+Clavulanate|Amoxicillin+Clavulanate
C0799530|T201|COMP|16367-5|LNC|Amphetamine/Methamphetamine|Amphetamine/Methamphetamine
C0799531|T201|COMP|16369-1|LNC|Amphetamines|Amphetamines
C0799532|T201|COMP|16370-9|LNC|Amphotericin B|Amphotericin B
C0799533|T201|COMP|16373-3|LNC|Amyl ether|Amyl ether
C0799534|T201|COMP|16374-1|LNC|Amyl nitrite|Amyl nitrite
C0799535|T201|COMP|16378-2|LNC|Androstenedione^2nd specimen post XXX challenge|Androstenedione^2nd specimen post XXX challenge
C0799536|T201|COMP|16379-0|LNC|Androstenedione^3rd specimen post XXX challenge|Androstenedione^3rd specimen post XXX challenge
C0799537|T201|COMP|16380-8|LNC|Androstenedione^4th specimen post XXX challenge|Androstenedione^4th specimen post XXX challenge
C0799538|T201|COMP|16381-6|LNC|Androstenedione^5th specimen post XXX challenge|Androstenedione^5th specimen post XXX challenge
C0799539|T201|COMP|16382-4|LNC|Androstenedione^6th specimen post XXX challenge|Androstenedione^6th specimen post XXX challenge
C0799540|T201|COMP|16383-2|LNC|Androstenedione^7th specimen post XXX challenge|Androstenedione^7th specimen post XXX challenge
C0799541|T201|COMP|16384-0|LNC|Androstenedione^8th specimen post XXX challenge|Androstenedione^8th specimen post XXX challenge
C0799542|T201|COMP|16385-7|LNC|Androstenedione^9th specimen post XXX challenge|Androstenedione^9th specimen post XXX challenge
C0799543|T201|COMP|16100-0|LNC|Rifabutin|Rifabutin
C0799544|T201|COMP|16387-3|LNC|Rifabutin+Ethambutol|Rifabutin+Ethambutol
C0799545|T201|COMP|16388-1|LNC|Anticonvulsants|Anticonvulsants
C0799546|T201|COMP|16389-9|LNC|Antidepressants|Antidepressants
C0799547|T201|COMP|16390-7|LNC|Antidiuretics|Antidiuretics
C0799548|T201|COMP|16391-5|LNC|Antimony|Antimony
C0799549|T201|COMP|16392-3|LNC|Nuclear Ab|Nuclear Ab
C0799550|T201|COMP|16393-1|LNC|Nuclear Ab|Nuclear Ab
C0799551|T201|COMP|16394-9|LNC|Nuclear Ab|Nuclear Ab
C0799552|T201|COMP|16395-6|LNC|Antipsychotics|Antipsychotics
C0799553|T201|COMP|16400-4|LNC|Appearance|Appearance
C0799554|T201|COMP|16401-2|LNC|Arginine|Arginine
C0799555|T201|COMP|16402-0|LNC|Aromatic solvents|Aromatic solvents
C0799556|T201|COMP|16403-8|LNC|Arsenic|Arsenic
C0799557|T201|COMP|16404-6|LNC|Arsenic|Arsenic
C0799558|T201|COMP|16405-3|LNC|Arylamidase|Arylamidase
C0799559|T201|COMP|16406-1|LNC|Arylamidase|Arylamidase
C0799560|T201|COMP|16407-9|LNC|Asbestos identified|Asbestos identified
C0799561|T201|COMP|16408-7|LNC|Ascorbate|Ascorbate
C0799562|T201|COMP|16409-5|LNC|Ascorbate^post dose|Ascorbate^post dose
C0799563|T201|COMP|16410-3|LNC|Asparagine|Asparagine
C0799564|T201|COMP|16411-1|LNC|Aspartate|Aspartate
C0799565|T201|COMP|16412-9|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0799566|T201|COMP|16414-5|LNC|Aspergillus amstelodami Ab|Aspergillus amstelodami Ab
C0799567|T201|COMP|16415-2|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C0799568|T201|COMP|16416-0|LNC|Aspergillus terreus Ab|Aspergillus terreus Ab
C0799569|T201|COMP|16417-8|LNC|Aspergillus versicolor Ab|Aspergillus versicolor Ab
C0799570|T201|COMP|16418-6|LNC|Azatadine|Azatadine
C0799571|T201|COMP|16419-4|LNC|azaTHIOprine|azaTHIOprine
C0799572|T201|COMP|16420-2|LNC|Azithromycin|Azithromycin
C0799573|T201|COMP|16421-0|LNC|Azithromycin+Ethambutol|Azithromycin+Ethambutol
C0799574|T201|COMP|16422-8|LNC|Azlocillin|Azlocillin
C0799575|T201|COMP|16423-6|LNC|Aztreonam|Aztreonam
C0799576|T201|COMP|16424-4|LNC|Salicylazosulfapyridine|Salicylazosulfapyridine
C0799577|T201|COMP|16425-1|LNC|Babesia sp Ab.IgM|Babesia sp Ab.IgM
C0799578|T201|COMP|16426-9|LNC|Babesia sp Ab.IgM|Babesia sp Ab.IgM
C0799579|T201|COMP|16427-7|LNC|Babesia microti Ab|Babesia microti Ab
C0799580|T201|COMP|16428-5|LNC|Bacitracin|Bacitracin
C0799581|T201|COMP|16429-3|LNC|Barbiturates|Barbiturates
C0799582|T201|COMP|16430-1|LNC|Barbiturates|Barbiturates
C0799583|T201|COMP|16431-9|LNC|Barium|Barium
C0799584|T201|COMP|16432-7|LNC|Barium|Barium
C0799585|T201|COMP|16433-5|LNC|Basement membrane Ab|Basement membrane Ab
C0799586|T201|COMP|16434-3|LNC|Basement membrane Ab|Basement membrane Ab
C0799587|T201|COMP|16435-0|LNC|Bean white Ab.IgE|Bean white Ab.IgE
C0799589|T201|COMP|16437-6|LNC|Bendroflumethiazide|Bendroflumethiazide
C0799590|T201|COMP|16438-4|LNC|Benzaldehyde|Benzaldehyde
C0799591|T201|COMP|16439-2|LNC|Benzene|Benzene
C0799592|T201|COMP|16440-0|LNC|Benzene ring Ab.IgE|Benzene ring Ab.IgE
C0799593|T201|COMP|16441-8|LNC|Benzene ring Ab.IgG|Benzene ring Ab.IgG
C0799594|T201|COMP|16442-6|LNC|Benzene ring Ab.IgM|Benzene ring Ab.IgM
C0799595|T201|COMP|16443-4|LNC|Benzonatate|Benzonatate
C0799596|T201|COMP|16444-2|LNC|Benzophenone|Benzophenone
C0799597|T201|COMP|16446-7|LNC|Benzoylecgonine|Benzoylecgonine
C0799598|T201|COMP|16447-5|LNC|Cocaine|Cocaine
C0799599|T201|COMP|16448-3|LNC|Cocaine|Cocaine
C0799600|T201|COMP|16449-1|LNC|Benzthiazide|Benzthiazide
C0799601|T201|COMP|16450-9|LNC|Benzylhydrazine|Benzylhydrazine
C0799602|T201|COMP|16451-7|LNC|Beryllium|Beryllium
C0799603|T201|COMP|16452-5|LNC|Beta alanine|Beta alanine
C0799604|T201|COMP|16453-3|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0799605|T201|COMP|16454-1|LNC|Beta galactosidase|Beta galactosidase
C0799606|T201|COMP|16455-8|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C0799607|T201|COMP|16456-6|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C0799608|T201|COMP|16457-4|LNC|Beta-N-acetylhexosaminidase.A|Beta-N-acetylhexosaminidase.A
C0799609|T201|COMP|16458-2|LNC|Bethanechol|Bethanechol
C0799610|T201|COMP|16459-0|LNC|Bicarbonate|Bicarbonate
C0799611|T201|COMP|16460-8|LNC|Bicarbonate|Bicarbonate
C0799612|T201|COMP|16461-6|LNC|Bicarbonate|Bicarbonate
C0799613|T201|COMP|16462-4|LNC|Bicarbonate|Bicarbonate
C0799614|T201|COMP|16463-2|LNC|Bile acid.dihydroxy|Bile acid.dihydroxy
C0799615|T201|COMP|16464-0|LNC|Bile acid|Bile acid
C0799616|T201|COMP|16465-7|LNC|Bile acid|Bile acid
C0799617|T201|COMP|16466-5|LNC|Bile acid.trihydroxy|Bile acid.trihydroxy
C0799618|T201|COMP|16467-3|LNC|Bismuth|Bismuth
C0799619|T201|COMP|16468-1|LNC|Bismuth|Bismuth
C0799620|T201|COMP|16469-9|LNC|Bismuth/Creatinine|Bismuth/Creatinine
C0799621|T201|COMP|16470-7|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0799622|T201|COMP|16471-5|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0799623|T201|COMP|16472-3|LNC|Blastomyces dermatitidis rRNA|Blastomyces dermatitidis rRNA
C0799624|T201|COMP|16473-1|LNC|Bordetella parapertussis Ab|Bordetella parapertussis Ab
C0799625|T201|COMP|16474-9|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C0799626|T201|COMP|16475-6|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0799627|T201|COMP|16476-4|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0799628|T201|COMP|16477-2|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0799629|T201|COMP|16478-0|LNC|Borrelia burgdorferi Ab.IgA|Borrelia burgdorferi Ab.IgA
C0799630|T201|COMP|16479-8|LNC|Borrelia burgdorferi Ab.IgA|Borrelia burgdorferi Ab.IgA
C0799631|T201|COMP|16480-6|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0799632|T201|COMP|16481-4|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0799633|T201|COMP|16482-2|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0799634|T201|COMP|16483-0|LNC|Borrelia hermsii|Borrelia hermsii
C0799635|T201|COMP|16484-8|LNC|Boysenberry Ab.IgE|Boysenberry Ab.IgE
C0799636|T201|COMP|16485-5|LNC|Bromodiphenhydramine|Bromodiphenhydramine
C0799637|T201|COMP|16486-3|LNC|Brucella abortus Ab.IgA+IgG+IgM|Brucella abortus Ab.IgA+IgG+IgM
C0799638|T201|COMP|16487-1|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C0799639|T201|COMP|16488-9|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C0799640|T201|COMP|16489-7|LNC|Brucella melitensis Ab|Brucella melitensis Ab
C0799641|T201|COMP|16490-5|LNC|Brucella suis Ab|Brucella suis Ab
C0799642|T201|COMP|16491-3|LNC|Brush border Ab|Brush border Ab
C0799643|T201|COMP|16492-1|LNC|Bufotenine|Bufotenine
C0799644|T201|COMP|16493-9|LNC|Bufotenine|Bufotenine
C0799645|T201|COMP|16494-7|LNC|Bumetanide|Bumetanide
C0799646|T201|COMP|16495-4|LNC|Buprenorphine|Buprenorphine
C0799647|T201|COMP|16496-2|LNC|Buprenorphine|Buprenorphine
C0799648|T201|COMP|16497-0|LNC|Butabarbital|Butabarbital
C0799649|T201|COMP|16498-8|LNC|Butalbital|Butalbital
C0799650|T201|COMP|16499-6|LNC|Butorphanol|Butorphanol
C0799651|T201|COMP|16500-1|LNC|Butyrate|Butyrate
C0799652|T201|COMP|16501-9|LNC|C peptide^7th specimen post XXX challenge|C peptide^7th specimen post XXX challenge
C0799653|T201|COMP|16502-7|LNC|C peptide^8th specimen post XXX challenge|C peptide^8th specimen post XXX challenge
C0799654|T201|COMP|16503-5|LNC|C reactive protein|C reactive protein
C0799655|T201|COMP|16504-3|LNC|Calcitonin^1.5M post XXX challenge|Calcitonin^1.5M post XXX challenge
C0799656|T201|COMP|16505-0|LNC|Calcitonin^10M post XXX challenge|Calcitonin^10M post XXX challenge
C0799657|T201|COMP|16506-8|LNC|Calcitonin^3H post XXX challenge|Calcitonin^3H post XXX challenge
C0799658|T201|COMP|16507-6|LNC|Calcitonin^4H post XXX challenge|Calcitonin^4H post XXX challenge
C0799659|T201|COMP|16508-4|LNC|Calcitonin^5M post XXX challenge|Calcitonin^5M post XXX challenge
C0799660|T201|COMP|16509-2|LNC|Calcitonin^7th specimen post XXX challenge|Calcitonin^7th specimen post XXX challenge
C0799661|T201|COMP|16510-0|LNC|Calcitonin^8th specimen post XXX challenge|Calcitonin^8th specimen post XXX challenge
C0799662|T201|COMP|16511-8|LNC|Calcitonin^9th specimen post XXX challenge|Calcitonin^9th specimen post XXX challenge
C0799663|T201|COMP|16512-6|LNC|Calcium.ionized^2nd specimen post XXX challenge|Calcium.ionized^2nd specimen post XXX challenge
C0799664|T201|COMP|16513-4|LNC|Calcium.ionized^3rd specimen post XXX challenge|Calcium.ionized^3rd specimen post XXX challenge
C0799665|T201|COMP|16514-2|LNC|Calcium.ionized^4th specimen post XXX challenge|Calcium.ionized^4th specimen post XXX challenge
C0799666|T201|COMP|16515-9|LNC|Calcium.ionized^5th specimen post XXX challenge|Calcium.ionized^5th specimen post XXX challenge
C0799667|T201|COMP|16516-7|LNC|Calcium.ionized^6th specimen post XXX challenge|Calcium.ionized^6th specimen post XXX challenge
C0799668|T201|COMP|16517-5|LNC|Calcium.ionized^7th specimen post XXX challenge|Calcium.ionized^7th specimen post XXX challenge
C0799669|T201|COMP|16518-3|LNC|Calcium|Calcium
C0799670|T201|COMP|16519-1|LNC|Calcium^10M post XXX challenge|Calcium^10M post XXX challenge
C0799671|T201|COMP|16520-9|LNC|Calcium^2nd specimen post XXX challenge|Calcium^2nd specimen post XXX challenge
C0799672|T201|COMP|16521-7|LNC|Calcium^3rd specimen post XXX challenge|Calcium^3rd specimen post XXX challenge
C0799673|T201|COMP|16522-5|LNC|Calcium^4th specimen post XXX challenge|Calcium^4th specimen post XXX challenge
C0799674|T201|COMP|16523-3|LNC|Calcium^5M post XXX challenge|Calcium^5M post XXX challenge
C0799675|T201|COMP|16524-1|LNC|Calcium^6H post XXX challenge|Calcium^6H post XXX challenge
C0799676|T201|COMP|16525-8|LNC|Calcium/Phosphate|Calcium/Phosphate
C0799677|T201|COMP|16526-6|LNC|Calcium/Protein|Calcium/Protein
C0799678|T201|COMP|16527-4|LNC|Calcium/Sodium|Calcium/Sodium
C0799679|T201|COMP|16528-2|LNC|Campylobacter coli rRNA|Campylobacter coli rRNA
C0799680|T201|COMP|16529-0|LNC|Campylobacter jejuni rRNA|Campylobacter jejuni rRNA
C0799681|T201|COMP|16530-8|LNC|Campylobacter jejuni rRNA|Campylobacter jejuni rRNA
C0799682|T201|COMP|16531-6|LNC|Campylobacter lari rRNA|Campylobacter lari rRNA
C0799683|T201|COMP|16532-4|LNC|Campylobacter lari rRNA|Campylobacter lari rRNA
C0799684|T201|COMP|16533-2|LNC|Helicobacter pylori Ab|Helicobacter pylori Ab
C0799685|T201|COMP|16534-0|LNC|Campylobacter sp rRNA|Campylobacter sp rRNA
C0799686|T201|COMP|16535-7|LNC|Canary droppings Ab.IgE|Canary droppings Ab.IgE
C0799687|T201|COMP|16536-5|LNC|Canary serum proteins Ab|Canary serum proteins Ab
C0799688|T201|COMP|16538-1|LNC|Candida sp Ab.IgA|Candida sp Ab.IgA
C0799689|T201|COMP|16539-9|LNC|Candida sp Ag|Candida sp Ag
C0799691|T201|COMP|16542-3|LNC|Cannabinoids|Cannabinoids
C0799692|T201|COMP|16543-1|LNC|Cannabinoids|Cannabinoids
C0799693|T201|COMP|16544-9|LNC|Canrenone|Canrenone
C0799694|T201|COMP|16545-6|LNC|Capreomycin|Capreomycin
C0799695|T201|COMP|16546-4|LNC|Captopril|Captopril
C0799696|T201|COMP|16547-2|LNC|Carbamate pesticides|Carbamate pesticides
C0799697|T201|COMP|16548-0|LNC|carBAMazepine|carBAMazepine
C0799698|T201|COMP|16549-8|LNC|Carbinoxamine|Carbinoxamine
C0799699|T201|COMP|16550-6|LNC|Carbohydrates|Carbohydrates
C0799700|T201|COMP|16551-4|LNC|Carbon dioxide|Carbon dioxide
C0799701|T201|COMP|16553-0|LNC|Carnitine|Carnitine
C0799702|T201|COMP|16555-5|LNC|Carnitine|Carnitine
C0799703|T201|COMP|16556-3|LNC|Carnitine|Carnitine
C0799704|T201|COMP|16557-1|LNC|Carnosine|Carnosine
C0799705|T201|COMP|16558-9|LNC|Catecholamines^2H post XXX challenge|Catecholamines^2H post XXX challenge
C0799706|T201|COMP|16559-7|LNC|Catecholamines^3H post XXX challenge|Catecholamines^3H post XXX challenge
C0799707|T201|COMP|16560-5|LNC|Catecholamines^5th specimen post XXX challenge|Catecholamines^5th specimen post XXX challenge
C0799708|T201|COMP|16561-3|LNC|Catecholamines^6th specimen post XXX challenge|Catecholamines^6th specimen post XXX challenge
C0799709|T201|COMP|16562-1|LNC|Cathartic laxatives|Cathartic laxatives
C0799710|T201|COMP|16563-9|LNC|Cathepsin D|Cathepsin D
C0799711|T201|COMP|16564-7|LNC|Cefaclor|Cefaclor
C0799712|T201|COMP|16565-4|LNC|Cefadroxil|Cefadroxil
C0799713|T201|COMP|16566-2|LNC|ceFAZolin|ceFAZolin
C0799714|T201|COMP|16567-0|LNC|Cefixime|Cefixime
C0799715|T201|COMP|16568-8|LNC|Cefuroxime Ab.IgE|Cefuroxime Ab.IgE
C0799716|T201|COMP|16569-6|LNC|cefTRIAXone Ab.IgE|cefTRIAXone Ab.IgE
C0799717|T201|COMP|16570-4|LNC|Centromere Ab|Centromere Ab
C0799718|T201|COMP|16571-2|LNC|Cephadrine|Cephadrine
C0799719|T201|COMP|16572-0|LNC|Cephaloridine|Cephaloridine
C0799722|T201|COMP|16575-3|LNC|Cerebroside sulfatase B|Cerebroside sulfatase B
C0799723|T201|COMP|16576-1|LNC|Cerebroside sulfatase B|Cerebroside sulfatase B
C0799724|T201|COMP|16577-9|LNC|Cerebroside sulfatase B|Cerebroside sulfatase B
C0799725|T201|COMP|16578-7|LNC|Cerebroside sulfatase B|Cerebroside sulfatase B
C0799726|T201|COMP|16579-5|LNC|Cerebroside sulfatase B|Cerebroside sulfatase B
C0799727|T201|COMP|16580-3|LNC|Cerebroside sulfatase B|Cerebroside sulfatase B
C0799728|T201|COMP|16581-1|LNC|Chlamydophila pneumoniae Ab.IgA|Chlamydophila pneumoniae Ab.IgA
C0799729|T201|COMP|16582-9|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C0799730|T201|COMP|16583-7|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C0799731|T201|COMP|16584-5|LNC|Chlamydophila pneumoniae rRNA|Chlamydophila pneumoniae rRNA
C0799732|T201|COMP|16585-2|LNC|Chlamydophila pneumoniae rRNA|Chlamydophila pneumoniae rRNA
C0799733|T201|COMP|16586-0|LNC|Chlamydophila psittaci Ab.IgA|Chlamydophila psittaci Ab.IgA
C0799734|T201|COMP|16587-8|LNC|Chlamydophila psittaci Ab.IgG|Chlamydophila psittaci Ab.IgG
C0799735|T201|COMP|16588-6|LNC|Chlamydophila psittaci Ab.IgM|Chlamydophila psittaci Ab.IgM
C0799736|T201|COMP|16589-4|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0799737|T201|COMP|16590-2|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0799738|T201|COMP|16591-0|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C0799739|T201|COMP|16592-8|LNC|Chlamydia sp Ab.IgM|Chlamydia sp Ab.IgM
C0799740|T201|COMP|16593-6|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0799741|T201|COMP|16594-4|LNC|Chlamydia trachomatis Ab.IgA|Chlamydia trachomatis Ab.IgA
C0799742|T201|COMP|16595-1|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C0799743|T201|COMP|16596-9|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C0799744|T201|COMP|16597-7|LNC|Chlamydia trachomatis B Ab.IgG|Chlamydia trachomatis B Ab.IgG
C0799745|T201|COMP|16598-5|LNC|Chlamydia trachomatis C Ab.IgG|Chlamydia trachomatis C Ab.IgG
C0799746|T201|COMP|16599-3|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0799747|T201|COMP|16600-9|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C0799748|T201|COMP|16601-7|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C0799749|T201|COMP|16602-5|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C0799750|T201|COMP|16603-3|LNC|Chloramphenicol^peak|Chloramphenicol^peak
C0799751|T201|COMP|16604-1|LNC|Chloramphenicol^trough|Chloramphenicol^trough
C0799752|T201|COMP|16605-8|LNC|Chlorocycline|Chlorocycline
C0799753|T201|COMP|16606-6|LNC|Chlorine|Chlorine
C0799754|T201|COMP|16607-4|LNC|Chlorine|Chlorine
C0799755|T201|COMP|16608-2|LNC|Chlorpheniramine|Chlorpheniramine
C0799756|T201|COMP|16609-0|LNC|Chlorphentermine|Chlorphentermine
C0799757|T201|COMP|16610-8|LNC|Chlorphentermine|Chlorphentermine
C0799758|T201|COMP|16611-6|LNC|Chlorpyrifos|Chlorpyrifos
C0799759|T201|COMP|16612-4|LNC|Chlorthalidone|Chlorthalidone
C0799760|T201|COMP|16613-2|LNC|Cholesterol crystals|Cholesterol crystals
C0799761|T201|COMP|16614-0|LNC|Cholesterol crystals|Cholesterol crystals
C0799762|T201|COMP|16615-7|LNC|Cholesterol.total/Cholesterol.in LDL|Cholesterol.total/Cholesterol.in LDL
C0799763|T201|COMP|16616-5|LNC|Cholesterol.in HDL/Cholesterol.in LDL|Cholesterol.in HDL/Cholesterol.in LDL
C0799764|T201|COMP|16617-3|LNC|Choriogonadotropin.intact|Choriogonadotropin.intact
C0799765|T201|COMP|16618-1|LNC|Cladosporium herbarum Ab|Cladosporium herbarum Ab
C0799766|T201|COMP|16619-9|LNC|Clarithromycin|Clarithromycin
C0799767|T201|COMP|16620-7|LNC|Clarithromycin+Ethambutol|Clarithromycin+Ethambutol
C0799768|T201|COMP|16621-5|LNC|Clindamycin^peak|Clindamycin^peak
C0799769|T201|COMP|16622-3|LNC|Clindamycin^trough|Clindamycin^trough
C0799770|T201|COMP|16623-1|LNC|Clofazimine|Clofazimine
C0799771|T201|COMP|16624-9|LNC|clomiPRAMINE|clomiPRAMINE
C0799772|T201|COMP|16625-6|LNC|clomiPRAMINE|clomiPRAMINE
C0799773|T201|COMP|16626-4|LNC|Clostridium tetani Ab^1st specimen|Clostridium tetani Ab^1st specimen
C0799774|T201|COMP|16627-2|LNC|Clostridium tetani Ab^2nd specimen|Clostridium tetani Ab^2nd specimen
C0799775|T201|COMP|16628-0|LNC|Cloxacillin|Cloxacillin
C0799776|T201|COMP|12185-5|LNC|Coagulation surface induced|Coagulation surface induced
C0799777|T201|COMP|16630-6|LNC|Coagulation surface induced|Coagulation surface induced
C0799778|T201|COMP|16631-4|LNC|Coagulation surface induced|Coagulation surface induced
C0799779|T201|COMP|16632-2|LNC|Cocaethylene|Cocaethylene
C0799780|T201|COMP|16633-0|LNC|Cocaine|Cocaine
C0799781|T201|COMP|16634-8|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0799782|T201|COMP|16635-5|LNC|Coccidioides immitis Ab.IgA|Coccidioides immitis Ab.IgA
C0799783|T201|COMP|16636-3|LNC|Coccidioides immitis Ab.IgA|Coccidioides immitis Ab.IgA
C0799784|T201|COMP|16637-1|LNC|Coccidioides immitis Ab.IgE|Coccidioides immitis Ab.IgE
C0799785|T201|COMP|16638-9|LNC|Coccidioides immitis Ab.IgG|Coccidioides immitis Ab.IgG
C0799786|T201|COMP|16639-7|LNC|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C0799787|T201|COMP|16640-5|LNC|Coccidioides reaction wheal|Coccidioides reaction wheal
C0799788|T201|COMP|16641-3|LNC|Cockatiel droppings Ab|Cockatiel droppings Ab
C0799789|T201|COMP|16642-1|LNC|Cockatiel droppings Ab.IgG|Cockatiel droppings Ab.IgG
C0799790|T201|COMP|16643-9|LNC|Cockatoo droppings Ab|Cockatoo droppings Ab
C0799791|T201|COMP|16644-7|LNC|Codeine.free|Codeine.free
C0799792|T201|COMP|16645-4|LNC|Colistin|Colistin
C0799793|T201|COMP|16647-0|LNC|Collagen Ab|Collagen Ab
C0799794|T201|COMP|16648-8|LNC|Copper|Copper
C0799795|T201|COMP|16649-6|LNC|Coproporphyrinogen oxidase|Coproporphyrinogen oxidase
C0799796|T201|COMP|16650-4|LNC|Coriandrum sativum Ab.IgE|Coriandrum sativum Ab.IgE
C0799797|T201|COMP|16651-2|LNC|Corticosterone^post XXX challenge|Corticosterone^post XXX challenge
C0799798|T201|COMP|16652-0|LNC|Corticotropin|Corticotropin
C0799799|T201|COMP|16653-8|LNC|Corticotropin.canine|Corticotropin.canine
C0799800|T201|COMP|16654-6|LNC|Corticotropin^1.5H post XXX challenge|Corticotropin^1.5H post XXX challenge
C0799801|T201|COMP|16655-3|LNC|Corticotropin^10M post XXX challenge|Corticotropin^10M post XXX challenge
C0799802|T201|COMP|16656-1|LNC|Corticotropin^15M post XXX challenge|Corticotropin^15M post XXX challenge
C0799803|T201|COMP|16657-9|LNC|Corticotropin^1H post XXX challenge|Corticotropin^1H post XXX challenge
C0799804|T201|COMP|16658-7|LNC|Corticotropin^1M post XXX challenge|Corticotropin^1M post XXX challenge
C0799805|T201|COMP|16659-5|LNC|Corticotropin^2.5H post XXX challenge|Corticotropin^2.5H post XXX challenge
C0799806|T201|COMP|16660-3|LNC|Corticotropin^20M post XXX challenge|Corticotropin^20M post XXX challenge
C0799807|T201|COMP|16661-1|LNC|Corticotropin^2H post XXX challenge|Corticotropin^2H post XXX challenge
C0799808|T201|COMP|16662-9|LNC|Corticotropin^30M post XXX challenge|Corticotropin^30M post XXX challenge
C0799809|T201|COMP|16663-7|LNC|Corticotropin^3H post XXX challenge|Corticotropin^3H post XXX challenge
C0799810|T201|COMP|16664-5|LNC|Corticotropin^45M post XXX challenge|Corticotropin^45M post XXX challenge
C0799811|T201|COMP|16665-2|LNC|Corticotropin^5M post XXX challenge|Corticotropin^5M post XXX challenge
C0799812|T201|COMP|16666-0|LNC|Corticotropin^9th specimen post XXX challenge|Corticotropin^9th specimen post XXX challenge
C0799813|T201|COMP|16667-8|LNC|Cortisol.free|Cortisol.free
C0799814|T201|COMP|16668-6|LNC|Cortisol.free|Cortisol.free
C0799815|T201|COMP|16669-4|LNC|Cortisol^10M post XXX challenge|Cortisol^10M post XXX challenge
C0799816|T201|COMP|16670-2|LNC|Cortisol^15M post XXX challenge|Cortisol^15M post XXX challenge
C0799817|T201|COMP|16671-0|LNC|Cortisol^1M post XXX challenge|Cortisol^1M post XXX challenge
C0799818|T201|COMP|16672-8|LNC|Cortisol^40M post XXX challenge|Cortisol^40M post XXX challenge
C0799819|T201|COMP|16673-6|LNC|Cortisol^50M post XXX challenge|Cortisol^50M post XXX challenge
C0799820|T201|COMP|16674-4|LNC|Cortisol^70M post XXX challenge|Cortisol^70M post XXX challenge
C0799821|T201|COMP|16675-1|LNC|Cortisol^80M post XXX challenge|Cortisol^80M post XXX challenge
C0799822|T201|COMP|16676-9|LNC|Corynebacterium diphtheriae|Corynebacterium diphtheriae
C0799823|T201|COMP|16677-7|LNC|Coxiella burnetii Ab.IgG|Coxiella burnetii Ab.IgG
C0799824|T201|COMP|16678-5|LNC|Coxiella burnetii Ab.IgM|Coxiella burnetii Ab.IgM
C0799825|T201|COMP|16679-3|LNC|Coxsackievirus A Ab|Coxsackievirus A Ab
C0799826|T201|COMP|16680-1|LNC|Coxsackievirus A Ab.IgG|Coxsackievirus A Ab.IgG
C0799827|T201|COMP|16681-9|LNC|Coxsackievirus A Ab.IgM|Coxsackievirus A Ab.IgM
C0799828|T201|COMP|16682-7|LNC|Coxsackievirus A2 Ab|Coxsackievirus A2 Ab
C0799829|T201|COMP|16683-5|LNC|Coxsackievirus A4 Ab|Coxsackievirus A4 Ab
C0799830|T201|COMP|16684-3|LNC|Coxsackievirus B Ab|Coxsackievirus B Ab
C0799831|T201|COMP|16685-0|LNC|Coxsackievirus B Ab.IgG|Coxsackievirus B Ab.IgG
C0799832|T201|COMP|16686-8|LNC|Coxsackievirus B Ab.IgM|Coxsackievirus B Ab.IgM
C0799833|T201|COMP|16687-6|LNC|Creatine|Creatine
C0799834|T201|COMP|16688-4|LNC|Creatine kinase|Creatine kinase
C0799835|T201|COMP|16689-2|LNC|Creatinine|Creatinine
C0799836|T201|COMP|16690-0|LNC|Creatinine|Creatinine
C0799837|T201|COMP|16691-8|LNC|Cresols|Cresols
C0799838|T201|COMP|16692-6|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C0799839|T201|COMP|16693-4|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C0799840|T201|COMP|16694-2|LNC|Cumene|Cumene
C0799841|T201|COMP|16695-9|LNC|Cobalamins|Cobalamins
C0799842|T201|COMP|16696-7|LNC|Cobalamins^post XXX challenge|Cobalamins^post XXX challenge
C0799843|T201|COMP|16697-5|LNC|Cyclohexane|Cyclohexane
C0799844|T201|COMP|16698-3|LNC|Cyclohexanol|Cyclohexanol
C0799845|T201|COMP|16699-1|LNC|Cyclohexanol|Cyclohexanol
C0799846|T201|COMP|16700-7|LNC|Cyclohexanol/Creatinine|Cyclohexanol/Creatinine
C0799847|T201|COMP|16701-5|LNC|Cyclopropane|Cyclopropane
C0799848|T201|COMP|16702-3|LNC|cycloSERINE|cycloSERINE
C0799849|T201|COMP|16703-1|LNC|cycloSPORINE|cycloSPORINE
C0799850|T201|COMP|16704-9|LNC|Cyproheptadine|Cyproheptadine
C0799851|T201|COMP|16705-6|LNC|Cystathionine|Cystathionine
C0799852|T201|COMP|16706-4|LNC|Taenia solium larva Ab.IgM|Taenia solium larva Ab.IgM
C0799853|T201|COMP|16707-2|LNC|Taenia solium larva Ab.IgM|Taenia solium larva Ab.IgM
C0799855|T201|COMP|16709-8|LNC|Cystine|Cystine
C0799856|T201|COMP|16710-6|LNC|Cystine crystals|Cystine crystals
C0799857|T201|COMP|16711-4|LNC|Cystine+Homocystine|Cystine+Homocystine
C0799858|T201|COMP|16712-2|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0799859|T201|COMP|16713-0|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0799860|T201|COMP|16714-8|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0799861|T201|COMP|16715-5|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0799862|T201|COMP|16716-3|LNC|Cytomegalovirus Ab.IgG^2nd specimen|Cytomegalovirus Ab.IgG^2nd specimen
C0799863|T201|COMP|16717-1|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0799864|T201|COMP|16718-9|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C0799865|T201|COMP|16719-7|LNC|Cytomegalovirus inclusion bodies|Cytomegalovirus inclusion bodies
C0799866|T201|COMP|16720-5|LNC|Dechlorane|Dechlorane
C0799867|T201|COMP|16721-3|LNC|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C0799877|T201|COMP|16731-2|LNC|Dehydroepiandrosterone.unconjugated|Dehydroepiandrosterone.unconjugated
C0799880|T201|COMP|16734-6|LNC|Dehydroepiandrosterone^baseline|Dehydroepiandrosterone^baseline
C0799881|T201|COMP|16735-3|LNC|Dehydroepiandrosterone^post XXX challenge|Dehydroepiandrosterone^post XXX challenge
C0799882|T201|COMP|16736-1|LNC|Dengue virus 1 Ab|Dengue virus 1 Ab
C0799883|T201|COMP|16737-9|LNC|Dengue virus 2 Ab|Dengue virus 2 Ab
C0799884|T201|COMP|16738-7|LNC|Dengue virus 3 Ab|Dengue virus 3 Ab
C0799885|T201|COMP|16739-5|LNC|Dengue virus 4 Ab|Dengue virus 4 Ab
C0799886|T201|COMP|16740-3|LNC|Dengue virus Ab|Dengue virus Ab
C0799887|T201|COMP|16741-1|LNC|Dermatophagoides farinae Ab.IgG|Dermatophagoides farinae Ab.IgG
C0799888|T201|COMP|16742-9|LNC|Dermatophagoides pteronyssinus Ab.IgG|Dermatophagoides pteronyssinus Ab.IgG
C0799889|T201|COMP|16745-2|LNC|Desmethylmethsuximide|Desmethylmethsuximide
C0799890|T201|COMP|16746-0|LNC|Nortrimipramine|Nortrimipramine
C0799891|T201|COMP|16747-8|LNC|Dextromoramide|Dextromoramide
C0799892|T201|COMP|16748-6|LNC|Propoxyphene|Propoxyphene
C0799893|T201|COMP|16749-4|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C0799894|T201|COMP|16750-2|LNC|Dezocine|Dezocine
C0799895|T201|COMP|16751-0|LNC|Dezocine|Dezocine
C0799896|T201|COMP|16752-8|LNC|Diacetate|Diacetate
C0799897|T201|COMP|16753-6|LNC|Dialtrazene|Dialtrazene
C0799898|T201|COMP|16754-4|LNC|Diamorphine|Diamorphine
C0799899|T201|COMP|16755-1|LNC|Diamorphine|Diamorphine
C0799900|T201|COMP|16756-9|LNC|Diamorphine|Diamorphine
C0799901|T201|COMP|16757-7|LNC|Diazepam+Nordiazepam|Diazepam+Nordiazepam
C0799902|T201|COMP|16758-5|LNC|Dicamba|Dicamba
C0799903|T201|COMP|16759-3|LNC|Dicamba|Dicamba
C0799904|T201|COMP|16760-1|LNC|Dicarboxylporphyrin|Dicarboxylporphyrin
C0799905|T201|COMP|16761-9|LNC|Protoporphyrin|Protoporphyrin
C0799906|T201|COMP|16762-7|LNC|Dichlorobenzene|Dichlorobenzene
C0799907|T201|COMP|16763-5|LNC|Dichlorodiphenyldichloroethylene|Dichlorodiphenyldichloroethylene
C0799908|T201|COMP|16764-3|LNC|Dichlorodiphenyldichloroethylene|Dichlorodiphenyldichloroethylene
C0799909|T201|COMP|16765-0|LNC|Dichlorodiphenyltrichloroethane|Dichlorodiphenyltrichloroethane
C0799910|T201|COMP|16766-8|LNC|Dichloroethane|Dichloroethane
C0799911|T201|COMP|16767-6|LNC|2,4-Dichlorophenoxyacetate|2,4-Dichlorophenoxyacetate
C0799912|T201|COMP|16768-4|LNC|Dichlorvos|Dichlorvos
C0799913|T201|COMP|16769-2|LNC|Dicloxacillin|Dicloxacillin
C0799914|T201|COMP|16770-0|LNC|Dicoumarol|Dicoumarol
C0799915|T201|COMP|16771-8|LNC|Dicyclomine|Dicyclomine
C0799916|T201|COMP|16772-6|LNC|Dieldrin|Dieldrin
C0799917|T201|COMP|16773-4|LNC|Dieldrin|Dieldrin
C0799918|T201|COMP|16774-2|LNC|Diethylcarbamazepine|Diethylcarbamazepine
C0799919|T201|COMP|16775-9|LNC|Dihydrocodeine.free|Dihydrocodeine.free
C0799920|T201|COMP|16776-7|LNC|dilTIAZem|dilTIAZem
C0799921|T201|COMP|16777-5|LNC|Dimethylacetamide|Dimethylacetamide
C0799922|T201|COMP|16778-3|LNC|Dinitrophenol|Dinitrophenol
C0799923|T201|COMP|16779-1|LNC|Dinitrophenol|Dinitrophenol
C0799924|T201|COMP|16780-9|LNC|Disopyramide|Disopyramide
C0799925|T201|COMP|16781-7|LNC|Disulfiram|Disulfiram
C0799926|T201|COMP|16782-5|LNC|DNA double strand Ab|DNA double strand Ab
C0799927|T201|COMP|16784-1|LNC|DOPamine^2nd specimen post XXX challenge|DOPamine^2nd specimen post XXX challenge
C0799928|T201|COMP|16785-8|LNC|DOPamine^3rd specimen post XXX challenge|DOPamine^3rd specimen post XXX challenge
C0799929|T201|COMP|16786-6|LNC|DOPamine^4th specimen post XXX challenge|DOPamine^4th specimen post XXX challenge
C0799930|T201|COMP|16787-4|LNC|DOPamine^5th specimen post XXX challenge|DOPamine^5th specimen post XXX challenge
C0799931|T201|COMP|16788-2|LNC|DOPamine^6th specimen post XXX challenge|DOPamine^6th specimen post XXX challenge
C0799932|T201|COMP|16789-0|LNC|DOPamine^7th specimen post XXX challenge|DOPamine^7th specimen post XXX challenge
C0799934|T201|COMP|16791-6|LNC|Doxylamine|Doxylamine
C0799935|T201|COMP|16792-4|LNC|Doxylamine|Doxylamine
C0799936|T201|COMP|16793-2|LNC|Drugs identified|Drugs identified
C0799937|T201|COMP|16794-0|LNC|Echinococcus sp Ab.IgM|Echinococcus sp Ab.IgM
C0799939|T201|COMP|16796-5|LNC|Echovirus Ab|Echovirus Ab
C0799940|T201|COMP|16797-3|LNC|Echovirus 1 Ab|Echovirus 1 Ab
C0799941|T201|COMP|16798-1|LNC|Echovirus 14 Ab|Echovirus 14 Ab
C0799942|T201|COMP|16799-9|LNC|Echovirus 140 Ab|Echovirus 140 Ab
C0799943|T201|COMP|16800-5|LNC|Echovirus 19 Ab|Echovirus 19 Ab
C0799944|T201|COMP|16801-3|LNC|Echovirus 3 Ab|Echovirus 3 Ab
C0799945|T201|COMP|16802-1|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C0799946|T201|COMP|16803-9|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C0799947|T201|COMP|16804-7|LNC|Echovirus 40 Ab|Echovirus 40 Ab
C0799948|T201|COMP|16805-4|LNC|Echovirus 6 Ab|Echovirus 6 Ab
C0799949|T201|COMP|16806-2|LNC|Echovirus 6+18+30 Ab|Echovirus 6+18+30 Ab
C0799950|T201|COMP|16807-0|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C0799951|T201|COMP|16808-8|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C0799952|T201|COMP|16809-6|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C0799953|T201|COMP|16811-2|LNC|Arachidate|Arachidate
C0799954|T201|COMP|16812-0|LNC|Emetine|Emetine
C0799955|T201|COMP|16813-8|LNC|Emetine|Emetine
C0799956|T201|COMP|16814-6|LNC|Endomysium Ab|Endomysium Ab
C0799957|T201|COMP|16815-3|LNC|Endomysium Ab|Endomysium Ab
C0799958|T201|COMP|16816-1|LNC|Enoxacin|Enoxacin
C0799959|T201|COMP|16817-9|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0799960|T201|COMP|16818-7|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0799961|T201|COMP|16819-5|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0799962|T201|COMP|16820-3|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0799963|T201|COMP|16821-1|LNC|EPINEPHrine^4H post XXX challenge|EPINEPHrine^4H post XXX challenge
C0799964|T201|COMP|16822-9|LNC|Epithelial cells|Epithelial cells
C0799965|T201|COMP|16823-7|LNC|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C0799966|T201|COMP|16824-5|LNC|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C0799967|T201|COMP|16825-2|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0799968|T201|COMP|16826-0|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0799970|T201|COMP|16828-6|LNC|Erythrocytes|Erythrocytes
C0799971|T201|COMP|16829-4|LNC|Erythromycin|Erythromycin
C0799972|T201|COMP|16830-2|LNC|Erythromycin+Ethambutol|Erythromycin+Ethambutol
C0799973|T201|COMP|16832-8|LNC|Escherichia coli enterotoxic identified|Escherichia coli enterotoxic identified
C0799974|T201|COMP|16833-6|LNC|Escherichia coli K1 Ag|Escherichia coli K1 Ag
C0799975|T201|COMP|16834-4|LNC|Escherichia coli K1 Ag|Escherichia coli K1 Ag
C0799976|T201|COMP|16835-1|LNC|Escherichia coli shiga-like toxin identified|Escherichia coli shiga-like toxin identified
C0799977|T201|COMP|16836-9|LNC|Escherichia coli verotoxic identified|Escherichia coli verotoxic identified
C0799978|T201|COMP|16838-5|LNC|Estriol|Estriol
C0799979|T201|COMP|16840-1|LNC|Ethacrynate|Ethacrynate
C0799980|T201|COMP|16841-9|LNC|Ethambutol+rifAMPin|Ethambutol+rifAMPin
C0799981|T201|COMP|16842-7|LNC|Ethanol|Ethanol
C0799982|T201|COMP|16843-5|LNC|Ethanol|Ethanol
C0799983|T201|COMP|16844-3|LNC|Ethinamate|Ethinamate
C0799984|T201|COMP|16845-0|LNC|Ethionamide|Ethionamide
C0799985|T201|COMP|16847-6|LNC|Ethoheptazine|Ethoheptazine
C0799986|T201|COMP|16848-4|LNC|Ethoheptazine|Ethoheptazine
C0799987|T201|COMP|16849-2|LNC|Ethyl benzene|Ethyl benzene
C0799988|T201|COMP|16850-0|LNC|Ethylene oxide|Ethylene oxide
C0799989|T201|COMP|16851-8|LNC|Ethylmorphine|Ethylmorphine
C0799990|T201|COMP|16852-6|LNC|Etodolac|Etodolac
C0799993|T201|COMP|16856-7|LNC|Fat.microscopic observation|Fat.microscopic observation
C0799994|T201|COMP|16857-5|LNC|Fenclorvos|Fenclorvos
C0799995|T201|COMP|16858-3|LNC|fentaNYL|fentaNYL
C0799996|T201|COMP|16859-1|LNC|Fibrinogen|Fibrinogen
C0799997|T201|COMP|16860-9|LNC|Fibrinopeptide A Ag|Fibrinopeptide A Ag
C0799998|T201|COMP|16861-7|LNC|Fibrinopeptide A Ag|Fibrinopeptide A Ag
C0799999|T201|COMP|16862-5|LNC|Fibrinopeptide B Ag|Fibrinopeptide B Ag
C0800000|T201|COMP|16863-3|LNC|Fibrinopeptide B beta (1-14) Ag|Fibrinopeptide B beta (1-14) Ag
C0800001|T201|COMP|16864-1|LNC|Fibrinopeptide B beta (1-42) Ag|Fibrinopeptide B beta (1-42) Ag
C0800002|T201|COMP|16865-8|LNC|Fibrinopeptide B beta (15-42) Ag|Fibrinopeptide B beta (15-42) Ag
C0800003|T201|COMP|16866-6|LNC|Fibrinopeptide B beta (43-47) Ag|Fibrinopeptide B beta (43-47) Ag
C0800004|T201|COMP|16867-4|LNC|Fibronectin aggregate Ab.IgG|Fibronectin aggregate Ab.IgG
C0800005|T201|COMP|16868-2|LNC|Finch droppings Ab.IgE|Finch droppings Ab.IgE
C0800006|T201|COMP|16869-0|LNC|Flubiprofen|Flubiprofen
C0800007|T201|COMP|16870-8|LNC|Fluconazole|Fluconazole
C0800008|T201|COMP|16871-6|LNC|Fluoride|Fluoride
C0800009|T201|COMP|16872-4|LNC|Fluorocarbons|Fluorocarbons
C0800010|T201|COMP|16873-2|LNC|Follitropin^105M post XXX challenge|Follitropin^105M post XXX challenge
C0800011|T201|COMP|16874-0|LNC|Formate+Formaldehyde|Formate+Formaldehyde
C0800012|T201|COMP|16875-7|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C0800013|T201|COMP|16876-5|LNC|Francisella tularensis Ab.IgA|Francisella tularensis Ab.IgA
C0800014|T201|COMP|16877-3|LNC|Francisella tularensis Ab.IgG|Francisella tularensis Ab.IgG
C0800015|T201|COMP|16878-1|LNC|Francisella tularensis Ab.IgM|Francisella tularensis Ab.IgM
C0800016|T201|COMP|16879-9|LNC|Francisella tularensis Ag|Francisella tularensis Ag
C0800017|T201|COMP|16881-5|LNC|Gallium|Gallium
C0800018|T201|COMP|16882-3|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0800023|T201|COMP|16887-2|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0800024|T201|COMP|16888-0|LNC|Gamma chlordane|Gamma chlordane
C0800025|T201|COMP|16890-6|LNC|Gastrin^10M post XXX challenge|Gastrin^10M post XXX challenge
C0800026|T201|COMP|16891-4|LNC|Gastrin^11th specimen post XXX challenge|Gastrin^11th specimen post XXX challenge
C0800027|T201|COMP|16892-2|LNC|Gastrin^15M post XXX challenge|Gastrin^15M post XXX challenge
C0800028|T201|COMP|16893-0|LNC|Gastrin^20M post XXX challenge|Gastrin^20M post XXX challenge
C0800029|T201|COMP|16894-8|LNC|Gastrin^25M post XXX challenge|Gastrin^25M post XXX challenge
C0800030|T201|COMP|16895-5|LNC|Gastrin^30M post XXX challenge|Gastrin^30M post XXX challenge
C0800031|T201|COMP|16896-3|LNC|Gastrin^5M post XXX challenge|Gastrin^5M post XXX challenge
C0800032|T201|COMP|16898-9|LNC|Giardia lamblia 65 Ag|Giardia lamblia 65 Ag
C0800033|T201|COMP|16899-7|LNC|Giardia lamblia Ag|Giardia lamblia Ag
C0800034|T201|COMP|16900-3|LNC|Gliadin Ab|Gliadin Ab
C0800035|T201|COMP|16901-1|LNC|Gliadin Ab.IgA|Gliadin Ab.IgA
C0800036|T201|COMP|16902-9|LNC|Gliadin Ab.IgG|Gliadin Ab.IgG
C0800037|T201|COMP|16903-7|LNC|Glucose|Glucose
C0800038|T201|COMP|16904-5|LNC|Glucose^1st specimen post XXX challenge|Glucose^1st specimen post XXX challenge
C0800039|T201|COMP|16905-2|LNC|Glucose^2nd specimen post XXX challenge|Glucose^2nd specimen post XXX challenge
C0800040|T201|COMP|16906-0|LNC|Glucose^3rd specimen post XXX challenge|Glucose^3rd specimen post XXX challenge
C0800041|T201|COMP|16907-8|LNC|Glucose^4th specimen post XXX challenge|Glucose^4th specimen post XXX challenge
C0800042|T201|COMP|16908-6|LNC|Glucose^5th specimen post XXX challenge|Glucose^5th specimen post XXX challenge
C0800043|T201|COMP|16909-4|LNC|Glucose^6th specimen post XXX challenge|Glucose^6th specimen post XXX challenge
C0800044|T201|COMP|16910-2|LNC|Glucose^7th specimen post XXX challenge|Glucose^7th specimen post XXX challenge
C0800045|T201|COMP|16911-0|LNC|Glucose^8th specimen post XXX challenge|Glucose^8th specimen post XXX challenge
C0800046|T201|COMP|16912-8|LNC|Glucose^9th specimen post XXX challenge|Glucose^9th specimen post XXX challenge
C0800047|T201|COMP|16913-6|LNC|Glucose^post CFst|Glucose^post CFst
C0800048|T201|COMP|16914-4|LNC|Glucose^post XXX challenge|Glucose^post XXX challenge
C0800049|T201|COMP|16915-1|LNC|Glucose^post meal|Glucose^post meal
C0800050|T201|COMP|16916-9|LNC|Glutamate|Glutamate
C0800051|T201|COMP|16917-7|LNC|Glutamine|Glutamine
C0800052|T201|COMP|16918-5|LNC|Glutathione|Glutathione
C0800053|T201|COMP|16919-3|LNC|Glycine|Glycine
C0800054|T201|COMP|16920-1|LNC|Glycoproteins|Glycoproteins
C0800055|T201|COMP|16921-9|LNC|Stenotaphrum secundatum Ab.IgE|Stenotaphrum secundatum Ab.IgE
C0800057|T201|COMP|16923-5|LNC|guaiFENesin|guaiFENesin
C0800058|T201|COMP|16924-3|LNC|Haemophilus influenzae Ab.IgG|Haemophilus influenzae Ab.IgG
C0800059|T201|COMP|16925-0|LNC|Haemophilus influenzae A Ag|Haemophilus influenzae A Ag
C0800060|T201|COMP|16926-8|LNC|Haemophilus influenzae A Ag|Haemophilus influenzae A Ag
C0800061|T201|COMP|16927-6|LNC|Haemophilus influenzae B Ab.IgG|Haemophilus influenzae B Ab.IgG
C0800062|T201|COMP|16928-4|LNC|Hantavirus puumala Ab.IgG+IgM|Hantavirus puumala Ab.IgG+IgM
C0800063|T201|COMP|16929-2|LNC|Helicobacter pylori Ab|Helicobacter pylori Ab
C0800064|T201|COMP|16930-0|LNC|Helminth Ab.IgE|Helminth Ab.IgE
C0800065|T201|COMP|16931-8|LNC|Hematocrit/Hemoglobin|Hematocrit/Hemoglobin
C0800066|T201|COMP|16932-6|LNC|Hemoglobin A3/Hemoglobin.total|Hemoglobin A3/Hemoglobin.total
C0800067|T201|COMP|16933-4|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C0800068|T201|COMP|16934-2|LNC|Hepatitis B virus polymerase DNA|Hepatitis B virus polymerase DNA
C0800069|T201|COMP|16935-9|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0800070|T201|COMP|16936-7|LNC|Hepatitis C virus Ab.IgG|Hepatitis C virus Ab.IgG
C0800071|T201|COMP|16937-5|LNC|Hepatitis G virus RNA|Hepatitis G virus RNA
C0800072|T201|COMP|16938-3|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C0800073|T201|COMP|16939-1|LNC|Heptachlor|Heptachlor
C0800074|T201|COMP|16940-9|LNC|Heptachlorepoxide|Heptachlorepoxide
C0800076|T201|COMP|16942-5|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C0800077|T201|COMP|16943-3|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C0800078|T201|COMP|16944-1|LNC|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C0800079|T201|COMP|16945-8|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C0800080|T201|COMP|16947-4|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C0800081|T201|COMP|16948-2|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C0800082|T201|COMP|16949-0|LNC|Herpes simplex virus 1 Ab.IgG^1st specimen|Herpes simplex virus 1 Ab.IgG^1st specimen
C0800083|T201|COMP|16950-8|LNC|Herpes simplex virus 1 Ab.IgG^2nd specimen|Herpes simplex virus 1 Ab.IgG^2nd specimen
C0800084|T201|COMP|16952-4|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C0800085|T201|COMP|16953-2|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C0800086|T201|COMP|16954-0|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C0800087|T201|COMP|16955-7|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0800088|T201|COMP|16956-5|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0800089|T201|COMP|16957-3|LNC|Herpes simplex virus 2 Ab.IgG^1st specimen|Herpes simplex virus 2 Ab.IgG^1st specimen
C0800090|T201|COMP|16958-1|LNC|Herpes simplex virus 2 Ab.IgG^2nd specimen|Herpes simplex virus 2 Ab.IgG^2nd specimen
C0800091|T201|COMP|16959-9|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C0800092|T201|COMP|16960-7|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C0800093|T201|COMP|16962-3|LNC|Heterophile Ab|Heterophile Ab
C0800094|T201|COMP|16963-1|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C0800095|T201|COMP|16964-9|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C0800096|T201|COMP|16965-6|LNC|Lindane|Lindane
C0800097|T201|COMP|16966-4|LNC|Hexachloroethane|Hexachloroethane
C0800098|T201|COMP|16967-2|LNC|Hexokinase 1|Hexokinase 1
C0800099|T201|COMP|16968-0|LNC|Hexokinase 3|Hexokinase 3
C0800100|T201|COMP|16969-8|LNC|Histone H2a+H2b Ab|Histone H2a+H2b Ab
C0800101|T201|COMP|16970-6|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0800102|T201|COMP|16971-4|LNC|Histoplasma capsulatum Ab.IgA|Histoplasma capsulatum Ab.IgA
C0800103|T201|COMP|16972-2|LNC|Histoplasma capsulatum Ab.IgE|Histoplasma capsulatum Ab.IgE
C0800104|T201|COMP|16973-0|LNC|Histoplasma capsulatum Ab.IgM|Histoplasma capsulatum Ab.IgM
C0800105|T201|COMP|16974-8|LNC|HIV 1 Ab|HIV 1 Ab
C0800106|T201|COMP|16975-5|LNC|HIV 1 Ab.IgG|HIV 1 Ab.IgG
C0800107|T201|COMP|16976-3|LNC|HIV 1 Ag|HIV 1 Ag
C0800108|T201|COMP|16977-1|LNC|HIV 1 Ag|HIV 1 Ag
C0800109|T201|COMP|16978-9|LNC|HIV 1 p24 Ab|HIV 1 p24 Ab
C0800110|T201|COMP|16979-7|LNC|HIV 1 p24 Ag|HIV 1 p24 Ag
C0800111|T201|COMP|16980-5|LNC|HTLV II DNA|HTLV II DNA
C0800112|T201|COMP|16981-3|LNC|HTLV I DNA|HTLV I DNA
C0800113|T201|COMP|16982-1|LNC|HTLV I+II Ab|HTLV I+II Ab
C0800114|T201|COMP|16983-9|LNC|hydrALAZINE|hydrALAZINE
C0800115|T201|COMP|16984-7|LNC|Hydrastine|Hydrastine
C0800116|T201|COMP|16985-4|LNC|Hydrogen/Expired gas^1.5H post dose glucose|Hydrogen/Expired gas^1.5H post dose glucose
C0800117|T201|COMP|16986-2|LNC|Hydrogen/Expired gas^1H post dose glucose|Hydrogen/Expired gas^1H post dose glucose
C0800118|T201|COMP|16987-0|LNC|Hydrogen/Expired gas^2.5H post dose glucose|Hydrogen/Expired gas^2.5H post dose glucose
C0800119|T201|COMP|16988-8|LNC|Hydrogen/Expired gas^2H post dose glucose|Hydrogen/Expired gas^2H post dose glucose
C0800120|T201|COMP|16989-6|LNC|Hydrogen/Expired gas^3.5H post dose glucose|Hydrogen/Expired gas^3.5H post dose glucose
C0800121|T201|COMP|16990-4|LNC|Hydrogen/Expired gas^3H post dose glucose|Hydrogen/Expired gas^3H post dose glucose
C0800122|T201|COMP|16991-2|LNC|Hydrogen/Expired gas^4.5H post dose glucose|Hydrogen/Expired gas^4.5H post dose glucose
C0800123|T201|COMP|16992-0|LNC|Hydrogen/Expired gas^4H post dose glucose|Hydrogen/Expired gas^4H post dose glucose
C0800124|T201|COMP|16993-8|LNC|Hydrogen/Expired gas^5.5H post dose glucose|Hydrogen/Expired gas^5.5H post dose glucose
C0800125|T201|COMP|16994-6|LNC|Hydrogen/Expired gas^5H post dose glucose|Hydrogen/Expired gas^5H post dose glucose
C0800126|T201|COMP|16995-3|LNC|Hydrogen/Expired gas^6H post dose glucose|Hydrogen/Expired gas^6H post dose glucose
C0800127|T201|COMP|16996-1|LNC|Hydrogen/Expired gas^pre dose glucose|Hydrogen/Expired gas^pre dose glucose
C0800128|T201|COMP|16997-9|LNC|Hydrogen/Expired gas^post dose glucose|Hydrogen/Expired gas^post dose glucose
C0800129|T201|COMP|16998-7|LNC|HYDROmorphone|HYDROmorphone
C0800130|T201|COMP|16999-5|LNC|Hydroquinone|Hydroquinone
C0800131|T201|COMP|17000-1|LNC|Hydroxylysine|Hydroxylysine
C0800132|T201|COMP|17001-9|LNC|Hydroxyproline|Hydroxyproline
C0800133|T201|COMP|17002-7|LNC|Hydroxytriazolam|Hydroxytriazolam
C0800135|T201|COMP|17004-3|LNC|Hypoxanthine|Hypoxanthine
C0800136|T201|COMP|17005-0|LNC|IgA subclass 1|IgA subclass 1
C0800137|T201|COMP|17006-8|LNC|IgA subclass 2|IgA subclass 2
C0800138|T201|COMP|17007-6|LNC|IgG|IgG
C0800139|T201|COMP|17008-4|LNC|IgG/Beta tubulin|IgG/Beta tubulin
C0800140|T201|COMP|17009-2|LNC|IgM|IgM
C0800141|T201|COMP|17010-0|LNC|Imipenem|Imipenem
C0800142|T201|COMP|17012-6|LNC|Influenza virus A Ab|Influenza virus A Ab
C0800143|T201|COMP|17013-4|LNC|Influenza virus A+B Ab|Influenza virus A+B Ab
C0800144|T201|COMP|17014-2|LNC|Influenza virus B Ab|Influenza virus B Ab
C0800145|T201|COMP|17015-9|LNC|Influenza virus B Ab.IgG|Influenza virus B Ab.IgG
C0800146|T201|COMP|17016-7|LNC|Influenza virus B Ab.IgM|Influenza virus B Ab.IgM
C0800147|T201|COMP|17017-5|LNC|Insulin^10M post XXX challenge|Insulin^10M post XXX challenge
C0800148|T201|COMP|17018-3|LNC|Insulin^20M post XXX challenge|Insulin^20M post XXX challenge
C0800150|T201|COMP|17020-9|LNC|Intercellular substance Ab|Intercellular substance Ab
C0800151|T201|COMP|17021-7|LNC|Intercellular substance Ab|Intercellular substance Ab
C0800152|T201|COMP|17022-5|LNC|Interleukin 1+2|Interleukin 1+2
C0800153|T201|COMP|17024-1|LNC|Iodine.inorganic|Iodine.inorganic
C0800154|T201|COMP|17025-8|LNC|Iron|Iron
C0800155|T201|COMP|17026-6|LNC|Isocyanate Ab.IgE|Isocyanate Ab.IgE
C0800156|T201|COMP|17027-4|LNC|Isocyanate Ab.IgG|Isocyanate Ab.IgG
C0800157|T201|COMP|17028-2|LNC|Isocyanate Ab.IgM|Isocyanate Ab.IgM
C0800158|T201|COMP|17029-0|LNC|Isoleucine|Isoleucine
C0800159|T201|COMP|17030-8|LNC|Isopropyl ether|Isopropyl ether
C0800160|T201|COMP|17031-6|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C0800161|T201|COMP|17032-4|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C0800162|T201|COMP|17033-2|LNC|Ketamine|Ketamine
C0800163|T201|COMP|17034-0|LNC|Ketoprofen|Ketoprofen
C0800164|T201|COMP|17035-7|LNC|Ketorolac|Ketorolac
C0800165|T201|COMP|17036-5|LNC|La Crosse virus Ab|La Crosse virus Ab
C0800166|T201|COMP|17037-3|LNC|La Crosse virus Ab|La Crosse virus Ab
C0800169|T201|COMP|17040-7|LNC|Labetalol|Labetalol
C0800170|T201|COMP|17041-5|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C0800171|T201|COMP|17042-3|LNC|Lactoglobulin Ab.IgE|Lactoglobulin Ab.IgE
C0800172|T201|COMP|17043-1|LNC|Lactose|Lactose
C0800173|T201|COMP|17044-9|LNC|Lamellar bodies|Lamellar bodies
C0800174|T201|COMP|17045-6|LNC|Latex Ab.IgE|Latex Ab.IgE
C0800175|T201|COMP|17046-4|LNC|Latex Ab.IgG|Latex Ab.IgG
C0800176|T201|COMP|17047-2|LNC|Latex Bencard Ab.IgE|Latex Bencard Ab.IgE
C0800177|T201|COMP|17048-0|LNC|Latex glove extract Ab.IgE|Latex glove extract Ab.IgE
C0800178|T201|COMP|17049-8|LNC|Latex glove extract ammoniated Ab.IgE|Latex glove extract ammoniated Ab.IgE
C0800179|T201|COMP|17050-6|LNC|Latex glove extract buffered Ab.IgE|Latex glove extract buffered Ab.IgE
C0800180|T201|COMP|17051-4|LNC|Laxatives|Laxatives
C0800181|T201|COMP|17052-2|LNC|Lead|Lead
C0800182|T201|COMP|17053-0|LNC|Legionella longbeachae 1 Ab.IgG|Legionella longbeachae 1 Ab.IgG
C0800183|T201|COMP|17054-8|LNC|Legionella longbeachae 1 Ab.IgM|Legionella longbeachae 1 Ab.IgM
C0800184|T201|COMP|17055-5|LNC|Legionella longbeachae 2 Ab.IgG|Legionella longbeachae 2 Ab.IgG
C0800185|T201|COMP|17056-3|LNC|Legionella longbeachae 2 Ab.IgM|Legionella longbeachae 2 Ab.IgM
C0800186|T201|COMP|17057-1|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C0800187|T201|COMP|17058-9|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C0800188|T201|COMP|17059-7|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C0800189|T201|COMP|17060-5|LNC|Legionella pneumophila 1 Ab|Legionella pneumophila 1 Ab
C0800190|T201|COMP|17061-3|LNC|Legionella pneumophila 1 Ab.IgM|Legionella pneumophila 1 Ab.IgM
C0800191|T201|COMP|17062-1|LNC|Legionella pneumophila 2 Ab|Legionella pneumophila 2 Ab
C0800192|T201|COMP|17063-9|LNC|Legionella pneumophila 2 Ab.IgM|Legionella pneumophila 2 Ab.IgM
C0800193|T201|COMP|17064-7|LNC|Legionella pneumophila 3 Ab|Legionella pneumophila 3 Ab
C0800194|T201|COMP|17065-4|LNC|Legionella pneumophila 3 Ab.IgM|Legionella pneumophila 3 Ab.IgM
C0800195|T201|COMP|17066-2|LNC|Legionella pneumophila 4 Ab|Legionella pneumophila 4 Ab
C0800196|T201|COMP|17067-0|LNC|Legionella pneumophila 4 Ab.IgM|Legionella pneumophila 4 Ab.IgM
C0800197|T201|COMP|17068-8|LNC|Legionella pneumophila 5 Ab|Legionella pneumophila 5 Ab
C0800198|T201|COMP|17069-6|LNC|Legionella pneumophila 5 Ab.IgM|Legionella pneumophila 5 Ab.IgM
C0800199|T201|COMP|17070-4|LNC|Legionella pneumophila 6 Ab|Legionella pneumophila 6 Ab
C0800200|T201|COMP|17071-2|LNC|Legionella pneumophila 7 Ab|Legionella pneumophila 7 Ab
C0800201|T201|COMP|17072-0|LNC|Legionella pneumophila 8 Ab|Legionella pneumophila 8 Ab
C0800202|T201|COMP|17073-8|LNC|Legionella pneumophila 9 Ab|Legionella pneumophila 9 Ab
C0800203|T201|COMP|17074-6|LNC|Leucine|Leucine
C0800204|T201|COMP|17075-3|LNC|Lidocaine|Lidocaine
C0800205|T201|COMP|17076-1|LNC|Lidocaine|Lidocaine
C0800207|T201|COMP|17078-7|LNC|Fatty acids.esterified|Fatty acids.esterified
C0800208|T201|COMP|17079-5|LNC|Fatty acids.long chain|Fatty acids.long chain
C0800209|T201|COMP|17080-3|LNC|Fatty acids.very long chain|Fatty acids.very long chain
C0800210|T201|COMP|17081-1|LNC|Triglyceride^post CFst|Triglyceride^post CFst
C0800211|T201|COMP|17082-9|LNC|Lipoprotein.alpha|Lipoprotein.alpha
C0800212|T201|COMP|17083-7|LNC|Lipoprotein.beta|Lipoprotein.beta
C0800213|T201|COMP|17084-5|LNC|Lipoprotein.pre-beta|Lipoprotein.pre-beta
C0800214|T201|COMP|17085-2|LNC|Lipoprotein|Lipoprotein
C0800215|T201|COMP|17086-0|LNC|Lithium|Lithium
C0800216|T201|COMP|17087-8|LNC|Loperamide|Loperamide
C0800217|T201|COMP|17088-6|LNC|LORazepam|LORazepam
C0800218|T201|COMP|17089-4|LNC|Lorcainide|Lorcainide
C0800219|T201|COMP|17090-2|LNC|Loxapine+8-Hydroxyloxapine|Loxapine+8-Hydroxyloxapine
C0800220|T201|COMP|17091-0|LNC|Lumpfish roe Ab.IgE|Lumpfish roe Ab.IgE
C0800221|T201|COMP|17092-8|LNC|Lupus erythematosus factor|Lupus erythematosus factor
C0800222|T201|COMP|17094-4|LNC|Lutropin^105M post XXX challenge|Lutropin^105M post XXX challenge
C0800223|T201|COMP|17095-1|LNC|Lutropin^75M post XXX challenge|Lutropin^75M post XXX challenge
C0800224|T201|COMP|17096-9|LNC|Lymphocytes.kappa/100 lymphocytes|Lymphocytes.kappa/100 lymphocytes
C0800225|T201|COMP|33596-8|LNC|Cells.CD10+CD20+|Cells.CD10+CD20+
C0800226|T201|COMP|17098-5|LNC|Cells.CD100/100 cells|Cells.CD100/100 cells
C0800227|T201|COMP|17099-3|LNC|Cells.CD102/100 cells|Cells.CD102/100 cells
C0800228|T201|COMP|17100-9|LNC|Cells.CD103/100 cells|Cells.CD103/100 cells
C0800229|T201|COMP|17101-7|LNC|Cells.CD104/100 cells|Cells.CD104/100 cells
C0800230|T201|COMP|17102-5|LNC|Cells.CD105/100 cells|Cells.CD105/100 cells
C0800231|T201|COMP|17103-3|LNC|Cells.CD106/100 cells|Cells.CD106/100 cells
C0800232|T201|COMP|17104-1|LNC|Cells.CD107a/100 cells|Cells.CD107a/100 cells
C0800233|T201|COMP|17105-8|LNC|Cells.CD107b/100 cells|Cells.CD107b/100 cells
C0800234|T201|COMP|17106-6|LNC|Cells.CD115/100 cells|Cells.CD115/100 cells
C0800235|T201|COMP|17107-4|LNC|Cells.CD117/100 cells|Cells.CD117/100 cells
C0800236|T201|COMP|17108-2|LNC|Cells.CD118/100 cells|Cells.CD118/100 cells
C0800237|T201|COMP|17109-0|LNC|Cells.CD11a/100 cells|Cells.CD11a/100 cells
C0800238|T201|COMP|17110-8|LNC|Cells.CD11b/100 cells|Cells.CD11b/100 cells
C0800239|T201|COMP|17111-6|LNC|Cells.CD12/100 cells|Cells.CD12/100 cells
C0800240|T201|COMP|17112-4|LNC|Cells.CD120a/100 cells|Cells.CD120a/100 cells
C0800241|T201|COMP|17113-2|LNC|Cells.CD120b/100 cells|Cells.CD120b/100 cells
C0800242|T201|COMP|17114-0|LNC|Cells.CD122/100 cells|Cells.CD122/100 cells
C0800243|T201|COMP|17115-7|LNC|Cells.CD126/100 cells|Cells.CD126/100 cells
C0800244|T201|COMP|17116-5|LNC|Cells.CD128/100 cells|Cells.CD128/100 cells
C0800245|T201|COMP|17117-3|LNC|Cells.CD15/100 cells|Cells.CD15/100 cells
C0800246|T201|COMP|17118-1|LNC|Cells.CD16b/100 cells|Cells.CD16b/100 cells
C0800247|T201|COMP|17119-9|LNC|Cells.CD16-CD34+/100 cells|Cells.CD16-CD34+/100 cells
C0800248|T201|COMP|17120-7|LNC|Cells.CD17/100 cells|Cells.CD17/100 cells
C0800249|T201|COMP|17121-5|LNC|Cells.CD18/100 cells|Cells.CD18/100 cells
C0800250|T201|COMP|17122-3|LNC|Cells.CD19+Kappa+/100 cells|Cells.CD19+Kappa+/100 cells
C0800251|T201|COMP|17123-1|LNC|Cells.CD19+Lambda+/100 cells|Cells.CD19+Lambda+/100 cells
C0800252|T201|COMP|17124-9|LNC|Cells.CD2+CD20+/100 cells|Cells.CD2+CD20+/100 cells
C0800253|T201|COMP|17125-6|LNC|Cells.CD22+CD19+/100 cells|Cells.CD22+CD19+/100 cells
C0800254|T201|COMP|17126-4|LNC|Cells.CD24/100 cells|Cells.CD24/100 cells
C0800255|T201|COMP|17127-2|LNC|Cells.CD26/100 cells|Cells.CD26/100 cells
C0800256|T201|COMP|17128-0|LNC|Cells.CD27/100 cells|Cells.CD27/100 cells
C0800257|T201|COMP|17129-8|LNC|Cells.CD28/100 cells|Cells.CD28/100 cells
C0800258|T201|COMP|17130-6|LNC|Cells.CD29/100 cells|Cells.CD29/100 cells
C0800259|T201|COMP|17131-4|LNC|Cells.CD3+CD69+/100 cells|Cells.CD3+CD69+/100 cells
C0800260|T201|COMP|17132-2|LNC|Cells.CD3+IL2R1+/100 cells|Cells.CD3+IL2R1+/100 cells
C0800261|T201|COMP|17133-0|LNC|Cells.CD3+CD16+/100 cells|Cells.CD3+CD16+/100 cells
C0800262|T201|COMP|17135-5|LNC|Cells.CD3+CD56+/100 cells|Cells.CD3+CD56+/100 cells
C0800263|T201|COMP|17136-3|LNC|Cells.CD3+DR+/100 cells|Cells.CD3+DR+/100 cells
C0800264|T201|COMP|17137-1|LNC|Cells.CD30/100 cells|Cells.CD30/100 cells
C0800265|T201|COMP|17138-9|LNC|Cells.CD31/100 cells|Cells.CD31/100 cells
C0800266|T201|COMP|17139-7|LNC|Cells.CD32/100 cells|Cells.CD32/100 cells
C0800267|T201|COMP|17140-5|LNC|Cells.CD34+DR+/100 cells|Cells.CD34+DR+/100 cells
C0800268|T201|COMP|17141-3|LNC|Cells.CD36/100 cells|Cells.CD36/100 cells
C0800269|T201|COMP|17142-1|LNC|Cells.CD37/100 cells|Cells.CD37/100 cells
C0800270|T201|COMP|17143-9|LNC|Cells.CD39/100 cells|Cells.CD39/100 cells
C0800271|T201|COMP|17144-7|LNC|Cells.CD4+CD69+/100 cells|Cells.CD4+CD69+/100 cells
C0800272|T201|COMP|17145-4|LNC|Cells.CD4+2H4/100 cells|Cells.CD4+2H4/100 cells
C0800273|T201|COMP|17146-2|LNC|Cells.CD4+CD8+/100 cells|Cells.CD4+CD8+/100 cells
C0800274|T201|COMP|17147-0|LNC|Cells.CD40/100 cells|Cells.CD40/100 cells
C0800275|T201|COMP|17148-8|LNC|Cells.CD41/100 cells|Cells.CD41/100 cells
C0800276|T201|COMP|17149-6|LNC|Cells.CD42a/100 cells|Cells.CD42a/100 cells
C0800277|T201|COMP|17150-4|LNC|Cells.CD42b/100 cells|Cells.CD42b/100 cells
C0800278|T201|COMP|17151-2|LNC|Cells.CD42c/100 cells|Cells.CD42c/100 cells
C0800279|T201|COMP|17152-0|LNC|Cells.CD42d/100 cells|Cells.CD42d/100 cells
C0800280|T201|COMP|17153-8|LNC|Cells.CD4+CD45RA+/Cells.CD8|Cells.CD4+CD45RA+/Cells.CD8
C0800281|T201|COMP|17154-6|LNC|Cells.CD43/100 cells|Cells.CD43/100 cells
C0800282|T201|COMP|17155-3|LNC|Cells.CD44/100 cells|Cells.CD44/100 cells
C0800283|T201|COMP|17156-1|LNC|Cells.CD44R/100 cells|Cells.CD44R/100 cells
C0800284|T201|COMP|17157-9|LNC|Cells.CD45RA/100 cells|Cells.CD45RA/100 cells
C0800285|T201|COMP|17158-7|LNC|Cells.CD45RB/100 cells|Cells.CD45RB/100 cells
C0800286|T201|COMP|17159-5|LNC|Cells.CD45RO/100 cells|Cells.CD45RO/100 cells
C0800287|T201|COMP|17160-3|LNC|Cells.CD46/100 cells|Cells.CD46/100 cells
C0800288|T201|COMP|17161-1|LNC|Cells.CD47/100 cells|Cells.CD47/100 cells
C0800289|T201|COMP|17162-9|LNC|Cells.CD48/100 cells|Cells.CD48/100 cells
C0800290|T201|COMP|17163-7|LNC|Cells.CD49a/100 cells|Cells.CD49a/100 cells
C0800291|T201|COMP|17164-5|LNC|Cells.CD49b/100 cells|Cells.CD49b/100 cells
C0800292|T201|COMP|17165-2|LNC|Cells.CD49c/100 cells|Cells.CD49c/100 cells
C0800293|T201|COMP|17166-0|LNC|Cells.CD49d/100 cells|Cells.CD49d/100 cells
C0800294|T201|COMP|17167-8|LNC|Cells.CD49e/100 cells|Cells.CD49e/100 cells
C0800295|T201|COMP|17168-6|LNC|Cells.CD49f/100 cells|Cells.CD49f/100 cells
C0800296|T201|COMP|17169-4|LNC|Cells.CD5+CD2-/100 cells|Cells.CD5+CD2-/100 cells
C0800297|T201|COMP|17170-2|LNC|Cells.CD50/100 cells|Cells.CD50/100 cells
C0800298|T201|COMP|17171-0|LNC|Cells.CD51/100 cells|Cells.CD51/100 cells
C0800299|T201|COMP|17172-8|LNC|Cells.CD52/100 cells|Cells.CD52/100 cells
C0800300|T201|COMP|17173-6|LNC|Cells.CD53/100 cells|Cells.CD53/100 cells
C0800301|T201|COMP|17174-4|LNC|Cells.CD54/100 cells|Cells.CD54/100 cells
C0800302|T201|COMP|17175-1|LNC|Cells.CD55/100 cells|Cells.CD55/100 cells
C0800303|T201|COMP|17176-9|LNC|Cells.CD58/100 cells|Cells.CD58/100 cells
C0800304|T201|COMP|17177-7|LNC|Cells.CD59/100 cells|Cells.CD59/100 cells
C0800305|T201|COMP|17178-5|LNC|Cells.CD6/100 cells|Cells.CD6/100 cells
C0800306|T201|COMP|17179-3|LNC|Cells.CD62E/100 cells|Cells.CD62E/100 cells
C0800307|T201|COMP|17180-1|LNC|Cells.CD62L/100 cells|Cells.CD62L/100 cells
C0800308|T201|COMP|17181-9|LNC|Cells.CD62P/100 cells|Cells.CD62P/100 cells
C0800309|T201|COMP|17182-7|LNC|Cells.CD63/100 cells|Cells.CD63/100 cells
C0800310|T201|COMP|17183-5|LNC|Cells.CD64/100 cells|Cells.CD64/100 cells
C0800311|T201|COMP|17184-3|LNC|Cells.CD66a/100 cells|Cells.CD66a/100 cells
C0800312|T201|COMP|17185-0|LNC|Cells.CD66b/100 cells|Cells.CD66b/100 cells
C0800313|T201|COMP|17186-8|LNC|Cells.CD66c/100 cells|Cells.CD66c/100 cells
C0800314|T201|COMP|17187-6|LNC|Cells.CD66d/100 cells|Cells.CD66d/100 cells
C0800315|T201|COMP|17188-4|LNC|Cells.CD66e/100 cells|Cells.CD66e/100 cells
C0800316|T201|COMP|17189-2|LNC|Cells.CD68/100 cells|Cells.CD68/100 cells
C0800317|T201|COMP|17190-0|LNC|Cells.CD69/100 cells|Cells.CD69/100 cells
C0800318|T201|COMP|17191-8|LNC|Cells.CD3-CD7+/100 cells|Cells.CD3-CD7+/100 cells
C0800319|T201|COMP|17192-6|LNC|Cells.CD72/100 cells|Cells.CD72/100 cells
C0800320|T201|COMP|17193-4|LNC|Cells.CD73/100 cells|Cells.CD73/100 cells
C0800321|T201|COMP|17194-2|LNC|Cells.CD74/100 cells|Cells.CD74/100 cells
C0800322|T201|COMP|17195-9|LNC|Cells.CD77/100 cells|Cells.CD77/100 cells
C0800323|T201|COMP|17196-7|LNC|Cells.CD79a/100 cells|Cells.CD79a/100 cells
C0800324|T201|COMP|17197-5|LNC|Cells.CD79b/100 cells|Cells.CD79b/100 cells
C0800325|T201|COMP|17198-3|LNC|Cells.CD8+CD28+/100 cells|Cells.CD8+CD28+/100 cells
C0800326|T201|COMP|17199-1|LNC|Cells.CD80/100 cells|Cells.CD80/100 cells
C0800327|T201|COMP|17200-7|LNC|Cells.CD82/100 cells|Cells.CD82/100 cells
C0800328|T201|COMP|17201-5|LNC|Cells.CD83/100 cells|Cells.CD83/100 cells
C0800329|T201|COMP|17202-3|LNC|Cells.CD85/100 cells|Cells.CD85/100 cells
C0800330|T201|COMP|17203-1|LNC|Cells.CD86/100 cells|Cells.CD86/100 cells
C0800331|T201|COMP|17204-9|LNC|Cells.CD87/100 cells|Cells.CD87/100 cells
C0800332|T201|COMP|17205-6|LNC|Cells.CD88/100 cells|Cells.CD88/100 cells
C0800333|T201|COMP|17206-4|LNC|Cells.CD9/100 cells|Cells.CD9/100 cells
C0800334|T201|COMP|17207-2|LNC|Cells.CD91/100 cells|Cells.CD91/100 cells
C0800335|T201|COMP|17208-0|LNC|Cells.CD93/100 cells|Cells.CD93/100 cells
C0800336|T201|COMP|17209-8|LNC|Cells.CD94/100 cells|Cells.CD94/100 cells
C0800337|T201|COMP|17210-6|LNC|Cells.CD95/100 cells|Cells.CD95/100 cells
C0800338|T201|COMP|17211-4|LNC|Cells.CD96/100 cells|Cells.CD96/100 cells
C0800339|T201|COMP|17212-2|LNC|Cells.CD97/100 cells|Cells.CD97/100 cells
C0800340|T201|COMP|17213-0|LNC|Cells.CD98/100 cells|Cells.CD98/100 cells
C0800341|T201|COMP|17214-8|LNC|Cells.CD99/100 cells|Cells.CD99/100 cells
C0800342|T201|COMP|17215-5|LNC|Lymphocytes.CV/100 lymphocytes|Lymphocytes.CV/100 lymphocytes
C0800343|T201|COMP|17216-3|LNC|Cells.cytoplasmic CD3/100 cells|Cells.cytoplasmic CD3/100 cells
C0800344|T201|COMP|17217-1|LNC|Cells.cytoplasmic CD79/100 cells|Cells.cytoplasmic CD79/100 cells
C0800345|T201|COMP|17218-9|LNC|Cells.cytoplasmic Ig mu/100 cells|Cells.cytoplasmic Ig mu/100 cells
C0800346|T201|COMP|17219-7|LNC|Cells.cytoplasmic Ig/100 cells|Cells.cytoplasmic Ig/100 cells
C0800347|T201|COMP|17220-5|LNC|Cells.FMC7/100 cells|Cells.FMC7/100 cells
C0800349|T201|COMP|17222-1|LNC|Lymphocytes.HLE/100 lymphocytes|Lymphocytes.HLE/100 lymphocytes
C0800351|T201|COMP|17224-7|LNC|Lymphocytes.lambda/100 lymphocytes|Lymphocytes.lambda/100 lymphocytes
C0800352|T201|COMP|17225-4|LNC|Lymphocytes.SmIg/100 lymphocytes|Lymphocytes.SmIg/100 lymphocytes
C0800353|T201|COMP|17226-2|LNC|Cells.SmIg-CD79/100 cells|Cells.SmIg-CD79/100 cells
C0800354|T201|COMP|17227-0|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0800355|T201|COMP|17228-8|LNC|Lymphocytic choriomeningitis virus Ab|Lymphocytic choriomeningitis virus Ab
C0800356|T201|COMP|17229-6|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C0800357|T201|COMP|17230-4|LNC|Lysine|Lysine
C0800358|T201|COMP|17231-2|LNC|Lysosomal enzymes|Lysosomal enzymes
C0800359|T201|COMP|17232-0|LNC|Lysozyme|Lysozyme
C0800360|T201|COMP|17234-6|LNC|Magnesium.plasma/Magnesium.RBC|Magnesium.plasma/Magnesium.RBC
C0800361|T201|COMP|17235-3|LNC|Magnesium|Magnesium
C0800362|T201|COMP|17236-1|LNC|Magnesium|Magnesium
C0800363|T201|COMP|17237-9|LNC|Magnesium|Magnesium
C0800364|T201|COMP|17238-7|LNC|Malignin Ab|Malignin Ab
C0800365|T201|COMP|17241-1|LNC|Prolactin^3H post XXX challenge|Prolactin^3H post XXX challenge
C0800366|T201|COMP|17242-9|LNC|Prolactin^40M post XXX challenge|Prolactin^40M post XXX challenge
C0800367|T201|COMP|17243-7|LNC|Prolactin^pre XXX challenge|Prolactin^pre XXX challenge
C0800368|T201|COMP|17244-5|LNC|Manganese|Manganese
C0800369|T201|COMP|13904-8|LNC|Meclizine|Meclizine
C0800370|T201|COMP|17246-0|LNC|Mefenamate|Mefenamate
C0800371|T201|COMP|17247-8|LNC|Melanin|Melanin
C0800372|T201|COMP|17248-6|LNC|Melanin|Melanin
C0800373|T201|COMP|17249-4|LNC|Menthol|Menthol
C0800374|T201|COMP|17250-2|LNC|Mephobarbital|Mephobarbital
C0800375|T201|COMP|17251-0|LNC|Mepivacaine|Mepivacaine
C0800376|T201|COMP|17252-8|LNC|Mercaptopurine|Mercaptopurine
C0800377|T201|COMP|17253-6|LNC|Mercury|Mercury
C0800378|T201|COMP|17254-4|LNC|Mercury|Mercury
C0800379|T201|COMP|17255-1|LNC|Mercury|Mercury
C0800380|T201|COMP|17256-9|LNC|Mesoridazine|Mesoridazine
C0800381|T201|COMP|17257-7|LNC|Mesothelial cells|Mesothelial cells
C0800382|T201|COMP|17258-5|LNC|Metandienone|Metandienone
C0800383|T201|COMP|17259-3|LNC|Methadone.long acting metabolite|Methadone.long acting metabolite
C0800384|T201|COMP|17260-1|LNC|Methamphetamine|Methamphetamine
C0800385|T201|COMP|17261-9|LNC|Methapyrilene|Methapyrilene
C0800386|T201|COMP|17263-5|LNC|Methemalbumin|Methemalbumin
C0800387|T201|COMP|17264-3|LNC|Methionine|Methionine
C0800388|T201|COMP|17265-0|LNC|Methocarbamol|Methocarbamol
C0800389|T201|COMP|17266-8|LNC|Methotrexate|Methotrexate
C0800390|T201|COMP|17267-6|LNC|Methoxychlor|Methoxychlor
C0800391|T201|COMP|10543-7|LNC|Methsuximide+Normethsuximide|Methsuximide+Normethsuximide
C0800392|T201|COMP|17269-2|LNC|Methyl isobutyl ketone|Methyl isobutyl ketone
C0800393|T201|COMP|17270-0|LNC|Methylacrylate|Methylacrylate
C0800394|T201|COMP|17271-8|LNC|1,1,1-Trichloroethane|1,1,1-Trichloroethane
C0800395|T201|COMP|17272-6|LNC|Methylenedianiline|Methylenedianiline
C0800396|T201|COMP|17273-4|LNC|MethylePHEDrine|MethylePHEDrine
C0800397|T201|COMP|17274-2|LNC|Methylergonovine|Methylergonovine
C0800398|T201|COMP|17275-9|LNC|Methylfentanyl|Methylfentanyl
C0800399|T201|COMP|17276-7|LNC|2-Methylpentane|2-Methylpentane
C0800400|T201|COMP|17277-5|LNC|metOLazone|metOLazone
C0800401|T201|COMP|17278-3|LNC|Miconazole|Miconazole
C0800402|T201|COMP|17279-1|LNC|Bacteria identified|Bacteria identified
C0800403|T201|COMP|17280-9|LNC|Plasmodium sp identified|Plasmodium sp identified
C0800405|T201|COMP|17282-5|LNC|Minoxidil|Minoxidil
C0800406|T201|COMP|17283-3|LNC|Mirtazapine|Mirtazapine
C0800407|T201|COMP|17284-1|LNC|Mitochondria Ab|Mitochondria Ab
C0800408|T201|COMP|17285-8|LNC|Mitochondria Ab|Mitochondria Ab
C0800409|T201|COMP|17286-6|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0800410|T201|COMP|17287-4|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0800411|T201|COMP|17288-2|LNC|Ganglioside GM1 Ab|Ganglioside GM1 Ab
C0800412|T201|COMP|17289-0|LNC|Monosodium glutamate Ab.IgE|Monosodium glutamate Ab.IgE
C0800413|T201|COMP|17290-8|LNC|Morphine|Morphine
C0800415|T201|COMP|17292-4|LNC|Mumps virus Ab|Mumps virus Ab
C0800416|T201|COMP|17293-2|LNC|Mumps virus Ab.IgG+IgM|Mumps virus Ab.IgG+IgM
C0800417|T201|COMP|17294-0|LNC|Mushroom toxins|Mushroom toxins
C0800418|T201|COMP|17296-5|LNC|Mycobacterium tuberculosis complex rRNA|Mycobacterium tuberculosis complex rRNA
C0800421|T201|COMP|17299-9|LNC|Mycoplasma fermentans Ab|Mycoplasma fermentans Ab
C0800422|T201|COMP|17300-5|LNC|Mycoplasma hominis Ab|Mycoplasma hominis Ab
C0800423|T201|COMP|17301-3|LNC|Mycoplasma hominis Ab|Mycoplasma hominis Ab
C0800424|T201|COMP|17302-1|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C0800425|T201|COMP|17303-9|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C0800426|T201|COMP|17304-7|LNC|Mycoplasma pneumoniae Ab.IgG+IgM|Mycoplasma pneumoniae Ab.IgG+IgM
C0800427|T201|COMP|17305-4|LNC|Myelin Ab.IgA|Myelin Ab.IgA
C0800428|T201|COMP|17306-2|LNC|Myelin Ab.IgG|Myelin Ab.IgG
C0800429|T201|COMP|17307-0|LNC|Myelin Ab.IgM|Myelin Ab.IgM
C0800430|T201|COMP|17308-8|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C0800431|T201|COMP|17310-4|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C0800432|T201|COMP|17311-2|LNC|Myelin associated glycoprotein Ab.IgA|Myelin associated glycoprotein Ab.IgA
C0800433|T201|COMP|17312-0|LNC|Myelin associated glycoprotein Ab.IgG|Myelin associated glycoprotein Ab.IgG
C0800434|T201|COMP|17313-8|LNC|Myelin associated glycoprotein Ab.IgG|Myelin associated glycoprotein Ab.IgG
C0800435|T201|COMP|17314-6|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C0800436|T201|COMP|17315-3|LNC|Myelin basic protein Ab|Myelin basic protein Ab
C0800437|T201|COMP|17316-1|LNC|Myeloperoxidase Ab|Myeloperoxidase Ab
C0800438|T201|COMP|17317-9|LNC|N-acetylprocainamide|N-acetylprocainamide
C0800439|T201|COMP|17318-7|LNC|Nalbuphine|Nalbuphine
C0800440|T201|COMP|17319-5|LNC|Nalidixate|Nalidixate
C0800441|T201|COMP|17320-3|LNC|Nefazodone|Nefazodone
C0800442|T201|COMP|17321-1|LNC|Neisseria meningitidis serogroups A+Y Ag|Neisseria meningitidis serogroups A+Y Ag
C0800443|T201|COMP|17322-9|LNC|Neisseria meningitidis Ab|Neisseria meningitidis Ab
C0800444|T201|COMP|17323-7|LNC|Neisseria meningitidis Ag|Neisseria meningitidis Ag
C0800445|T201|COMP|17324-5|LNC|Neisseria meningitidis Ag|Neisseria meningitidis Ag
C0800446|T201|COMP|17325-2|LNC|Neisseria meningitidis serogroups C+w135 Ag|Neisseria meningitidis serogroups C+w135 Ag
C0800447|T201|COMP|17326-0|LNC|Neisseria meningitidis serogroup A Ag|Neisseria meningitidis serogroup A Ag
C0800448|T201|COMP|17327-8|LNC|Neisseria meningitidis serogroup B Ab|Neisseria meningitidis serogroup B Ab
C0800449|T201|COMP|17328-6|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C0800450|T201|COMP|17329-4|LNC|Neisseria meningitidis serogroup C Ag|Neisseria meningitidis serogroup C Ag
C0800451|T201|COMP|17330-2|LNC|Neisseria meningitidis serogroup Y Ag|Neisseria meningitidis serogroup Y Ag
C0800452|T201|COMP|17331-0|LNC|Neisseria meningitidis polyvalent Ab|Neisseria meningitidis polyvalent Ab
C0800453|T201|COMP|17332-8|LNC|Neisseria meningitidis polyvalent Ag|Neisseria meningitidis polyvalent Ag
C0800454|T201|COMP|17333-6|LNC|Neisseria meningitidis serogroup w135 Ag|Neisseria meningitidis serogroup w135 Ag
C0800455|T201|COMP|17334-4|LNC|Neopterin/Creatinine|Neopterin/Creatinine
C0800456|T201|COMP|17335-1|LNC|Neostigmine|Neostigmine
C0800457|T201|COMP|17336-9|LNC|Neuronal Ab|Neuronal Ab
C0800458|T201|COMP|17337-7|LNC|Neuronal Ab|Neuronal Ab
C0800459|T201|COMP|17338-5|LNC|Neuronal Ab|Neuronal Ab
C0800460|T201|COMP|17339-3|LNC|Neuronal Ab|Neuronal Ab
C0800461|T201|COMP|17340-1|LNC|Neuronal Ab.IgG|Neuronal Ab.IgG
C0800462|T201|COMP|17341-9|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C0800463|T201|COMP|17342-7|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C0800464|T201|COMP|17343-5|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C0800465|T201|COMP|17344-3|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C0800466|T201|COMP|5171-4|LNC|Neutrophil Ab|Neutrophil Ab
C0800467|T201|COMP|17346-8|LNC|Neutrophil Ab|Neutrophil Ab
C0800468|T201|COMP|17347-6|LNC|Neutrophil Ab|Neutrophil Ab
C0800469|T201|COMP|17348-4|LNC|Neutrophil Ab.IgA|Neutrophil Ab.IgA
C0800470|T201|COMP|17349-2|LNC|Neutrophil Ab.IgG|Neutrophil Ab.IgG
C0800471|T201|COMP|17350-0|LNC|Neutrophil Ab.IgM|Neutrophil Ab.IgM
C0800472|T201|COMP|17351-8|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C0800473|T201|COMP|17352-6|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C0800474|T201|COMP|17353-4|LNC|Neutrophil cytoplasmic Ab.classic|Neutrophil cytoplasmic Ab.classic
C0800475|T201|COMP|17354-2|LNC|Neutrophil cytoplasmic Ab.IgA|Neutrophil cytoplasmic Ab.IgA
C0800476|T201|COMP|17355-9|LNC|Neutrophil cytoplasmic Ab.IgG|Neutrophil cytoplasmic Ab.IgG
C0800477|T201|COMP|17356-7|LNC|Neutrophil cytoplasmic Ab.IgM|Neutrophil cytoplasmic Ab.IgM
C0800478|T201|COMP|17357-5|LNC|Neutrophil cytoplasmic Ab.perinuclear|Neutrophil cytoplasmic Ab.perinuclear
C0800479|T201|COMP|17358-3|LNC|Neutrophil cytoplasmic Ab.atypical|Neutrophil cytoplasmic Ab.atypical
C0800480|T201|COMP|17359-1|LNC|Neutrophils|Neutrophils
C0800481|T201|COMP|17360-9|LNC|Heptane|Heptane
C0800482|T201|COMP|9475-5|LNC|Hexane|Hexane
C0800483|T201|COMP|17362-5|LNC|Nicotinamide|Nicotinamide
C0800484|T201|COMP|17363-3|LNC|Nitrazepam|Nitrazepam
C0800485|T201|COMP|17364-1|LNC|Nitrophenol|Nitrophenol
C0800486|T201|COMP|17365-8|LNC|Nitroprusside|Nitroprusside
C0800487|T201|COMP|17366-6|LNC|Nizatidine|Nizatidine
C0800488|T201|COMP|17367-4|LNC|Nomifensine|Nomifensine
C0800489|T201|COMP|17368-2|LNC|Norepinephrine^standing|Norepinephrine^standing
C0800490|T201|COMP|17369-0|LNC|Norepinephrine^2nd specimen post XXX challenge|Norepinephrine^2nd specimen post XXX challenge
C0800491|T201|COMP|17370-8|LNC|Norepinephrine^3rd specimen post XXX challenge|Norepinephrine^3rd specimen post XXX challenge
C0800492|T201|COMP|17371-6|LNC|Norepinephrine^4th specimen post XXX challenge|Norepinephrine^4th specimen post XXX challenge
C0800493|T201|COMP|17372-4|LNC|Norepinephrine^5th specimen post XXX challenge|Norepinephrine^5th specimen post XXX challenge
C0800494|T201|COMP|17373-2|LNC|Norepinephrine^6th specimen post XXX challenge|Norepinephrine^6th specimen post XXX challenge
C0800495|T201|COMP|17374-0|LNC|Norepinephrine^7th specimen post XXX challenge|Norepinephrine^7th specimen post XXX challenge
C0800496|T201|COMP|17375-7|LNC|Norflunitrazepam|Norflunitrazepam
C0800497|T201|COMP|17376-5|LNC|Norpropoxyphene|Norpropoxyphene
C0800498|T201|COMP|17377-3|LNC|Norpropoxyphene|Norpropoxyphene
C0800499|T201|COMP|17378-1|LNC|Novobiocin|Novobiocin
C0800500|T201|COMP|17379-9|LNC|Propanol|Propanol
C0800501|T201|COMP|17380-7|LNC|Nuclear Ab.histone reactive|Nuclear Ab.histone reactive
C0800502|T201|COMP|17381-5|LNC|Uroporphyrin|Uroporphyrin
C0800503|T201|COMP|17382-3|LNC|Octadecanoate|Octadecanoate
C0800504|T201|COMP|17384-9|LNC|Opiates|Opiates
C0800505|T201|COMP|17385-6|LNC|Organic acids|Organic acids
C0800506|T201|COMP|17386-4|LNC|Organic acids|Organic acids
C0800507|T201|COMP|17387-2|LNC|Organic acids|Organic acids
C0800508|T201|COMP|17388-0|LNC|Organochlorine pesticides|Organochlorine pesticides
C0800509|T201|COMP|17389-8|LNC|Ornithine|Ornithine
C0800510|T201|COMP|17390-6|LNC|Orphenadrine|Orphenadrine
C0800511|T201|COMP|17391-4|LNC|Orthocresol|Orthocresol
C0800512|T201|COMP|17392-2|LNC|Osmium|Osmium
C0800513|T201|COMP|17393-0|LNC|Ovary Ab|Ovary Ab
C0800514|T201|COMP|17394-8|LNC|Oxychlordane|Oxychlordane
C0800515|T201|COMP|17395-5|LNC|oxyMORphone|oxyMORphone
C0800516|T201|COMP|17396-3|LNC|Oxytetracycline|Oxytetracycline
C0800517|T201|COMP|17397-1|LNC|Oxytriphylline|Oxytriphylline
C0800518|T201|COMP|17398-9|LNC|Human papilloma virus 11 Ag|Human papilloma virus 11 Ag
C0800519|T201|COMP|17399-7|LNC|Human papilloma virus 16 Ag|Human papilloma virus 16 Ag
C0800520|T201|COMP|17400-3|LNC|Human papilloma virus 16+18 Ag|Human papilloma virus 16+18 Ag
C0800521|T201|COMP|17401-1|LNC|Human papilloma virus 18 Ag|Human papilloma virus 18 Ag
C0800522|T201|COMP|17402-9|LNC|Human papilloma virus 31 Ag|Human papilloma virus 31 Ag
C0800523|T201|COMP|17403-7|LNC|Human papilloma virus 31+33+35 Ag|Human papilloma virus 31+33+35 Ag
C0800524|T201|COMP|17404-5|LNC|Human papilloma virus 33 Ag|Human papilloma virus 33 Ag
C0800525|T201|COMP|17405-2|LNC|Human papilloma virus 42 Ag|Human papilloma virus 42 Ag
C0800526|T201|COMP|17406-0|LNC|Human papilloma virus 43 Ag|Human papilloma virus 43 Ag
C0800527|T201|COMP|17407-8|LNC|Human papilloma virus 44 Ag|Human papilloma virus 44 Ag
C0800528|T201|COMP|17408-6|LNC|Human papilloma virus 45 Ag|Human papilloma virus 45 Ag
C0800529|T201|COMP|17409-4|LNC|Human papilloma virus 5 Ag|Human papilloma virus 5 Ag
C0800530|T201|COMP|17410-2|LNC|Human papilloma virus 51 Ag|Human papilloma virus 51 Ag
C0800531|T201|COMP|17411-0|LNC|Human papilloma virus 6 Ag|Human papilloma virus 6 Ag
C0800532|T201|COMP|17412-8|LNC|Human papilloma virus 6+11 Ag|Human papilloma virus 6+11 Ag
C0800533|T201|COMP|17413-6|LNC|Papova virus SV40 Ab|Papova virus SV40 Ab
C0800534|T201|COMP|17414-4|LNC|Parainfluenza virus 1+2+3 Ag|Parainfluenza virus 1+2+3 Ag
C0800535|T201|COMP|17415-1|LNC|Parainfluenza virus A Ab|Parainfluenza virus A Ab
C0800536|T201|COMP|17416-9|LNC|Parakeet droppings Ab|Parakeet droppings Ab
C0800537|T201|COMP|17417-7|LNC|Parakeet droppings Ab.IgG|Parakeet droppings Ab.IgG
C0800538|T201|COMP|17418-5|LNC|Parakeet serum Ab|Parakeet serum Ab
C0800539|T201|COMP|17419-3|LNC|Parathion|Parathion
C0800540|T201|COMP|17420-1|LNC|Parrot droppings Ab|Parrot droppings Ab
C0800541|T201|COMP|17421-9|LNC|Parrot serum Ab|Parrot serum Ab
C0800542|T201|COMP|17422-7|LNC|Parvovirus B19 Ab.IgG+IgM|Parvovirus B19 Ab.IgG+IgM
C0800544|T201|COMP|17424-3|LNC|1,4-Dichlorobenzene|1,4-Dichlorobenzene
C0800545|T201|COMP|17426-8|LNC|Penicillium roqueforti Ab.IgE|Penicillium roqueforti Ab.IgE
C0800546|T201|COMP|17427-6|LNC|Penicillium sp Ab|Penicillium sp Ab
C0800547|T201|COMP|17428-4|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C0800548|T201|COMP|17429-2|LNC|Pentachlorophenol|Pentachlorophenol
C0800549|T201|COMP|17430-0|LNC|Pentane|Pentane
C0800550|T201|COMP|17431-8|LNC|PENTobarbital|PENTobarbital
C0800551|T201|COMP|17432-6|LNC|Tetrachloroethylene|Tetrachloroethylene
C0800553|T201|COMP|17434-2|LNC|Phenazopyridine|Phenazopyridine
C0800554|T201|COMP|17435-9|LNC|Pheniramine|Pheniramine
C0800555|T201|COMP|17436-7|LNC|PHENobarbital|PHENobarbital
C0800556|T201|COMP|17437-5|LNC|Phenolphthalein|Phenolphthalein
C0800557|T201|COMP|17438-3|LNC|Phenolphthalein|Phenolphthalein
C0800558|T201|COMP|17439-1|LNC|Phenols|Phenols
C0800559|T201|COMP|17440-9|LNC|Phenothiazines|Phenothiazines
C0800560|T201|COMP|17441-7|LNC|Phenothiazines|Phenothiazines
C0800561|T201|COMP|17442-5|LNC|Phenylephrine|Phenylephrine
C0800562|T201|COMP|17443-3|LNC|Phenylpropanolamine|Phenylpropanolamine
C0800563|T201|COMP|17444-1|LNC|Phenytoin|Phenytoin
C0800564|T201|COMP|17445-8|LNC|Phoma herbarum Ab.IgG|Phoma herbarum Ab.IgG
C0800565|T201|COMP|17446-6|LNC|Phoma sp Ab.IgE|Phoma sp Ab.IgE
C0800566|T201|COMP|17447-4|LNC|Phosphate|Phosphate
C0800567|T201|COMP|17448-2|LNC|Phosphatidylethanolamine Ab.IgA|Phosphatidylethanolamine Ab.IgA
C0800568|T201|COMP|17449-0|LNC|Phosphatidylethanolamine Ab.IgG|Phosphatidylethanolamine Ab.IgG
C0800569|T201|COMP|17450-8|LNC|Phosphatidylethanolamine Ab.IgM|Phosphatidylethanolamine Ab.IgM
C0800570|T201|COMP|17451-6|LNC|Phosphatidylglycerol Ab.IgA|Phosphatidylglycerol Ab.IgA
C0800571|T201|COMP|17452-4|LNC|Phosphatidylglycerol Ab.IgG|Phosphatidylglycerol Ab.IgG
C0800572|T201|COMP|17453-2|LNC|Phosphatidylglycerol Ab.IgM|Phosphatidylglycerol Ab.IgM
C0800573|T201|COMP|17454-0|LNC|Phosphatidylinositol Ab.IgA|Phosphatidylinositol Ab.IgA
C0800574|T201|COMP|17455-7|LNC|Phosphatidylinositol Ab.IgG|Phosphatidylinositol Ab.IgG
C0800575|T201|COMP|17456-5|LNC|Phosphatidylinositol Ab.IgM|Phosphatidylinositol Ab.IgM
C0800576|T201|COMP|17457-3|LNC|Phosphoethanolamine|Phosphoethanolamine
C0800577|T201|COMP|17458-1|LNC|Phosphoethanolamine|Phosphoethanolamine
C0800578|T201|COMP|17459-9|LNC|Phospholipid Ab.IgA|Phospholipid Ab.IgA
C0800579|T201|COMP|17460-7|LNC|Phosphoserine|Phosphoserine
C0800580|T201|COMP|17461-5|LNC|Phosphoserine|Phosphoserine
C0800581|T201|COMP|17462-3|LNC|Picloram|Picloram
C0800582|T201|COMP|17463-1|LNC|Pigeon droppings Ab|Pigeon droppings Ab
C0800583|T201|COMP|17464-9|LNC|Pigeon feather Ab.IgE|Pigeon feather Ab.IgE
C0800584|T201|COMP|17465-6|LNC|Pigeon serum Ab.IgE|Pigeon serum Ab.IgE
C0800585|T201|COMP|17466-4|LNC|Plasminogen activator inhibitor 1 Ag|Plasminogen activator inhibitor 1 Ag
C0800586|T201|COMP|17467-2|LNC|Plasminogen activator inhibitor 2 Ag|Plasminogen activator inhibitor 2 Ag
C0800587|T201|COMP|17468-0|LNC|Plutonium|Plutonium
C0800588|T201|COMP|17469-8|LNC|PM-1 Ab|PM-1 Ab
C0800589|T201|COMP|17470-6|LNC|PM-1 Ab|PM-1 Ab
C0800590|T201|COMP|17471-4|LNC|PM-1 Ab|PM-1 Ab
C0800591|T201|COMP|17472-2|LNC|Polybrominated biphenyl|Polybrominated biphenyl
C0800592|T201|COMP|17473-0|LNC|Polymyxin B|Polymyxin B
C0800593|T201|COMP|17474-8|LNC|Porphobilinogen|Porphobilinogen
C0800594|T201|COMP|17475-5|LNC|Porphyrins|Porphyrins
C0800595|T201|COMP|17476-3|LNC|Porphyrins|Porphyrins
C0800596|T201|COMP|17477-1|LNC|Porphyrins|Porphyrins
C0800597|T201|COMP|17478-9|LNC|Porphyrins|Porphyrins
C0800598|T201|COMP|17479-7|LNC|Prazepam|Prazepam
C0800599|T201|COMP|17480-5|LNC|Pregnenolone|Pregnenolone
C0800600|T201|COMP|17481-3|LNC|Probenecid|Probenecid
C0800601|T201|COMP|17482-1|LNC|Procainamide|Procainamide
C0800602|T201|COMP|17483-9|LNC|Progesterone|Progesterone
C0800603|T201|COMP|17484-7|LNC|Progesterone^1.5H post XXX challenge|Progesterone^1.5H post XXX challenge
C0800604|T201|COMP|17485-4|LNC|Progesterone^15M post XXX challenge|Progesterone^15M post XXX challenge
C0800605|T201|COMP|17486-2|LNC|Progesterone^2H post XXX challenge|Progesterone^2H post XXX challenge
C0800606|T201|COMP|17487-0|LNC|Progesterone^45M post XXX challenge|Progesterone^45M post XXX challenge
C0800607|T201|COMP|17488-8|LNC|Progesterone^7th specimen post XXX challenge|Progesterone^7th specimen post XXX challenge
C0800608|T201|COMP|17489-6|LNC|Progesterone^8th specimen post XXX challenge|Progesterone^8th specimen post XXX challenge
C0800609|T201|COMP|17490-4|LNC|Progesterone^9th specimen post XXX challenge|Progesterone^9th specimen post XXX challenge
C0800610|T201|COMP|17491-2|LNC|Proinsulin^baseline|Proinsulin^baseline
C0800611|T201|COMP|17492-0|LNC|Proline|Proline
C0800612|T201|COMP|17493-8|LNC|Prostaglandin E|Prostaglandin E
C0800613|T201|COMP|17494-6|LNC|Prostaglandin F2 alpha|Prostaglandin F2 alpha
C0800614|T201|COMP|17495-3|LNC|Prostaglandins|Prostaglandins
C0800615|T201|COMP|17496-1|LNC|Alpha 1 globulin|Alpha 1 globulin
C0800616|T201|COMP|17497-9|LNC|Alpha 2 globulin|Alpha 2 globulin
C0800617|T201|COMP|17498-7|LNC|Beta globulin|Beta globulin
C0800618|T201|COMP|17499-5|LNC|Gamma globulin|Gamma globulin
C0800619|T201|COMP|17501-8|LNC|Protoporphyrin|Protoporphyrin
C0800620|T201|COMP|17502-6|LNC|Pseudomonas aeruginosa Ab|Pseudomonas aeruginosa Ab
C0800621|T201|COMP|17504-2|LNC|Psilocybin|Psilocybin
C0800622|T201|COMP|17505-9|LNC|Psilocybin/Psilocin|Psilocybin/Psilocin
C0800623|T201|COMP|17506-7|LNC|Quinacrine|Quinacrine
C0800624|T201|COMP|17507-5|LNC|quiNIDine|quiNIDine
C0800625|T201|COMP|17508-3|LNC|quiNINE|quiNINE
C0800626|T201|COMP|17509-1|LNC|Ragweed marsh Ab.IgE|Ragweed marsh Ab.IgE
C0800627|T201|COMP|17510-9|LNC|Raisin Ab.IgE|Raisin Ab.IgE
C0800628|T201|COMP|17511-7|LNC|Red dye Ab.IgE|Red dye Ab.IgE
C0800629|T201|COMP|17512-5|LNC|Redfish Ab.IgE|Redfish Ab.IgE
C0800630|T201|COMP|17513-3|LNC|Renin^5H post XXX challenge|Renin^5H post XXX challenge
C0800631|T201|COMP|17514-1|LNC|Renin^9th specimen post XXX challenge|Renin^9th specimen post XXX challenge
C0800632|T201|COMP|17515-8|LNC|Renin^baseline|Renin^baseline
C0800633|T201|COMP|17516-6|LNC|Renin^supine|Renin^supine
C0800634|T201|COMP|17517-4|LNC|Respiratory syncytial virus Ab.IgG|Respiratory syncytial virus Ab.IgG
C0800635|T201|COMP|17518-2|LNC|Respiratory syncytial virus Ab.IgG|Respiratory syncytial virus Ab.IgG
C0800636|T201|COMP|17519-0|LNC|Respiratory syncytial virus Ab.IgM|Respiratory syncytial virus Ab.IgM
C0800637|T201|COMP|17520-8|LNC|Respiratory syncytial virus identified|Respiratory syncytial virus identified
C0800638|T201|COMP|17521-6|LNC|Reticulin Ab|Reticulin Ab
C0800639|T201|COMP|17522-4|LNC|Reticulin Ab.IgA|Reticulin Ab.IgA
C0800640|T201|COMP|17523-2|LNC|Reticulin Ab.IgG|Reticulin Ab.IgG
C0800641|T201|COMP|17524-0|LNC|Reticulin Ab.IgG|Reticulin Ab.IgG
C0800642|T201|COMP|17525-7|LNC|Retinoate esters|Retinoate esters
C0800643|T201|COMP|17526-5|LNC|Retinyl esters|Retinyl esters
C0800644|T201|COMP|17527-3|LNC|Retinol.free|Retinol.free
C0800645|T201|COMP|17528-1|LNC|Retinol^3H post dose|Retinol^3H post dose
C0800646|T201|COMP|17529-9|LNC|Retinol^6H post dose|Retinol^6H post dose
C0800647|T201|COMP|17530-7|LNC|Retrovirus identified|Retrovirus identified
C0800648|T201|COMP|17531-5|LNC|Rh|Rh
C0800649|T201|COMP|17532-3|LNC|Rheumatoid arthritis nuclear Ab|Rheumatoid arthritis nuclear Ab
C0800650|T201|COMP|17533-1|LNC|Rheumatoid arthritis nuclear Ab|Rheumatoid arthritis nuclear Ab
C0800651|T201|COMP|17534-9|LNC|Rheumatoid factor|Rheumatoid factor
C0800652|T201|COMP|17535-6|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0800653|T201|COMP|17536-4|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0800654|T201|COMP|17537-2|LNC|Rickettsia spotted fever group RNA|Rickettsia spotted fever group RNA
C0800655|T201|COMP|17538-0|LNC|Rickettsia spotted fever group RNA|Rickettsia spotted fever group RNA
C0800656|T201|COMP|17539-8|LNC|Rickettsia typhi Ab|Rickettsia typhi Ab
C0800657|T201|COMP|17540-6|LNC|Rickettsia typhi Ab.IgA|Rickettsia typhi Ab.IgA
C0800658|T201|COMP|17541-4|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C0800659|T201|COMP|17544-8|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C0800660|T201|COMP|17545-5|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C0800661|T201|COMP|17546-3|LNC|Bartonella quintana rRNA|Bartonella quintana rRNA
C0800662|T201|COMP|17547-1|LNC|Rotavirus Ag|Rotavirus Ag
C0800663|T201|COMP|17548-9|LNC|Rotavirus RNA|Rotavirus RNA
C0800664|T201|COMP|17549-7|LNC|Rubella virus Ab|Rubella virus Ab
C0800665|T201|COMP|17550-5|LNC|Rubella virus Ab|Rubella virus Ab
C0800666|T201|COMP|17551-3|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0800667|T201|COMP|17552-1|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C0800668|T201|COMP|17553-9|LNC|Measles virus Ab|Measles virus Ab
C0800669|T201|COMP|17554-7|LNC|Measles virus Ab.IgA|Measles virus Ab.IgA
C0800670|T201|COMP|17555-4|LNC|Measles virus Ab^1st specimen|Measles virus Ab^1st specimen
C0800671|T201|COMP|17556-2|LNC|Measles virus Ab^2nd specimen|Measles virus Ab^2nd specimen
C0800672|T201|COMP|17557-0|LNC|Saccharomonospora viridis Ab.IgG|Saccharomonospora viridis Ab.IgG
C0800673|T201|COMP|17558-8|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0800674|T201|COMP|17559-6|LNC|Salicylates|Salicylates
C0800675|T201|COMP|17560-4|LNC|Salicylates|Salicylates
C0800676|T201|COMP|17561-2|LNC|Salmo salar roe Ab.IgE|Salmo salar roe Ab.IgE
C0800677|T201|COMP|17562-0|LNC|Salmonella sp Ab|Salmonella sp Ab
C0800679|T201|COMP|17564-6|LNC|Salmonella typhi O D Ab|Salmonella typhi O D Ab
C0800680|T201|COMP|17565-3|LNC|Salmonella typhi H D Ab|Salmonella typhi H D Ab
C0800681|T201|COMP|17566-1|LNC|Salmonella typhi O Ab|Salmonella typhi O Ab
C0800682|T201|COMP|17567-9|LNC|Sasapyrine|Sasapyrine
C0800683|T201|COMP|17568-7|LNC|Sarcosine|Sarcosine
C0800684|T201|COMP|17569-5|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C0800685|T201|COMP|17570-3|LNC|SCL-70 extractable nuclear Ab.IgG|SCL-70 extractable nuclear Ab.IgG
C0800686|T201|COMP|17571-1|LNC|Scopolamine|Scopolamine
C0800687|T201|COMP|17572-9|LNC|2-Butanol|2-Butanol
C0800688|T201|COMP|17573-7|LNC|Secobarbital|Secobarbital
C0800689|T201|COMP|17574-5|LNC|Selenium|Selenium
C0800690|T201|COMP|17575-2|LNC|Serine|Serine
C0800691|T201|COMP|17576-0|LNC|Shigella sp identified|Shigella sp identified
C0800692|T201|COMP|17577-8|LNC|Ganglioside GQ1a Ab.IgM|Ganglioside GQ1a Ab.IgM
C0800693|T201|COMP|17578-6|LNC|Ganglioside GQ1b Ab|Ganglioside GQ1b Ab
C0800694|T201|COMP|17579-4|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C0800695|T201|COMP|17580-2|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C0800696|T201|COMP|17581-0|LNC|Ganglioside GQ1b Ab.IgM|Ganglioside GQ1b Ab.IgM
C0800697|T201|COMP|17582-8|LNC|Silver|Silver
C0800698|T201|COMP|17583-6|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C0800699|T201|COMP|17584-4|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C0800700|T201|COMP|17585-1|LNC|Sjogrens syndrome-A extractable nuclear Ab.IgG|Sjogrens syndrome-A extractable nuclear Ab.IgG
C0800701|T201|COMP|17586-9|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C0800702|T201|COMP|17587-7|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C0800703|T201|COMP|17588-5|LNC|Sjogrens syndrome-B extractable nuclear Ab.IgG|Sjogrens syndrome-B extractable nuclear Ab.IgG
C0800704|T201|COMP|17589-3|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0800705|T201|COMP|17590-1|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0800706|T201|COMP|17591-9|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0800707|T201|COMP|17592-7|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0800708|T201|COMP|17593-5|LNC|Smooth muscle Ab|Smooth muscle Ab
C0800709|T201|COMP|17594-3|LNC|Somatotropin^1.5H post XXX challenge|Somatotropin^1.5H post XXX challenge
C0800710|T201|COMP|17595-0|LNC|Somatotropin^1H post XXX challenge|Somatotropin^1H post XXX challenge
C0800711|T201|COMP|17597-6|LNC|Somatotropin^52H post XXX challenge|Somatotropin^52H post XXX challenge
C0800712|T201|COMP|17598-4|LNC|Specific gravity|Specific gravity
C0800713|T201|COMP|17599-2|LNC|Specimen volume|Specimen volume
C0800714|T201|COMP|17600-8|LNC|Specimen volume|Specimen volume
C0800715|T201|COMP|17601-6|LNC|Specimen volume|Specimen volume
C0800716|T201|COMP|17602-4|LNC|Specimen volume|Specimen volume
C0800717|T201|COMP|17603-2|LNC|Specimen volume|Specimen volume
C0800718|T201|COMP|17604-0|LNC|Specimen volume|Specimen volume
C0800719|T201|COMP|17605-7|LNC|Specimen volume|Specimen volume
C0800720|T201|COMP|17606-5|LNC|Specimen volume|Specimen volume
C0800721|T201|COMP|17607-3|LNC|Specimen volume|Specimen volume
C0800722|T201|COMP|17608-1|LNC|Specimen weight|Specimen weight
C0800723|T201|COMP|17609-9|LNC|Specimen weight|Specimen weight
C0800724|T201|COMP|17610-7|LNC|Spermatozoa.motile^30M post collection|Spermatozoa.motile^30M post collection
C0800725|T201|COMP|17611-5|LNC|Stimulants|Stimulants
C0800726|T201|COMP|13139-1|LNC|Streptococcus pneumoniae 1 Ab^1st specimen|Streptococcus pneumoniae 1 Ab^1st specimen
C0800727|T201|COMP|13140-9|LNC|Streptococcus pneumoniae 1 Ab^2nd specimen|Streptococcus pneumoniae 1 Ab^2nd specimen
C0800728|T201|COMP|17614-9|LNC|Streptococcus pneumoniae 12 Ab|Streptococcus pneumoniae 12 Ab
C0800729|T201|COMP|13153-2|LNC|Streptococcus pneumoniae 12 Ab^1st specimen|Streptococcus pneumoniae 12 Ab^1st specimen
C0800731|T201|COMP|17617-2|LNC|Streptococcus pneumoniae 14 Ab^1st specimen|Streptococcus pneumoniae 14 Ab^1st specimen
C0800732|T201|COMP|17618-0|LNC|Streptococcus pneumoniae 14 Ab^2nd specimen|Streptococcus pneumoniae 14 Ab^2nd specimen
C0800736|T201|COMP|17622-2|LNC|Streptococcus pneumoniae 18 Ab^1st specimen|Streptococcus pneumoniae 18 Ab^1st specimen
C0800737|T201|COMP|13160-7|LNC|Streptococcus pneumoniae 19 Ab^2nd specimen|Streptococcus pneumoniae 19 Ab^2nd specimen
C0800738|T201|COMP|13161-5|LNC|Streptococcus pneumoniae 23 Ab^1st specimen|Streptococcus pneumoniae 23 Ab^1st specimen
C0800739|T201|COMP|13162-3|LNC|Streptococcus pneumoniae 23 Ab^2nd specimen|Streptococcus pneumoniae 23 Ab^2nd specimen
C0800740|T201|COMP|13141-7|LNC|Streptococcus pneumoniae 3 Ab^1st specimen|Streptococcus pneumoniae 3 Ab^1st specimen
C0800741|T201|COMP|17627-1|LNC|Streptococcus pneumoniae 3 Ab^1st specimen|Streptococcus pneumoniae 3 Ab^1st specimen
C0800742|T201|COMP|13142-5|LNC|Streptococcus pneumoniae 3 Ab^2nd specimen|Streptococcus pneumoniae 3 Ab^2nd specimen
C0800743|T201|COMP|17629-7|LNC|Streptococcus pneumoniae 3 Ab^2nd specimen|Streptococcus pneumoniae 3 Ab^2nd specimen
C0800745|T201|COMP|17631-3|LNC|Streptococcus pneumoniae 36a+6b Ab.IgG|Streptococcus pneumoniae 36a+6b Ab.IgG
C0800746|T201|COMP|17632-1|LNC|Streptococcus pneumoniae 4 Ab.IgG|Streptococcus pneumoniae 4 Ab.IgG
C0800747|T201|COMP|13143-3|LNC|Streptococcus pneumoniae 4 Ab^1st specimen|Streptococcus pneumoniae 4 Ab^1st specimen
C0800748|T201|COMP|13144-1|LNC|Streptococcus pneumoniae 4 Ab^2nd specimen|Streptococcus pneumoniae 4 Ab^2nd specimen
C0800755|T201|COMP|17641-2|LNC|Streptococcus pneumoniae 8 Ab|Streptococcus pneumoniae 8 Ab
C0800756|T201|COMP|17642-0|LNC|Streptococcus pneumoniae 8 Ab|Streptococcus pneumoniae 8 Ab
C0800757|T201|COMP|17643-8|LNC|Streptococcus pneumoniae 9 Ab|Streptococcus pneumoniae 9 Ab
C0800759|T201|COMP|17645-3|LNC|Streptococcus pneumoniae 9 Ab^1st specimen|Streptococcus pneumoniae 9 Ab^1st specimen
C0800760|T201|COMP|17646-1|LNC|Streptococcus pneumoniae 9 Ab^2nd specimen|Streptococcus pneumoniae 9 Ab^2nd specimen
C0800761|T201|COMP|17647-9|LNC|Streptococcus pneumoniae Ab|Streptococcus pneumoniae Ab
C0800762|T201|COMP|17648-7|LNC|Streptococcus pneumoniae Ab|Streptococcus pneumoniae Ab
C0800764|T201|COMP|17650-3|LNC|Streptococcus pneumoniae Ab.IgG^1st specimen|Streptococcus pneumoniae Ab.IgG^1st specimen
C0800765|T201|COMP|17651-1|LNC|Streptococcus pneumoniae Ab.IgG^2nd specimen|Streptococcus pneumoniae Ab.IgG^2nd specimen
C0800766|T201|COMP|17652-9|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C0800767|T201|COMP|17653-7|LNC|Streptococcus pneumoniae group A Ag|Streptococcus pneumoniae group A Ag
C0800768|T201|COMP|17654-5|LNC|Streptococcus pneumoniae group B Ab|Streptococcus pneumoniae group B Ab
C0800769|T201|COMP|17655-2|LNC|Streptococcus pneumoniae group B Ag|Streptococcus pneumoniae group B Ag
C0800770|T201|COMP|17656-0|LNC|Streptococcus pyogenes|Streptococcus pyogenes
C0800771|T201|COMP|17657-8|LNC|Streptolysin O Ab|Streptolysin O Ab
C0800772|T201|COMP|17658-6|LNC|Strontium/Creatinine|Strontium/Creatinine
C0800773|T201|COMP|17659-4|LNC|Strychnine|Strychnine
C0800774|T201|COMP|17660-2|LNC|Strychnine|Strychnine
C0800775|T201|COMP|17661-0|LNC|Succinylcholine|Succinylcholine
C0800776|T201|COMP|17662-8|LNC|Succinylpurines|Succinylpurines
C0800777|T201|COMP|17663-6|LNC|sulfADIAZINE Ab.IgE|sulfADIAZINE Ab.IgE
C0800778|T201|COMP|17664-4|LNC|Sulfalazine Ab.IgE|Sulfalazine Ab.IgE
C0800779|T201|COMP|17665-1|LNC|Sulfamedraxozole Ab.IgE|Sulfamedraxozole Ab.IgE
C0800780|T201|COMP|17666-9|LNC|Sulfate|Sulfate
C0800781|T201|COMP|17667-7|LNC|Sulfate.organic/Sulfate.total|Sulfate.organic/Sulfate.total
C0800782|T201|COMP|17668-5|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C0800783|T201|COMP|17669-3|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C0800784|T201|COMP|17670-1|LNC|Sulfatide Ab.IgM|Sulfatide Ab.IgM
C0800785|T201|COMP|17671-9|LNC|Sulfatide Ab.IgM|Sulfatide Ab.IgM
C0800786|T201|COMP|17672-7|LNC|Sulfide|Sulfide
C0800787|T201|COMP|17673-5|LNC|sulfiSOXAZOLE Ab.IgE|sulfiSOXAZOLE Ab.IgE
C0800788|T201|COMP|17674-3|LNC|Sulfonamide|Sulfonamide
C0800789|T201|COMP|17675-0|LNC|Sulfonamide|Sulfonamide
C0800790|T201|COMP|17676-8|LNC|Sulindac sulfide metabolite|Sulindac sulfide metabolite
C0800791|T201|COMP|17677-6|LNC|Helianthus annuus Ab.IgE|Helianthus annuus Ab.IgE
C0800792|T201|COMP|17678-4|LNC|Taurine|Taurine
C0800793|T201|COMP|17679-2|LNC|Taurine|Taurine
C0800794|T201|COMP|17681-8|LNC|Tellurium|Tellurium
C0800795|T201|COMP|17682-6|LNC|Terpineol|Terpineol
C0800796|T201|COMP|17683-4|LNC|2-Methyl-2-Propanol|2-Methyl-2-Propanol
C0800797|T201|COMP|17685-9|LNC|Testosterone.free|Testosterone.free
C0800798|T201|COMP|17686-7|LNC|Testosterone.weakly bound|Testosterone.weakly bound
C0800799|T201|COMP|17687-5|LNC|Testosterone/Epitestosterone|Testosterone/Epitestosterone
C0800800|T201|COMP|17688-3|LNC|Testosterone^1.5H post XXX challenge|Testosterone^1.5H post XXX challenge
C0800801|T201|COMP|17689-1|LNC|Testosterone^15M post XXX challenge|Testosterone^15M post XXX challenge
C0800802|T201|COMP|17690-9|LNC|Testosterone^2H post XXX challenge|Testosterone^2H post XXX challenge
C0800803|T201|COMP|17691-7|LNC|Testosterone^30M post XXX challenge|Testosterone^30M post XXX challenge
C0800804|T201|COMP|17692-5|LNC|Testosterone^45M post XXX challenge|Testosterone^45M post XXX challenge
C0800805|T201|COMP|17693-3|LNC|Testosterone^4D post XXX challenge|Testosterone^4D post XXX challenge
C0800807|T201|COMP|17695-8|LNC|Tetrachlorodiphenylethane|Tetrachlorodiphenylethane
C0800808|T201|COMP|17696-6|LNC|Tetrachlorodiphenylethane|Tetrachlorodiphenylethane
C0800809|T201|COMP|17697-4|LNC|Tetrachloroethane|Tetrachloroethane
C0800810|T201|COMP|17698-2|LNC|Tetraethyl lead|Tetraethyl lead
C0800811|T201|COMP|17699-0|LNC|Thebaine|Thebaine
C0800812|T201|COMP|17700-6|LNC|Theophylline|Theophylline
C0800813|T201|COMP|17701-4|LNC|Thiazides|Thiazides
C0800814|T201|COMP|17703-0|LNC|Thorium|Thorium
C0800815|T201|COMP|17704-8|LNC|Threonine|Threonine
C0800816|T201|COMP|17705-5|LNC|Thyroglobulin Ab.IgM|Thyroglobulin Ab.IgM
C0800817|T201|COMP|17706-3|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C0800818|T201|COMP|17707-1|LNC|Thyroperoxidase Ab.IgM|Thyroperoxidase Ab.IgM
C0800819|T201|COMP|17708-9|LNC|Thyroid stimulating immunoglobulins|Thyroid stimulating immunoglobulins
C0800820|T201|COMP|17709-7|LNC|Ticlopidine|Ticlopidine
C0800821|T201|COMP|17710-5|LNC|Tin/Creatinine|Tin/Creatinine
C0800822|T201|COMP|17712-1|LNC|Toluene diisocyanate|Toluene diisocyanate
C0800823|T201|COMP|17713-9|LNC|Topiramate|Topiramate
C0800824|T201|COMP|17714-7|LNC|Toxaphene|Toxaphene
C0800825|T201|COMP|17715-4|LNC|Toxocara canis Ab|Toxocara canis Ab
C0800826|T201|COMP|17716-2|LNC|Toxoplasma gondii Ab.IgE|Toxoplasma gondii Ab.IgE
C0800827|T201|COMP|17717-0|LNC|Toxoplasma gondii Ab.IgG+IgM|Toxoplasma gondii Ab.IgG+IgM
C0800828|T201|COMP|17718-8|LNC|traMADol|traMADol
C0800829|T201|COMP|17719-6|LNC|traMADol|traMADol
C0800830|T201|COMP|17720-4|LNC|Trans nonachlor|Trans nonachlor
C0800831|T201|COMP|17721-2|LNC|Trans nonachlor|Trans nonachlor
C0800832|T201|COMP|17723-8|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0800833|T201|COMP|17724-6|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0800834|T201|COMP|17725-3|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0800835|T201|COMP|17726-1|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C0800836|T201|COMP|17727-9|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C0800837|T201|COMP|17728-7|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C0800838|T201|COMP|17729-5|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C0800839|T201|COMP|17730-3|LNC|Triamterene|Triamterene
C0800840|T201|COMP|17732-9|LNC|Trichinella spiralis Ab|Trichinella spiralis Ab
C0800841|T201|COMP|17733-7|LNC|Trichinella spiralis Ab.IgA|Trichinella spiralis Ab.IgA
C0800842|T201|COMP|17734-5|LNC|Trichinella spiralis Ab.IgG|Trichinella spiralis Ab.IgG
C0800843|T201|COMP|17735-2|LNC|Trichinella spiralis Ab.IgM|Trichinella spiralis Ab.IgM
C0800844|T201|COMP|17736-0|LNC|Trichloroacetate|Trichloroacetate
C0800845|T201|COMP|17737-8|LNC|Trichloroethane|Trichloroethane
C0800847|T201|COMP|17739-4|LNC|Chloral hydrate|Chloral hydrate
C0800848|T201|COMP|17740-2|LNC|Trichlorophenoxyacetate|Trichlorophenoxyacetate
C0800849|T201|COMP|17741-0|LNC|Trichlorophenoxyacetate|Trichlorophenoxyacetate
C0800850|T201|COMP|17742-8|LNC|Trichlorothiazide|Trichlorothiazide
C0800852|T201|COMP|17744-4|LNC|Trimellitic anhydride Ab.IgG|Trimellitic anhydride Ab.IgG
C0800853|T201|COMP|17745-1|LNC|Trimellitic anhydride Ab.IgM|Trimellitic anhydride Ab.IgM
C0800854|T201|COMP|17746-9|LNC|Trimeprazine|Trimeprazine
C0800855|T201|COMP|17747-7|LNC|Trimethoprim|Trimethoprim
C0800856|T201|COMP|17748-5|LNC|Trimethylamine|Trimethylamine
C0800857|T201|COMP|17749-3|LNC|Tromethamine|Tromethamine
C0800858|T201|COMP|17750-1|LNC|Trypsinogen|Trypsinogen
C0800859|T201|COMP|17751-9|LNC|Tryptamine|Tryptamine
C0800860|T201|COMP|17752-7|LNC|Tryptophan|Tryptophan
C0800861|T201|COMP|17753-5|LNC|Tungsten|Tungsten
C0800862|T201|COMP|17754-3|LNC|Tyrosine|Tyrosine
C0800863|T201|COMP|17755-0|LNC|Urate|Urate
C0800864|T201|COMP|17756-8|LNC|Urate|Urate
C0800865|T201|COMP|17757-6|LNC|Urea nitrogen|Urea nitrogen
C0800866|T201|COMP|17758-4|LNC|Urea nitrogen|Urea nitrogen
C0800867|T201|COMP|17759-2|LNC|Urea nitrogen^post dialysis|Urea nitrogen^post dialysis
C0800868|T201|COMP|17760-0|LNC|Urea nitrogen^pre dialysis|Urea nitrogen^pre dialysis
C0800869|T201|COMP|17761-8|LNC|Urobilinogen|Urobilinogen
C0800870|T201|COMP|17762-6|LNC|Valproate|Valproate
C0800871|T201|COMP|17763-4|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0800872|T201|COMP|17764-2|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0800873|T201|COMP|17765-9|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0800874|T201|COMP|17766-7|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0800875|T201|COMP|17767-5|LNC|Verapamil|Verapamil
C0800876|T201|COMP|17768-3|LNC|Vinyl chloride|Vinyl chloride
C0800877|T201|COMP|17769-1|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0800879|T201|COMP|17771-7|LNC|Whitefish roe Ab.IgE|Whitefish roe Ab.IgE
C0800880|T201|COMP|17772-5|LNC|Dimethylbenzene|Dimethylbenzene
C0800881|T201|COMP|17773-3|LNC|Yeast|Yeast
C0800882|T201|COMP|17774-1|LNC|Yellow dye Ab.IgE|Yellow dye Ab.IgE
C0800883|T201|COMP|17775-8|LNC|Yersinia sp Ab.IgA|Yersinia sp Ab.IgA
C0800884|T201|COMP|17776-6|LNC|Yersinia sp Ab.IgG|Yersinia sp Ab.IgG
C0800885|T201|COMP|17777-4|LNC|Yersinia sp Ab.IgM|Yersinia sp Ab.IgM
C0800886|T201|COMP|17778-2|LNC|Zinc|Zinc
C0800887|T201|COMP|17780-8|LNC|Helicobacter pylori Ag|Helicobacter pylori Ag
C0800888|T201|COMP|17781-6|LNC|21-Hydroxylase Ab|21-Hydroxylase Ab
C0800889|T201|COMP|17782-4|LNC|Lipoprotein.beta.subparticle|Lipoprotein.beta.subparticle
C0800890|T201|COMP|17783-2|LNC|Hemosiderin|Hemosiderin
C0800891|T201|COMP|17784-0|LNC|Parasite identified|Parasite identified
C0800893|T201|COMP|17786-5|LNC|Thyrotropin^post dose TRH|Thyrotropin^post dose TRH
C0800895|T201|COMP|17788-1|LNC|Large unstained cells/100 leukocytes|Large unstained cells/100 leukocytes
C0800896|T201|COMP|17789-9|LNC|Large unstained cells|Large unstained cells
C0800897|T201|COMP|17790-7|LNC|Leukocytes.left shift|Leukocytes.left shift
C0800898|T201|COMP|17791-5|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C0800899|T201|COMP|17792-3|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C0800900|T201|COMP|17793-1|LNC|Immunoglobulin light chains|Immunoglobulin light chains
C0800901|T201|COMP|17794-9|LNC|Osmolality|Osmolality
C0800902|T201|COMP|17795-6|LNC|Potassium|Potassium
C0800903|T201|COMP|17796-4|LNC|Sodium|Sodium
C0800904|T201|COMP|17797-2|LNC|Thyroid colloidal Ab|Thyroid colloidal Ab
C0800905|T201|COMP|17798-0|LNC|Amikacin|Amikacin
C0800906|T201|COMP|17799-8|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C0800907|T201|COMP|17800-4|LNC|Myelocytes/100 leukocytes|Myelocytes/100 leukocytes
C0800908|T201|COMP|17801-2|LNC|Metamyelocytes/100 leukocytes|Metamyelocytes/100 leukocytes
C0800909|T201|COMP|17802-0|LNC|Prolymphocytes/100 leukocytes|Prolymphocytes/100 leukocytes
C0800910|T201|COMP|17803-8|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C0800911|T201|COMP|17804-6|LNC|Promonocytes/100 leukocytes|Promonocytes/100 leukocytes
C0800912|T201|COMP|17805-3|LNC|Procainamide|Procainamide
C0800913|T201|COMP|17806-1|LNC|N-acetylprocainamide|N-acetylprocainamide
C0800914|T201|COMP|17807-9|LNC|cycloSPORINE|cycloSPORINE
C0800915|T201|COMP|17808-7|LNC|Tobramycin|Tobramycin
C0800916|T201|COMP|17809-5|LNC|Hematocrit|Hematocrit
C0800917|T201|COMP|17810-3|LNC|Prealbumin/Protein.total|Prealbumin/Protein.total
C0800918|T201|COMP|17811-1|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0800919|T201|COMP|17812-9|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0800920|T201|COMP|17813-7|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0800921|T201|COMP|17814-5|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0800922|T201|COMP|17815-2|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C0800923|T201|COMP|17816-0|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C0800924|T201|COMP|17817-8|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0800925|T201|COMP|17818-6|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0800926|T201|COMP|17819-4|LNC|Albumin/Protein.total|Albumin/Protein.total
C0800927|T201|COMP|17820-2|LNC|Albumin/Protein.total|Albumin/Protein.total
C0800928|T201|COMP|17821-0|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C0800929|T201|COMP|17822-8|LNC|Cells.CD3+CD4+/100 cells|Cells.CD3+CD4+/100 cells
C0800930|T201|COMP|17823-6|LNC|Cells.CD45/100 cells|Cells.CD45/100 cells
C0800931|T201|COMP|17824-4|LNC|Cells.CD3+CD8+/100 cells|Cells.CD3+CD8+/100 cells
C0800932|T201|COMP|17825-1|LNC|Cells.CD41a/100 cells|Cells.CD41a/100 cells
C0800933|T201|COMP|17826-9|LNC|Cells.CD3/100 cells|Cells.CD3/100 cells
C0800934|T201|COMP|17827-7|LNC|Cells.CD2/100 cells|Cells.CD2/100 cells
C0800935|T201|COMP|17828-5|LNC|Cells.CD16/100 cells|Cells.CD16/100 cells
C0800936|T201|COMP|17829-3|LNC|Cells.CD19/100 cells|Cells.CD19/100 cells
C0800937|T201|COMP|17830-1|LNC|Centromere Ab|Centromere Ab
C0800940|T201|COMP|17833-5|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0800941|T201|COMP|17834-3|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0800942|T201|COMP|17835-0|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0800943|T201|COMP|17836-8|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0800944|T201|COMP|17837-6|LNC|Acid phosphatase.tartrate resistant|Acid phosphatase.tartrate resistant
C0800945|T201|COMP|17838-4|LNC|Alkaline phosphatase.bone|Alkaline phosphatase.bone
C0800946|T201|COMP|17839-2|LNC|Alpha fucosidase|Alpha fucosidase
C0800947|T201|COMP|17840-0|LNC|Alpha-L-iduronidase|Alpha-L-iduronidase
C0800948|T201|COMP|17841-8|LNC|Amylase|Amylase
C0800949|T201|COMP|17842-6|LNC|Cancer Ag 27-29|Cancer Ag 27-29
C0800950|T201|COMP|17843-4|LNC|Cancer Ag 72-4|Cancer Ag 72-4
C0800951|T201|COMP|17844-2|LNC|Estradiol.albumin bound|Estradiol.albumin bound
C0800952|T201|COMP|17845-9|LNC|Lipoprotein.alpha|Lipoprotein.alpha
C0800953|T201|COMP|17846-7|LNC|Lipoprotein.beta|Lipoprotein.beta
C0800954|T201|COMP|17847-5|LNC|Lipoprotein.pre-beta|Lipoprotein.pre-beta
C0800955|T201|COMP|17848-3|LNC|Reticulocytes/1000 erythrocytes|Reticulocytes/1000 erythrocytes
C0800956|T201|COMP|17849-1|LNC|Reticulocytes/100 erythrocytes|Reticulocytes/100 erythrocytes
C0800957|T201|COMP|17850-9|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C0800958|T201|COMP|17851-7|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0800959|T201|COMP|17852-5|LNC|Ureaplasma urealyticum|Ureaplasma urealyticum
C0800960|T201|COMP|17853-3|LNC|Ganglioside GM1b Ab.IgG|Ganglioside GM1b Ab.IgG
C0800961|T201|COMP|17854-1|LNC|Ganglioside GM1b Ab.IgM|Ganglioside GM1b Ab.IgM
C0800962|T201|COMP|17855-8|LNC|Hemoglobin A1c/Hemoglobin.total|Hemoglobin A1c/Hemoglobin.total
C0800963|T201|COMP|17856-6|LNC|Hemoglobin A1c/Hemoglobin.total|Hemoglobin A1c/Hemoglobin.total
C0800964|T201|COMP|17857-4|LNC|Rheumatoid factor|Rheumatoid factor
C0800965|T201|COMP|17858-2|LNC|Gamma glutamyl transferase|Gamma glutamyl transferase
C0800966|T201|COMP|17859-0|LNC|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C0800967|T201|COMP|17860-8|LNC|3-Methylhistidine|3-Methylhistidine
C0800968|T201|COMP|17861-6|LNC|Calcium|Calcium
C0800969|T201|COMP|17862-4|LNC|Calcium|Calcium
C0800970|T201|COMP|17863-2|LNC|Calcium.ionized|Calcium.ionized
C0800971|T201|COMP|17864-0|LNC|Calcium.ionized|Calcium.ionized
C0800972|T201|COMP|17865-7|LNC|Glucose^post 8H CFst|Glucose^post 8H CFst
C0800973|T201|COMP|17866-5|LNC|Carnitine/Creatinine|Carnitine/Creatinine
C0800974|T201|COMP|17867-3|LNC|Carnitine.free (C0)/Creatinine|Carnitine.free (C0)/Creatinine
C0800975|T201|COMP|17868-1|LNC|Acylcarnitine/Creatinine|Acylcarnitine/Creatinine
C0800976|T201|COMP|17869-9|LNC|Orotate/Creatinine|Orotate/Creatinine
C0800977|T201|COMP|17870-7|LNC|Orotidine/Creatinine|Orotidine/Creatinine
C0800978|T201|COMP|17871-5|LNC|Hemoglobin H|Hemoglobin H
C0800979|T201|COMP|17872-3|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0800980|T201|COMP|17898-8|LNC|Bacteria identified|Bacteria identified
C0800981|T201|COMP|17899-6|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0800982|T201|COMP|17900-2|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0800983|T201|COMP|17901-0|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C0800984|T201|COMP|17902-8|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C0800985|T201|COMP|17903-6|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0800986|T201|COMP|17909-3|LNC|Bacteria identified|Bacteria identified
C0800987|T201|COMP|17910-1|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0800988|T201|COMP|17911-9|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0800989|T201|COMP|17912-7|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C0800990|T201|COMP|17913-5|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C0800991|T201|COMP|17914-3|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0800992|T201|COMP|17915-0|LNC|Bacteria identified|Bacteria identified
C0800993|T201|COMP|17916-8|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0800994|T201|COMP|17917-6|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0800995|T201|COMP|17918-4|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C0800996|T201|COMP|17919-2|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C0800997|T201|COMP|17920-0|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0800998|T201|COMP|17921-8|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0800999|T201|COMP|17922-6|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0801000|T201|COMP|17925-9|LNC|Bacteria identified|Bacteria identified
C0801001|T201|COMP|17926-7|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0801002|T201|COMP|17927-5|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0801003|T201|COMP|17928-3|LNC|Bacteria identified|Bacteria identified
C0801004|T201|COMP|17929-1|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0801005|T201|COMP|17930-9|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0801006|T201|COMP|17931-7|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C0801007|T201|COMP|17932-5|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C0801008|T201|COMP|17933-3|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0801009|T201|COMP|17934-1|LNC|Bacteria identified|Bacteria identified
C0801010|T201|COMP|17935-8|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0801011|T201|COMP|17936-6|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0801012|T201|COMP|17950-7|LNC|Microorganism identified|Microorganism identified
C0801013|T201|COMP|17951-5|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0801014|T201|COMP|17952-3|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0801015|T201|COMP|17953-1|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C0801016|T201|COMP|17954-9|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C0801017|T201|COMP|17955-6|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0801018|T201|COMP|17956-4|LNC|Bacteria identified|Bacteria identified
C0801019|T201|COMP|17957-2|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0801020|T201|COMP|17958-0|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0801021|T201|COMP|17969-7|LNC|Bacteria identified|Bacteria identified
C0801022|T201|COMP|17970-5|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C0801023|T201|COMP|17971-3|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C0801024|T201|COMP|17972-1|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C0801025|T201|COMP|17973-9|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C0801026|T201|COMP|17974-7|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C0801229|T201|COMP|18180-0|LNC|Albumin|Albumin
C0801230|T201|COMP|18182-6|LNC|Osmolality|Osmolality
C0801231|T201|COMP|18183-4|LNC|Melatonin|Melatonin
C0801232|T201|COMP|18184-2|LNC|Erythrocyte sedimentation rate|Erythrocyte sedimentation rate
C0801234|T201|COMP|18186-7|LNC|Calcium|Calcium
C0801235|T201|COMP|18187-5|LNC|LORazepam|LORazepam
C0801236|T201|COMP|18188-3|LNC|Acebutolol|Acebutolol
C0801237|T201|COMP|18189-1|LNC|Acetone|Acetone
C0801238|T201|COMP|18190-9|LNC|Acid phosphatase.tartrate resistant|Acid phosphatase.tartrate resistant
C0801239|T201|COMP|18191-7|LNC|Amino acids|Amino acids
C0801240|T201|COMP|18192-5|LNC|Bacteria|Bacteria
C0801241|T201|COMP|18194-1|LNC|Barium|Barium
C0801242|T201|COMP|18195-8|LNC|Glucosylceramidase|Glucosylceramidase
C0801243|T201|COMP|18196-6|LNC|Beta-N-acetylhexosaminidase.A|Beta-N-acetylhexosaminidase.A
C0801244|T201|COMP|18197-4|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0801245|T201|COMP|18198-2|LNC|Blastomyces dermatitidis Ab.IgE|Blastomyces dermatitidis Ab.IgE
C0801246|T201|COMP|18199-0|LNC|Blastomyces dermatitidis Ab.IgG|Blastomyces dermatitidis Ab.IgG
C0801247|T201|COMP|18200-6|LNC|Blastomyces dermatitidis Ab.IgM|Blastomyces dermatitidis Ab.IgM
C0801248|T201|COMP|18201-4|LNC|Borrelia burgdorferi Ab.IgA|Borrelia burgdorferi Ab.IgA
C0801249|T201|COMP|18202-2|LNC|Borrelia burgdorferi Ab.IgA|Borrelia burgdorferi Ab.IgA
C0801250|T201|COMP|18203-0|LNC|Borrelia burgdorferi Ab.IgG+IgM|Borrelia burgdorferi Ab.IgG+IgM
C0801251|T201|COMP|18204-8|LNC|Caffeine renal clearance|Caffeine renal clearance
C0801252|T201|COMP|18205-5|LNC|Carbon disulfide|Carbon disulfide
C0801253|T201|COMP|18206-3|LNC|Catecholamines^7th specimen post XXX challenge|Catecholamines^7th specimen post XXX challenge
C0801254|T201|COMP|18208-9|LNC|Cocaine|Cocaine
C0801255|T201|COMP|18209-7|LNC|Ubiquinone 10|Ubiquinone 10
C0801256|T201|COMP|18210-5|LNC|Complement C1 esterase inhibitor bound Ab.IgG|Complement C1 esterase inhibitor bound Ab.IgG
C0801257|T201|COMP|18211-3|LNC|Complement C1 esterase inhibitor bound Ab.IgM|Complement C1 esterase inhibitor bound Ab.IgM
C0801258|T201|COMP|18212-1|LNC|Complement C1 esterase inhibitor free Ab.IgG|Complement C1 esterase inhibitor free Ab.IgG
C0801259|T201|COMP|18213-9|LNC|Complement C1 esterase inhibitor free Ab.IgM|Complement C1 esterase inhibitor free Ab.IgM
C0801260|T201|COMP|18214-7|LNC|Delta 5-Pregnanetriol|Delta 5-Pregnanetriol
C0801261|T201|COMP|18215-4|LNC|Delta alanine|Delta alanine
C0801262|T201|COMP|18216-2|LNC|Dezocine|Dezocine
C0801263|T201|COMP|18217-0|LNC|Epidermis Ab.IgA|Epidermis Ab.IgA
C0801264|T201|COMP|18218-8|LNC|Epidermis Ab.IgM|Epidermis Ab.IgM
C0801265|T201|COMP|18219-6|LNC|EPINEPHrine^2nd specimen post XXX challenge|EPINEPHrine^2nd specimen post XXX challenge
C0801266|T201|COMP|18220-4|LNC|EPINEPHrine^3rd specimen post XXX challenge|EPINEPHrine^3rd specimen post XXX challenge
C0801267|T201|COMP|18221-2|LNC|EPINEPHrine^4th specimen post XXX challenge|EPINEPHrine^4th specimen post XXX challenge
C0801268|T201|COMP|18222-0|LNC|EPINEPHrine^5th specimen post XXX challenge|EPINEPHrine^5th specimen post XXX challenge
C0801269|T201|COMP|18223-8|LNC|EPINEPHrine^6th specimen post XXX challenge|EPINEPHrine^6th specimen post XXX challenge
C0801270|T201|COMP|18224-6|LNC|EPINEPHrine^7th specimen post XXX challenge|EPINEPHrine^7th specimen post XXX challenge
C0801271|T201|COMP|18225-3|LNC|Erythrocyte shape|Erythrocyte shape
C0801272|T201|COMP|18226-1|LNC|Erythrocyte size|Erythrocyte size
C0801273|T201|COMP|18227-9|LNC|Glucose|Glucose
C0801274|T201|COMP|18228-7|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C0801275|T201|COMP|18229-5|LNC|Heparan sulfate|Heparan sulfate
C0801276|T201|COMP|18230-3|LNC|Histone H2a+H2b Ab|Histone H2a+H2b Ab
C0801277|T201|COMP|18231-1|LNC|Histone H2a+H2b Ab|Histone H2a+H2b Ab
C0801278|T201|COMP|18232-9|LNC|Hydrocorticosterone|Hydrocorticosterone
C0801279|T201|COMP|18233-7|LNC|Influenza virus Ab|Influenza virus Ab
C0801280|T201|COMP|18234-5|LNC|Insulin|Insulin
C0801281|T201|COMP|18235-2|LNC|Ketone solvents|Ketone solvents
C0801282|T201|COMP|18236-0|LNC|Lead|Lead
C0801283|T201|COMP|18237-8|LNC|Legionella pneumophila atypical Ab.IgM|Legionella pneumophila atypical Ab.IgM
C0801284|T201|COMP|18238-6|LNC|Lithium|Lithium
C0801285|T201|COMP|18239-4|LNC|Lupus erythematosus factor|Lupus erythematosus factor
C0801286|T201|COMP|18240-2|LNC|1,3-Dichlorobenzene|1,3-Dichlorobenzene
C0801287|T201|COMP|18241-0|LNC|cefOXitin Ab.IgE|cefOXitin Ab.IgE
C0801288|T201|COMP|18242-8|LNC|Methyprylon|Methyprylon
C0801289|T201|COMP|18243-6|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C0801290|T201|COMP|18244-4|LNC|Niacin|Niacin
C0801291|T201|COMP|18245-1|LNC|Nickel|Nickel
C0801292|T201|COMP|18246-9|LNC|Nitrogen|Nitrogen
C0801293|T201|COMP|18247-7|LNC|Nitrogen|Nitrogen
C0801294|T201|COMP|18248-5|LNC|Nordiazepam|Nordiazepam
C0801295|T201|COMP|18249-3|LNC|Para aminobenzoate|Para aminobenzoate
C0801296|T201|COMP|18250-1|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C0801297|T201|COMP|18251-9|LNC|Polychlorinated biphenyl|Polychlorinated biphenyl
C0801298|T201|COMP|18252-7|LNC|predniSONE|predniSONE
C0801299|T201|COMP|18253-5|LNC|Serotonin|Serotonin
C0801300|T201|COMP|18254-3|LNC|Silicate|Silicate
C0801301|T201|COMP|18255-0|LNC|Sulfonylurea|Sulfonylurea
C0801302|T201|COMP|18256-8|LNC|Sulfonylurea|Sulfonylurea
C0801303|T201|COMP|18257-6|LNC|Coproporphyrin|Coproporphyrin
C0801304|T201|COMP|18258-4|LNC|Trimethoprim Ab.IgE|Trimethoprim Ab.IgE
C0801305|T201|COMP|18259-2|LNC|Vasoactive intestinal peptide|Vasoactive intestinal peptide
C0801306|T201|COMP|18260-0|LNC|Zinc|Zinc
C0801307|T201|COMP|18261-8|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C0801308|T201|COMP|18262-6|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C0801309|T201|COMP|18263-4|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C0801310|T201|COMP|18264-2|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C0801311|T201|COMP|18265-9|LNC|Acetaminophen|Acetaminophen
C0801312|T201|COMP|18266-7|LNC|Cells.CD3+CD4+/Cells.CD3+CD8+|Cells.CD3+CD4+/Cells.CD3+CD8+
C0801313|T201|COMP|18267-5|LNC|Cells.CD16+CD56+/100 cells|Cells.CD16+CD56+/100 cells
C0801314|T201|COMP|18268-3|LNC|Cells.CD16+CD56+/100 cells|Cells.CD16+CD56+/100 cells
C0801315|T201|COMP|18269-1|LNC|Immune complex|Immune complex
C0801316|T201|COMP|18270-9|LNC|carBAMazepine 10,11-Epoxide|carBAMazepine 10,11-Epoxide
C0801317|T201|COMP|18271-7|LNC|Alpha 1 antitrypsin fecal clearance|Alpha 1 antitrypsin fecal clearance
C0801318|T201|COMP|18272-5|LNC|RNA Ab|RNA Ab
C0801319|T201|COMP|18273-3|LNC|Blood group antibody screen|Blood group antibody screen
C0801320|T201|COMP|18274-1|LNC|Blood group antibody screen|Blood group antibody screen
C0801321|T201|COMP|18275-8|LNC|Blood group antigens present|Blood group antigens present
C0801322|T201|COMP|18276-6|LNC|Blood group antigens absent|Blood group antigens absent
C0801323|T201|COMP|18277-4|LNC|Hemoglobin F|Hemoglobin F
C0801324|T201|COMP|18278-2|LNC|Hemoglobin F|Hemoglobin F
C0801325|T201|COMP|18279-0|LNC|Hemoglobin F|Hemoglobin F
C0801326|T201|COMP|18280-8|LNC|Background stain|Background stain
C0801327|T201|COMP|18281-6|LNC|Calcium^^corrected for total protein|Calcium^^corrected for total protein
C0801328|T201|COMP|18282-4|LNC|Cannabinoids|Cannabinoids
C0801329|T201|COMP|18283-2|LNC|Cells.CD11/100 cells|Cells.CD11/100 cells
C0801330|T201|COMP|18284-0|LNC|Cells.CD198/100 cells|Cells.CD198/100 cells
C0801331|T201|COMP|18285-7|LNC|Cells.CDA/100 cells|Cells.CDA/100 cells
C0801332|T201|COMP|18286-5|LNC|Donath Landsteiner Ab|Donath Landsteiner Ab
C0801333|T201|COMP|18287-3|LNC|Donath Landsteiner Ab|Donath Landsteiner Ab
C0801334|T201|COMP|18288-1|LNC|Donath Landsteiner Ab|Donath Landsteiner Ab
C0801335|T201|COMP|18289-9|LNC|Erythrocytes|Erythrocytes
C0801336|T201|COMP|18290-7|LNC|Erythrocytes|Erythrocytes
C0801337|T201|COMP|18291-5|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C0801339|T201|COMP|18293-1|LNC|Hemoglobin.fetal/Hemoglobin.total^post partum|Hemoglobin.fetal/Hemoglobin.total^post partum
C0801341|T201|COMP|18295-6|LNC|Hemoglobin.fetal/Hemoglobin.total^pre partum|Hemoglobin.fetal/Hemoglobin.total^pre partum
C0801342|T201|COMP|18296-4|LNC|Glucose^post dose glucose|Glucose^post dose glucose
C0801343|T201|COMP|18297-2|LNC|Acid hemolysis|Acid hemolysis
C0801344|T201|COMP|18298-0|LNC|High titer low avidity Ab|High titer low avidity Ab
C0801345|T201|COMP|18299-8|LNC|IgA|IgA
C0801346|T201|COMP|18300-4|LNC|IgA|IgA
C0801347|T201|COMP|18301-2|LNC|IgG|IgG
C0801348|T201|COMP|18302-0|LNC|IgG|IgG
C0801349|T201|COMP|18303-8|LNC|IgM|IgM
C0801350|T201|COMP|18304-6|LNC|IgM|IgM
C0801351|T201|COMP|18305-3|LNC|Amoeba identified|Amoeba identified
C0801352|T201|COMP|18306-1|LNC|Hydatid cyst identified|Hydatid cyst identified
C0801353|T201|COMP|18307-9|LNC|Ova & parasites identified|Ova & parasites identified
C0801354|T201|COMP|18308-7|LNC|Pneumocystis sp identified|Pneumocystis sp identified
C0801355|T201|COMP|18309-5|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C0801356|T201|COMP|18310-3|LNC|Hemoglobin.other/Hemoglobin.total|Hemoglobin.other/Hemoglobin.total
C0801357|T201|COMP|18311-1|LNC|Pelger Huet cells|Pelger Huet cells
C0801358|T201|COMP|18312-9|LNC|Platelet satellitism|Platelet satellitism
C0801359|T201|COMP|18313-7|LNC|Coagulation|Coagulation
C0801360|T201|COMP|18314-5|LNC|Morphology|Morphology
C0801361|T201|COMP|18319-4|LNC|Neutrophils.vacuolated|Neutrophils.vacuolated
C0801362|T201|COMP|18320-2|LNC|Globulin|Globulin
C0801363|T201|COMP|18321-0|LNC|Benzidine|Benzidine
C0801364|T201|COMP|18322-8|LNC|Norketamine|Norketamine
C0801365|T201|COMP|18323-6|LNC|Smith extractable nuclear Ab.IgG|Smith extractable nuclear Ab.IgG
C0801366|T201|COMP|18324-4|LNC|Cockatiel serum Ab.IgE|Cockatiel serum Ab.IgE
C0801367|T201|COMP|18325-1|LNC|oxyMORphone|oxyMORphone
C0801371|T201|COMP|18329-3|LNC|Neutrophil cytoplasmic Ab.IgA|Neutrophil cytoplasmic Ab.IgA
C0801372|T201|COMP|18330-1|LNC|Neutrophil cytoplasmic Ab.IgG|Neutrophil cytoplasmic Ab.IgG
C0801373|T201|COMP|18331-9|LNC|Neutrophil cytoplasmic Ab.IgM|Neutrophil cytoplasmic Ab.IgM
C0801374|T201|COMP|18332-7|LNC|Thyroperoxidase Ab.IgG|Thyroperoxidase Ab.IgG
C0801375|T201|COMP|18333-5|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C0801376|T201|COMP|18334-3|LNC|Naltrexone|Naltrexone
C0801377|T201|COMP|18335-0|LNC|Antihistamines|Antihistamines
C0801378|T201|COMP|18336-8|LNC|Methyl tert-butyl ether|Methyl tert-butyl ether
C0801379|T201|COMP|18337-6|LNC|Hydroxyitraconazole|Hydroxyitraconazole
C0801380|T201|COMP|18338-4|LNC|Nortramadol|Nortramadol
C0801381|T201|COMP|18339-2|LNC|Nortramadol|Nortramadol
C0801382|T201|COMP|18340-0|LNC|Nortramadol|Nortramadol
C0801383|T201|COMP|18341-8|LNC|Propylene glycol|Propylene glycol
C0801384|T201|COMP|18342-6|LNC|Glucose^3H post XXX challenge|Glucose^3H post XXX challenge
C0801385|T201|COMP|18343-4|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0801386|T201|COMP|18344-2|LNC|Beta-N-acetylhexosaminidase|Beta-N-acetylhexosaminidase
C0801387|T201|COMP|18345-9|LNC|Protein S Ag/Coagulation factor VII Ag|Protein S Ag/Coagulation factor VII Ag
C0801388|T201|COMP|18346-7|LNC|Streptococcus pneumoniae 18c Ab.IgG|Streptococcus pneumoniae 18c Ab.IgG
C0801389|T201|COMP|18347-5|LNC|Streptococcus pneumoniae 12 Ab^2nd specimen|Streptococcus pneumoniae 12 Ab^2nd specimen
C0801390|T201|COMP|18348-3|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0801391|T201|COMP|18349-1|LNC|Cells.CD8+CD25+|Cells.CD8+CD25+
C0801392|T201|COMP|18350-9|LNC|Cells.CD8+CD57+|Cells.CD8+CD57+
C0801393|T201|COMP|18351-7|LNC|11-Deoxycortisol^2nd specimen post XXX challenge|11-Deoxycortisol^2nd specimen post XXX challenge
C0801394|T201|COMP|18352-5|LNC|Specimen volume|Specimen volume
C0801395|T201|COMP|18353-3|LNC|Glucose^6H post 50 g lactose PO|Glucose^6H post 50 g lactose PO
C0801396|T201|COMP|18354-1|LNC|Glucose^12H post 50 g lactose PO|Glucose^12H post 50 g lactose PO
C0801397|T201|COMP|18355-8|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0801398|T201|COMP|18356-6|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0801399|T201|COMP|18357-4|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0801400|T201|COMP|18358-2|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0801401|T201|COMP|18359-0|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0801402|T201|COMP|18360-8|LNC|8-Hydroxyamoxapine|8-Hydroxyamoxapine
C0801403|T201|COMP|18361-6|LNC|Adenosine monophosphate.cyclic/Creatinine|Adenosine monophosphate.cyclic/Creatinine
C0801404|T201|COMP|18362-4|LNC|Alpha-2-Retinol binding protein|Alpha-2-Retinol binding protein
C0801405|T201|COMP|18363-2|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C0801406|T201|COMP|18364-0|LNC|Chondroitin sulfate|Chondroitin sulfate
C0801407|T201|COMP|18365-7|LNC|Cortisol.free|Cortisol.free
C0801408|T201|COMP|18366-5|LNC|Cytochrome C oxidase|Cytochrome C oxidase
C0801409|T201|COMP|18367-3|LNC|Iodine.free|Iodine.free
C0801410|T201|COMP|18368-1|LNC|Magnesium|Magnesium
C0801411|T201|COMP|18369-9|LNC|Magnesium|Magnesium
C0801412|T201|COMP|18370-7|LNC|Nitrite|Nitrite
C0801413|T201|COMP|18371-5|LNC|Methyl parathion|Methyl parathion
C0801414|T201|COMP|18372-3|LNC|Potassium|Potassium
C0801415|T201|COMP|18373-1|LNC|Protein|Protein
C0801416|T201|COMP|18374-9|LNC|Riboflavin|Riboflavin
C0801417|T201|COMP|17003-5|LNC|Serotonin|Serotonin
C0801418|T201|COMP|18376-4|LNC|Sodium|Sodium
C0801419|T201|COMP|18377-2|LNC|Sodium|Sodium
C0801420|T201|COMP|18378-0|LNC|Transcortin|Transcortin
C0801421|T201|COMP|18379-8|LNC|Urate|Urate
C0801422|T201|COMP|18380-6|LNC|Uroporphyrinogen decarboxylase|Uroporphyrinogen decarboxylase
C0801423|T201|COMP|18381-4|LNC|Uroporphyrinogen decarboxylase|Uroporphyrinogen decarboxylase
C0801424|T201|COMP|18382-2|LNC|Specimen.dry weight|Specimen.dry weight
C0801425|T201|COMP|18383-0|LNC|Alfentanil|Alfentanil
C0801426|T201|COMP|18384-8|LNC|Butabarbital|Butabarbital
C0801427|T201|COMP|18385-5|LNC|Butalbital|Butalbital
C0801428|T201|COMP|18386-3|LNC|Chlorothiazide|Chlorothiazide
C0801429|T201|COMP|18387-1|LNC|Diamorphine|Diamorphine
C0801430|T201|COMP|18388-9|LNC|diazePAM|diazePAM
C0801431|T201|COMP|18389-7|LNC|Methaqualone|Methaqualone
C0801432|T201|COMP|18390-5|LNC|Opiates|Opiates
C0801433|T201|COMP|18391-3|LNC|Paraldehyde|Paraldehyde
C0801434|T201|COMP|18392-1|LNC|Phencyclidine|Phencyclidine
C0801435|T201|COMP|18393-9|LNC|quiNIDine+Quinine|quiNIDine+Quinine
C0801436|T201|COMP|18394-7|LNC|HLA-A24(9)|HLA-A24(9)
C0801437|T201|COMP|18395-4|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C0801438|T201|COMP|18396-2|LNC|HIV 1 p24 Ag|HIV 1 p24 Ag
C0801439|T201|COMP|18397-0|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C0801440|T201|COMP|18398-8|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C0801441|T201|COMP|18399-6|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C0801442|T201|COMP|18400-2|LNC|Spermatozoa Ab.IgA|Spermatozoa Ab.IgA
C0801443|T201|COMP|18401-0|LNC|Spermatozoa Ab.IgG|Spermatozoa Ab.IgG
C0801444|T201|COMP|18402-8|LNC|Spermatozoa Ab.IgA|Spermatozoa Ab.IgA
C0801445|T201|COMP|18403-6|LNC|Spermatozoa Ab.IgG|Spermatozoa Ab.IgG
C0801446|T201|COMP|18404-4|LNC|Spermatozoa Ab.IgM|Spermatozoa Ab.IgM
C0801447|T201|COMP|18405-1|LNC|Arsenate|Arsenate
C0801448|T201|COMP|18406-9|LNC|Arsenic trioxide|Arsenic trioxide
C0801449|T201|COMP|18407-7|LNC|Leukocytes|Leukocytes
C0801450|T201|COMP|18408-5|LNC|Cells.CD3+HLA-DR+/100 cells|Cells.CD3+HLA-DR+/100 cells
C0801451|T201|COMP|18409-3|LNC|Curvularia lunata Ab.IgG|Curvularia lunata Ab.IgG
C0801452|T201|COMP|18410-1|LNC|Epicoccum purpurascens Ab.IgG|Epicoccum purpurascens Ab.IgG
C0801453|T201|COMP|18411-9|LNC|Rhizopus nigricans Ab.IgG|Rhizopus nigricans Ab.IgG
C0801454|T201|COMP|18412-7|LNC|Stemphylium botryosum Ab.IgG|Stemphylium botryosum Ab.IgG
C0801455|T201|COMP|18413-5|LNC|HLA-DR16|HLA-DR16
C0801456|T201|COMP|18414-3|LNC|Psilocin|Psilocin
C0801457|T201|COMP|18415-0|LNC|Psilocin|Psilocin
C0801458|T201|COMP|18416-8|LNC|Aspergillus nidulans Ab.IgG|Aspergillus nidulans Ab.IgG
C0801459|T201|COMP|18417-6|LNC|Bean black Ab.IgG|Bean black Ab.IgG
C0801460|T201|COMP|18418-4|LNC|Casein Ab.IgA|Casein Ab.IgA
C0801461|T201|COMP|18419-2|LNC|Cephalosporine mold Ab.IgG|Cephalosporine mold Ab.IgG
C0801462|T201|COMP|18420-0|LNC|Chaetomium globosum Ab.IgG|Chaetomium globosum Ab.IgG
C0801463|T201|COMP|18421-8|LNC|Fusarium oxysporum Ab.IgG|Fusarium oxysporum Ab.IgG
C0801464|T201|COMP|18422-6|LNC|Microcytes|Microcytes
C0801465|T201|COMP|18423-4|LNC|Phthalic anhydride Ab.IgG|Phthalic anhydride Ab.IgG
C0801466|T201|COMP|18424-2|LNC|Phthalic anhydride Ab.IgM|Phthalic anhydride Ab.IgM
C0801467|T201|COMP|18425-9|LNC|Squash zucchini Ab.IgG|Squash zucchini Ab.IgG
C0801468|T201|COMP|18426-7|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C0801469|T201|COMP|18427-5|LNC|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C0801470|T201|COMP|18428-3|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0801471|T201|COMP|18429-1|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C0801472|T201|COMP|18430-9|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C0801473|T201|COMP|18431-7|LNC|Amphetamines|Amphetamines
C0801474|T201|COMP|18432-5|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0801476|T201|COMP|18434-1|LNC|1,2-Dichlorobenzene|1,2-Dichlorobenzene
C0801477|T201|COMP|18435-8|LNC|SUFentanil|SUFentanil
C0801478|T201|COMP|18436-6|LNC|Acetylcarnitine (C2)|Acetylcarnitine (C2)
C0801479|T201|COMP|18437-4|LNC|Acrylylcarnitine (C3:1)|Acrylylcarnitine (C3:1)
C0801480|T201|COMP|18438-2|LNC|Propionylcarnitine (C3)|Propionylcarnitine (C3)
C0801481|T201|COMP|18439-0|LNC|Butyrylcarnitine (C4)|Butyrylcarnitine (C4)
C0801482|T201|COMP|18440-8|LNC|Crotonylcarnitine (C4:1)|Crotonylcarnitine (C4:1)
C0801483|T201|COMP|18441-6|LNC|Isovalerylcarnitine (C5)|Isovalerylcarnitine (C5)
C0801484|T201|COMP|18442-4|LNC|3-Hydroxybutyrylcarnitine (C4-OH)|3-Hydroxybutyrylcarnitine (C4-OH)
C0801485|T201|COMP|18443-2|LNC|Hexanoylcarnitine (C6)|Hexanoylcarnitine (C6)
C0801486|T201|COMP|18444-0|LNC|3-Hydroxyisovalerylcarnitine (C5-OH)|3-Hydroxyisovalerylcarnitine (C5-OH)
C0801487|T201|COMP|18445-7|LNC|Benzoylcarnitine (BzCn)|Benzoylcarnitine (BzCn)
C0801488|T201|COMP|18446-5|LNC|Methylmalonylcarnitine (C4-DC)|Methylmalonylcarnitine (C4-DC)
C0801489|T201|COMP|18447-3|LNC|Octenoylcarnitine (C8:1)|Octenoylcarnitine (C8:1)
C0801490|T201|COMP|18448-1|LNC|Octanoylcarnitine (C8)|Octanoylcarnitine (C8)
C0801491|T201|COMP|18449-9|LNC|Glutarylcarnitine (C5-DC)|Glutarylcarnitine (C5-DC)
C0801492|T201|COMP|18450-7|LNC|Adipoylcarnitine (C6-DC)|Adipoylcarnitine (C6-DC)
C0801493|T201|COMP|18451-5|LNC|Cis-4-decenoylcarnitine (Cis 4 C10:1)|Cis-4-decenoylcarnitine (Cis 4 C10:1)
C0801494|T201|COMP|18452-3|LNC|Decanoylcarnitine (C10)|Decanoylcarnitine (C10)
C0801495|T201|COMP|18453-1|LNC|Suberylcarnitine (C8-DC)|Suberylcarnitine (C8-DC)
C0801496|T201|COMP|18454-9|LNC|Dodecenoylcarnitine (C12:1)|Dodecenoylcarnitine (C12:1)
C0801497|T201|COMP|18455-6|LNC|Dodecanoylcarnitine (C12)|Dodecanoylcarnitine (C12)
C0801498|T201|COMP|18456-4|LNC|Tetradecadienoylcarnitine (C14:2)|Tetradecadienoylcarnitine (C14:2)
C0801499|T201|COMP|18457-2|LNC|Tetradecenoylcarnitine (C14:1)|Tetradecenoylcarnitine (C14:1)
C0801500|T201|COMP|18458-0|LNC|3-Hydroxytetradecadienoylcarnitine (C14:2-OH)|3-Hydroxytetradecadienoylcarnitine (C14:2-OH)
C0801501|T201|COMP|18459-8|LNC|3-Hydroxytetradecenoylcarnitine (C14:1-OH)|3-Hydroxytetradecenoylcarnitine (C14:1-OH)
C0801502|T201|COMP|18460-6|LNC|Palmitoylcarnitine (C16)|Palmitoylcarnitine (C16)
C0801503|T201|COMP|18461-4|LNC|3-Hydroxypalmitoylcarnitine (C16-OH)|3-Hydroxypalmitoylcarnitine (C16-OH)
C0801504|T201|COMP|18462-2|LNC|Linoleoylcarnitine (C18:2)|Linoleoylcarnitine (C18:2)
C0801505|T201|COMP|18463-0|LNC|Oleoylcarnitine (C18:1)|Oleoylcarnitine (C18:1)
C0801506|T201|COMP|18464-8|LNC|3-Hydroxylinoleoylcarnitine (C18:2-OH)|3-Hydroxylinoleoylcarnitine (C18:2-OH)
C0801507|T201|COMP|18465-5|LNC|3-Hydroxyoleoylcarnitine (C18:1-OH)|3-Hydroxyoleoylcarnitine (C18:1-OH)
C0801508|T201|COMP|18466-3|LNC|Dicarboxyoleylcarnitine (C18:1-DC)|Dicarboxyoleylcarnitine (C18:1-DC)
C0801509|T201|COMP|18467-1|LNC|Venlafaxine|Venlafaxine
C0801510|T201|COMP|18468-9|LNC|Aspergillus fumigatus Ab|Aspergillus fumigatus Ab
C0801511|T201|COMP|18469-7|LNC|Methyclothiazide|Methyclothiazide
C0801512|T201|COMP|18470-5|LNC|Norclomipramine|Norclomipramine
C0801513|T201|COMP|18471-3|LNC|Metoclopramide|Metoclopramide
C0801514|T201|COMP|18472-1|LNC|Organophosphate pesticides|Organophosphate pesticides
C0801515|T201|COMP|18473-9|LNC|HYDROmorphone|HYDROmorphone
C0801516|T201|COMP|18475-4|LNC|Phenylalanine/Creatinine|Phenylalanine/Creatinine
C0801517|T201|COMP|18476-2|LNC|Uroporphyrinogen decarboxylase|Uroporphyrinogen decarboxylase
C0801518|T201|COMP|18477-0|LNC|Lithium|Lithium
C0801519|T201|COMP|18478-8|LNC|Human papilloma virus 16+18 DNA|Human papilloma virus 16+18 DNA
C0801520|T201|COMP|18479-6|LNC|Human papilloma virus 31+35+51 DNA|Human papilloma virus 31+35+51 DNA
C0801521|T201|COMP|18480-4|LNC|Human papilloma virus 6+11 DNA|Human papilloma virus 6+11 DNA
C0801522|T201|COMP|18481-2|LNC|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C0801523|T201|COMP|18482-0|LNC|Yeast|Yeast
C0801524|T201|COMP|18483-8|LNC|Yeast|Yeast
C0801525|T201|COMP|18484-6|LNC|Ku Ab|Ku Ab
C0801526|T201|COMP|18485-3|LNC|Mi-2 Ab|Mi-2 Ab
C0801527|T201|COMP|18486-1|LNC|Methylenediamine|Methylenediamine
C0801528|T201|COMP|18487-9|LNC|Broad casts|Broad casts
C0801529|T201|COMP|18488-7|LNC|Calcium|Calcium
C0801530|T201|COMP|18489-5|LNC|Valproate.protein bound|Valproate.protein bound
C0801531|T201|COMP|18490-3|LNC|Chlamydia trachomatis G+F+K Ab.IgA|Chlamydia trachomatis G+F+K Ab.IgA
C0801532|T201|COMP|18491-1|LNC|Chlamydia trachomatis G+F+K Ab.IgG|Chlamydia trachomatis G+F+K Ab.IgG
C0801533|T201|COMP|18492-9|LNC|Chlamydia trachomatis G+F+K Ab.IgM|Chlamydia trachomatis G+F+K Ab.IgM
C0801534|T201|COMP|18493-7|LNC|Ova & parasites identified^3rd specimen|Ova & parasites identified^3rd specimen
C0801535|T201|COMP|18494-5|LNC|Ova & parasites identified^2nd specimen|Ova & parasites identified^2nd specimen
C0801536|T201|COMP|18495-2|LNC|Ova & parasites identified^3rd specimen|Ova & parasites identified^3rd specimen
C0801537|T201|COMP|18496-0|LNC|Ova & parasites identified^2nd specimen|Ova & parasites identified^2nd specimen
C0801851|T201|COMP|18857-3|LNC|Almecillin|Almecillin
C0801853|T201|COMP|18860-7|LNC|Amikacin|Amikacin
C0801854|T201|COMP|18861-5|LNC|Amoxicillin|Amoxicillin
C0801855|T201|COMP|18862-3|LNC|Amoxicillin+Clavulanate|Amoxicillin+Clavulanate
C0801856|T201|COMP|18863-1|LNC|Amphotericin B|Amphotericin B
C0801857|T201|COMP|18864-9|LNC|Ampicillin|Ampicillin
C0801858|T201|COMP|18865-6|LNC|Ampicillin+Sulbactam|Ampicillin+Sulbactam
C0801859|T201|COMP|18866-4|LNC|Azithromycin|Azithromycin
C0801860|T201|COMP|18867-2|LNC|Azlocillin|Azlocillin
C0801861|T201|COMP|18868-0|LNC|Aztreonam|Aztreonam
C0801862|T201|COMP|18869-8|LNC|Bacampicillin|Bacampicillin
C0801863|T201|COMP|18870-6|LNC|Bacitracin|Bacitracin
C0801864|T201|COMP|18871-4|LNC|Butirosin|Butirosin
C0801865|T201|COMP|18872-2|LNC|Capreomycin|Capreomycin
C0801866|T201|COMP|18873-0|LNC|Carbenicillin|Carbenicillin
C0801867|T201|COMP|18874-8|LNC|Cefaclor|Cefaclor
C0801868|T201|COMP|18875-5|LNC|Cefadroxil|Cefadroxil
C0801869|T201|COMP|18876-3|LNC|Cefamandole|Cefamandole
C0801870|T201|COMP|18877-1|LNC|Cefatrizine|Cefatrizine
C0801871|T201|COMP|18878-9|LNC|ceFAZolin|ceFAZolin
C0801872|T201|COMP|18879-7|LNC|Cefepime|Cefepime
C0801873|T201|COMP|18880-5|LNC|Cefixime|Cefixime
C0801874|T201|COMP|18881-3|LNC|Cefmetazole|Cefmetazole
C0801875|T201|COMP|18882-1|LNC|Cefodizime|Cefodizime
C0801876|T201|COMP|18883-9|LNC|Cefonicid|Cefonicid
C0801877|T201|COMP|18884-7|LNC|Cefoperazone|Cefoperazone
C0801878|T201|COMP|18885-4|LNC|Ceforanide|Ceforanide
C0801879|T201|COMP|18886-2|LNC|Cefotaxime|Cefotaxime
C0801880|T201|COMP|18887-0|LNC|cefoTEtan|cefoTEtan
C0801881|T201|COMP|18888-8|LNC|cefOXitin|cefOXitin
C0801882|T201|COMP|18889-6|LNC|Cefpirome|Cefpirome
C0801883|T201|COMP|18890-4|LNC|Cefpodoxime|Cefpodoxime
C0801884|T201|COMP|18891-2|LNC|Cefprozil|Cefprozil
C0801885|T201|COMP|18892-0|LNC|Cefsulodin|Cefsulodin
C0801886|T201|COMP|18893-8|LNC|cefTAZidime|cefTAZidime
C0801887|T201|COMP|18894-6|LNC|Ceftizoxime|Ceftizoxime
C0801888|T201|COMP|18895-3|LNC|cefTRIAXone|cefTRIAXone
C0801889|T201|COMP|18896-1|LNC|Cefuroxime.parenteral|Cefuroxime.parenteral
C0801890|T201|COMP|18897-9|LNC|Cephalexin|Cephalexin
C0801891|T201|COMP|18898-7|LNC|Cephaloglycin|Cephaloglycin
C0801892|T201|COMP|18899-5|LNC|Cephaloridine|Cephaloridine
C0801893|T201|COMP|18900-1|LNC|Cephalothin|Cephalothin
C0801894|T201|COMP|18901-9|LNC|Cephapirin|Cephapirin
C0801895|T201|COMP|18902-7|LNC|Cephradine|Cephradine
C0801896|T201|COMP|18903-5|LNC|Chloramphenicol|Chloramphenicol
C0801897|T201|COMP|18904-3|LNC|Chlortetracycline|Chlortetracycline
C0801898|T201|COMP|18905-0|LNC|Cinoxacin|Cinoxacin
C0801899|T201|COMP|18906-8|LNC|Ciprofloxacin|Ciprofloxacin
C0801900|T201|COMP|18907-6|LNC|Clarithromycin|Clarithromycin
C0801901|T201|COMP|18908-4|LNC|Clindamycin|Clindamycin
C0801902|T201|COMP|18909-2|LNC|Clotrimazole|Clotrimazole
C0801903|T201|COMP|18910-0|LNC|Cloxacillin|Cloxacillin
C0801904|T201|COMP|18911-8|LNC|Colistimethate|Colistimethate
C0801905|T201|COMP|18912-6|LNC|Colistin|Colistin
C0801906|T201|COMP|18913-4|LNC|Cyclacillin|Cyclacillin
C0801907|T201|COMP|18914-2|LNC|cycloSERINE|cycloSERINE
C0801908|T201|COMP|18915-9|LNC|Demeclocycline|Demeclocycline
C0801910|T201|COMP|18917-5|LNC|Doxycycline|Doxycycline
C0801911|T201|COMP|18918-3|LNC|Enoxacin|Enoxacin
C0801912|T201|COMP|18919-1|LNC|Erythromycin|Erythromycin
C0801913|T201|COMP|18920-9|LNC|Erythromycin+sulfiSOXAZOLE|Erythromycin+sulfiSOXAZOLE
C0801914|T201|COMP|18921-7|LNC|Ethambutol|Ethambutol
C0801915|T201|COMP|18922-5|LNC|Ethionamide|Ethionamide
C0801916|T201|COMP|18923-3|LNC|Floxacillin|Floxacillin
C0801917|T201|COMP|18924-1|LNC|Fluconazole|Fluconazole
C0801918|T201|COMP|18855-7|LNC|5-Fluorocytosine|5-Fluorocytosine
C0801919|T201|COMP|18926-6|LNC|Framycetin|Framycetin
C0801920|T201|COMP|18927-4|LNC|Fusidate|Fusidate
C0801921|T201|COMP|18928-2|LNC|Gentamicin|Gentamicin
C0801922|T201|COMP|18929-0|LNC|Gentamicin.high potency|Gentamicin.high potency
C0801923|T201|COMP|18930-8|LNC|Gramicidin D|Gramicidin D
C0801924|T201|COMP|18931-6|LNC|Hetacillin|Hetacillin
C0801925|T201|COMP|18932-4|LNC|Imipenem|Imipenem
C0801926|T201|COMP|18933-2|LNC|Imipenem+Cilastatin|Imipenem+Cilastatin
C0801927|T201|COMP|18934-0|LNC|Isoniazid|Isoniazid
C0801928|T201|COMP|18935-7|LNC|Kanamycin|Kanamycin
C0801929|T201|COMP|18936-5|LNC|Kanamycin.high potency|Kanamycin.high potency
C0801930|T201|COMP|18937-3|LNC|Ketoconazole|Ketoconazole
C0801931|T201|COMP|18938-1|LNC|Lincomycin|Lincomycin
C0801932|T201|COMP|18939-9|LNC|Lomefloxacin|Lomefloxacin
C0801933|T201|COMP|18940-7|LNC|Loracarbef|Loracarbef
C0801934|T201|COMP|18941-5|LNC|Lymecycline|Lymecycline
C0801935|T201|COMP|18942-3|LNC|Meclocycline|Meclocycline
C0801936|T201|COMP|18943-1|LNC|Meropenem|Meropenem
C0801937|T201|COMP|18944-9|LNC|Methacycline|Methacycline
C0801938|T201|COMP|18945-6|LNC|Methicillin|Methicillin
C0801939|T201|COMP|18946-4|LNC|metroNIDAZOLE|metroNIDAZOLE
C0801940|T201|COMP|18947-2|LNC|Mezlocillin|Mezlocillin
C0801941|T201|COMP|18948-0|LNC|Minocycline|Minocycline
C0801942|T201|COMP|18949-8|LNC|Miocamycin|Miocamycin
C0801943|T201|COMP|18950-6|LNC|Moxalactam|Moxalactam
C0801944|T201|COMP|18951-4|LNC|Nafcillin|Nafcillin
C0801945|T201|COMP|18952-2|LNC|Nalidixate|Nalidixate
C0801946|T201|COMP|18953-0|LNC|Neomycin|Neomycin
C0801947|T201|COMP|18954-8|LNC|Netilmicin|Netilmicin
C0801948|T201|COMP|18955-5|LNC|Nitrofurantoin|Nitrofurantoin
C0801949|T201|COMP|18956-3|LNC|Norfloxacin|Norfloxacin
C0801950|T201|COMP|18957-1|LNC|Novobiocin|Novobiocin
C0801951|T201|COMP|18958-9|LNC|Nystatin|Nystatin
C0801952|T201|COMP|18959-7|LNC|Ofloxacin|Ofloxacin
C0801953|T201|COMP|18960-5|LNC|Oleandomycin|Oleandomycin
C0801954|T201|COMP|18961-3|LNC|Oxacillin|Oxacillin
C0801955|T201|COMP|18962-1|LNC|Oxytetracycline|Oxytetracycline
C0801956|T201|COMP|18963-9|LNC|Pefloxacin|Pefloxacin
C0801957|T201|COMP|18964-7|LNC|Penicillin|Penicillin
C0801958|T201|COMP|18965-4|LNC|Penicillin G|Penicillin G
C0801959|T201|COMP|18966-2|LNC|Penicillin V|Penicillin V
C0801960|T201|COMP|18967-0|LNC|Phenethicillin|Phenethicillin
C0801961|T201|COMP|18968-8|LNC|Pipemidate|Pipemidate
C0801962|T201|COMP|18969-6|LNC|Piperacillin|Piperacillin
C0801963|T201|COMP|18970-4|LNC|Piperacillin+Tazobactam|Piperacillin+Tazobactam
C0801964|T201|COMP|18971-2|LNC|Pivampicillin|Pivampicillin
C0801965|T201|COMP|18972-0|LNC|Polymyxin B|Polymyxin B
C0801966|T201|COMP|18973-8|LNC|Pyrazinamide|Pyrazinamide
C0801967|T201|COMP|18974-6|LNC|rifAMPin|rifAMPin
C0801968|T201|COMP|18975-3|LNC|Ristocetin|Ristocetin
C0801969|T201|COMP|18976-1|LNC|Rolitetracycline|Rolitetracycline
C0801970|T201|COMP|18977-9|LNC|Rosoxacin|Rosoxacin
C0801971|T201|COMP|18978-7|LNC|Roxithromycin|Roxithromycin
C0801972|T201|COMP|18979-5|LNC|Sisomicin|Sisomicin
C0801973|T201|COMP|18980-3|LNC|Spectinomycin|Spectinomycin
C0801974|T201|COMP|18981-1|LNC|Spiramycin|Spiramycin
C0801975|T201|COMP|18982-9|LNC|Streptomycin|Streptomycin
C0801976|T201|COMP|18983-7|LNC|Streptomycin.high potency|Streptomycin.high potency
C0801977|T201|COMP|18984-5|LNC|sulfADIAZINE|sulfADIAZINE
C0801978|T201|COMP|18985-2|LNC|Sulfamethoxazole|Sulfamethoxazole
C0801979|T201|COMP|18986-0|LNC|sulfiSOXAZOLE|sulfiSOXAZOLE
C0801980|T201|COMP|18987-8|LNC|Sulfonamide|Sulfonamide
C0801981|T201|COMP|18988-6|LNC|Talampicillin|Talampicillin
C0801982|T201|COMP|18989-4|LNC|Teicoplanin|Teicoplanin
C0801983|T201|COMP|18990-2|LNC|Temafloxacin|Temafloxacin
C0801984|T201|COMP|18991-0|LNC|Temocillin|Temocillin
C0801985|T201|COMP|18992-8|LNC|Terbinafine|Terbinafine
C0801986|T201|COMP|18993-6|LNC|Tetracycline|Tetracycline
C0801987|T201|COMP|18994-4|LNC|Ticarcillin|Ticarcillin
C0801988|T201|COMP|18995-1|LNC|Ticarcillin+Clavulanate|Ticarcillin+Clavulanate
C0801989|T201|COMP|18996-9|LNC|Tobramycin|Tobramycin
C0801990|T201|COMP|18997-7|LNC|Trimethoprim|Trimethoprim
C0801991|T201|COMP|18998-5|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0801992|T201|COMP|18999-3|LNC|Troleandomycin|Troleandomycin
C0801993|T201|COMP|19000-9|LNC|Vancomycin|Vancomycin
C0801994|T201|COMP|19001-7|LNC|Viomycin|Viomycin
C0802011|T201|COMP|19022-3|LNC|Neisseria meningitidis serogroups C+w135 Ag|Neisseria meningitidis serogroups C+w135 Ag
C0802012|T201|COMP|19023-1|LNC|Granulocytes/100 leukocytes|Granulocytes/100 leukocytes
C0802013|T201|COMP|19057-9|LNC|ABO & Rh group|ABO & Rh group
C0802014|T201|COMP|19058-7|LNC|Allergens identified|Allergens identified
C0802015|T201|COMP|19059-5|LNC|Amphetamines cutoff|Amphetamines cutoff
C0802016|T201|COMP|888-8|LNC|Blood group antibodies identified|Blood group antibodies identified
C0802017|T201|COMP|19064-5|LNC|Benzodiazepines cutoff|Benzodiazepines cutoff
C0802018|T201|COMP|19065-2|LNC|Benzoylecgonine cutoff|Benzoylecgonine cutoff
C0802019|T201|COMP|19066-0|LNC|Blood bank comment|Blood bank comment
C0802020|T201|COMP|19071-0|LNC|Blood removed from patient|Blood removed from patient
C0802021|T201|COMP|19073-6|LNC|Cannabinoids cutoff|Cannabinoids cutoff
C0802022|T201|COMP|19074-4|LNC|Carnitine esters|Carnitine esters
C0802023|T201|COMP|19075-1|LNC|Cells counted.total|Cells counted.total
C0802024|T201|COMP|19076-9|LNC|Cells counted.total|Cells counted.total
C0802025|T201|COMP|19077-7|LNC|Cells identified|Cells identified
C0802027|T201|COMP|19079-3|LNC|Cells.CD43/100 cells|Cells.CD43/100 cells
C0802028|T201|COMP|19080-1|LNC|Choriogonadotropin|Choriogonadotropin
C0802029|T201|COMP|13362-9|LNC|Collection duration|Collection duration
C0802030|T201|COMP|19086-8|LNC|Collection end date|Collection end date
C0802031|T201|COMP|19087-6|LNC|Collection end time|Collection end time
C0802032|T201|COMP|19088-4|LNC|Collection start date|Collection start date
C0802033|T201|COMP|19089-2|LNC|Collection start time|Collection start time
C0802034|T201|COMP|19090-0|LNC|Colony count|Colony count
C0802035|T201|COMP|19091-8|LNC|Colony count|Colony count
C0802036|T201|COMP|19092-6|LNC|Cotinine cutoff|Cotinine cutoff
C0802037|T201|COMP|19096-7|LNC|Electrolytes|Electrolytes
C0802038|T201|COMP|19098-3|LNC|Erythrocytes|Erythrocytes
C0802039|T201|COMP|19099-1|LNC|Events counted|Events counted
C0802040|T201|COMP|19101-5|LNC|Fungus colony count|Fungus colony count
C0802041|T201|COMP|19102-3|LNC|Genetic screen|Genetic screen
C0802042|T201|COMP|19104-9|LNC|Glucose^1H post dose glucose|Glucose^1H post dose glucose
C0802043|T201|COMP|19105-6|LNC|Glucose^3H post dose glucose|Glucose^3H post dose glucose
C0802044|T201|COMP|19106-4|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C0802045|T201|COMP|19107-2|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C0802046|T201|COMP|19108-0|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C0802047|T201|COMP|19109-8|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C0802048|T201|COMP|19110-6|LNC|HIV 1 gp41+gp43 Ab|HIV 1 gp41+gp43 Ab
C0802050|T201|COMP|19113-0|LNC|IgE|IgE
C0802051|T201|COMP|19114-8|LNC|Lamellar bodies|Lamellar bodies
C0802052|T201|COMP|19122-1|LNC|Cells.CD42/100 cells|Cells.CD42/100 cells
C0802053|T201|COMP|19123-9|LNC|Magnesium|Magnesium
C0802054|T201|COMP|19124-7|LNC|Magnesium|Magnesium
C0802055|T201|COMP|19125-4|LNC|Meconium|Meconium
C0802056|T201|COMP|19126-2|LNC|Bacteria identified|Bacteria identified
C0802057|T201|COMP|19127-0|LNC|Bacteria identified|Bacteria identified
C0802058|T201|COMP|19128-8|LNC|Bacteria identified|Bacteria identified
C0802061|T201|COMP|19133-8|LNC|Neisseria meningitidis serogroups A+C+w135+Y Ag|Neisseria meningitidis serogroups A+C+w135+Y Ag
C0802063|T201|COMP|19137-9|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C0802064|T201|COMP|19138-7|LNC|Opiates cutoff|Opiates cutoff
C0802066|T201|COMP|19140-3|LNC|Phospholipid Ab|Phospholipid Ab
C0802068|T201|COMP|19144-5|LNC|Reason for drug test|Reason for drug test
C0802069|T201|COMP|19145-2|LNC|Reference lab test name|Reference lab test name
C0802070|T201|COMP|19146-0|LNC|Reference lab test results|Reference lab test results
C0802071|T201|COMP|19147-8|LNC|Reference lab test reference range|Reference lab test reference range
C0802072|T201|COMP|19148-6|LNC|Rh immune globulin candidate (yes/no)|Rh immune globulin candidate (yes/no)
C0802073|T201|COMP|19149-4|LNC|Rifabutin|Rifabutin
C0802074|T201|COMP|19150-2|LNC|Specimen creatinine acceptable|Specimen creatinine acceptable
C0802075|T201|COMP|19151-0|LNC|Specimen drawn|Specimen drawn
C0802076|T201|COMP|19152-8|LNC|Specimen specific gravity acceptable|Specimen specific gravity acceptable
C0802077|T201|COMP|19153-6|LNC|Specimen volume|Specimen volume
C0802078|T201|COMP|19156-9|LNC|Susceptibility method|Susceptibility method
C0802079|T201|COMP|19157-7|LNC|Tube number|Tube number
C0802080|T201|COMP|19158-5|LNC|Urea nitrogen comment|Urea nitrogen comment
C0802081|T201|COMP|19159-3|LNC|Urinalysis specimen collection method|Urinalysis specimen collection method
C0802082|T201|COMP|19161-9|LNC|Urobilinogen|Urobilinogen
C0802083|T201|COMP|19162-7|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0802084|T201|COMP|19163-5|LNC|Cancer Ag 19-9|Cancer Ag 19-9
C0802085|T201|COMP|19164-3|LNC|Cancer Ag 72-4|Cancer Ag 72-4
C0802086|T201|COMP|19165-0|LNC|Cancer Ag 125|Cancer Ag 125
C0802087|T201|COMP|19166-8|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0802088|T201|COMP|19167-6|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0802089|T201|COMP|19168-4|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0802090|T201|COMP|19169-2|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0802091|T201|COMP|19170-0|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C0802092|T201|COMP|19171-8|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0802093|T201|COMP|19172-6|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0802094|T201|COMP|19173-4|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0802095|T201|COMP|19174-2|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0802096|T201|COMP|19175-9|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0802097|T201|COMP|19176-7|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0802098|T201|COMP|19177-5|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0802099|T201|COMP|19178-3|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C0802100|T201|COMP|19179-1|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C0802101|T201|COMP|19180-9|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C0802102|T201|COMP|19182-5|LNC|Cytokeratin 19|Cytokeratin 19
C0802103|T201|COMP|19183-3|LNC|Cytokeratin 19|Cytokeratin 19
C0802104|T201|COMP|19184-1|LNC|Tissue polypeptide specific Ag|Tissue polypeptide specific Ag
C0802105|T201|COMP|19185-8|LNC|Tissue polypeptide specific Ag|Tissue polypeptide specific Ag
C0802106|T201|COMP|19186-6|LNC|Cancer Ag 15-3|Cancer Ag 15-3
C0802107|T201|COMP|19187-4|LNC|Cancer Ag 27-29|Cancer Ag 27-29
C0802108|T201|COMP|19188-2|LNC|Mucin-like carcinoma associated Ag|Mucin-like carcinoma associated Ag
C0802109|T201|COMP|19189-0|LNC|Cancer Ag 549|Cancer Ag 549
C0802110|T201|COMP|19190-8|LNC|Cancer Ag 549|Cancer Ag 549
C0802111|T201|COMP|19193-2|LNC|Enolase.neuron specific|Enolase.neuron specific
C0802112|T201|COMP|19194-0|LNC|Enolase.neuron specific|Enolase.neuron specific
C0802113|T201|COMP|19195-7|LNC|Prostate specific Ag|Prostate specific Ag
C0802114|T201|COMP|19197-3|LNC|Prostate specific Ag|Prostate specific Ag
C0802115|T201|COMP|19198-1|LNC|Prostate specific Ag|Prostate specific Ag
C0802116|T201|COMP|19199-9|LNC|Prostate specific Ag|Prostate specific Ag
C0802117|T201|COMP|19200-5|LNC|Prostate specific Ag|Prostate specific Ag
C0802118|T201|COMP|19201-3|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C0802119|T201|COMP|19203-9|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C0802120|T201|COMP|19204-7|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C0802121|T201|COMP|19205-4|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C0802122|T201|COMP|19206-2|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C0802123|T201|COMP|19207-0|LNC|Squamous cell carcinoma Ag|Squamous cell carcinoma Ag
C0802124|T201|COMP|19208-8|LNC|Squamous cell carcinoma Ag|Squamous cell carcinoma Ag
C0802125|T201|COMP|19209-6|LNC|Squamous cell carcinoma Ag|Squamous cell carcinoma Ag
C0802126|T201|COMP|19210-4|LNC|Squamous cell carcinoma Ag|Squamous cell carcinoma Ag
C0802127|T201|COMP|19211-2|LNC|Oxygen|Oxygen
C0802128|T201|COMP|19212-0|LNC|Carbon dioxide|Carbon dioxide
C0802130|T201|COMP|19217-9|LNC|Oxygen^^saturation adjusted to 0.5|Oxygen^^saturation adjusted to 0.5
C0802131|T201|COMP|19218-7|LNC|Oxygen content|Oxygen content
C0802132|T201|COMP|19219-5|LNC|Oxygen content|Oxygen content
C0802133|T201|COMP|19220-3|LNC|Oxygen content|Oxygen content
C0802134|T201|COMP|19221-1|LNC|Oxygen content|Oxygen content
C0802135|T201|COMP|19223-7|LNC|Carbon dioxide|Carbon dioxide
C0802137|T201|COMP|19225-2|LNC|Deoxyhemoglobin/Hemoglobin.total|Deoxyhemoglobin/Hemoglobin.total
C0802138|T201|COMP|19226-0|LNC|Deoxyhemoglobin/Hemoglobin.total|Deoxyhemoglobin/Hemoglobin.total
C0802139|T201|COMP|19227-8|LNC|Deoxyhemoglobin/Hemoglobin.total|Deoxyhemoglobin/Hemoglobin.total
C0802140|T201|COMP|19228-6|LNC|Deoxyhemoglobin/Hemoglobin.total|Deoxyhemoglobin/Hemoglobin.total
C0802141|T201|COMP|19229-4|LNC|Bicarbonate|Bicarbonate
C0802142|T201|COMP|19232-8|LNC|Bicarbonate^^standard|Bicarbonate^^standard
C0802143|T201|COMP|19234-4|LNC|Base excess|Base excess
C0802144|T201|COMP|19239-3|LNC|Lactate|Lactate
C0802145|T201|COMP|19240-1|LNC|Lactate|Lactate
C0802146|T201|COMP|19242-7|LNC|Corticotropin^post XXX challenge|Corticotropin^post XXX challenge
C0802147|T201|COMP|19243-5|LNC|Brucella abortus Ab|Brucella abortus Ab
C0802148|T201|COMP|19244-3|LNC|Character|Character
C0802149|T201|COMP|19245-0|LNC|clonazePAM|clonazePAM
C0802150|T201|COMP|19247-6|LNC|Doxepin+Metabolites|Doxepin+Metabolites
C0802151|T201|COMP|19248-4|LNC|Lactate dehydrogenase 2|Lactate dehydrogenase 2
C0802152|T201|COMP|19249-2|LNC|Lactose^3H post 50 g lactose PO|Lactose^3H post 50 g lactose PO
C0802153|T201|COMP|19250-0|LNC|Lipoprotein.alpha|Lipoprotein.alpha
C0802154|T201|COMP|19251-8|LNC|Prolactin^post XXX challenge|Prolactin^post XXX challenge
C0802155|T201|COMP|19252-6|LNC|Megakaryocytes/100 leukocytes|Megakaryocytes/100 leukocytes
C0802156|T201|COMP|19253-4|LNC|Trichinella spiralis Ab|Trichinella spiralis Ab
C0802157|T201|COMP|19254-2|LNC|Oxygen^^adjusted to patient's actual temperature|Oxygen^^adjusted to patient's actual temperature
C0802158|T201|COMP|19257-5|LNC|Oxygen^^adjusted to patient's actual temperature|Oxygen^^adjusted to patient's actual temperature
C0802159|T201|COMP|19259-1|LNC|Neisseria meningitidis serogroups A+C+w135+Y Ag|Neisseria meningitidis serogroups A+C+w135+Y Ag
C0802161|T201|COMP|19261-7|LNC|Amphetamines|Amphetamines
C0802162|T201|COMP|19262-5|LNC|Amphetamines tested for|Amphetamines tested for
C0802163|T201|COMP|19263-3|LNC|Amphetamines tested for|Amphetamines tested for
C0802164|T201|COMP|19265-8|LNC|Amphetamines positive|Amphetamines positive
C0802165|T201|COMP|19266-6|LNC|Amphetamines cutoff|Amphetamines cutoff
C0802166|T201|COMP|19267-4|LNC|Amphetamines cutoff|Amphetamines cutoff
C0802167|T201|COMP|19268-2|LNC|Amphetamines screen method|Amphetamines screen method
C0802168|T201|COMP|19269-0|LNC|Amphetamines confirm method|Amphetamines confirm method
C0802169|T201|COMP|19270-8|LNC|Barbiturates|Barbiturates
C0802170|T201|COMP|19271-6|LNC|Barbiturates tested for|Barbiturates tested for
C0802171|T201|COMP|19272-4|LNC|Barbiturates tested for|Barbiturates tested for
C0802172|T201|COMP|19274-0|LNC|Barbiturates positive|Barbiturates positive
C0802173|T201|COMP|19275-7|LNC|Barbiturates cutoff|Barbiturates cutoff
C0802174|T201|COMP|19276-5|LNC|Barbiturates cutoff|Barbiturates cutoff
C0802175|T201|COMP|19277-3|LNC|Barbiturates screen method|Barbiturates screen method
C0802176|T201|COMP|19278-1|LNC|Barbiturates confirm method|Barbiturates confirm method
C0802177|T201|COMP|19279-9|LNC|Benzodiazepines tested for|Benzodiazepines tested for
C0802179|T201|COMP|19282-3|LNC|Benzodiazepines positive|Benzodiazepines positive
C0802180|T201|COMP|19283-1|LNC|Benzodiazepines cutoff|Benzodiazepines cutoff
C0802181|T201|COMP|19284-9|LNC|Benzodiazepines cutoff|Benzodiazepines cutoff
C0802182|T201|COMP|19285-6|LNC|Benzodiazepines screen method|Benzodiazepines screen method
C0802183|T201|COMP|19286-4|LNC|Benzodiazepines confirm method|Benzodiazepines confirm method
C0802184|T201|COMP|19287-2|LNC|Cannabinoids tested for|Cannabinoids tested for
C0802185|T201|COMP|19288-0|LNC|Cannabinoids tested for|Cannabinoids tested for
C0802186|T201|COMP|19289-8|LNC|Cannabinoids|Cannabinoids
C0802187|T201|COMP|19290-6|LNC|Cannabinoids positive|Cannabinoids positive
C0802188|T201|COMP|19291-4|LNC|Cannabinoids cutoff|Cannabinoids cutoff
C0802189|T201|COMP|19292-2|LNC|Cannabinoids cutoff|Cannabinoids cutoff
C0802190|T201|COMP|19293-0|LNC|Cannabinoids screen method|Cannabinoids screen method
C0802191|T201|COMP|19294-8|LNC|Cannabinoids confirm method|Cannabinoids confirm method
C0802192|T201|COMP|19295-5|LNC|Opiates|Opiates
C0802193|T201|COMP|19296-3|LNC|Opiates tested for|Opiates tested for
C0802195|T201|COMP|19298-9|LNC|Opiates positive|Opiates positive
C0802196|T201|COMP|19299-7|LNC|Opiates cutoff|Opiates cutoff
C0802197|T201|COMP|19300-3|LNC|Opiates cutoff|Opiates cutoff
C0802198|T201|COMP|19301-1|LNC|Opiates screen method|Opiates screen method
C0802199|T201|COMP|19302-9|LNC|Opiates confirm method|Opiates confirm method
C0802200|T201|COMP|19303-7|LNC|Thiazides|Thiazides
C0802201|T201|COMP|19304-5|LNC|Thiazides tested for|Thiazides tested for
C0802202|T201|COMP|19305-2|LNC|Thiazides tested for|Thiazides tested for
C0802203|T201|COMP|19306-0|LNC|Thiazides|Thiazides
C0802204|T201|COMP|19307-8|LNC|Thiazides positive|Thiazides positive
C0802205|T201|COMP|19308-6|LNC|Thiazides cutoff|Thiazides cutoff
C0802206|T201|COMP|19309-4|LNC|Thiazides cutoff|Thiazides cutoff
C0802207|T201|COMP|19310-2|LNC|Thiazides screen method|Thiazides screen method
C0802208|T201|COMP|19311-0|LNC|Thiazides confirm method|Thiazides confirm method
C0802209|T201|COMP|19312-8|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0802210|T201|COMP|19313-6|LNC|Tricyclic antidepressants tested for|Tricyclic antidepressants tested for
C0802211|T201|COMP|19314-4|LNC|Tricyclic antidepressants tested for|Tricyclic antidepressants tested for
C0802212|T201|COMP|19315-1|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0802213|T201|COMP|19316-9|LNC|Tricyclic antidepressants positive|Tricyclic antidepressants positive
C0802214|T201|COMP|19317-7|LNC|Tricyclic antidepressants cutoff|Tricyclic antidepressants cutoff
C0802215|T201|COMP|19318-5|LNC|Tricyclic antidepressants cutoff|Tricyclic antidepressants cutoff
C0802216|T201|COMP|19319-3|LNC|Tricyclic antidepressants screen method|Tricyclic antidepressants screen method
C0802217|T201|COMP|19320-1|LNC|Tricyclic antidepressants confirm method|Tricyclic antidepressants confirm method
C0802218|T201|COMP|19321-9|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0802219|T201|COMP|19322-7|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0802220|T201|COMP|19323-5|LNC|6-Monoacetylmorphine cutoff|6-Monoacetylmorphine cutoff
C0802221|T201|COMP|19324-3|LNC|6-Monoacetylmorphine cutoff|6-Monoacetylmorphine cutoff
C0802222|T201|COMP|19325-0|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C0802223|T201|COMP|19326-8|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C0802224|T201|COMP|19328-4|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C0802225|T201|COMP|19329-2|LNC|Alpha hydroxyalprazolam cutoff|Alpha hydroxyalprazolam cutoff
C0802226|T201|COMP|19330-0|LNC|Alpha hydroxyalprazolam cutoff|Alpha hydroxyalprazolam cutoff
C0802227|T201|COMP|19331-8|LNC|Amitriptyline|Amitriptyline
C0802228|T201|COMP|19333-4|LNC|Amitriptyline cutoff|Amitriptyline cutoff
C0802229|T201|COMP|19334-2|LNC|Amitriptyline cutoff|Amitriptyline cutoff
C0802230|T201|COMP|19335-9|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C0802231|T201|COMP|19336-7|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C0802232|T201|COMP|19337-5|LNC|Amitriptyline+Nortriptyline cutoff|Amitriptyline+Nortriptyline cutoff
C0802233|T201|COMP|19338-3|LNC|Amitriptyline+Nortriptyline cutoff|Amitriptyline+Nortriptyline cutoff
C0802234|T201|COMP|19339-1|LNC|Amobarbital|Amobarbital
C0802235|T201|COMP|19341-7|LNC|Amobarbital cutoff|Amobarbital cutoff
C0802236|T201|COMP|19342-5|LNC|Amobarbital cutoff|Amobarbital cutoff
C0802237|T201|COMP|19343-3|LNC|Amphetamine|Amphetamine
C0802238|T201|COMP|19344-1|LNC|Amphetamine|Amphetamine
C0802239|T201|COMP|19346-6|LNC|Amphetamine|Amphetamine
C0802240|T201|COMP|19347-4|LNC|Amphetamine cutoff|Amphetamine cutoff
C0802241|T201|COMP|19348-2|LNC|Amphetamine cutoff|Amphetamine cutoff
C0802242|T201|COMP|19349-0|LNC|Aprobarbital|Aprobarbital
C0802243|T201|COMP|19350-8|LNC|Aprobarbital|Aprobarbital
C0802244|T201|COMP|19351-6|LNC|Aprobarbital cutoff|Aprobarbital cutoff
C0802245|T201|COMP|19352-4|LNC|Aprobarbital cutoff|Aprobarbital cutoff
C0802246|T201|COMP|19353-2|LNC|Barbital|Barbital
C0802247|T201|COMP|19354-0|LNC|Barbital|Barbital
C0802248|T201|COMP|19355-7|LNC|Barbital cutoff|Barbital cutoff
C0802249|T201|COMP|19356-5|LNC|Barbital cutoff|Barbital cutoff
C0802250|T201|COMP|19357-3|LNC|Benzoylecgonine cutoff|Benzoylecgonine cutoff
C0802251|T201|COMP|19358-1|LNC|Benzoylecgonine cutoff|Benzoylecgonine cutoff
C0802252|T201|COMP|19359-9|LNC|Cocaine|Cocaine
C0802253|T201|COMP|19360-7|LNC|Cocaine|Cocaine
C0802254|T201|COMP|3398-5|LNC|Cocaine|Cocaine
C0802255|T201|COMP|19362-3|LNC|Cocaine cutoff|Cocaine cutoff
C0802256|T201|COMP|19363-1|LNC|Cocaine cutoff|Cocaine cutoff
C0802257|T201|COMP|19364-9|LNC|Bromazepam|Bromazepam
C0802258|T201|COMP|19365-6|LNC|Bromazepam|Bromazepam
C0802259|T201|COMP|19366-4|LNC|Bromazepam cutoff|Bromazepam cutoff
C0802260|T201|COMP|19367-2|LNC|Bromazepam cutoff|Bromazepam cutoff
C0802261|T201|COMP|19368-0|LNC|Butabarbital|Butabarbital
C0802262|T201|COMP|19370-6|LNC|Butabarbital|Butabarbital
C0802263|T201|COMP|19371-4|LNC|Butabarbital cutoff|Butabarbital cutoff
C0802264|T201|COMP|19372-2|LNC|Butabarbital cutoff|Butabarbital cutoff
C0802265|T201|COMP|19373-0|LNC|Butalbital|Butalbital
C0802266|T201|COMP|19375-5|LNC|Butalbital cutoff|Butalbital cutoff
C0802267|T201|COMP|19376-3|LNC|Butalbital cutoff|Butalbital cutoff
C0802268|T201|COMP|19377-1|LNC|Butorphanol|Butorphanol
C0802269|T201|COMP|19378-9|LNC|Butorphanol|Butorphanol
C0802270|T201|COMP|19379-7|LNC|Butorphanol cutoff|Butorphanol cutoff
C0802271|T201|COMP|19380-5|LNC|Butorphanol cutoff|Butorphanol cutoff
C0802272|T201|COMP|19381-3|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0802273|T201|COMP|19382-1|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0802274|T201|COMP|19383-9|LNC|Carboxy tetrahydrocannabinol cutoff|Carboxy tetrahydrocannabinol cutoff
C0802275|T201|COMP|19384-7|LNC|Carboxy tetrahydrocannabinol cutoff|Carboxy tetrahydrocannabinol cutoff
C0802276|T201|COMP|19385-4|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0802277|T201|COMP|19386-2|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0802278|T201|COMP|19387-0|LNC|chlordiazePOXIDE cutoff|chlordiazePOXIDE cutoff
C0802279|T201|COMP|19388-8|LNC|chlordiazePOXIDE cutoff|chlordiazePOXIDE cutoff
C0802280|T201|COMP|19389-6|LNC|Chlorpheniramine|Chlorpheniramine
C0802281|T201|COMP|19391-2|LNC|Chlorpheniramine|Chlorpheniramine
C0802282|T201|COMP|19392-0|LNC|Chlorpheniramine|Chlorpheniramine
C0802283|T201|COMP|19393-8|LNC|Chlorpheniramine cutoff|Chlorpheniramine cutoff
C0802284|T201|COMP|19394-6|LNC|Chlorpheniramine cutoff|Chlorpheniramine cutoff
C0802285|T201|COMP|19395-3|LNC|chlorproMAZINE|chlorproMAZINE
C0802286|T201|COMP|19396-1|LNC|chlorproMAZINE|chlorproMAZINE
C0802287|T201|COMP|19397-9|LNC|chlorproMAZINE cutoff|chlorproMAZINE cutoff
C0802288|T201|COMP|19398-7|LNC|chlorproMAZINE cutoff|chlorproMAZINE cutoff
C0802289|T201|COMP|19399-5|LNC|clonazePAM|clonazePAM
C0802290|T201|COMP|19402-7|LNC|clonazePAM|clonazePAM
C0802291|T201|COMP|19403-5|LNC|clonazePAM cutoff|clonazePAM cutoff
C0802292|T201|COMP|19404-3|LNC|clonazePAM cutoff|clonazePAM cutoff
C0802293|T201|COMP|19405-0|LNC|Cocaethylene|Cocaethylene
C0802294|T201|COMP|19406-8|LNC|Cocaethylene|Cocaethylene
C0802295|T201|COMP|19408-4|LNC|Cocaethylene|Cocaethylene
C0802296|T201|COMP|19409-2|LNC|Cocaethylene cutoff|Cocaethylene cutoff
C0802297|T201|COMP|19410-0|LNC|Cocaethylene cutoff|Cocaethylene cutoff
C0802298|T201|COMP|19411-8|LNC|Codeine|Codeine
C0802299|T201|COMP|19413-4|LNC|Codeine cutoff|Codeine cutoff
C0802300|T201|COMP|19414-2|LNC|Codeine cutoff|Codeine cutoff
C0802301|T201|COMP|19415-9|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0802302|T201|COMP|19416-7|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0802303|T201|COMP|19417-5|LNC|Tetrahydrocannabinol cutoff|Tetrahydrocannabinol cutoff
C0802304|T201|COMP|19418-3|LNC|Tetrahydrocannabinol cutoff|Tetrahydrocannabinol cutoff
C0802305|T201|COMP|19419-1|LNC|Dextroamphetamine|Dextroamphetamine
C0802306|T201|COMP|19420-9|LNC|Dextroamphetamine|Dextroamphetamine
C0802307|T201|COMP|19421-7|LNC|Dextroamphetamine cutoff|Dextroamphetamine cutoff
C0802308|T201|COMP|19422-5|LNC|Dextroamphetamine cutoff|Dextroamphetamine cutoff
C0802309|T201|COMP|19423-3|LNC|Dextromethamphetamine|Dextromethamphetamine
C0802310|T201|COMP|19424-1|LNC|Dextromethamphetamine|Dextromethamphetamine
C0802311|T201|COMP|19425-8|LNC|Dextromethamphetamine|Dextromethamphetamine
C0802312|T201|COMP|12477-6|LNC|Dextromethamphetamine|Dextromethamphetamine
C0802313|T201|COMP|19427-4|LNC|Dextromethamphetamine cutoff|Dextromethamphetamine cutoff
C0802314|T201|COMP|19428-2|LNC|Dextromethamphetamine cutoff|Dextromethamphetamine cutoff
C0802315|T201|COMP|19429-0|LNC|Propoxyphene|Propoxyphene
C0802316|T201|COMP|19431-6|LNC|Propoxyphene cutoff|Propoxyphene cutoff
C0802317|T201|COMP|19432-4|LNC|Propoxyphene cutoff|Propoxyphene cutoff
C0802318|T201|COMP|19433-2|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C0802319|T201|COMP|19434-0|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C0802320|T201|COMP|19435-7|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C0802321|T201|COMP|19436-5|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C0802322|T201|COMP|19437-3|LNC|Propoxyphene+Norpropoxyphene cutoff|Propoxyphene+Norpropoxyphene cutoff
C0802323|T201|COMP|19438-1|LNC|Propoxyphene+Norpropoxyphene cutoff|Propoxyphene+Norpropoxyphene cutoff
C0802324|T201|COMP|19439-9|LNC|Diamorphine|Diamorphine
C0802325|T201|COMP|19441-5|LNC|Diamorphine cutoff|Diamorphine cutoff
C0802326|T201|COMP|19442-3|LNC|Diamorphine cutoff|Diamorphine cutoff
C0802327|T201|COMP|19443-1|LNC|diazePAM|diazePAM
C0802328|T201|COMP|19444-9|LNC|diazePAM cutoff|diazePAM cutoff
C0802329|T201|COMP|19445-6|LNC|diazePAM cutoff|diazePAM cutoff
C0802330|T201|COMP|19446-4|LNC|Dihydrocodeine|Dihydrocodeine
C0802331|T201|COMP|19448-0|LNC|Dihydrocodeine|Dihydrocodeine
C0802332|T201|COMP|19449-8|LNC|Dihydrocodeine|Dihydrocodeine
C0802333|T201|COMP|19450-6|LNC|Dihydrocodeine cutoff|Dihydrocodeine cutoff
C0802334|T201|COMP|19451-4|LNC|Dihydrocodeine cutoff|Dihydrocodeine cutoff
C0802335|T201|COMP|19452-2|LNC|Dimetamphetamine|Dimetamphetamine
C0802336|T201|COMP|19453-0|LNC|Dimetamphetamine|Dimetamphetamine
C0802337|T201|COMP|19454-8|LNC|Dimetamphetamine cutoff|Dimetamphetamine cutoff
C0802338|T201|COMP|19455-5|LNC|Dimetamphetamine cutoff|Dimetamphetamine cutoff
C0802339|T201|COMP|19456-3|LNC|Ethylamphetamine|Ethylamphetamine
C0802340|T201|COMP|19458-9|LNC|Ethylamphetamine|Ethylamphetamine
C0802341|T201|COMP|19459-7|LNC|Ethylamphetamine|Ethylamphetamine
C0802342|T201|COMP|19460-5|LNC|Ethylamphetamine cutoff|Ethylamphetamine cutoff
C0802343|T201|COMP|19461-3|LNC|Ethylamphetamine cutoff|Ethylamphetamine cutoff
C0802344|T201|COMP|19462-1|LNC|Ethylmorphine|Ethylmorphine
C0802345|T201|COMP|19463-9|LNC|Ethylmorphine|Ethylmorphine
C0802346|T201|COMP|19464-7|LNC|Ethylmorphine cutoff|Ethylmorphine cutoff
C0802347|T201|COMP|19465-4|LNC|Ethylmorphine cutoff|Ethylmorphine cutoff
C0802348|T201|COMP|19466-2|LNC|Flunitrazepam|Flunitrazepam
C0802349|T201|COMP|19467-0|LNC|Flunitrazepam|Flunitrazepam
C0802350|T201|COMP|19468-8|LNC|Flunitrazepam cutoff|Flunitrazepam cutoff
C0802351|T201|COMP|19469-6|LNC|Flunitrazepam cutoff|Flunitrazepam cutoff
C0802352|T201|COMP|19470-4|LNC|FLUoxetine|FLUoxetine
C0802353|T201|COMP|19471-2|LNC|FLUoxetine|FLUoxetine
C0802354|T201|COMP|19472-0|LNC|FLUoxetine cutoff|FLUoxetine cutoff
C0802355|T201|COMP|19473-8|LNC|FLUoxetine cutoff|FLUoxetine cutoff
C0802356|T201|COMP|19474-6|LNC|Flurazepam|Flurazepam
C0802357|T201|COMP|19475-3|LNC|Flurazepam|Flurazepam
C0802358|T201|COMP|19476-1|LNC|Flurazepam cutoff|Flurazepam cutoff
C0802359|T201|COMP|19477-9|LNC|Flurazepam cutoff|Flurazepam cutoff
C0802360|T201|COMP|19478-7|LNC|Haloperidol|Haloperidol
C0802361|T201|COMP|19479-5|LNC|Haloperidol|Haloperidol
C0802362|T201|COMP|19480-3|LNC|Haloperidol cutoff|Haloperidol cutoff
C0802363|T201|COMP|19481-1|LNC|Haloperidol cutoff|Haloperidol cutoff
C0802364|T201|COMP|19482-9|LNC|HYDROcodone|HYDROcodone
C0802365|T201|COMP|19483-7|LNC|HYDROcodone|HYDROcodone
C0802366|T201|COMP|19484-5|LNC|HYDROcodone cutoff|HYDROcodone cutoff
C0802367|T201|COMP|19485-2|LNC|HYDROcodone cutoff|HYDROcodone cutoff
C0802368|T201|COMP|19486-0|LNC|HYDROmorphone|HYDROmorphone
C0802369|T201|COMP|19487-8|LNC|HYDROmorphone cutoff|HYDROmorphone cutoff
C0802370|T201|COMP|19488-6|LNC|HYDROmorphone cutoff|HYDROmorphone cutoff
C0802371|T201|COMP|19489-4|LNC|Hydroxyalprazolam|Hydroxyalprazolam
C0802372|T201|COMP|19490-2|LNC|Hydroxyalprazolam|Hydroxyalprazolam
C0802373|T201|COMP|19491-0|LNC|Hydroxyalprazolam cutoff|Hydroxyalprazolam cutoff
C0802374|T201|COMP|19492-8|LNC|Hydroxyalprazolam cutoff|Hydroxyalprazolam cutoff
C0802375|T201|COMP|19493-6|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C0802376|T201|COMP|19494-4|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C0802377|T201|COMP|19495-1|LNC|Hydroxyethylflurazepam cutoff|Hydroxyethylflurazepam cutoff
C0802378|T201|COMP|19496-9|LNC|Hydroxyethylflurazepam cutoff|Hydroxyethylflurazepam cutoff
C0802379|T201|COMP|19497-7|LNC|Hydroxytriazolam|Hydroxytriazolam
C0802380|T201|COMP|19499-3|LNC|Ketamine|Ketamine
C0802381|T201|COMP|19500-8|LNC|Ketamine cutoff|Ketamine cutoff
C0802382|T201|COMP|19501-6|LNC|Ketamine cutoff|Ketamine cutoff
C0802383|T201|COMP|19502-4|LNC|Methotrimeprazine|Methotrimeprazine
C0802384|T201|COMP|19503-2|LNC|Methotrimeprazine|Methotrimeprazine
C0802385|T201|COMP|19504-0|LNC|Methotrimeprazine cutoff|Methotrimeprazine cutoff
C0802386|T201|COMP|19505-7|LNC|Methotrimeprazine cutoff|Methotrimeprazine cutoff
C0802387|T201|COMP|19506-5|LNC|Levomepromazine|Levomepromazine
C0802388|T201|COMP|19507-3|LNC|Levomepromazine|Levomepromazine
C0802389|T201|COMP|19508-1|LNC|Levomepromazine cutoff|Levomepromazine cutoff
C0802390|T201|COMP|19509-9|LNC|Levomepromazine cutoff|Levomepromazine cutoff
C0802391|T201|COMP|19510-7|LNC|Levomethamphetamine|Levomethamphetamine
C0802392|T201|COMP|19511-5|LNC|Levomethamphetamine|Levomethamphetamine
C0802393|T201|COMP|19512-3|LNC|Levomethamphetamine|Levomethamphetamine
C0802394|T201|COMP|19514-9|LNC|Levomethamphetamine cutoff|Levomethamphetamine cutoff
C0802395|T201|COMP|19515-6|LNC|Levomethamphetamine cutoff|Levomethamphetamine cutoff
C0802396|T201|COMP|19516-4|LNC|Levorphanol|Levorphanol
C0802397|T201|COMP|19518-0|LNC|Levorphanol cutoff|Levorphanol cutoff
C0802398|T201|COMP|19519-8|LNC|Levorphanol cutoff|Levorphanol cutoff
C0802399|T201|COMP|19520-6|LNC|LORazepam|LORazepam
C0802400|T201|COMP|19522-2|LNC|LORazepam cutoff|LORazepam cutoff
C0802401|T201|COMP|19523-0|LNC|LORazepam cutoff|LORazepam cutoff
C0802402|T201|COMP|19524-8|LNC|Lormetazepam|Lormetazepam
C0802403|T201|COMP|19525-5|LNC|Lormetazepam|Lormetazepam
C0802404|T201|COMP|19526-3|LNC|Lormetazepam cutoff|Lormetazepam cutoff
C0802405|T201|COMP|19527-1|LNC|Lormetazepam cutoff|Lormetazepam cutoff
C0802406|T201|COMP|19528-9|LNC|Lysergate diethylamide|Lysergate diethylamide
C0802407|T201|COMP|19530-5|LNC|Lysergate diethylamide cutoff|Lysergate diethylamide cutoff
C0802408|T201|COMP|19531-3|LNC|Lysergate diethylamide cutoff|Lysergate diethylamide cutoff
C0802409|T201|COMP|19532-1|LNC|Meperidine|Meperidine
C0802410|T201|COMP|19534-7|LNC|Meperidine cutoff|Meperidine cutoff
C0802411|T201|COMP|19535-4|LNC|Meperidine cutoff|Meperidine cutoff
C0802412|T201|COMP|19536-2|LNC|Mephobarbital|Mephobarbital
C0802413|T201|COMP|19537-0|LNC|Mephobarbital|Mephobarbital
C0802414|T201|COMP|19539-6|LNC|Mephobarbital|Mephobarbital
C0802415|T201|COMP|19540-4|LNC|Mephobarbital cutoff|Mephobarbital cutoff
C0802416|T201|COMP|19541-2|LNC|Mephobarbital cutoff|Mephobarbital cutoff
C0802417|T201|COMP|19542-0|LNC|Mescaline|Mescaline
C0802418|T201|COMP|19543-8|LNC|Mescaline|Mescaline
C0802419|T201|COMP|19544-6|LNC|Mescaline cutoff|Mescaline cutoff
C0802420|T201|COMP|19545-3|LNC|Mescaline cutoff|Mescaline cutoff
C0802421|T201|COMP|19546-1|LNC|Mesoridazine|Mesoridazine
C0802422|T201|COMP|19547-9|LNC|Mesoridazine|Mesoridazine
C0802423|T201|COMP|19548-7|LNC|Mesoridazine cutoff|Mesoridazine cutoff
C0802424|T201|COMP|19549-5|LNC|Mesoridazine cutoff|Mesoridazine cutoff
C0802425|T201|COMP|19550-3|LNC|Methadone|Methadone
C0802426|T201|COMP|19552-9|LNC|Methadone cutoff|Methadone cutoff
C0802427|T201|COMP|19553-7|LNC|Methadone cutoff|Methadone cutoff
C0802428|T201|COMP|19554-5|LNC|Methamphetamine|Methamphetamine
C0802429|T201|COMP|19555-2|LNC|Methamphetamine|Methamphetamine
C0802430|T201|COMP|19556-0|LNC|Methamphetamine cutoff|Methamphetamine cutoff
C0802431|T201|COMP|19557-8|LNC|Methamphetamine cutoff|Methamphetamine cutoff
C0802432|T201|COMP|19558-6|LNC|Methaqualone|Methaqualone
C0802433|T201|COMP|19559-4|LNC|Methaqualone cutoff|Methaqualone cutoff
C0802434|T201|COMP|19560-2|LNC|Methaqualone cutoff|Methaqualone cutoff
C0802435|T201|COMP|19561-0|LNC|Methylenediamine|Methylenediamine
C0802436|T201|COMP|19562-8|LNC|Methylenediamine|Methylenediamine
C0802437|T201|COMP|19563-6|LNC|Methylenediamine cutoff|Methylenediamine cutoff
C0802438|T201|COMP|19564-4|LNC|Methylenediamine cutoff|Methylenediamine cutoff
C0802439|T201|COMP|19565-1|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0802440|T201|COMP|19566-9|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0802441|T201|COMP|19567-7|LNC|Methylenedioxyamphetamine cutoff|Methylenedioxyamphetamine cutoff
C0802442|T201|COMP|19568-5|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0802443|T201|COMP|19569-3|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0802444|T201|COMP|19570-1|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0802445|T201|COMP|19571-9|LNC|Methylenedioxymethamphetamine cutoff|Methylenedioxymethamphetamine cutoff
C0802446|T201|COMP|19572-7|LNC|Methylenedioxymethamphetamine cutoff|Methylenedioxymethamphetamine cutoff
C0802447|T201|COMP|19573-5|LNC|MethylePHEDrine|MethylePHEDrine
C0802448|T201|COMP|19575-0|LNC|MethylePHEDrine cutoff|MethylePHEDrine cutoff
C0802449|T201|COMP|19576-8|LNC|MethylePHEDrine cutoff|MethylePHEDrine cutoff
C0802450|T201|COMP|19577-6|LNC|Methylphenidate|Methylphenidate
C0802451|T201|COMP|19578-4|LNC|Methylphenidate|Methylphenidate
C0802452|T201|COMP|19579-2|LNC|Methylphenidate cutoff|Methylphenidate cutoff
C0802453|T201|COMP|19580-0|LNC|Methylphenidate cutoff|Methylphenidate cutoff
C0802454|T201|COMP|19581-8|LNC|Methyprylon|Methyprylon
C0802455|T201|COMP|19583-4|LNC|Methyprylon cutoff|Methyprylon cutoff
C0802456|T201|COMP|19584-2|LNC|Methyprylon cutoff|Methyprylon cutoff
C0802457|T201|COMP|19585-9|LNC|Midazolam|Midazolam
C0802458|T201|COMP|19586-7|LNC|Midazolam|Midazolam
C0802459|T201|COMP|19588-3|LNC|Midazolam|Midazolam
C0802460|T201|COMP|19589-1|LNC|Midazolam cutoff|Midazolam cutoff
C0802461|T201|COMP|19590-9|LNC|Midazolam cutoff|Midazolam cutoff
C0802462|T201|COMP|19591-7|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0802463|T201|COMP|19592-5|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0802464|T201|COMP|19593-3|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0802465|T201|COMP|21050-0|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0802466|T201|COMP|19595-8|LNC|6-Monoacetylmorphine cutoff|6-Monoacetylmorphine cutoff
C0802467|T201|COMP|19596-6|LNC|6-Monoacetylmorphine cutoff|6-Monoacetylmorphine cutoff
C0802468|T201|COMP|19597-4|LNC|Morphine|Morphine
C0802469|T201|COMP|19599-0|LNC|Morphine cutoff|Morphine cutoff
C0802470|T201|COMP|19600-6|LNC|Morphine cutoff|Morphine cutoff
C0802471|T201|COMP|19601-4|LNC|Morphine.free|Morphine.free
C0802472|T201|COMP|19602-2|LNC|Morphine.free|Morphine.free
C0802473|T201|COMP|19603-0|LNC|Morphine.free cutoff|Morphine.free cutoff
C0802474|T201|COMP|19604-8|LNC|Morphine.free cutoff|Morphine.free cutoff
C0802475|T201|COMP|19605-5|LNC|Nalbuphine|Nalbuphine
C0802476|T201|COMP|19607-1|LNC|Nalbuphine cutoff|Nalbuphine cutoff
C0802477|T201|COMP|19608-9|LNC|Nalbuphine cutoff|Nalbuphine cutoff
C0802478|T201|COMP|19609-7|LNC|Naltrexone|Naltrexone
C0802479|T201|COMP|19610-5|LNC|Naltrexone|Naltrexone
C0802480|T201|COMP|19611-3|LNC|Naltrexone|Naltrexone
C0802481|T201|COMP|19612-1|LNC|Naltrexone cutoff|Naltrexone cutoff
C0802482|T201|COMP|19613-9|LNC|Naltrexone cutoff|Naltrexone cutoff
C0802483|T201|COMP|19614-7|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0802484|T201|COMP|19615-4|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0802485|T201|COMP|19617-0|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0802486|T201|COMP|19618-8|LNC|N-desalkylflurazepam cutoff|N-desalkylflurazepam cutoff
C0802487|T201|COMP|19619-6|LNC|N-desalkylflurazepam cutoff|N-desalkylflurazepam cutoff
C0802488|T201|COMP|19620-4|LNC|Nitrazepam|Nitrazepam
C0802489|T201|COMP|19621-2|LNC|Nitrazepam|Nitrazepam
C0802490|T201|COMP|19622-0|LNC|Nitrazepam cutoff|Nitrazepam cutoff
C0802491|T201|COMP|19623-8|LNC|Nitrazepam cutoff|Nitrazepam cutoff
C0802492|T201|COMP|19624-6|LNC|Nordiazepam|Nordiazepam
C0802493|T201|COMP|19626-1|LNC|Nordiazepam cutoff|Nordiazepam cutoff
C0802494|T201|COMP|19627-9|LNC|Nordiazepam cutoff|Nordiazepam cutoff
C0802495|T201|COMP|19628-7|LNC|Norfluoxetine|Norfluoxetine
C0802496|T201|COMP|19629-5|LNC|Norfluoxetine|Norfluoxetine
C0802497|T201|COMP|19630-3|LNC|Norfluoxetine cutoff|Norfluoxetine cutoff
C0802498|T201|COMP|19631-1|LNC|Norfluoxetine cutoff|Norfluoxetine cutoff
C0802499|T201|COMP|19632-9|LNC|Norpropoxyphene|Norpropoxyphene
C0802500|T201|COMP|19635-2|LNC|Norpropoxyphene|Norpropoxyphene
C0802501|T201|COMP|19636-0|LNC|Norpropoxyphene cutoff|Norpropoxyphene cutoff
C0802502|T201|COMP|19637-8|LNC|Norpropoxyphene cutoff|Norpropoxyphene cutoff
C0802503|T201|COMP|19638-6|LNC|Oxazepam|Oxazepam
C0802504|T201|COMP|19639-4|LNC|Oxazepam|Oxazepam
C0802505|T201|COMP|19640-2|LNC|Oxazepam cutoff|Oxazepam cutoff
C0802506|T201|COMP|19641-0|LNC|Oxazepam cutoff|Oxazepam cutoff
C0802507|T201|COMP|19642-8|LNC|oxyCODONE|oxyCODONE
C0802508|T201|COMP|19643-6|LNC|oxyCODONE|oxyCODONE
C0802509|T201|COMP|19644-4|LNC|oxyCODONE cutoff|oxyCODONE cutoff
C0802510|T201|COMP|19645-1|LNC|oxyCODONE cutoff|oxyCODONE cutoff
C0802511|T201|COMP|19646-9|LNC|oxyMORphone|oxyMORphone
C0802512|T201|COMP|19648-5|LNC|oxyMORphone|oxyMORphone
C0802513|T201|COMP|19649-3|LNC|oxyMORphone cutoff|oxyMORphone cutoff
C0802514|T201|COMP|19650-1|LNC|oxyMORphone cutoff|oxyMORphone cutoff
C0802515|T201|COMP|19651-9|LNC|Para hydroxyamphetamine|Para hydroxyamphetamine
C0802516|T201|COMP|19652-7|LNC|Para hydroxyamphetamine|Para hydroxyamphetamine
C0802517|T201|COMP|19653-5|LNC|Para hydroxyamphetamine cutoff|Para hydroxyamphetamine cutoff
C0802518|T201|COMP|19654-3|LNC|Para hydroxyamphetamine cutoff|Para hydroxyamphetamine cutoff
C0802519|T201|COMP|19655-0|LNC|PENTobarbital|PENTobarbital
C0802520|T201|COMP|19657-6|LNC|PENTobarbital cutoff|PENTobarbital cutoff
C0802521|T201|COMP|19658-4|LNC|PENTobarbital cutoff|PENTobarbital cutoff
C0802522|T201|COMP|19659-2|LNC|Phencyclidine|Phencyclidine
C0802523|T201|COMP|19660-0|LNC|Phencyclidine cutoff|Phencyclidine cutoff
C0802524|T201|COMP|19661-8|LNC|Phencyclidine cutoff|Phencyclidine cutoff
C0802525|T201|COMP|19662-6|LNC|Phenmetrazine|Phenmetrazine
C0802526|T201|COMP|19664-2|LNC|Phenmetrazine cutoff|Phenmetrazine cutoff
C0802527|T201|COMP|19665-9|LNC|Phenmetrazine cutoff|Phenmetrazine cutoff
C0802528|T201|COMP|19666-7|LNC|PHENobarbital|PHENobarbital
C0802529|T201|COMP|19668-3|LNC|PHENobarbital cutoff|PHENobarbital cutoff
C0802530|T201|COMP|19669-1|LNC|PHENobarbital cutoff|PHENobarbital cutoff
C0802531|T201|COMP|19670-9|LNC|Phenothiazines|Phenothiazines
C0802532|T201|COMP|19672-5|LNC|Phenothiazines cutoff|Phenothiazines cutoff
C0802533|T201|COMP|19673-3|LNC|Phenothiazines cutoff|Phenothiazines cutoff
C0802534|T201|COMP|19674-1|LNC|Phentermine|Phentermine
C0802535|T201|COMP|19676-6|LNC|Phentermine cutoff|Phentermine cutoff
C0802536|T201|COMP|19677-4|LNC|Phentermine cutoff|Phentermine cutoff
C0802537|T201|COMP|19678-2|LNC|Prazepam|Prazepam
C0802538|T201|COMP|19679-0|LNC|Prazepam|Prazepam
C0802539|T201|COMP|19680-8|LNC|Prazepam cutoff|Prazepam cutoff
C0802540|T201|COMP|19681-6|LNC|Prazepam cutoff|Prazepam cutoff
C0802541|T201|COMP|19682-4|LNC|Psilocin|Psilocin
C0802542|T201|COMP|19683-2|LNC|Psilocin|Psilocin
C0802543|T201|COMP|19684-0|LNC|Psilocin cutoff|Psilocin cutoff
C0802544|T201|COMP|19685-7|LNC|Psilocin cutoff|Psilocin cutoff
C0802545|T201|COMP|19686-5|LNC|Psilocybin|Psilocybin
C0802546|T201|COMP|19687-3|LNC|Psilocybin|Psilocybin
C0802547|T201|COMP|19688-1|LNC|Psilocybin|Psilocybin
C0802548|T201|COMP|6930-2|LNC|Psilocybin|Psilocybin
C0802549|T201|COMP|19690-7|LNC|Psilocybin cutoff|Psilocybin cutoff
C0802550|T201|COMP|19691-5|LNC|Psilocybin cutoff|Psilocybin cutoff
C0802551|T201|COMP|19692-3|LNC|Secobarbital|Secobarbital
C0802552|T201|COMP|19695-6|LNC|Secobarbital|Secobarbital
C0802553|T201|COMP|19696-4|LNC|Secobarbital cutoff|Secobarbital cutoff
C0802554|T201|COMP|19697-2|LNC|Secobarbital cutoff|Secobarbital cutoff
C0802555|T201|COMP|19698-0|LNC|Temazepam|Temazepam
C0802556|T201|COMP|19700-4|LNC|Temazepam cutoff|Temazepam cutoff
C0802557|T201|COMP|19701-2|LNC|Temazepam cutoff|Temazepam cutoff
C0802558|T201|COMP|19702-0|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0802559|T201|COMP|19703-8|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0802560|T201|COMP|19704-6|LNC|Tetrahydrocannabinol cutoff|Tetrahydrocannabinol cutoff
C0802561|T201|COMP|19705-3|LNC|Tetrahydrocannabinol cutoff|Tetrahydrocannabinol cutoff
C0802562|T201|COMP|19706-1|LNC|Thioridazine|Thioridazine
C0802563|T201|COMP|19707-9|LNC|Thioridazine|Thioridazine
C0802564|T201|COMP|19708-7|LNC|Thioridazine cutoff|Thioridazine cutoff
C0802565|T201|COMP|19709-5|LNC|Thioridazine cutoff|Thioridazine cutoff
C0802566|T201|COMP|19710-3|LNC|traMADol|traMADol
C0802567|T201|COMP|19712-9|LNC|traMADol cutoff|traMADol cutoff
C0802568|T201|COMP|19713-7|LNC|traMADol cutoff|traMADol cutoff
C0802569|T201|COMP|19714-5|LNC|Triazolam|Triazolam
C0802570|T201|COMP|19716-0|LNC|Triazolam cutoff|Triazolam cutoff
C0802571|T201|COMP|19717-8|LNC|Triazolam cutoff|Triazolam cutoff
C0802572|T201|COMP|19718-6|LNC|Trichlorothiazide|Trichlorothiazide
C0802573|T201|COMP|19719-4|LNC|Trichlorothiazide|Trichlorothiazide
C0802574|T201|COMP|19720-2|LNC|Trichlorothiazide|Trichlorothiazide
C0802575|T201|COMP|19721-0|LNC|Trichlorothiazide|Trichlorothiazide
C0802576|T201|COMP|19722-8|LNC|Trichlorothiazide cutoff|Trichlorothiazide cutoff
C0802577|T201|COMP|19723-6|LNC|Trichlorothiazide cutoff|Trichlorothiazide cutoff
C0802578|T201|COMP|19762-4|LNC|General categories|General categories
C0802579|T201|COMP|19763-2|LNC|Specimen source|Specimen source
C0802580|T201|COMP|19764-0|LNC|Statement of adequacy|Statement of adequacy
C0802583|T201|COMP|19767-3|LNC|Cytologist|Cytologist
C0802584|T201|COMP|19768-1|LNC|Reviewing cytologist|Reviewing cytologist
C0802585|T201|COMP|19769-9|LNC|Pathologist|Pathologist
C0802586|T201|COMP|19771-5|LNC|Screen techniques|Screen techniques
C0802587|T201|COMP|19772-3|LNC|Preparation techniques|Preparation techniques
C0802588|T201|COMP|19773-1|LNC|Recommended follow-up|Recommended follow-up
C0802589|T201|COMP|19774-9|LNC|Cytology study comment|Cytology study comment
C0803188|T201|COMP|20373-7|LNC|Amikacin|Amikacin
C0803189|T201|COMP|20374-5|LNC|Ampicillin+Sulbactam|Ampicillin+Sulbactam
C0803190|T201|COMP|20375-2|LNC|Clarithromycin|Clarithromycin
C0803191|T201|COMP|20376-0|LNC|Clofazimine|Clofazimine
C0803192|T201|COMP|20377-8|LNC|Ciprofloxacin|Ciprofloxacin
C0803193|T201|COMP|20378-6|LNC|Ceftizoxime|Ceftizoxime
C0803194|T201|COMP|20379-4|LNC|Doxycycline|Doxycycline
C0803195|T201|COMP|20380-2|LNC|Erythromycin|Erythromycin
C0803196|T201|COMP|20381-0|LNC|Ethambutol|Ethambutol
C0803197|T201|COMP|20382-8|LNC|Ethionamide|Ethionamide
C0803198|T201|COMP|20383-6|LNC|Isoniazid|Isoniazid
C0803199|T201|COMP|20384-4|LNC|Ofloxacin|Ofloxacin
C0803200|T201|COMP|20385-1|LNC|rifAMPin|rifAMPin
C0803201|T201|COMP|20386-9|LNC|Rifabutin|Rifabutin
C0803202|T201|COMP|20387-7|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0803203|T201|COMP|20388-5|LNC|Nitrofurazone|Nitrofurazone
C0803204|T201|COMP|20389-3|LNC|Mupirocin|Mupirocin
C0803205|T201|COMP|20390-1|LNC|Silver sulfADIAZINE|Silver sulfADIAZINE
C0803206|T201|COMP|20391-9|LNC|Mafenide|Mafenide
C0803207|T201|COMP|20392-7|LNC|Sample icteric|Sample icteric
C0803208|T201|COMP|20393-5|LNC|Sample hemolyzed|Sample hemolyzed
C0803209|T201|COMP|20394-3|LNC|Sample lipemic|Sample lipemic
C0803210|T201|COMP|20395-0|LNC|Sample integrity|Sample integrity
C0803211|T201|COMP|20396-8|LNC|levoFLOXacin|levoFLOXacin
C0803212|T201|COMP|20397-6|LNC|Sparfloxacin|Sparfloxacin
C0803213|T201|COMP|20398-4|LNC|Nuclear Ab pattern.homogeneous|Nuclear Ab pattern.homogeneous
C0803214|T201|COMP|20399-2|LNC|Nuclear Ab pattern.nucleolar|Nuclear Ab pattern.nucleolar
C0803215|T201|COMP|20400-8|LNC|Nuclear Ab pattern.rim|Nuclear Ab pattern.rim
C0803216|T201|COMP|20401-6|LNC|Nuclear Ab pattern.speckled|Nuclear Ab pattern.speckled
C0803217|T201|COMP|20402-4|LNC|Cells.CD16+CD56+|Cells.CD16+CD56+
C0803218|T201|COMP|20403-2|LNC|Fibronectin.fetal|Fibronectin.fetal
C0803219|T201|COMP|20404-0|LNC|Fibronectin.fetal|Fibronectin.fetal
C0803220|T201|COMP|20405-7|LNC|Urobilinogen|Urobilinogen
C0803221|T201|COMP|20406-5|LNC|Glucose|Glucose
C0803222|T201|COMP|20407-3|LNC|Nitrite|Nitrite
C0803223|T201|COMP|20408-1|LNC|Leukocytes|Leukocytes
C0803224|T201|COMP|20409-9|LNC|Erythrocytes|Erythrocytes
C0803225|T201|COMP|20410-7|LNC|Amphetamines|Amphetamines
C0803226|T201|COMP|20411-5|LNC|Barbiturates|Barbiturates
C0803227|T201|COMP|20412-3|LNC|Benzodiazepines|Benzodiazepines
C0803228|T201|COMP|20413-1|LNC|Cannabinoids|Cannabinoids
C0803229|T201|COMP|20414-9|LNC|Thiazides|Thiazides
C0803230|T201|COMP|20415-6|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0803231|T201|COMP|20416-4|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C0803232|T201|COMP|20417-2|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C0803233|T201|COMP|20418-0|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C0803234|T201|COMP|20419-8|LNC|Lutropin|Lutropin
C0803235|T201|COMP|20420-6|LNC|Acid phosphatase.prostatic|Acid phosphatase.prostatic
C0803236|T201|COMP|20421-4|LNC|Barbiturates|Barbiturates
C0803237|T201|COMP|1825-9|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C0803238|T201|COMP|20423-0|LNC|Beta lactamase organism identified|Beta lactamase organism identified
C0803239|T201|COMP|20424-8|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C0803240|T201|COMP|20425-5|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C0803241|T201|COMP|20426-3|LNC|Alkaline phosphatase.bile|Alkaline phosphatase.bile
C0803242|T201|COMP|20427-1|LNC|Acetylcholine receptor Ab|Acetylcholine receptor Ab
C0803243|T201|COMP|20428-9|LNC|Phospholipid Ab.IgG|Phospholipid Ab.IgG
C0803244|T201|COMP|20429-7|LNC|Phospholipid Ab.IgM|Phospholipid Ab.IgM
C0803245|T201|COMP|20430-5|LNC|Culture medium|Culture medium
C0803247|T201|COMP|20432-1|LNC|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C0803248|T201|COMP|20433-9|LNC|Follitropin|Follitropin
C0803249|T201|COMP|20434-7|LNC|Prolactin|Prolactin
C0803250|T201|COMP|20435-4|LNC|Unidentified extractable nuclear Ab|Unidentified extractable nuclear Ab
C0803251|T201|COMP|20436-2|LNC|Glucose^2H post dose glucose|Glucose^2H post dose glucose
C0803252|T201|COMP|20437-0|LNC|Glucose^3H post dose glucose|Glucose^3H post dose glucose
C0803253|T201|COMP|20438-8|LNC|Glucose^1H post dose glucose|Glucose^1H post dose glucose
C0803254|T201|COMP|20439-6|LNC|Glucose^30M post dose glucose|Glucose^30M post dose glucose
C0803255|T201|COMP|20440-4|LNC|Glucose^1.5H post dose glucose|Glucose^1.5H post dose glucose
C0803256|T201|COMP|20441-2|LNC|Glucose^post 50 g glucose|Glucose^post 50 g glucose
C0803257|T201|COMP|20442-0|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C0803258|T201|COMP|20444-6|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C0803259|T201|COMP|20445-3|LNC|Herpes virus identified|Herpes virus identified
C0803260|T201|COMP|20446-1|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C0803261|T201|COMP|20447-9|LNC|HIV 1 RNA|HIV 1 RNA
C0803262|T201|COMP|20448-7|LNC|Insulin|Insulin
C0803263|T201|COMP|20449-5|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0803264|T201|COMP|20450-3|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0803265|T201|COMP|20451-1|LNC|Thyroxine|Thyroxine
C0803266|T201|COMP|20452-9|LNC|Thyrotropin|Thyrotropin
C0803267|T201|COMP|20453-7|LNC|Epithelial cells|Epithelial cells
C0803268|T201|COMP|20454-5|LNC|Protein|Protein
C0803269|T201|COMP|20455-2|LNC|Leukocytes|Leukocytes
C0803270|T201|COMP|20456-0|LNC|Fungi.yeastlike|Fungi.yeastlike
C0803271|T201|COMP|20457-8|LNC|Fungi.filamentous|Fungi.filamentous
C0803272|T201|COMP|20458-6|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0803273|T201|COMP|20459-4|LNC|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C0803274|T201|COMP|20460-2|LNC|Cefuroxime.oral|Cefuroxime.oral
C0803275|T201|COMP|20461-0|LNC|Pyrazinamide|Pyrazinamide
C0803276|T201|COMP|20462-8|LNC|Streptomycin|Streptomycin
C0803277|T201|COMP|20463-6|LNC|Mycobacterium avium complex rRNA|Mycobacterium avium complex rRNA
C0803278|T201|COMP|20464-4|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C0803279|T201|COMP|20465-1|LNC|Choriogonadotropin|Choriogonadotropin
C0803280|T201|COMP|20466-9|LNC|Estriol.unconjugated|Estriol.unconjugated
C0803281|T201|COMP|20467-7|LNC|Blood bank alert|Blood bank alert
C0803282|T201|COMP|20468-5|LNC|Thiamine|Thiamine
C0803283|T201|COMP|20469-3|LNC|Acetone|Acetone
C0803284|T201|COMP|20470-1|LNC|Ethanol|Ethanol
C0803285|T201|COMP|20471-9|LNC|Isopropanol|Isopropanol
C0803286|T201|COMP|20472-7|LNC|Eosinophils|Eosinophils
C0803287|T201|COMP|20473-5|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C0803288|T201|COMP|20474-3|LNC|Bacteria identified|Bacteria identified
C0803289|T201|COMP|20475-0|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0803290|T201|COMP|20476-8|LNC|Cells.CD1a/100 cells|Cells.CD1a/100 cells
C0803291|T201|COMP|20477-6|LNC|Cells.CD33+CD44+/100 cells|Cells.CD33+CD44+/100 cells
C0803292|T201|COMP|20478-4|LNC|Cells.CD61/100 cells|Cells.CD61/100 cells
C0803293|T201|COMP|20479-2|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0803294|T201|COMP|20482-6|LNC|Granulocytes|Granulocytes
C0803295|T201|COMP|20483-4|LNC|Mitochondria Ab|Mitochondria Ab
C0803296|T201|COMP|20484-2|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C0803297|T201|COMP|20485-9|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C0803298|T201|COMP|20486-7|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C0803299|T201|COMP|20487-5|LNC|Neisseria meningitidis serogroups A+Y Ag|Neisseria meningitidis serogroups A+Y Ag
C0803300|T201|COMP|20488-3|LNC|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C0803301|T201|COMP|20489-1|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C0803302|T201|COMP|20490-9|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0803303|T201|COMP|20491-7|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0803304|T201|COMP|20492-5|LNC|Hemoglobin pattern imp|Hemoglobin pattern imp
C0803305|T201|COMP|20493-3|LNC|Histiocytes/100 cells|Histiocytes/100 cells
C0803306|T201|COMP|20495-8|LNC|Gliadin Ab.IgA|Gliadin Ab.IgA
C0803307|T201|COMP|20496-6|LNC|Gliadin Ab.IgG|Gliadin Ab.IgG
C0803308|T201|COMP|20497-4|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C0803309|T201|COMP|20498-2|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C0803310|T201|COMP|20499-0|LNC|Phosphatidylglycerol/Surfactant.total|Phosphatidylglycerol/Surfactant.total
C0803311|T201|COMP|20500-5|LNC|Hydroxyalprazolam|Hydroxyalprazolam
C0803312|T201|COMP|20501-3|LNC|Hydroxytriazolam|Hydroxytriazolam
C0803313|T201|COMP|20502-1|LNC|Clue cells|Clue cells
C0803314|T201|COMP|20503-9|LNC|Cells.CD22+CD11c+/100 cells|Cells.CD22+CD11c+/100 cells
C0803315|T201|COMP|20504-7|LNC|Histiocytes/100 cells|Histiocytes/100 cells
C0803316|T201|COMP|20505-4|LNC|Bilirubin|Bilirubin
C0803317|T201|COMP|20506-2|LNC|Specimen drawn from|Specimen drawn from
C0803318|T201|COMP|20507-0|LNC|Reagin Ab|Reagin Ab
C0803319|T201|COMP|20508-8|LNC|Reagin Ab|Reagin Ab
C0803320|T201|COMP|20509-6|LNC|Hemoglobin|Hemoglobin
C0803321|T201|COMP|20510-4|LNC|Lipoprotein pattern|Lipoprotein pattern
C0803322|T201|COMP|20511-2|LNC|Creatinine|Creatinine
C0803323|T201|COMP|20512-0|LNC|Turbidity|Turbidity
C0803324|T201|COMP|20513-8|LNC|Turbidity|Turbidity
C0803325|T201|COMP|20514-6|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0803326|T201|COMP|20515-3|LNC|Amitriptyline|Amitriptyline
C0803327|T201|COMP|20516-1|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C0803328|T201|COMP|20517-9|LNC|Aprobarbital|Aprobarbital
C0803329|T201|COMP|20518-7|LNC|Barbital|Barbital
C0803330|T201|COMP|20519-5|LNC|Cocaine|Cocaine
C0803331|T201|COMP|20520-3|LNC|Bromazepam|Bromazepam
C0803332|T201|COMP|20521-1|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0803333|T201|COMP|20522-9|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0803334|T201|COMP|20523-7|LNC|chlorproMAZINE|chlorproMAZINE
C0803335|T201|COMP|20524-5|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0803336|T201|COMP|20525-2|LNC|Dextroamphetamine|Dextroamphetamine
C0803337|T201|COMP|20526-0|LNC|Dimetamphetamine|Dimetamphetamine
C0803338|T201|COMP|20527-8|LNC|Ethylmorphine|Ethylmorphine
C0803339|T201|COMP|20528-6|LNC|Flunitrazepam|Flunitrazepam
C0803340|T201|COMP|20529-4|LNC|FLUoxetine|FLUoxetine
C0803341|T201|COMP|20530-2|LNC|Haloperidol|Haloperidol
C0803342|T201|COMP|20532-8|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C0803343|T201|COMP|20533-6|LNC|Hydroxytriazolam|Hydroxytriazolam
C0803344|T201|COMP|20535-1|LNC|Hydroxytriazolam cutoff|Hydroxytriazolam cutoff
C0803345|T201|COMP|20536-9|LNC|Hydroxytriazolam cutoff|Hydroxytriazolam cutoff
C0803346|T201|COMP|20537-7|LNC|Ketamine|Ketamine
C0803347|T201|COMP|20538-5|LNC|Methotrimeprazine|Methotrimeprazine
C0803348|T201|COMP|20539-3|LNC|Levomepromazine|Levomepromazine
C0803349|T201|COMP|20540-1|LNC|Levorphanol|Levorphanol
C0803350|T201|COMP|20541-9|LNC|Lormetazepam|Lormetazepam
C0803351|T201|COMP|20542-7|LNC|Lysergate diethylamide|Lysergate diethylamide
C0803352|T201|COMP|20543-5|LNC|Mescaline|Mescaline
C0803353|T201|COMP|20544-3|LNC|Mesoridazine|Mesoridazine
C0803354|T201|COMP|20545-0|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0803355|T201|COMP|20546-8|LNC|Methylenedioxyamphetamine cutoff|Methylenedioxyamphetamine cutoff
C0803356|T201|COMP|20547-6|LNC|MethylePHEDrine|MethylePHEDrine
C0803357|T201|COMP|20548-4|LNC|Methylphenidate|Methylphenidate
C0803358|T201|COMP|20549-2|LNC|Methyprylon|Methyprylon
C0803359|T201|COMP|20550-0|LNC|Morphine.free|Morphine.free
C0803360|T201|COMP|20551-8|LNC|Nalbuphine|Nalbuphine
C0803361|T201|COMP|20552-6|LNC|Nitrazepam|Nitrazepam
C0803362|T201|COMP|20553-4|LNC|Norfluoxetine|Norfluoxetine
C0803363|T201|COMP|20554-2|LNC|Para hydroxyamphetamine|Para hydroxyamphetamine
C0803364|T201|COMP|20555-9|LNC|Phenmetrazine|Phenmetrazine
C0803365|T201|COMP|20556-7|LNC|Phenothiazines|Phenothiazines
C0803366|T201|COMP|20557-5|LNC|Phentermine|Phentermine
C0803367|T201|COMP|20558-3|LNC|Psilocin|Psilocin
C0803368|T201|COMP|20559-1|LNC|Temazepam|Temazepam
C0803369|T201|COMP|20560-9|LNC|Thioridazine|Thioridazine
C0803370|T201|COMP|20561-7|LNC|traMADol|traMADol
C0803372|T201|COMP|20563-3|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C0803374|T201|COMP|20565-8|LNC|Carbon dioxide|Carbon dioxide
C0803375|T201|COMP|20566-6|LNC|Colony count|Colony count
C0803376|T201|COMP|20567-4|LNC|Ferritin|Ferritin
C0803377|T201|COMP|20568-2|LNC|Prolactin|Prolactin
C0803378|T201|COMP|20569-0|LNC|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C0803379|T201|COMP|20570-8|LNC|Hematocrit|Hematocrit
C0803380|T201|COMP|20571-6|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C0803381|T201|COMP|20572-4|LNC|Hemoglobin A/Hemoglobin.total|Hemoglobin A/Hemoglobin.total
C0803382|T201|COMP|20573-2|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C0803383|T201|COMP|20574-0|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C0803384|T201|COMP|20575-7|LNC|Hepatitis A virus Ab|Hepatitis A virus Ab
C0803385|T201|COMP|20576-5|LNC|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C0803386|T201|COMP|20577-3|LNC|Protein|Protein
C0803387|T201|COMP|20578-1|LNC|Vancomycin|Vancomycin
C0803388|T201|COMP|20579-9|LNC|Methanol|Methanol
C0803389|T201|COMP|20584-9|LNC|Leukocytes|Leukocytes
C0803390|T201|COMP|20585-6|LNC|Lymphocytes|Lymphocytes
C0803391|T201|COMP|20586-4|LNC|Cells.CD1/100 cells|Cells.CD1/100 cells
C0803392|T201|COMP|20587-2|LNC|Cells.CD10/100 cells|Cells.CD10/100 cells
C0803393|T201|COMP|20588-0|LNC|Cells.CD13/100 cells|Cells.CD13/100 cells
C0803394|T201|COMP|20589-8|LNC|Cells.CD14/100 cells|Cells.CD14/100 cells
C0803395|T201|COMP|20590-6|LNC|Cells.CD15/100 cells|Cells.CD15/100 cells
C0803396|T201|COMP|20591-4|LNC|Cells.CD16+CD57-/100 cells|Cells.CD16+CD57-/100 cells
C0803397|T201|COMP|20592-2|LNC|Cells.CD19|Cells.CD19
C0803398|T201|COMP|20593-0|LNC|Cells.CD19/100 cells|Cells.CD19/100 cells
C0803399|T201|COMP|20594-8|LNC|Cells.CD2/100 cells|Cells.CD2/100 cells
C0803400|T201|COMP|20595-5|LNC|Cells.CD20/100 cells|Cells.CD20/100 cells
C0803401|T201|COMP|20596-3|LNC|Cells.CD22/100 cells|Cells.CD22/100 cells
C0803402|T201|COMP|20597-1|LNC|Cells.CD24/100 cells|Cells.CD24/100 cells
C0803403|T201|COMP|20598-9|LNC|Cells.CD3|Cells.CD3
C0803404|T201|COMP|20599-7|LNC|Cells.CD3/100 cells|Cells.CD3/100 cells
C0803405|T201|COMP|20600-3|LNC|Cells.CD30/100 cells|Cells.CD30/100 cells
C0803406|T201|COMP|20601-1|LNC|Cells.CD33/100 cells|Cells.CD33/100 cells
C0803407|T201|COMP|20602-9|LNC|Cells.CD34/100 cells|Cells.CD34/100 cells
C0803408|T201|COMP|20603-7|LNC|Cells.CD38/100 cells|Cells.CD38/100 cells
C0803409|T201|COMP|20604-5|LNC|Cells.CD3-CD16+CD56+|Cells.CD3-CD16+CD56+
C0803410|T201|COMP|20605-2|LNC|Cells.CD4|Cells.CD4
C0803411|T201|COMP|20606-0|LNC|Cells.CD4/100 cells|Cells.CD4/100 cells
C0803412|T201|COMP|20607-8|LNC|Cells.CD3+CD4+/Cells.CD3+CD8+|Cells.CD3+CD4+/Cells.CD3+CD8+
C0803413|T201|COMP|20608-6|LNC|Cells.CD41/100 cells|Cells.CD41/100 cells
C0803414|T201|COMP|20609-4|LNC|Cells.CD42/100 cells|Cells.CD42/100 cells
C0803415|T201|COMP|20610-2|LNC|Cells.CD45/100 cells|Cells.CD45/100 cells
C0803416|T201|COMP|20611-0|LNC|Cells.CD5/100 cells|Cells.CD5/100 cells
C0803417|T201|COMP|20612-8|LNC|Cells.CD7/100 cells|Cells.CD7/100 cells
C0803418|T201|COMP|20613-6|LNC|Cells.CD8|Cells.CD8
C0803419|T201|COMP|20614-4|LNC|Cells.CD8/100 cells|Cells.CD8/100 cells
C0803420|T201|COMP|20615-1|LNC|Lymphocytes.IgD/100 lymphocytes|Lymphocytes.IgD/100 lymphocytes
C0803421|T201|COMP|20616-9|LNC|Lymphocytes.IgM/100 lymphocytes|Lymphocytes.IgM/100 lymphocytes
C0803422|T201|COMP|20617-7|LNC|Lymphocytes.kappa/100 lymphocytes|Lymphocytes.kappa/100 lymphocytes
C0803423|T201|COMP|20618-5|LNC|Lymphocytes.lambda/100 lymphocytes|Lymphocytes.lambda/100 lymphocytes
C0803424|T201|COMP|20619-3|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0803425|T201|COMP|20620-1|LNC|Cells.CD16+CD56+/100 cells|Cells.CD16+CD56+/100 cells
C0803426|T201|COMP|20621-9|LNC|Albumin/Creatinine|Albumin/Creatinine
C0803427|T201|COMP|20622-7|LNC|Cortisol|Cortisol
C0803428|T201|COMP|20623-5|LNC|Coproporphyrin|Coproporphyrin
C0803429|T201|COMP|20624-3|LNC|Creatinine|Creatinine
C0803430|T201|COMP|20625-0|LNC|Lead|Lead
C0803431|T201|COMP|20626-8|LNC|Reducing substances|Reducing substances
C0803432|T201|COMP|20627-6|LNC|Turbidity|Turbidity
C0803434|T201|COMP|20629-2|LNC|levoFLOXacin|levoFLOXacin
C0803437|T201|COMP|20633-4|LNC|1-Methylhistidine|1-Methylhistidine
C0803438|T201|COMP|20634-2|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0803439|T201|COMP|20635-9|LNC|3-Methylhistidine|3-Methylhistidine
C0803440|T201|COMP|20636-7|LNC|Alanine|Alanine
C0803441|T201|COMP|20637-5|LNC|Arginine|Arginine
C0803442|T201|COMP|20638-3|LNC|Asparagine|Asparagine
C0803443|T201|COMP|20639-1|LNC|Aspartate|Aspartate
C0803444|T201|COMP|20640-9|LNC|Citrulline|Citrulline
C0803445|T201|COMP|20641-7|LNC|Cysteine|Cysteine
C0803447|T201|COMP|20643-3|LNC|Glutamine|Glutamine
C0803448|T201|COMP|20644-1|LNC|Glycine|Glycine
C0803449|T201|COMP|20645-8|LNC|Histidine|Histidine
C0803451|T201|COMP|20647-4|LNC|Hydroxyproline|Hydroxyproline
C0803452|T201|COMP|20648-2|LNC|Isoleucine|Isoleucine
C0803453|T201|COMP|20649-0|LNC|Leucine|Leucine
C0803454|T201|COMP|20650-8|LNC|Lysine|Lysine
C0803455|T201|COMP|20651-6|LNC|Methionine|Methionine
C0803456|T201|COMP|20652-4|LNC|Ornithine|Ornithine
C0803457|T201|COMP|20654-0|LNC|Phosphoserine|Phosphoserine
C0803458|T201|COMP|20655-7|LNC|Proline|Proline
C0803459|T201|COMP|20656-5|LNC|Serine|Serine
C0803460|T201|COMP|20657-3|LNC|Taurine|Taurine
C0803461|T201|COMP|20658-1|LNC|Threonine|Threonine
C0803463|T201|COMP|20660-7|LNC|Tyrosine|Tyrosine
C0803464|T201|COMP|20661-5|LNC|Valine|Valine
C0803465|T201|COMP|20662-3|LNC|Allergens tested for|Allergens tested for
C0803466|T201|COMP|20663-1|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0803467|T201|COMP|20664-9|LNC|Barbiturates|Barbiturates
C0803468|T201|COMP|20665-6|LNC|Echovirus 14 Ab|Echovirus 14 Ab
C0803469|T201|COMP|20666-4|LNC|Echovirus Ab|Echovirus Ab
C0803470|T201|COMP|20669-8|LNC|Cardiolipin Ab.IgA|Cardiolipin Ab.IgA
C0803471|T201|COMP|20671-4|LNC|Amino acids|Amino acids
C0803472|T201|COMP|20672-2|LNC|Actinobacillus pleuropneumoniae serotype|Actinobacillus pleuropneumoniae serotype
C0803473|T201|COMP|20673-0|LNC|Actinobacillus pleuropneumoniae Ab|Actinobacillus pleuropneumoniae Ab
C0803474|T201|COMP|20674-8|LNC|Avian adenovirus 2 Ag|Avian adenovirus 2 Ag
C0803475|T201|COMP|20675-5|LNC|Bovine adenovirus 3 Ag|Bovine adenovirus 3 Ag
C0803476|T201|COMP|20676-3|LNC|Bovine adenovirus 5 Ag|Bovine adenovirus 5 Ag
C0803477|T201|COMP|20677-1|LNC|Equine adenovirus Ag|Equine adenovirus Ag
C0803478|T201|COMP|20678-9|LNC|Alkaloid identified|Alkaloid identified
C0803479|T201|COMP|20679-7|LNC|Alkaloid identified|Alkaloid identified
C0803480|T201|COMP|20680-5|LNC|Alkaloid identified|Alkaloid identified
C0803481|T201|COMP|20681-3|LNC|Alpha tocopherol|Alpha tocopherol
C0803482|T201|COMP|20682-1|LNC|Ammonia|Ammonia
C0803483|T201|COMP|20683-9|LNC|Ammonia|Ammonia
C0803484|T201|COMP|20684-7|LNC|Ammonia|Ammonia
C0803485|T201|COMP|20685-4|LNC|Anaplasma marginale Ab|Anaplasma marginale Ab
C0803486|T201|COMP|20686-2|LNC|Anaplasma marginale Ab|Anaplasma marginale Ab
C0803487|T201|COMP|20687-0|LNC|Arsenic|Arsenic
C0803488|T201|COMP|20688-8|LNC|Aspergillus sp identified|Aspergillus sp identified
C0803489|T201|COMP|20689-6|LNC|Babesia caballi Ab|Babesia caballi Ab
C0803490|T201|COMP|20690-4|LNC|Theileria equi Ab|Theileria equi Ab
C0803491|T201|COMP|20691-2|LNC|Bacillus anthracis|Bacillus anthracis
C0803492|T201|COMP|20692-0|LNC|Bacillus cereus|Bacillus cereus
C0803493|T201|COMP|20693-8|LNC|Bacteria identified|Bacteria identified
C0803494|T201|COMP|20694-6|LNC|Bacteria identified|Bacteria identified
C0803495|T201|COMP|20695-3|LNC|Bacteria|Bacteria
C0803496|T201|COMP|20696-1|LNC|Bifidobacterium sp|Bifidobacterium sp
C0803497|T201|COMP|20697-9|LNC|Amines.biogenic|Amines.biogenic
C0803498|T201|COMP|20698-7|LNC|Bluetongue virus serotype|Bluetongue virus serotype
C0803499|T201|COMP|20699-5|LNC|Bluetongue virus Ab|Bluetongue virus Ab
C0803500|T201|COMP|20700-1|LNC|Bluetongue virus RNA|Bluetongue virus RNA
C0803501|T201|COMP|20701-9|LNC|Bluetongue virus Ag|Bluetongue virus Ag
C0803502|T201|COMP|20702-7|LNC|Bluetongue virus|Bluetongue virus
C0803503|T201|COMP|20703-5|LNC|Border disease virus Ag|Border disease virus Ag
C0803504|T201|COMP|20704-3|LNC|Border disease virus Ag|Border disease virus Ag
C0803505|T201|COMP|20705-0|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C0803506|T201|COMP|20706-8|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C0803507|T201|COMP|20707-6|LNC|Bovine leukosis virus Ab|Bovine leukosis virus Ab
C0803508|T201|COMP|20708-4|LNC|Bovine papular stomatitis virus Ag|Bovine papular stomatitis virus Ag
C0803509|T201|COMP|20709-2|LNC|Bovine diarrhea virus RNA|Bovine diarrhea virus RNA
C0803510|T201|COMP|20710-0|LNC|Bovine diarrhea virus RNA|Bovine diarrhea virus RNA
C0803511|T201|COMP|20711-8|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C0803512|T201|COMP|20712-6|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C0803513|T201|COMP|20713-4|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C0803514|T201|COMP|20714-2|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C0803515|T201|COMP|20715-9|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C0803516|T201|COMP|20716-7|LNC|Bovine diarrhea virus|Bovine diarrhea virus
C0803517|T201|COMP|20717-5|LNC|Bovine diarrhea virus 2 Ag|Bovine diarrhea virus 2 Ag
C0803518|T201|COMP|20718-3|LNC|Bromide|Bromide
C0803519|T201|COMP|20719-1|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803520|T201|COMP|20720-9|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803521|T201|COMP|20721-7|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803522|T201|COMP|20722-5|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803523|T201|COMP|20723-3|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803524|T201|COMP|20724-1|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803525|T201|COMP|20725-8|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803526|T201|COMP|20726-6|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803527|T201|COMP|20727-4|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803528|T201|COMP|20728-2|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803529|T201|COMP|20729-0|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803530|T201|COMP|20730-8|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803531|T201|COMP|20731-6|LNC|Brucella abortus Ab|Brucella abortus Ab
C0803532|T201|COMP|20732-4|LNC|Brucella ovis Ab|Brucella ovis Ab
C0803533|T201|COMP|20733-2|LNC|Brucella ovis Ab|Brucella ovis Ab
C0803534|T201|COMP|20734-0|LNC|Brucella sp identified|Brucella sp identified
C0803535|T201|COMP|20735-7|LNC|Brucella sp identified|Brucella sp identified
C0803536|T201|COMP|20736-5|LNC|Cache valley virus Ab|Cache valley virus Ab
C0803537|T201|COMP|20737-3|LNC|Cadmium|Cadmium
C0803538|T201|COMP|20738-1|LNC|Campylobacter sp identified|Campylobacter sp identified
C0803539|T201|COMP|20739-9|LNC|Campylobacter sp identified|Campylobacter sp identified
C0803540|T201|COMP|20740-7|LNC|Campylobacter sp identified|Campylobacter sp identified
C0803541|T201|COMP|20741-5|LNC|Canarypox virus Ag|Canarypox virus Ag
C0803542|T201|COMP|20742-3|LNC|Canine distemper virus Ag|Canine distemper virus Ag
C0803543|T201|COMP|15465-8|LNC|Caprine arthritis encephalitis virus Ab|Caprine arthritis encephalitis virus Ab
C0803544|T201|COMP|15464-1|LNC|Caprine arthritis encephalitis virus Ab|Caprine arthritis encephalitis virus Ab
C0803545|T201|COMP|20745-6|LNC|Carbamates|Carbamates
C0803546|T201|COMP|20746-4|LNC|Carbamates|Carbamates
C0803547|T201|COMP|20747-2|LNC|Carbamates|Carbamates
C0803548|T201|COMP|20748-0|LNC|Carbamates|Carbamates
C0803549|T201|COMP|20749-8|LNC|Carbamates|Carbamates
C0803550|T201|COMP|20750-6|LNC|Chicken anemia virus Ab|Chicken anemia virus Ab
C0803551|T201|COMP|20751-4|LNC|Chicken anemia virus Ab|Chicken anemia virus Ab
C0803552|T201|COMP|20752-2|LNC|Chlamydophila psittaci|Chlamydophila psittaci
C0803553|T201|COMP|20753-0|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C0803554|T201|COMP|20754-8|LNC|Chlamydophila psittaci Ab|Chlamydophila psittaci Ab
C0803555|T201|COMP|20755-5|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0803556|T201|COMP|20756-3|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0803557|T201|COMP|20757-1|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C0803558|T201|COMP|20758-9|LNC|Cholinesterase|Cholinesterase
C0803559|T201|COMP|20759-7|LNC|Chromium|Chromium
C0803560|T201|COMP|20760-5|LNC|Clostridium chauvoei Ag|Clostridium chauvoei Ag
C0803561|T201|COMP|20761-3|LNC|Clostridioides difficile|Clostridioides difficile
C0803562|T201|COMP|20762-1|LNC|Clostridioides difficile|Clostridioides difficile
C0803563|T201|COMP|20763-9|LNC|Clostridium novyii Ag|Clostridium novyii Ag
C0803564|T201|COMP|20764-7|LNC|Clostridium perfringens genotype|Clostridium perfringens genotype
C0803565|T201|COMP|20765-4|LNC|Clostridium septicum Ag|Clostridium septicum Ag
C0803566|T201|COMP|20766-2|LNC|Clostridium sordellii Ag|Clostridium sordellii Ag
C0803567|T201|COMP|20767-0|LNC|Coccidioides immitis|Coccidioides immitis
C0803568|T201|COMP|20768-8|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0803569|T201|COMP|20769-6|LNC|Coliform bacteria|Coliform bacteria
C0803570|T201|COMP|20770-4|LNC|Coliform bacteria|Coliform bacteria
C0803571|T201|COMP|20771-2|LNC|Coliform bacteria|Coliform bacteria
C0803572|T201|COMP|20772-0|LNC|Coliform colony count|Coliform colony count
C0803573|T201|COMP|20773-8|LNC|Colony count|Colony count
C0803574|T201|COMP|20774-6|LNC|Colony count|Colony count
C0803575|T201|COMP|20775-3|LNC|Colony count|Colony count
C0803576|T201|COMP|20776-1|LNC|Caprine parapoxvirus Ab|Caprine parapoxvirus Ab
C0803577|T201|COMP|20777-9|LNC|Caprine parapoxvirus Ab|Caprine parapoxvirus Ab
C0803578|T201|COMP|20778-7|LNC|Copper|Copper
C0803579|T201|COMP|20779-5|LNC|Bovine coronavirus Ag|Bovine coronavirus Ag
C0803580|T201|COMP|20780-3|LNC|Cryptosporidium sp|Cryptosporidium sp
C0803581|T201|COMP|20781-1|LNC|Cryptosporidium sp|Cryptosporidium sp
C0803582|T201|COMP|20782-9|LNC|Cyanide|Cyanide
C0803583|T201|COMP|20783-7|LNC|Cyanide|Cyanide
C0803584|T201|COMP|20784-5|LNC|Cyanide|Cyanide
C0803585|T201|COMP|20785-2|LNC|Drugs identified|Drugs identified
C0803586|T201|COMP|20786-0|LNC|Drugs identified|Drugs identified
C0803587|T201|COMP|20787-8|LNC|Drugs identified|Drugs identified
C0803588|T201|COMP|20788-6|LNC|Duck enteritis virus Ab|Duck enteritis virus Ab
C0803589|T201|COMP|20789-4|LNC|Escherichia coli serotype|Escherichia coli serotype
C0803590|T201|COMP|20790-2|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0803591|T201|COMP|20791-0|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0803592|T201|COMP|20792-8|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0803593|T201|COMP|20793-6|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0803594|T201|COMP|20794-4|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0803595|T201|COMP|20795-1|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0803596|T201|COMP|20796-9|LNC|Endophyte identified|Endophyte identified
C0803597|T201|COMP|20797-7|LNC|Endotoxin identified|Endotoxin identified
C0803598|T201|COMP|20798-5|LNC|Clostridium perfringens enterotoxin|Clostridium perfringens enterotoxin
C0803599|T201|COMP|20799-3|LNC|Clostridium perfringens enterotoxin|Clostridium perfringens enterotoxin
C0803600|T201|COMP|20800-9|LNC|Clostridium perfringens enterotoxin|Clostridium perfringens enterotoxin
C0803601|T201|COMP|20801-7|LNC|Encephalitozoon cuniculi Ab|Encephalitozoon cuniculi Ab
C0803602|T201|COMP|20802-5|LNC|Epizootic hemorrhagic disease virus Ab|Epizootic hemorrhagic disease virus Ab
C0803603|T201|COMP|20803-3|LNC|Epizootic hemorrhagic disease virus Ab|Epizootic hemorrhagic disease virus Ab
C0803604|T201|COMP|20804-1|LNC|Epizootic hemorrhagic disease virus Ag|Epizootic hemorrhagic disease virus Ag
C0803605|T201|COMP|20805-8|LNC|Epizootic hemorrhagic disease virus Ag|Epizootic hemorrhagic disease virus Ag
C0803606|T201|COMP|20806-6|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0803607|T201|COMP|20807-4|LNC|Equine arteritis virus|Equine arteritis virus
C0803608|T201|COMP|20808-2|LNC|Ergot alkaloid|Ergot alkaloid
C0803609|T201|COMP|20809-0|LNC|Ergot alkaloid|Ergot alkaloid
C0803611|T201|COMP|20811-6|LNC|Escherichia coli|Escherichia coli
C0803612|T201|COMP|20812-4|LNC|Escherichia coli 987P|Escherichia coli 987P
C0803613|T201|COMP|20813-2|LNC|Escherichia coli F41|Escherichia coli F41
C0803614|T201|COMP|20814-0|LNC|Escherichia coli F41|Escherichia coli F41
C0803615|T201|COMP|20815-7|LNC|Escherichia coli K88|Escherichia coli K88
C0803616|T201|COMP|20816-5|LNC|Escherichia coli K88|Escherichia coli K88
C0803617|T201|COMP|20817-3|LNC|Escherichia coli K88|Escherichia coli K88
C0803618|T201|COMP|20818-1|LNC|Escherichia coli K99|Escherichia coli K99
C0803619|T201|COMP|20819-9|LNC|Escherichia coli K99|Escherichia coli K99
C0803621|T201|COMP|20821-5|LNC|Escherichia coli K99|Escherichia coli K99
C0803622|T201|COMP|20822-3|LNC|Escherichia coli K99|Escherichia coli K99
C0803623|T201|COMP|20823-1|LNC|Escherichia coli O157:H7|Escherichia coli O157:H7
C0803624|T201|COMP|20824-9|LNC|Freezing point|Freezing point
C0803625|T201|COMP|20825-6|LNC|Fumonisin|Fumonisin
C0803626|T201|COMP|20826-4|LNC|Gallotannin|Gallotannin
C0803627|T201|COMP|20827-2|LNC|Gallotannin|Gallotannin
C0803628|T201|COMP|20828-0|LNC|Gallotannin|Gallotannin
C0803629|T201|COMP|20829-8|LNC|Glycol|Glycol
C0803630|T201|COMP|20830-6|LNC|Glycol|Glycol
C0803631|T201|COMP|20831-4|LNC|Glycolate|Glycolate
C0803632|T201|COMP|20832-2|LNC|Gossypol|Gossypol
C0803633|T201|COMP|20833-0|LNC|Haemophilus paragallinarum serotype|Haemophilus paragallinarum serotype
C0803634|T201|COMP|16941-7|LNC|Herbicide|Herbicide
C0803635|T201|COMP|20835-5|LNC|Herbicide|Herbicide
C0803636|T201|COMP|20836-3|LNC|Herbicide|Herbicide
C0803637|T201|COMP|20837-1|LNC|Herbicide|Herbicide
C0803638|T201|COMP|20838-9|LNC|Herbicide|Herbicide
C0803639|T201|COMP|20839-7|LNC|Herbicide|Herbicide
C0803640|T201|COMP|20840-5|LNC|Herbicide|Herbicide
C0803641|T201|COMP|20841-3|LNC|Herbicide|Herbicide
C0803642|T201|COMP|20842-1|LNC|Herbicide|Herbicide
C0803643|T201|COMP|20843-9|LNC|Avian infectious laryngotracheitis virus Ag|Avian infectious laryngotracheitis virus Ag
C0803644|T201|COMP|20844-7|LNC|Avian infectious laryngotracheitis virus Ag|Avian infectious laryngotracheitis virus Ag
C0803645|T201|COMP|20845-4|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C0803646|T201|COMP|20846-2|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C0803647|T201|COMP|20847-0|LNC|Bovine herpesvirus 2 Ag|Bovine herpesvirus 2 Ag
C0803648|T201|COMP|20848-8|LNC|Bovine herpesvirus 2 Ag|Bovine herpesvirus 2 Ag
C0803649|T201|COMP|20849-6|LNC|Bovine herpesvirus 4 Ag|Bovine herpesvirus 4 Ag
C0803650|T201|COMP|20850-4|LNC|Bovine herpesvirus 4 Ag|Bovine herpesvirus 4 Ag
C0803651|T201|COMP|20851-2|LNC|Bovine herpesvirus 5 Ag|Bovine herpesvirus 5 Ag
C0803652|T201|COMP|20852-0|LNC|Duck enteritis virus Ag|Duck enteritis virus Ag
C0803653|T201|COMP|20853-8|LNC|Equine herpesvirus 1 Ag|Equine herpesvirus 1 Ag
C0803654|T201|COMP|20854-6|LNC|Equine herpesvirus 1 Ag|Equine herpesvirus 1 Ag
C0803655|T201|COMP|20855-3|LNC|IgG.bovine|IgG.bovine
C0803656|T201|COMP|20856-1|LNC|IgG.equine|IgG.equine
C0803657|T201|COMP|20857-9|LNC|IgG.equine|IgG.equine
C0803658|T201|COMP|20858-7|LNC|Infectious bronchitis virus genotype|Infectious bronchitis virus genotype
C0803659|T201|COMP|20859-5|LNC|Infectious bronchitis virus serotype|Infectious bronchitis virus serotype
C0803660|T201|COMP|20860-3|LNC|Infectious bronchitis virus|Infectious bronchitis virus
C0803661|T201|COMP|20861-1|LNC|Infectious bronchitis virus genotype|Infectious bronchitis virus genotype
C0803662|T201|COMP|20862-9|LNC|Influenza virus A Ab|Influenza virus A Ab
C0803663|T201|COMP|20863-7|LNC|Iodine|Iodine
C0803664|T201|COMP|20864-5|LNC|Iodine|Iodine
C0803665|T201|COMP|20865-2|LNC|Iodine|Iodine
C0803666|T201|COMP|20866-0|LNC|Lactobacillus acidophilus colony count|Lactobacillus acidophilus colony count
C0803667|T201|COMP|20867-8|LNC|Lead|Lead
C0803668|T201|COMP|20868-6|LNC|Leptospira sp|Leptospira sp
C0803669|T201|COMP|20869-4|LNC|Leptospira sp|Leptospira sp
C0803670|T201|COMP|20870-2|LNC|Listeria sp|Listeria sp
C0803671|T201|COMP|20871-0|LNC|Listeria sp|Listeria sp
C0803672|T201|COMP|20872-8|LNC|Magnesium|Magnesium
C0803673|T201|COMP|20873-6|LNC|Alcelaphine herpesvirus 1 Ab|Alcelaphine herpesvirus 1 Ab
C0803674|T201|COMP|20874-4|LNC|Manganese|Manganese
C0803675|T201|COMP|20875-1|LNC|Manganese|Manganese
C0803676|T201|COMP|20876-9|LNC|Mercury|Mercury
C0803677|T201|COMP|20877-7|LNC|Bacteria identified|Bacteria identified
C0803678|T201|COMP|20878-5|LNC|Bacteria identified|Bacteria identified
C0803679|T201|COMP|20879-3|LNC|Bacteria identified|Bacteria identified
C0803685|T201|COMP|20886-8|LNC|Molybdenum|Molybdenum
C0803686|T201|COMP|20887-6|LNC|Molybdenum|Molybdenum
C0803687|T201|COMP|20888-4|LNC|Molybdenum|Molybdenum
C0803688|T201|COMP|20889-2|LNC|Monensin|Monensin
C0803689|T201|COMP|20890-0|LNC|Monensin|Monensin
C0803690|T201|COMP|20891-8|LNC|Mushroom identified|Mushroom identified
C0803691|T201|COMP|20892-6|LNC|Mycobacterium avium subspecies paratuberculosis|Mycobacterium avium subspecies paratuberculosis
C0803692|T201|COMP|20893-4|LNC|Mycobacterium avium subspecies paratuberculosis|Mycobacterium avium subspecies paratuberculosis
C0803694|T201|COMP|20895-9|LNC|Mycoplasma gallisepticum Ag|Mycoplasma gallisepticum Ag
C0803695|T201|COMP|20896-7|LNC|Mycoplasma sp|Mycoplasma sp
C0803696|T201|COMP|20897-5|LNC|Mycoplasma sp serotype|Mycoplasma sp serotype
C0803697|T201|COMP|20898-3|LNC|Mycoplasma sp|Mycoplasma sp
C0803698|T201|COMP|20899-1|LNC|Mycoplasma sp|Mycoplasma sp
C0803699|T201|COMP|20900-7|LNC|Mycoplasma sp Ab|Mycoplasma sp Ab
C0803700|T201|COMP|20901-5|LNC|Mycoplasma sp Ag|Mycoplasma sp Ag
C0803701|T201|COMP|20902-3|LNC|Mycoplasma sp+Ureaplasma sp|Mycoplasma sp+Ureaplasma sp
C0803702|T201|COMP|20903-1|LNC|Mycotoxin identified|Mycotoxin identified
C0803703|T201|COMP|20904-9|LNC|Neospora caninum Ab|Neospora caninum Ab
C0803704|T201|COMP|20905-6|LNC|Oleandrin|Oleandrin
C0803705|T201|COMP|20906-4|LNC|Oleandrin|Oleandrin
C0803706|T201|COMP|20907-2|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803707|T201|COMP|20908-0|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803708|T201|COMP|20909-8|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803709|T201|COMP|20910-6|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803710|T201|COMP|20911-4|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803711|T201|COMP|20912-2|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803712|T201|COMP|20913-0|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803713|T201|COMP|20914-8|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803714|T201|COMP|20915-5|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803715|T201|COMP|20916-3|LNC|Organochlorine pesticides|Organochlorine pesticides
C0803716|T201|COMP|20917-1|LNC|Organophosphate pesticides|Organophosphate pesticides
C0803717|T201|COMP|20918-9|LNC|Organophosphate pesticides|Organophosphate pesticides
C0803718|T201|COMP|20919-7|LNC|Organophosphate pesticides|Organophosphate pesticides
C0803719|T201|COMP|20920-5|LNC|Organophosphate pesticides|Organophosphate pesticides
C0803720|T201|COMP|20921-3|LNC|Organophosphate pesticides|Organophosphate pesticides
C0803721|T201|COMP|20922-1|LNC|Organophosphate pesticides|Organophosphate pesticides
C0803722|T201|COMP|20923-9|LNC|Organophosphate pesticides|Organophosphate pesticides
C0803723|T201|COMP|20924-7|LNC|Ova & parasites identified|Ova & parasites identified
C0803724|T201|COMP|20925-4|LNC|Ova & parasites identified|Ova & parasites identified
C0803725|T201|COMP|20926-2|LNC|Ova & parasites identified|Ova & parasites identified
C0803726|T201|COMP|20927-0|LNC|Oxalate|Oxalate
C0803727|T201|COMP|20928-8|LNC|Oxalate|Oxalate
C0803728|T201|COMP|20929-6|LNC|Paraquat|Paraquat
C0803729|T201|COMP|20930-4|LNC|Paraquat|Paraquat
C0803730|T201|COMP|20931-2|LNC|Parasites|Parasites
C0803731|T201|COMP|20932-0|LNC|Parasite identified|Parasite identified
C0803732|T201|COMP|20933-8|LNC|Parasite identified|Parasite identified
C0803733|T201|COMP|20934-6|LNC|Bovine parvovirus Ag|Bovine parvovirus Ag
C0803734|T201|COMP|20935-3|LNC|Pasteurella multocida serotype|Pasteurella multocida serotype
C0803735|T201|COMP|20936-1|LNC|Pentachlorophenol|Pentachlorophenol
C0803736|T201|COMP|20937-9|LNC|Pentachlorophenol|Pentachlorophenol
C0803737|T201|COMP|20938-7|LNC|Phenols|Phenols
C0803738|T201|COMP|20939-5|LNC|Phosphide|Phosphide
C0803739|T201|COMP|20940-3|LNC|Phosphide|Phosphide
C0803740|T201|COMP|20941-1|LNC|Phosphate|Phosphate
C0803742|T201|COMP|20943-7|LNC|Bovine respiratory syncytial virus Ag|Bovine respiratory syncytial virus Ag
C0803743|T201|COMP|20944-5|LNC|Bovine respiratory syncytial virus Ag|Bovine respiratory syncytial virus Ag
C0803744|T201|COMP|20945-2|LNC|Bovine respiratory syncytial virus Ag|Bovine respiratory syncytial virus Ag
C0803745|T201|COMP|20946-0|LNC|Retinol|Retinol
C0803746|T201|COMP|20947-8|LNC|Retinol|Retinol
C0803747|T201|COMP|20948-6|LNC|Retinol|Retinol
C0803748|T201|COMP|20949-4|LNC|Rickettsia sp|Rickettsia sp
C0803749|T201|COMP|20950-2|LNC|Bovine rotavirus Ag|Bovine rotavirus Ag
C0803750|T201|COMP|20951-0|LNC|Salmonella sp serotype|Salmonella sp serotype
C0803751|T201|COMP|20952-8|LNC|Salmonella sp identified|Salmonella sp identified
C0803752|T201|COMP|20953-6|LNC|Salmonella sp identified|Salmonella sp identified
C0803753|T201|COMP|17563-8|LNC|Salmonella sp identified|Salmonella sp identified
C0803754|T201|COMP|20955-1|LNC|Salmonella sp identified|Salmonella sp identified
C0803755|T201|COMP|20956-9|LNC|Sarcocystis neurona Ab|Sarcocystis neurona Ab
C0803756|T201|COMP|20957-7|LNC|Sarcocystis neurona Ab|Sarcocystis neurona Ab
C0803757|T201|COMP|20958-5|LNC|Sarcocystis neurona Ab|Sarcocystis neurona Ab
C0803758|T201|COMP|20959-3|LNC|Sarcocystis neurona Ag|Sarcocystis neurona Ag
C0803759|T201|COMP|20960-1|LNC|Selenium|Selenium
C0803760|T201|COMP|20961-9|LNC|Selenium|Selenium
C0803761|T201|COMP|20962-7|LNC|Serpulina hyodysenteria|Serpulina hyodysenteria
C0803762|T201|COMP|20963-5|LNC|Serpulina hyodysenteria|Serpulina hyodysenteria
C0803763|T201|COMP|20964-3|LNC|Shigella sp identified|Shigella sp identified
C0803764|T201|COMP|20965-0|LNC|Somatic cells|Somatic cells
C0803765|T201|COMP|20966-8|LNC|Staphylococcus sp identified|Staphylococcus sp identified
C0803766|T201|COMP|20967-6|LNC|Staphylococcus sp identified|Staphylococcus sp identified
C0803767|T201|COMP|20968-4|LNC|Staphylococcus sp identified|Staphylococcus sp identified
C0803768|T201|COMP|20969-2|LNC|Strychnine|Strychnine
C0803769|T201|COMP|20970-0|LNC|Strychnine|Strychnine
C0803770|T201|COMP|20972-6|LNC|Strychnine|Strychnine
C0803771|T201|COMP|20973-4|LNC|Sulfate|Sulfate
C0803772|T201|COMP|20974-2|LNC|Sulfate|Sulfate
C0803773|T201|COMP|20975-9|LNC|Thallium|Thallium
C0803774|T201|COMP|20976-7|LNC|Tritrichomonas foetus|Tritrichomonas foetus
C0803775|T201|COMP|20977-5|LNC|Urea|Urea
C0803776|T201|COMP|20978-3|LNC|Urea|Urea
C0803777|T201|COMP|20979-1|LNC|Urea|Urea
C0803778|T201|COMP|20980-9|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C0803779|T201|COMP|20981-7|LNC|Verotoxin identified|Verotoxin identified
C0803780|T201|COMP|20982-5|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0803781|T201|COMP|20983-3|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0803782|T201|COMP|20984-1|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0803783|T201|COMP|20985-8|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0803784|T201|COMP|20986-6|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0803785|T201|COMP|20987-4|LNC|Yersinia sp identified|Yersinia sp identified
C0803786|T201|COMP|20988-2|LNC|Zinc phosphide|Zinc phosphide
C0803787|T201|COMP|20989-0|LNC|Zinc phosphide|Zinc phosphide
C0803788|T201|COMP|20990-8|LNC|APC gene targeted mutation analysis|APC gene targeted mutation analysis
C0803789|T201|COMP|20991-6|LNC|Antithrombin|Antithrombin
C0803790|T201|COMP|20992-4|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C0803791|T201|COMP|6358-6|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C0803792|T201|COMP|20994-0|LNC|Choriogonadotropin|Choriogonadotropin
C0803793|T201|COMP|20995-7|LNC|Cortisol^1H post dose corticotropin|Cortisol^1H post dose corticotropin
C0803794|T201|COMP|20996-5|LNC|Coxsackievirus B1+B2+B3+B4+B5+B6 Ab|Coxsackievirus B1+B2+B3+B4+B5+B6 Ab
C0803795|T201|COMP|20998-1|LNC|Cell fractions|Cell fractions
C0803796|T201|COMP|20999-9|LNC|Cell fractions|Cell fractions
C0803797|T201|COMP|21000-5|LNC|Erythrocyte distribution width|Erythrocyte distribution width
C0803798|T201|COMP|21001-3|LNC|Coagulation factor VIII|Coagulation factor VIII
C0803799|T201|COMP|21002-1|LNC|Fibrinogen|Fibrinogen
C0803800|T201|COMP|21003-9|LNC|Fungus identified|Fungus identified
C0803801|T201|COMP|21004-7|LNC|Glucose tolerance|Glucose tolerance
C0803802|T201|COMP|21005-4|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C0803803|T201|COMP|21006-2|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0803804|T201|COMP|21007-0|LNC|HIV 1 Ab|HIV 1 Ab
C0803805|T201|COMP|21008-8|LNC|HIV 1 RNA|HIV 1 RNA
C0803806|T201|COMP|21009-6|LNC|HIV 1|HIV 1
C0803807|T201|COMP|21010-4|LNC|Cells.CD1|Cells.CD1
C0803808|T201|COMP|21011-2|LNC|Cells.CD13|Cells.CD13
C0803809|T201|COMP|21012-0|LNC|Cells.CD15|Cells.CD15
C0803810|T201|COMP|21013-8|LNC|Cells.CD22|Cells.CD22
C0803811|T201|COMP|21014-6|LNC|Cells.CD24|Cells.CD24
C0803812|T201|COMP|21015-3|LNC|Cells.CD33|Cells.CD33
C0803813|T201|COMP|21016-1|LNC|Cells.CD41|Cells.CD41
C0803814|T201|COMP|21017-9|LNC|Cells.CD57|Cells.CD57
C0803815|T201|COMP|21018-7|LNC|Cells.CD61|Cells.CD61
C0803816|T201|COMP|19050-4|LNC|Metanephrines|Metanephrines
C0803817|T201|COMP|21020-3|LNC|Bacteria identified|Bacteria identified
C0803820|T201|COMP|21023-7|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C0803821|T201|COMP|21024-5|LNC|Pathologist interpretation|Pathologist interpretation
C0803822|T201|COMP|21025-2|LNC|Pathologist interpretation|Pathologist interpretation
C0803823|T201|COMP|21026-0|LNC|Pathologist interpretation|Pathologist interpretation
C0803824|T201|COMP|21027-8|LNC|Platelet aggregation|Platelet aggregation
C0803825|T201|COMP|21028-6|LNC|Protein|Protein
C0803826|T201|COMP|21030-2|LNC|Reagin Ab|Reagin Ab
C0803827|T201|COMP|21031-0|LNC|Saint Louis encephalitis virus|Saint Louis encephalitis virus
C0803828|T201|COMP|21032-8|LNC|Coagulation thrombin induced|Coagulation thrombin induced
C0803829|T201|COMP|21033-6|LNC|Yeast.budding|Yeast.budding
C0803830|T201|COMP|21034-4|LNC|11-Deoxycortisol^evening specimen|11-Deoxycortisol^evening specimen
C0803831|T201|COMP|21035-1|LNC|11-Deoxycortisol^morning specimen|11-Deoxycortisol^morning specimen
C0803832|T201|COMP|21036-9|LNC|17-Hydroxycorticosteroids|17-Hydroxycorticosteroids
C0803833|T201|COMP|21037-7|LNC|17-Hydroxypregnenolone|17-Hydroxypregnenolone
C0803834|T201|COMP|21038-5|LNC|17-Ketosteroids|17-Ketosteroids
C0803835|T201|COMP|21039-3|LNC|18-Hydroxycortisol|18-Hydroxycortisol
C0803837|T201|COMP|21041-9|LNC|3-Hydroxydodecanedioate/Creatinine|3-Hydroxydodecanedioate/Creatinine
C0803838|T201|COMP|21042-7|LNC|3-Hydroxydodecanoate/Creatinine|3-Hydroxydodecanoate/Creatinine
C0803839|T201|COMP|21043-5|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C0803840|T201|COMP|21044-3|LNC|5-Alpha tetrahydrocortisol|5-Alpha tetrahydrocortisol
C0803841|T201|COMP|21045-0|LNC|5-Hydroxytryptophan|5-Hydroxytryptophan
C0803842|T201|COMP|21046-8|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C0803843|T201|COMP|21047-6|LNC|8-Hydroxyloxapine|8-Hydroxyloxapine
C0803844|T201|COMP|21048-4|LNC|Acetaldehyde|Acetaldehyde
C0803845|T201|COMP|21049-2|LNC|Acetone|Acetone
C0803847|T201|COMP|21051-8|LNC|Acrylaldehyde|Acrylaldehyde
C0803848|T201|COMP|21052-6|LNC|Adenosine monophosphate.cyclic.nephrogenous|Adenosine monophosphate.cyclic.nephrogenous
C0803849|T201|COMP|21053-4|LNC|Adenovirus Ab.IgG|Adenovirus Ab.IgG
C0803850|T201|COMP|21054-2|LNC|Adenovirus Ab.IgM|Adenovirus Ab.IgM
C0803851|T201|COMP|21055-9|LNC|Adenovirus DNA|Adenovirus DNA
C0803853|T201|COMP|21057-5|LNC|Alanine+Histidine+Leucine+Phenylalanine+Tyrosine|Alanine+Histidine+Leucine+Phenylalanine+Tyrosine
C0803854|T201|COMP|21058-3|LNC|Albumin^2H post peritoneal dialysis|Albumin^2H post peritoneal dialysis
C0803855|T201|COMP|21059-1|LNC|Albumin|Albumin
C0803856|T201|COMP|21060-9|LNC|Alnus incana Ab.IgE.RAST class|Alnus incana Ab.IgE.RAST class
C0803857|T201|COMP|21061-7|LNC|Medicago sativa Ab.IgG.RAST class|Medicago sativa Ab.IgG.RAST class
C0803858|T201|COMP|21062-5|LNC|Allobarbital|Allobarbital
C0803859|T201|COMP|21063-3|LNC|Prunus dulcis Ab.IgG.RAST class|Prunus dulcis Ab.IgG.RAST class
C0803860|T201|COMP|21064-1|LNC|Acid alpha glucosidase|Acid alpha glucosidase
C0803861|T201|COMP|21065-8|LNC|Alternaria alternata Ab.IgG.RAST class|Alternaria alternata Ab.IgG.RAST class
C0803862|T201|COMP|21066-6|LNC|Ampicillin|Ampicillin
C0803863|T201|COMP|21067-4|LNC|Monomorium minimum Ab.IgE.RAST class|Monomorium minimum Ab.IgE.RAST class
C0803864|T201|COMP|21068-2|LNC|Pogonomyrmex barbatus Ab.IgE.RAST class|Pogonomyrmex barbatus Ab.IgE.RAST class
C0803865|T201|COMP|21070-8|LNC|Antibiotic XXX|Antibiotic XXX
C0803866|T201|COMP|21071-6|LNC|Antimony|Antimony
C0803867|T201|COMP|21072-4|LNC|Malus sylvestris Ab.IgG.RAST class|Malus sylvestris Ab.IgG.RAST class
C0803868|T201|COMP|21073-2|LNC|Prunus armeniaca Ab.IgG.RAST class|Prunus armeniaca Ab.IgG.RAST class
C0803869|T201|COMP|21074-0|LNC|Arsenic|Arsenic
C0803870|T201|COMP|21075-7|LNC|Ascaris lumbricoides Ab.IgE|Ascaris lumbricoides Ab.IgE
C0803871|T201|COMP|21076-5|LNC|Ascaris lumbricoides Ab.IgE.RAST class|Ascaris lumbricoides Ab.IgE.RAST class
C0803872|T201|COMP|21077-3|LNC|Fraxinus nigra Ab.IgE|Fraxinus nigra Ab.IgE
C0803873|T201|COMP|21078-1|LNC|Fraxinus pennsylvanica Ab.IgE|Fraxinus pennsylvanica Ab.IgE
C0803874|T201|COMP|21079-9|LNC|Fraxinus pennsylvanica Ab.IgE.RAST class|Fraxinus pennsylvanica Ab.IgE.RAST class
C0803875|T201|COMP|21080-7|LNC|Asialoganglioside GM1 Ab|Asialoganglioside GM1 Ab
C0803876|T201|COMP|21081-5|LNC|ASPA gene targeted mutation analysis|ASPA gene targeted mutation analysis
C0803877|T201|COMP|21082-3|LNC|Asparagus officinalis Ab.IgG.RAST class|Asparagus officinalis Ab.IgG.RAST class
C0803878|T201|COMP|15548-1|LNC|Populus tremula Ab.IgE.RAST class|Populus tremula Ab.IgE.RAST class
C0803879|T201|COMP|21084-9|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C0803880|T201|COMP|21085-6|LNC|Aspergillus fumigatus Ab|Aspergillus fumigatus Ab
C0803881|T201|COMP|21086-4|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C0803882|T201|COMP|21087-2|LNC|Aspergillus terreus Ab.IgE.RAST class|Aspergillus terreus Ab.IgE.RAST class
C0803883|T201|COMP|21088-0|LNC|Azinphos-methyl|Azinphos-methyl
C0803884|T201|COMP|21089-8|LNC|Babesia microti DNA|Babesia microti DNA
C0803885|T201|COMP|21090-6|LNC|Musa spp Ab.IgG.RAST class|Musa spp Ab.IgG.RAST class
C0803886|T201|COMP|21091-4|LNC|Barbiturates present|Barbiturates present
C0803887|T201|COMP|21092-2|LNC|Hordeum vulgare Ab.IgG.RAST class|Hordeum vulgare Ab.IgG.RAST class
C0803888|T201|COMP|21093-0|LNC|Basement membrane Ab.IgG|Basement membrane Ab.IgG
C0803889|T201|COMP|21094-8|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0803891|T201|COMP|21096-3|LNC|Bean black Ab.IgE|Bean black Ab.IgE
C0803892|T201|COMP|21097-1|LNC|Bean black Ab.IgE.RAST class|Bean black Ab.IgE.RAST class
C0803893|T201|COMP|21098-9|LNC|Bean green Ab.IgG.RAST class|Bean green Ab.IgG.RAST class
C0803894|T201|COMP|21099-7|LNC|Bean kidney red Ab.IgG.RAST class|Bean kidney red Ab.IgG.RAST class
C0803895|T201|COMP|21100-3|LNC|Vigna radiata Ab.IgG.RAST class|Vigna radiata Ab.IgG.RAST class
C0803896|T201|COMP|21101-1|LNC|Bean pinto Ab.IgG.RAST class|Bean pinto Ab.IgG.RAST class
C0803897|T201|COMP|21102-9|LNC|Glycine max Ab.IgG.RAST class|Glycine max Ab.IgG.RAST class
C0803898|T201|COMP|21104-5|LNC|Glycine max dust Ab.IgE.RAST class|Glycine max dust Ab.IgE.RAST class
C0803899|T201|COMP|21105-2|LNC|Bean yellow Ab.IgG.RAST class|Bean yellow Ab.IgG.RAST class
C0803900|T201|COMP|21106-0|LNC|Beef Ab.IgG.RAST class|Beef Ab.IgG.RAST class
C0803901|T201|COMP|21107-8|LNC|Bendiocarb|Bendiocarb
C0803902|T201|COMP|21108-6|LNC|Beta 2 glycoprotein 1 Ab.IgA|Beta 2 glycoprotein 1 Ab.IgA
C0803903|T201|COMP|21109-4|LNC|Beta lactoglobulin Ab.IgG.RAST class|Beta lactoglobulin Ab.IgG.RAST class
C0803906|T201|COMP|21112-8|LNC|Birth date|Birth date
C0803907|T201|COMP|21113-6|LNC|Bismuth|Bismuth
C0803908|T201|COMP|21114-4|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C0803909|T201|COMP|21115-1|LNC|Vaccinium myrtillus Ab.IgG.RAST class|Vaccinium myrtillus Ab.IgG.RAST class
C0803910|T201|COMP|21116-9|LNC|Borrelia burgdorferi 66kD Ab.IgM|Borrelia burgdorferi 66kD Ab.IgM
C0803911|T201|COMP|21117-7|LNC|Borrelia burgdorferi 93kD Ab.IgM|Borrelia burgdorferi 93kD Ab.IgM
C0803912|T201|COMP|21118-5|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0803913|T201|COMP|21119-3|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0803914|T201|COMP|21120-1|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C0803915|T201|COMP|21121-9|LNC|Borrelia hermsii Ab.IgG|Borrelia hermsii Ab.IgG
C0803916|T201|COMP|21122-7|LNC|Borrelia hermsii Ab.IgM|Borrelia hermsii Ab.IgM
C0803917|T201|COMP|21123-5|LNC|Bran wheat Ab.IgE.RAST class|Bran wheat Ab.IgE.RAST class
C0803918|T201|COMP|21124-3|LNC|Brassica oleracea var italica Ab.IgG.RAST class|Brassica oleracea var italica Ab.IgG.RAST class
C0803919|T201|COMP|21125-0|LNC|Brush border Ab|Brush border Ab
C0803920|T201|COMP|21126-8|LNC|Brassica oleracea var gemmifera Ab.IgG.RAST class|Brassica oleracea var gemmifera Ab.IgG.RAST class
C0803921|T201|COMP|21127-6|LNC|Brassica oleracea var capitata Ab.IgG.RAST class|Brassica oleracea var capitata Ab.IgG.RAST class
C0803922|T201|COMP|21128-4|LNC|Cadmium|Cadmium
C0803923|T201|COMP|21129-2|LNC|Cadmium|Cadmium
C0803924|T201|COMP|21130-0|LNC|Cadmium|Cadmium
C0803925|T201|COMP|21131-8|LNC|Calcitonin^10M post 0.5 ug/kg pentagastrin IV|Calcitonin^10M post 0.5 ug/kg pentagastrin IV
C0803926|T201|COMP|21132-6|LNC|Calcitonin^1M post 0.5 ug/kg pentagastrin IV|Calcitonin^1M post 0.5 ug/kg pentagastrin IV
C0803927|T201|COMP|21133-4|LNC|Calcitonin^2M post 0.5 ug/kg pentagastrin IV|Calcitonin^2M post 0.5 ug/kg pentagastrin IV
C0803928|T201|COMP|21134-2|LNC|Calcitonin^3M post 0.5 ug/kg pentagastrin IV|Calcitonin^3M post 0.5 ug/kg pentagastrin IV
C0803929|T201|COMP|21135-9|LNC|Canrenone|Canrenone
C0803930|T201|COMP|21136-7|LNC|Cucumis melo spp Ab.IgG.RAST class|Cucumis melo spp Ab.IgG.RAST class
C0803931|T201|COMP|21137-5|LNC|Carageenan Ab.IgE.RAST class|Carageenan Ab.IgE.RAST class
C0803932|T201|COMP|21138-3|LNC|Carbaryl|Carbaryl
C0803933|T201|COMP|21139-1|LNC|Carbofuran|Carbofuran
C0803934|T201|COMP|21140-9|LNC|Carbophenothion|Carbophenothion
C0803935|T201|COMP|21141-7|LNC|Elettaria cardamomum Ab.IgE.RAST class|Elettaria cardamomum Ab.IgE.RAST class
C0803936|T201|COMP|21142-5|LNC|Carisoprodol|Carisoprodol
C0803937|T201|COMP|21143-3|LNC|Carp Ab.IgE|Carp Ab.IgE
C0803938|T201|COMP|21144-1|LNC|Carp Ab.IgE.RAST class|Carp Ab.IgE.RAST class
C0803939|T201|COMP|21145-8|LNC|Daucus carota Ab.IgG.RAST class|Daucus carota Ab.IgG.RAST class
C0803940|T201|COMP|21146-6|LNC|Casein Ab.IgG.RAST class|Casein Ab.IgG.RAST class
C0803941|T201|COMP|21147-4|LNC|Brassica oleracea var botrytis Ab.IgG.RAST class|Brassica oleracea var botrytis Ab.IgG.RAST class
C0803942|T201|COMP|21148-2|LNC|Cedar white Ab.IgE|Cedar white Ab.IgE
C0803943|T201|COMP|19733-5|LNC|Cefaclor Ab.IgE|Cefaclor Ab.IgE
C0803944|T201|COMP|21150-8|LNC|Cefaclor Ab.IgE.RAST class|Cefaclor Ab.IgE.RAST class
C0803945|T201|COMP|21151-6|LNC|cefTAZidime|cefTAZidime
C0803946|T201|COMP|21152-4|LNC|Apium graveolens Ab.IgG.RAST class|Apium graveolens Ab.IgG.RAST class
C0803947|T201|COMP|21153-2|LNC|Cells.CD10/Gated cells.total|Cells.CD10/Gated cells.total
C0803948|T201|COMP|21154-0|LNC|Cells.CD11c/100 cells|Cells.CD11c/100 cells
C0803949|T201|COMP|21155-7|LNC|Cells.CD13/Gated cells.total|Cells.CD13/Gated cells.total
C0803950|T201|COMP|21156-5|LNC|Cells.CD14/Gated cells.total|Cells.CD14/Gated cells.total
C0803951|T201|COMP|21157-3|LNC|Cells.CD19/Gated cells.total|Cells.CD19/Gated cells.total
C0803952|T201|COMP|21158-1|LNC|Cells.CD20/Gated cells.total|Cells.CD20/Gated cells.total
C0803953|T201|COMP|21159-9|LNC|Cells.CD23/Gated cells.total|Cells.CD23/Gated cells.total
C0803954|T201|COMP|21160-7|LNC|Cells.CD3/Gated cells.total|Cells.CD3/Gated cells.total
C0803955|T201|COMP|21161-5|LNC|Cells.CD33/Gated cells.total|Cells.CD33/Gated cells.total
C0803956|T201|COMP|21162-3|LNC|Cells.CD34/Gated cells.total|Cells.CD34/Gated cells.total
C0803957|T201|COMP|21163-1|LNC|Cells.CD38/Gated cells.total|Cells.CD38/Gated cells.total
C0803958|T201|COMP|21164-9|LNC|Cells.CD4/Gated cells.total|Cells.CD4/Gated cells.total
C0803959|T201|COMP|21165-6|LNC|Cells.CD5/Gated cells.total|Cells.CD5/Gated cells.total
C0803961|T201|COMP|21167-2|LNC|Cells.CD61/100 cells|Cells.CD61/100 cells
C0803962|T201|COMP|21168-0|LNC|Cells.CD7/Gated cells.total|Cells.CD7/Gated cells.total
C0803963|T201|COMP|21169-8|LNC|Cells.CD71/100 cells|Cells.CD71/100 cells
C0803964|T201|COMP|21170-6|LNC|Cells.CD8/Gated cells.total|Cells.CD8/Gated cells.total
C0803965|T201|COMP|21171-4|LNC|Cells.FMC7/100 cells|Cells.FMC7/100 cells
C0803966|T201|COMP|21172-2|LNC|Cells.XXX/100 cells|Cells.XXX/100 cells
C0803967|T201|COMP|21173-0|LNC|Cephaeline|Cephaeline
C0803968|T201|COMP|21174-8|LNC|Cephaeline|Cephaeline
C0803969|T201|COMP|21175-5|LNC|Cephalexin|Cephalexin
C0803970|T201|COMP|21176-3|LNC|Cerebroventricular lining cells|Cerebroventricular lining cells
C0803971|T201|COMP|21654-9|LNC|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C0803972|T201|COMP|21178-9|LNC|Cheese cheddar type Ab.IgG.RAST class|Cheese cheddar type Ab.IgG.RAST class
C0803973|T201|COMP|21179-7|LNC|Cheese cream Ab.IgE.RAST class|Cheese cream Ab.IgE.RAST class
C0803974|T201|COMP|21180-5|LNC|Cheese roquefort Ab.IgE.RAST class|Cheese roquefort Ab.IgE.RAST class
C0803975|T201|COMP|21181-3|LNC|Prunus avium Ab.IgG.RAST class|Prunus avium Ab.IgG.RAST class
C0803976|T201|COMP|21182-1|LNC|Chicken Ab.IgG.RAST class|Chicken Ab.IgG.RAST class
C0803977|T201|COMP|21183-9|LNC|Chicken meat Ab.IgG.RAST class|Chicken meat Ab.IgG.RAST class
C0803978|T201|COMP|21184-7|LNC|Chlamydophila pneumoniae|Chlamydophila pneumoniae
C0803979|T201|COMP|21185-4|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C0803980|T201|COMP|21186-2|LNC|Chlamydia sp Ab.IgM|Chlamydia sp Ab.IgM
C0803981|T201|COMP|21187-0|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0803982|T201|COMP|21188-8|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C0803983|T201|COMP|21189-6|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0803984|T201|COMP|21190-4|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0803985|T201|COMP|21191-2|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0803986|T201|COMP|21192-0|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C0803987|T201|COMP|21193-8|LNC|Chlordiazepoxide+Norchlordiazepoxide|Chlordiazepoxide+Norchlordiazepoxide
C0803988|T201|COMP|21194-6|LNC|Chloride|Chloride
C0803989|T201|COMP|21195-3|LNC|Chlorzoxazone|Chlorzoxazone
C0803990|T201|COMP|21196-1|LNC|Chocolate Ab.IgG.RAST class|Chocolate Ab.IgG.RAST class
C0803991|T201|COMP|21197-9|LNC|Cholesterol esters/Cholesterol.total|Cholesterol esters/Cholesterol.total
C0803992|T201|COMP|21198-7|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0803993|T201|COMP|21199-5|LNC|Chromium|Chromium
C0803994|T201|COMP|21200-1|LNC|Chromium|Chromium
C0803995|T201|COMP|21201-9|LNC|Chromium|Chromium
C0803996|T201|COMP|21202-7|LNC|Cinnamomum spp Ab.IgG.RAST class|Cinnamomum spp Ab.IgG.RAST class
C0803997|T201|COMP|21203-5|LNC|Citrate|Citrate
C0803998|T201|COMP|21204-3|LNC|Ruditapes spp Ab.IgG.RAST class|Ruditapes spp Ab.IgG.RAST class
C0803999|T201|COMP|21205-0|LNC|Syzygium aromaticum Ab.IgG.RAST class|Syzygium aromaticum Ab.IgG.RAST class
C0804000|T201|COMP|21206-8|LNC|Clover sweet Ab.IgE|Clover sweet Ab.IgE
C0804001|T201|COMP|21207-6|LNC|CCR5 gene targeted mutation analysis|CCR5 gene targeted mutation analysis
C0804002|T201|COMP|21208-4|LNC|Cobalt|Cobalt
C0804003|T201|COMP|21209-2|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0804004|T201|COMP|21210-0|LNC|Cockatiel droppings Ab.IgE.RAST class|Cockatiel droppings Ab.IgE.RAST class
C0804005|T201|COMP|21211-8|LNC|Cockatiel feather Ab.IgE.RAST class|Cockatiel feather Ab.IgE.RAST class
C0804006|T201|COMP|21212-6|LNC|Cocos nucifera Ab.IgG.RAST class|Cocos nucifera Ab.IgG.RAST class
C0804007|T201|COMP|21213-4|LNC|Gadus morhua Ab.IgG.RAST class|Gadus morhua Ab.IgG.RAST class
C0804008|T201|COMP|21214-2|LNC|Coffea spp Ab.IgG.RAST class|Coffea spp Ab.IgG.RAST class
C0804009|T201|COMP|21215-9|LNC|Collagen crosslinked N-telopeptide|Collagen crosslinked N-telopeptide
C0804010|T201|COMP|21216-7|LNC|Collagen crosslinked N-telopeptide/Creatinine|Collagen crosslinked N-telopeptide/Creatinine
C0804011|T201|COMP|21217-5|LNC|Complement C4d|Complement C4d
C0804012|T201|COMP|21218-3|LNC|Complement total hemolytic CH50|Complement total hemolytic CH50
C0804013|T201|COMP|21219-1|LNC|Copper|Copper
C0804014|T201|COMP|21220-9|LNC|Coriandrum sativum Ab.IgE.RAST class|Coriandrum sativum Ab.IgE.RAST class
C0804015|T201|COMP|21221-7|LNC|Zea mays Ab.IgG.RAST class|Zea mays Ab.IgG.RAST class
C0804016|T201|COMP|21222-5|LNC|Cortisol^11 PM specimen|Cortisol^11 PM specimen
C0804017|T201|COMP|21223-3|LNC|Cortisol^1st specimen post XXX challenge|Cortisol^1st specimen post XXX challenge
C0804018|T201|COMP|21224-1|LNC|Cortisol^2H post XXX challenge|Cortisol^2H post XXX challenge
C0804019|T201|COMP|21225-8|LNC|Cortisol^3H post XXX challenge|Cortisol^3H post XXX challenge
C0804020|T201|COMP|21226-6|LNC|Cortisol^4 PM specimen|Cortisol^4 PM specimen
C0804021|T201|COMP|21227-4|LNC|Cotton linters Ab.IgE.RAST class|Cotton linters Ab.IgE.RAST class
C0804022|T201|COMP|21228-2|LNC|Cottonseed Ab.IgG.RAST class|Cottonseed Ab.IgG.RAST class
C0804023|T201|COMP|21229-0|LNC|Coumaphos|Coumaphos
C0804024|T201|COMP|21230-8|LNC|Cow milk Ab.IgG.RAST class|Cow milk Ab.IgG.RAST class
C0804025|T201|COMP|21231-6|LNC|Cancer pagurus Ab.IgG.RAST class|Cancer pagurus Ab.IgG.RAST class
C0804026|T201|COMP|21232-4|LNC|Creatinine|Creatinine
C0804027|T201|COMP|21233-2|LNC|Cryptosporidium sp Ag|Cryptosporidium sp Ag
C0804028|T201|COMP|21234-0|LNC|Cucumis sativus Ab.IgG.RAST class|Cucumis sativus Ab.IgG.RAST class
C0804029|T201|COMP|21235-7|LNC|Cuminum cyminum Ab.IgE.RAST class|Cuminum cyminum Ab.IgE.RAST class
C0804030|T201|COMP|21236-5|LNC|Cyclohexanone|Cyclohexanone
C0804031|T201|COMP|21237-3|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0804032|T201|COMP|21238-1|LNC|Deer hair Ab.IgE.RAST class|Deer hair Ab.IgE.RAST class
C0804033|T201|COMP|21239-9|LNC|Desalkylhalazepam|Desalkylhalazepam
C0804034|T201|COMP|21240-7|LNC|Dextromethorphan|Dextromethorphan
C0804035|T201|COMP|21241-5|LNC|Diazepam+Nordiazepam|Diazepam+Nordiazepam
C0804036|T201|COMP|21242-3|LNC|Protoporphyrin|Protoporphyrin
C0804037|T201|COMP|21243-1|LNC|Diethyl ether|Diethyl ether
C0804038|T201|COMP|16366-7|LNC|Diethylpropion|Diethylpropion
C0804039|T201|COMP|21245-6|LNC|Diisobutylketone|Diisobutylketone
C0804040|T201|COMP|21246-4|LNC|Dimethoate|Dimethoate
C0804041|T201|COMP|21247-2|LNC|DMD gene targeted mutation analysis|DMD gene targeted mutation analysis
C0804042|T201|COMP|21248-0|LNC|DOBUTamine|DOBUTamine
C0804043|T201|COMP|21249-8|LNC|Dolichol|Dolichol
C0804044|T201|COMP|21250-6|LNC|Doxycycline|Doxycycline
C0804045|T201|COMP|21251-4|LNC|Echinococcus granulosus Ab.IgE.RAST class|Echinococcus granulosus Ab.IgE.RAST class
C0804046|T201|COMP|21252-2|LNC|Echinococcus granulosus Ab.IgG|Echinococcus granulosus Ab.IgG
C0804047|T201|COMP|21253-0|LNC|Egg white Ab.IgG.RAST class|Egg white Ab.IgG.RAST class
C0804048|T201|COMP|21254-8|LNC|Egg yolk Ab.IgG.RAST class|Egg yolk Ab.IgG.RAST class
C0804049|T201|COMP|21255-5|LNC|Solanum melongena Ab.IgG.RAST class|Solanum melongena Ab.IgG.RAST class
C0804052|T201|COMP|21258-9|LNC|Cichorium endivia Ab.IgG.RAST class|Cichorium endivia Ab.IgG.RAST class
C0804053|T201|COMP|21259-7|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0804054|T201|COMP|21260-5|LNC|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C0804055|T201|COMP|21261-3|LNC|Erythromycin Ab.IgE.RAST class|Erythromycin Ab.IgE.RAST class
C0804056|T201|COMP|21262-1|LNC|Escherichia coli shiga-like toxin|Escherichia coli shiga-like toxin
C0804057|T201|COMP|21263-9|LNC|Estradiol|Estradiol
C0804058|T201|COMP|21264-7|LNC|Estriol.unconjugated^^adjusted|Estriol.unconjugated^^adjusted
C0804059|T201|COMP|21265-4|LNC|Estriol.unconjugated^^unadjusted|Estriol.unconjugated^^unadjusted
C0804060|T201|COMP|21266-2|LNC|Ethion|Ethion
C0804061|T201|COMP|21267-0|LNC|O-Ethyl O-(p-nitrophenyl) phenylphosphonothionate|O-Ethyl O-(p-nitrophenyl) phenylphosphonothionate
C0804062|T201|COMP|21268-8|LNC|Fenchlorphos|Fenchlorphos
C0804063|T201|COMP|21269-6|LNC|Fenthion|Fenthion
C0804064|T201|COMP|21270-4|LNC|Ficus carica Ab.IgE.RAST class|Ficus carica Ab.IgE.RAST class
C0804065|T201|COMP|21271-2|LNC|Chamerion angustifolium Ab.IgE|Chamerion angustifolium Ab.IgE
C0804066|T201|COMP|21272-0|LNC|Chamerion angustifolium Ab.IgE.RAST class|Chamerion angustifolium Ab.IgE.RAST class
C0804067|T201|COMP|21273-8|LNC|Linum usitatissimum Ab.IgE.RAST class|Linum usitatissimum Ab.IgE.RAST class
C0804068|T201|COMP|21274-6|LNC|Flounder Ab.IgG.RAST class|Flounder Ab.IgG.RAST class
C0804070|T201|COMP|21276-1|LNC|Follitropin^1H post XXX challenge|Follitropin^1H post XXX challenge
C0804073|T201|COMP|21279-5|LNC|Follitropin^1.5H post XXX challenge|Follitropin^1.5H post XXX challenge
C0804074|T201|COMP|21280-3|LNC|Fonofos|Fonofos
C0804075|T201|COMP|21281-1|LNC|Fusarium oxysporum Ab.IgE.RAST class|Fusarium oxysporum Ab.IgE.RAST class
C0804076|T201|COMP|21282-9|LNC|Ganglioside GD1a Ab.IgM|Ganglioside GD1a Ab.IgM
C0804077|T201|COMP|21283-7|LNC|Ganglioside GD1a Ab.IgG|Ganglioside GD1a Ab.IgG
C0804078|T201|COMP|21284-5|LNC|Gardnerella vaginalis|Gardnerella vaginalis
C0804079|T201|COMP|21285-2|LNC|Allium sativum Ab.IgG.RAST class|Allium sativum Ab.IgG.RAST class
C0804080|T201|COMP|21286-0|LNC|Gastrin^1.5H post 0.2 U/kg secretin|Gastrin^1.5H post 0.2 U/kg secretin
C0804081|T201|COMP|21287-8|LNC|Gastrin^1H post 0.2 U/kg secretin|Gastrin^1H post 0.2 U/kg secretin
C0804082|T201|COMP|21288-6|LNC|Gastrin^2.5H post 0.2 U/kg secretin|Gastrin^2.5H post 0.2 U/kg secretin
C0804083|T201|COMP|21289-4|LNC|Gastrin^2H post 0.2 U/kg secretin|Gastrin^2H post 0.2 U/kg secretin
C0804084|T201|COMP|21290-2|LNC|Gastrin^3.5H post 0.2 U/kg secretin|Gastrin^3.5H post 0.2 U/kg secretin
C0804085|T201|COMP|21291-0|LNC|Gastrin^3H post 0.2 U/kg secretin|Gastrin^3H post 0.2 U/kg secretin
C0804086|T201|COMP|21292-8|LNC|Gastrin^40M post 0.2 U/kg secretin|Gastrin^40M post 0.2 U/kg secretin
C0804087|T201|COMP|21293-6|LNC|Gastrin^45M post 0.2 U/kg secretin|Gastrin^45M post 0.2 U/kg secretin
C0804088|T201|COMP|21294-4|LNC|Gastrin^4H post 0.2 U/kg secretin|Gastrin^4H post 0.2 U/kg secretin
C0804089|T201|COMP|21295-1|LNC|Gastrin^50M post 0.2 U/kg secretin|Gastrin^50M post 0.2 U/kg secretin
C0804090|T201|COMP|21296-9|LNC|Gastrin^7M post 0.2 U/kg secretin|Gastrin^7M post 0.2 U/kg secretin
C0804091|T201|COMP|21297-7|LNC|Gelatin bovine Ab.IgE.RAST class|Gelatin bovine Ab.IgE.RAST class
C0804092|T201|COMP|21298-5|LNC|Gelatin porcine Ab.IgE.RAST class|Gelatin porcine Ab.IgE.RAST class
C0804094|T201|COMP|21300-9|LNC|Giardia lamblia Ab.IgA|Giardia lamblia Ab.IgA
C0804095|T201|COMP|21301-7|LNC|Giardia lamblia Ab.IgM|Giardia lamblia Ab.IgM
C0804096|T201|COMP|21302-5|LNC|Giardia lamblia Ag^2nd specimen|Giardia lamblia Ag^2nd specimen
C0804097|T201|COMP|21303-3|LNC|Giardia lamblia Ag^3rd specimen|Giardia lamblia Ag^3rd specimen
C0804098|T201|COMP|21304-1|LNC|Zingiber officinale Ab.IgG.RAST class|Zingiber officinale Ab.IgG.RAST class
C0804099|T201|COMP|21305-8|LNC|Glucose|Glucose
C0804100|T201|COMP|21306-6|LNC|Glucose|Glucose
C0804101|T201|COMP|21307-4|LNC|Glucose|Glucose
C0804102|T201|COMP|21308-2|LNC|Glucose^105M post XXX challenge|Glucose^105M post XXX challenge
C0804103|T201|COMP|21309-0|LNC|Glucose^45M post XXX challenge|Glucose^45M post XXX challenge
C0804104|T201|COMP|21310-8|LNC|Glucose^75M post XXX challenge|Glucose^75M post XXX challenge
C0804105|T201|COMP|21311-6|LNC|Gluten Ab.IgG.RAST class|Gluten Ab.IgG.RAST class
C0804106|T201|COMP|21312-4|LNC|Gold|Gold
C0804107|T201|COMP|21313-2|LNC|Grain elevator dust Ab.IgE.RAST class|Grain elevator dust Ab.IgE.RAST class
C0804108|T201|COMP|21314-0|LNC|Vitis vinifera Ab.IgG.RAST class|Vitis vinifera Ab.IgG.RAST class
C0804109|T201|COMP|21315-7|LNC|Citrus paradisis Ab.IgG.RAST class|Citrus paradisis Ab.IgG.RAST class
C0804110|T201|COMP|21316-5|LNC|Grepafloxacin|Grepafloxacin
C0804112|T201|COMP|15552-3|LNC|Baccharis spp Ab.IgE.RAST class|Baccharis spp Ab.IgE.RAST class
C0804113|T201|COMP|21319-9|LNC|Melanogrammus aeglefinus Ab.IgG.RAST class|Melanogrammus aeglefinus Ab.IgG.RAST class
C0804114|T201|COMP|21320-7|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C0804115|T201|COMP|21321-5|LNC|Hippoglossus hippoglossus Ab.IgG.RAST class|Hippoglossus hippoglossus Ab.IgG.RAST class
C0804116|T201|COMP|21322-3|LNC|Hantavirus puumala Ab.IgG|Hantavirus puumala Ab.IgG
C0804117|T201|COMP|21323-1|LNC|Hantavirus puumala Ab.IgM|Hantavirus puumala Ab.IgM
C0804118|T201|COMP|21324-9|LNC|Helminthosporium sativum Ab.IgE.RAST class|Helminthosporium sativum Ab.IgE.RAST class
C0804119|T201|COMP|15768-5|LNC|Helminthosporium sp Ab.IgE.RAST class|Helminthosporium sp Ab.IgE.RAST class
C0804120|T201|COMP|21326-4|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C0804121|T201|COMP|21327-2|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C0804122|T201|COMP|21328-0|LNC|Beta-N-acetylhexosaminidase A & B|Beta-N-acetylhexosaminidase A & B
C0804123|T201|COMP|21329-8|LNC|Carya ovata Ab.IgE.RAST class|Carya ovata Ab.IgE.RAST class
C0804124|T201|COMP|21330-6|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0804125|T201|COMP|21331-4|LNC|HIV 1 p24 Ab|HIV 1 p24 Ab
C0804126|T201|COMP|21332-2|LNC|HIV 1 p41 Ab|HIV 1 p41 Ab
C0804127|T201|COMP|21333-0|LNC|HIV 1 RNA|HIV 1 RNA
C0804128|T201|COMP|21334-8|LNC|HIV 2 gp105 Ab|HIV 2 gp105 Ab
C0804129|T201|COMP|21335-5|LNC|HIV 2 gp120 Ab|HIV 2 gp120 Ab
C0804130|T201|COMP|21336-3|LNC|HIV 2 gp15 Ab|HIV 2 gp15 Ab
C0804131|T201|COMP|21337-1|LNC|HIV 2 gp34 Ab|HIV 2 gp34 Ab
C0804132|T201|COMP|21338-9|LNC|HIV 2 p31 Ab|HIV 2 p31 Ab
C0804133|T201|COMP|21339-7|LNC|HIV 2 p55 Ab|HIV 2 p55 Ab
C0804134|T201|COMP|21340-5|LNC|HIV 2 p58 Ab|HIV 2 p58 Ab
C0804135|T201|COMP|21341-3|LNC|HLA-DR locus|HLA-DR locus
C0804136|T201|COMP|21342-1|LNC|HLA-DR locus 2|HLA-DR locus 2
C0804137|T201|COMP|21343-9|LNC|HLA-DR+DQ|HLA-DR+DQ
C0804138|T201|COMP|21344-7|LNC|House dust Greer Ab.IgG.RAST class|House dust Greer Ab.IgG.RAST class
C0804139|T201|COMP|21345-4|LNC|HTLV I+II Ab|HTLV I+II Ab
C0804140|T201|COMP|21346-2|LNC|HTLV I+II Ab band pattern|HTLV I+II Ab band pattern
C0804141|T201|COMP|21347-0|LNC|HTLV I+II Ab band pattern|HTLV I+II Ab band pattern
C0804142|T201|COMP|21348-8|LNC|HTLV I+II Ab.IgG|HTLV I+II Ab.IgG
C0804143|T201|COMP|21349-6|LNC|IgA|IgA
C0804144|T201|COMP|21350-4|LNC|IgG|IgG
C0804145|T201|COMP|21351-2|LNC|IgM|IgM
C0804146|T201|COMP|21352-0|LNC|Intercellular substance Ab.IgG|Intercellular substance Ab.IgG
C0804147|T201|COMP|21353-8|LNC|Juniperus occidentalis Ab.IgE.RAST class|Juniperus occidentalis Ab.IgE.RAST class
C0804148|T201|COMP|21354-6|LNC|Karaya gum Ab.IgE.RAST class|Karaya gum Ab.IgE.RAST class
C0804149|T201|COMP|21355-3|LNC|Ketones^2.5H post XXX challenge|Ketones^2.5H post XXX challenge
C0804150|T201|COMP|21356-1|LNC|Ketones^3.5H post XXX challenge|Ketones^3.5H post XXX challenge
C0804151|T201|COMP|21357-9|LNC|Ketones^1.5H post XXX challenge|Ketones^1.5H post XXX challenge
C0804152|T201|COMP|21358-7|LNC|Lactalbumin alpha Ab.IgG.RAST class|Lactalbumin alpha Ab.IgG.RAST class
C0804153|T201|COMP|21359-5|LNC|Beta galactosidase Ab.IgE.RAST class|Beta galactosidase Ab.IgE.RAST class
C0804154|T201|COMP|21360-3|LNC|Lamb Ab.IgG.RAST class|Lamb Ab.IgG.RAST class
C0804155|T201|COMP|21361-1|LNC|Laxatives present|Laxatives present
C0804156|T201|COMP|21362-9|LNC|Legionella pneumophila Ab.IgG|Legionella pneumophila Ab.IgG
C0804157|T201|COMP|21363-7|LNC|Legionella pneumophila DNA|Legionella pneumophila DNA
C0804158|T201|COMP|21364-5|LNC|Citrus limon Ab.IgG.RAST class|Citrus limon Ab.IgG.RAST class
C0804159|T201|COMP|21365-2|LNC|Leptin|Leptin
C0804160|T201|COMP|21366-0|LNC|Lactuca sativa Ab.IgG.RAST class|Lactuca sativa Ab.IgG.RAST class
C0804161|T201|COMP|21367-8|LNC|levoFLOXacin|levoFLOXacin
C0804162|T201|COMP|21368-6|LNC|levoFLOXacin|levoFLOXacin
C0804163|T201|COMP|21369-4|LNC|Glycyrrhiza lepidota Ab.IgE.RAST class|Glycyrrhiza lepidota Ab.IgE.RAST class
C0804164|T201|COMP|21370-2|LNC|Citrus aurantifolia Ab.IgG.RAST class|Citrus aurantifolia Ab.IgG.RAST class
C0804165|T201|COMP|21371-0|LNC|Homarus gammarus Ab.IgG.RAST class|Homarus gammarus Ab.IgG.RAST class
C0804166|T201|COMP|21372-8|LNC|Lymphocytes.abnormal/100 leukocytes|Lymphocytes.abnormal/100 leukocytes
C0804167|T201|COMP|21373-6|LNC|Lymphocytes.abnormal/100 leukocytes|Lymphocytes.abnormal/100 leukocytes
C0804168|T201|COMP|21374-4|LNC|Cells.CD8+CD38+|Cells.CD8+CD38+
C0804169|T201|COMP|21375-1|LNC|Lymphocytes.kappa/Lymphocytes.lambda|Lymphocytes.kappa/Lymphocytes.lambda
C0804170|T201|COMP|21376-9|LNC|Macadamia spp Ab.IgE.RAST class|Macadamia spp Ab.IgE.RAST class
C0804171|T201|COMP|21377-7|LNC|Magnesium|Magnesium
C0804172|T201|COMP|21378-5|LNC|Malathion|Malathion
C0804173|T201|COMP|21379-3|LNC|Malt Ab.IgG.RAST class|Malt Ab.IgG.RAST class
C0804174|T201|COMP|21380-1|LNC|Prolactin|Prolactin
C0804175|T201|COMP|21381-9|LNC|Prolactin^1.5H post XXX challenge|Prolactin^1.5H post XXX challenge
C0804176|T201|COMP|21382-7|LNC|Manganese|Manganese
C0804177|T201|COMP|21383-5|LNC|Mercury|Mercury
C0804178|T201|COMP|21384-3|LNC|Mesothelial cells|Mesothelial cells
C0804179|T201|COMP|21385-0|LNC|Metasystox|Metasystox
C0804180|T201|COMP|21386-8|LNC|Methamphetamine|Methamphetamine
C0804181|T201|COMP|21387-6|LNC|Methylhippurate|Methylhippurate
C0804182|T201|COMP|21388-4|LNC|Mevinphos|Mevinphos
C0804183|T201|COMP|21389-2|LNC|Saccharopolyspora rectivirgula Ab.IgE|Saccharopolyspora rectivirgula Ab.IgE
C0804184|T201|COMP|21390-0|LNC|Saccharopolyspora rectivirgula Ab.IgE.RAST class|Saccharopolyspora rectivirgula Ab.IgE.RAST class
C0804186|T201|COMP|15849-3|LNC|Panicum milliaceum Ab.IgE.RAST class|Panicum milliaceum Ab.IgE.RAST class
C0804187|T201|COMP|21393-4|LNC|Monkey epithelium Ab.IgE.RAST class|Monkey epithelium Ab.IgE.RAST class
C0804188|T201|COMP|21394-2|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C0804189|T201|COMP|21395-9|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C0804190|T201|COMP|21396-7|LNC|Mononuclear cells|Mononuclear cells
C0804191|T201|COMP|21397-5|LNC|Mononuclear cells|Mononuclear cells
C0804192|T201|COMP|21398-3|LNC|Mononuclear cells|Mononuclear cells
C0804193|T201|COMP|21399-1|LNC|Broussonetia papyrifera Ab.IgE.RAST class|Broussonetia papyrifera Ab.IgE.RAST class
C0804194|T201|COMP|21400-7|LNC|Morus rubra Ab.IgE.RAST class|Morus rubra Ab.IgE.RAST class
C0804195|T201|COMP|21401-5|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0804196|T201|COMP|21402-3|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C0804197|T201|COMP|21403-1|LNC|Agaricus hortensis Ab.IgG.RAST class|Agaricus hortensis Ab.IgG.RAST class
C0804198|T201|COMP|21404-9|LNC|Mustard Ab.IgG.RAST class|Mustard Ab.IgG.RAST class
C0804199|T201|COMP|21405-6|LNC|Mycobacterium sp DNA|Mycobacterium sp DNA
C0804200|T201|COMP|21406-4|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C0804201|T201|COMP|21407-2|LNC|Myelin Ab.IgA|Myelin Ab.IgA
C0804202|T201|COMP|21408-0|LNC|Myelin Ab.IgG|Myelin Ab.IgG
C0804203|T201|COMP|21409-8|LNC|Myelin Ab.IgM|Myelin Ab.IgM
C0804204|T201|COMP|21410-6|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C0804205|T201|COMP|21411-4|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C0804206|T201|COMP|21412-2|LNC|Myocardium Ab pattern|Myocardium Ab pattern
C0804207|T201|COMP|21413-0|LNC|N-Acetylgalactosamine-4-Sulfatase|N-Acetylgalactosamine-4-Sulfatase
C0804208|T201|COMP|21414-8|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C0804209|T201|COMP|21415-5|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C0804210|T201|COMP|21416-3|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C0804211|T201|COMP|21417-1|LNC|Neurokinin A|Neurokinin A
C0804212|T201|COMP|21418-9|LNC|Neutrophil Ab|Neutrophil Ab
C0804213|T201|COMP|21419-7|LNC|Neutrophil cytoplasmic Ab pattern|Neutrophil cytoplasmic Ab pattern
C0804214|T201|COMP|21420-5|LNC|Nitrate|Nitrate
C0804215|T201|COMP|21421-3|LNC|Norketamine|Norketamine
C0804216|T201|COMP|21422-1|LNC|Normetanephrine|Normetanephrine
C0804217|T201|COMP|21423-9|LNC|Nuclear Ab|Nuclear Ab
C0804218|T201|COMP|21424-7|LNC|Nuclear Ab.IgG|Nuclear Ab.IgG
C0804219|T201|COMP|21425-4|LNC|Nutmeg Ab.IgG.RAST class|Nutmeg Ab.IgG.RAST class
C0804220|T201|COMP|21426-2|LNC|Avena sativa Ab.IgG.RAST class|Avena sativa Ab.IgG.RAST class
C0804221|T201|COMP|15885-7|LNC|Avena sativa Ab.IgE.RAST class|Avena sativa Ab.IgE.RAST class
C0804222|T201|COMP|21428-8|LNC|Olea europaea Ab.IgE|Olea europaea Ab.IgE
C0804223|T201|COMP|21429-6|LNC|Olea europaea Ab.IgE.RAST class|Olea europaea Ab.IgE.RAST class
C0804224|T201|COMP|21430-4|LNC|Allium cepa Ab.IgG.RAST class|Allium cepa Ab.IgG.RAST class
C0804225|T201|COMP|21431-2|LNC|Opiates|Opiates
C0804226|T201|COMP|21432-0|LNC|Citrus sinensis Ab.IgG.RAST class|Citrus sinensis Ab.IgG.RAST class
C0804227|T201|COMP|21433-8|LNC|Citrus sinensis tree Ab.IgE.RAST class|Citrus sinensis tree Ab.IgE.RAST class
C0804228|T201|COMP|21434-6|LNC|Origanum vulgare Ab.IgG.RAST class|Origanum vulgare Ab.IgG.RAST class
C0804229|T201|COMP|21435-3|LNC|Osteocalcin.bovine|Osteocalcin.bovine
C0804230|T201|COMP|21436-1|LNC|Ovary Ab|Ovary Ab
C0804231|T201|COMP|21437-9|LNC|Oxychlordane|Oxychlordane
C0804232|T201|COMP|21438-7|LNC|Ostrea edulis Ab.IgG.RAST class|Ostrea edulis Ab.IgG.RAST class
C0804233|T201|COMP|21439-5|LNC|Papain Ab.IgE.RAST class|Papain Ab.IgE.RAST class
C0804235|T201|COMP|21441-1|LNC|Human papilloma virus 6+11+42+43+44 DNA|Human papilloma virus 6+11+42+43+44 DNA
C0804236|T201|COMP|21442-9|LNC|Parainfluenza virus identified|Parainfluenza virus identified
C0804237|T201|COMP|21443-7|LNC|Paraoxon|Paraoxon
C0804238|T201|COMP|21444-5|LNC|Petroselinum crispum Ab.IgG.RAST class|Petroselinum crispum Ab.IgG.RAST class
C0804239|T201|COMP|21445-2|LNC|Pisum sativum Ab.IgG.RAST class|Pisum sativum Ab.IgG.RAST class
C0804240|T201|COMP|21446-0|LNC|Prunus persica Ab.IgG.RAST class|Prunus persica Ab.IgG.RAST class
C0804241|T201|COMP|21447-8|LNC|Arachis hypogaea Ab.IgG.RAST class|Arachis hypogaea Ab.IgG.RAST class
C0804242|T201|COMP|21448-6|LNC|Pyrus communis Ab.IgG.RAST class|Pyrus communis Ab.IgG.RAST class
C0804243|T201|COMP|21449-4|LNC|Piper nigrum Ab.IgG.RAST class|Piper nigrum Ab.IgG.RAST class
C0804244|T201|COMP|21450-2|LNC|Pepper cayenne Ab.IgG.RAST class|Pepper cayenne Ab.IgG.RAST class
C0804245|T201|COMP|21451-0|LNC|Capsicum frutescens Ab.IgG.RAST class|Capsicum frutescens Ab.IgG.RAST class
C0804246|T201|COMP|21452-8|LNC|Pepper green Ab.IgG.RAST class|Pepper green Ab.IgG.RAST class
C0804247|T201|COMP|21453-6|LNC|Pepper jalapeno Ab.IgE.RAST class|Pepper jalapeno Ab.IgE.RAST class
C0804248|T201|COMP|21454-4|LNC|Pepper white Ab.IgG.RAST class|Pepper white Ab.IgG.RAST class
C0804249|T201|COMP|21455-1|LNC|Mentha piperita Ab.IgE.RAST class|Mentha piperita Ab.IgE.RAST class
C0804250|T201|COMP|21456-9|LNC|Pheasant Ab.IgE.RAST class|Pheasant Ab.IgE.RAST class
C0804251|T201|COMP|21457-7|LNC|Phorate|Phorate
C0804252|T201|COMP|21458-5|LNC|Phosphate|Phosphate
C0804253|T201|COMP|21459-3|LNC|Salicornia spp Ab.IgE.RAST class|Salicornia spp Ab.IgE.RAST class
C0804254|T201|COMP|21460-1|LNC|Stizostedion vitreum Ab.IgE.RAST class|Stizostedion vitreum Ab.IgE.RAST class
C0804255|T201|COMP|21461-9|LNC|(Pinus contorta+Pinus ponderosa ) Ab.IgE|(Pinus contorta+Pinus ponderosa ) Ab.IgE
C0804257|T201|COMP|21463-5|LNC|Ananas comosus Ab.IgG.RAST class|Ananas comosus Ab.IgG.RAST class
C0804258|T201|COMP|21464-3|LNC|Plasminogen activator urokinase type|Plasminogen activator urokinase type
C0804259|T201|COMP|21465-0|LNC|Plasmodium falciparum Ab|Plasmodium falciparum Ab
C0804260|T201|COMP|21466-8|LNC|Plasmodium malariae Ab|Plasmodium malariae Ab
C0804261|T201|COMP|21467-6|LNC|Plasmodium ovale Ab|Plasmodium ovale Ab
C0804262|T201|COMP|21468-4|LNC|Plasmodium vivax Ab|Plasmodium vivax Ab
C0804263|T201|COMP|21469-2|LNC|Prunus domestica Ab.IgG.RAST class|Prunus domestica Ab.IgG.RAST class
C0804264|T201|COMP|21470-0|LNC|Pollachius virens Ab.IgE.RAST class|Pollachius virens Ab.IgE.RAST class
C0804265|T201|COMP|21471-8|LNC|Punica granatum Ab.IgE|Punica granatum Ab.IgE
C0804266|T201|COMP|21472-6|LNC|Punica granatum Ab.IgE.RAST class|Punica granatum Ab.IgE.RAST class
C0804267|T201|COMP|21473-4|LNC|Populus alba Ab.IgE|Populus alba Ab.IgE
C0804268|T201|COMP|21474-2|LNC|Populus alba Ab.IgE.RAST class|Populus alba Ab.IgE.RAST class
C0804269|T201|COMP|21475-9|LNC|Pork Ab.IgG.RAST class|Pork Ab.IgG.RAST class
C0804270|T201|COMP|21476-7|LNC|Potassium|Potassium
C0804271|T201|COMP|6220-8|LNC|Solanum tuberosum Ab.IgE|Solanum tuberosum Ab.IgE
C0804272|T201|COMP|15957-4|LNC|Solanum tuberosum Ab.IgE.RAST class|Solanum tuberosum Ab.IgE.RAST class
C0804273|T201|COMP|21479-1|LNC|Solanum tuberosum Ab.IgG.RAST class|Solanum tuberosum Ab.IgG.RAST class
C0804274|T201|COMP|21480-9|LNC|Propoxur|Propoxur
C0804275|T201|COMP|21481-7|LNC|Propranolol|Propranolol
C0804276|T201|COMP|21482-5|LNC|Protein|Protein
C0804277|T201|COMP|21483-3|LNC|quiNIDine^peak|quiNIDine^peak
C0804279|T201|COMP|21485-8|LNC|Raphanus sativus Ab.IgG.RAST class|Raphanus sativus Ab.IgG.RAST class
C0804280|T201|COMP|21486-6|LNC|Brassica napus pollen Ab.IgE.RAST class|Brassica napus pollen Ab.IgE.RAST class
C0804281|T201|COMP|21487-4|LNC|Ribosomal P Ab|Ribosomal P Ab
C0804282|T201|COMP|21488-2|LNC|Oryza sativa Ab.IgG.RAST class|Oryza sativa Ab.IgG.RAST class
C0804283|T201|COMP|21489-0|LNC|Rickettsia (Proteus OX19) Ab|Rickettsia (Proteus OX19) Ab
C0804284|T201|COMP|21490-8|LNC|Rickettsia (Proteus OX2) Ab|Rickettsia (Proteus OX2) Ab
C0804285|T201|COMP|21491-6|LNC|Rickettsia (Proteus OXK) Ab|Rickettsia (Proteus OXK) Ab
C0804286|T201|COMP|21492-4|LNC|Rickettsia conorii Ab.IgG|Rickettsia conorii Ab.IgG
C0804287|T201|COMP|21493-2|LNC|Rickettsia conorii Ab.IgM|Rickettsia conorii Ab.IgM
C0804288|T201|COMP|21494-0|LNC|Rickettsia spotted fever group Ab.IgG|Rickettsia spotted fever group Ab.IgG
C0804289|T201|COMP|21495-7|LNC|Rickettsia spotted fever group Ab.IgM|Rickettsia spotted fever group Ab.IgM
C0804290|T201|COMP|21496-5|LNC|Rickettsia typhus group Ab.IgG|Rickettsia typhus group Ab.IgG
C0804291|T201|COMP|21497-3|LNC|Rickettsia typhus group Ab.IgM|Rickettsia typhus group Ab.IgM
C0804292|T201|COMP|21498-1|LNC|Orientia tsutsugamushi Ab.IgG|Orientia tsutsugamushi Ab.IgG
C0804293|T201|COMP|21499-9|LNC|Hoplostethus atlanticus Ab.IgE.RAST class|Hoplostethus atlanticus Ab.IgE.RAST class
C0804294|T201|COMP|21500-4|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0804295|T201|COMP|21501-2|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0804296|T201|COMP|21502-0|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C0804297|T201|COMP|21503-8|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C0804298|T201|COMP|21505-3|LNC|Secale cereale Ab.IgG.RAST class|Secale cereale Ab.IgG.RAST class
C0804300|T201|COMP|21506-1|LNC|Carthamus tinctorius Ab.IgG.RAST class|Carthamus tinctorius Ab.IgG.RAST class
C0804301|T201|COMP|21507-9|LNC|Salvia officinalis Ab.IgG.RAST class|Salvia officinalis Ab.IgG.RAST class
C0804302|T201|COMP|21508-7|LNC|Artemisia californica Ab.IgE.RAST class|Artemisia californica Ab.IgE.RAST class
C0804303|T201|COMP|21509-5|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C0804304|T201|COMP|21510-3|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C0804305|T201|COMP|21511-1|LNC|Salmonella paratyphi A H Ab|Salmonella paratyphi A H Ab
C0804306|T201|COMP|21512-9|LNC|Salmonella paratyphi A H Ab|Salmonella paratyphi A H Ab
C0804307|T201|COMP|21513-7|LNC|Salmonella paratyphi B H Ab|Salmonella paratyphi B H Ab
C0804308|T201|COMP|21514-5|LNC|Salmonella paratyphi B H Ab|Salmonella paratyphi B H Ab
C0804309|T201|COMP|21515-2|LNC|Saltbush annual Ab.IgE.RAST class|Saltbush annual Ab.IgE.RAST class
C0804310|T201|COMP|21516-0|LNC|Pecten spp Ab.IgG.RAST class|Pecten spp Ab.IgG.RAST class
C0804311|T201|COMP|21517-8|LNC|Schistosoma sp Ab.IgE.RAST class|Schistosoma sp Ab.IgE.RAST class
C0804312|T201|COMP|21518-6|LNC|SCL-70 extractable nuclear Ab.IgG|SCL-70 extractable nuclear Ab.IgG
C0804313|T201|COMP|21519-4|LNC|Sesamum indicum Ab.IgG.RAST class|Sesamum indicum Ab.IgG.RAST class
C0804314|T201|COMP|21520-2|LNC|Shark Ab.IgE.RAST class|Shark Ab.IgE.RAST class
C0804315|T201|COMP|21521-0|LNC|Pandalus borealis Ab.IgG.RAST class|Pandalus borealis Ab.IgG.RAST class
C0804317|T201|COMP|21523-6|LNC|Smith extractable nuclear Ab.IgG|Smith extractable nuclear Ab.IgG
C0804318|T201|COMP|21524-4|LNC|Snapper red Ab.IgG.RAST class|Snapper red Ab.IgG.RAST class
C0804319|T201|COMP|21525-1|LNC|Sodium|Sodium
C0804320|T201|COMP|21526-9|LNC|Sodium|Sodium
C0804321|T201|COMP|21527-7|LNC|Sodium|Sodium
C0804322|T201|COMP|21528-5|LNC|Solea solea Ab.IgG.RAST class|Solea solea Ab.IgG.RAST class
C0804323|T201|COMP|21529-3|LNC|Specimen volume|Specimen volume
C0804324|T201|COMP|21530-1|LNC|Specimen volume|Specimen volume
C0804330|T201|COMP|21536-8|LNC|Acid sphingomyelinase|Acid sphingomyelinase
C0804331|T201|COMP|21537-6|LNC|Spinacia oleracea Ab.IgG.RAST class|Spinacia oleracea Ab.IgG.RAST class
C0804332|T201|COMP|21538-4|LNC|Picea pungens Ab.IgE.RAST class|Picea pungens Ab.IgE.RAST class
C0804333|T201|COMP|21539-2|LNC|Squash summer Ab.IgE.RAST class|Squash summer Ab.IgE.RAST class
C0804334|T201|COMP|21540-0|LNC|Squash zucchini Ab.IgE.RAST class|Squash zucchini Ab.IgE.RAST class
C0804335|T201|COMP|21541-8|LNC|Squash zucchini Ab.IgG.RAST class|Squash zucchini Ab.IgG.RAST class
C0804336|T201|COMP|21542-6|LNC|Fragaria vesca Ab.IgG.RAST class|Fragaria vesca Ab.IgG.RAST class
C0804337|T201|COMP|21543-4|LNC|Saccharum officinarum Ab.IgG.RAST class|Saccharum officinarum Ab.IgG.RAST class
C0804338|T201|COMP|21544-2|LNC|Sulfamethoxazole Ab.IgE.RAST class|Sulfamethoxazole Ab.IgE.RAST class
C0804339|T201|COMP|21545-9|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C0804340|T201|COMP|21546-7|LNC|Sulfatide Ab.IgM|Sulfatide Ab.IgM
C0804341|T201|COMP|21547-5|LNC|Helianthus annuus seed Ab.IgG.RAST class|Helianthus annuus seed Ab.IgG.RAST class
C0804342|T201|COMP|21548-3|LNC|Ipomoea batatas Ab.IgG.RAST class|Ipomoea batatas Ab.IgG.RAST class
C0804343|T201|COMP|15761-0|LNC|Liquidambar styraciflua Ab.IgE.RAST class|Liquidambar styraciflua Ab.IgE.RAST class
C0804344|T201|COMP|21550-9|LNC|Synovial lining cells|Synovial lining cells
C0804345|T201|COMP|21551-7|LNC|t(15;17)(q24.1;q21.1)(PML,RARA) fusion transcript|t(15;17)(q24.1;q21.1)(PML,RARA) fusion transcript
C0804346|T201|COMP|21552-5|LNC|Citrus reticulata Ab.IgG.RAST class|Citrus reticulata Ab.IgG.RAST class
C0804347|T201|COMP|21553-3|LNC|Camellia sinensis Ab.IgG.RAST class|Camellia sinensis Ab.IgG.RAST class
C0804348|T201|COMP|21554-1|LNC|Terbufos|Terbufos
C0804350|T201|COMP|21556-6|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0804351|T201|COMP|21557-4|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0804352|T201|COMP|21558-2|LNC|Thallium|Thallium
C0804353|T201|COMP|21559-0|LNC|Theophylline|Theophylline
C0804354|T201|COMP|21560-8|LNC|Thermoactinomyces candidus Ab|Thermoactinomyces candidus Ab
C0804355|T201|COMP|21561-6|LNC|Thermoactinomyces sacchari Ab|Thermoactinomyces sacchari Ab
C0804356|T201|COMP|21562-4|LNC|Thiocyanate/Creatinine|Thiocyanate/Creatinine
C0804357|T201|COMP|21563-2|LNC|Thiopurine methyltransferase|Thiopurine methyltransferase
C0804358|T201|COMP|21564-0|LNC|Thiosulfate|Thiosulfate
C0804359|T201|COMP|21565-7|LNC|tiaGABine|tiaGABine
C0804360|T201|COMP|21566-5|LNC|TOLAZamide|TOLAZamide
C0804361|T201|COMP|21567-3|LNC|TOLBUTamide|TOLBUTamide
C0804362|T201|COMP|21568-1|LNC|Lycopersicon lycopersicum Ab.IgG.RAST class|Lycopersicon lycopersicum Ab.IgG.RAST class
C0804363|T201|COMP|21569-9|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0804364|T201|COMP|21570-7|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0804365|T201|COMP|21571-5|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0804372|T201|COMP|21578-0|LNC|Ailanthus altissima Ab.IgE.RAST class|Ailanthus altissima Ab.IgE.RAST class
C0804373|T201|COMP|21579-8|LNC|Trichloroethylene|Trichloroethylene
C0804374|T201|COMP|21580-6|LNC|Trimethobenzamide|Trimethobenzamide
C0804375|T201|COMP|21581-4|LNC|Oncorhynchus mykiss Ab.IgG.RAST class|Oncorhynchus mykiss Ab.IgG.RAST class
C0804376|T201|COMP|21582-2|LNC|Tryptase|Tryptase
C0804377|T201|COMP|21583-0|LNC|Turkey Ab.IgG.RAST class|Turkey Ab.IgG.RAST class
C0804378|T201|COMP|21584-8|LNC|Turkey feather Ab.IgE.RAST class|Turkey feather Ab.IgE.RAST class
C0804379|T201|COMP|21585-5|LNC|Uranium|Uranium
C0804380|T201|COMP|21586-3|LNC|Uranium|Uranium
C0804381|T201|COMP|21587-1|LNC|Urate|Urate
C0804382|T201|COMP|21588-9|LNC|Urobilinogen|Urobilinogen
C0804383|T201|COMP|21589-7|LNC|Ustilago nuda+Ustilago tritici Ab.IgE.RAST class|Ustilago nuda+Ustilago tritici Ab.IgE.RAST class
C0804384|T201|COMP|21590-5|LNC|Valproate.bound/Valproate.total|Valproate.bound/Valproate.total
C0804385|T201|COMP|21591-3|LNC|Vanilla planifolia Ab.IgG.RAST class|Vanilla planifolia Ab.IgG.RAST class
C0804386|T201|COMP|21592-1|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C0804387|T201|COMP|21594-7|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C0804388|T201|COMP|21595-4|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0804389|T201|COMP|21596-2|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0804390|T201|COMP|21597-0|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0804391|T201|COMP|21598-8|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C0804392|T201|COMP|21599-6|LNC|Venison Ab.IgE.RAST class|Venison Ab.IgE.RAST class
C0804393|T201|COMP|21600-2|LNC|Juglans regia Ab.IgE.RAST class|Juglans regia Ab.IgE.RAST class
C0804394|T201|COMP|21601-0|LNC|Citrullus lanatus Ab.IgG.RAST class|Citrullus lanatus Ab.IgG.RAST class
C0804395|T201|COMP|21602-8|LNC|Triticum aestivum Ab.IgG.RAST class|Triticum aestivum Ab.IgG.RAST class
C0804396|T201|COMP|21603-6|LNC|Wheat dust Ab.IgE|Wheat dust Ab.IgE
C0804397|T201|COMP|21604-4|LNC|Wheat dust Ab.IgE.RAST class|Wheat dust Ab.IgE.RAST class
C0804398|T201|COMP|21605-1|LNC|Whitefish Ab.IgG.RAST class|Whitefish Ab.IgG.RAST class
C0804399|T201|COMP|21606-9|LNC|Xylose^2nd specimen post XXX challenge|Xylose^2nd specimen post XXX challenge
C0804400|T201|COMP|21607-7|LNC|Saccharomyces cerevisiae Ab.IgG.RAST class|Saccharomyces cerevisiae Ab.IgG.RAST class
C0804401|T201|COMP|21608-5|LNC|Yeast brewer's Ab.IgG.RAST class|Yeast brewer's Ab.IgG.RAST class
C0804402|T201|COMP|21609-3|LNC|Yogurt Ab.IgE.RAST class|Yogurt Ab.IgE.RAST class
C0804403|T201|COMP|21610-1|LNC|Zinc|Zinc
C0804404|T201|COMP|21611-9|LNC|Age|Age
C0804405|T201|COMP|21612-7|LNC|Age|Age
C0804406|T201|COMP|21613-5|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0804407|T201|COMP|21614-3|LNC|CDKN2A gene deletion|CDKN2A gene deletion
C0804408|T201|COMP|21615-0|LNC|CDKN2B gene deletion|CDKN2B gene deletion
C0804409|T201|COMP|21617-6|LNC|APC gene.p.Ile1307Lys|APC gene.p.Ile1307Lys
C0804410|T201|COMP|21618-4|LNC|APC gene mutations tested for|APC gene mutations tested for
C0804411|T201|COMP|21619-2|LNC|APOE gene targeted mutation analysis|APOE gene targeted mutation analysis
C0804412|T201|COMP|21620-0|LNC|STS gene deletion|STS gene deletion
C0804413|T201|COMP|21622-6|LNC|ASPA gene.p.Glu285Ala|ASPA gene.p.Glu285Ala
C0804414|T201|COMP|21623-4|LNC|ASPA gene mutations tested for|ASPA gene mutations tested for
C0804415|T201|COMP|21624-2|LNC|ATM gene targeted mutation analysis|ATM gene targeted mutation analysis
C0804416|T201|COMP|21625-9|LNC|ATM gene mutations tested for|ATM gene mutations tested for
C0804417|T201|COMP|21626-7|LNC|ATP7B gene targeted mutation analysis|ATP7B gene targeted mutation analysis
C0804418|T201|COMP|21627-5|LNC|ATP7B gene.c.2010_2016del|ATP7B gene.c.2010_2016del
C0804419|T201|COMP|21628-3|LNC|ATP7B gene.c.2337delC|ATP7B gene.c.2337delC
C0804420|T201|COMP|21629-1|LNC|ATP7B gene.c.2487insT|ATP7B gene.c.2487insT
C0804421|T201|COMP|21630-9|LNC|ATP7B gene.c.1711G>C|ATP7B gene.c.1711G>C
C0804422|T201|COMP|21631-7|LNC|ATP7B gene.p.Gly1267Arg|ATP7B gene.p.Gly1267Arg
C0804423|T201|COMP|21632-5|LNC|ATP7B gene.p.His1070Gln|ATP7B gene.p.His1070Gln
C0804424|T201|COMP|21633-3|LNC|ATP7B gene.p.His714Gln|ATP7B gene.p.His714Gln
C0804425|T201|COMP|21634-1|LNC|ATP7B gene.p.Asn915Ser|ATP7B gene.p.Asn915Ser
C0804426|T201|COMP|21635-8|LNC|ATP7B gene.p.Arg778Leu|ATP7B gene.p.Arg778Leu
C0804427|T201|COMP|21636-6|LNC|BRCA1 gene targeted mutation analysis|BRCA1 gene targeted mutation analysis
C0804428|T201|COMP|21637-4|LNC|BRCA1 gene.c.185delAG|BRCA1 gene.c.185delAG
C0804429|T201|COMP|21638-2|LNC|BRCA1 gene.c.5382insC|BRCA1 gene.c.5382insC
C0804430|T201|COMP|21639-0|LNC|BRCA1 gene mutations tested for|BRCA1 gene mutations tested for
C0804431|T201|COMP|21640-8|LNC|BRCA2 gene.c.6174delT|BRCA2 gene.c.6174delT
C0804432|T201|COMP|21641-6|LNC|CACNA1S gene targeted mutation analysis|CACNA1S gene targeted mutation analysis
C0804433|T201|COMP|21642-4|LNC|CACNA1S gene.p.Arg1239Gly|CACNA1S gene.p.Arg1239Gly
C0804434|T201|COMP|21643-2|LNC|CACNA1S gene.p.Arg1239His|CACNA1S gene.p.Arg1239His
C0804435|T201|COMP|21644-0|LNC|CACNA1S gene.p.Arg528His|CACNA1S gene.p.Arg528His
C0804436|T201|COMP|21645-7|LNC|CACNA1S gene mutations tested for|CACNA1S gene mutations tested for
C0804437|T201|COMP|21646-5|LNC|CBS gene targeted mutation analysis|CBS gene targeted mutation analysis
C0804438|T201|COMP|21647-3|LNC|CBS gene.p.G307S|CBS gene.p.G307S
C0804439|T201|COMP|21648-1|LNC|CBS gene.p.I278T|CBS gene.p.I278T
C0804440|T201|COMP|21649-9|LNC|CBS gene mutations tested for|CBS gene mutations tested for
C0804441|T201|COMP|21650-7|LNC|CCR5 gene mutation analysis|CCR5 gene mutation analysis
C0804442|T201|COMP|21651-5|LNC|CCR5 gene mutations tested for|CCR5 gene mutations tested for
C0804443|T201|COMP|21652-3|LNC|CDH1 gene targeted mutation analysis|CDH1 gene targeted mutation analysis
C0804444|T201|COMP|21653-1|LNC|CDH1 gene mutations tested for|CDH1 gene mutations tested for
C0804445|T201|COMP|21655-6|LNC|CFTR gene.p.Phe508del|CFTR gene.p.Phe508del
C0804446|T201|COMP|21656-4|LNC|CFTR gene mutations tested for|CFTR gene mutations tested for
C0804447|T201|COMP|21657-2|LNC|COL2A1 gene targeted mutation analysis|COL2A1 gene targeted mutation analysis
C0804448|T201|COMP|21658-0|LNC|COL2A1 gene mutations tested for|COL2A1 gene mutations tested for
C0804449|T201|COMP|21659-8|LNC|CTNNB1 gene targeted mutation analysis|CTNNB1 gene targeted mutation analysis
C0804450|T201|COMP|21660-6|LNC|CTNNB1 gene mutations tested for|CTNNB1 gene mutations tested for
C0804451|T201|COMP|21661-4|LNC|CYP2D6 gene deletion|CYP2D6 gene deletion
C0804452|T201|COMP|21662-2|LNC|CYP2D6 gene.c.2637delA|CYP2D6 gene.c.2637delA
C0804453|T201|COMP|21663-0|LNC|CYP2D6 gene mutation analysis G-A NT1 X4|CYP2D6 gene mutation analysis G-A NT1 X4
C0804454|T201|COMP|21664-8|LNC|CYP2D6 gene.p.Gly169Ter|CYP2D6 gene.p.Gly169Ter
C0804455|T201|COMP|21665-5|LNC|EGFR gene targeted mutation analysis|EGFR gene targeted mutation analysis
C0804456|T201|COMP|21666-3|LNC|EGFR gene mutations tested for|EGFR gene mutations tested for
C0804457|T201|COMP|21667-1|LNC|F5 gene targeted mutation analysis|F5 gene targeted mutation analysis
C0804458|T201|COMP|21668-9|LNC|F5 gene.p.Arg506Gln|F5 gene.p.Arg506Gln
C0804459|T201|COMP|21669-7|LNC|F5 gene mutations tested for|F5 gene mutations tested for
C0804460|T201|COMP|21670-5|LNC|F7 gene targeted mutation analysis|F7 gene targeted mutation analysis
C0804461|T201|COMP|21671-3|LNC|F7 gene mutations tested for|F7 gene mutations tested for
C0804462|T201|COMP|21672-1|LNC|F8 gene targeted mutation analysis|F8 gene targeted mutation analysis
C0804463|T201|COMP|21673-9|LNC|F8 gene mutations tested for|F8 gene mutations tested for
C0804464|T201|COMP|21674-7|LNC|FGFR2 gene targeted mutation analysis|FGFR2 gene targeted mutation analysis
C0804465|T201|COMP|21675-4|LNC|FGFR2 gene mutations tested for|FGFR2 gene mutations tested for
C0804466|T201|COMP|21676-2|LNC|FGFR3 gene targeted mutation analysis|FGFR3 gene targeted mutation analysis
C0804467|T201|COMP|21677-0|LNC|FGFR3 gene.p.Gly375Cys|FGFR3 gene.p.Gly375Cys
C0804468|T201|COMP|21678-8|LNC|FGFR3 gene.p.Gly380Arg|FGFR3 gene.p.Gly380Arg
C0804469|T201|COMP|21679-6|LNC|FGFR3 gene.p.Lys650Glu|FGFR3 gene.p.Lys650Glu
C0804470|T201|COMP|21680-4|LNC|G6PD gene targeted mutation analysis|G6PD gene targeted mutation analysis
C0804471|T201|COMP|21681-2|LNC|G6PD gene mutations tested for|G6PD gene mutations tested for
C0804472|T201|COMP|21682-0|LNC|Gauchers disease type 1 gene mutations tested for|Gauchers disease type 1 gene mutations tested for
C0804473|T201|COMP|21683-8|LNC|Gauchers disease type 2 gene mutations tested for|Gauchers disease type 2 gene mutations tested for
C0804474|T201|COMP|21684-6|LNC|Gauchers disease type 3 gene mutations tested for|Gauchers disease type 3 gene mutations tested for
C0804475|T201|COMP|21685-3|LNC|HADHB gene targeted mutation analysis|HADHB gene targeted mutation analysis
C0804476|T201|COMP|21686-1|LNC|HADHB gene mutations tested for|HADHB gene mutations tested for
C0804477|T201|COMP|21687-9|LNC|HBA1 gene targeted mutation analysis|HBA1 gene targeted mutation analysis
C0804478|T201|COMP|21688-7|LNC|HBA1 gene mutations tested for|HBA1 gene mutations tested for
C0804479|T201|COMP|21689-5|LNC|HBB gene targeted mutation analysis|HBB gene targeted mutation analysis
C0804480|T201|COMP|21690-3|LNC|HBB gene.p.Glu6Val|HBB gene.p.Glu6Val
C0804481|T201|COMP|21691-1|LNC|HBB gene mutations tested for|HBB gene mutations tested for
C0804482|T201|COMP|21692-9|LNC|PRSS1 gene targeted mutation analysis|PRSS1 gene targeted mutation analysis
C0804483|T201|COMP|21693-7|LNC|Hereditary pancreatitis gene mutations tested for|Hereditary pancreatitis gene mutations tested for
C0804485|T201|COMP|21695-2|LNC|HFE gene.p.Cys282Tyr|HFE gene.p.Cys282Tyr
C0804486|T201|COMP|21696-0|LNC|HFE gene.p.His63Asp|HFE gene.p.His63Asp
C0804487|T201|COMP|21697-8|LNC|HFE gene mutations tested for|HFE gene mutations tested for
C0804488|T201|COMP|21698-6|LNC|HRAS gene targeted mutation analysis|HRAS gene targeted mutation analysis
C0804489|T201|COMP|21699-4|LNC|HRAS gene mutations tested for|HRAS gene mutations tested for
C0804490|T201|COMP|21700-0|LNC|Kallmann syndrome gene targeted mutation analysis|Kallmann syndrome gene targeted mutation analysis
C0804491|T201|COMP|21701-8|LNC|Kallmann syndrome gene mutations tested for|Kallmann syndrome gene mutations tested for
C0804492|T201|COMP|21702-6|LNC|KRAS gene targeted mutation analysis|KRAS gene targeted mutation analysis
C0804493|T201|COMP|21703-4|LNC|KRAS gene mutations tested for|KRAS gene mutations tested for
C0804494|T201|COMP|21704-2|LNC|MT-ATP6 gene targeted mutation analysis|MT-ATP6 gene targeted mutation analysis
C0804495|T201|COMP|21705-9|LNC|MT-ND4 gene.m.11696G>A|MT-ND4 gene.m.11696G>A
C0804496|T201|COMP|21706-7|LNC|MT-ND4 gene.p.R304H|MT-ND4 gene.p.R304H
C0804497|T201|COMP|21707-5|LNC|MT-ND4 gene.p.Thr109Ala|MT-ND4 gene.p.Thr109Ala
C0804498|T201|COMP|21708-3|LNC|MT-ATP6 gene.p.L156R|MT-ATP6 gene.p.L156R
C0804499|T201|COMP|21709-1|LNC|MTHFR gene targeted mutation analysis|MTHFR gene targeted mutation analysis
C0804500|T201|COMP|21710-9|LNC|MTHFR gene.p.Ala677Val|MTHFR gene.p.Ala677Val
C0804501|T201|COMP|21711-7|LNC|MTHFR gene.p.Cys677Glu|MTHFR gene.p.Cys677Glu
C0804502|T201|COMP|21712-5|LNC|MTHFR gene mutations tested for|MTHFR gene mutations tested for
C0804503|T201|COMP|21713-3|LNC|MT-TK gene.m.8344A>G|MT-TK gene.m.8344A>G
C0804504|T201|COMP|21714-1|LNC|MT-TL1 gene.m.3243A>G|MT-TL1 gene.m.3243A>G
C0804505|T201|COMP|21715-8|LNC|MXI1 gene targeted mutation analysis|MXI1 gene targeted mutation analysis
C0804506|T201|COMP|21716-6|LNC|NB gene targeted mutation analysis|NB gene targeted mutation analysis
C0804507|T201|COMP|21717-4|LNC|NF1 gene targeted mutation analysis|NF1 gene targeted mutation analysis
C0804508|T201|COMP|21718-2|LNC|NF1 gene mutations tested for|NF1 gene mutations tested for
C0804509|T201|COMP|21719-0|LNC|NRAS gene targeted mutation analysis|NRAS gene targeted mutation analysis
C0804510|T201|COMP|21720-8|LNC|NRAS gene mutations tested for|NRAS gene mutations tested for
C0804511|T201|COMP|21721-6|LNC|OTC gene targeted mutation analysis|OTC gene targeted mutation analysis
C0804512|T201|COMP|21722-4|LNC|OTC gene mutations tested for|OTC gene mutations tested for
C0804513|T201|COMP|21723-2|LNC|SERPINA1 gene targeted mutation analysis|SERPINA1 gene targeted mutation analysis
C0804514|T201|COMP|21724-0|LNC|SERPINA1 gene.p.Glu264Val|SERPINA1 gene.p.Glu264Val
C0804515|T201|COMP|21725-7|LNC|SERPINA1 gene.p.Glu342Lys|SERPINA1 gene.p.Glu342Lys
C0804516|T201|COMP|21726-5|LNC|SERPINA1 gene mutations tested for|SERPINA1 gene mutations tested for
C0804517|T201|COMP|21727-3|LNC|PMP22 gene targeted mutation analysis|PMP22 gene targeted mutation analysis
C0804518|T201|COMP|21728-1|LNC|PMP22 gene mutations tested for|PMP22 gene mutations tested for
C0804519|T201|COMP|21729-9|LNC|PSAP gene targeted mutation analysis|PSAP gene targeted mutation analysis
C0804520|T201|COMP|21730-7|LNC|PSAP gene mutations tested for|PSAP gene mutations tested for
C0804521|T201|COMP|21731-5|LNC|RB1 gene targeted mutation analysis|RB1 gene targeted mutation analysis
C0804522|T201|COMP|21732-3|LNC|RB1 gene mutations tested for|RB1 gene mutations tested for
C0804523|T201|COMP|21733-1|LNC|RET gene targeted mutation analysis|RET gene targeted mutation analysis
C0804524|T201|COMP|21734-9|LNC|RET gene mutations tested for|RET gene mutations tested for
C0804525|T201|COMP|21735-6|LNC|SNCA gene targeted mutation analysis|SNCA gene targeted mutation analysis
C0804526|T201|COMP|21736-4|LNC|SNCA gene.p.Ala30Pro|SNCA gene.p.Ala30Pro
C0804527|T201|COMP|21737-2|LNC|SNCA gene.p.Ala53Thr|SNCA gene.p.Ala53Thr
C0804528|T201|COMP|21738-0|LNC|SNCA gene mutations tested for|SNCA gene mutations tested for
C0804529|T201|COMP|21739-8|LNC|TP53 gene targeted mutation analysis|TP53 gene targeted mutation analysis
C0804530|T201|COMP|21740-6|LNC|TRAF3 gene targeted mutation analysis|TRAF3 gene targeted mutation analysis
C0804531|T201|COMP|21741-4|LNC|TRAF3 gene mutations tested for|TRAF3 gene mutations tested for
C0804532|T201|COMP|21742-2|LNC|WT1 gene targeted mutation analysis|WT1 gene targeted mutation analysis
C0804533|T201|COMP|21743-0|LNC|WT1 gene mutations tested for|WT1 gene mutations tested for
C0804534|T201|COMP|21744-8|LNC|CCND1 gene rearrangements|CCND1 gene rearrangements
C0804535|T201|COMP|21095-5|LNC|BCL2 gene rearrangements|BCL2 gene rearrangements
C0804536|T201|COMP|21746-3|LNC|BCL6 gene rearrangements|BCL6 gene rearrangements
C0804537|T201|COMP|21747-1|LNC|Immunoglobulin heavy chain gene rearrangements|Immunoglobulin heavy chain gene rearrangements
C0804540|T201|COMP|21750-5|LNC|MYC gene rearrangements|MYC gene rearrangements
C0804541|T201|COMP|21751-3|LNC|TCRB gene rearrangements|TCRB gene rearrangements
C0804542|T201|COMP|21752-1|LNC|TCRD gene rearrangements|TCRD gene rearrangements
C0804543|T201|COMP|21753-9|LNC|TCRG gene rearrangements|TCRG gene rearrangements
C0804544|T201|COMP|21754-7|LNC|AR gene.CAG repeats|AR gene.CAG repeats
C0804545|T201|COMP|21755-4|LNC|CACNA1A gene.CAG repeats|CACNA1A gene.CAG repeats
C0804546|T201|COMP|21756-2|LNC|ATN1 gene.CAG repeats|ATN1 gene.CAG repeats
C0804547|T201|COMP|21757-0|LNC|DMPK gene.CTG repeats|DMPK gene.CTG repeats
C0804548|T201|COMP|21759-6|LNC|FMR1 gene.CGG repeats|FMR1 gene.CGG repeats
C0804549|T201|COMP|21760-4|LNC|FRAXE gene.CGG repeats|FRAXE gene.CGG repeats
C0804550|T201|COMP|21761-2|LNC|FRAXE gene.CGG repeats|FRAXE gene.CGG repeats
C0804551|T201|COMP|21762-0|LNC|FXN gene.GAA repeats|FXN gene.GAA repeats
C0804552|T201|COMP|21763-8|LNC|HTT gene.CAG repeats|HTT gene.CAG repeats
C0804553|T201|COMP|21764-6|LNC|MJD gene.CAG repeats|MJD gene.CAG repeats
C0804554|T201|COMP|21765-3|LNC|SCA1 gene.CAG repeats|SCA1 gene.CAG repeats
C0804555|T201|COMP|21766-1|LNC|SCA2 gene.CAG repeats|SCA2 gene.CAG repeats
C0804556|T201|COMP|21767-9|LNC|SCA7 gene.CAG repeats|SCA7 gene.CAG repeats
C0804557|T201|COMP|21768-7|LNC|Spinocerebellar ataxia gene mutations tested for|Spinocerebellar ataxia gene mutations tested for
C0804558|T201|COMP|21769-5|LNC|Spinocerebellar ataxia genes.CAG repeats|Spinocerebellar ataxia genes.CAG repeats
C0804559|T201|COMP|21770-3|LNC|Chromosome 12 trisomy|Chromosome 12 trisomy
C0804560|T201|COMP|21771-1|LNC|Chromosome 21 trisomy|Chromosome 21 trisomy
C0804561|T201|COMP|21772-9|LNC|Chromosome 7 trisomy|Chromosome 7 trisomy
C0804562|T201|COMP|21773-7|LNC|Chromosome 8 trisomy|Chromosome 8 trisomy
C0804563|T201|COMP|21774-5|LNC|Chromosome 9 trisomy|Chromosome 9 trisomy
C0804565|T201|COMP|21776-0|LNC|Cells.t(1;19)(q23.3;p13.3)(PBX1,TCF3)/Cells.total|Cells.t(1;19)(q23.3;p13.3)(PBX1,TCF3)/Cells.total
C0804566|T201|COMP|21777-8|LNC|Cells.t(11;14)(q13;q32)(CCND1,IGH)/Cells.total|Cells.t(11;14)(q13;q32)(CCND1,IGH)/Cells.total
C0804567|T201|COMP|21778-6|LNC|Cells.t(11;19)(q23;p13.3)(MLL,MLLT1)/Cells.total|Cells.t(11;19)(q23;p13.3)(MLL,MLLT1)/Cells.total
C0804568|T201|COMP|21779-4|LNC|Cells.t(11;22)(q24;q12.2)(FLI1,EWSR1)/Cells.total|Cells.t(11;22)(q24;q12.2)(FLI1,EWSR1)/Cells.total
C0804569|T201|COMP|21780-2|LNC|Cells.t(11;22)(p13;q12.2)(WT1,EWSR1)/Cells.total|Cells.t(11;22)(p13;q12.2)(WT1,EWSR1)/Cells.total
C0804570|T201|COMP|21781-0|LNC|Cells.t(12;16)(q13;p11.2)(DDIT3,FUS)/Cells.total|Cells.t(12;16)(q13;p11.2)(DDIT3,FUS)/Cells.total
C0804571|T201|COMP|21782-8|LNC|Cells.t(12;21)(p13;q22.3)(ETV6,RUNX1)/Cells.total|Cells.t(12;21)(p13;q22.3)(ETV6,RUNX1)/Cells.total
C0804572|T201|COMP|21783-6|LNC|Cells.t(12;22)(q13;q12.2)(ATF1,EWSR1)/Cells.total|Cells.t(12;22)(q13;q12.2)(ATF1,EWSR1)/Cells.total
C0804573|T201|COMP|21784-4|LNC|Cells.t(14;18)(q32;q21.3)(IGH,BCL2)/Cells.total|Cells.t(14;18)(q32;q21.3)(IGH,BCL2)/Cells.total
C0804574|T201|COMP|21785-1|LNC|Cells.t(15;17)(q24.1;q21.1)(PML,RARA)/Cells.total|Cells.t(15;17)(q24.1;q21.1)(PML,RARA)/Cells.total
C0804576|T201|COMP|21787-7|LNC|Cells.t(2;5)(p23;q35.1)(ALK,NPM1)/Cells.total|Cells.t(2;5)(p23;q35.1)(ALK,NPM1)/Cells.total
C0804578|T201|COMP|21789-3|LNC|Cells.t(4;11)(q21.3;q23)(AFF1,MLL)/Cells.total|Cells.t(4;11)(q21.3;q23)(AFF1,MLL)/Cells.total
C0804579|T201|COMP|21790-1|LNC|Cells.t(5;12)(q33.1;p13)(PDGFRB,ETV6)/Cells.total|Cells.t(5;12)(q33.1;p13)(PDGFRB,ETV6)/Cells.total
C0804580|T201|COMP|21791-9|LNC|Cells.t(6;9)(p22;q34)(DEK,NUP214)/Cells.total|Cells.t(6;9)(p22;q34)(DEK,NUP214)/Cells.total
C0804581|T201|COMP|21792-7|LNC|Cells.t(8;14)(q24;q32)(MYC,IGH)/Cells.total|Cells.t(8;14)(q24;q32)(MYC,IGH)/Cells.total
C0804583|T201|COMP|21794-3|LNC|Cells.t(9;11)(p22;q23)(MLLT3,MLL)/Cells.total|Cells.t(9;11)(p22;q23)(MLLT3,MLL)/Cells.total
C0804584|T201|COMP|21795-0|LNC|Cells.t(9;22)(q34.1;q11)(ABL1,BCR)/Cells.total|Cells.t(9;22)(q34.1;q11)(ABL1,BCR)/Cells.total
C0804585|T201|COMP|21796-8|LNC|Cells.t(9;22)(q22;q12.2)(NR4A3,EWSR1)/Cells.total|Cells.t(9;22)(q22;q12.2)(NR4A3,EWSR1)/Cells.total
C0804589|T201|COMP|21800-8|LNC|t(1;19)(q23.3;p13.3)(PBX1,TCF3) fusion transcript|t(1;19)(q23.3;p13.3)(PBX1,TCF3) fusion transcript
C0804590|T201|COMP|21801-6|LNC|t(11;14)(q13;q32)(CCND1,IGH) fusion transcript|t(11;14)(q13;q32)(CCND1,IGH) fusion transcript
C0804591|T201|COMP|21802-4|LNC|t(11;19)(q23;p13.3)(MLL,MLLT1) fusion transcript|t(11;19)(q23;p13.3)(MLL,MLLT1) fusion transcript
C0804592|T201|COMP|21803-2|LNC|t(11;22)(q24;q12.2)(FLI1,EWSR1) fusion transcript|t(11;22)(q24;q12.2)(FLI1,EWSR1) fusion transcript
C0804593|T201|COMP|21804-0|LNC|t(11;22)(p13;q12.2)(WT1,EWSR1) fusion transcript|t(11;22)(p13;q12.2)(WT1,EWSR1) fusion transcript
C0804594|T201|COMP|21805-7|LNC|t(12;16)(q13;p11.2)(DDIT3,FUS) fusion transcript|t(12;16)(q13;p11.2)(DDIT3,FUS) fusion transcript
C0804595|T201|COMP|21806-5|LNC|t(12;21)(p13;q22.3)(ETV6,RUNX1) fusion transcript|t(12;21)(p13;q22.3)(ETV6,RUNX1) fusion transcript
C0804596|T201|COMP|21807-3|LNC|t(12;22)(q13;q12.2)(ATF1,EWSR1) fusion transcript|t(12;22)(q13;q12.2)(ATF1,EWSR1) fusion transcript
C0804597|T201|COMP|21808-1|LNC|t(14;18)(q32;q21.3)(IGH,BCL2) fusion transcript|t(14;18)(q32;q21.3)(IGH,BCL2) fusion transcript
C0804601|T201|COMP|21813-1|LNC|t(2;5)(p23;q35.1)(ALK,NPM1) fusion transcript|t(2;5)(p23;q35.1)(ALK,NPM1) fusion transcript
C0804603|T201|COMP|21815-6|LNC|t(4;11)(q21.3;q23)(AFF1,MLL) fusion transcript|t(4;11)(q21.3;q23)(AFF1,MLL) fusion transcript
C0804604|T201|COMP|21816-4|LNC|t(5;12)(q33.1;p13)(PDGFRB,ETV6) fusion transcript|t(5;12)(q33.1;p13)(PDGFRB,ETV6) fusion transcript
C0804605|T201|COMP|21817-2|LNC|t(6;9)(p22;q34)(DEK,NUP214) fusion transcript|t(6;9)(p22;q34)(DEK,NUP214) fusion transcript
C0804606|T201|COMP|21818-0|LNC|t(8;14)(q24;q32)(MYC,IGH) fusion transcript|t(8;14)(q24;q32)(MYC,IGH) fusion transcript
C0804608|T201|COMP|21820-6|LNC|t(9;11)(p22;q23)(MLLT3,MLL) fusion transcript|t(9;11)(p22;q23)(MLLT3,MLL) fusion transcript
C0804609|T201|COMP|21821-4|LNC|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript
C0804612|T201|COMP|21824-8|LNC|t(9;22)(q22;q12.2)(NR4A3,EWSR1) fusion transcript|t(9;22)(q22;q12.2)(NR4A3,EWSR1) fusion transcript
C0804851|T201|COMP|22064-0|LNC|Alpha 1 globulin|Alpha 1 globulin
C0804853|T201|COMP|22066-5|LNC|PRSS1 gene mutations tested for|PRSS1 gene mutations tested for
C0804854|T201|COMP|22067-3|LNC|NB gene mutations tested for|NB gene mutations tested for
C0804855|T201|COMP|22068-1|LNC|MXI1 gene mutations tested for|MXI1 gene mutations tested for
C0804856|T201|COMP|22069-9|LNC|MT-ATP6 gene mutations tested for|MT-ATP6 gene mutations tested for
C0804861|T201|COMP|22074-9|LNC|FGFR3 gene mutations tested for|FGFR3 gene mutations tested for
C0804862|T201|COMP|22075-6|LNC|DMD gene mutations tested for|DMD gene mutations tested for
C0804863|T201|COMP|22076-4|LNC|CMKBR5 gene mutations tested for|CMKBR5 gene mutations tested for
C0804864|T201|COMP|66-1|LNC|Cefadroxil|Cefadroxil
C0812452|T201|COMP|19238-5|LNC|Base excess^^standard|Base excess^^standard
C0812457|T201|COMP|19235-1|LNC|Base excess^^standard|Base excess^^standard
C0812458|T201|COMP|19236-9|LNC|Base excess^^standard|Base excess^^standard
C0812459|T201|COMP|19237-7|LNC|Base excess^^standard|Base excess^^standard
C0812460|T201|COMP|19230-2|LNC|Bicarbonate^^standard|Bicarbonate^^standard
C0812461|T201|COMP|19231-0|LNC|Bicarbonate^^standard|Bicarbonate^^standard
C0812462|T201|COMP|19072-8|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C0812463|T201|COMP|5917-0|LNC|???lead|???lead
C0877808|T201|COMP|1005-8|LNC|Indirect antiglobulin test.IgG specific reagent|Indirect antiglobulin test.IgG specific reagent
C0877809|T201|COMP|1008-2|LNC|Indirect antiglobulin test.poly specific reagent|Indirect antiglobulin test.poly specific reagent
C0877892|T201|COMP|16827-8|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0879639|T201|COMP|19044-7|LNC|Artemia salina Ab.IgE.RAST class|Artemia salina Ab.IgE.RAST class
C0879640|T201|COMP|19045-4|LNC|Salmo salar Ab.IgG.RAST class|Salmo salar Ab.IgG.RAST class
C0879641|T201|COMP|19047-0|LNC|Thunnus albacares Ab.IgG.RAST class|Thunnus albacares Ab.IgG.RAST class
C0879643|T201|COMP|19051-2|LNC|Saquinavir|Saquinavir
C0879644|T201|COMP|19052-0|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C0879645|T201|COMP|19053-8|LNC|Brucella sp Ab|Brucella sp Ab
C0879646|T201|COMP|19054-6|LNC|Mycoplasma pneumoniae|Mycoplasma pneumoniae
C0879647|T201|COMP|19055-3|LNC|Carboxy tetrahydrocannabinol/Creatinine|Carboxy tetrahydrocannabinol/Creatinine
C0879648|T201|COMP|19056-1|LNC|Mercury|Mercury
C0879649|T201|COMP|19724-4|LNC|Triplochiton scleroxylon Ab.IgE|Triplochiton scleroxylon Ab.IgE
C0879650|T201|COMP|19726-9|LNC|Aspergillus fumigatus Ab.IgG|Aspergillus fumigatus Ab.IgG
C0879651|T201|COMP|19727-7|LNC|Aspergillus niger Ab.IgG|Aspergillus niger Ab.IgG
C0879652|T201|COMP|19728-5|LNC|Beet Ab.IgE|Beet Ab.IgE
C0879653|T201|COMP|19729-3|LNC|Lathyrus sativus Ab.IgE|Lathyrus sativus Ab.IgE
C0879654|T201|COMP|19730-1|LNC|Budgerigar droppings Ab.IgE|Budgerigar droppings Ab.IgE
C0879655|T201|COMP|19731-9|LNC|Budgerigar serum proteins Ab.IgE|Budgerigar serum proteins Ab.IgE
C0879656|T201|COMP|19732-7|LNC|Cat serum albumin Ab.IgE|Cat serum albumin Ab.IgE
C0879657|T201|COMP|19734-3|LNC|Chicken droppings Ab.IgE|Chicken droppings Ab.IgE
C0879659|T201|COMP|19736-8|LNC|Coralbumin Ab.IgE|Coralbumin Ab.IgE
C0879660|T201|COMP|19737-6|LNC|Cotton fibers Ab.IgE|Cotton fibers Ab.IgE
C0879661|T201|COMP|19739-2|LNC|Trigonella foenum-graecum Ab.IgE|Trigonella foenum-graecum Ab.IgE
C0879662|T201|COMP|19740-0|LNC|Fox epithelium Ab.IgE|Fox epithelium Ab.IgE
C0879663|T201|COMP|19741-8|LNC|Merluccius merluccius Ab.IgE|Merluccius merluccius Ab.IgE
C0879664|T201|COMP|19743-4|LNC|Horse meat Ab.IgE|Horse meat Ab.IgE
C0879665|T201|COMP|19744-2|LNC|Artocarpus heterophyllus Ab.IgE|Artocarpus heterophyllus Ab.IgE
C0879667|T201|COMP|19746-7|LNC|Maleic anhydride Ab.IgE|Maleic anhydride Ab.IgE
C0879668|T201|COMP|19747-5|LNC|Tenebrio mollitor Ab.IgE|Tenebrio mollitor Ab.IgE
C0879669|T201|COMP|19748-3|LNC|Methyltetrahydrophthalic anhydride Ab.IgE|Methyltetrahydrophthalic anhydride Ab.IgE
C0879670|T201|COMP|19749-1|LNC|Saccharopolyspora rectivirgula Ab.IgG|Saccharopolyspora rectivirgula Ab.IgG
C0879671|T201|COMP|19750-9|LNC|Mentha piperita Ab.IgE|Mentha piperita Ab.IgE
C0879673|T201|COMP|19752-5|LNC|Pigeon serum Ab.IgG|Pigeon serum Ab.IgG
C0879675|T201|COMP|19754-1|LNC|Ribes sylvestre Ab.IgE|Ribes sylvestre Ab.IgE
C0879676|T201|COMP|19755-8|LNC|Crocus sativus Ab.IgE|Crocus sativus Ab.IgE
C0879677|T201|COMP|19756-6|LNC|Sheep milk Ab.IgE|Sheep milk Ab.IgE
C0879678|T201|COMP|19757-4|LNC|Sheep whey Ab.IgE|Sheep whey Ab.IgE
C0879679|T201|COMP|19758-2|LNC|Silk waste Ab.IgE|Silk waste Ab.IgE
C0879680|T201|COMP|19759-0|LNC|Swine serum albumin Ab.IgE|Swine serum albumin Ab.IgE
C0879681|T201|COMP|19760-8|LNC|Clostridium tetani toxoid Ab.IgE|Clostridium tetani toxoid Ab.IgE
C0879682|T201|COMP|19761-6|LNC|Thermoactinomyces vulgaris Ab.IgG|Thermoactinomyces vulgaris Ab.IgG
C0879683|T201|COMP|22077-2|LNC|Acanthamoeba sp Ab|Acanthamoeba sp Ab
C0879684|T201|COMP|22078-0|LNC|Acanthamoeba sp Ab|Acanthamoeba sp Ab
C0879685|T201|COMP|22080-6|LNC|Adenovirus Ab|Adenovirus Ab
C0879686|T201|COMP|22081-4|LNC|Afipia felis Ab.IgG|Afipia felis Ab.IgG
C0879687|T201|COMP|22082-2|LNC|Afipia felis Ab.IgM|Afipia felis Ab.IgM
C0879688|T201|COMP|22084-8|LNC|Anaplasma marginale Ab|Anaplasma marginale Ab
C0879689|T201|COMP|22085-5|LNC|Aspergillus fumigatus 3 Ab|Aspergillus fumigatus 3 Ab
C0879690|T201|COMP|22086-3|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C0879691|T201|COMP|22087-1|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C0879692|T201|COMP|22089-7|LNC|Avian adenovirus Ab|Avian adenovirus Ab
C0879693|T201|COMP|22091-3|LNC|Avian hemorrhagic enteritis virus Ab|Avian hemorrhagic enteritis virus Ab
C0879694|T201|COMP|22093-9|LNC|Infectious bronchitis virus Conn-42 Ab|Infectious bronchitis virus Conn-42 Ab
C0879695|T201|COMP|22094-7|LNC|Infectious bronchitis virus Mass-41 Ab|Infectious bronchitis virus Mass-41 Ab
C0879696|T201|COMP|22096-2|LNC|Influenza virus A Ab|Influenza virus A Ab
C0879697|T201|COMP|22097-0|LNC|Avian paramyxovirus 1 Ab|Avian paramyxovirus 1 Ab
C0879698|T201|COMP|22098-8|LNC|Avian paramyxovirus 1 Ab|Avian paramyxovirus 1 Ab
C0879699|T201|COMP|22099-6|LNC|Avian paramyxovirus 2 Ab|Avian paramyxovirus 2 Ab
C0879700|T201|COMP|22100-2|LNC|Avian paramyxovirus 3 Ab|Avian paramyxovirus 3 Ab
C0879701|T201|COMP|22101-0|LNC|Avian pox virus Ab|Avian pox virus Ab
C0879702|T201|COMP|22102-8|LNC|Avian reovirus Ab|Avian reovirus Ab
C0879703|T201|COMP|22103-6|LNC|Reticuloendotheliosis virus Ab|Reticuloendotheliosis virus Ab
C0879704|T201|COMP|22105-1|LNC|Theileria equi Ab|Theileria equi Ab
C0879705|T201|COMP|22106-9|LNC|Babesia sp Ab|Babesia sp Ab
C0879706|T201|COMP|22107-7|LNC|Babesia sp Ab.IgG|Babesia sp Ab.IgG
C0879707|T201|COMP|22108-5|LNC|Babesia sp Ab.IgM|Babesia sp Ab.IgM
C0879708|T201|COMP|22109-3|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0879709|T201|COMP|22110-1|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C0879710|T201|COMP|22111-9|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C0879711|T201|COMP|22112-7|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0879712|T201|COMP|22113-5|LNC|Bluetongue virus Ab|Bluetongue virus Ab
C0879713|T201|COMP|22114-3|LNC|Bordetella avium Ab|Bordetella avium Ab
C0879714|T201|COMP|22115-0|LNC|Bordetella avium Ab|Bordetella avium Ab
C0879715|T201|COMP|22116-8|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C0879716|T201|COMP|22117-6|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C0879717|T201|COMP|22118-4|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0879718|T201|COMP|22119-2|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0879719|T201|COMP|22120-0|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0879720|T201|COMP|22121-8|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0879721|T201|COMP|22122-6|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0879722|T201|COMP|22123-4|LNC|Borrelia burgdorferi Ab.IgA|Borrelia burgdorferi Ab.IgA
C0879723|T201|COMP|22124-2|LNC|Borrelia burgdorferi Ab.IgA|Borrelia burgdorferi Ab.IgA
C0879724|T201|COMP|22126-7|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0879725|T201|COMP|22127-5|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0879726|T201|COMP|22129-1|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0879727|T201|COMP|22130-9|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0879728|T201|COMP|22131-7|LNC|Borrelia burgdorferi Ab.IgG+IgM|Borrelia burgdorferi Ab.IgG+IgM
C0879729|T201|COMP|22132-5|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0879730|T201|COMP|22134-1|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0879731|T201|COMP|22135-8|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0879732|T201|COMP|22136-6|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0879733|T201|COMP|22137-4|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0879734|T201|COMP|22139-0|LNC|Borrelia hermsii Ab.IgM|Borrelia hermsii Ab.IgM
C0879735|T201|COMP|22140-8|LNC|Bovine diarrhea virus 1 Ab|Bovine diarrhea virus 1 Ab
C0879736|T201|COMP|22141-6|LNC|Bovine diarrhea virus 2 Ab|Bovine diarrhea virus 2 Ab
C0879737|T201|COMP|22143-2|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C0879738|T201|COMP|22144-0|LNC|Bovine leukemia virus Ab|Bovine leukemia virus Ab
C0879739|T201|COMP|22145-7|LNC|Bovine leukosis virus Ab|Bovine leukosis virus Ab
C0879740|T201|COMP|22146-5|LNC|Brucella abortus Ab|Brucella abortus Ab
C0879741|T201|COMP|22148-1|LNC|Brucella abortus Ab|Brucella abortus Ab
C0879742|T201|COMP|22149-9|LNC|Brucella abortus Ab|Brucella abortus Ab
C0879743|T201|COMP|22150-7|LNC|Brucella abortus Ab|Brucella abortus Ab
C0879744|T201|COMP|22152-3|LNC|Brucella canis Ab|Brucella canis Ab
C0879745|T201|COMP|22153-1|LNC|Brucella canis Ab.IgG|Brucella canis Ab.IgG
C0879746|T201|COMP|22154-9|LNC|Brucella canis Ab.IgG|Brucella canis Ab.IgG
C0879747|T201|COMP|22155-6|LNC|Brucella canis Ab.IgM|Brucella canis Ab.IgM
C0879748|T201|COMP|22156-4|LNC|Brucella canis Ab.IgM|Brucella canis Ab.IgM
C0879749|T201|COMP|22157-2|LNC|Brucella melitensis Ab|Brucella melitensis Ab
C0879750|T201|COMP|22158-0|LNC|Brucella ovis Ab|Brucella ovis Ab
C0879751|T201|COMP|22159-8|LNC|Brucella sp Ab|Brucella sp Ab
C0879752|T201|COMP|22160-6|LNC|Brucella suis Ab|Brucella suis Ab
C0879753|T201|COMP|22161-4|LNC|Cache valley virus Ab|Cache valley virus Ab
C0879754|T201|COMP|22162-2|LNC|Candida albicans Ab|Candida albicans Ab
C0879755|T201|COMP|22163-0|LNC|Candida albicans Ab|Candida albicans Ab
C0879756|T201|COMP|22164-8|LNC|Caprine arthritis encephalitis virus Ab|Caprine arthritis encephalitis virus Ab
C0879757|T201|COMP|22166-3|LNC|Caprine parapoxvirus Ab|Caprine parapoxvirus Ab
C0879758|T201|COMP|22167-1|LNC|Caprine parapoxvirus Ab|Caprine parapoxvirus Ab
C0879759|T201|COMP|22168-9|LNC|Chicken anemia virus Ab|Chicken anemia virus Ab
C0879760|T201|COMP|22169-7|LNC|Chlamydophila pneumoniae Ab.IgA|Chlamydophila pneumoniae Ab.IgA
C0879761|T201|COMP|22170-5|LNC|Chlamydophila pneumoniae Ab.IgA|Chlamydophila pneumoniae Ab.IgA
C0879762|T201|COMP|22171-3|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C0879763|T201|COMP|22172-1|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C0879764|T201|COMP|22173-9|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C0879765|T201|COMP|22174-7|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C0879766|T201|COMP|22175-4|LNC|Chlamydophila psittaci Ab|Chlamydophila psittaci Ab
C0879767|T201|COMP|22176-2|LNC|Chlamydophila psittaci Ab|Chlamydophila psittaci Ab
C0879768|T201|COMP|22177-0|LNC|Chlamydophila psittaci Ab.IgA|Chlamydophila psittaci Ab.IgA
C0879769|T201|COMP|22178-8|LNC|Chlamydophila psittaci Ab.IgA|Chlamydophila psittaci Ab.IgA
C0879770|T201|COMP|22180-4|LNC|Chlamydophila psittaci Ab.IgG|Chlamydophila psittaci Ab.IgG
C0879771|T201|COMP|22181-2|LNC|Chlamydophila psittaci Ab.IgM|Chlamydophila psittaci Ab.IgM
C0879772|T201|COMP|22182-0|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0879773|T201|COMP|22183-8|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C0879774|T201|COMP|22184-6|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C0879775|T201|COMP|22185-3|LNC|Chlamydia sp Ab.IgM|Chlamydia sp Ab.IgM
C0879776|T201|COMP|22186-1|LNC|Chlamydia sp Ab.IgM|Chlamydia sp Ab.IgM
C0879777|T201|COMP|22188-7|LNC|Chlamydia trachomatis Ab.IgA|Chlamydia trachomatis Ab.IgA
C0879778|T201|COMP|22189-5|LNC|Chlamydia trachomatis Ab.IgA|Chlamydia trachomatis Ab.IgA
C0879779|T201|COMP|22190-3|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C0879780|T201|COMP|22192-9|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C0879781|T201|COMP|22193-7|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C0879782|T201|COMP|22194-5|LNC|Chlamydia trachomatis B Ab.IgA|Chlamydia trachomatis B Ab.IgA
C0879783|T201|COMP|22195-2|LNC|Chlamydia trachomatis B Ab.IgG|Chlamydia trachomatis B Ab.IgG
C0879784|T201|COMP|22197-8|LNC|Chlamydia trachomatis C Ab.IgA|Chlamydia trachomatis C Ab.IgA
C0879785|T201|COMP|22198-6|LNC|Chlamydia trachomatis C Ab.IgG|Chlamydia trachomatis C Ab.IgG
C0879786|T201|COMP|22199-4|LNC|Chlamydia trachomatis C Ab.IgM|Chlamydia trachomatis C Ab.IgM
C0879787|T201|COMP|22200-0|LNC|Chlamydia trachomatis G+F+K Ab.IgA|Chlamydia trachomatis G+F+K Ab.IgA
C0879788|T201|COMP|22201-8|LNC|Chlamydia trachomatis G+F+K Ab.IgG|Chlamydia trachomatis G+F+K Ab.IgG
C0879789|T201|COMP|22202-6|LNC|Chlamydia trachomatis G+F+K Ab.IgM|Chlamydia trachomatis G+F+K Ab.IgM
C0879790|T201|COMP|22204-2|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0879791|T201|COMP|22205-9|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0879792|T201|COMP|22206-7|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0879793|T201|COMP|22207-5|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0879794|T201|COMP|22209-1|LNC|Coccidioides immitis Ab.IgG|Coccidioides immitis Ab.IgG
C0879795|T201|COMP|22210-9|LNC|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C0879796|T201|COMP|22213-3|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C0879797|T201|COMP|22214-1|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C0879798|T201|COMP|22215-8|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C0879799|T201|COMP|22216-6|LNC|Coxsackievirus A2 Ab|Coxsackievirus A2 Ab
C0879800|T201|COMP|22218-2|LNC|Coxsackievirus A4 Ab|Coxsackievirus A4 Ab
C0879801|T201|COMP|22219-0|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C0879802|T201|COMP|22220-8|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C0879803|T201|COMP|22221-6|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C0879804|T201|COMP|22222-4|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C0879805|T201|COMP|22223-2|LNC|Coxsackievirus B Ab.IgG|Coxsackievirus B Ab.IgG
C0879806|T201|COMP|22224-0|LNC|Coxsackievirus B Ab.IgM|Coxsackievirus B Ab.IgM
C0879807|T201|COMP|22225-7|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C0879808|T201|COMP|22226-5|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C0879809|T201|COMP|22227-3|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C0879810|T201|COMP|22228-1|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C0879811|T201|COMP|22229-9|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C0879812|T201|COMP|22230-7|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C0879813|T201|COMP|22231-5|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C0879814|T201|COMP|22232-3|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C0879815|T201|COMP|22233-1|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C0879816|T201|COMP|22234-9|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C0879817|T201|COMP|22235-6|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C0879818|T201|COMP|22236-4|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C0879819|T201|COMP|22238-0|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C0879820|T201|COMP|22239-8|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0879821|T201|COMP|22240-6|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0879823|T201|COMP|22241-4|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C0879824|T201|COMP|22243-0|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0879825|T201|COMP|22244-8|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0879826|T201|COMP|22245-5|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0879827|T201|COMP|22246-3|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0879828|T201|COMP|22247-1|LNC|Cytomegalovirus Ab.IgG^2nd specimen|Cytomegalovirus Ab.IgG^2nd specimen
C0879829|T201|COMP|22248-9|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0879830|T201|COMP|22249-7|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0879831|T201|COMP|22251-3|LNC|Dengue virus 2 Ab|Dengue virus 2 Ab
C0879832|T201|COMP|22252-1|LNC|Dengue virus 3 Ab|Dengue virus 3 Ab
C0879833|T201|COMP|22253-9|LNC|Dengue virus 4 Ab|Dengue virus 4 Ab
C0879834|T201|COMP|22254-7|LNC|Duck enteritis virus Ab|Duck enteritis virus Ab
C0879835|T201|COMP|22256-2|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0879837|T201|COMP|22258-8|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C0879838|T201|COMP|22259-6|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C0879839|T201|COMP|22260-4|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C0879840|T201|COMP|22261-2|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C0879841|T201|COMP|22257-0|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0879842|T201|COMP|22263-8|LNC|Ebola virus Ab|Ebola virus Ab
C0879843|T201|COMP|22265-3|LNC|Echinococcus sp Ab.IgG|Echinococcus sp Ab.IgG
C0879844|T201|COMP|22266-1|LNC|Echovirus 1 Ab|Echovirus 1 Ab
C0879845|T201|COMP|22267-9|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C0879846|T201|COMP|22268-7|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C0879847|T201|COMP|22270-3|LNC|Echovirus 140 Ab|Echovirus 140 Ab
C0879848|T201|COMP|22271-1|LNC|Echovirus 16 Ab|Echovirus 16 Ab
C0879849|T201|COMP|22272-9|LNC|Echovirus 18 Ab|Echovirus 18 Ab
C0879850|T201|COMP|22274-5|LNC|Echovirus 3 Ab|Echovirus 3 Ab
C0879851|T201|COMP|22275-2|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C0879852|T201|COMP|22276-0|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C0879853|T201|COMP|22278-6|LNC|Echovirus 6 Ab|Echovirus 6 Ab
C0879854|T201|COMP|22279-4|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C0879855|T201|COMP|22280-2|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C0879856|T201|COMP|22282-8|LNC|Echovirus NOS Ab|Echovirus NOS Ab
C0879857|T201|COMP|22283-6|LNC|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C0879858|T201|COMP|22284-4|LNC|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C0879859|T201|COMP|22285-1|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0879860|T201|COMP|22286-9|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0879861|T201|COMP|22287-7|LNC|Entamoeba histolytica Ab.IgA|Entamoeba histolytica Ab.IgA
C0879862|T201|COMP|22288-5|LNC|Entamoeba histolytica Ab.IgG|Entamoeba histolytica Ab.IgG
C0879863|T201|COMP|22289-3|LNC|Entamoeba histolytica Ab.IgM|Entamoeba histolytica Ab.IgM
C0879864|T201|COMP|22290-1|LNC|Epstein Barr virus capsid Ab.IgA|Epstein Barr virus capsid Ab.IgA
C0879865|T201|COMP|22291-9|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0879866|T201|COMP|22292-7|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0879867|T201|COMP|22294-3|LNC|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C0879868|T201|COMP|22295-0|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C0879869|T201|COMP|22296-8|LNC|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C0879870|T201|COMP|22297-6|LNC|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C0879871|T201|COMP|22298-4|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0879872|T201|COMP|22299-2|LNC|Equine arteritis virus Ab|Equine arteritis virus Ab
C0879873|T201|COMP|22300-8|LNC|Equine herpesvirus 1 Ab|Equine herpesvirus 1 Ab
C0879874|T201|COMP|22301-6|LNC|Equine infectious anemia virus Ab|Equine infectious anemia virus Ab
C0879875|T201|COMP|22302-4|LNC|Equine influenza virus A1 Ab|Equine influenza virus A1 Ab
C0879876|T201|COMP|22303-2|LNC|Equine influenza virus A2 Ab|Equine influenza virus A2 Ab
C0879877|T201|COMP|22304-0|LNC|Giardia lamblia Ab|Giardia lamblia Ab
C0879878|T201|COMP|22305-7|LNC|Giardia lamblia Ab.IgA|Giardia lamblia Ab.IgA
C0879879|T201|COMP|22306-5|LNC|Giardia lamblia Ab.IgG|Giardia lamblia Ab.IgG
C0879880|T201|COMP|22307-3|LNC|Giardia lamblia Ab.IgM|Giardia lamblia Ab.IgM
C0879881|T201|COMP|22308-1|LNC|Hantavirus puumala Ab.IgG|Hantavirus puumala Ab.IgG
C0879882|T201|COMP|22309-9|LNC|Hantavirus puumala Ab.IgM|Hantavirus puumala Ab.IgM
C0879883|T201|COMP|22310-7|LNC|Helicobacter pylori Ab|Helicobacter pylori Ab
C0879884|T201|COMP|22313-1|LNC|Hepatitis A virus Ab.IgG|Hepatitis A virus Ab.IgG
C0879885|T201|COMP|22314-9|LNC|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C0879886|T201|COMP|22315-6|LNC|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C0879887|T201|COMP|22316-4|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C0879888|T201|COMP|22318-0|LNC|Hepatitis B virus core Ab.IgG|Hepatitis B virus core Ab.IgG
C0879889|T201|COMP|22319-8|LNC|Hepatitis B virus core Ab.IgM|Hepatitis B virus core Ab.IgM
C0879890|T201|COMP|22320-6|LNC|Hepatitis B virus little e Ab|Hepatitis B virus little e Ab
C0879891|T201|COMP|22322-2|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0879892|T201|COMP|22323-0|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0879893|T201|COMP|22325-5|LNC|Hepatitis C virus 22-3 Ab|Hepatitis C virus 22-3 Ab
C0879894|T201|COMP|22327-1|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C0879895|T201|COMP|22328-9|LNC|Hepatitis C virus superoxide dismutase Ab|Hepatitis C virus superoxide dismutase Ab
C0879896|T201|COMP|22329-7|LNC|Hepatitis C virus c33c Ab|Hepatitis C virus c33c Ab
C0879897|T201|COMP|22330-5|LNC|Hepatitis D virus Ab|Hepatitis D virus Ab
C0879898|T201|COMP|22332-1|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C0879899|T201|COMP|22333-9|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C0879900|T201|COMP|22334-7|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C0879901|T201|COMP|22335-4|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C0879902|T201|COMP|22337-0|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0879903|T201|COMP|22338-8|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C0879904|T201|COMP|22339-6|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C0879905|T201|COMP|22341-2|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C0879906|T201|COMP|22342-0|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C0879907|T201|COMP|22343-8|LNC|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C0879908|T201|COMP|22344-6|LNC|Heterophile Ab after absorption|Heterophile Ab after absorption
C0879909|T201|COMP|22345-3|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0879910|T201|COMP|22346-1|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0879911|T201|COMP|22347-9|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0879912|T201|COMP|22348-7|LNC|Histoplasma capsulatum Ab.IgA|Histoplasma capsulatum Ab.IgA
C0879913|T201|COMP|22350-3|LNC|Histoplasma capsulatum Ab.IgE|Histoplasma capsulatum Ab.IgE
C0879914|T201|COMP|22351-1|LNC|Histoplasma capsulatum Ab.IgG|Histoplasma capsulatum Ab.IgG
C0879915|T201|COMP|22352-9|LNC|Histoplasma capsulatum Ab.IgM|Histoplasma capsulatum Ab.IgM
C0879916|T201|COMP|22353-7|LNC|Histoplasma capsulatum Ab.IgM|Histoplasma capsulatum Ab.IgM
C0879917|T201|COMP|22354-5|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C0879918|T201|COMP|22355-2|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C0879919|T201|COMP|22356-0|LNC|HIV 1 Ab|HIV 1 Ab
C0879920|T201|COMP|22357-8|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C0879921|T201|COMP|22358-6|LNC|HIV 2 Ab|HIV 2 Ab
C0879922|T201|COMP|22359-4|LNC|HTLV I Ab|HTLV I Ab
C0879923|T201|COMP|22360-2|LNC|HTLV I Ab.IgG|HTLV I Ab.IgG
C0879924|T201|COMP|22361-0|LNC|HTLV I+II Ab|HTLV I+II Ab
C0879925|T201|COMP|22362-8|LNC|HTLV I+II Ab|HTLV I+II Ab
C0879926|T201|COMP|22363-6|LNC|HTLV I+II Ab|HTLV I+II Ab
C0879927|T201|COMP|22364-4|LNC|Infectious bursal disease virus Ab|Infectious bursal disease virus Ab
C0879928|T201|COMP|22365-1|LNC|Influenza virus A Ab|Influenza virus A Ab
C0879929|T201|COMP|22366-9|LNC|Influenza virus A+B Ab|Influenza virus A+B Ab
C0879930|T201|COMP|22367-7|LNC|Influenza virus B Ab|Influenza virus B Ab
C0879931|T201|COMP|22368-5|LNC|Influenza virus C Ab|Influenza virus C Ab
C0879932|T201|COMP|22369-3|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0879933|T201|COMP|22370-1|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0879934|T201|COMP|22371-9|LNC|Junin virus Ab|Junin virus Ab
C0879935|T201|COMP|22372-7|LNC|La Crosse virus Ab|La Crosse virus Ab
C0879936|T201|COMP|22373-5|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C0879937|T201|COMP|22375-0|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C0879938|T201|COMP|17039-9|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C0879939|T201|COMP|22377-6|LNC|Lassa virus Ab.IgG|Lassa virus Ab.IgG
C0879940|T201|COMP|22379-2|LNC|Lassa virus Ab.IgM|Lassa virus Ab.IgM
C0879941|T201|COMP|22380-0|LNC|Lassa virus Ab.IgM|Lassa virus Ab.IgM
C0879942|T201|COMP|22381-8|LNC|Legionella pneumophila 1 Ab.IgG|Legionella pneumophila 1 Ab.IgG
C0879943|T201|COMP|22383-4|LNC|Legionella pneumophila 2 Ab.IgG|Legionella pneumophila 2 Ab.IgG
C0879944|T201|COMP|22384-2|LNC|Legionella pneumophila 2 Ab.IgM|Legionella pneumophila 2 Ab.IgM
C0879945|T201|COMP|22385-9|LNC|Legionella pneumophila 3 Ab.IgG|Legionella pneumophila 3 Ab.IgG
C0879946|T201|COMP|22386-7|LNC|Legionella pneumophila 3 Ab.IgM|Legionella pneumophila 3 Ab.IgM
C0879947|T201|COMP|22388-3|LNC|Legionella pneumophila 4 Ab.IgM|Legionella pneumophila 4 Ab.IgM
C0879948|T201|COMP|22389-1|LNC|Legionella pneumophila 5 Ab.IgG|Legionella pneumophila 5 Ab.IgG
C0879949|T201|COMP|22390-9|LNC|Legionella pneumophila 5 Ab.IgM|Legionella pneumophila 5 Ab.IgM
C0879950|T201|COMP|22391-7|LNC|Legionella pneumophila 6 Ab.IgG|Legionella pneumophila 6 Ab.IgG
C0879951|T201|COMP|22393-3|LNC|Legionella pneumophila 7 Ab|Legionella pneumophila 7 Ab
C0879952|T201|COMP|22394-1|LNC|Legionella pneumophila 8 Ab|Legionella pneumophila 8 Ab
C0879953|T201|COMP|22395-8|LNC|Legionella pneumophila 9 Ab|Legionella pneumophila 9 Ab
C0879954|T201|COMP|22396-6|LNC|Legionella pneumophila Ab|Legionella pneumophila Ab
C0879955|T201|COMP|22398-2|LNC|Legionella pneumophila Ab.IgM|Legionella pneumophila Ab.IgM
C0879956|T201|COMP|22399-0|LNC|Legionella sp Ab|Legionella sp Ab
C0879957|T201|COMP|22401-4|LNC|Leptospira interrogans serovar Canicola Ab|Leptospira interrogans serovar Canicola Ab
C0879958|T201|COMP|22402-2|LNC|Leptospira interrogans serovar Grippotyphosa Ab|Leptospira interrogans serovar Grippotyphosa Ab
C0879959|T201|COMP|22403-0|LNC|Leptospira interrogans serovar Hardjo Ab|Leptospira interrogans serovar Hardjo Ab
C0879961|T201|COMP|22405-5|LNC|Leptospira interrogans serovar Pomona Ab|Leptospira interrogans serovar Pomona Ab
C0879962|T201|COMP|22406-3|LNC|Listeria monocytogenes Ab|Listeria monocytogenes Ab
C0879963|T201|COMP|22407-1|LNC|little d little s DNA (Crithidia lucilia) Ab|little d little s DNA (Crithidia lucilia) Ab
C0879964|T201|COMP|22408-9|LNC|Lymphocytic choriomeningitis virus Ab|Lymphocytic choriomeningitis virus Ab
C0879965|T201|COMP|22410-5|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C0879966|T201|COMP|22411-3|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C0879967|T201|COMP|22412-1|LNC|Saccharopolyspora rectivirgula Ab|Saccharopolyspora rectivirgula Ab
C0879968|T201|COMP|22413-9|LNC|Mumps virus Ab|Mumps virus Ab
C0879969|T201|COMP|22414-7|LNC|Mumps virus Ab|Mumps virus Ab
C0879970|T201|COMP|22415-4|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0879971|T201|COMP|22416-2|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0879972|T201|COMP|22417-0|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0879973|T201|COMP|22418-8|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C0879974|T201|COMP|22419-6|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C0879975|T201|COMP|22420-4|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C0879977|T201|COMP|22422-0|LNC|Mycoplasma gallisepticum Ab|Mycoplasma gallisepticum Ab
C0879978|T201|COMP|22423-8|LNC|Mycoplasma hominis Ab|Mycoplasma hominis Ab
C0879979|T201|COMP|22424-6|LNC|Mycoplasma meleagridis Ab|Mycoplasma meleagridis Ab
C0879980|T201|COMP|22425-3|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C0879981|T201|COMP|22426-1|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C0879982|T201|COMP|22427-9|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C0879983|T201|COMP|22428-7|LNC|Mycoplasma sp Ab|Mycoplasma sp Ab
C0879984|T201|COMP|22429-5|LNC|Mycoplasma synoviae Ab|Mycoplasma synoviae Ab
C0879985|T201|COMP|22430-3|LNC|Neisseria gonorrhoeae Ab|Neisseria gonorrhoeae Ab
C0879986|T201|COMP|22431-1|LNC|Neisseria meningitidis serogroup Y Ab|Neisseria meningitidis serogroup Y Ab
C0879987|T201|COMP|22432-9|LNC|Neospora caninum Ab|Neospora caninum Ab
C0879988|T201|COMP|22434-5|LNC|Human papilloma virus Ab|Human papilloma virus Ab
C0879989|T201|COMP|22435-2|LNC|Paracoccidioides brasiliensis Ab|Paracoccidioides brasiliensis Ab
C0879990|T201|COMP|22436-0|LNC|Paragonimus sp Ab|Paragonimus sp Ab
C0879991|T201|COMP|22438-6|LNC|Parainfluenza virus 2 Ab|Parainfluenza virus 2 Ab
C0879992|T201|COMP|22439-4|LNC|Parainfluenza virus 3 Ab|Parainfluenza virus 3 Ab
C0879993|T201|COMP|22440-2|LNC|Pasteurella multocida Ab|Pasteurella multocida Ab
C0879994|T201|COMP|22443-6|LNC|Plasmodium ovale Ab|Plasmodium ovale Ab
C0879995|T201|COMP|22444-4|LNC|Plasmodium vivax Ab|Plasmodium vivax Ab
C0879996|T201|COMP|22445-1|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C0879997|T201|COMP|22447-7|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C0879998|T201|COMP|22448-5|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C0879999|T201|COMP|22449-3|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C0880001|T201|COMP|22452-7|LNC|Pseudorabies virus Ab|Pseudorabies virus Ab
C0880002|T201|COMP|22453-5|LNC|Pseudorabies virus Ab|Pseudorabies virus Ab
C0880003|T201|COMP|22455-0|LNC|Pseudorabies virus.HerdCheck gene deletion Ab|Pseudorabies virus.HerdCheck gene deletion Ab
C0880004|T201|COMP|22456-8|LNC|Pseudorabies virus.OmniMark gene deletion Ab|Pseudorabies virus.OmniMark gene deletion Ab
C0880005|T201|COMP|22457-6|LNC|Pseudorabies virus.Tolvid gene deletion Ab|Pseudorabies virus.Tolvid gene deletion Ab
C0880006|T201|COMP|22458-4|LNC|Rabies virus Ab|Rabies virus Ab
C0880007|T201|COMP|22459-2|LNC|Reagin Ab|Reagin Ab
C0880008|T201|COMP|22460-0|LNC|Reagin Ab|Reagin Ab
C0880009|T201|COMP|22461-8|LNC|Reagin Ab|Reagin Ab
C0880010|T201|COMP|22462-6|LNC|Reagin Ab|Reagin Ab
C0880011|T201|COMP|22463-4|LNC|Reagin Ab|Reagin Ab
C0880012|T201|COMP|22465-9|LNC|Reovirus Ab|Reovirus Ab
C0880013|T201|COMP|22466-7|LNC|Respiratory syncytial virus Ab|Respiratory syncytial virus Ab
C0880014|T201|COMP|22467-5|LNC|Respiratory syncytial virus Ab.IgM|Respiratory syncytial virus Ab.IgM
C0880015|T201|COMP|22468-3|LNC|Rickettsia (Proteus OX19) Ab|Rickettsia (Proteus OX19) Ab
C0880016|T201|COMP|22469-1|LNC|Rickettsia (Proteus OX19) Ab|Rickettsia (Proteus OX19) Ab
C0880017|T201|COMP|22470-9|LNC|Rickettsia (Proteus OX2) Ab|Rickettsia (Proteus OX2) Ab
C0880018|T201|COMP|22471-7|LNC|Rickettsia (Proteus OX2) Ab|Rickettsia (Proteus OX2) Ab
C0880019|T201|COMP|22472-5|LNC|Rickettsia (Proteus OXK) Ab|Rickettsia (Proteus OXK) Ab
C0880020|T201|COMP|22473-3|LNC|Rickettsia (Proteus OXK) Ab|Rickettsia (Proteus OXK) Ab
C0880021|T201|COMP|22474-1|LNC|Rickettsia spotted fever group Ab|Rickettsia spotted fever group Ab
C0880022|T201|COMP|22475-8|LNC|Rickettsia spotted fever group Ab|Rickettsia spotted fever group Ab
C0880023|T201|COMP|22476-6|LNC|Rickettsia spotted fever group Ab.IgG|Rickettsia spotted fever group Ab.IgG
C0880024|T201|COMP|22477-4|LNC|Rickettsia spotted fever group Ab.IgG|Rickettsia spotted fever group Ab.IgG
C0880025|T201|COMP|22478-2|LNC|Rickettsia spotted fever group Ab.IgM|Rickettsia spotted fever group Ab.IgM
C0880026|T201|COMP|22479-0|LNC|Rickettsia spotted fever group Ab.IgM|Rickettsia spotted fever group Ab.IgM
C0880027|T201|COMP|22481-6|LNC|Rickettsia typhus group Ab.IgM|Rickettsia typhus group Ab.IgM
C0880028|T201|COMP|22482-4|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C0880029|T201|COMP|22483-2|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C0880030|T201|COMP|22484-0|LNC|Rickettsia sp Ab|Rickettsia sp Ab
C0880031|T201|COMP|22485-7|LNC|Orientia tsutsugamushi Ab|Orientia tsutsugamushi Ab
C0880032|T201|COMP|22486-5|LNC|Rickettsia typhi Ab|Rickettsia typhi Ab
C0880033|T201|COMP|22487-3|LNC|Rickettsia typhi Ab.IgA|Rickettsia typhi Ab.IgA
C0880034|T201|COMP|22488-1|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C0880035|T201|COMP|22489-9|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C0880036|T201|COMP|22490-7|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C0880037|T201|COMP|22491-5|LNC|Rickettsia typhus group Ab|Rickettsia typhus group Ab
C0880038|T201|COMP|22492-3|LNC|Rickettsia typhus group Ab|Rickettsia typhus group Ab
C0880039|T201|COMP|22493-1|LNC|Rickettsia typhus group Ab.IgG|Rickettsia typhus group Ab.IgG
C0880040|T201|COMP|22494-9|LNC|Rickettsia typhus group Ab.IgM|Rickettsia typhus group Ab.IgM
C0880041|T201|COMP|22495-6|LNC|Rotavirus Ab|Rotavirus Ab
C0880042|T201|COMP|22496-4|LNC|Rubella virus Ab|Rubella virus Ab
C0880043|T201|COMP|22497-2|LNC|Rubella virus Ab|Rubella virus Ab
C0880044|T201|COMP|22498-0|LNC|Measles virus Ab|Measles virus Ab
C0880045|T201|COMP|22500-3|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0880046|T201|COMP|22501-1|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0880047|T201|COMP|22503-7|LNC|Measles virus Ab.IgG^1st specimen|Measles virus Ab.IgG^1st specimen
C0880048|T201|COMP|22504-5|LNC|Measles virus Ab.IgG^2nd specimen|Measles virus Ab.IgG^2nd specimen
C0880049|T201|COMP|22505-2|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C0880050|T201|COMP|22507-8|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0880051|T201|COMP|22509-4|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0880052|T201|COMP|22511-0|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C0880053|T201|COMP|22512-8|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C0880054|T201|COMP|22513-6|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C0880055|T201|COMP|22514-4|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C0880056|T201|COMP|22515-1|LNC|Salmonella arizonae Ab|Salmonella arizonae Ab
C0880057|T201|COMP|22518-5|LNC|Salmonella paratyphi A H Ab|Salmonella paratyphi A H Ab
C0880058|T201|COMP|22519-3|LNC|Salmonella paratyphi A O Ab|Salmonella paratyphi A O Ab
C0880059|T201|COMP|22521-9|LNC|Salmonella paratyphi B H Ab|Salmonella paratyphi B H Ab
C0880060|T201|COMP|22522-7|LNC|Salmonella paratyphi B H Ab|Salmonella paratyphi B H Ab
C0880061|T201|COMP|22523-5|LNC|Salmonella paratyphi B O Ab|Salmonella paratyphi B O Ab
C0880062|T201|COMP|22524-3|LNC|Salmonella paratyphi C H Ab|Salmonella paratyphi C H Ab
C0880063|T201|COMP|22526-8|LNC|Salmonella pullorum Ab|Salmonella pullorum Ab
C0880064|T201|COMP|22527-6|LNC|Salmonella sp Ab|Salmonella sp Ab
C0880065|T201|COMP|22528-4|LNC|Salmonella typhi D Ab|Salmonella typhi D Ab
C0880066|T201|COMP|22529-2|LNC|Salmonella typhi H Ab|Salmonella typhi H Ab
C0880067|T201|COMP|22530-0|LNC|Salmonella typhi little d Ab|Salmonella typhi little d Ab
C0880068|T201|COMP|22531-8|LNC|Salmonella typhimurium Ab|Salmonella typhimurium Ab
C0880069|T201|COMP|22532-6|LNC|Sarcocystis neurona Ab|Sarcocystis neurona Ab
C0880070|T201|COMP|22533-4|LNC|Sarcocystis neurona Ab|Sarcocystis neurona Ab
C0880071|T201|COMP|22535-9|LNC|Schistosoma japonicum Ab|Schistosoma japonicum Ab
C0880072|T201|COMP|22536-7|LNC|Schistosoma mansoni Ab|Schistosoma mansoni Ab
C0880073|T201|COMP|22537-5|LNC|Shigella boydii Ab|Shigella boydii Ab
C0880074|T201|COMP|22538-3|LNC|Shigella dysenteriae Ab|Shigella dysenteriae Ab
C0880075|T201|COMP|22539-1|LNC|Shigella flexneri Ab|Shigella flexneri Ab
C0880076|T201|COMP|22540-9|LNC|Shigella sonnei Ab|Shigella sonnei Ab
C0880077|T201|COMP|22541-7|LNC|Streptococcus pneumoniae 1 Ab.IgG|Streptococcus pneumoniae 1 Ab.IgG
C0880078|T201|COMP|22542-5|LNC|Streptococcus pneumoniae 12 Ab.IgG|Streptococcus pneumoniae 12 Ab.IgG
C0880079|T201|COMP|22543-3|LNC|Streptococcus pneumoniae 14 Ab.IgG|Streptococcus pneumoniae 14 Ab.IgG
C0880080|T201|COMP|13155-7|LNC|Streptococcus pneumoniae 14 Ab^1st specimen|Streptococcus pneumoniae 14 Ab^1st specimen
C0880081|T201|COMP|22545-8|LNC|Streptococcus pneumoniae 14 Ab^2nd specimen|Streptococcus pneumoniae 14 Ab^2nd specimen
C0880083|T201|COMP|22547-4|LNC|Streptococcus pneumoniae 19 Ab.IgG|Streptococcus pneumoniae 19 Ab.IgG
C0880084|T201|COMP|22548-2|LNC|Streptococcus pneumoniae 23 Ab.IgG|Streptococcus pneumoniae 23 Ab.IgG
C0880085|T201|COMP|22549-0|LNC|Streptococcus pneumoniae 3 Ab.IgG|Streptococcus pneumoniae 3 Ab.IgG
C0880086|T201|COMP|22550-8|LNC|Streptococcus pneumoniae 6+26 Ab.IgG|Streptococcus pneumoniae 6+26 Ab.IgG
C0880087|T201|COMP|22551-6|LNC|Streptococcus pneumoniae 7 Ab.IgG|Streptococcus pneumoniae 7 Ab.IgG
C0880092|T201|COMP|22556-5|LNC|Streptococcus pneumoniae 8 Ab.IgG|Streptococcus pneumoniae 8 Ab.IgG
C0880093|T201|COMP|22557-3|LNC|Streptococcus pneumoniae 9 Ab|Streptococcus pneumoniae 9 Ab
C0880094|T201|COMP|22558-1|LNC|Streptococcus pneumoniae 9 Ab.IgG|Streptococcus pneumoniae 9 Ab.IgG
C0880095|T201|COMP|13151-6|LNC|Streptococcus pneumoniae 9 Ab^1st specimen|Streptococcus pneumoniae 9 Ab^1st specimen
C0880097|T201|COMP|13152-4|LNC|Streptococcus pneumoniae 9 Ab^2nd specimen|Streptococcus pneumoniae 9 Ab^2nd specimen
C0880098|T201|COMP|22562-3|LNC|Streptococcus pneumoniae Ab.IgG^1st specimen|Streptococcus pneumoniae Ab.IgG^1st specimen
C0880099|T201|COMP|22565-6|LNC|Streptococcus pneumoniae group B Ab|Streptococcus pneumoniae group B Ab
C0880100|T201|COMP|22566-4|LNC|Streptococcus pyogenes enzyme Ab|Streptococcus pyogenes enzyme Ab
C0880101|T201|COMP|22567-2|LNC|Streptococcus pyogenes enzyme Ab|Streptococcus pyogenes enzyme Ab
C0880102|T201|COMP|22568-0|LNC|Streptolysin O Ab|Streptolysin O Ab
C0880103|T201|COMP|22569-8|LNC|Strongyloides sp Ab|Strongyloides sp Ab
C0880104|T201|COMP|22571-4|LNC|Teichoate Ab|Teichoate Ab
C0880106|T201|COMP|22573-0|LNC|Thermoactinomyces vulgaris Ab|Thermoactinomyces vulgaris Ab
C0880107|T201|COMP|13276-1|LNC|Toxocara canis Ab.IgA|Toxocara canis Ab.IgA
C0880108|T201|COMP|13275-3|LNC|Toxocara canis Ab.IgM|Toxocara canis Ab.IgM
C0880109|T201|COMP|22577-1|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C0880110|T201|COMP|22578-9|LNC|Toxoplasma gondii Ab.IgA|Toxoplasma gondii Ab.IgA
C0880111|T201|COMP|22579-7|LNC|Toxoplasma gondii Ab.IgA+IgE|Toxoplasma gondii Ab.IgA+IgE
C0880112|T201|COMP|22580-5|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0880113|T201|COMP|22581-3|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0880114|T201|COMP|22582-1|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0880115|T201|COMP|22584-7|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0880116|T201|COMP|22585-4|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0880117|T201|COMP|22586-2|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0880118|T201|COMP|22587-0|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0880119|T201|COMP|22588-8|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0880120|T201|COMP|22589-6|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0880121|T201|COMP|22590-4|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0880122|T201|COMP|22591-2|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C0880123|T201|COMP|22592-0|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C0880124|T201|COMP|22593-8|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C0880125|T201|COMP|22594-6|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C0880126|T201|COMP|22595-3|LNC|Trichinella spiralis Ab|Trichinella spiralis Ab
C0880127|T201|COMP|22599-5|LNC|Trypanosoma cruzi Ab|Trypanosoma cruzi Ab
C0880128|T201|COMP|22600-1|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C0880129|T201|COMP|22601-9|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0880130|T201|COMP|22602-7|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0880131|T201|COMP|22603-5|LNC|Varicella zoster virus Ab.IgG^1st specimen|Varicella zoster virus Ab.IgG^1st specimen
C0880132|T201|COMP|22604-3|LNC|Varicella zoster virus Ab.IgG^2nd specimen|Varicella zoster virus Ab.IgG^2nd specimen
C0880133|T201|COMP|22605-0|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0880134|T201|COMP|22606-8|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0880135|T201|COMP|22607-6|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C0880136|T201|COMP|22608-4|LNC|Escherichia coli verotoxin 1 Ab|Escherichia coli verotoxin 1 Ab
C0880137|T201|COMP|22609-2|LNC|Escherichia coli verotoxin 2 Ab|Escherichia coli verotoxin 2 Ab
C0880138|T201|COMP|22610-0|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0880139|T201|COMP|22611-8|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0880140|T201|COMP|17770-9|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0880141|T201|COMP|22613-4|LNC|Western equine encephalitis virus Ab.IgG|Western equine encephalitis virus Ab.IgG
C0880142|T201|COMP|22614-2|LNC|Western equine encephalitis virus Ab.IgG|Western equine encephalitis virus Ab.IgG
C0880143|T201|COMP|22615-9|LNC|Western equine encephalitis virus Ab.IgM|Western equine encephalitis virus Ab.IgM
C0880144|T201|COMP|22616-7|LNC|Western equine encephalitis virus Ab.IgM|Western equine encephalitis virus Ab.IgM
C0880145|T201|COMP|22617-5|LNC|Wuchereria bancrofti Ab|Wuchereria bancrofti Ab
C0880146|T201|COMP|22619-1|LNC|Yersinia enterocolitica Ab.IgA|Yersinia enterocolitica Ab.IgA
C0880147|T201|COMP|22620-9|LNC|Yersinia enterocolitica Ab.IgG|Yersinia enterocolitica Ab.IgG
C0880148|T201|COMP|22621-7|LNC|Yersinia enterocolitica Ab.IgM|Yersinia enterocolitica Ab.IgM
C0880149|T201|COMP|22624-1|LNC|Xylose^2H post 5 g xylose PO|Xylose^2H post 5 g xylose PO
C0880150|T201|COMP|22626-6|LNC|Xylose^post 25 g xylose PO|Xylose^post 25 g xylose PO
C0880151|T201|COMP|22628-2|LNC|Xylose^post 25 g xylose PO|Xylose^post 25 g xylose PO
C0880152|T201|COMP|22629-0|LNC|Xylose^post 5 g xylose PO|Xylose^post 5 g xylose PO
C0880153|T201|COMP|22630-8|LNC|Xylose/Xylose.dose^post 25 g xylose PO|Xylose/Xylose.dose^post 25 g xylose PO
C0880154|T201|COMP|22632-4|LNC|Xylose/Xylose.dose^post dose xylose PO|Xylose/Xylose.dose^post dose xylose PO
C0880161|T201|COMP|22641-5|LNC|Glutamine|Glutamine
C0880162|T201|COMP|22642-3|LNC|Tyrosine|Tyrosine
C0880163|T201|COMP|22643-1|LNC|Threonine|Threonine
C0880164|T201|COMP|22644-9|LNC|Serine|Serine
C0880165|T201|COMP|22646-4|LNC|Phenylalanine|Phenylalanine
C0880166|T201|COMP|22647-2|LNC|Ornithine|Ornithine
C0880167|T201|COMP|22648-0|LNC|Methionine|Methionine
C0880168|T201|COMP|22649-8|LNC|Valine|Valine
C0880169|T201|COMP|22650-6|LNC|Glycine|Glycine
C0880170|T201|COMP|22651-4|LNC|Lysine|Lysine
C0880171|T201|COMP|22652-2|LNC|Glutamate|Glutamate
C0880172|T201|COMP|22653-0|LNC|Cystine|Cystine
C0880173|T201|COMP|22654-8|LNC|Citrulline|Citrulline
C0880174|T201|COMP|22655-5|LNC|Aspartate|Aspartate
C0880175|T201|COMP|22656-3|LNC|Arginine|Arginine
C0880176|T201|COMP|22657-1|LNC|Alanine|Alanine
C0880177|T201|COMP|22658-9|LNC|Alloisoleucine|Alloisoleucine
C0880178|T201|COMP|22659-7|LNC|Isoleucine|Isoleucine
C0880179|T201|COMP|22660-5|LNC|Homocystine|Homocystine
C0880180|T201|COMP|22661-3|LNC|Coproporphyrin|Coproporphyrin
C0880181|T201|COMP|22662-1|LNC|Uroporphyrin|Uroporphyrin
C0880182|T201|COMP|22663-9|LNC|Estrone|Estrone
C0880183|T201|COMP|22665-4|LNC|Bilirubin.albumin bound|Bilirubin.albumin bound
C0880184|T201|COMP|22666-2|LNC|Busulfan|Busulfan
C0880185|T201|COMP|15066-4|LNC|Fatty acids.nonesterified|Fatty acids.nonesterified
C0880186|T201|COMP|22668-8|LNC|Propylene glycol|Propylene glycol
C0880187|T201|COMP|20642-5|LNC|Glutamate|Glutamate
C0880188|T201|COMP|22670-4|LNC|Alloisoleucine|Alloisoleucine
C0880189|T201|COMP|22671-2|LNC|Phytanate|Phytanate
C0880190|T201|COMP|22672-0|LNC|Cystine|Cystine
C0880191|T201|COMP|20646-6|LNC|Homocystine|Homocystine
C0880192|T201|COMP|22674-6|LNC|Transferrin|Transferrin
C0880193|T201|COMP|22675-3|LNC|Angiotensin converting enzyme|Angiotensin converting enzyme
C0880194|T201|COMP|22676-1|LNC|7-Dehydrocholesterol|7-Dehydrocholesterol
C0880195|T201|COMP|22678-7|LNC|Ethylene glycol|Ethylene glycol
C0880196|T201|COMP|22679-5|LNC|Lysine/Creatinine|Lysine/Creatinine
C0880197|T201|COMP|22681-1|LNC|Methionine/Creatinine|Methionine/Creatinine
C0880198|T201|COMP|22682-9|LNC|Ornithine/Creatinine|Ornithine/Creatinine
C0880199|T201|COMP|22685-2|LNC|Tyrosine/Creatinine|Tyrosine/Creatinine
C0880200|T201|COMP|22686-0|LNC|Protoporphyrin|Protoporphyrin
C0880201|T201|COMP|22687-8|LNC|Cystine/Creatinine|Cystine/Creatinine
C0880202|T201|COMP|22688-6|LNC|Threonine/Creatinine|Threonine/Creatinine
C0880203|T201|COMP|22691-0|LNC|Aspartate/Creatinine|Aspartate/Creatinine
C0880204|T201|COMP|22693-6|LNC|Leucine/Creatinine|Leucine/Creatinine
C0880205|T201|COMP|22694-4|LNC|Citrulline/Creatinine|Citrulline/Creatinine
C0880206|T201|COMP|22695-1|LNC|Carnitine/Creatinine|Carnitine/Creatinine
C0880207|T201|COMP|22696-9|LNC|Cadmium/Creatinine|Cadmium/Creatinine
C0880208|T201|COMP|22698-5|LNC|Alanine/Creatinine|Alanine/Creatinine
C0880209|T201|COMP|22699-3|LNC|Alloisoleucine/Creatinine|Alloisoleucine/Creatinine
C0880210|T201|COMP|22700-9|LNC|Urea|Urea
C0880211|T201|COMP|22701-7|LNC|Salicylates|Salicylates
C0880212|T201|COMP|22702-5|LNC|Ketones|Ketones
C0880213|T201|COMP|22703-3|LNC|Histidine/Creatinine|Histidine/Creatinine
C0880214|T201|COMP|22705-8|LNC|Glucose|Glucose
C0880215|T201|COMP|22706-6|LNC|Isoleucine/Creatinine|Isoleucine/Creatinine
C0880216|T201|COMP|22707-4|LNC|Homocystine/Creatinine|Homocystine/Creatinine
C0880217|T201|COMP|22709-0|LNC|Glycine/Creatinine|Glycine/Creatinine
C0880218|T201|COMP|22710-8|LNC|Glutamine/Creatinine|Glutamine/Creatinine
C0880219|T201|COMP|22711-6|LNC|Glutamate/Creatinine|Glutamate/Creatinine
C0880220|T201|COMP|22713-2|LNC|Lysine|Lysine
C0880221|T201|COMP|22714-0|LNC|Isoleucine|Isoleucine
C0880222|T201|COMP|22715-7|LNC|Homocystine|Homocystine
C0880223|T201|COMP|22716-5|LNC|Methionine|Methionine
C0880224|T201|COMP|22717-3|LNC|Histidine|Histidine
C0880225|T201|COMP|22718-1|LNC|Glycine|Glycine
C0880226|T201|COMP|22719-9|LNC|Leucine|Leucine
C0880227|T201|COMP|22720-7|LNC|Glutamine|Glutamine
C0880228|T201|COMP|22721-5|LNC|Glutamate|Glutamate
C0880229|T201|COMP|22722-3|LNC|Citrulline|Citrulline
C0880230|T201|COMP|22723-1|LNC|Aspartate|Aspartate
C0880231|T201|COMP|22724-9|LNC|Alanine|Alanine
C0880232|T201|COMP|22725-6|LNC|Ornithine|Ornithine
C0880233|T201|COMP|22727-2|LNC|Arginine|Arginine
C0880234|T201|COMP|22728-0|LNC|Cystine|Cystine
C0880235|T201|COMP|22729-8|LNC|Valine|Valine
C0880236|T201|COMP|22730-6|LNC|Alloisoleucine|Alloisoleucine
C0880237|T201|COMP|22731-4|LNC|Triglyceride|Triglyceride
C0880238|T201|COMP|22732-2|LNC|Salicylates|Salicylates
C0880239|T201|COMP|22733-0|LNC|Phosphate|Phosphate
C0880240|T201|COMP|22734-8|LNC|Ethylene glycol|Ethylene glycol
C0880241|T201|COMP|22735-5|LNC|Bicarbonate|Bicarbonate
C0880242|T201|COMP|22736-3|LNC|Acetaminophen|Acetaminophen
C0880243|T201|COMP|22737-1|LNC|Phenylalanine|Phenylalanine
C0880244|T201|COMP|22738-9|LNC|Urea|Urea
C0880245|T201|COMP|22739-7|LNC|Tyrosine|Tyrosine
C0880246|T201|COMP|22740-5|LNC|Threonine|Threonine
C0880247|T201|COMP|22741-3|LNC|Serine|Serine
C0880248|T201|COMP|22742-1|LNC|Propylene glycol|Propylene glycol
C0880249|T201|COMP|22743-9|LNC|Proline|Proline
C0880250|T201|COMP|22744-7|LNC|Copper|Copper
C0880251|T201|COMP|22745-4|LNC|Ethanol|Ethanol
C0880252|T201|COMP|22746-2|LNC|Gentamicin^peak|Gentamicin^peak
C0880253|T201|COMP|22748-8|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C0880254|T201|COMP|22749-6|LNC|Amylase.pancreatic|Amylase.pancreatic
C0880255|T201|COMP|22750-4|LNC|Tobramycin^random|Tobramycin^random
C0880256|T201|COMP|22753-8|LNC|Iron binding capacity.unsaturated|Iron binding capacity.unsaturated
C0880257|T201|COMP|22754-6|LNC|Dibucaine number|Dibucaine number
C0880258|T201|COMP|22756-1|LNC|HLA-DR|HLA-DR
C0880259|T201|COMP|22758-7|LNC|Plasminogen activator inhibitor 1 Ag|Plasminogen activator inhibitor 1 Ag
C0880260|T201|COMP|22759-5|LNC|Platelet Ab|Platelet Ab
C0880261|T201|COMP|22761-1|LNC|Pristanate|Pristanate
C0880263|T201|COMP|22763-7|LNC|Ammonia|Ammonia
C0880264|T201|COMP|22765-2|LNC|Adult fly identified|Adult fly identified
C0880265|T201|COMP|22766-0|LNC|African horse sickness virus Ab|African horse sickness virus Ab
C0880266|T201|COMP|22767-8|LNC|African horse sickness virus Ab|African horse sickness virus Ab
C0880267|T201|COMP|22768-6|LNC|African horse sickness virus Ab|African horse sickness virus Ab
C0880268|T201|COMP|22769-4|LNC|African horse sickness virus Ab|African horse sickness virus Ab
C0880269|T201|COMP|22770-2|LNC|African horse sickness virus Ab|African horse sickness virus Ab
C0880270|T201|COMP|22771-0|LNC|African horse sickness virus Ab|African horse sickness virus Ab
C0880271|T201|COMP|22772-8|LNC|African horse sickness virus Ag|African horse sickness virus Ag
C0880272|T201|COMP|22774-4|LNC|African horse sickness virus RNA|African horse sickness virus RNA
C0880273|T201|COMP|22775-1|LNC|African horse sickness virus serotype|African horse sickness virus serotype
C0880274|T201|COMP|22776-9|LNC|African horse sickness virus serotype|African horse sickness virus serotype
C0880275|T201|COMP|22777-7|LNC|African swine fever virus Ab|African swine fever virus Ab
C0880276|T201|COMP|22779-3|LNC|African swine fever virus Ab|African swine fever virus Ab
C0880277|T201|COMP|22780-1|LNC|African swine fever virus Ab|African swine fever virus Ab
C0880278|T201|COMP|22781-9|LNC|African swine fever virus Ag|African swine fever virus Ag
C0880279|T201|COMP|22782-7|LNC|African swine fever virus Ag|African swine fever virus Ag
C0880280|T201|COMP|22783-5|LNC|African swine fever virus Ag|African swine fever virus Ag
C0880281|T201|COMP|22784-3|LNC|African swine fever virus Ag|African swine fever virus Ag
C0880282|T201|COMP|22785-0|LNC|African swine fever virus DNA|African swine fever virus DNA
C0880283|T201|COMP|22786-8|LNC|Alcelaphine herpesvirus 1 Ab|Alcelaphine herpesvirus 1 Ab
C0880284|T201|COMP|22787-6|LNC|Alcelaphine herpesvirus 1 Ab|Alcelaphine herpesvirus 1 Ab
C0880285|T201|COMP|22788-4|LNC|Alcelaphine herpesvirus 1 Ab|Alcelaphine herpesvirus 1 Ab
C0880286|T201|COMP|22789-2|LNC|Alcelaphine herpesvirus 1 Ag|Alcelaphine herpesvirus 1 Ag
C0880287|T201|COMP|22790-0|LNC|Alcelaphine herpesvirus 1 Ag|Alcelaphine herpesvirus 1 Ag
C0880288|T201|COMP|22792-6|LNC|Aleutian disease virus Ab|Aleutian disease virus Ab
C0880289|T201|COMP|22793-4|LNC|Aleutian disease virus Ab|Aleutian disease virus Ab
C0880290|T201|COMP|22794-2|LNC|Anaplasma marginale Ab|Anaplasma marginale Ab
C0880291|T201|COMP|22795-9|LNC|Anaplasma marginale Ab|Anaplasma marginale Ab
C0880292|T201|COMP|22796-7|LNC|Anaplasma marginale Ag|Anaplasma marginale Ag
C0880293|T201|COMP|22797-5|LNC|Anaplasma marginale DNA|Anaplasma marginale DNA
C0880294|T201|COMP|22798-3|LNC|Anaplasma marginale rRNA|Anaplasma marginale rRNA
C0880295|T201|COMP|22799-1|LNC|Anaplasma sp identified|Anaplasma sp identified
C0880296|T201|COMP|22800-7|LNC|Anaplasma sp identified|Anaplasma sp identified
C0880297|T201|COMP|22801-5|LNC|Infectious bronchitis virus Ab|Infectious bronchitis virus Ab
C0880298|T201|COMP|22802-3|LNC|Infectious bronchitis virus Ab|Infectious bronchitis virus Ab
C0880299|T201|COMP|22803-1|LNC|Infectious bronchitis virus Ab|Infectious bronchitis virus Ab
C0880300|T201|COMP|22804-9|LNC|Infectious bronchitis virus Ab|Infectious bronchitis virus Ab
C0880301|T201|COMP|22805-6|LNC|Infectious bronchitis virus Ag|Infectious bronchitis virus Ag
C0880302|T201|COMP|22806-4|LNC|Infectious bronchitis virus Ag|Infectious bronchitis virus Ag
C0880303|T201|COMP|22807-2|LNC|Infectious bronchitis virus Ag|Infectious bronchitis virus Ag
C0880304|T201|COMP|22808-0|LNC|Infectious bronchitis virus|Infectious bronchitis virus
C0880305|T201|COMP|22809-8|LNC|Infectious bronchitis virus RNA|Infectious bronchitis virus RNA
C0880306|T201|COMP|22810-6|LNC|Infectious bronchitis virus RNA|Infectious bronchitis virus RNA
C0880307|T201|COMP|22811-4|LNC|Avian infectious laryngotracheitis virus|Avian infectious laryngotracheitis virus
C0880308|T201|COMP|22812-2|LNC|Avian infectious laryngotracheitis virus|Avian infectious laryngotracheitis virus
C0880309|T201|COMP|22813-0|LNC|Avian infectious laryngotracheitis virus Ab|Avian infectious laryngotracheitis virus Ab
C0880310|T201|COMP|22815-5|LNC|Avian infectious laryngotracheitis virus Ab|Avian infectious laryngotracheitis virus Ab
C0880311|T201|COMP|22816-3|LNC|Avian infectious laryngotracheitis virus Ag|Avian infectious laryngotracheitis virus Ag
C0880312|T201|COMP|22817-1|LNC|Avian infectious laryngotracheitis virus Ag|Avian infectious laryngotracheitis virus Ag
C0880313|T201|COMP|22818-9|LNC|Avian infectious laryngotracheitis virus Ag|Avian infectious laryngotracheitis virus Ag
C0880314|T201|COMP|22820-5|LNC|Avian orthoreovirus Ag|Avian orthoreovirus Ag
C0880315|T201|COMP|22821-3|LNC|Influenza virus A Ab|Influenza virus A Ab
C0880316|T201|COMP|22822-1|LNC|Influenza virus A Ab|Influenza virus A Ab
C0880317|T201|COMP|22823-9|LNC|Influenza virus A Ab|Influenza virus A Ab
C0880318|T201|COMP|22825-4|LNC|Influenza virus A Ag|Influenza virus A Ag
C0880319|T201|COMP|22827-0|LNC|Influenza virus A subtype|Influenza virus A subtype
C0880320|T201|COMP|22828-8|LNC|Influenza virus A subtype|Influenza virus A subtype
C0880321|T201|COMP|22830-4|LNC|Avian paramyxovirus 1 Ab|Avian paramyxovirus 1 Ab
C0880322|T201|COMP|22831-2|LNC|Avian paramyxovirus 1 Ag|Avian paramyxovirus 1 Ag
C0880323|T201|COMP|22832-0|LNC|Avian paramyxovirus 1 identified|Avian paramyxovirus 1 identified
C0880324|T201|COMP|22833-8|LNC|Avian paramyxovirus 1|Avian paramyxovirus 1
C0880325|T201|COMP|22836-1|LNC|Avian pox virus|Avian pox virus
C0880326|T201|COMP|22837-9|LNC|Avian pox virus Ab|Avian pox virus Ab
C0880327|T201|COMP|22838-7|LNC|Avian pox virus Ab|Avian pox virus Ab
C0880328|T201|COMP|22839-5|LNC|Avian pox virus Ab|Avian pox virus Ab
C0880329|T201|COMP|22840-3|LNC|Avian pox virus Ab|Avian pox virus Ab
C0880330|T201|COMP|22841-1|LNC|Avian pox virus Ab|Avian pox virus Ab
C0880331|T201|COMP|22842-9|LNC|Avian pox virus DNA|Avian pox virus DNA
C0880332|T201|COMP|22843-7|LNC|Avian pox virus DNA|Avian pox virus DNA
C0880333|T201|COMP|22845-2|LNC|Babesia bigemina Ab|Babesia bigemina Ab
C0880334|T201|COMP|22846-0|LNC|Babesia bigemina Ab|Babesia bigemina Ab
C0880335|T201|COMP|22847-8|LNC|Babesia bovis Ab|Babesia bovis Ab
C0880336|T201|COMP|22848-6|LNC|Babesia bovis Ab|Babesia bovis Ab
C0880337|T201|COMP|22849-4|LNC|Babesia bovis Ab|Babesia bovis Ab
C0880338|T201|COMP|22850-2|LNC|Babesia caballi Ab|Babesia caballi Ab
C0880339|T201|COMP|22851-0|LNC|Babesia caballi Ab|Babesia caballi Ab
C0880340|T201|COMP|22104-4|LNC|Babesia caballi Ab|Babesia caballi Ab
C0880341|T201|COMP|22853-6|LNC|Babesia caballi rRNA|Babesia caballi rRNA
C0880342|T201|COMP|22854-4|LNC|Babesia divergens Ab|Babesia divergens Ab
C0880343|T201|COMP|22855-1|LNC|Babesia divergens Ab|Babesia divergens Ab
C0880344|T201|COMP|22856-9|LNC|Babesia sp rRNA|Babesia sp rRNA
C0880345|T201|COMP|22857-7|LNC|Babesia sp DNA|Babesia sp DNA
C0880346|T201|COMP|22858-5|LNC|Babesia sp identified|Babesia sp identified
C0880347|T201|COMP|22859-3|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0880348|T201|COMP|22860-1|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0880349|T201|COMP|22861-9|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0880350|T201|COMP|22862-7|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0880351|T201|COMP|22863-5|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0880352|T201|COMP|22864-3|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0880353|T201|COMP|22865-0|LNC|Bacillus anthracis Ab|Bacillus anthracis Ab
C0880354|T201|COMP|22866-8|LNC|Bacillus anthracis Ag|Bacillus anthracis Ag
C0880355|T201|COMP|22867-6|LNC|Bacillus anthracis Ag|Bacillus anthracis Ag
C0880356|T201|COMP|22869-2|LNC|Bluetongue virus Ag|Bluetongue virus Ag
C0880357|T201|COMP|22870-0|LNC|Bluetongue virus Ag|Bluetongue virus Ag
C0880358|T201|COMP|22871-8|LNC|Bluetongue virus Ag|Bluetongue virus Ag
C0880359|T201|COMP|22874-2|LNC|Bluetongue virus serotype|Bluetongue virus serotype
C0880360|T201|COMP|22875-9|LNC|Border disease virus Ab|Border disease virus Ab
C0880361|T201|COMP|22876-7|LNC|Border disease virus Ab|Border disease virus Ab
C0880362|T201|COMP|22878-3|LNC|Border disease virus Ab|Border disease virus Ab
C0880363|T201|COMP|22879-1|LNC|Border disease virus Ag|Border disease virus Ag
C0880364|T201|COMP|22880-9|LNC|Border disease virus Ag|Border disease virus Ag
C0880365|T201|COMP|22882-5|LNC|Border disease virus Ag|Border disease virus Ag
C0880366|T201|COMP|22883-3|LNC|Border disease virus RNA|Border disease virus RNA
C0880367|T201|COMP|22884-1|LNC|Border disease virus RNA|Border disease virus RNA
C0880368|T201|COMP|22885-8|LNC|Border disease virus RNA|Border disease virus RNA
C0880369|T201|COMP|22887-4|LNC|Bordetella bronchiseptica Ab|Bordetella bronchiseptica Ab
C0880370|T201|COMP|22888-2|LNC|Bordetella bronchiseptica Ag|Bordetella bronchiseptica Ag
C0880371|T201|COMP|22889-0|LNC|Bovine diarrhea virus Ab|Bovine diarrhea virus Ab
C0880372|T201|COMP|22891-6|LNC|Bovine diarrhea virus Ab|Bovine diarrhea virus Ab
C0880373|T201|COMP|22892-4|LNC|Bovine diarrhea virus Ab|Bovine diarrhea virus Ab
C0880374|T201|COMP|22893-2|LNC|Bovine diarrhea virus Ab|Bovine diarrhea virus Ab
C0880375|T201|COMP|22894-0|LNC|Bovine diarrhea virus Ab|Bovine diarrhea virus Ab
C0880376|T201|COMP|22896-5|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C0880377|T201|COMP|22897-3|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C0880378|T201|COMP|22898-1|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C0880379|T201|COMP|22899-9|LNC|Bovine diarrhea virus RNA|Bovine diarrhea virus RNA
C0880380|T201|COMP|22900-5|LNC|Bovine diarrhea virus RNA|Bovine diarrhea virus RNA
C0880381|T201|COMP|22901-3|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C0880382|T201|COMP|22902-1|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C0880383|T201|COMP|22903-9|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C0880384|T201|COMP|22904-7|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C0880385|T201|COMP|22905-4|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C0880386|T201|COMP|22906-2|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C0880387|T201|COMP|22907-0|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C0880388|T201|COMP|22908-8|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C0880389|T201|COMP|22909-6|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C0880390|T201|COMP|22910-4|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C0880391|T201|COMP|22911-2|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C0880392|T201|COMP|22912-0|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C0880393|T201|COMP|22913-8|LNC|Bovine herpesvirus 1 DNA|Bovine herpesvirus 1 DNA
C0880394|T201|COMP|22914-6|LNC|Bovine herpesvirus 1 DNA|Bovine herpesvirus 1 DNA
C0880395|T201|COMP|22915-3|LNC|Bovine leukemia virus Ab|Bovine leukemia virus Ab
C0880396|T201|COMP|22916-1|LNC|Bovine leukemia virus Ab|Bovine leukemia virus Ab
C0880397|T201|COMP|22917-9|LNC|Bovine leukemia virus Ag|Bovine leukemia virus Ag
C0880398|T201|COMP|22918-7|LNC|Bovine leukemia virus RNA|Bovine leukemia virus RNA
C0880399|T201|COMP|22919-5|LNC|Bovine leukemia virus RNA|Bovine leukemia virus RNA
C0880400|T201|COMP|22920-3|LNC|Brucella abortus Ab|Brucella abortus Ab
C0880401|T201|COMP|22921-1|LNC|Brucella abortus Ab|Brucella abortus Ab
C0880402|T201|COMP|22922-9|LNC|Brucella abortus Ab.IgG1|Brucella abortus Ab.IgG1
C0880403|T201|COMP|22923-7|LNC|Brucella abortus Ab.IgG1|Brucella abortus Ab.IgG1
C0880404|T201|COMP|22925-2|LNC|Brucella abortus Ab.IgG1|Brucella abortus Ab.IgG1
C0880405|T201|COMP|22926-0|LNC|Brucella abortus rRNA|Brucella abortus rRNA
C0880406|T201|COMP|22927-8|LNC|Brucella abortus DNA|Brucella abortus DNA
C0880407|T201|COMP|22928-6|LNC|Brucella canis Ab|Brucella canis Ab
C0880408|T201|COMP|22929-4|LNC|Brucella canis Ab|Brucella canis Ab
C0880409|T201|COMP|22930-2|LNC|Brucella canis Ab|Brucella canis Ab
C0880410|T201|COMP|22931-0|LNC|Brucella melitensis Ab|Brucella melitensis Ab
C0880411|T201|COMP|22933-6|LNC|Brucella melitensis Ab|Brucella melitensis Ab
C0880412|T201|COMP|22934-4|LNC|Brucella melitensis Ab|Brucella melitensis Ab
C0880413|T201|COMP|22935-1|LNC|Brucella melitensis Ab|Brucella melitensis Ab
C0880414|T201|COMP|22936-9|LNC|Brucella melitensis DNA|Brucella melitensis DNA
C0880415|T201|COMP|22938-5|LNC|Brucella ovis Ab|Brucella ovis Ab
C0880416|T201|COMP|22939-3|LNC|Brucella ovis Ab|Brucella ovis Ab
C0880419|T201|COMP|22943-5|LNC|Brucella sp Ag|Brucella sp Ag
C0880420|T201|COMP|22944-3|LNC|Brucella sp Ag|Brucella sp Ag
C0880421|T201|COMP|22946-8|LNC|Brucella sp Ag|Brucella sp Ag
C0880422|T201|COMP|22947-6|LNC|Brucella sp Ag|Brucella sp Ag
C0880423|T201|COMP|22948-4|LNC|Brucella sp Ag|Brucella sp Ag
C0880424|T201|COMP|22949-2|LNC|Brucella sp Ag|Brucella sp Ag
C0880425|T201|COMP|22950-0|LNC|Brucella suis Ab|Brucella suis Ab
C0880426|T201|COMP|22951-8|LNC|Brucella suis Ab|Brucella suis Ab
C0880427|T201|COMP|22952-6|LNC|Brucella suis Ab|Brucella suis Ab
C0880428|T201|COMP|22954-2|LNC|Brucella suis rRNA|Brucella suis rRNA
C0880429|T201|COMP|22955-9|LNC|Brucella suis DNA|Brucella suis DNA
C0880431|T201|COMP|22959-1|LNC|Burkholderia mallei Ab|Burkholderia mallei Ab
C0880434|T201|COMP|22962-5|LNC|Campylobacter fetus Ab|Campylobacter fetus Ab
C0880435|T201|COMP|22963-3|LNC|Campylobacter fetus Ab|Campylobacter fetus Ab
C0880436|T201|COMP|22964-1|LNC|Campylobacter fetus Ag|Campylobacter fetus Ag
C0880437|T201|COMP|22965-8|LNC|Campylobacter fetus Ag|Campylobacter fetus Ag
C0880438|T201|COMP|22966-6|LNC|Campylobacter fetus Ag|Campylobacter fetus Ag
C0880439|T201|COMP|22967-4|LNC|Campylobacter fetus subspecies venerealis Ab|Campylobacter fetus subspecies venerealis Ab
C0880440|T201|COMP|22968-2|LNC|Campylobacter fetus subspecies venerealis Ab|Campylobacter fetus subspecies venerealis Ab
C0880441|T201|COMP|22970-8|LNC|Campylobacter fetus subspecies venerealis Ab.IgA|Campylobacter fetus subspecies venerealis Ab.IgA
C0880442|T201|COMP|22971-6|LNC|Caprine arthritis encephalitis virus|Caprine arthritis encephalitis virus
C0880443|T201|COMP|22972-4|LNC|Caprine arthritis encephalitis virus Ab|Caprine arthritis encephalitis virus Ab
C0880444|T201|COMP|22973-2|LNC|Caprine arthritis encephalitis virus Ab|Caprine arthritis encephalitis virus Ab
C0880445|T201|COMP|22974-0|LNC|Caprine arthritis encephalitis virus Ab|Caprine arthritis encephalitis virus Ab
C0880446|T201|COMP|22975-7|LNC|Caprine arthritis encephalitis virus Ag|Caprine arthritis encephalitis virus Ag
C0880447|T201|COMP|22976-5|LNC|Caprine arthritis encephalitis virus Ag|Caprine arthritis encephalitis virus Ag
C0880448|T201|COMP|22977-3|LNC|Caprine arthritis encephalitis virus DNA|Caprine arthritis encephalitis virus DNA
C0880449|T201|COMP|22978-1|LNC|Caprine arthritis encephalitis virus DNA|Caprine arthritis encephalitis virus DNA
C0880450|T201|COMP|22979-9|LNC|Caprine herpesvirus 1 Ab|Caprine herpesvirus 1 Ab
C0880451|T201|COMP|22980-7|LNC|Caprine herpesvirus 1 Ab|Caprine herpesvirus 1 Ab
C0880452|T201|COMP|22981-5|LNC|Capripox virus|Capripox virus
C0880453|T201|COMP|22983-1|LNC|Capripox virus Ab|Capripox virus Ab
C0880454|T201|COMP|22984-9|LNC|Capripox virus Ab|Capripox virus Ab
C0880455|T201|COMP|22982-3|LNC|Capripox virus Ab|Capripox virus Ab
C0880456|T201|COMP|22986-4|LNC|Capripox virus Ag|Capripox virus Ag
C0880457|T201|COMP|22987-2|LNC|Capripox virus Ag|Capripox virus Ag
C0880458|T201|COMP|22988-0|LNC|Capripox virus Ag|Capripox virus Ag
C0880459|T201|COMP|22989-8|LNC|Capripox virus Ag|Capripox virus Ag
C0880460|T201|COMP|22990-6|LNC|Capripox virus Ag|Capripox virus Ag
C0880461|T201|COMP|22991-4|LNC|Capripox virus DNA|Capripox virus DNA
C0880462|T201|COMP|22993-0|LNC|Chlamydophila psittaci|Chlamydophila psittaci
C0880463|T201|COMP|22994-8|LNC|Chlamydophila psittaci Ab|Chlamydophila psittaci Ab
C0880464|T201|COMP|22995-5|LNC|Chlamydophila psittaci Ab|Chlamydophila psittaci Ab
C0880465|T201|COMP|22996-3|LNC|Chlamydophila psittaci Ab|Chlamydophila psittaci Ab
C0880466|T201|COMP|22997-1|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C0880467|T201|COMP|22999-7|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C0880468|T201|COMP|23001-1|LNC|Chlamydophila psittaci DNA|Chlamydophila psittaci DNA
C0880469|T201|COMP|23002-9|LNC|Classical swine fever virus Ab|Classical swine fever virus Ab
C0880470|T201|COMP|23003-7|LNC|Classical swine fever virus Ab|Classical swine fever virus Ab
C0880471|T201|COMP|23005-2|LNC|Classical swine fever virus Ag|Classical swine fever virus Ag
C0880472|T201|COMP|23007-8|LNC|Classical swine fever virus Ag|Classical swine fever virus Ag
C0880473|T201|COMP|23008-6|LNC|Classical swine fever virus RNA|Classical swine fever virus RNA
C0880474|T201|COMP|23009-4|LNC|Cowdria ruminantium|Cowdria ruminantium
C0880475|T201|COMP|23011-0|LNC|Cowdria ruminantium Ab|Cowdria ruminantium Ab
C0880476|T201|COMP|23012-8|LNC|Cowdria ruminantium Ab|Cowdria ruminantium Ab
C0880477|T201|COMP|23013-6|LNC|Cowdria ruminantium Ab|Cowdria ruminantium Ab
C0880478|T201|COMP|23014-4|LNC|Cowdria ruminantium DNA|Cowdria ruminantium DNA
C0880479|T201|COMP|23015-1|LNC|Cowdria ruminantium rRNA|Cowdria ruminantium rRNA
C0880480|T201|COMP|23016-9|LNC|Coxiella burnetii|Coxiella burnetii
C0880481|T201|COMP|23017-7|LNC|Coxiella burnetii Ab|Coxiella burnetii Ab
C0880482|T201|COMP|23019-3|LNC|Coxiella burnetii Ab|Coxiella burnetii Ab
C0880483|T201|COMP|23020-1|LNC|Coxiella burnetii Ab|Coxiella burnetii Ab
C0880484|T201|COMP|23021-9|LNC|Coxiella burnetii Ag|Coxiella burnetii Ag
C0880485|T201|COMP|23022-7|LNC|Coxiella burnetii Ag|Coxiella burnetii Ag
C0880486|T201|COMP|23023-5|LNC|Coxiella burnetii Ag|Coxiella burnetii Ag
C0880487|T201|COMP|23024-3|LNC|Coxiella burnetii DNA|Coxiella burnetii DNA
C0880488|T201|COMP|23025-0|LNC|Dermatophilus congolensis|Dermatophilus congolensis
C0880489|T201|COMP|23026-8|LNC|Dermatophilus congolensis Ab|Dermatophilus congolensis Ab
C0880490|T201|COMP|23027-6|LNC|Dermatophilus congolensis Ab|Dermatophilus congolensis Ab
C0880491|T201|COMP|23028-4|LNC|Dermatophilus congolensis Ag|Dermatophilus congolensis Ag
C0880492|T201|COMP|23029-2|LNC|Dirofilaria immitis Ag|Dirofilaria immitis Ag
C0880493|T201|COMP|23030-0|LNC|Duck enteritis virus|Duck enteritis virus
C0880494|T201|COMP|23031-8|LNC|Duck enteritis virus Ag|Duck enteritis virus Ag
C0880495|T201|COMP|23032-6|LNC|Duck enteritis virus Ag|Duck enteritis virus Ag
C0880496|T201|COMP|23033-4|LNC|Duck hepatitis virus 1 Ab|Duck hepatitis virus 1 Ab
C0880497|T201|COMP|23034-2|LNC|Duck hepatitis virus 1 Ab|Duck hepatitis virus 1 Ab
C0880498|T201|COMP|23035-9|LNC|Duck hepatitis virus 1 Ag|Duck hepatitis virus 1 Ag
C0880499|T201|COMP|23036-7|LNC|Duck hepatitis virus 2 Ab|Duck hepatitis virus 2 Ab
C0880500|T201|COMP|23037-5|LNC|Duck hepatitis virus 2 Ab|Duck hepatitis virus 2 Ab
C0880501|T201|COMP|23038-3|LNC|Duck hepatitis virus 2 Ag|Duck hepatitis virus 2 Ag
C0880502|T201|COMP|23039-1|LNC|Duck hepatitis virus 3 Ab|Duck hepatitis virus 3 Ab
C0880503|T201|COMP|23040-9|LNC|Duck hepatitis virus 3 Ab|Duck hepatitis virus 3 Ab
C0880504|T201|COMP|23041-7|LNC|Duck hepatitis virus 3 Ag|Duck hepatitis virus 3 Ag
C0880505|T201|COMP|23042-5|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0880506|T201|COMP|23043-3|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0880507|T201|COMP|23044-1|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0880508|T201|COMP|23045-8|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C0880509|T201|COMP|23048-2|LNC|Eastern equine encephalitis virus Ag|Eastern equine encephalitis virus Ag
C0880510|T201|COMP|23049-0|LNC|Eastern equine encephalitis virus Ag|Eastern equine encephalitis virus Ag
C0880511|T201|COMP|23050-8|LNC|Eastern equine encephalitis virus Ag|Eastern equine encephalitis virus Ag
C0880512|T201|COMP|23051-6|LNC|Eastern equine encephalitis virus RNA|Eastern equine encephalitis virus RNA
C0880513|T201|COMP|23053-2|LNC|Echinococcus sp Ag|Echinococcus sp Ag
C0880514|T201|COMP|23054-0|LNC|Ehrlichia canis Ab|Ehrlichia canis Ab
C0880515|T201|COMP|23055-7|LNC|Ehrlichia risticii Ab|Ehrlichia risticii Ab
C0880516|T201|COMP|23056-5|LNC|Ehrlichia risticii Ab|Ehrlichia risticii Ab
C0880517|T201|COMP|23057-3|LNC|Ephemeral fever virus Ab|Ephemeral fever virus Ab
C0880518|T201|COMP|23059-9|LNC|Epizootic hemorrhagic disease virus Ab|Epizootic hemorrhagic disease virus Ab
C0880519|T201|COMP|23060-7|LNC|Epizootic hemorrhagic disease virus Ab|Epizootic hemorrhagic disease virus Ab
C0880520|T201|COMP|23061-5|LNC|Epizootic hemorrhagic disease virus Ag|Epizootic hemorrhagic disease virus Ag
C0880521|T201|COMP|23063-1|LNC|Epizootic hemorrhagic disease virus Alberta Ab|Epizootic hemorrhagic disease virus Alberta Ab
C0880522|T201|COMP|23064-9|LNC|Epizootic hemorrhagic disease virus Alberta Ab|Epizootic hemorrhagic disease virus Alberta Ab
C0880523|T201|COMP|23065-6|LNC|Epizootic hemorrhagic disease virus New Jersey Ab|Epizootic hemorrhagic disease virus New Jersey Ab
C0880524|T201|COMP|23066-4|LNC|Epizootic hemorrhagic disease virus New Jersey Ab|Epizootic hemorrhagic disease virus New Jersey Ab
C0880525|T201|COMP|23068-0|LNC|Equine arteritis virus Ab|Equine arteritis virus Ab
C0880526|T201|COMP|23069-8|LNC|Equine arteritis virus Ab|Equine arteritis virus Ab
C0880527|T201|COMP|23070-6|LNC|Equine arteritis virus Ab|Equine arteritis virus Ab
C0880528|T201|COMP|23071-4|LNC|Equine arteritis virus Ab|Equine arteritis virus Ab
C0880529|T201|COMP|23072-2|LNC|Equine arteritis virus Ab|Equine arteritis virus Ab
C0880530|T201|COMP|23073-0|LNC|Equine arteritis virus Ab|Equine arteritis virus Ab
C0880531|T201|COMP|23075-5|LNC|Equine arteritis virus Ag|Equine arteritis virus Ag
C0880532|T201|COMP|23076-3|LNC|Equine arteritis virus Ag|Equine arteritis virus Ag
C0880533|T201|COMP|23077-1|LNC|Equine arteritis virus Ag|Equine arteritis virus Ag
C0880534|T201|COMP|23078-9|LNC|Equine arteritis virus Ag|Equine arteritis virus Ag
C0880535|T201|COMP|23079-7|LNC|Equine arteritis virus RNA|Equine arteritis virus RNA
C0880536|T201|COMP|23080-5|LNC|Equine herpesvirus 1 Ag|Equine herpesvirus 1 Ag
C0880537|T201|COMP|23081-3|LNC|Equine herpesvirus 1 Ag|Equine herpesvirus 1 Ag
C0880538|T201|COMP|23082-1|LNC|Equine herpesvirus 1 DNA|Equine herpesvirus 1 DNA
C0880539|T201|COMP|23083-9|LNC|Equine herpesvirus 1 DNA|Equine herpesvirus 1 DNA
C0880540|T201|COMP|23084-7|LNC|Equine herpesvirus 1 DNA|Equine herpesvirus 1 DNA
C0880541|T201|COMP|23085-4|LNC|Equine herpesvirus 1+4 Ab|Equine herpesvirus 1+4 Ab
C0880542|T201|COMP|23086-2|LNC|Equine herpesvirus 1+4 Ab|Equine herpesvirus 1+4 Ab
C0880543|T201|COMP|23087-0|LNC|Equine herpesvirus 1+4 Ab|Equine herpesvirus 1+4 Ab
C0880544|T201|COMP|23088-8|LNC|Equine herpesvirus 1+4 Ab|Equine herpesvirus 1+4 Ab
C0880545|T201|COMP|23089-6|LNC|Equine herpesvirus 1+4 Ab|Equine herpesvirus 1+4 Ab
C0880546|T201|COMP|23090-4|LNC|Equine herpesvirus 1+4 Ab|Equine herpesvirus 1+4 Ab
C0880547|T201|COMP|23091-2|LNC|Equine herpesvirus 1+4 Ag|Equine herpesvirus 1+4 Ag
C0880548|T201|COMP|23092-0|LNC|Equine herpesvirus 4 Ag|Equine herpesvirus 4 Ag
C0880549|T201|COMP|23093-8|LNC|Equine herpesvirus 4 DNA|Equine herpesvirus 4 DNA
C0880550|T201|COMP|23094-6|LNC|Equine herpesvirus 4 DNA|Equine herpesvirus 4 DNA
C0880551|T201|COMP|23095-3|LNC|Equine herpesvirus 4 DNA|Equine herpesvirus 4 DNA
C0880552|T201|COMP|23096-1|LNC|Equine infectious anemia virus Ab|Equine infectious anemia virus Ab
C0880553|T201|COMP|23097-9|LNC|Equine infectious anemia virus Ab|Equine infectious anemia virus Ab
C0880554|T201|COMP|23098-7|LNC|Equine infectious anemia virus Ag|Equine infectious anemia virus Ag
C0880555|T201|COMP|23099-5|LNC|Equine infectious anemia virus Ag|Equine infectious anemia virus Ag
C0880556|T201|COMP|23100-1|LNC|Equine influenza virus A1 Ab|Equine influenza virus A1 Ab
C0880557|T201|COMP|23101-9|LNC|Equine influenza virus A1 Ab|Equine influenza virus A1 Ab
C0880558|T201|COMP|23103-5|LNC|Equine influenza virus A2 Ab|Equine influenza virus A2 Ab
C0880559|T201|COMP|23104-3|LNC|Equine influenza virus A2 Ag|Equine influenza virus A2 Ag
C0880560|T201|COMP|23106-8|LNC|Foot and mouth disease virus Ab|Foot and mouth disease virus Ab
C0880561|T201|COMP|23107-6|LNC|Foot and mouth disease virus Ab|Foot and mouth disease virus Ab
C0880562|T201|COMP|23108-4|LNC|Foot and mouth disease virus Ab|Foot and mouth disease virus Ab
C0880563|T201|COMP|23109-2|LNC|Foot and mouth disease virus Ab|Foot and mouth disease virus Ab
C0880564|T201|COMP|23110-0|LNC|Foot and mouth disease virus Ag|Foot and mouth disease virus Ag
C0880565|T201|COMP|23111-8|LNC|Foot and mouth disease virus Ag|Foot and mouth disease virus Ag
C0880566|T201|COMP|23112-6|LNC|Foot and mouth disease virus Ag|Foot and mouth disease virus Ag
C0880567|T201|COMP|23113-4|LNC|Foot and mouth disease virus Ag|Foot and mouth disease virus Ag
C0880568|T201|COMP|23115-9|LNC|Foot and mouth disease virus serotype|Foot and mouth disease virus serotype
C0880569|T201|COMP|23116-7|LNC|Foot and mouth disease virus serotype|Foot and mouth disease virus serotype
C0880570|T201|COMP|23117-5|LNC|Foot and mouth disease virus serotype|Foot and mouth disease virus serotype
C0880571|T201|COMP|23118-3|LNC|Foot and mouth disease virus serotype|Foot and mouth disease virus serotype
C0880572|T201|COMP|23119-1|LNC|Foot and mouth disease virus serotype|Foot and mouth disease virus serotype
C0880573|T201|COMP|23120-9|LNC|Foot and mouth disease virus serotype|Foot and mouth disease virus serotype
C0880574|T201|COMP|23121-7|LNC|Foot and mouth disease virus serotype|Foot and mouth disease virus serotype
C0880575|T201|COMP|23122-5|LNC|Francisella tularensis A DNA|Francisella tularensis A DNA
C0880576|T201|COMP|23124-1|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C0880577|T201|COMP|23125-8|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C0880578|T201|COMP|23126-6|LNC|Francisella tularensis Ag|Francisella tularensis Ag
C0880579|T201|COMP|23127-4|LNC|Francisella tularensis Ag|Francisella tularensis Ag
C0880580|T201|COMP|23128-2|LNC|Francisella tularensis B DNA|Francisella tularensis B DNA
C0880581|T201|COMP|23129-0|LNC|Francisella tularensis B rRNA|Francisella tularensis B rRNA
C0880582|T201|COMP|23130-8|LNC|Francisella tularensis DNA|Francisella tularensis DNA
C0880583|T201|COMP|23131-6|LNC|Francisella tularensis rRNA|Francisella tularensis rRNA
C0880584|T201|COMP|23132-4|LNC|Histoplasma capsulatum farciminosum Ab|Histoplasma capsulatum farciminosum Ab
C0880585|T201|COMP|23133-2|LNC|Histoplasma capsulatum farciminosum Ab|Histoplasma capsulatum farciminosum Ab
C0880586|T201|COMP|23134-0|LNC|Histoplasma capsulatum farciminosum Ab|Histoplasma capsulatum farciminosum Ab
C0880587|T201|COMP|23135-7|LNC|Histoplasma capsulatum farciminosum Ab|Histoplasma capsulatum farciminosum Ab
C0880590|T201|COMP|23139-9|LNC|Infectious bursal disease virus Ab|Infectious bursal disease virus Ab
C0880591|T201|COMP|23140-7|LNC|Infectious bursal disease virus Ab|Infectious bursal disease virus Ab
C0880592|T201|COMP|23141-5|LNC|Infectious bursal disease virus Ab|Infectious bursal disease virus Ab
C0880593|T201|COMP|23142-3|LNC|Infectious bursal disease virus Ag|Infectious bursal disease virus Ag
C0880594|T201|COMP|23143-1|LNC|Infectious bursal disease virus Ag|Infectious bursal disease virus Ag
C0880595|T201|COMP|23144-9|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0880596|T201|COMP|23145-6|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0880597|T201|COMP|23146-4|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0880598|T201|COMP|23147-2|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C0880599|T201|COMP|23148-0|LNC|Japanese encephalitis virus Ag|Japanese encephalitis virus Ag
C0880600|T201|COMP|23149-8|LNC|Japanese encephalitis virus Ag|Japanese encephalitis virus Ag
C0880601|T201|COMP|23150-6|LNC|Leishmania donovani Ag|Leishmania donovani Ag
C0880603|T201|COMP|23152-2|LNC|Leishmania sp Ab|Leishmania sp Ab
C0880604|T201|COMP|23153-0|LNC|Leishmania sp Ab|Leishmania sp Ab
C0880605|T201|COMP|23154-8|LNC|Leishmania sp Ab|Leishmania sp Ab
C0880606|T201|COMP|23155-5|LNC|Leishmania sp Ab|Leishmania sp Ab
C0880607|T201|COMP|23156-3|LNC|Leishmania sp Ab|Leishmania sp Ab
C0880608|T201|COMP|23157-1|LNC|Leishmania sp Ab|Leishmania sp Ab
C0880609|T201|COMP|23158-9|LNC|Leishmania sp rRNA|Leishmania sp rRNA
C0880610|T201|COMP|23159-7|LNC|Leishmania sp DNA|Leishmania sp DNA
C0880611|T201|COMP|23160-5|LNC|Leishmania sp identified|Leishmania sp identified
C0880612|T201|COMP|23161-3|LNC|Leishmania sp identified|Leishmania sp identified
C0880613|T201|COMP|23162-1|LNC|Leishmania sp identified|Leishmania sp identified
C0880614|T201|COMP|23164-7|LNC|Leptospira interrogans serovar Australis Ab|Leptospira interrogans serovar Australis Ab
C0880615|T201|COMP|23165-4|LNC|Leptospira interrogans serovar Autumnalis Ab|Leptospira interrogans serovar Autumnalis Ab
C0880616|T201|COMP|23166-2|LNC|Leptospira interrogans serovar Autumnalis Ab|Leptospira interrogans serovar Autumnalis Ab
C0880617|T201|COMP|23167-0|LNC|Leptospira borgpetersenii serovar Ballum Ab|Leptospira borgpetersenii serovar Ballum Ab
C0880618|T201|COMP|23168-8|LNC|Leptospira borgpetersenii serovar Ballum Ab|Leptospira borgpetersenii serovar Ballum Ab
C0880619|T201|COMP|23170-4|LNC|Leptospira interrogans serovar Bataviae Ab|Leptospira interrogans serovar Bataviae Ab
C0880620|T201|COMP|23171-2|LNC|Leptospira interrogans serovar Bratislava Ab|Leptospira interrogans serovar Bratislava Ab
C0880621|T201|COMP|23173-8|LNC|Leptospira interrogans serovar Canicola Ab|Leptospira interrogans serovar Canicola Ab
C0880622|T201|COMP|23175-3|LNC|Leptospira interrogans serovar Copenhageni Ab|Leptospira interrogans serovar Copenhageni Ab
C0880623|T201|COMP|23176-1|LNC|Leptospira interrogans serovar Copenhageni Ab|Leptospira interrogans serovar Copenhageni Ab
C0880624|T201|COMP|23177-9|LNC|Leptospira interrogans serovar Grippotyphosa Ab|Leptospira interrogans serovar Grippotyphosa Ab
C0880625|T201|COMP|23178-7|LNC|Leptospira interrogans serovar Grippotyphosa Ab|Leptospira interrogans serovar Grippotyphosa Ab
C0880626|T201|COMP|23179-5|LNC|Leptospira interrogans serovar Hardjo Ab|Leptospira interrogans serovar Hardjo Ab
C0880627|T201|COMP|23180-3|LNC|Leptospira interrogans serovar Hardjo Ab|Leptospira interrogans serovar Hardjo Ab
C0880628|T201|COMP|23181-1|LNC|Leptospira interrogans serovar Hardjo Ab|Leptospira interrogans serovar Hardjo Ab
C0880629|T201|COMP|23182-9|LNC|Leptospira interrogans serovar Hebdomadis Ab|Leptospira interrogans serovar Hebdomadis Ab
C0880630|T201|COMP|23183-7|LNC|Leptospira interrogans serovar Hebdomadis Ab|Leptospira interrogans serovar Hebdomadis Ab
C0880633|T201|COMP|23186-0|LNC|Leptospira interrogans Ab|Leptospira interrogans Ab
C0880634|T201|COMP|23187-8|LNC|Leptospira interrogans Ab|Leptospira interrogans Ab
C0880635|T201|COMP|23188-6|LNC|Leptospira interrogans Ab|Leptospira interrogans Ab
C0880636|T201|COMP|23189-4|LNC|Leptospira interrogans serovar Mitis Ab|Leptospira interrogans serovar Mitis Ab
C0880637|T201|COMP|23190-2|LNC|Leptospira interrogans serovar Mitis Ab|Leptospira interrogans serovar Mitis Ab
C0880638|T201|COMP|23191-0|LNC|Leptospira interrogans serovar Pomona Ab|Leptospira interrogans serovar Pomona Ab
C0880639|T201|COMP|23192-8|LNC|Leptospira interrogans serovar Pomona Ab|Leptospira interrogans serovar Pomona Ab
C0880640|T201|COMP|23193-6|LNC|Leptospira borgpetersenii serovar Sejroe Ab|Leptospira borgpetersenii serovar Sejroe Ab
C0880641|T201|COMP|23194-4|LNC|Leptospira borgpetersenii serovar Sejroe Ab|Leptospira borgpetersenii serovar Sejroe Ab
C0880642|T201|COMP|23195-1|LNC|Leptospira sp Ab|Leptospira sp Ab
C0880643|T201|COMP|23196-9|LNC|Leptospira sp Ab|Leptospira sp Ab
C0880644|T201|COMP|23197-7|LNC|Leptospira sp Ab|Leptospira sp Ab
C0880645|T201|COMP|23198-5|LNC|Leptospira sp Ab|Leptospira sp Ab
C0880646|T201|COMP|23199-3|LNC|Leptospira sp Ab.IgG|Leptospira sp Ab.IgG
C0880647|T201|COMP|23200-9|LNC|Leptospira sp Ab.IgG|Leptospira sp Ab.IgG
C0880648|T201|COMP|23201-7|LNC|Leptospira sp Ab.IgM|Leptospira sp Ab.IgM
C0880649|T201|COMP|23202-5|LNC|Leptospira sp Ab.IgM|Leptospira sp Ab.IgM
C0880650|T201|COMP|23203-3|LNC|Leptospira sp Ag|Leptospira sp Ag
C0880651|T201|COMP|23204-1|LNC|Leptospira sp Ag|Leptospira sp Ag
C0880652|T201|COMP|23205-8|LNC|Leptospira sp DNA|Leptospira sp DNA
C0880653|T201|COMP|23206-6|LNC|Leptospira sp DNA|Leptospira sp DNA
C0880654|T201|COMP|23207-4|LNC|Leptospira sp subtype|Leptospira sp subtype
C0880655|T201|COMP|23208-2|LNC|Leptospira borgpetersenii serovar Tarrasovi Ab|Leptospira borgpetersenii serovar Tarrasovi Ab
C0880656|T201|COMP|23209-0|LNC|Leptospira borgpetersenii serovar Tarrasovi Ab|Leptospira borgpetersenii serovar Tarrasovi Ab
C0880657|T201|COMP|23210-8|LNC|Listeria sp Ab|Listeria sp Ab
C0880658|T201|COMP|23211-6|LNC|Listeria sp Ab|Listeria sp Ab
C0880659|T201|COMP|23212-4|LNC|Lumpy skin disease virus|Lumpy skin disease virus
C0880660|T201|COMP|23213-2|LNC|Lumpy skin disease virus Ab|Lumpy skin disease virus Ab
C0880661|T201|COMP|23215-7|LNC|Lumpy skin disease virus Ab|Lumpy skin disease virus Ab
C0880662|T201|COMP|23216-5|LNC|Lumpy skin disease virus Ab|Lumpy skin disease virus Ab
C0880663|T201|COMP|23217-3|LNC|Lumpy skin disease virus Ab|Lumpy skin disease virus Ab
C0880664|T201|COMP|23218-1|LNC|Lumpy skin disease virus Ag|Lumpy skin disease virus Ag
C0880665|T201|COMP|23220-7|LNC|Lumpy skin disease virus Ag|Lumpy skin disease virus Ag
C0880666|T201|COMP|23221-5|LNC|Lumpy skin disease virus Ag|Lumpy skin disease virus Ag
C0880667|T201|COMP|23222-3|LNC|Lumpy skin disease virus Ag|Lumpy skin disease virus Ag
C0880668|T201|COMP|23223-1|LNC|Lumpy skin disease virus DNA|Lumpy skin disease virus DNA
C0880669|T201|COMP|23225-6|LNC|Mareks disease virus Ab|Mareks disease virus Ab
C0880670|T201|COMP|23226-4|LNC|Mareks disease virus Ab|Mareks disease virus Ab
C0880671|T201|COMP|23229-8|LNC|Mareks disease virus Ag|Mareks disease virus Ag
C0880672|T201|COMP|23230-6|LNC|Mareks disease virus Ag|Mareks disease virus Ag
C0880673|T201|COMP|23231-4|LNC|Mareks disease virus DNA|Mareks disease virus DNA
C0880674|T201|COMP|23232-2|LNC|Mite identified|Mite identified
C0880675|T201|COMP|23234-8|LNC|Mycobacterium avium subspecies avium Ab|Mycobacterium avium subspecies avium Ab
C0880676|T201|COMP|23235-5|LNC|Mycobacterium avium subspecies avium Ab|Mycobacterium avium subspecies avium Ab
C0880677|T201|COMP|23236-3|LNC|Mycobacterium avium subspecies avium rRNA|Mycobacterium avium subspecies avium rRNA
C0880678|T201|COMP|23237-1|LNC|Mycobacterium avium subspecies avium identified|Mycobacterium avium subspecies avium identified
C0880679|T201|COMP|23239-7|LNC|Mycobacterium bovis Ab|Mycobacterium bovis Ab
C0880680|T201|COMP|23240-5|LNC|Mycobacterium bovis Ab|Mycobacterium bovis Ab
C0880681|T201|COMP|23241-3|LNC|Mycobacterium bovis Ag|Mycobacterium bovis Ag
C0880682|T201|COMP|23242-1|LNC|Mycobacterium bovis Ag|Mycobacterium bovis Ag
C0880683|T201|COMP|23243-9|LNC|Mycobacterium avium subspecies paratuberculosis|Mycobacterium avium subspecies paratuberculosis
C0880684|T201|COMP|23244-7|LNC|Mycobacterium avium subspecies paratuberculosis|Mycobacterium avium subspecies paratuberculosis
C0880687|T201|COMP|23247-0|LNC|Mycobacterium sp DNA|Mycobacterium sp DNA
C0880688|T201|COMP|23248-8|LNC|Mycoplasma agalactiae Ab|Mycoplasma agalactiae Ab
C0880689|T201|COMP|23249-6|LNC|Mycoplasma agalactiae Ab|Mycoplasma agalactiae Ab
C0880690|T201|COMP|23250-4|LNC|Mycoplasma agalactiae Ab|Mycoplasma agalactiae Ab
C0880691|T201|COMP|23251-2|LNC|Mycoplasma agalactiae Ab|Mycoplasma agalactiae Ab
C0880692|T201|COMP|23252-0|LNC|Mycoplasma agalactiae DNA|Mycoplasma agalactiae DNA
C0880693|T201|COMP|23253-8|LNC|Mycoplasma arginini Ab|Mycoplasma arginini Ab
C0880694|T201|COMP|23254-6|LNC|Mycoplasma arginini Ab|Mycoplasma arginini Ab
C0880695|T201|COMP|23256-1|LNC|Mycoplasma bovis Ab|Mycoplasma bovis Ab
C0880696|T201|COMP|23257-9|LNC|Mycoplasma capricolum subspecies capricolum Ab|Mycoplasma capricolum subspecies capricolum Ab
C0880697|T201|COMP|23258-7|LNC|Mycoplasma capricolum subspecies capricolum Ab|Mycoplasma capricolum subspecies capricolum Ab
C0880698|T201|COMP|23259-5|LNC|Mycoplasma capricolum subspecies capricolum Ab|Mycoplasma capricolum subspecies capricolum Ab
C0880711|T201|COMP|23273-6|LNC|Mycoplasma gallisepticum Ab|Mycoplasma gallisepticum Ab
C0880712|T201|COMP|23275-1|LNC|Mycoplasma gallisepticum Ab|Mycoplasma gallisepticum Ab
C0880713|T201|COMP|23276-9|LNC|Mycoplasma gallisepticum Ag|Mycoplasma gallisepticum Ag
C0880714|T201|COMP|23277-7|LNC|Mycoplasma gallisepticum Ag|Mycoplasma gallisepticum Ag
C0880715|T201|COMP|23278-5|LNC|Mycoplasma gallisepticum Ag|Mycoplasma gallisepticum Ag
C0880716|T201|COMP|23279-3|LNC|Mycoplasma gallisepticum DNA|Mycoplasma gallisepticum DNA
C0880717|T201|COMP|23280-1|LNC|Mycoplasma meleagridis Ab|Mycoplasma meleagridis Ab
C0880718|T201|COMP|23281-9|LNC|Mycoplasma mycoides subspecies capri Ab|Mycoplasma mycoides subspecies capri Ab
C0880719|T201|COMP|23282-7|LNC|Mycoplasma mycoides subspecies capri Ab|Mycoplasma mycoides subspecies capri Ab
C0880729|T201|COMP|23294-2|LNC|Mycoplasma putrefaciens Ab|Mycoplasma putrefaciens Ab
C0880730|T201|COMP|23295-9|LNC|Mycoplasma putrefaciens Ab|Mycoplasma putrefaciens Ab
C0880731|T201|COMP|23296-7|LNC|Mycoplasma putrefaciens Ab|Mycoplasma putrefaciens Ab
C0880732|T201|COMP|23297-5|LNC|Mycoplasma sp Ab|Mycoplasma sp Ab
C0880733|T201|COMP|23298-3|LNC|Mycoplasma sp Ag|Mycoplasma sp Ag
C0880734|T201|COMP|23299-1|LNC|Mycoplasma sp Ag|Mycoplasma sp Ag
C0880735|T201|COMP|23300-7|LNC|Mycoplasma sp rRNA|Mycoplasma sp rRNA
C0880736|T201|COMP|23301-5|LNC|Mycoplasma sp DNA|Mycoplasma sp DNA
C0880737|T201|COMP|23302-3|LNC|Mycoplasma synoviae Ab|Mycoplasma synoviae Ab
C0880738|T201|COMP|23303-1|LNC|Myxoma virus Ab|Myxoma virus Ab
C0880739|T201|COMP|23304-9|LNC|Myxoma virus Ab|Myxoma virus Ab
C0880740|T201|COMP|23305-6|LNC|Myxoma virus Ab|Myxoma virus Ab
C0880741|T201|COMP|23306-4|LNC|Myxoma virus Ab|Myxoma virus Ab
C0880742|T201|COMP|23307-2|LNC|Myxoma virus Ab|Myxoma virus Ab
C0880743|T201|COMP|23308-0|LNC|Myxoma virus Ab|Myxoma virus Ab
C0880744|T201|COMP|23309-8|LNC|Myxoma virus Ab|Myxoma virus Ab
C0880745|T201|COMP|23310-6|LNC|Myxoma virus Ag|Myxoma virus Ag
C0880746|T201|COMP|23311-4|LNC|Myxoma virus Ag|Myxoma virus Ag
C0880747|T201|COMP|23316-3|LNC|Nairobi sheep disease virus Ab|Nairobi sheep disease virus Ab
C0880748|T201|COMP|23313-0|LNC|Nairobi sheep disease virus Ab|Nairobi sheep disease virus Ab
C0880749|T201|COMP|23314-8|LNC|Nairobi sheep disease virus Ab|Nairobi sheep disease virus Ab
C0880750|T201|COMP|23315-5|LNC|Nairobi sheep disease virus Ab|Nairobi sheep disease virus Ab
C0880751|T201|COMP|23318-9|LNC|Nairobi sheep disease virus Ag|Nairobi sheep disease virus Ag
C0880752|T201|COMP|23319-7|LNC|Nairobi sheep disease virus Ag|Nairobi sheep disease virus Ag
C0880753|T201|COMP|23320-5|LNC|Nairobi sheep disease virus Ag|Nairobi sheep disease virus Ag
C0880754|T201|COMP|23322-1|LNC|Ovine herpesvirus 2 Ab|Ovine herpesvirus 2 Ab
C0880755|T201|COMP|23324-7|LNC|Ovine herpesvirus 2 Ab|Ovine herpesvirus 2 Ab
C0880756|T201|COMP|23325-4|LNC|Ovine herpesvirus 2 Ab|Ovine herpesvirus 2 Ab
C0880757|T201|COMP|23326-2|LNC|Ovine herpesvirus 2 Ab|Ovine herpesvirus 2 Ab
C0880758|T201|COMP|23327-0|LNC|Ovine herpesvirus 2 DNA|Ovine herpesvirus 2 DNA
C0880759|T201|COMP|23330-4|LNC|Ovine progressive pneumonia virus Ab|Ovine progressive pneumonia virus Ab
C0880760|T201|COMP|23329-6|LNC|Ovine progressive pneumonia virus Ab|Ovine progressive pneumonia virus Ab
C0880761|T201|COMP|23332-0|LNC|Ovine progressive pneumonia virus Ab|Ovine progressive pneumonia virus Ab
C0880762|T201|COMP|23334-6|LNC|Ovine progressive pneumonia virus Ag|Ovine progressive pneumonia virus Ag
C0880763|T201|COMP|23335-3|LNC|Ovine progressive pneumonia virus Ag|Ovine progressive pneumonia virus Ag
C0880764|T201|COMP|23336-1|LNC|Ovine progressive pneumonia virus DNA|Ovine progressive pneumonia virus DNA
C0880765|T201|COMP|23337-9|LNC|Ovine progressive pneumonia virus DNA|Ovine progressive pneumonia virus DNA
C0880768|T201|COMP|23341-1|LNC|Pasteurella multocida Ab|Pasteurella multocida Ab
C0880769|T201|COMP|23342-9|LNC|Pasteurella multocida Ab|Pasteurella multocida Ab
C0880770|T201|COMP|23343-7|LNC|Pasteurella multocida Ag|Pasteurella multocida Ag
C0880771|T201|COMP|23346-0|LNC|Pasteurella multocida serotype|Pasteurella multocida serotype
C0880772|T201|COMP|23347-8|LNC|Pasteurella multocida serotype|Pasteurella multocida serotype
C0880773|T201|COMP|23345-2|LNC|Pasteurella multocida serotype|Pasteurella multocida serotype
C0880774|T201|COMP|23350-2|LNC|Peste des petits ruminants virus Ab|Peste des petits ruminants virus Ab
C0880775|T201|COMP|23352-8|LNC|Peste des petits ruminants virus Ab|Peste des petits ruminants virus Ab
C0880776|T201|COMP|23351-0|LNC|Peste des petits ruminants virus Ab|Peste des petits ruminants virus Ab
C0880777|T201|COMP|23354-4|LNC|Peste des petits ruminants virus Ab|Peste des petits ruminants virus Ab
C0880778|T201|COMP|23355-1|LNC|Peste des petits ruminants virus Ag|Peste des petits ruminants virus Ag
C0880779|T201|COMP|23356-9|LNC|Peste des petits ruminants virus Ag|Peste des petits ruminants virus Ag
C0880780|T201|COMP|23357-7|LNC|Peste des petits ruminants virus Ag|Peste des petits ruminants virus Ag
C0880781|T201|COMP|23358-5|LNC|Peste des petits ruminants virus RNA|Peste des petits ruminants virus RNA
C0880782|T201|COMP|23359-3|LNC|Peste des petits ruminants virus RNA|Peste des petits ruminants virus RNA
C0880783|T201|COMP|23360-1|LNC|Porcine enterovirus Ag|Porcine enterovirus Ag
C0880784|T201|COMP|23361-9|LNC|Porcine enterovirus Ab|Porcine enterovirus Ab
C0880785|T201|COMP|23362-7|LNC|Porcine enterovirus Ab|Porcine enterovirus Ab
C0880786|T201|COMP|23363-5|LNC|Porcine enterovirus Ab|Porcine enterovirus Ab
C0880787|T201|COMP|23364-3|LNC|Porcine enterovirus Ag|Porcine enterovirus Ag
C0880788|T201|COMP|23365-0|LNC|Porcine parvovirus Ab|Porcine parvovirus Ab
C0880789|T201|COMP|23366-8|LNC|Porcine parvovirus Ab|Porcine parvovirus Ab
C0880795|T201|COMP|23372-6|LNC|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C0880796|T201|COMP|23374-2|LNC|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C0880797|T201|COMP|23376-7|LNC|Porcine respiratory coronavirus Ag|Porcine respiratory coronavirus Ag
C0880798|T201|COMP|23377-5|LNC|Porcine respiratory coronavirus Ag|Porcine respiratory coronavirus Ag
C0880799|T201|COMP|23378-3|LNC|Porcine respiratory coronavirus RNA|Porcine respiratory coronavirus RNA
C0880800|T201|COMP|23379-1|LNC|Prion protein.abnormal|Prion protein.abnormal
C0880801|T201|COMP|23380-9|LNC|Prion protein.abnormal|Prion protein.abnormal
C0880802|T201|COMP|23381-7|LNC|Prion protein.abnormal|Prion protein.abnormal
C0880803|T201|COMP|23383-3|LNC|Pseudorabies virus Ag|Pseudorabies virus Ag
C0880804|T201|COMP|23384-1|LNC|Pseudorabies virus Ag|Pseudorabies virus Ag
C0880805|T201|COMP|23385-8|LNC|Pseudorabies virus Ag|Pseudorabies virus Ag
C0880806|T201|COMP|23386-6|LNC|Pseudorabies virus Ag|Pseudorabies virus Ag
C0880807|T201|COMP|23388-2|LNC|Rabies virus|Rabies virus
C0880808|T201|COMP|23389-0|LNC|Rabies virus Ag|Rabies virus Ag
C0880809|T201|COMP|23390-8|LNC|Rabies virus Ag|Rabies virus Ag
C0880810|T201|COMP|23391-6|LNC|Rabies virus Ag|Rabies virus Ag
C0880811|T201|COMP|23393-2|LNC|Rabies virus DNA|Rabies virus DNA
C0880812|T201|COMP|23396-5|LNC|Rift valley fever virus Ab|Rift valley fever virus Ab
C0880813|T201|COMP|23398-1|LNC|Rift valley fever virus Ab|Rift valley fever virus Ab
C0880814|T201|COMP|23399-9|LNC|Rift valley fever virus Ab|Rift valley fever virus Ab
C0880815|T201|COMP|23401-3|LNC|Rift valley fever virus Ag|Rift valley fever virus Ag
C0880816|T201|COMP|23402-1|LNC|Rift valley fever virus Ag|Rift valley fever virus Ag
C0880817|T201|COMP|23403-9|LNC|Rift valley fever virus Ag|Rift valley fever virus Ag
C0880818|T201|COMP|23404-7|LNC|Rift valley fever virus Ag|Rift valley fever virus Ag
C0880819|T201|COMP|23406-2|LNC|Rift valley fever virus Ag|Rift valley fever virus Ag
C0880820|T201|COMP|23407-0|LNC|Rinderpest virus Ab|Rinderpest virus Ab
C0880821|T201|COMP|23408-8|LNC|Rinderpest virus Ab|Rinderpest virus Ab
C0880822|T201|COMP|23409-6|LNC|Rinderpest virus Ab|Rinderpest virus Ab
C0880823|T201|COMP|23410-4|LNC|Rinderpest virus Ab|Rinderpest virus Ab
C0880824|T201|COMP|23411-2|LNC|Rinderpest virus Ab|Rinderpest virus Ab
C0880825|T201|COMP|23412-0|LNC|Rinderpest virus Ag|Rinderpest virus Ag
C0880826|T201|COMP|23413-8|LNC|Rinderpest virus Ag|Rinderpest virus Ag
C0880827|T201|COMP|23414-6|LNC|Rinderpest virus Ag|Rinderpest virus Ag
C0880828|T201|COMP|23415-3|LNC|Rinderpest virus Ag|Rinderpest virus Ag
C0880829|T201|COMP|23416-1|LNC|Rinderpest virus Ag|Rinderpest virus Ag
C0880830|T201|COMP|23417-9|LNC|Rinderpest virus RNA|Rinderpest virus RNA
C0880831|T201|COMP|23418-7|LNC|Salmonella abortus equi Ab|Salmonella abortus equi Ab
C0880832|T201|COMP|23419-5|LNC|Salmonella abortus equi Ab|Salmonella abortus equi Ab
C0880833|T201|COMP|23421-1|LNC|Salmonella abortus ovis Ab|Salmonella abortus ovis Ab
C0880834|T201|COMP|23422-9|LNC|Salmonella enteritidis Ab.IgG|Salmonella enteritidis Ab.IgG
C0880835|T201|COMP|23423-7|LNC|Salmonella enteritidis Ab.IgG|Salmonella enteritidis Ab.IgG
C0880836|T201|COMP|23424-5|LNC|Salmonella enteritidis Ab.IgG|Salmonella enteritidis Ab.IgG
C0880837|T201|COMP|23425-2|LNC|Salmonella enteritidis Ab.IgG|Salmonella enteritidis Ab.IgG
C0880838|T201|COMP|23426-0|LNC|Salmonella gallinarum Ab|Salmonella gallinarum Ab
C0880839|T201|COMP|23427-8|LNC|Salmonella gallinarum Ab|Salmonella gallinarum Ab
C0880840|T201|COMP|23428-6|LNC|Salmonella gallinarum Ab|Salmonella gallinarum Ab
C0880841|T201|COMP|23429-4|LNC|Salmonella gallinarum Ab|Salmonella gallinarum Ab
C0880842|T201|COMP|23431-0|LNC|Salmonella gallinarum DNA|Salmonella gallinarum DNA
C0880843|T201|COMP|23432-8|LNC|Salmonella gallinarum rRNA|Salmonella gallinarum rRNA
C0880844|T201|COMP|23433-6|LNC|Salmonella pullorum Ab|Salmonella pullorum Ab
C0880845|T201|COMP|23434-4|LNC|Salmonella pullorum Ab|Salmonella pullorum Ab
C0880846|T201|COMP|23435-1|LNC|Salmonella pullorum DNA|Salmonella pullorum DNA
C0880847|T201|COMP|23436-9|LNC|Salmonella pullorum rRNA|Salmonella pullorum rRNA
C0880848|T201|COMP|23437-7|LNC|Swine influenza virus Ab|Swine influenza virus Ab
C0880849|T201|COMP|23438-5|LNC|Swine influenza virus Ab|Swine influenza virus Ab
C0880850|T201|COMP|23440-1|LNC|Swine vesicular disease virus Ab|Swine vesicular disease virus Ab
C0880851|T201|COMP|23441-9|LNC|Swine vesicular disease virus Ab|Swine vesicular disease virus Ab
C0880852|T201|COMP|23442-7|LNC|Swine vesicular disease virus Ab|Swine vesicular disease virus Ab
C0880853|T201|COMP|23444-3|LNC|Swine vesicular disease virus Ag|Swine vesicular disease virus Ag
C0880854|T201|COMP|23445-0|LNC|Swine vesicular disease virus Ag|Swine vesicular disease virus Ag
C0880855|T201|COMP|23446-8|LNC|Swine vesicular disease virus Ag|Swine vesicular disease virus Ag
C0880856|T201|COMP|23447-6|LNC|Swine vesicular disease virus Ag|Swine vesicular disease virus Ag
C0880857|T201|COMP|23448-4|LNC|Swine vesicular disease virus RNA|Swine vesicular disease virus RNA
C0880858|T201|COMP|23450-0|LNC|Taenia sp Ag|Taenia sp Ag
C0880859|T201|COMP|23451-8|LNC|Taenia sp eggs|Taenia sp eggs
C0880860|T201|COMP|23454-2|LNC|Taylorella equigenitalis Ab|Taylorella equigenitalis Ab
C0880861|T201|COMP|23455-9|LNC|Taylorella equigenitalis Ag|Taylorella equigenitalis Ag
C0880862|T201|COMP|23456-7|LNC|Taylorella equigenitalis Ag|Taylorella equigenitalis Ag
C0880863|T201|COMP|23459-1|LNC|Theileria annulata Ab|Theileria annulata Ab
C0880864|T201|COMP|23460-9|LNC|Theileria annulata Ab|Theileria annulata Ab
C0880865|T201|COMP|23461-7|LNC|Theileria annulata Ab|Theileria annulata Ab
C0880866|T201|COMP|23462-5|LNC|Theileria annulata Ab|Theileria annulata Ab
C0880867|T201|COMP|23464-1|LNC|Theileria equi Ab|Theileria equi Ab
C0880868|T201|COMP|23465-8|LNC|Theileria equi rRNA|Theileria equi rRNA
C0880869|T201|COMP|23466-6|LNC|Theileria equi Ab|Theileria equi Ab
C0880870|T201|COMP|23467-4|LNC|Theileria mutans Ab|Theileria mutans Ab
C0880871|T201|COMP|23468-2|LNC|Theileria mutans Ab|Theileria mutans Ab
C0880872|T201|COMP|23469-0|LNC|Theileria mutans Ab|Theileria mutans Ab
C0880873|T201|COMP|23470-8|LNC|Theileria mutans Ab|Theileria mutans Ab
C0880874|T201|COMP|23471-6|LNC|Theileria mutans Ab|Theileria mutans Ab
C0880875|T201|COMP|23472-4|LNC|Theileria mutans rRNA|Theileria mutans rRNA
C0880876|T201|COMP|23473-2|LNC|Theileria mutans DNA|Theileria mutans DNA
C0880877|T201|COMP|23474-0|LNC|Theileria parva Ab|Theileria parva Ab
C0880878|T201|COMP|23475-7|LNC|Theileria parva Ab|Theileria parva Ab
C0880879|T201|COMP|23476-5|LNC|Theileria parva Ab|Theileria parva Ab
C0880880|T201|COMP|23477-3|LNC|Theileria parva Ab|Theileria parva Ab
C0880881|T201|COMP|23478-1|LNC|Theileria parva Ab|Theileria parva Ab
C0880882|T201|COMP|23479-9|LNC|Theileria parva rRNA|Theileria parva rRNA
C0880883|T201|COMP|23480-7|LNC|Theileria parva DNA|Theileria parva DNA
C0880884|T201|COMP|23481-5|LNC|Theileria parva rRNA|Theileria parva rRNA
C0880885|T201|COMP|23482-3|LNC|Theileria sp|Theileria sp
C0880886|T201|COMP|23483-1|LNC|Theileria sp|Theileria sp
C0880887|T201|COMP|23484-9|LNC|Toxoplasma sp Ab|Toxoplasma sp Ab
C0880888|T201|COMP|23485-6|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C0880889|T201|COMP|23486-4|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C0880890|T201|COMP|23488-0|LNC|Transmissible gastroenteritis virus Ab|Transmissible gastroenteritis virus Ab
C0880891|T201|COMP|23489-8|LNC|Transmissible gastroenteritis virus Ab|Transmissible gastroenteritis virus Ab
C0880892|T201|COMP|23487-2|LNC|Transmissible gastroenteritis virus Ab|Transmissible gastroenteritis virus Ab
C0880893|T201|COMP|23492-2|LNC|Transmissible gastroenteritis virus Ab|Transmissible gastroenteritis virus Ab
C0880894|T201|COMP|23493-0|LNC|Transmissible gastroenteritis virus Ag|Transmissible gastroenteritis virus Ag
C0880895|T201|COMP|23494-8|LNC|Transmissible gastroenteritis virus Ag|Transmissible gastroenteritis virus Ag
C0880896|T201|COMP|23495-5|LNC|Transmissible gastroenteritis virus Ag|Transmissible gastroenteritis virus Ag
C0880897|T201|COMP|23497-1|LNC|Transmissible gastroenteritis virus Ag|Transmissible gastroenteritis virus Ag
C0880898|T201|COMP|23498-9|LNC|Transmissible gastroenteritis virus RNA|Transmissible gastroenteritis virus RNA
C0880899|T201|COMP|23499-7|LNC|Trichinella spiralis|Trichinella spiralis
C0880900|T201|COMP|23501-0|LNC|Tritrichomonas foetus Ab|Tritrichomonas foetus Ab
C0880901|T201|COMP|23502-8|LNC|Tritrichomonas foetus Ag|Tritrichomonas foetus Ag
C0880902|T201|COMP|23503-6|LNC|Tritrichomonas foetus Ag|Tritrichomonas foetus Ag
C0880903|T201|COMP|23504-4|LNC|Tritrichomonas foetus DNA|Tritrichomonas foetus DNA
C0880905|T201|COMP|23507-7|LNC|Trypanosoma brucei DNA|Trypanosoma brucei DNA
C0880906|T201|COMP|23508-5|LNC|Trypanosoma congolense DNA|Trypanosoma congolense DNA
C0880907|T201|COMP|23509-3|LNC|Trypanosoma equiperdum|Trypanosoma equiperdum
C0880908|T201|COMP|23511-9|LNC|Trypanosoma equiperdum Ab|Trypanosoma equiperdum Ab
C0880909|T201|COMP|23512-7|LNC|Trypanosoma equiperdum Ab|Trypanosoma equiperdum Ab
C0880910|T201|COMP|23513-5|LNC|Trypanosoma equiperdum Ab|Trypanosoma equiperdum Ab
C0880911|T201|COMP|23514-3|LNC|Trypanosoma equiperdum Ab|Trypanosoma equiperdum Ab
C0880913|T201|COMP|23517-6|LNC|Trypanosoma equiperdum Ab|Trypanosoma equiperdum Ab
C0880914|T201|COMP|23518-4|LNC|Trypanosoma evansi|Trypanosoma evansi
C0880915|T201|COMP|23519-2|LNC|Trypanosoma evansi|Trypanosoma evansi
C0880916|T201|COMP|23520-0|LNC|Trypanosoma evansi|Trypanosoma evansi
C0880917|T201|COMP|23521-8|LNC|Trypanosoma evansi Ab|Trypanosoma evansi Ab
C0880918|T201|COMP|23523-4|LNC|Trypanosoma evansi Ab|Trypanosoma evansi Ab
C0880919|T201|COMP|23522-6|LNC|Trypanosoma evansi Ab|Trypanosoma evansi Ab
C0880920|T201|COMP|23526-7|LNC|Trypanosoma evansi Ab|Trypanosoma evansi Ab
C0880921|T201|COMP|23527-5|LNC|Trypanosoma evansi Ag|Trypanosoma evansi Ag
C0880922|T201|COMP|23528-3|LNC|Trypanosoma evansi Ag|Trypanosoma evansi Ag
C0880923|T201|COMP|23529-1|LNC|Trypanosoma evansi DNA|Trypanosoma evansi DNA
C0880924|T201|COMP|23530-9|LNC|Trypanosoma evansi rRNA|Trypanosoma evansi rRNA
C0880925|T201|COMP|23531-7|LNC|Trypanosoma sp Ab|Trypanosoma sp Ab
C0880926|T201|COMP|23532-5|LNC|Trypanosoma sp Ab|Trypanosoma sp Ab
C0880927|T201|COMP|23533-3|LNC|Trypanosoma sp Ab|Trypanosoma sp Ab
C0880928|T201|COMP|23534-1|LNC|Trypanosoma sp Ab|Trypanosoma sp Ab
C0880929|T201|COMP|23535-8|LNC|Trypanosoma sp Ag|Trypanosoma sp Ag
C0880930|T201|COMP|23536-6|LNC|Trypanosoma sp identified|Trypanosoma sp identified
C0880934|T201|COMP|23540-8|LNC|Turkey enteritis coronavirus|Turkey enteritis coronavirus
C0880935|T201|COMP|23541-6|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C0880936|T201|COMP|23542-4|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C0880937|T201|COMP|23543-2|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C0880938|T201|COMP|23544-0|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C0880939|T201|COMP|23545-7|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C0880940|T201|COMP|23546-5|LNC|Venezuelan equine encephalitis virus Ab.IgM|Venezuelan equine encephalitis virus Ab.IgM
C0880941|T201|COMP|23547-3|LNC|Venezuelan equine encephalitis virus Ab.IgM|Venezuelan equine encephalitis virus Ab.IgM
C0880942|T201|COMP|23548-1|LNC|Venezuelan equine encephalitis virus Ag|Venezuelan equine encephalitis virus Ag
C0880943|T201|COMP|23549-9|LNC|Venezuelan equine encephalitis virus Ag|Venezuelan equine encephalitis virus Ag
C0880944|T201|COMP|23550-7|LNC|Venezuelan equine encephalitis virus Ag|Venezuelan equine encephalitis virus Ag
C0880945|T201|COMP|23551-5|LNC|Venezuelan equine encephalitis virus Ag|Venezuelan equine encephalitis virus Ag
C0880946|T201|COMP|23552-3|LNC|Venezuelan equine encephalitis virus subtype|Venezuelan equine encephalitis virus subtype
C0880947|T201|COMP|23553-1|LNC|Venezuelan equine encephalitis virus subtype|Venezuelan equine encephalitis virus subtype
C0880948|T201|COMP|23554-9|LNC|Venezuelan equine encephalitis virus subtype|Venezuelan equine encephalitis virus subtype
C0880949|T201|COMP|23555-6|LNC|Vesicular stomatitis virus Ab|Vesicular stomatitis virus Ab
C0880950|T201|COMP|23558-0|LNC|Vesicular stomatitis virus Ag|Vesicular stomatitis virus Ag
C0880951|T201|COMP|23559-8|LNC|Vesicular stomatitis virus Ag|Vesicular stomatitis virus Ag
C0880952|T201|COMP|23560-6|LNC|Vesicular stomatitis virus Ag|Vesicular stomatitis virus Ag
C0880953|T201|COMP|23561-4|LNC|Vesicular stomatitis Indiana virus Ab|Vesicular stomatitis Indiana virus Ab
C0880954|T201|COMP|23563-0|LNC|Vesicular stomatitis Indiana virus Ab|Vesicular stomatitis Indiana virus Ab
C0880955|T201|COMP|23564-8|LNC|Vesicular stomatitis Indiana virus Ab|Vesicular stomatitis Indiana virus Ab
C0880956|T201|COMP|23565-5|LNC|Vesicular stomatitis New Jersey virus Ab|Vesicular stomatitis New Jersey virus Ab
C0880957|T201|COMP|23566-3|LNC|Vesicular stomatitis New Jersey virus Ab|Vesicular stomatitis New Jersey virus Ab
C0880958|T201|COMP|23568-9|LNC|Vesicular stomatitis New Jersey virus Ab|Vesicular stomatitis New Jersey virus Ab
C0880959|T201|COMP|23570-5|LNC|Vesicular stomatitis virus serotype|Vesicular stomatitis virus serotype
C0880960|T201|COMP|23571-3|LNC|Vesicular stomatitis virus serotype|Vesicular stomatitis virus serotype
C0880961|T201|COMP|23573-9|LNC|Viral hemorrhagic disease virus|Viral hemorrhagic disease virus
C0880962|T201|COMP|23574-7|LNC|Viral hemorrhagic disease virus Ab|Viral hemorrhagic disease virus Ab
C0880963|T201|COMP|23575-4|LNC|Viral hemorrhagic disease virus Ab|Viral hemorrhagic disease virus Ab
C0880964|T201|COMP|23576-2|LNC|Viral hemorrhagic disease virus Ab|Viral hemorrhagic disease virus Ab
C0880965|T201|COMP|23577-0|LNC|Viral hemorrhagic disease virus Ab|Viral hemorrhagic disease virus Ab
C0880966|T201|COMP|23579-6|LNC|Viral hemorrhagic disease virus Ag|Viral hemorrhagic disease virus Ag
C0880967|T201|COMP|23580-4|LNC|Viral hemorrhagic disease virus Ag|Viral hemorrhagic disease virus Ag
C0880968|T201|COMP|23581-2|LNC|Viral hemorrhagic disease virus Ag|Viral hemorrhagic disease virus Ag
C0880969|T201|COMP|23582-0|LNC|Viral hemorrhagic disease virus Ag|Viral hemorrhagic disease virus Ag
C0880970|T201|COMP|23583-8|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0880971|T201|COMP|23584-6|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0880972|T201|COMP|23585-3|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0880973|T201|COMP|23586-1|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0880974|T201|COMP|23587-9|LNC|Western equine encephalitis virus Ab.IgM|Western equine encephalitis virus Ab.IgM
C0880975|T201|COMP|23588-7|LNC|Western equine encephalitis virus Ab.IgM|Western equine encephalitis virus Ab.IgM
C0880976|T201|COMP|23589-5|LNC|Western equine encephalitis virus Ag|Western equine encephalitis virus Ag
C0880977|T201|COMP|23590-3|LNC|Western equine encephalitis virus Ag|Western equine encephalitis virus Ag
C0880978|T201|COMP|23591-1|LNC|Western equine encephalitis virus Ag|Western equine encephalitis virus Ag
C0880979|T201|COMP|23592-9|LNC|African swine fever virus Ab|African swine fever virus Ab
C0880980|T201|COMP|23593-7|LNC|Bovine leukemia virus|Bovine leukemia virus
C0880981|T201|COMP|23594-5|LNC|Brucella sp identified|Brucella sp identified
C0880982|T201|COMP|23595-2|LNC|Dermatophilus congolensis|Dermatophilus congolensis
C0880983|T201|COMP|23596-0|LNC|Dermatophilus congolensis|Dermatophilus congolensis
C0880984|T201|COMP|23597-8|LNC|Dermatophilus congolensis|Dermatophilus congolensis
C0880985|T201|COMP|23598-6|LNC|Dermatophilus congolensis Ag|Dermatophilus congolensis Ag
C0880986|T201|COMP|23599-4|LNC|Leptospira sp identified|Leptospira sp identified
C0880987|T201|COMP|23600-0|LNC|Leptospira sp identified|Leptospira sp identified
C0880988|T201|COMP|23601-8|LNC|Mareks disease virus serotype|Mareks disease virus serotype
C0880989|T201|COMP|23602-6|LNC|Salmonella enteritidis|Salmonella enteritidis
C0880990|T201|COMP|23603-4|LNC|Taylorella equigenitalis|Taylorella equigenitalis
C0880991|T201|COMP|23604-2|LNC|Tritrichomonas foetus|Tritrichomonas foetus
C0880992|T201|COMP|23605-9|LNC|Tritrichomonas foetus|Tritrichomonas foetus
C0880993|T201|COMP|23606-7|LNC|Tritrichomonas foetus|Tritrichomonas foetus
C0880994|T201|COMP|23607-5|LNC|Capreomycin|Capreomycin
C0880995|T201|COMP|23608-3|LNC|cycloSERINE|cycloSERINE
C0880996|T201|COMP|23609-1|LNC|Kanamycin|Kanamycin
C0880997|T201|COMP|23610-9|LNC|Sparfloxacin|Sparfloxacin
C0880998|T201|COMP|23612-5|LNC|Azithromycin|Azithromycin
C0880999|T201|COMP|23613-3|LNC|Imipenem|Imipenem
C0881000|T201|COMP|23614-1|LNC|Trimethoprim|Trimethoprim
C0881001|T201|COMP|23615-8|LNC|Vancomycin|Vancomycin
C0881002|T201|COMP|23616-6|LNC|Viomycin|Viomycin
C0881003|T201|COMP|23618-2|LNC|Ampicillin+Sulbactam|Ampicillin+Sulbactam
C0881004|T201|COMP|23619-0|LNC|Clarithromycin|Clarithromycin
C0881005|T201|COMP|23621-6|LNC|Ciprofloxacin|Ciprofloxacin
C0881006|T201|COMP|23622-4|LNC|Ceftizoxime|Ceftizoxime
C0881007|T201|COMP|23623-2|LNC|Doxycycline|Doxycycline
C0881008|T201|COMP|23624-0|LNC|Amikacin|Amikacin
C0881009|T201|COMP|23626-5|LNC|Streptomycin|Streptomycin
C0881010|T201|COMP|23627-3|LNC|Clofazimine|Clofazimine
C0881011|T201|COMP|23628-1|LNC|Sparfloxacin|Sparfloxacin
C0881012|T201|COMP|23629-9|LNC|Para aminosalicylate|Para aminosalicylate
C0881013|T201|COMP|23630-7|LNC|Rifabutin|Rifabutin
C0881014|T201|COMP|23631-5|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0881015|T201|COMP|23632-3|LNC|Pyrazinamide|Pyrazinamide
C0881016|T201|COMP|23634-9|LNC|Erythropoietin given|Erythropoietin given
C0881017|T201|COMP|23636-4|LNC|Cefdinir|Cefdinir
C0881018|T201|COMP|23637-2|LNC|Cefdinir|Cefdinir
C0881019|T201|COMP|23639-8|LNC|Grepafloxacin|Grepafloxacin
C0881020|T201|COMP|23640-6|LNC|Quinupristin+Dalfopristin|Quinupristin+Dalfopristin
C0881021|T201|COMP|23641-4|LNC|Quinupristin+Dalfopristin|Quinupristin+Dalfopristin
C0881022|T201|COMP|23642-2|LNC|Trovafloxacin|Trovafloxacin
C0881023|T201|COMP|23643-0|LNC|Trovafloxacin|Trovafloxacin
C0881024|T201|COMP|23644-8|LNC|Actinobacillus pleuropneumoniae serotype 1 Ab|Actinobacillus pleuropneumoniae serotype 1 Ab
C0881025|T201|COMP|23645-5|LNC|Actinobacillus pleuropneumoniae serotype 3 Ab|Actinobacillus pleuropneumoniae serotype 3 Ab
C0881026|T201|COMP|23646-3|LNC|Actinobacillus pleuropneumoniae serotype 5 Ab|Actinobacillus pleuropneumoniae serotype 5 Ab
C0881027|T201|COMP|23647-1|LNC|Actinobacillus pleuropneumoniae serotype 7 Ab|Actinobacillus pleuropneumoniae serotype 7 Ab
C0881028|T201|COMP|23648-9|LNC|Actinobacillus pleuropneumoniae Ab|Actinobacillus pleuropneumoniae Ab
C0881029|T201|COMP|23650-5|LNC|Actinobacillus pleuropneumoniae serotype|Actinobacillus pleuropneumoniae serotype
C0881030|T201|COMP|23651-3|LNC|Actinobacillus suis serotype|Actinobacillus suis serotype
C0881031|T201|COMP|23652-1|LNC|Aeromonas salmonicida DNA|Aeromonas salmonicida DNA
C0881032|T201|COMP|23653-9|LNC|Aflatoxin|Aflatoxin
C0881033|T201|COMP|23654-7|LNC|Aflatoxin|Aflatoxin
C0881034|T201|COMP|23655-4|LNC|Aflatoxin|Aflatoxin
C0881035|T201|COMP|23656-2|LNC|Ammonia|Ammonia
C0881036|T201|COMP|23657-0|LNC|Anaplasma marginale Ab|Anaplasma marginale Ab
C0881037|T201|COMP|23658-8|LNC|Antibiotic XXX|Antibiotic XXX
C0881038|T201|COMP|23659-6|LNC|Apramycin|Apramycin
C0881039|T201|COMP|23660-4|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C0881040|T201|COMP|23661-2|LNC|Avian paramyxovirus 1 Ab|Avian paramyxovirus 1 Ab
C0881041|T201|COMP|23662-0|LNC|Babesia bigemina Ab|Babesia bigemina Ab
C0881042|T201|COMP|23663-8|LNC|Babesia bovis Ab|Babesia bovis Ab
C0881043|T201|COMP|23664-6|LNC|Babesia canis Ab|Babesia canis Ab
C0881044|T201|COMP|23665-3|LNC|Babesia divergens Ab|Babesia divergens Ab
C0881045|T201|COMP|23666-1|LNC|Babesia sp Ab|Babesia sp Ab
C0881046|T201|COMP|23667-9|LNC|Bacteria identified|Bacteria identified
C0881047|T201|COMP|23668-7|LNC|Bartonella henselae Ab|Bartonella henselae Ab
C0881048|T201|COMP|23669-5|LNC|Biochanin A|Biochanin A
C0881049|T201|COMP|23670-3|LNC|Blastomyces sp Ab|Blastomyces sp Ab
C0881050|T201|COMP|23671-1|LNC|Bluetongue virus 10 Ab|Bluetongue virus 10 Ab
C0881051|T201|COMP|23672-9|LNC|Bluetongue virus 11 Ab|Bluetongue virus 11 Ab
C0881052|T201|COMP|23673-7|LNC|Bluetongue virus 13 Ab|Bluetongue virus 13 Ab
C0881053|T201|COMP|23675-2|LNC|Bluetongue virus 2 Ab|Bluetongue virus 2 Ab
C0881054|T201|COMP|23676-0|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0881055|T201|COMP|23677-8|LNC|Bovine leukemia virus Ab|Bovine leukemia virus Ab
C0881056|T201|COMP|23678-6|LNC|Bovine parainfluenza virus 3 Ag|Bovine parainfluenza virus 3 Ag
C0881057|T201|COMP|23679-4|LNC|Bovine respiratory syncytial virus Ag|Bovine respiratory syncytial virus Ag
C0881058|T201|COMP|23680-2|LNC|Bromide|Bromide
C0881059|T201|COMP|23681-0|LNC|Brucella canis Ab|Brucella canis Ab
C0881060|T201|COMP|23682-8|LNC|Brucella canis Ab|Brucella canis Ab
C0881061|T201|COMP|23683-6|LNC|Brucella canis Ab|Brucella canis Ab
C0881062|T201|COMP|23685-1|LNC|Canine adenovirus 1 Ab|Canine adenovirus 1 Ab
C0881063|T201|COMP|23686-9|LNC|Canine adenovirus Ag|Canine adenovirus Ag
C0881064|T201|COMP|23689-3|LNC|Canine distemper virus Ab|Canine distemper virus Ab
C0881065|T201|COMP|23690-1|LNC|Canine distemper virus Ab|Canine distemper virus Ab
C0881066|T201|COMP|23691-9|LNC|Canine distemper virus Ab.IgG|Canine distemper virus Ab.IgG
C0881067|T201|COMP|23693-5|LNC|Canine distemper virus Ab.IgM|Canine distemper virus Ab.IgM
C0881068|T201|COMP|23694-3|LNC|Canine distemper virus Ab.IgM|Canine distemper virus Ab.IgM
C0881069|T201|COMP|23695-0|LNC|Canine distemper virus Ag|Canine distemper virus Ag
C0881070|T201|COMP|23696-8|LNC|Canine distemper virus Ag|Canine distemper virus Ag
C0881071|T201|COMP|23698-4|LNC|Canine herpesvirus Ag|Canine herpesvirus Ag
C0881072|T201|COMP|23699-2|LNC|Canine parainfluenza virus 2 Ag|Canine parainfluenza virus 2 Ag
C0881073|T201|COMP|23700-8|LNC|Canine parvovirus Ab|Canine parvovirus Ab
C0881074|T201|COMP|23701-6|LNC|Canine parvovirus Ab|Canine parvovirus Ab
C0881075|T201|COMP|23702-4|LNC|Canine parvovirus Ab|Canine parvovirus Ab
C0881076|T201|COMP|23703-2|LNC|Canine parvovirus Ab.IgG|Canine parvovirus Ab.IgG
C0881077|T201|COMP|23704-0|LNC|Canine parvovirus Ab.IgM|Canine parvovirus Ab.IgM
C0881078|T201|COMP|23705-7|LNC|Canine parvovirus Ag|Canine parvovirus Ag
C0881079|T201|COMP|23706-5|LNC|Canine parvovirus Ag|Canine parvovirus Ag
C0881080|T201|COMP|23707-3|LNC|Canine parvovirus DNA|Canine parvovirus DNA
C0881081|T201|COMP|23708-1|LNC|Caprine arthritis encephalitis virus Ag|Caprine arthritis encephalitis virus Ag
C0881082|T201|COMP|23710-7|LNC|Dirofilaria immitis Ag|Dirofilaria immitis Ag
C0881083|T201|COMP|23711-5|LNC|Ehrlichia canis Ab|Ehrlichia canis Ab
C0881084|T201|COMP|23712-3|LNC|Enrofloxacin|Enrofloxacin
C0881085|T201|COMP|23713-1|LNC|Ethylene glycol|Ethylene glycol
C0881087|T201|COMP|23715-6|LNC|Feline calicivirus Ab|Feline calicivirus Ab
C0881088|T201|COMP|23716-4|LNC|Feline coronavirus Ab|Feline coronavirus Ab
C0881089|T201|COMP|23717-2|LNC|Feline coronavirus Ab|Feline coronavirus Ab
C0881090|T201|COMP|23718-0|LNC|Feline coronavirus Ab|Feline coronavirus Ab
C0881091|T201|COMP|23719-8|LNC|Feline herpesvirus 1 Ab|Feline herpesvirus 1 Ab
C0881092|T201|COMP|23720-6|LNC|Feline herpesvirus 1 Ag|Feline herpesvirus 1 Ag
C0881093|T201|COMP|23721-4|LNC|Feline herpesvirus 1 DNA|Feline herpesvirus 1 DNA
C0881094|T201|COMP|23722-2|LNC|Feline herpesvirus Ab|Feline herpesvirus Ab
C0881095|T201|COMP|23723-0|LNC|Feline immunodeficiency virus Ab|Feline immunodeficiency virus Ab
C0881096|T201|COMP|23724-8|LNC|Feline immunodeficiency virus Ab|Feline immunodeficiency virus Ab
C0881097|T201|COMP|23725-5|LNC|Feline immunodeficiency virus Ab|Feline immunodeficiency virus Ab
C0881098|T201|COMP|23726-3|LNC|Feline infectious peritonitis virus Ab|Feline infectious peritonitis virus Ab
C0881099|T201|COMP|23727-1|LNC|Feline infectious peritonitis virus Ab|Feline infectious peritonitis virus Ab
C0881100|T201|COMP|23728-9|LNC|Feline infectious peritonitis virus Ab|Feline infectious peritonitis virus Ab
C0881101|T201|COMP|23729-7|LNC|Feline infectious peritonitis virus Ag|Feline infectious peritonitis virus Ag
C0881102|T201|COMP|23730-5|LNC|Feline infectious peritonitis virus Ag|Feline infectious peritonitis virus Ag
C0881103|T201|COMP|23731-3|LNC|Feline leukemia provirus|Feline leukemia provirus
C0881104|T201|COMP|23733-9|LNC|Feline leukemia virus Ab|Feline leukemia virus Ab
C0881105|T201|COMP|23734-7|LNC|Feline leukemia virus Ab|Feline leukemia virus Ab
C0881106|T201|COMP|23736-2|LNC|Feline leukemia virus Ag|Feline leukemia virus Ag
C0881107|T201|COMP|23737-0|LNC|Feline panleukopenia virus Ab|Feline panleukopenia virus Ab
C0881108|T201|COMP|23739-6|LNC|Feline syncytial virus Ab|Feline syncytial virus Ab
C0881109|T201|COMP|23740-4|LNC|Florfenicol|Florfenicol
C0881110|T201|COMP|23741-2|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C0881111|T201|COMP|23743-8|LNC|Genistein|Genistein
C0881112|T201|COMP|23744-6|LNC|Giardia lamblia Ag|Giardia lamblia Ag
C0881113|T201|COMP|23745-3|LNC|Gossypol|Gossypol
C0881114|T201|COMP|23747-9|LNC|Heavy metals|Heavy metals
C0881115|T201|COMP|23748-7|LNC|Histoplasma sp Ab|Histoplasma sp Ab
C0881116|T201|COMP|23749-5|LNC|Lead|Lead
C0881117|T201|COMP|23751-1|LNC|Metaldehyde|Metaldehyde
C0881118|T201|COMP|23752-9|LNC|Mite identified|Mite identified
C0881119|T201|COMP|23753-7|LNC|Mycoplasma hyopneumoniae Ab|Mycoplasma hyopneumoniae Ab
C0881120|T201|COMP|23755-2|LNC|Mycoplasma synoviae Ab|Mycoplasma synoviae Ab
C0881121|T201|COMP|23756-0|LNC|Neospora caninum Ab|Neospora caninum Ab
C0881122|T201|COMP|23757-8|LNC|Neospora caninum Ab|Neospora caninum Ab
C0881123|T201|COMP|23758-6|LNC|Neospora caninum Ab|Neospora caninum Ab
C0881124|T201|COMP|23760-2|LNC|Neospora caninum Ag|Neospora caninum Ag
C0881125|T201|COMP|23761-0|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0881126|T201|COMP|23762-8|LNC|Nitrate+Nitrite|Nitrate+Nitrite
C0881127|T201|COMP|23763-6|LNC|Pasteurella multocida serotype|Pasteurella multocida serotype
C0881128|T201|COMP|23764-4|LNC|Pesticides|Pesticides
C0881129|T201|COMP|23765-1|LNC|Porcine adenovirus Ag|Porcine adenovirus Ag
C0881130|T201|COMP|23766-9|LNC|Porcine circovirus Ag|Porcine circovirus Ag
C0881131|T201|COMP|23767-7|LNC|Porcine circovirus Ag|Porcine circovirus Ag
C0881132|T201|COMP|23768-5|LNC|Porcine influenza virus A Ab|Porcine influenza virus A Ab
C0881133|T201|COMP|23769-3|LNC|Porcine influenza virus A Ag|Porcine influenza virus A Ag
C0881134|T201|COMP|23770-1|LNC|Porcine parvovirus Ab|Porcine parvovirus Ab
C0881136|T201|COMP|23773-5|LNC|Porcine rotavirus Ag|Porcine rotavirus Ag
C0881137|T201|COMP|23774-3|LNC|Pseudorabies virus Ag|Pseudorabies virus Ag
C0881138|T201|COMP|23775-0|LNC|Rhodococcus equi Ab|Rhodococcus equi Ab
C0881139|T201|COMP|23776-8|LNC|Rickettsia spotted fever group Ab|Rickettsia spotted fever group Ab
C0881140|T201|COMP|23777-6|LNC|Salmonella pullorum Ab|Salmonella pullorum Ab
C0881141|T201|COMP|23778-4|LNC|Salmonella typhimurium Ab|Salmonella typhimurium Ab
C0881142|T201|COMP|23779-2|LNC|Selenium|Selenium
C0881143|T201|COMP|23780-0|LNC|Strychnine|Strychnine
C0881144|T201|COMP|23781-8|LNC|Swine influenza virus Ag|Swine influenza virus Ag
C0881145|T201|COMP|23782-6|LNC|Swine influenza virus Ag|Swine influenza virus Ag
C0881146|T201|COMP|23783-4|LNC|Taylorella equigenitalis Ab|Taylorella equigenitalis Ab
C0881147|T201|COMP|23784-2|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C0881148|T201|COMP|23785-9|LNC|Trypanosoma cruzi Ab|Trypanosoma cruzi Ab
C0881149|T201|COMP|23786-7|LNC|Urea|Urea
C0881150|T201|COMP|23787-5|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C0881151|T201|COMP|23788-3|LNC|Vesicular stomatitis Indiana virus Ab|Vesicular stomatitis Indiana virus Ab
C0881152|T201|COMP|23789-1|LNC|Vesicular stomatitis Indiana virus Ab|Vesicular stomatitis Indiana virus Ab
C0881153|T201|COMP|23790-9|LNC|Vesicular stomatitis New Jersey virus Ab|Vesicular stomatitis New Jersey virus Ab
C0881154|T201|COMP|23791-7|LNC|Vesicular stomatitis New Jersey virus Ab|Vesicular stomatitis New Jersey virus Ab
C0881155|T201|COMP|23792-5|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C0881156|T201|COMP|23793-3|LNC|Canine parvovirus Ag|Canine parvovirus Ag
C0881165|T201|COMP|23805-5|LNC|5-Fluorocytosine|5-Fluorocytosine
C0881166|T201|COMP|23806-3|LNC|Albumin^2H post peritoneal dialysis|Albumin^2H post peritoneal dialysis
C0881167|T201|COMP|23807-1|LNC|Albumin^4H post peritoneal dialysis|Albumin^4H post peritoneal dialysis
C0881168|T201|COMP|23808-9|LNC|Aldosterone.free|Aldosterone.free
C0881169|T201|COMP|23809-7|LNC|Alloisoleucine|Alloisoleucine
C0881170|T201|COMP|23810-5|LNC|Alpha fucosidase|Alpha fucosidase
C0881171|T201|COMP|23811-3|LNC|Alpha-1-Fetoprotein^^adjusted|Alpha-1-Fetoprotein^^adjusted
C0881172|T201|COMP|23812-1|LNC|Alpha-1-Fetoprotein^^unadjusted|Alpha-1-Fetoprotein^^unadjusted
C0881173|T201|COMP|23813-9|LNC|Alternaria sp Ab.IgE.RAST class|Alternaria sp Ab.IgE.RAST class
C0881174|T201|COMP|23815-4|LNC|Androstanediol|Androstanediol
C0881175|T201|COMP|23816-2|LNC|Antibiotic XXX|Antibiotic XXX
C0881176|T201|COMP|23817-0|LNC|Antibiotic XXX^peak|Antibiotic XXX^peak
C0881177|T201|COMP|23819-6|LNC|Antibody coated bacteria|Antibody coated bacteria
C0881178|T201|COMP|23820-4|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C0881179|T201|COMP|23821-2|LNC|Aspergillus fumigatus Ab|Aspergillus fumigatus Ab
C0881180|T201|COMP|23822-0|LNC|Azinphos-methyl|Azinphos-methyl
C0881181|T201|COMP|23823-8|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0881184|T201|COMP|23826-1|LNC|Bordetella pertussis DNA|Bordetella pertussis DNA
C0881188|T201|COMP|23830-3|LNC|Bordetella pertussis.pertussis toxin Ab.IgA|Bordetella pertussis.pertussis toxin Ab.IgA
C0881189|T201|COMP|23831-1|LNC|Bordetella pertussis.pertussis toxin Ab.IgG|Bordetella pertussis.pertussis toxin Ab.IgG
C0881190|T201|COMP|23832-9|LNC|Bordetella pertussis.pertussis toxin Ab.IgM|Bordetella pertussis.pertussis toxin Ab.IgM
C0881191|T201|COMP|23833-7|LNC|Borrelia burgdorferi Ab index|Borrelia burgdorferi Ab index
C0881192|T201|COMP|23834-5|LNC|Canary droppings Ab.IgE.RAST class|Canary droppings Ab.IgE.RAST class
C0881193|T201|COMP|23835-2|LNC|Carbon disulfide|Carbon disulfide
C0881194|T201|COMP|23836-0|LNC|Carbon disulfide|Carbon disulfide
C0881195|T201|COMP|23837-8|LNC|Chicken serum proteins Ab.IgE.RAST class|Chicken serum proteins Ab.IgE.RAST class
C0881196|T201|COMP|23838-6|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C0881197|T201|COMP|23839-4|LNC|Cholinesterase|Cholinesterase
C0881198|T201|COMP|23840-2|LNC|Choriogonadotropin.beta subunit^^unadjusted|Choriogonadotropin.beta subunit^^unadjusted
C0881199|T201|COMP|23841-0|LNC|Choriogonadotropin.beta subunit^^adjusted|Choriogonadotropin.beta subunit^^adjusted
C0881200|T201|COMP|23842-8|LNC|Cobalt|Cobalt
C0881201|T201|COMP|23843-6|LNC|Cockatiel droppings Ab|Cockatiel droppings Ab
C0881202|T201|COMP|23844-4|LNC|C3 nephritic factor|C3 nephritic factor
C0881203|T201|COMP|23845-1|LNC|Coproporphyrin 1|Coproporphyrin 1
C0881204|T201|COMP|23846-9|LNC|Coproporphyrin 3|Coproporphyrin 3
C0881205|T201|COMP|23850-1|LNC|Creosol|Creosol
C0881206|T201|COMP|23852-7|LNC|Deuteroporphyrin|Deuteroporphyrin
C0881207|T201|COMP|23853-5|LNC|Dimethylformamide/Creatinine|Dimethylformamide/Creatinine
C0881208|T201|COMP|23854-3|LNC|Dioxin|Dioxin
C0881209|T201|COMP|23855-0|LNC|Echinococcus granulosus Ab.IgE|Echinococcus granulosus Ab.IgE
C0881210|T201|COMP|23857-6|LNC|Epidermis Ab|Epidermis Ab
C0881211|T201|COMP|23858-4|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C0881212|T201|COMP|23859-2|LNC|Erythrocytes|Erythrocytes
C0881213|T201|COMP|23860-0|LNC|Erythrocytes|Erythrocytes
C0881214|T201|COMP|23861-8|LNC|Ethanol|Ethanol
C0881215|T201|COMP|23862-6|LNC|Famotidine|Famotidine
C0881216|T201|COMP|23864-2|LNC|Flunitrazepam|Flunitrazepam
C0881217|T201|COMP|23865-9|LNC|Fluoxetine+Norfluoxetine|Fluoxetine+Norfluoxetine
C0881218|T201|COMP|23866-7|LNC|Glutaraldehyde|Glutaraldehyde
C0881219|T201|COMP|23867-5|LNC|Hantavirus sin nombre Ab.IgG|Hantavirus sin nombre Ab.IgG
C0881220|T201|COMP|23868-3|LNC|Hantavirus sin nombre Ab.IgM|Hantavirus sin nombre Ab.IgM
C0881221|T201|COMP|23870-9|LNC|Hepatitis C virus 100+5-1-1 Ab|Hepatitis C virus 100+5-1-1 Ab
C0881222|T201|COMP|23871-7|LNC|Hepatitis C virus NS5 Ab|Hepatitis C virus NS5 Ab
C0881223|T201|COMP|23872-5|LNC|Heptacarboxylporphyrin I|Heptacarboxylporphyrin I
C0881224|T201|COMP|23874-1|LNC|Hexacarboxylporphyrin I|Hexacarboxylporphyrin I
C0881225|T201|COMP|23875-8|LNC|Hexacarboxylporphyrin III|Hexacarboxylporphyrin III
C0881226|T201|COMP|23876-6|LNC|HIV 1 RNA|HIV 1 RNA
C0881227|T201|COMP|23877-4|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C0881228|T201|COMP|23878-2|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C0881229|T201|COMP|23879-0|LNC|Immune complex|Immune complex
C0881230|T201|COMP|23880-8|LNC|Immune complex|Immune complex
C0881231|T201|COMP|23881-6|LNC|Immune complex|Immune complex
C0881232|T201|COMP|23882-4|LNC|Immune complex|Immune complex
C0881233|T201|COMP|23883-2|LNC|Inhibin A|Inhibin A
C0881234|T201|COMP|23884-0|LNC|Interleukin 2 receptor|Interleukin 2 receptor
C0881235|T201|COMP|23885-7|LNC|Isoheptacarboxylporphyrin|Isoheptacarboxylporphyrin
C0881236|T201|COMP|23886-5|LNC|Isohexacarboxylporphyrin|Isohexacarboxylporphyrin
C0881237|T201|COMP|23887-3|LNC|Isopentacarboxylporphyrin|Isopentacarboxylporphyrin
C0881238|T201|COMP|23888-1|LNC|Isopropanol|Isopropanol
C0881239|T201|COMP|23889-9|LNC|Kanamycin|Kanamycin
C0881240|T201|COMP|23891-5|LNC|Magnesium|Magnesium
C0881241|T201|COMP|23892-3|LNC|Magnesium|Magnesium
C0881242|T201|COMP|23893-1|LNC|Malaoxon|Malaoxon
C0881243|T201|COMP|23894-9|LNC|Maple Ab.IgE.RAST class|Maple Ab.IgE.RAST class
C0881244|T201|COMP|23895-6|LNC|Mattress dust Ab.IgE.RAST class|Mattress dust Ab.IgE.RAST class
C0881245|T201|COMP|23896-4|LNC|Mercury|Mercury
C0881246|T201|COMP|23897-2|LNC|Mesothelial cells|Mesothelial cells
C0881247|T201|COMP|23898-0|LNC|Mesothelial cells|Mesothelial cells
C0881248|T201|COMP|23899-8|LNC|Methanol|Methanol
C0881249|T201|COMP|23900-4|LNC|Methanol|Methanol
C0881251|T201|COMP|23903-8|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C0881252|T201|COMP|23904-6|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C0881253|T201|COMP|23905-3|LNC|Mycophenolate|Mycophenolate
C0881254|T201|COMP|23906-1|LNC|Mycophenolate glucuronide|Mycophenolate glucuronide
C0881256|T201|COMP|23909-5|LNC|Trisetum paniceum Ab.IgE.RAST class|Trisetum paniceum Ab.IgE.RAST class
C0881257|T201|COMP|23910-3|LNC|Osmotic fragility^0.0% sodium chloride|Osmotic fragility^0.0% sodium chloride
C0881258|T201|COMP|23911-1|LNC|Osmotic fragility^0.30% sodium chloride|Osmotic fragility^0.30% sodium chloride
C0881259|T201|COMP|23913-7|LNC|Osmotic fragility^0.40% sodium chloride|Osmotic fragility^0.40% sodium chloride
C0881260|T201|COMP|23914-5|LNC|Osmotic fragility^0.45% sodium chloride|Osmotic fragility^0.45% sodium chloride
C0881261|T201|COMP|23916-0|LNC|Osmotic fragility^0.55% sodium chloride|Osmotic fragility^0.55% sodium chloride
C0881262|T201|COMP|23917-8|LNC|Osmotic fragility^0.60% sodium chloride|Osmotic fragility^0.60% sodium chloride
C0881263|T201|COMP|23919-4|LNC|Osmotic fragility^0.65% sodium chloride|Osmotic fragility^0.65% sodium chloride
C0881266|T201|COMP|23922-8|LNC|Osmotic fragility^0.85% sodium chloride|Osmotic fragility^0.85% sodium chloride
C0881267|T201|COMP|23924-4|LNC|Parakeet serum Ab.IgE.RAST class|Parakeet serum Ab.IgE.RAST class
C0881268|T201|COMP|23925-1|LNC|Penicillin|Penicillin
C0881269|T201|COMP|23926-9|LNC|Pepper bell Ab.IgE.RAST class|Pepper bell Ab.IgE.RAST class
C0881270|T201|COMP|23927-7|LNC|Pepper white Ab.IgE.RAST class|Pepper white Ab.IgE.RAST class
C0881271|T201|COMP|23930-1|LNC|Salmonella typhi O D Ab|Salmonella typhi O D Ab
C0881272|T201|COMP|23931-9|LNC|Salmonella typhi O D|Salmonella typhi O D
C0881273|T201|COMP|23932-7|LNC|Squash zucchini Ab.IgE.RAST class|Squash zucchini Ab.IgE.RAST class
C0881274|T201|COMP|23934-3|LNC|Staphylococcus aureus enterotoxin B Ab|Staphylococcus aureus enterotoxin B Ab
C0881277|T201|COMP|23937-6|LNC|Trans nonachlor|Trans nonachlor
C0881278|T201|COMP|23938-4|LNC|Trapa natans Ab.IgE.RAST class|Trapa natans Ab.IgE.RAST class
C0881279|T201|COMP|23939-2|LNC|Xylose^1H post 5 g xylose PO|Xylose^1H post 5 g xylose PO
C0881280|T201|COMP|23940-0|LNC|Xylose^1H post dose xylose PO|Xylose^1H post dose xylose PO
C0881281|T201|COMP|23942-6|LNC|Xylose^2H post 5 g xylose PO|Xylose^2H post 5 g xylose PO
C0881282|T201|COMP|23943-4|LNC|Xylose^2H post dose xylose PO|Xylose^2H post dose xylose PO
C0881283|T201|COMP|23945-9|LNC|Xylose^1H post 5 g xylose PO|Xylose^1H post 5 g xylose PO
C0881284|T201|COMP|23946-7|LNC|Xylose^1H post dose xylose PO|Xylose^1H post dose xylose PO
C0881285|T201|COMP|23947-5|LNC|Isoniazid|Isoniazid
C0881286|T201|COMP|23948-3|LNC|Ofloxacin|Ofloxacin
C0881287|T201|COMP|23949-1|LNC|rifAMPin|rifAMPin
C0881288|T201|COMP|23950-9|LNC|Adenovirus Ab|Adenovirus Ab
C0881289|T201|COMP|23951-7|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C0881290|T201|COMP|23952-5|LNC|Asialoganglioside GM1 Ab.IgM|Asialoganglioside GM1 Ab.IgM
C0881291|T201|COMP|23953-3|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C0881292|T201|COMP|23954-1|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C0881293|T201|COMP|23955-8|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C0881294|T201|COMP|23956-6|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C0881295|T201|COMP|23957-4|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C0881296|T201|COMP|23958-2|LNC|Dengue virus Ab.IgG|Dengue virus Ab.IgG
C0881297|T201|COMP|23959-0|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0881298|T201|COMP|23960-8|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C0881299|T201|COMP|23961-6|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C0881300|T201|COMP|23962-4|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C0881301|T201|COMP|23963-2|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C0881302|T201|COMP|23964-0|LNC|Brucella abortus Ab.IgM|Brucella abortus Ab.IgM
C0881303|T201|COMP|23966-5|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0881304|T201|COMP|23967-3|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0881305|T201|COMP|23968-1|LNC|Dengue virus Ab.IgM|Dengue virus Ab.IgM
C0881306|T201|COMP|23969-9|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C0881307|T201|COMP|23970-7|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0881308|T201|COMP|23971-5|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C0881309|T201|COMP|23972-3|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C0881310|T201|COMP|23973-1|LNC|Burkholderia pseudomallei Ab.IgM|Burkholderia pseudomallei Ab.IgM
C0881311|T201|COMP|23975-6|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C0881312|T201|COMP|23976-4|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0881313|T201|COMP|23977-2|LNC|Borrelia burgdorferi Ag|Borrelia burgdorferi Ag
C0881314|T201|COMP|23978-0|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0881315|T201|COMP|23980-6|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0881316|T201|COMP|23981-4|LNC|Borrelia burgdorferi Ab.IgG band pattern|Borrelia burgdorferi Ab.IgG band pattern
C0881317|T201|COMP|23982-2|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0881318|T201|COMP|23983-0|LNC|Borrelia burgdorferi Ab.IgM band pattern|Borrelia burgdorferi Ab.IgM band pattern
C0881319|T201|COMP|23985-5|LNC|Borrelia burgdorferi Ab.IgM band pattern|Borrelia burgdorferi Ab.IgM band pattern
C0881320|T201|COMP|23986-3|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C0881321|T201|COMP|23987-1|LNC|Brucella abortus Ab.IgM|Brucella abortus Ab.IgM
C0881322|T201|COMP|23988-9|LNC|Burkholderia pseudomallei Ab.IgG|Burkholderia pseudomallei Ab.IgG
C0881323|T201|COMP|23990-5|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0881324|T201|COMP|23991-3|LNC|Dengue virus Ab.IgG|Dengue virus Ab.IgG
C0881325|T201|COMP|23992-1|LNC|Dengue virus Ab.IgM|Dengue virus Ab.IgM
C0881326|T201|COMP|23994-7|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0881327|T201|COMP|23995-4|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C0881328|T201|COMP|23996-2|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C0881329|T201|COMP|23997-0|LNC|Ganglioside GD1a Ab.IgG|Ganglioside GD1a Ab.IgG
C0881330|T201|COMP|23998-8|LNC|Ganglioside GD1a Ab.IgM|Ganglioside GD1a Ab.IgM
C0881331|T201|COMP|23999-6|LNC|Ganglioside GD1b Ab.IgG|Ganglioside GD1b Ab.IgG
C0881332|T201|COMP|24000-2|LNC|Ganglioside GD1b Ab.IgM|Ganglioside GD1b Ab.IgM
C0881333|T201|COMP|24001-0|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C0881335|T201|COMP|24003-6|LNC|Brucella sp identified|Brucella sp identified
C0881336|T201|COMP|24004-4|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C0881337|T201|COMP|24005-1|LNC|Chlamydia sp identified|Chlamydia sp identified
C0881338|T201|COMP|24006-9|LNC|Eastern equine encephalitis virus Ab.IgG & IgM|Eastern equine encephalitis virus Ab.IgG & IgM
C0881339|T201|COMP|24007-7|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C0881340|T201|COMP|24008-5|LNC|Echovirus 14 Ab|Echovirus 14 Ab
C0881341|T201|COMP|24009-3|LNC|Fungus identified|Fungus identified
C0881342|T201|COMP|24010-1|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C0881343|T201|COMP|24012-7|LNC|HIV 1 Ag|HIV 1 Ag
C0881344|T201|COMP|24013-5|LNC|HIV 1 RNA|HIV 1 RNA
C0881345|T201|COMP|24014-3|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0881346|T201|COMP|24015-0|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C0881347|T201|COMP|24016-8|LNC|La Crosse virus Ab|La Crosse virus Ab
C0881348|T201|COMP|24017-6|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C0881349|T201|COMP|24018-4|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C0881350|T201|COMP|24019-2|LNC|Neisseria meningitdis B Ag|Neisseria meningitdis B Ag
C0881351|T201|COMP|24020-0|LNC|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C0881352|T201|COMP|24021-8|LNC|Streptococcus pneumoniae 12 Ab|Streptococcus pneumoniae 12 Ab
C0881353|T201|COMP|24022-6|LNC|Streptococcus pneumoniae 14 Ab|Streptococcus pneumoniae 14 Ab
C0881354|T201|COMP|24023-4|LNC|Streptococcus pneumoniae 3 Ab|Streptococcus pneumoniae 3 Ab
C0881355|T201|COMP|24025-9|LNC|Streptococcus pneumoniae 8 Ab|Streptococcus pneumoniae 8 Ab
C0881356|T201|COMP|24027-5|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C0881357|T201|COMP|24028-3|LNC|Toxocara canis Ab.IgA|Toxocara canis Ab.IgA
C0881358|T201|COMP|24029-1|LNC|Toxocara canis Ab.IgG|Toxocara canis Ab.IgG
C0881359|T201|COMP|24030-9|LNC|Toxocara canis Ab.IgM|Toxocara canis Ab.IgM
C0881360|T201|COMP|24031-7|LNC|14-3-3 Ag|14-3-3 Ag
C0881361|T201|COMP|24032-5|LNC|Rifabutin|Rifabutin
C0881364|T201|COMP|24036-6|LNC|Borrelia sp Ag|Borrelia sp Ag
C0881365|T201|COMP|24037-4|LNC|Coccidioides immitis rRNA|Coccidioides immitis rRNA
C0881366|T201|COMP|24038-2|LNC|Cryoglobulin type|Cryoglobulin type
C0881367|T201|COMP|24039-0|LNC|Taenia solium larva Ab.IgG band pattern|Taenia solium larva Ab.IgG band pattern
C0881368|T201|COMP|24040-8|LNC|Taenia solium larva Ab.IgG band pattern|Taenia solium larva Ab.IgG band pattern
C0881369|T201|COMP|24041-6|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C0881370|T201|COMP|24042-4|LNC|Ehrlichia chaffeensis DNA|Ehrlichia chaffeensis DNA
C0881371|T201|COMP|24044-0|LNC|Acetyl-CoA:glucosamine acetyltransferase|Acetyl-CoA:glucosamine acetyltransferase
C0881372|T201|COMP|24045-7|LNC|Alpha fucosidase|Alpha fucosidase
C0881373|T201|COMP|24046-5|LNC|Alpha fucosidase|Alpha fucosidase
C0881374|T201|COMP|24047-3|LNC|Alpha fucosidase|Alpha fucosidase
C0881375|T201|COMP|24050-7|LNC|Acid alpha glucosidase|Acid alpha glucosidase
C0881376|T201|COMP|24051-5|LNC|Acid alpha glucosidase|Acid alpha glucosidase
C0881377|T201|COMP|24053-1|LNC|Alpha mannosidase|Alpha mannosidase
C0881378|T201|COMP|24054-9|LNC|Alpha-N-acetylgalactosaminidase|Alpha-N-acetylgalactosaminidase
C0881379|T201|COMP|24055-6|LNC|Alpha-N-acetylgalactosaminidase|Alpha-N-acetylgalactosaminidase
C0881380|T201|COMP|24056-4|LNC|Alpha-L-iduronidase|Alpha-L-iduronidase
C0881381|T201|COMP|24058-0|LNC|Aspartylglucosaminidase|Aspartylglucosaminidase
C0881382|T201|COMP|24059-8|LNC|Aspartylglucosaminidase|Aspartylglucosaminidase
C0881383|T201|COMP|24060-6|LNC|Beta galactosidase|Beta galactosidase
C0881384|T201|COMP|24061-4|LNC|Beta galactosidase|Beta galactosidase
C0881385|T201|COMP|24064-8|LNC|Beta glucuronidase|Beta glucuronidase
C0881386|T201|COMP|24066-3|LNC|Beta mannosidase|Beta mannosidase
C0881387|T201|COMP|24067-1|LNC|Beta mannosidase|Beta mannosidase
C0881388|T201|COMP|24068-9|LNC|Beta mannosidase|Beta mannosidase
C0881392|T201|COMP|24072-1|LNC|Beta-N-acetylhexosaminidase.B|Beta-N-acetylhexosaminidase.B
C0881393|T201|COMP|24073-9|LNC|Beta-N-acetylhexosaminidase.B|Beta-N-acetylhexosaminidase.B
C0881394|T201|COMP|24074-7|LNC|Beta-N-acetylhexosaminidase|Beta-N-acetylhexosaminidase
C0881395|T201|COMP|24075-4|LNC|Beta-N-acetylhexosaminidase|Beta-N-acetylhexosaminidase
C0881396|T201|COMP|24076-2|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C0881397|T201|COMP|24077-0|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C0881398|T201|COMP|24078-8|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C0881399|T201|COMP|24079-6|LNC|Cholesterol esterase|Cholesterol esterase
C0881400|T201|COMP|24080-4|LNC|Cholesterol esterase|Cholesterol esterase
C0881402|T201|COMP|24082-0|LNC|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C0881403|T201|COMP|24083-8|LNC|Galactosylceramidase|Galactosylceramidase
C0881404|T201|COMP|24084-6|LNC|Galactosylceramidase|Galactosylceramidase
C0881405|T201|COMP|24085-3|LNC|Heparan-N-sulfatase|Heparan-N-sulfatase
C0881406|T201|COMP|24086-1|LNC|Heparan-N-sulfatase|Heparan-N-sulfatase
C0881407|T201|COMP|24087-9|LNC|Iduronate-2-Sulfatase|Iduronate-2-Sulfatase
C0881408|T201|COMP|24088-7|LNC|Iduronate-2-Sulfatase|Iduronate-2-Sulfatase
C0881409|T201|COMP|24089-5|LNC|Iduronate-2-Sulfatase|Iduronate-2-Sulfatase
C0881410|T201|COMP|1837-4|LNC|Alpha-N-acetylglucosaminidase|Alpha-N-acetylglucosaminidase
C0881411|T201|COMP|24093-7|LNC|N-Acetylgalactosamine-4-Sulfatase|N-Acetylgalactosamine-4-Sulfatase
C0881412|T201|COMP|24094-5|LNC|N-Acetylgalactosamine-4-Sulfatase|N-Acetylgalactosamine-4-Sulfatase
C0881413|T201|COMP|24095-2|LNC|N-Acetylgalactosamine-6-Sulfatase|N-Acetylgalactosamine-6-Sulfatase
C0881414|T201|COMP|24097-8|LNC|N-Acetylglucosamine-6-Sulfatase|N-Acetylglucosamine-6-Sulfatase
C0881415|T201|COMP|24098-6|LNC|N-Acetylglucosamine-6-Sulfatase|N-Acetylglucosamine-6-Sulfatase
C0881416|T201|COMP|24099-4|LNC|Sialidase|Sialidase
C0881417|T201|COMP|24100-0|LNC|Acid sphingomyelinase|Acid sphingomyelinase
C0881418|T201|COMP|24101-8|LNC|Acid sphingomyelinase|Acid sphingomyelinase
C0881419|T201|COMP|24102-6|LNC|Corynebacterium spp toxin|Corynebacterium spp toxin
C0881420|T201|COMP|24104-2|LNC|Lymphoma cells/100 leukocytes|Lymphoma cells/100 leukocytes
C0881421|T201|COMP|24105-9|LNC|Lymphoma cells|Lymphoma cells
C0881422|T201|COMP|24106-7|LNC|Hairy cells/100 leukocytes|Hairy cells/100 leukocytes
C0881423|T201|COMP|24107-5|LNC|Hairy cells|Hairy cells
C0881424|T201|COMP|24109-1|LNC|Progesterone|Progesterone
C0881425|T201|COMP|24110-9|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0881426|T201|COMP|24111-7|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C0881427|T201|COMP|24113-3|LNC|Hepatitis B virus core Ab.IgM|Hepatitis B virus core Ab.IgM
C0881428|T201|COMP|24114-1|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0881429|T201|COMP|24115-8|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0881430|T201|COMP|24116-6|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C0881431|T201|COMP|24118-2|LNC|Barmah forest virus Ab.IgM|Barmah forest virus Ab.IgM
C0881432|T201|COMP|24119-0|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0881433|T201|COMP|24120-8|LNC|Ross river virus Ab.IgM|Ross river virus Ab.IgM
C0881434|T201|COMP|24121-6|LNC|Barmah forest virus Ab.IgG|Barmah forest virus Ab.IgG
C0881436|T201|COMP|24123-2|LNC|Epithelial cells|Epithelial cells
C0881437|T201|COMP|24124-0|LNC|Casts|Casts
C0881438|T201|COMP|24125-7|LNC|Androgen.free index|Androgen.free index
C0881439|T201|COMP|24126-5|LNC|Adenovirus type|Adenovirus type
C0881440|T201|COMP|24127-3|LNC|Bordetella pertussis.pertussis toxin Ab.IgG|Bordetella pertussis.pertussis toxin Ab.IgG
C0881441|T201|COMP|24128-1|LNC|Bordetella pertussis.pertussis toxin Ab.IgA|Bordetella pertussis.pertussis toxin Ab.IgA
C0881442|T201|COMP|24129-9|LNC|Bordetella pertussis.pertussis toxin Ab.IgM|Bordetella pertussis.pertussis toxin Ab.IgM
C0881443|T201|COMP|24130-7|LNC|Bordetella pertussis.secretory Ab.IgA|Bordetella pertussis.secretory Ab.IgA
C0881449|T201|COMP|24136-4|LNC|Juglans nigra Ab.IgG|Juglans nigra Ab.IgG
C0881450|T201|COMP|24137-2|LNC|Carya tomentosa Ab.IgG|Carya tomentosa Ab.IgG
C0881451|T201|COMP|24138-0|LNC|Sorghum halepense Ab.IgG|Sorghum halepense Ab.IgG
C0881452|T201|COMP|24139-8|LNC|Blatella germanica Ab.IgG|Blatella germanica Ab.IgG
C0881453|T201|COMP|24141-4|LNC|Iva ciliata Ab.IgG|Iva ciliata Ab.IgG
C0881454|T201|COMP|24142-2|LNC|Morus rubra Ab.IgG|Morus rubra Ab.IgG
C0881455|T201|COMP|24143-0|LNC|Rumex acetosella Ab.IgG|Rumex acetosella Ab.IgG
C0881456|T201|COMP|24144-8|LNC|Bromus inermis Ab.IgG|Bromus inermis Ab.IgG
C0881457|T201|COMP|24145-5|LNC|Platanus occidentalis Ab.IgG|Platanus occidentalis Ab.IgG
C0881458|T201|COMP|24146-3|LNC|Acnida tamariscina Ab.IgG|Acnida tamariscina Ab.IgG
C0881460|T201|COMP|24148-9|LNC|Poa pratensis Ab.IgG|Poa pratensis Ab.IgG
C0881462|T201|COMP|24150-5|LNC|Acer rubrum Ab.IgG|Acer rubrum Ab.IgG
C0881463|T201|COMP|24151-3|LNC|Ambrosia trifida Ab.IgG|Ambrosia trifida Ab.IgG
C0881464|T201|COMP|24152-1|LNC|Alternaria alternata Ab.IgG|Alternaria alternata Ab.IgG
C0881464|T201|COMP|25306-2|LNC|Alternaria alternata Ab.IgG|Alternaria alternata Ab.IgG
C0881464|T201|COMP|7076-3|LNC|Alternaria alternata Ab.IgG|Alternaria alternata Ab.IgG
C0881465|T201|COMP|24153-9|LNC|Kamut flour Ab.IgG|Kamut flour Ab.IgG
C0881466|T201|COMP|24154-7|LNC|Chenopodium album Ab.IgG|Chenopodium album Ab.IgG
C0881467|T201|COMP|24156-2|LNC|Maple syrup Ab.IgG|Maple syrup Ab.IgG
C0881468|T201|COMP|6164-8|LNC|Quercus virginiana Ab.IgE|Quercus virginiana Ab.IgE
C0881469|T201|COMP|24158-8|LNC|Pepper white+Pepper black Ab.IgG|Pepper white+Pepper black Ab.IgG
C0881470|T201|COMP|24160-4|LNC|Bean wax Ab.IgE|Bean wax Ab.IgE
C0881470|T201|COMP|16436-8|LNC|Bean wax Ab.IgE|Bean wax Ab.IgE
C0881472|T201|COMP|24162-0|LNC|Aspergillus fumigatus Ab.IgG.RAST class|Aspergillus fumigatus Ab.IgG.RAST class
C0881474|T201|COMP|24165-3|LNC|Beta vulgaris seed Ab.IgE|Beta vulgaris seed Ab.IgE
C0881475|T201|COMP|7609-1|LNC|Pinus radiata Ab.IgE|Pinus radiata Ab.IgE
C0881476|T201|COMP|24168-7|LNC|Cat hair+Cat dander Ab.IgG|Cat hair+Cat dander Ab.IgG
C0881477|T201|COMP|24170-3|LNC|Polio virus 1 Ab^2nd specimen|Polio virus 1 Ab^2nd specimen
C0881478|T201|COMP|24171-1|LNC|Polio virus 2 Ab^1st specimen|Polio virus 2 Ab^1st specimen
C0881479|T201|COMP|24172-9|LNC|Polio virus 2 Ab^2nd specimen|Polio virus 2 Ab^2nd specimen
C0881480|T201|COMP|24174-5|LNC|Polio virus 3 Ab^2nd specimen|Polio virus 3 Ab^2nd specimen
C0881481|T201|COMP|24175-2|LNC|Adenovirus Ab^1st specimen|Adenovirus Ab^1st specimen
C0881482|T201|COMP|24176-0|LNC|Adenovirus Ab^2nd specimen|Adenovirus Ab^2nd specimen
C0881483|T201|COMP|24177-8|LNC|Coxsackievirus B1 Ab^1st specimen|Coxsackievirus B1 Ab^1st specimen
C0881484|T201|COMP|24178-6|LNC|Coxsackievirus B1 Ab^2nd specimen|Coxsackievirus B1 Ab^2nd specimen
C0881485|T201|COMP|24180-2|LNC|Coxsackievirus B1 Ab^2nd specimen|Coxsackievirus B1 Ab^2nd specimen
C0881486|T201|COMP|24181-0|LNC|Coxsackievirus B2 Ab^1st specimen|Coxsackievirus B2 Ab^1st specimen
C0881487|T201|COMP|24182-8|LNC|Coxsackievirus B2 Ab^2nd specimen|Coxsackievirus B2 Ab^2nd specimen
C0881488|T201|COMP|24183-6|LNC|Coxsackievirus B2 Ab^1st specimen|Coxsackievirus B2 Ab^1st specimen
C0881489|T201|COMP|24184-4|LNC|Coxsackievirus B2 Ab^2nd specimen|Coxsackievirus B2 Ab^2nd specimen
C0881490|T201|COMP|24185-1|LNC|Coxsackievirus B3 Ab^1st specimen|Coxsackievirus B3 Ab^1st specimen
C0881491|T201|COMP|24186-9|LNC|Coxsackievirus B3 Ab^2nd specimen|Coxsackievirus B3 Ab^2nd specimen
C0881492|T201|COMP|24187-7|LNC|Coxsackievirus B3 Ab^1st specimen|Coxsackievirus B3 Ab^1st specimen
C0881493|T201|COMP|24188-5|LNC|Coxsackievirus B3 Ab^2nd specimen|Coxsackievirus B3 Ab^2nd specimen
C0881494|T201|COMP|24189-3|LNC|Coxsackievirus B4 Ab^1st specimen|Coxsackievirus B4 Ab^1st specimen
C0881495|T201|COMP|24190-1|LNC|Coxsackievirus B4 Ab^2nd specimen|Coxsackievirus B4 Ab^2nd specimen
C0881496|T201|COMP|24191-9|LNC|Coxsackievirus B4 Ab^1st specimen|Coxsackievirus B4 Ab^1st specimen
C0881497|T201|COMP|24192-7|LNC|Coxsackievirus B4 Ab^2nd specimen|Coxsackievirus B4 Ab^2nd specimen
C0881498|T201|COMP|24193-5|LNC|Coxsackievirus B5 Ab^1st specimen|Coxsackievirus B5 Ab^1st specimen
C0881499|T201|COMP|24194-3|LNC|Coxsackievirus B5 Ab^2nd specimen|Coxsackievirus B5 Ab^2nd specimen
C0881500|T201|COMP|24195-0|LNC|Coxsackievirus B5 Ab^1st specimen|Coxsackievirus B5 Ab^1st specimen
C0881501|T201|COMP|24196-8|LNC|Coxsackievirus B5 Ab^2nd specimen|Coxsackievirus B5 Ab^2nd specimen
C0881502|T201|COMP|24197-6|LNC|Coxsackievirus B6 Ab^1st specimen|Coxsackievirus B6 Ab^1st specimen
C0881503|T201|COMP|24198-4|LNC|Coxsackievirus B6 Ab^2nd specimen|Coxsackievirus B6 Ab^2nd specimen
C0881504|T201|COMP|24199-2|LNC|Coxsackievirus B6 Ab^1st specimen|Coxsackievirus B6 Ab^1st specimen
C0881505|T201|COMP|24200-8|LNC|Coxsackievirus B6 Ab^2nd specimen|Coxsackievirus B6 Ab^2nd specimen
C0881506|T201|COMP|24201-6|LNC|Saint Louis encephalitis virus Ab^1st specimen|Saint Louis encephalitis virus Ab^1st specimen
C0881507|T201|COMP|24202-4|LNC|Saint Louis encephalitis virus Ab^2nd specimen|Saint Louis encephalitis virus Ab^2nd specimen
C0881508|T201|COMP|24203-2|LNC|Legionella pneumophila Ab^1st specimen|Legionella pneumophila Ab^1st specimen
C0881509|T201|COMP|24204-0|LNC|Legionella pneumophila Ab^2nd specimen|Legionella pneumophila Ab^2nd specimen
C0881510|T201|COMP|24205-7|LNC|Rickettsia typhi Ab.IgG^1st specimen|Rickettsia typhi Ab.IgG^1st specimen
C0881511|T201|COMP|24206-5|LNC|Rickettsia typhi Ab.IgG^2nd specimen|Rickettsia typhi Ab.IgG^2nd specimen
C0881514|T201|COMP|24209-9|LNC|La Crosse virus Ab^1st specimen|La Crosse virus Ab^1st specimen
C0881515|T201|COMP|24210-7|LNC|La Crosse virus Ab^2nd specimen|La Crosse virus Ab^2nd specimen
C0881516|T201|COMP|24211-5|LNC|Western equine encephalitis virus Ab^1st specimen|Western equine encephalitis virus Ab^1st specimen
C0881517|T201|COMP|24213-1|LNC|Eastern equine encephalitis virus Ab^1st specimen|Eastern equine encephalitis virus Ab^1st specimen
C0881518|T201|COMP|24214-9|LNC|Eastern equine encephalitis virus Ab^2nd specimen|Eastern equine encephalitis virus Ab^2nd specimen
C0881519|T201|COMP|24215-6|LNC|Influenza virus A Ab^1st specimen|Influenza virus A Ab^1st specimen
C0881520|T201|COMP|24216-4|LNC|Influenza virus A Ab^2nd specimen|Influenza virus A Ab^2nd specimen
C0881521|T201|COMP|24217-2|LNC|Influenza virus B Ab^1st specimen|Influenza virus B Ab^1st specimen
C0881522|T201|COMP|24219-8|LNC|Parainfluenza virus 1 Ab^1st specimen|Parainfluenza virus 1 Ab^1st specimen
C0881523|T201|COMP|24220-6|LNC|Parainfluenza virus 2 Ab^1st specimen|Parainfluenza virus 2 Ab^1st specimen
C0881524|T201|COMP|24221-4|LNC|Parainfluenza virus 2 Ab^2nd specimen|Parainfluenza virus 2 Ab^2nd specimen
C0881525|T201|COMP|24222-2|LNC|Parainfluenza virus 3 Ab^1st specimen|Parainfluenza virus 3 Ab^1st specimen
C0881526|T201|COMP|24224-8|LNC|Respiratory syncytial virus Ab^1st specimen|Respiratory syncytial virus Ab^1st specimen
C0881527|T201|COMP|24225-5|LNC|Respiratory syncytial virus Ab^2nd specimen|Respiratory syncytial virus Ab^2nd specimen
C0881528|T201|COMP|24226-3|LNC|Coxsackievirus A10 Ab^1st specimen|Coxsackievirus A10 Ab^1st specimen
C0881529|T201|COMP|24227-1|LNC|Coxsackievirus A10 Ab^2nd specimen|Coxsackievirus A10 Ab^2nd specimen
C0881530|T201|COMP|24229-7|LNC|Coxsackievirus A16 Ab^2nd specimen|Coxsackievirus A16 Ab^2nd specimen
C0881531|T201|COMP|24231-3|LNC|Coxsackievirus A7 Ab^2nd specimen|Coxsackievirus A7 Ab^2nd specimen
C0881532|T201|COMP|24232-1|LNC|Coxsackievirus A9 Ab^1st specimen|Coxsackievirus A9 Ab^1st specimen
C0881533|T201|COMP|24234-7|LNC|Mycoplasma pneumoniae Ab.IgG^1st specimen|Mycoplasma pneumoniae Ab.IgG^1st specimen
C0881534|T201|COMP|24235-4|LNC|Mycoplasma pneumoniae Ab.IgG^2nd specimen|Mycoplasma pneumoniae Ab.IgG^2nd specimen
C0881535|T201|COMP|24236-2|LNC|Mycoplasma pneumoniae Ab^1st specimen|Mycoplasma pneumoniae Ab^1st specimen
C0881536|T201|COMP|24237-0|LNC|Mycoplasma pneumoniae Ab^2nd specimen|Mycoplasma pneumoniae Ab^2nd specimen
C0881537|T201|COMP|24238-8|LNC|Chlamydia sp Ab.IgG^1st specimen|Chlamydia sp Ab.IgG^1st specimen
C0881538|T201|COMP|24239-6|LNC|Chlamydia sp Ab.IgG^2nd specimen|Chlamydia sp Ab.IgG^2nd specimen
C0881539|T201|COMP|24240-4|LNC|Mumps virus Ab.IgG^1st specimen|Mumps virus Ab.IgG^1st specimen
C0881540|T201|COMP|24241-2|LNC|Mumps virus Ab.IgG^2nd specimen|Mumps virus Ab.IgG^2nd specimen
C0881541|T201|COMP|24242-0|LNC|Toxoplasma gondii Ab.IgG^1st specimen|Toxoplasma gondii Ab.IgG^1st specimen
C0881542|T201|COMP|24243-8|LNC|Polio virus 1 Ab^1st specimen|Polio virus 1 Ab^1st specimen
C0881543|T201|COMP|24244-6|LNC|Polio virus 1 Ab^2nd specimen|Polio virus 1 Ab^2nd specimen
C0881544|T201|COMP|24245-3|LNC|Polio virus 2 Ab^1st specimen|Polio virus 2 Ab^1st specimen
C0881545|T201|COMP|24246-1|LNC|Polio virus 2 Ab^2nd specimen|Polio virus 2 Ab^2nd specimen
C0881546|T201|COMP|24247-9|LNC|Polio virus 3 Ab^1st specimen|Polio virus 3 Ab^1st specimen
C0881547|T201|COMP|24248-7|LNC|Polio virus 3 Ab^2nd specimen|Polio virus 3 Ab^2nd specimen
C0881548|T201|COMP|24249-5|LNC|Adenovirus Ab^1st specimen|Adenovirus Ab^1st specimen
C0881549|T201|COMP|24250-3|LNC|Adenovirus Ab^2nd specimen|Adenovirus Ab^2nd specimen
C0881550|T201|COMP|24251-1|LNC|Coxsackievirus B1 Ab^1st specimen|Coxsackievirus B1 Ab^1st specimen
C0881551|T201|COMP|24252-9|LNC|Coxsackievirus B1 Ab^2nd specimen|Coxsackievirus B1 Ab^2nd specimen
C0881552|T201|COMP|24255-2|LNC|Coxsackievirus B2 Ab^1st specimen|Coxsackievirus B2 Ab^1st specimen
C0881553|T201|COMP|24256-0|LNC|Coxsackievirus B2 Ab^2nd specimen|Coxsackievirus B2 Ab^2nd specimen
C0881554|T201|COMP|24259-4|LNC|Coxsackievirus B3 Ab^1st specimen|Coxsackievirus B3 Ab^1st specimen
C0881555|T201|COMP|24260-2|LNC|Coxsackievirus B3 Ab^2nd specimen|Coxsackievirus B3 Ab^2nd specimen
C0881556|T201|COMP|24263-6|LNC|Coxsackievirus B4 Ab^1st specimen|Coxsackievirus B4 Ab^1st specimen
C0881557|T201|COMP|24264-4|LNC|Coxsackievirus B4 Ab^2nd specimen|Coxsackievirus B4 Ab^2nd specimen
C0881558|T201|COMP|24267-7|LNC|Coxsackievirus B5 Ab^1st specimen|Coxsackievirus B5 Ab^1st specimen
C0881559|T201|COMP|24268-5|LNC|Coxsackievirus B5 Ab^2nd specimen|Coxsackievirus B5 Ab^2nd specimen
C0881560|T201|COMP|24271-9|LNC|Coxsackievirus B6 Ab^1st specimen|Coxsackievirus B6 Ab^1st specimen
C0881561|T201|COMP|24275-0|LNC|Saint Louis encephalitis virus Ab^1st specimen|Saint Louis encephalitis virus Ab^1st specimen
C0881562|T201|COMP|24276-8|LNC|Saint Louis encephalitis virus Ab^2nd specimen|Saint Louis encephalitis virus Ab^2nd specimen
C0881563|T201|COMP|24277-6|LNC|Legionella pneumophila Ab^1st specimen|Legionella pneumophila Ab^1st specimen
C0881564|T201|COMP|24278-4|LNC|Legionella pneumophila Ab^2nd specimen|Legionella pneumophila Ab^2nd specimen
C0881565|T201|COMP|24280-0|LNC|Rickettsia typhi Ab.IgG^2nd specimen|Rickettsia typhi Ab.IgG^2nd specimen
C0881568|T201|COMP|24283-4|LNC|La Crosse virus Ab^1st specimen|La Crosse virus Ab^1st specimen
C0881569|T201|COMP|24285-9|LNC|Western equine encephalitis virus Ab^1st specimen|Western equine encephalitis virus Ab^1st specimen
C0881570|T201|COMP|24286-7|LNC|Western equine encephalitis virus Ab^2nd specimen|Western equine encephalitis virus Ab^2nd specimen
C0881571|T201|COMP|24287-5|LNC|Eastern equine encephalitis virus Ab^1st specimen|Eastern equine encephalitis virus Ab^1st specimen
C0881572|T201|COMP|24288-3|LNC|Eastern equine encephalitis virus Ab^2nd specimen|Eastern equine encephalitis virus Ab^2nd specimen
C0881573|T201|COMP|24290-9|LNC|Influenza virus A Ab^2nd specimen|Influenza virus A Ab^2nd specimen
C0881574|T201|COMP|24291-7|LNC|Influenza virus B Ab^1st specimen|Influenza virus B Ab^1st specimen
C0881575|T201|COMP|24292-5|LNC|Influenza virus B Ab^2nd specimen|Influenza virus B Ab^2nd specimen
C0881576|T201|COMP|24294-1|LNC|Parainfluenza virus 2 Ab^1st specimen|Parainfluenza virus 2 Ab^1st specimen
C0881577|T201|COMP|24295-8|LNC|Parainfluenza virus 2 Ab^2nd specimen|Parainfluenza virus 2 Ab^2nd specimen
C0881578|T201|COMP|24296-6|LNC|Parainfluenza virus 3 Ab^1st specimen|Parainfluenza virus 3 Ab^1st specimen
C0881579|T201|COMP|24297-4|LNC|Parainfluenza virus 3 Ab^2nd specimen|Parainfluenza virus 3 Ab^2nd specimen
C0881580|T201|COMP|24298-2|LNC|Respiratory syncytial virus Ab^1st specimen|Respiratory syncytial virus Ab^1st specimen
C0881581|T201|COMP|24300-6|LNC|Coxsackievirus A10 Ab^1st specimen|Coxsackievirus A10 Ab^1st specimen
C0881582|T201|COMP|24301-4|LNC|Coxsackievirus A10 Ab^2nd specimen|Coxsackievirus A10 Ab^2nd specimen
C0881583|T201|COMP|24302-2|LNC|Coxsackievirus A16 Ab^1st specimen|Coxsackievirus A16 Ab^1st specimen
C0881584|T201|COMP|24304-8|LNC|Coxsackievirus A7 Ab^1st specimen|Coxsackievirus A7 Ab^1st specimen
C0881585|T201|COMP|24305-5|LNC|Coxsackievirus A7 Ab^2nd specimen|Coxsackievirus A7 Ab^2nd specimen
C0881586|T201|COMP|24306-3|LNC|Coxsackievirus A9 Ab^1st specimen|Coxsackievirus A9 Ab^1st specimen
C0881587|T201|COMP|24307-1|LNC|Coxsackievirus A9 Ab^2nd specimen|Coxsackievirus A9 Ab^2nd specimen
C0881588|T201|COMP|24310-5|LNC|Mycoplasma pneumoniae Ab^1st specimen|Mycoplasma pneumoniae Ab^1st specimen
C0881589|T201|COMP|24311-3|LNC|Mycoplasma pneumoniae Ab^2nd specimen|Mycoplasma pneumoniae Ab^2nd specimen
C0881590|T201|COMP|24312-1|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0881591|T201|COMP|24313-9|LNC|Hepatitis 1996 panel|Hepatitis 1996 panel
C0881592|T201|COMP|24314-7|LNC|TORCH 1996 panel|TORCH 1996 panel
C0881593|T201|COMP|24315-4|LNC|Cytomegalovirus Ab.IgG & IgM panel|Cytomegalovirus Ab.IgG & IgM panel
C0881594|T201|COMP|24316-2|LNC|Epstein Barr virus capsid Ab.IgG & IgM panel|Epstein Barr virus capsid Ab.IgG & IgM panel
C0881595|T201|COMP|24317-0|LNC|Hemogram & platelets WO differential panel|Hemogram & platelets WO differential panel
C0881596|T201|COMP|24318-8|LNC|Manual Differential panel|Manual Differential panel
C0881597|T201|COMP|24319-6|LNC|Cardiolipin Ab.IgG & IgM panel|Cardiolipin Ab.IgG & IgM panel
C0881598|T201|COMP|24320-4|LNC|Basic metabolic 1998 panel|Basic metabolic 1998 panel
C0881599|T201|COMP|24321-2|LNC|Basic metabolic 2000 panel|Basic metabolic 2000 panel
C0881600|T201|COMP|24322-0|LNC|Comprehensive metabolic 1998 panel|Comprehensive metabolic 1998 panel
C0881601|T201|COMP|24323-8|LNC|Comprehensive metabolic 2000 panel|Comprehensive metabolic 2000 panel
C0881602|T201|COMP|24324-6|LNC|Hepatic function 1996 panel|Hepatic function 1996 panel
C0881603|T201|COMP|24325-3|LNC|Hepatic function 2000 panel|Hepatic function 2000 panel
C0881604|T201|COMP|24326-1|LNC|Electrolytes 1998 panel|Electrolytes 1998 panel
C0881605|T201|COMP|24327-9|LNC|Electrolytes 3 panel|Electrolytes 3 panel
C0881606|T201|COMP|24328-7|LNC|Electrolytes 3 panel|Electrolytes 3 panel
C0881607|T201|COMP|24329-5|LNC|Electrolytes 3 panel|Electrolytes 3 panel
C0881608|T201|COMP|24331-1|LNC|Lipid 1996 panel|Lipid 1996 panel
C0881609|T201|COMP|24332-9|LNC|Alkaline phosphatase isoenz panel|Alkaline phosphatase isoenz panel
C0881610|T201|COMP|24333-7|LNC|Amylase isoenz 3 panel|Amylase isoenz 3 panel
C0881611|T201|COMP|24334-5|LNC|Amylase isoenz 7 panel|Amylase isoenz 7 panel
C0881612|T201|COMP|24335-2|LNC|Creatine kinase panel|Creatine kinase panel
C0881613|T201|COMP|24337-8|LNC|Gas panel|Gas panel
C0881614|T201|COMP|24339-4|LNC|Gas panel|Gas panel
C0881615|T201|COMP|24340-2|LNC|Gas panel|Gas panel
C0881616|T201|COMP|24342-8|LNC|Gas & CO panel|Gas & CO panel
C0881617|T201|COMP|24343-6|LNC|Gas & CO panel|Gas & CO panel
C0881618|T201|COMP|24344-4|LNC|Gas & CO panel|Gas & CO panel
C0881619|T201|COMP|24346-9|LNC|Parathyrin.intact & Calcium panel|Parathyrin.intact & Calcium panel
C0881620|T201|COMP|24347-7|LNC|Parathyrin.mid molecule & Calcium panel|Parathyrin.mid molecule & Calcium panel
C0881621|T201|COMP|24348-5|LNC|Free T4 & TSH panel|Free T4 & TSH panel
C0881622|T201|COMP|24349-3|LNC|Drugs of abuse 5 panel|Drugs of abuse 5 panel
C0881623|T201|COMP|24350-1|LNC|Volatiles panel|Volatiles panel
C0881624|T201|COMP|24351-9|LNC|Protein fractions panel|Protein fractions panel
C0881625|T201|COMP|24352-7|LNC|Protein fractions panel|Protein fractions panel
C0881626|T201|COMP|24355-0|LNC|Urinalysis macroscopic panel|Urinalysis macroscopic panel
C0881627|T201|COMP|24356-8|LNC|Urinalysis complete panel|Urinalysis complete panel
C0881628|T201|COMP|24357-6|LNC|Urinalysis macro (dipstick) panel|Urinalysis macro (dipstick) panel
C0881629|T201|COMP|24358-4|LNC|Hemogram WO platelets panel|Hemogram WO platelets panel
C0881630|T201|COMP|24360-0|LNC|Hemoglobin & Hematocrit panel|Hemoglobin & Hematocrit panel
C0881631|T201|COMP|24361-8|LNC|Hemogram, platelets & Differential panel|Hemogram, platelets & Differential panel
C0881632|T201|COMP|24362-6|LNC|Renal function 2000 panel|Renal function 2000 panel
C0881633|T201|COMP|24364-2|LNC|Obstetric 1996 panel|Obstetric 1996 panel
C0881634|T201|COMP|24365-9|LNC|Urinalysis microscopic panel|Urinalysis microscopic panel
C0881639|T201|COMP|24373-3|LNC|Ferritin|Ferritin
C0881640|T201|COMP|24374-1|LNC|Platelet associated Ab|Platelet associated Ab
C0881641|T201|COMP|24375-8|LNC|Platelet Ab|Platelet Ab
C0881642|T201|COMP|24376-6|LNC|von Willebrand factor multimers|von Willebrand factor multimers
C0881644|T201|COMP|24378-2|LNC|Platelet aggregation.EPINEPHrine induced|Platelet aggregation.EPINEPHrine induced
C0881645|T201|COMP|24379-0|LNC|Platelet aggregation.collagen induced|Platelet aggregation.collagen induced
C0881646|T201|COMP|24380-8|LNC|Platelet aggregation.ristocetin induced|Platelet aggregation.ristocetin induced
C0881647|T201|COMP|24381-6|LNC|Platelet aggregation.arachidonate induced|Platelet aggregation.arachidonate induced
C0881648|T201|COMP|24382-4|LNC|Neutrophil associated Ab|Neutrophil associated Ab
C0881649|T201|COMP|24383-2|LNC|Intrinsic factor Ab|Intrinsic factor Ab
C0881650|T201|COMP|24384-0|LNC|little c Ab|little c Ab
C0881651|T201|COMP|24386-5|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C0881652|T201|COMP|24387-3|LNC|Brucella sp Ab.IgG|Brucella sp Ab.IgG
C0881653|T201|COMP|24388-1|LNC|Brucella sp Ab.IgM|Brucella sp Ab.IgM
C0881654|T201|COMP|24389-9|LNC|Cortisol^pre 250 ug corticotropin IM|Cortisol^pre 250 ug corticotropin IM
C0881655|T201|COMP|24390-7|LNC|Cortisol^30M post 250 ug corticotropin IM|Cortisol^30M post 250 ug corticotropin IM
C0881656|T201|COMP|24391-5|LNC|Cortisol^1H post 250 ug corticotropin IM|Cortisol^1H post 250 ug corticotropin IM
C0881657|T201|COMP|24392-3|LNC|Cortisol^pre 1 mg dexamethasone PO overnight|Cortisol^pre 1 mg dexamethasone PO overnight
C0881658|T201|COMP|24393-1|LNC|Cortisol^10H post 1 mg dexamethasone PO overnight|Cortisol^10H post 1 mg dexamethasone PO overnight
C0881659|T201|COMP|24394-9|LNC|Cortisol^17H post 1 mg dexamethasone PO overnight|Cortisol^17H post 1 mg dexamethasone PO overnight
C0881660|T201|COMP|24395-6|LNC|Cortisol^24H post 1 mg dexamethasone PO overnight|Cortisol^24H post 1 mg dexamethasone PO overnight
C0881661|T201|COMP|24396-4|LNC|Brucella sp Ab.IgG|Brucella sp Ab.IgG
C0881662|T201|COMP|24397-2|LNC|Brucella sp Ab.IgM|Brucella sp Ab.IgM
C0881663|T201|COMP|24398-0|LNC|Toxoplasma sp Ab.IgM|Toxoplasma sp Ab.IgM
C0881664|T201|COMP|24399-8|LNC|Toxoplasma sp Ab.IgM|Toxoplasma sp Ab.IgM
C0881665|T201|COMP|24400-4|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C0881666|T201|COMP|24401-2|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C0881667|T201|COMP|24403-8|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C0881668|T201|COMP|24404-6|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C0881669|T201|COMP|24405-3|LNC|Aeromonas salmonicida|Aeromonas salmonicida
C0881670|T201|COMP|24406-1|LNC|Aeromonas salmonicida serotype|Aeromonas salmonicida serotype
C0881671|T201|COMP|24407-9|LNC|Androstenedione^baseline|Androstenedione^baseline
C0881672|T201|COMP|24408-7|LNC|Babesia canis|Babesia canis
C0881673|T201|COMP|24410-3|LNC|Brucella canis Ab|Brucella canis Ab
C0881674|T201|COMP|24411-1|LNC|Canine parvovirus Ab|Canine parvovirus Ab
C0881675|T201|COMP|24412-9|LNC|Coccidia identified|Coccidia identified
C0881676|T201|COMP|24415-2|LNC|Feline panleukopenia virus Ag|Feline panleukopenia virus Ag
C0881677|T201|COMP|24416-0|LNC|Filovirus Ab|Filovirus Ab
C0881678|T201|COMP|24417-8|LNC|Follitropin^1st specimen post XXX challenge|Follitropin^1st specimen post XXX challenge
C0881680|T201|COMP|24420-2|LNC|Haemophilus somnus Ab|Haemophilus somnus Ab
C0881681|T201|COMP|24421-0|LNC|Haemobartonella felis|Haemobartonella felis
C0881682|T201|COMP|24427-7|LNC|Mycobacterium avium subspecies paratuberculosis|Mycobacterium avium subspecies paratuberculosis
C0881683|T201|COMP|24428-5|LNC|Mycoplasma hyopneumoniae Ab|Mycoplasma hyopneumoniae Ab
C0881684|T201|COMP|24429-3|LNC|Parasite identified|Parasite identified
C0881685|T201|COMP|24431-9|LNC|IgA.canine|IgA.canine
C0881686|T201|COMP|24432-7|LNC|IgG.canine|IgG.canine
C0881687|T201|COMP|24433-5|LNC|IgG.equine|IgG.equine
C0881688|T201|COMP|24434-3|LNC|IgM.canine|IgM.canine
C0881689|T201|COMP|24435-0|LNC|2-Methylbutyrylglycine/Creatinine|2-Methylbutyrylglycine/Creatinine
C0881690|T201|COMP|24436-8|LNC|3-Methylcrotonylglycine/Creatinine|3-Methylcrotonylglycine/Creatinine
C0881691|T201|COMP|24437-6|LNC|Butyrylglycine/Creatinine|Butyrylglycine/Creatinine
C0881692|T201|COMP|24438-4|LNC|Hexanoylglycine/Creatinine|Hexanoylglycine/Creatinine
C0881693|T201|COMP|24439-2|LNC|Isobutyrylglycine/Creatinine|Isobutyrylglycine/Creatinine
C0881694|T201|COMP|24440-0|LNC|Isovalerylglycine/Creatinine|Isovalerylglycine/Creatinine
C0881695|T201|COMP|24441-8|LNC|Phenylpropionylglycine/Creatinine|Phenylpropionylglycine/Creatinine
C0881696|T201|COMP|24442-6|LNC|Propionylglycine/Creatinine|Propionylglycine/Creatinine
C0881697|T201|COMP|24443-4|LNC|Suberylglycine/Creatinine|Suberylglycine/Creatinine
C0881698|T201|COMP|24444-2|LNC|Tiglylglycine/Creatinine|Tiglylglycine/Creatinine
C0881699|T201|COMP|24445-9|LNC|Valerylglycine/Creatinine|Valerylglycine/Creatinine
C0881700|T201|COMP|24446-7|LNC|Porphobilinogen|Porphobilinogen
C0881701|T201|COMP|24447-5|LNC|Magnesium|Magnesium
C0881702|T201|COMP|24448-3|LNC|Carnitine|Carnitine
C0881703|T201|COMP|24449-1|LNC|Carnitine esters|Carnitine esters
C0881704|T201|COMP|24451-7|LNC|Carnitine|Carnitine
C0881705|T201|COMP|24452-5|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C0881706|T201|COMP|24453-3|LNC|Carnitine|Carnitine
C0881707|T201|COMP|24454-1|LNC|Collection duration|Collection duration
C0881708|T201|COMP|24456-6|LNC|Deoxypyridinoline/Creatinine|Deoxypyridinoline/Creatinine
C0881709|T201|COMP|20659-9|LNC|Tryptophan|Tryptophan
C0881710|T201|COMP|24458-2|LNC|Interleukin 2 receptor|Interleukin 2 receptor
C0881711|T201|COMP|24459-0|LNC|Thyrotropin^20M post dose TRH|Thyrotropin^20M post dose TRH
C0881712|T201|COMP|24461-6|LNC|Fatty acids|Fatty acids
C0881713|T201|COMP|24462-4|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C0881714|T201|COMP|24463-2|LNC|Keratan sulfate|Keratan sulfate
C0881715|T201|COMP|24464-0|LNC|Chondroitin sulfate|Chondroitin sulfate
C0881716|T201|COMP|21166-4|LNC|Cells.CD56/100 cells|Cells.CD56/100 cells
C0881717|T201|COMP|24467-3|LNC|Cells.CD3+CD4+|Cells.CD3+CD4+
C0881718|T201|COMP|24468-1|LNC|Cells.CD14+CD16+CD59+|Cells.CD14+CD16+CD59+
C0881719|T201|COMP|24469-9|LNC|Hemoglobin XXX/Hemoglobin.total|Hemoglobin XXX/Hemoglobin.total
C0881720|T201|COMP|24470-7|LNC|Hemoglobin A2+XXX/Hemoglobin.total|Hemoglobin A2+XXX/Hemoglobin.total
C0881721|T201|COMP|24471-5|LNC|Platelet function.collagen+EPINEPHrine induced|Platelet function.collagen+EPINEPHrine induced
C0881723|T201|COMP|24474-9|LNC|Cancer associated serum Ag|Cancer associated serum Ag
C0881724|T201|COMP|24475-6|LNC|F2 gene.c.20210G>A|F2 gene.c.20210G>A
C0881725|T201|COMP|24476-4|LNC|F2 gene targeted mutation analysis|F2 gene targeted mutation analysis
C0881726|T201|COMP|24477-2|LNC|F2 gene mutations tested for|F2 gene mutations tested for
C0881743|T201|COMP|24497-0|LNC|Canary serum proteins Ab|Canary serum proteins Ab
C0881744|T201|COMP|24498-8|LNC|Chicken serum Ab|Chicken serum Ab
C0881745|T201|COMP|24499-6|LNC|Cryptostroma corticale Ab|Cryptostroma corticale Ab
C0881746|T201|COMP|24500-1|LNC|Parrot serum Ab|Parrot serum Ab
C0881747|T201|COMP|24501-9|LNC|Parrot droppings Ab|Parrot droppings Ab
C0881748|T201|COMP|24502-7|LNC|Parakeet serum Ab|Parakeet serum Ab
C0881749|T201|COMP|24503-5|LNC|Parakeet droppings Ab|Parakeet droppings Ab
C0881750|T201|COMP|24504-3|LNC|Pullularia sp Ab|Pullularia sp Ab
C0881751|T201|COMP|24505-0|LNC|Pigeon droppings Ab|Pigeon droppings Ab
C0881753|T201|COMP|24507-6|LNC|Aspergillus clavatus Ab|Aspergillus clavatus Ab
C0881754|T201|COMP|24508-4|LNC|Aspergillus nidulans Ab|Aspergillus nidulans Ab
C0881755|T201|COMP|24509-2|LNC|Aspergillus terreus Ab|Aspergillus terreus Ab
C0881756|T201|COMP|24510-0|LNC|Vespa crabro Ab.IgE.RAST class|Vespa crabro Ab.IgE.RAST class
C0881757|T201|COMP|24511-8|LNC|Pascopyrum smithii Ab.IgE|Pascopyrum smithii Ab.IgE
C0881759|T201|COMP|24514-2|LNC|Maple syrup Ab.IgE.RAST class|Maple syrup Ab.IgE.RAST class
C0881761|T201|COMP|24516-7|LNC|Pascopyrum smithii Ab.IgE.RAST class|Pascopyrum smithii Ab.IgE.RAST class
C0881762|T201|COMP|24517-5|LNC|Phoma sp Ab.IgG|Phoma sp Ab.IgG
C0881763|T201|COMP|24518-3|LNC|Calcium/Creatinine|Calcium/Creatinine
C0881764|T201|COMP|24519-1|LNC|Phosphate|Phosphate
C0881765|T201|COMP|24521-7|LNC|EPINEPHrine|EPINEPHrine
C0881766|T201|COMP|24522-5|LNC|EPINEPHrine/Creatinine|EPINEPHrine/Creatinine
C0881767|T201|COMP|24523-3|LNC|Norepinephrine/Creatinine|Norepinephrine/Creatinine
C0881768|T201|COMP|24524-1|LNC|DOPamine/Creatinine|DOPamine/Creatinine
C0882230|T201|COMP|19725-1|LNC|Aspergillus flavus Ab.IgG|Aspergillus flavus Ab.IgG
C0882231|T201|COMP|19738-4|LNC|Dog serum albumin Ab.IgE|Dog serum albumin Ab.IgE
C0882232|T201|COMP|19742-6|LNC|Hexahydrophthalic anhydride Ab.IgE|Hexahydrophthalic anhydride Ab.IgE
C0882233|T201|COMP|22079-8|LNC|Actinomyces sp Ab|Actinomyces sp Ab
C0882234|T201|COMP|22083-0|LNC|Alcelaphine herpesvirus 1 Ab|Alcelaphine herpesvirus 1 Ab
C0882235|T201|COMP|22088-9|LNC|Avian adenovirus 2 Ab|Avian adenovirus 2 Ab
C0882236|T201|COMP|22090-5|LNC|Avian encephalomyelitis virus Ab|Avian encephalomyelitis virus Ab
C0882237|T201|COMP|22092-1|LNC|Infectious bronchitis virus Ark-99 Ab|Infectious bronchitis virus Ark-99 Ab
C0882238|T201|COMP|22095-4|LNC|Avian infectious laryngotracheitis virus Ab|Avian infectious laryngotracheitis virus Ab
C0882239|T201|COMP|22125-9|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0882240|T201|COMP|22128-3|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0882241|T201|COMP|22133-3|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0882242|T201|COMP|22138-2|LNC|Borrelia hermsii Ab.IgG|Borrelia hermsii Ab.IgG
C0882243|T201|COMP|22142-4|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C0882244|T201|COMP|22147-3|LNC|Brucella abortus Ab|Brucella abortus Ab
C0882245|T201|COMP|22151-5|LNC|Brucella abortus Ab.IgM|Brucella abortus Ab.IgM
C0882246|T201|COMP|22179-6|LNC|Chlamydophila psittaci Ab.IgG|Chlamydophila psittaci Ab.IgG
C0882247|T201|COMP|22187-9|LNC|Chlamydia trachomatis Ab|Chlamydia trachomatis Ab
C0882248|T201|COMP|22191-1|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C0882249|T201|COMP|22196-0|LNC|Chlamydia trachomatis B Ab.IgM|Chlamydia trachomatis B Ab.IgM
C0882250|T201|COMP|22203-4|LNC|Clostridium tetani Ab.IgG|Clostridium tetani Ab.IgG
C0882251|T201|COMP|22208-3|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0882252|T201|COMP|22211-7|LNC|Coxiella burnetii Ab|Coxiella burnetii Ab
C0882253|T201|COMP|22212-5|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C0882254|T201|COMP|22217-4|LNC|Coxsackievirus A21 Ab|Coxsackievirus A21 Ab
C0882255|T201|COMP|22237-2|LNC|Cryptococcus neoformans Ab|Cryptococcus neoformans Ab
C0882256|T201|COMP|22255-4|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C0882257|T201|COMP|22264-6|LNC|Echinococcus granulosus Ab.IgG|Echinococcus granulosus Ab.IgG
C0882258|T201|COMP|22269-5|LNC|Echovirus 14 Ab|Echovirus 14 Ab
C0882259|T201|COMP|22273-7|LNC|Echovirus 19 Ab|Echovirus 19 Ab
C0882260|T201|COMP|22281-0|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C0882261|T201|COMP|22293-5|LNC|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C0882262|T201|COMP|22312-3|LNC|Hepatitis A virus Ab|Hepatitis A virus Ab
C0882263|T201|COMP|22317-2|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C0882264|T201|COMP|22321-4|LNC|Hepatitis B virus little e Ab|Hepatitis B virus little e Ab
C0882265|T201|COMP|22324-8|LNC|Hepatitis C virus 100-3 Ab|Hepatitis C virus 100-3 Ab
C0882266|T201|COMP|22331-3|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C0882267|T201|COMP|22340-4|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C0882268|T201|COMP|22349-5|LNC|Histoplasma capsulatum Ab.IgA|Histoplasma capsulatum Ab.IgA
C0882269|T201|COMP|17038-1|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C0882270|T201|COMP|22378-4|LNC|Lassa virus Ab.IgG|Lassa virus Ab.IgG
C0882271|T201|COMP|22382-6|LNC|Legionella pneumophila 1 Ab.IgM|Legionella pneumophila 1 Ab.IgM
C0882272|T201|COMP|22387-5|LNC|Legionella pneumophila 4 Ab.IgG|Legionella pneumophila 4 Ab.IgG
C0882273|T201|COMP|22392-5|LNC|Legionella pneumophila 6 Ab.IgM|Legionella pneumophila 6 Ab.IgM
C0882274|T201|COMP|22400-6|LNC|Leptospira interrogans serovar Bratislava Ab|Leptospira interrogans serovar Bratislava Ab
C0882275|T201|COMP|22409-7|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C0882276|T201|COMP|22437-8|LNC|Parainfluenza virus 1 Ab|Parainfluenza virus 1 Ab
C0882277|T201|COMP|22441-0|LNC|Plasmodium falciparum Ab|Plasmodium falciparum Ab
C0882278|T201|COMP|22442-8|LNC|Plasmodium malariae Ab|Plasmodium malariae Ab
C0882279|T201|COMP|22446-9|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C0882280|T201|COMP|22450-1|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C0882281|T201|COMP|22454-3|LNC|Pseudorabies virus.ClinEase gene deletion Ab|Pseudorabies virus.ClinEase gene deletion Ab
C0882282|T201|COMP|22464-2|LNC|Reagin Ab|Reagin Ab
C0882283|T201|COMP|22480-8|LNC|Rickettsia typhus group Ab.IgG|Rickettsia typhus group Ab.IgG
C0882284|T201|COMP|22499-8|LNC|Measles virus Ab|Measles virus Ab
C0882285|T201|COMP|22502-9|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0882286|T201|COMP|22506-0|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C0882287|T201|COMP|22510-2|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C0882288|T201|COMP|22516-9|LNC|Salmonella paratyphi A Ab|Salmonella paratyphi A Ab
C0882289|T201|COMP|22517-7|LNC|Salmonella paratyphi A H Ab|Salmonella paratyphi A H Ab
C0882290|T201|COMP|22520-1|LNC|Salmonella paratyphi B Ab|Salmonella paratyphi B Ab
C0882291|T201|COMP|22525-0|LNC|Salmonella paratyphi C O Ab|Salmonella paratyphi C O Ab
C0882292|T201|COMP|22534-2|LNC|Sarcocystis neurona Ab|Sarcocystis neurona Ab
C0882294|T201|COMP|22564-9|LNC|Streptococcus pneumoniae Ab.IgG^2nd specimen|Streptococcus pneumoniae Ab.IgG^2nd specimen
C0882295|T201|COMP|22570-6|LNC|Taenia solium Ab|Taenia solium Ab
C0882296|T201|COMP|22575-5|LNC|Toxocara canis Ab.IgG|Toxocara canis Ab.IgG
C0882297|T201|COMP|22583-9|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0882298|T201|COMP|22596-1|LNC|Trichinella spiralis Ab|Trichinella spiralis Ab
C0882299|T201|COMP|22618-3|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C0882300|T201|COMP|22625-8|LNC|Xylose^2H post dose xylose PO|Xylose^2H post dose xylose PO
C0882301|T201|COMP|22631-6|LNC|Xylose/Xylose.dose^post 5 g xylose PO|Xylose/Xylose.dose^post 5 g xylose PO
C0882304|T201|COMP|22645-6|LNC|Proline|Proline
C0882305|T201|COMP|22664-7|LNC|Urea|Urea
C0882306|T201|COMP|22680-3|LNC|Mercury/Creatinine|Mercury/Creatinine
C0882307|T201|COMP|22684-5|LNC|Serine/Creatinine|Serine/Creatinine
C0882308|T201|COMP|22689-4|LNC|Zinc|Zinc
C0882309|T201|COMP|22690-2|LNC|Proline/Creatinine|Proline/Creatinine
C0882310|T201|COMP|22692-8|LNC|Valine/Creatinine|Valine/Creatinine
C0882311|T201|COMP|22697-7|LNC|Arginine/Creatinine|Arginine/Creatinine
C0882312|T201|COMP|22708-2|LNC|Homovanillate/Creatinine|Homovanillate/Creatinine
C0882313|T201|COMP|22712-4|LNC|Adenosine monophosphate.cyclic|Adenosine monophosphate.cyclic
C0882314|T201|COMP|22726-4|LNC|Creatinine|Creatinine
C0882315|T201|COMP|22747-0|LNC|Gentamicin^trough|Gentamicin^trough
C0882316|T201|COMP|22751-2|LNC|Tobramycin^peak|Tobramycin^peak
C0882317|T201|COMP|22752-0|LNC|Tobramycin^trough|Tobramycin^trough
C0882318|T201|COMP|22755-3|LNC|Haemophilus influenzae B Ab|Haemophilus influenzae B Ab
C0882319|T201|COMP|22760-3|LNC|Potassium|Potassium
C0882320|T201|COMP|22764-5|LNC|Actinobacillus pleuropneumoniae Ab|Actinobacillus pleuropneumoniae Ab
C0882321|T201|COMP|22773-6|LNC|African horse sickness virus Ag|African horse sickness virus Ag
C0882322|T201|COMP|22778-5|LNC|African swine fever virus Ab|African swine fever virus Ab
C0882323|T201|COMP|22791-8|LNC|Alcelaphine herpesvirus 1 DNA|Alcelaphine herpesvirus 1 DNA
C0882324|T201|COMP|22814-8|LNC|Avian infectious laryngotracheitis virus Ab|Avian infectious laryngotracheitis virus Ab
C0882325|T201|COMP|22819-7|LNC|Avian infectious laryngotracheitis virus Ag|Avian infectious laryngotracheitis virus Ag
C0882326|T201|COMP|22824-7|LNC|Influenza virus A Ab|Influenza virus A Ab
C0882327|T201|COMP|22826-2|LNC|Influenza virus A identified|Influenza virus A identified
C0882328|T201|COMP|22829-6|LNC|Avian paramyxovirus 1 Ab|Avian paramyxovirus 1 Ab
C0882329|T201|COMP|22834-6|LNC|Avian metapneumovirus Ab|Avian metapneumovirus Ab
C0882330|T201|COMP|22844-5|LNC|Babesia bigemina Ab|Babesia bigemina Ab
C0882331|T201|COMP|22868-4|LNC|Bluetongue virus Ab|Bluetongue virus Ab
C0882332|T201|COMP|22872-6|LNC|Bluetongue virus Ag|Bluetongue virus Ag
C0882333|T201|COMP|22873-4|LNC|Bluetongue virus Ag|Bluetongue virus Ag
C0882334|T201|COMP|22877-5|LNC|Border disease virus Ab|Border disease virus Ab
C0882335|T201|COMP|22881-7|LNC|Border disease virus Ag|Border disease virus Ag
C0882336|T201|COMP|22886-6|LNC|Bordetella bronchiseptica Ab|Bordetella bronchiseptica Ab
C0882337|T201|COMP|22890-8|LNC|Bovine diarrhea virus Ab|Bovine diarrhea virus Ab
C0882338|T201|COMP|22895-7|LNC|Bovine diarrhea virus Ab|Bovine diarrhea virus Ab
C0882339|T201|COMP|22924-5|LNC|Brucella abortus Ab.IgG1|Brucella abortus Ab.IgG1
C0882340|T201|COMP|22932-8|LNC|Brucella melitensis Ab|Brucella melitensis Ab
C0882341|T201|COMP|22937-7|LNC|Brucella ovis Ab|Brucella ovis Ab
C0882342|T201|COMP|22940-1|LNC|Brucella ovis Ab|Brucella ovis Ab
C0882343|T201|COMP|22945-0|LNC|Brucella sp Ag|Brucella sp Ag
C0882344|T201|COMP|22953-4|LNC|Brucella suis Ab|Brucella suis Ab
C0882345|T201|COMP|22956-7|LNC|Burkholderia mallei Ab|Burkholderia mallei Ab
C0882346|T201|COMP|22958-3|LNC|Burkholderia mallei Ab|Burkholderia mallei Ab
C0882347|T201|COMP|22969-0|LNC|Campylobacter fetus subspecies venerealis Ab.IgA|Campylobacter fetus subspecies venerealis Ab.IgA
C0882348|T201|COMP|22992-2|LNC|Chlamydophila psittaci|Chlamydophila psittaci
C0882349|T201|COMP|22998-9|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C0882350|T201|COMP|23000-3|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C0882351|T201|COMP|23004-5|LNC|Classical swine fever virus Ab|Classical swine fever virus Ab
C0882352|T201|COMP|23006-0|LNC|Classical swine fever virus Ag|Classical swine fever virus Ag
C0882353|T201|COMP|23010-2|LNC|Cowdria ruminantium Ab|Cowdria ruminantium Ab
C0882354|T201|COMP|23018-5|LNC|Coxiella burnetii Ab|Coxiella burnetii Ab
C0882355|T201|COMP|23046-6|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C0882356|T201|COMP|23047-4|LNC|Eastern equine encephalitis virus Ag|Eastern equine encephalitis virus Ag
C0882357|T201|COMP|23052-4|LNC|Eastern equine encephalitis virus RNA|Eastern equine encephalitis virus RNA
C0882358|T201|COMP|23058-1|LNC|Ephemeral fever virus Ab|Ephemeral fever virus Ab
C0882359|T201|COMP|23062-3|LNC|Epizootic hemorrhagic disease virus Ag|Epizootic hemorrhagic disease virus Ag
C0882360|T201|COMP|23067-2|LNC|Epizootic hemorrhagic disease virus RNA|Epizootic hemorrhagic disease virus RNA
C0882361|T201|COMP|23074-8|LNC|Equine arteritis virus Ag|Equine arteritis virus Ag
C0882362|T201|COMP|23102-7|LNC|Equine influenza virus A1 Ag|Equine influenza virus A1 Ag
C0882363|T201|COMP|23105-0|LNC|Fly larvae identified|Fly larvae identified
C0882364|T201|COMP|23114-2|LNC|Foot and mouth disease virus RNA|Foot and mouth disease virus RNA
C0882365|T201|COMP|23123-3|LNC|Francisella tularensis A rRNA|Francisella tularensis A rRNA
C0882367|T201|COMP|23163-9|LNC|Leptospira interrogans serovar Australis Ab|Leptospira interrogans serovar Australis Ab
C0882368|T201|COMP|23169-6|LNC|Leptospira interrogans serovar Bataviae Ab|Leptospira interrogans serovar Bataviae Ab
C0882369|T201|COMP|23172-0|LNC|Leptospira interrogans serovar Bratislava Ab|Leptospira interrogans serovar Bratislava Ab
C0882370|T201|COMP|23174-6|LNC|Leptospira interrogans serovar Canicola Ab|Leptospira interrogans serovar Canicola Ab
C0882371|T201|COMP|23214-0|LNC|Lumpy skin disease virus Ab|Lumpy skin disease virus Ab
C0882372|T201|COMP|23219-9|LNC|Lumpy skin disease virus Ag|Lumpy skin disease virus Ag
C0882373|T201|COMP|23224-9|LNC|Mareks disease virus Ab|Mareks disease virus Ab
C0882374|T201|COMP|23227-2|LNC|Mareks disease virus Ab|Mareks disease virus Ab
C0882375|T201|COMP|23228-0|LNC|Mareks disease virus Ab|Mareks disease virus Ab
C0882376|T201|COMP|23233-0|LNC|Mite identified|Mite identified
C0882377|T201|COMP|23238-9|LNC|Mycobacterium avium subspecies avium serotype|Mycobacterium avium subspecies avium serotype
C0882378|T201|COMP|23255-3|LNC|Mycoplasma bovis Ab|Mycoplasma bovis Ab
C0882379|T201|COMP|23274-4|LNC|Mycoplasma gallisepticum Ab|Mycoplasma gallisepticum Ab
C0882382|T201|COMP|23328-8|LNC|Ovine progressive pneumonia virus Ab|Ovine progressive pneumonia virus Ab
C0882383|T201|COMP|23333-8|LNC|Ovine progressive pneumonia virus Ab|Ovine progressive pneumonia virus Ab
C0882384|T201|COMP|23338-7|LNC|Ovine pulmonary adenomatosis retrovirus RNA|Ovine pulmonary adenomatosis retrovirus RNA
C0882385|T201|COMP|23344-5|LNC|Pasteurella multocida rRNA|Pasteurella multocida rRNA
C0882386|T201|COMP|23349-4|LNC|Pasteurella multocida toxin|Pasteurella multocida toxin
C0882387|T201|COMP|23373-4|LNC|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C0882388|T201|COMP|23382-5|LNC|Pseudorabies virus Ab|Pseudorabies virus Ab
C0882389|T201|COMP|23387-4|LNC|Pseudorabies virus DNA|Pseudorabies virus DNA
C0882390|T201|COMP|23392-4|LNC|Rabies virus DNA|Rabies virus DNA
C0882391|T201|COMP|23397-3|LNC|Rift valley fever virus Ab|Rift valley fever virus Ab
C0882392|T201|COMP|23400-5|LNC|Rift valley fever virus Ab|Rift valley fever virus Ab
C0882393|T201|COMP|23405-4|LNC|Rift valley fever virus Ag|Rift valley fever virus Ag
C0882394|T201|COMP|23443-5|LNC|Swine vesicular disease virus Ab|Swine vesicular disease virus Ab
C0882395|T201|COMP|23449-2|LNC|Taenia hydatigena Ag|Taenia hydatigena Ag
C0882396|T201|COMP|23452-6|LNC|Taenia sp eggs|Taenia sp eggs
C0882397|T201|COMP|23453-4|LNC|Taylorella equigenitalis Ab|Taylorella equigenitalis Ab
C0882398|T201|COMP|23458-3|LNC|Taylorella equigenitalis DNA|Taylorella equigenitalis DNA
C0882399|T201|COMP|23463-3|LNC|Theileria annulata rRNA|Theileria annulata rRNA
C0882400|T201|COMP|23491-4|LNC|Transmissible gastroenteritis virus Ab|Transmissible gastroenteritis virus Ab
C0882401|T201|COMP|23496-3|LNC|Transmissible gastroenteritis virus Ag|Transmissible gastroenteritis virus Ag
C0882402|T201|COMP|23500-2|LNC|Tritrichomonas foetus Ab|Tritrichomonas foetus Ab
C0882403|T201|COMP|23505-1|LNC|Tritrichomonas foetus DNA|Tritrichomonas foetus DNA
C0882404|T201|COMP|23510-1|LNC|Trypanosoma equiperdum Ab|Trypanosoma equiperdum Ab
C0882405|T201|COMP|23524-2|LNC|Trypanosoma evansi Ab|Trypanosoma evansi Ab
C0882406|T201|COMP|23557-2|LNC|Vesicular stomatitis virus Ag|Vesicular stomatitis virus Ag
C0882407|T201|COMP|23562-2|LNC|Vesicular stomatitis Indiana virus Ab|Vesicular stomatitis Indiana virus Ab
C0882408|T201|COMP|23567-1|LNC|Vesicular stomatitis New Jersey virus Ab|Vesicular stomatitis New Jersey virus Ab
C0882409|T201|COMP|23569-7|LNC|Vesicular stomatitis virus serotype|Vesicular stomatitis virus serotype
C0882410|T201|COMP|23572-1|LNC|Vesicular stomatitis virus serotype|Vesicular stomatitis virus serotype
C0882411|T201|COMP|23578-8|LNC|Viral hemorrhagic disease virus Ab|Viral hemorrhagic disease virus Ab
C0882412|T201|COMP|23611-7|LNC|Para aminosalicylate|Para aminosalicylate
C0882413|T201|COMP|23617-4|LNC|Ethionamide|Ethionamide
C0882414|T201|COMP|23620-8|LNC|Clofazimine|Clofazimine
C0882415|T201|COMP|23625-7|LNC|Ethambutol|Ethambutol
C0882416|T201|COMP|23633-1|LNC|Erythromycin|Erythromycin
C0882417|T201|COMP|23635-6|LNC|Erythropoietin given|Erythropoietin given
C0882418|T201|COMP|23638-0|LNC|Grepafloxacin|Grepafloxacin
C0882419|T201|COMP|23649-7|LNC|Actinobacillus pleuropneumoniae biovar 2 serotype|Actinobacillus pleuropneumoniae biovar 2 serotype
C0882420|T201|COMP|23674-5|LNC|Bluetongue virus 17 Ab|Bluetongue virus 17 Ab
C0882421|T201|COMP|23684-4|LNC|Brucella ovis Ab|Brucella ovis Ab
C0882422|T201|COMP|23687-7|LNC|Canine coronavirus Ab|Canine coronavirus Ab
C0882423|T201|COMP|23688-5|LNC|Canine coronavirus Ag|Canine coronavirus Ag
C0882424|T201|COMP|23692-7|LNC|Canine distemper virus Ab.IgG|Canine distemper virus Ab.IgG
C0882425|T201|COMP|23697-6|LNC|Canine herpesvirus Ab|Canine herpesvirus Ab
C0882426|T201|COMP|23709-9|LNC|Ceftiofur|Ceftiofur
C0882427|T201|COMP|23732-1|LNC|Feline leukemia virus Ab|Feline leukemia virus Ab
C0882428|T201|COMP|23735-4|LNC|Feline leukemia virus Ab|Feline leukemia virus Ab
C0882429|T201|COMP|23738-8|LNC|Feline herpesvirus 1 Ab|Feline herpesvirus 1 Ab
C0882430|T201|COMP|23742-0|LNC|Fumonisin|Fumonisin
C0882431|T201|COMP|23746-1|LNC|Gossypol.free|Gossypol.free
C0882432|T201|COMP|23750-3|LNC|Leptospira sp Ag|Leptospira sp Ag
C0882433|T201|COMP|23759-4|LNC|Neospora caninum Ag|Neospora caninum Ag
C0882434|T201|COMP|23771-9|LNC|Porcine parvovirus Ag|Porcine parvovirus Ag
C0882437|T201|COMP|23814-7|LNC|Amantadine|Amantadine
C0882438|T201|COMP|23818-8|LNC|Antibiotic XXX^trough|Antibiotic XXX^trough
C0882439|T201|COMP|23848-5|LNC|Creosol|Creosol
C0882440|T201|COMP|23849-3|LNC|Creosol|Creosol
C0882441|T201|COMP|23851-9|LNC|Cyclohexanone|Cyclohexanone
C0882442|T201|COMP|23856-8|LNC|Endrin|Endrin
C0882443|T201|COMP|23863-4|LNC|Finch droppings Ab.IgE.RAST class|Finch droppings Ab.IgE.RAST class
C0882444|T201|COMP|23869-1|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C0882445|T201|COMP|23873-3|LNC|Heptacarboxylporphyrin III|Heptacarboxylporphyrin III
C0882446|T201|COMP|23890-7|LNC|Lead|Lead
C0882448|T201|COMP|23915-2|LNC|Osmotic fragility^0.50% sodium chloride|Osmotic fragility^0.50% sodium chloride
C0882450|T201|COMP|23923-6|LNC|Parakeet droppings Ab.IgE.RAST class|Parakeet droppings Ab.IgE.RAST class
C0882451|T201|COMP|23929-3|LNC|Ribonucleoprotein extractable nuclear Ab.IgG|Ribonucleoprotein extractable nuclear Ab.IgG
C0882452|T201|COMP|23933-5|LNC|Staphylococcus aureus enterotoxin B|Staphylococcus aureus enterotoxin B
C0882453|T201|COMP|23965-7|LNC|Burkholderia pseudomallei Ab.IgG|Burkholderia pseudomallei Ab.IgG
C0882454|T201|COMP|23974-9|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C0882455|T201|COMP|23979-8|LNC|Borrelia burgdorferi Ab.IgG band pattern|Borrelia burgdorferi Ab.IgG band pattern
C0882456|T201|COMP|23984-8|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0882457|T201|COMP|23993-9|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C0882459|T201|COMP|24043-2|LNC|Acetyl-CoA:glucosamine acetyltransferase|Acetyl-CoA:glucosamine acetyltransferase
C0882460|T201|COMP|24048-1|LNC|Alpha galactosidase A|Alpha galactosidase A
C0882461|T201|COMP|24049-9|LNC|Alpha galactosidase A|Alpha galactosidase A
C0882462|T201|COMP|24052-3|LNC|Alpha mannosidase|Alpha mannosidase
C0882463|T201|COMP|24057-2|LNC|Alpha-L-iduronidase|Alpha-L-iduronidase
C0882464|T201|COMP|24065-5|LNC|Beta glucuronidase|Beta glucuronidase
C0882465|T201|COMP|24091-1|LNC|Alpha-N-acetylglucosaminidase|Alpha-N-acetylglucosaminidase
C0882466|T201|COMP|24092-9|LNC|Alpha-N-acetylglucosaminidase|Alpha-N-acetylglucosaminidase
C0882467|T201|COMP|24096-0|LNC|N-Acetylgalactosamine-6-Sulfatase|N-Acetylgalactosamine-6-Sulfatase
C0882468|T201|COMP|24103-4|LNC|Plasma cells|Plasma cells
C0882469|T201|COMP|24108-3|LNC|Cancer Ag 19-9|Cancer Ag 19-9
C0882470|T201|COMP|24112-5|LNC|Trichomonas vaginalis rRNA|Trichomonas vaginalis rRNA
C0882471|T201|COMP|24117-4|LNC|Ross river virus Ab.IgG|Ross river virus Ab.IgG
C0882472|T201|COMP|24140-6|LNC|Fraxinus americana Ab.IgG|Fraxinus americana Ab.IgG
C0882473|T201|COMP|24155-4|LNC|Mangifera indica Ab.IgG|Mangifera indica Ab.IgG
C0882474|T201|COMP|24159-6|LNC|Pepper white+Pepper black Ab.IgE|Pepper white+Pepper black Ab.IgE
C0882475|T201|COMP|24163-8|LNC|(Beef+Chicken+Pork) Ab.IgE|(Beef+Chicken+Pork) Ab.IgE
C0882476|T201|COMP|24169-5|LNC|Polio virus 1 Ab^1st specimen|Polio virus 1 Ab^1st specimen
C0882477|T201|COMP|24173-7|LNC|Polio virus 3 Ab^1st specimen|Polio virus 3 Ab^1st specimen
C0882478|T201|COMP|24179-4|LNC|Coxsackievirus B1 Ab^1st specimen|Coxsackievirus B1 Ab^1st specimen
C0882479|T201|COMP|24212-3|LNC|Western equine encephalitis virus Ab^2nd specimen|Western equine encephalitis virus Ab^2nd specimen
C0882480|T201|COMP|24218-0|LNC|Influenza virus B Ab^2nd specimen|Influenza virus B Ab^2nd specimen
C0882481|T201|COMP|24223-0|LNC|Parainfluenza virus 3 Ab^2nd specimen|Parainfluenza virus 3 Ab^2nd specimen
C0882482|T201|COMP|24228-9|LNC|Coxsackievirus A16 Ab^1st specimen|Coxsackievirus A16 Ab^1st specimen
C0882483|T201|COMP|24230-5|LNC|Coxsackievirus A7 Ab^1st specimen|Coxsackievirus A7 Ab^1st specimen
C0882484|T201|COMP|24233-9|LNC|Coxsackievirus A9 Ab^2nd specimen|Coxsackievirus A9 Ab^2nd specimen
C0882485|T201|COMP|24272-7|LNC|Coxsackievirus B6 Ab^2nd specimen|Coxsackievirus B6 Ab^2nd specimen
C0882486|T201|COMP|24279-2|LNC|Rickettsia typhi Ab.IgG^1st specimen|Rickettsia typhi Ab.IgG^1st specimen
C0882487|T201|COMP|24284-2|LNC|La Crosse virus Ab^2nd specimen|La Crosse virus Ab^2nd specimen
C0882488|T201|COMP|24289-1|LNC|Influenza virus A Ab^1st specimen|Influenza virus A Ab^1st specimen
C0882489|T201|COMP|24293-3|LNC|Parainfluenza virus 1 Ab^1st specimen|Parainfluenza virus 1 Ab^1st specimen
C0882490|T201|COMP|24299-0|LNC|Respiratory syncytial virus Ab^2nd specimen|Respiratory syncytial virus Ab^2nd specimen
C0882491|T201|COMP|24303-0|LNC|Coxsackievirus A16 Ab^2nd specimen|Coxsackievirus A16 Ab^2nd specimen
C0882492|T201|COMP|24336-0|LNC|Gas panel|Gas panel
C0882493|T201|COMP|24338-6|LNC|Gas panel|Gas panel
C0882494|T201|COMP|24341-0|LNC|Gas & CO panel|Gas & CO panel
C0882495|T201|COMP|24345-1|LNC|Gas & CO panel|Gas & CO panel
C0882496|T201|COMP|24353-5|LNC|Glucose tolerance 2H gestational panel|Glucose tolerance 2H gestational panel
C0882498|T201|COMP|24385-7|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C0882500|T201|COMP|24413-7|LNC|Eperythrozoon sp|Eperythrozoon sp
C0882501|T201|COMP|24414-5|LNC|Estradiol^baseline|Estradiol^baseline
C0882502|T201|COMP|24418-6|LNC|Formononetin|Formononetin
C0882503|T201|COMP|24422-8|LNC|Hydrocarbons.chlorinated|Hydrocarbons.chlorinated
C0882504|T201|COMP|24430-1|LNC|Streptococcus suis serotype|Streptococcus suis serotype
C0882505|T201|COMP|24450-9|LNC|Carnitine esters|Carnitine esters
C0882506|T201|COMP|24465-7|LNC|Urea nitrogen|Urea nitrogen
C0882507|T201|COMP|19078-5|LNC|Cells.CD23/100 cells|Cells.CD23/100 cells
C0882512|T201|COMP|24520-9|LNC|Phosphate|Phosphate
C0884099|T201|COMP|22250-5|LNC|Dengue virus 1 Ab|Dengue virus 1 Ab
C0884100|T201|COMP|22277-8|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C0884101|T201|COMP|22326-3|LNC|Hepatitis C virus 5-1-1 Ab|Hepatitis C virus 5-1-1 Ab
C0884102|T201|COMP|22397-4|LNC|Legionella pneumophila Ab.IgG|Legionella pneumophila Ab.IgG
C0884103|T201|COMP|22627-4|LNC|Xylose^post 5 g xylose PO|Xylose^post 5 g xylose PO
C0884104|T201|COMP|22704-1|LNC|Carnitine.free (C0)/Creatinine|Carnitine.free (C0)/Creatinine
C0884105|T201|COMP|23321-3|LNC|Ovine herpesvirus 2 Ab|Ovine herpesvirus 2 Ab
C0884106|T201|COMP|23754-5|LNC|Mycoplasma sp Ab|Mycoplasma sp Ab
C0884107|T201|COMP|23912-9|LNC|Osmotic fragility^0.35% sodium chloride|Osmotic fragility^0.35% sodium chloride
C0884108|T201|COMP|23989-7|LNC|Burkholderia pseudomallei Ab.IgM|Burkholderia pseudomallei Ab.IgM
C0884109|T201|COMP|24363-4|LNC|Acute hepatitis 2000 panel|Acute hepatitis 2000 panel
C0884110|T201|COMP|24409-5|LNC|Brachyspira sp identified|Brachyspira sp identified
C0884313|T201|COMP|23420-3|LNC|Salmonella abortus ovis Ab|Salmonella abortus ovis Ab
C0884314|T201|COMP|24011-9|LNC|Hepatitis C virus Ab band pattern|Hepatitis C virus Ab band pattern
C0941291|T201|COMP|18474-7|LNC|HER2 Ag|HER2 Ag
C0941292|T201|COMP|25082-9|LNC|2-Methyl-3-Hydroxybutyrate/Creatinine|2-Methyl-3-Hydroxybutyrate/Creatinine
C0941293|T201|COMP|25083-7|LNC|2-Oxo,3-Methylvalerate/Creatinine|2-Oxo,3-Methylvalerate/Creatinine
C0941294|T201|COMP|25084-5|LNC|2-Oxoisocaproate/Creatinine|2-Oxoisocaproate/Creatinine
C0941295|T201|COMP|25085-2|LNC|2-Oxoisovalerate/Creatinine|2-Oxoisovalerate/Creatinine
C0941296|T201|COMP|25086-0|LNC|Beta aminoisobutyrate/Creatinine|Beta aminoisobutyrate/Creatinine
C0941297|T201|COMP|25087-8|LNC|3-Methylglutaconate/Creatinine|3-Methylglutaconate/Creatinine
C0941298|T201|COMP|25089-4|LNC|4-Hydroxyphenyllactate/Creatinine|4-Hydroxyphenyllactate/Creatinine
C0941299|T201|COMP|25091-0|LNC|C peptide/Creatinine|C peptide/Creatinine
C0941300|T201|COMP|25092-8|LNC|Cystathionine/Creatinine|Cystathionine/Creatinine
C0941301|T201|COMP|25093-6|LNC|Decadienediate/Creatinine|Decadienediate/Creatinine
C0941302|T201|COMP|25094-4|LNC|Decenedioate/Creatinine|Decenedioate/Creatinine
C0941303|T201|COMP|25095-1|LNC|Deoxypyridinoline/Creatinine|Deoxypyridinoline/Creatinine
C0941304|T201|COMP|25096-9|LNC|Deoxypyridinoline/Creatinine|Deoxypyridinoline/Creatinine
C0941305|T201|COMP|25097-7|LNC|Dodecanedioate/Creatinine|Dodecanedioate/Creatinine
C0941306|T201|COMP|25098-5|LNC|Ethanolamine/Creatinine|Ethanolamine/Creatinine
C0941307|T201|COMP|25099-3|LNC|Ethylmalonate/Creatinine|Ethylmalonate/Creatinine
C0941308|T201|COMP|25100-9|LNC|Formate/Creatinine|Formate/Creatinine
C0941309|T201|COMP|25101-7|LNC|Fumarate/Creatinine|Fumarate/Creatinine
C0941310|T201|COMP|25102-5|LNC|Galactose/Creatinine|Galactose/Creatinine
C0941311|T201|COMP|25103-3|LNC|Glutaconate/Creatinine|Glutaconate/Creatinine
C0941312|T201|COMP|25104-1|LNC|Glutarate/Creatinine|Glutarate/Creatinine
C0941313|T201|COMP|25105-8|LNC|Glycerate/Creatinine|Glycerate/Creatinine
C0941314|T201|COMP|25106-6|LNC|Glycolate/Creatinine|Glycolate/Creatinine
C0941315|T201|COMP|25107-4|LNC|Glyoxylate/Creatinine|Glyoxylate/Creatinine
C0941316|T201|COMP|25108-2|LNC|Hydroxydecanedioate/Creatinine|Hydroxydecanedioate/Creatinine
C0941317|T201|COMP|25109-0|LNC|Hydroxylysine/Creatinine|Hydroxylysine/Creatinine
C0941318|T201|COMP|25110-8|LNC|Hydroxyproline/Creatinine|Hydroxyproline/Creatinine
C0941319|T201|COMP|25111-6|LNC|Isocitrate/Creatinine|Isocitrate/Creatinine
C0941320|T201|COMP|25113-2|LNC|Malate/Creatinine|Malate/Creatinine
C0941321|T201|COMP|25114-0|LNC|2-Methylcitrate/Creatinine|2-Methylcitrate/Creatinine
C0941322|T201|COMP|25115-7|LNC|Methylmalonate/Creatinine|Methylmalonate/Creatinine
C0941323|T201|COMP|25116-5|LNC|Methylmalonate/Creatinine|Methylmalonate/Creatinine
C0941324|T201|COMP|25118-1|LNC|Mevalonate/Creatinine|Mevalonate/Creatinine
C0941325|T201|COMP|25122-3|LNC|Phosphoethanolamine/Creatinine|Phosphoethanolamine/Creatinine
C0941326|T201|COMP|25123-1|LNC|Para nitrophenol/Creatinine|Para nitrophenol/Creatinine
C0941327|T201|COMP|25124-9|LNC|Phenylacetate/Creatinine|Phenylacetate/Creatinine
C0941328|T201|COMP|25125-6|LNC|Phenyllactate/Creatinine|Phenyllactate/Creatinine
C0941329|T201|COMP|25127-2|LNC|Phosphate/Creatinine|Phosphate/Creatinine
C0941330|T201|COMP|25128-0|LNC|Phosphoserine/Creatinine|Phosphoserine/Creatinine
C0941331|T201|COMP|25129-8|LNC|Pyridinoline/Creatinine|Pyridinoline/Creatinine
C0941332|T201|COMP|25131-4|LNC|Pyridinoline/Creatinine|Pyridinoline/Creatinine
C0941333|T201|COMP|25132-2|LNC|Pyruvate/Creatinine|Pyruvate/Creatinine
C0941334|T201|COMP|25133-0|LNC|Sarcosine/Creatinine|Sarcosine/Creatinine
C0941335|T201|COMP|25135-5|LNC|Suberate/Creatinine|Suberate/Creatinine
C0941336|T201|COMP|25136-3|LNC|Succinate/Creatinine|Succinate/Creatinine
C0941337|T201|COMP|25137-1|LNC|Succinylacetone/Creatinine|Succinylacetone/Creatinine
C0941338|T201|COMP|25138-9|LNC|Taurine/Creatinine|Taurine/Creatinine
C0941339|T201|COMP|25140-5|LNC|Uracil/Creatinine|Uracil/Creatinine
C0941340|T201|COMP|25141-3|LNC|Carnitine esters/Creatinine|Carnitine esters/Creatinine
C0941341|T201|COMP|25142-1|LNC|5-Fluorocytosine^peak|5-Fluorocytosine^peak
C0941342|T201|COMP|25143-9|LNC|5-Fluorocytosine^trough|5-Fluorocytosine^trough
C0941343|T201|COMP|25144-7|LNC|Ammonium urate crystals|Ammonium urate crystals
C0941344|T201|COMP|25145-4|LNC|Bacteria|Bacteria
C0941345|T201|COMP|25146-2|LNC|Bilirubin crystals|Bilirubin crystals
C0941346|T201|COMP|25148-8|LNC|Calcium oxalate crystals|Calcium oxalate crystals
C0941347|T201|COMP|25149-6|LNC|Calcium phosphate crystals|Calcium phosphate crystals
C0941348|T201|COMP|25150-4|LNC|Calcium sulfate crystals|Calcium sulfate crystals
C0941349|T201|COMP|25153-8|LNC|Cholesterol crystals|Cholesterol crystals
C0941350|T201|COMP|25154-6|LNC|Crystals.unidentified|Crystals.unidentified
C0941351|T201|COMP|25155-3|LNC|Cystine crystals|Cystine crystals
C0941352|T201|COMP|25157-9|LNC|Epithelial casts|Epithelial casts
C0941353|T201|COMP|25158-7|LNC|Oval fat bodies (globules)|Oval fat bodies (globules)
C0941354|T201|COMP|25159-5|LNC|Fatty casts|Fatty casts
C0941355|T201|COMP|25160-3|LNC|Granular casts|Granular casts
C0941356|T201|COMP|25161-1|LNC|Hippurate crystals|Hippurate crystals
C0941357|T201|COMP|25162-9|LNC|Hyaline casts|Hyaline casts
C0941358|T201|COMP|25163-7|LNC|Leucine crystals|Leucine crystals
C0941359|T201|COMP|25164-5|LNC|Cells.CD21|Cells.CD21
C0941360|T201|COMP|25165-2|LNC|Cells.CD23|Cells.CD23
C0941361|T201|COMP|25166-0|LNC|Uroporphyrin|Uroporphyrin
C0941362|T201|COMP|25167-8|LNC|Coproporphyrin|Coproporphyrin
C0941363|T201|COMP|25168-6|LNC|Perhexiline|Perhexiline
C0941364|T201|COMP|25169-4|LNC|Nickel|Nickel
C0941365|T201|COMP|25170-2|LNC|Mercury|Mercury
C0941366|T201|COMP|25171-0|LNC|Bromide|Bromide
C0941367|T201|COMP|25172-8|LNC|Fluoride|Fluoride
C0941368|T201|COMP|25173-6|LNC|Thallium|Thallium
C0941369|T201|COMP|25174-4|LNC|Amikacin 8.0 ug/mL|Amikacin 8.0 ug/mL
C0941370|T201|COMP|25175-1|LNC|Amikacin 16.0 ug/mL|Amikacin 16.0 ug/mL
C0941371|T201|COMP|25176-9|LNC|Amikacin 32.0 ug/mL|Amikacin 32.0 ug/mL
C0941372|T201|COMP|25177-7|LNC|Amikacin 12.0 ug/mL|Amikacin 12.0 ug/mL
C0941373|T201|COMP|25179-3|LNC|Amikacin 6.0 ug/mL|Amikacin 6.0 ug/mL
C0941374|T201|COMP|25180-1|LNC|Ciprofloxacin 2.0 ug/mL|Ciprofloxacin 2.0 ug/mL
C0941375|T201|COMP|25181-9|LNC|Ciprofloxacin 4.0 ug/mL|Ciprofloxacin 4.0 ug/mL
C0941376|T201|COMP|25183-5|LNC|Ethionamide 11.0 ug/mL|Ethionamide 11.0 ug/mL
C0941377|T201|COMP|25185-0|LNC|Streptomycin 6.0 ug/mL|Streptomycin 6.0 ug/mL
C0941378|T201|COMP|25186-8|LNC|Pyrazinamide 25.0 ug/mL|Pyrazinamide 25.0 ug/mL
C0941379|T201|COMP|25188-4|LNC|Ciprofloxacin 8.0 ug/mL|Ciprofloxacin 8.0 ug/mL
C0941380|T201|COMP|25189-2|LNC|Ciprofloxacin 5.0 ug/mL|Ciprofloxacin 5.0 ug/mL
C0941381|T201|COMP|25190-0|LNC|Clarithromycin 8.0 ug/mL|Clarithromycin 8.0 ug/mL
C0941382|T201|COMP|25192-6|LNC|Clarithromycin 32.0 ug/mL|Clarithromycin 32.0 ug/mL
C0941383|T201|COMP|25194-2|LNC|Ethambutol 5.0 ug/mL|Ethambutol 5.0 ug/mL
C0941384|T201|COMP|25195-9|LNC|Ethambutol 10.0 ug/mL|Ethambutol 10.0 ug/mL
C0941385|T201|COMP|25196-7|LNC|Ethionamide 5.0 ug/mL|Ethionamide 5.0 ug/mL
C0941386|T201|COMP|25198-3|LNC|Ethionamide 15.0 ug/mL|Ethionamide 15.0 ug/mL
C0941387|T201|COMP|25200-7|LNC|Rifabutin 2.0 ug/mL|Rifabutin 2.0 ug/mL
C0941388|T201|COMP|25201-5|LNC|Rifabutin 4.0 ug/mL|Rifabutin 4.0 ug/mL
C0941389|T201|COMP|25203-1|LNC|rifAMPin 2.0 ug/mL|rifAMPin 2.0 ug/mL
C0941390|T201|COMP|25204-9|LNC|rifAMPin 5.0 ug/mL|rifAMPin 5.0 ug/mL
C0941391|T201|COMP|25205-6|LNC|Streptomycin 2.0 ug/mL|Streptomycin 2.0 ug/mL
C0941392|T201|COMP|25206-4|LNC|Streptomycin 10.0 ug/mL|Streptomycin 10.0 ug/mL
C0941393|T201|COMP|25207-2|LNC|cycloSERINE 10.0 ug/mL|cycloSERINE 10.0 ug/mL
C0941394|T201|COMP|25208-0|LNC|cycloSERINE 20.0 ug/mL|cycloSERINE 20.0 ug/mL
C0941395|T201|COMP|25209-8|LNC|cycloSERINE 30.0 ug/mL|cycloSERINE 30.0 ug/mL
C0941396|T201|COMP|25210-6|LNC|Capreomycin 10.0 ug/mL|Capreomycin 10.0 ug/mL
C0941397|T201|COMP|25211-4|LNC|Capreomycin 20.0 ug/mL|Capreomycin 20.0 ug/mL
C0941398|T201|COMP|25212-2|LNC|Capreomycin 30.0 ug/mL|Capreomycin 30.0 ug/mL
C0941399|T201|COMP|25213-0|LNC|Kanamycin 6.0 ug/mL|Kanamycin 6.0 ug/mL
C0941400|T201|COMP|25214-8|LNC|Kanamycin 30.0 ug/mL|Kanamycin 30.0 ug/mL
C0941401|T201|COMP|25215-5|LNC|Para aminosalicylate 2.0 ug/mL|Para aminosalicylate 2.0 ug/mL
C0941402|T201|COMP|25216-3|LNC|Para aminosalicylate 8.0 ug/mL|Para aminosalicylate 8.0 ug/mL
C0941403|T201|COMP|25217-1|LNC|Isoniazid 0.1 ug/mL|Isoniazid 0.1 ug/mL
C0941404|T201|COMP|25218-9|LNC|Isoniazid 0.2 ug/mL|Isoniazid 0.2 ug/mL
C0941405|T201|COMP|25219-7|LNC|Isoniazid 1.0 ug/mL|Isoniazid 1.0 ug/mL
C0941406|T201|COMP|25220-5|LNC|cefOXitin 30.0 ug/mL|cefOXitin 30.0 ug/mL
C0941407|T201|COMP|25221-3|LNC|Imipenem 10.0 ug/mL|Imipenem 10.0 ug/mL
C0941408|T201|COMP|25222-1|LNC|Cefmetazole 30.0 ug/mL|Cefmetazole 30.0 ug/mL
C0941409|T201|COMP|25224-7|LNC|Erythromycin 15.0 ug/mL|Erythromycin 15.0 ug/mL
C0941410|T201|COMP|25225-4|LNC|Minocycline 30.0 ug/mL|Minocycline 30.0 ug/mL
C0941411|T201|COMP|25226-2|LNC|sulfiSOXAZOLE 300.0 ug/mL|sulfiSOXAZOLE 300.0 ug/mL
C0941412|T201|COMP|25227-0|LNC|Tobramycin 10.0 ug/mL|Tobramycin 10.0 ug/mL
C0941413|T201|COMP|25228-8|LNC|Vancomycin 30.0 ug/mL|Vancomycin 30.0 ug/mL
C0941414|T201|COMP|25229-6|LNC|Pyrazinamide 100.0 ug/mL|Pyrazinamide 100.0 ug/mL
C0941415|T201|COMP|25230-4|LNC|Ethambutol 2.5 ug/mL|Ethambutol 2.5 ug/mL
C0941416|T201|COMP|25231-2|LNC|Ethionamide 10.0 ug/mL|Ethionamide 10.0 ug/mL
C0941417|T201|COMP|25233-8|LNC|Azithromycin|Azithromycin
C0941418|T201|COMP|25234-6|LNC|Aztreonam|Aztreonam
C0941419|T201|COMP|25235-3|LNC|ceFAZolin|ceFAZolin
C0941420|T201|COMP|25236-1|LNC|Cefixime|Cefixime
C0941421|T201|COMP|25238-7|LNC|Cefotaxime|Cefotaxime
C0941422|T201|COMP|25239-5|LNC|cefoTEtan|cefoTEtan
C0941423|T201|COMP|25241-1|LNC|Cefpodoxime|Cefpodoxime
C0941424|T201|COMP|25242-9|LNC|Cefsulodin|Cefsulodin
C0941425|T201|COMP|25243-7|LNC|Ceftizoxime|Ceftizoxime
C0941426|T201|COMP|25245-2|LNC|Cefuroxime.parenteral|Cefuroxime.parenteral
C0941427|T201|COMP|25246-0|LNC|Cephalothin|Cephalothin
C0941428|T201|COMP|25247-8|LNC|Chloramphenicol|Chloramphenicol
C0941429|T201|COMP|25248-6|LNC|Ciprofloxacin|Ciprofloxacin
C0941430|T201|COMP|25250-2|LNC|Cloxacillin|Cloxacillin
C0941431|T201|COMP|25251-0|LNC|cycloSERINE|cycloSERINE
C0941432|T201|COMP|25253-6|LNC|Clarithromycin|Clarithromycin
C0941433|T201|COMP|25254-4|LNC|Ticarcillin|Ticarcillin
C0941434|T201|COMP|25255-1|LNC|Fluconazole|Fluconazole
C0941435|T201|COMP|25256-9|LNC|Ganciclovir|Ganciclovir
C0941436|T201|COMP|25258-5|LNC|Itraconazole|Itraconazole
C0941437|T201|COMP|25259-3|LNC|Ketoconazole|Ketoconazole
C0941438|T201|COMP|25262-7|LNC|Neomycin|Neomycin
C0941439|T201|COMP|25263-5|LNC|Netilmicin|Netilmicin
C0941440|T201|COMP|25266-8|LNC|Oxytetracycline|Oxytetracycline
C0941441|T201|COMP|25267-6|LNC|Penicillin|Penicillin
C0941442|T201|COMP|25268-4|LNC|Piperacillin|Piperacillin
C0941443|T201|COMP|25269-2|LNC|Polymyxin B|Polymyxin B
C0941444|T201|COMP|25270-0|LNC|Pyrazinamide|Pyrazinamide
C0941445|T201|COMP|25271-8|LNC|Sulfamethoxazole|Sulfamethoxazole
C0941446|T201|COMP|25272-6|LNC|Tetracycline|Tetracycline
C0941447|T201|COMP|25274-2|LNC|Amoxicillin|Amoxicillin
C0941448|T201|COMP|25275-9|LNC|Erythromycin|Erythromycin
C0941459|T201|COMP|25287-4|LNC|Streptococcus pneumoniae 19 Ab.IgG^1st specimen|Streptococcus pneumoniae 19 Ab.IgG^1st specimen
C0941460|T201|COMP|25288-2|LNC|Streptococcus pneumoniae 19 Ab.IgG^2nd specimen|Streptococcus pneumoniae 19 Ab.IgG^2nd specimen
C0941462|T201|COMP|25290-8|LNC|Streptococcus pneumoniae 14 Ab.IgG^1st specimen|Streptococcus pneumoniae 14 Ab.IgG^1st specimen
C0941463|T201|COMP|25291-6|LNC|Streptococcus pneumoniae 14 Ab.IgG^2nd specimen|Streptococcus pneumoniae 14 Ab.IgG^2nd specimen
C0941464|T201|COMP|25292-4|LNC|Streptococcus pneumoniae 12 Ab.IgG^1st specimen|Streptococcus pneumoniae 12 Ab.IgG^1st specimen
C0941465|T201|COMP|25293-2|LNC|Streptococcus pneumoniae 12 Ab.IgG^2nd specimen|Streptococcus pneumoniae 12 Ab.IgG^2nd specimen
C0941466|T201|COMP|25294-0|LNC|Streptococcus pneumoniae 1 Ab.IgG^2nd specimen|Streptococcus pneumoniae 1 Ab.IgG^2nd specimen
C0941469|T201|COMP|25297-3|LNC|Parainfluenza virus 1 Ab^2nd specimen|Parainfluenza virus 1 Ab^2nd specimen
C0941470|T201|COMP|25298-1|LNC|Rubella virus Ab.IgG^1st specimen/2nd specimen|Rubella virus Ab.IgG^1st specimen/2nd specimen
C0941471|T201|COMP|25299-9|LNC|Measles virus Ab.IgG^1st specimen/2nd specimen|Measles virus Ab.IgG^1st specimen/2nd specimen
C0941473|T201|COMP|25301-3|LNC|Alanine|Alanine
C0941474|T201|COMP|25302-1|LNC|Alanine aminotransferase|Alanine aminotransferase
C0941475|T201|COMP|25303-9|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C0941476|T201|COMP|25304-7|LNC|Alpha aminoadipate|Alpha aminoadipate
C0941477|T201|COMP|25305-4|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0941478|T201|COMP|25309-6|LNC|Amobarbital|Amobarbital
C0941479|T201|COMP|25310-4|LNC|Amoxicillin+Clavulanate|Amoxicillin+Clavulanate
C0941480|T201|COMP|25312-0|LNC|Amylase.pancreatic/Amylase.total|Amylase.pancreatic/Amylase.total
C0941481|T201|COMP|25313-8|LNC|Amylase.salivary/Amylase.total|Amylase.salivary/Amylase.total
C0941482|T201|COMP|25314-6|LNC|Androstenediol|Androstenediol
C0941483|T201|COMP|25316-1|LNC|17-Hydroxypregnenolone|17-Hydroxypregnenolone
C0941484|T201|COMP|25317-9|LNC|17-Ketosteroids|17-Ketosteroids
C0941485|T201|COMP|25318-7|LNC|1-Methylhistidine|1-Methylhistidine
C0941486|T201|COMP|25319-5|LNC|3-Methylhistidine|3-Methylhistidine
C0941487|T201|COMP|25320-3|LNC|Anserine|Anserine
C0941488|T201|COMP|25321-1|LNC|Antimony|Antimony
C0941489|T201|COMP|25322-9|LNC|Arginine|Arginine
C0941490|T201|COMP|25323-7|LNC|Arsenic|Arsenic
C0941491|T201|COMP|25326-0|LNC|Asparagine|Asparagine
C0941492|T201|COMP|25327-8|LNC|Aspartate|Aspartate
C0941493|T201|COMP|25328-6|LNC|Aspergillus versicolor Ab.IgE.RAST class|Aspergillus versicolor Ab.IgE.RAST class
C0941494|T201|COMP|25331-0|LNC|Bordetella pertussis Ab.IgG|Bordetella pertussis Ab.IgG
C0941495|T201|COMP|25332-8|LNC|Bordetella pertussis Ab.IgM|Bordetella pertussis Ab.IgM
C0941496|T201|COMP|25333-6|LNC|Campylobacter fetus Ab|Campylobacter fetus Ab
C0941497|T201|COMP|25335-1|LNC|Coxiella burnetii Ab.IgG|Coxiella burnetii Ab.IgG
C0941498|T201|COMP|25336-9|LNC|Coxiella burnetii Ab.IgM|Coxiella burnetii Ab.IgM
C0941499|T201|COMP|25337-7|LNC|Taenia solium larva Ab.IgG|Taenia solium larva Ab.IgG
C0941500|T201|COMP|25338-5|LNC|Dengue virus Ab.IgM|Dengue virus Ab.IgM
C0941501|T201|COMP|25339-3|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0941502|T201|COMP|25342-7|LNC|Fasciola sp Ab|Fasciola sp Ab
C0941503|T201|COMP|25343-5|LNC|Fasciola sp Ab.IgG|Fasciola sp Ab.IgG
C0941504|T201|COMP|25344-3|LNC|Filaria Ab|Filaria Ab
C0941505|T201|COMP|25345-0|LNC|Beet red Ab.IgE.RAST class|Beet red Ab.IgE.RAST class
C0941506|T201|COMP|25346-8|LNC|Beta alanine|Beta alanine
C0941507|T201|COMP|25348-4|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0941508|T201|COMP|25349-2|LNC|Betula verrucosa Ab.IgG|Betula verrucosa Ab.IgG
C0941509|T201|COMP|25350-0|LNC|Betula verrucosa Ab.IgG.RAST class|Betula verrucosa Ab.IgG.RAST class
C0941510|T201|COMP|25351-8|LNC|Bismuth|Bismuth
C0941511|T201|COMP|25352-6|LNC|Bordetella pertussis Ab.IgG|Bordetella pertussis Ab.IgG
C0941512|T201|COMP|25353-4|LNC|Bordetella pertussis Ab.IgM|Bordetella pertussis Ab.IgM
C0941513|T201|COMP|25354-2|LNC|Bran wheat Ab.IgG|Bran wheat Ab.IgG
C0941514|T201|COMP|25355-9|LNC|Bran wheat Ab.IgG.RAST class|Bran wheat Ab.IgG.RAST class
C0941515|T201|COMP|25356-7|LNC|Budgerigar droppings Ab.IgE.RAST class|Budgerigar droppings Ab.IgE.RAST class
C0941516|T201|COMP|25357-5|LNC|Butabarbital|Butabarbital
C0941517|T201|COMP|25358-3|LNC|C peptide|C peptide
C0941518|T201|COMP|25359-1|LNC|Cadmium|Cadmium
C0941519|T201|COMP|25360-9|LNC|Cadmium|Cadmium
C0941520|T201|COMP|25363-3|LNC|Campylobacter fetus Ab|Campylobacter fetus Ab
C0941521|T201|COMP|25364-1|LNC|Campylobacter jejuni Ab|Campylobacter jejuni Ab
C0941522|T201|COMP|25367-4|LNC|cefTRIAXone|cefTRIAXone
C0941523|T201|COMP|25368-2|LNC|Cheese blue Ab.IgE.RAST class|Cheese blue Ab.IgE.RAST class
C0941524|T201|COMP|25369-0|LNC|Chlamydia sp Ab.IgA|Chlamydia sp Ab.IgA
C0941525|T201|COMP|25371-6|LNC|Cholesterol.in VLDL|Cholesterol.in VLDL
C0941526|T201|COMP|25372-4|LNC|Choriogonadotropin|Choriogonadotropin
C0941527|T201|COMP|25373-2|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C0941528|T201|COMP|25374-0|LNC|Chromium|Chromium
C0941529|T201|COMP|25376-5|LNC|Citrulline|Citrulline
C0941530|T201|COMP|25377-3|LNC|Coagulation calcium ion induced|Coagulation calcium ion induced
C0941531|T201|COMP|25378-1|LNC|Cobalt|Cobalt
C0941532|T201|COMP|25381-5|LNC|Corticosterone|Corticosterone
C0941533|T201|COMP|25383-1|LNC|Cow milk Ab.IgE.RAST class|Cow milk Ab.IgE.RAST class
C0941534|T201|COMP|25384-9|LNC|Coxiella burnetii Ab.IgG|Coxiella burnetii Ab.IgG
C0941535|T201|COMP|25385-6|LNC|Coxiella burnetii Ab.IgM|Coxiella burnetii Ab.IgM
C0941536|T201|COMP|25386-4|LNC|Creatinine|Creatinine
C0941537|T201|COMP|25388-0|LNC|Cystathionine|Cystathionine
C0941538|T201|COMP|25389-8|LNC|Taenia solium larva Ab.IgG|Taenia solium larva Ab.IgG
C0941539|T201|COMP|25391-4|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C0941540|T201|COMP|25392-2|LNC|Dengue virus Ab.IgM|Dengue virus Ab.IgM
C0941541|T201|COMP|25393-0|LNC|Desethylamiodarone|Desethylamiodarone
C0941542|T201|COMP|25394-8|LNC|Nortrimipramine|Nortrimipramine
C0941543|T201|COMP|25395-5|LNC|Dog serum albumin Ab.IgE.RAST class|Dog serum albumin Ab.IgE.RAST class
C0941544|T201|COMP|25396-3|LNC|Duck meat Ab.IgE.RAST class|Duck meat Ab.IgE.RAST class
C0941545|T201|COMP|25397-1|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0941546|T201|COMP|25399-7|LNC|Endomysium Ab|Endomysium Ab
C0941547|T201|COMP|25400-3|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C0941548|T201|COMP|25401-1|LNC|Estradiol|Estradiol
C0941549|T201|COMP|25402-9|LNC|Estrogen|Estrogen
C0941550|T201|COMP|25403-7|LNC|Estrone|Estrone
C0941551|T201|COMP|25404-5|LNC|Ethambutol|Ethambutol
C0941552|T201|COMP|25405-2|LNC|Ethanolamine|Ethanolamine
C0941553|T201|COMP|25406-0|LNC|Fasciola sp Ab|Fasciola sp Ab
C0941554|T201|COMP|25407-8|LNC|Fasciola sp Ab.IgG|Fasciola sp Ab.IgG
C0941555|T201|COMP|25408-6|LNC|Trigonella foenum-graecum Ab.IgE.RAST class|Trigonella foenum-graecum Ab.IgE.RAST class
C0941556|T201|COMP|25409-4|LNC|Filaria Ab|Filaria Ab
C0941557|T201|COMP|25410-2|LNC|Filaria Ab.IgG|Filaria Ab.IgG
C0941558|T201|COMP|25411-0|LNC|Fleroxacin|Fleroxacin
C0941559|T201|COMP|25412-8|LNC|Flunitrazepam|Flunitrazepam
C0941560|T201|COMP|25413-6|LNC|Fluoride|Fluoride
C0941561|T201|COMP|25414-4|LNC|Gasterophilus intestinalis Ab.IgE.RAST class|Gasterophilus intestinalis Ab.IgE.RAST class
C0941562|T201|COMP|25415-1|LNC|Folate|Folate
C0941563|T201|COMP|25416-9|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C0941564|T201|COMP|25417-7|LNC|Herpes virus 6 Ab.IgM|Herpes virus 6 Ab.IgM
C0941565|T201|COMP|25418-5|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0941566|T201|COMP|25419-3|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C0941567|T201|COMP|25420-1|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C0941568|T201|COMP|25421-9|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C0941569|T201|COMP|25423-5|LNC|Trichinella spiralis Ab.IgG|Trichinella spiralis Ab.IgG
C0941570|T201|COMP|25425-0|LNC|Gabapentin|Gabapentin
C0941571|T201|COMP|25426-8|LNC|Galactose|Galactose
C0941572|T201|COMP|25428-4|LNC|Glucose|Glucose
C0941573|T201|COMP|25429-2|LNC|Glutamate|Glutamate
C0941574|T201|COMP|25430-0|LNC|Glutamine|Glutamine
C0941575|T201|COMP|25432-6|LNC|Haemophilus influenzae Ab|Haemophilus influenzae Ab
C0941576|T201|COMP|25433-4|LNC|Hemoglobin.free|Hemoglobin.free
C0941577|T201|COMP|25434-2|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C0941578|T201|COMP|25438-3|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C0941579|T201|COMP|25439-1|LNC|Histamine|Histamine
C0941580|T201|COMP|25440-9|LNC|Histidine|Histidine
C0941581|T201|COMP|25442-5|LNC|Horse meat Ab.IgE.RAST class|Horse meat Ab.IgE.RAST class
C0941582|T201|COMP|25443-3|LNC|Hydroxylysine|Hydroxylysine
C0941583|T201|COMP|25444-1|LNC|IgA|IgA
C0941584|T201|COMP|25445-8|LNC|IgG|IgG
C0941585|T201|COMP|25447-4|LNC|Insulin.free|Insulin.free
C0941586|T201|COMP|25448-2|LNC|Iodine|Iodine
C0941587|T201|COMP|25449-0|LNC|Iodine|Iodine
C0941588|T201|COMP|25450-8|LNC|Isoleucine|Isoleucine
C0941589|T201|COMP|25451-6|LNC|Isoniazid|Isoniazid
C0941590|T201|COMP|25452-4|LNC|Itraconazole|Itraconazole
C0941591|T201|COMP|25453-2|LNC|Lactalbumin alpha Ab.IgA|Lactalbumin alpha Ab.IgA
C0941592|T201|COMP|25454-0|LNC|Lactalbumin alpha Ab.IgA.RAST class|Lactalbumin alpha Ab.IgA.RAST class
C0941593|T201|COMP|25455-7|LNC|Lactoglobulin Ab.IgA|Lactoglobulin Ab.IgA
C0941594|T201|COMP|25457-3|LNC|Lactoglobulin Ab.IgE.RAST class|Lactoglobulin Ab.IgE.RAST class
C0941595|T201|COMP|25458-1|LNC|lamoTRIgine|lamoTRIgine
C0941596|T201|COMP|25459-9|LNC|Lead|Lead
C0941597|T201|COMP|25460-7|LNC|Leucine|Leucine
C0941598|T201|COMP|25461-5|LNC|Lithium|Lithium
C0941599|T201|COMP|25462-3|LNC|Lithium|Lithium
C0941600|T201|COMP|25463-1|LNC|Lithium|Lithium
C0941601|T201|COMP|25464-9|LNC|Lysine|Lysine
C0941602|T201|COMP|25465-6|LNC|Maleic anhydride Ab.IgE.RAST class|Maleic anhydride Ab.IgE.RAST class
C0941603|T201|COMP|25467-2|LNC|Manganese|Manganese
C0941604|T201|COMP|25468-0|LNC|Mephenytoin|Mephenytoin
C0941605|T201|COMP|25469-8|LNC|Meprobamate|Meprobamate
C0941606|T201|COMP|25470-6|LNC|Mercury|Mercury
C0941607|T201|COMP|25471-4|LNC|Mercury|Mercury
C0941608|T201|COMP|25472-2|LNC|Mesoridazine|Mesoridazine
C0941609|T201|COMP|25473-0|LNC|Metanephrine|Metanephrine
C0941610|T201|COMP|25474-8|LNC|Metanephrines|Metanephrines
C0941611|T201|COMP|25475-5|LNC|Methaqualone|Methaqualone
C0941612|T201|COMP|25476-3|LNC|Methionine|Methionine
C0941613|T201|COMP|25477-1|LNC|Methionine sulfoxide|Methionine sulfoxide
C0941614|T201|COMP|25478-9|LNC|Methyprylon|Methyprylon
C0941615|T201|COMP|25479-7|LNC|Saccharopolyspora rectivirgula Ab.IgG|Saccharopolyspora rectivirgula Ab.IgG
C0941616|T201|COMP|25480-5|LNC|Saccharopolyspora rectivirgula Ab.IgG.RAST class|Saccharopolyspora rectivirgula Ab.IgG.RAST class
C0941617|T201|COMP|25481-3|LNC|Molybdenum|Molybdenum
C0941618|T201|COMP|25485-4|LNC|Neurospora sitophila Ab.IgE.RAST class|Neurospora sitophila Ab.IgE.RAST class
C0941619|T201|COMP|25486-2|LNC|Nickel|Nickel
C0941620|T201|COMP|25487-0|LNC|Nickel|Nickel
C0941621|T201|COMP|25488-8|LNC|Nicotinamide|Nicotinamide
C0941622|T201|COMP|25489-6|LNC|Normetanephrine|Normetanephrine
C0941623|T201|COMP|25490-4|LNC|Olive green Ab.IgE.RAST class|Olive green Ab.IgE.RAST class
C0941624|T201|COMP|25491-2|LNC|Ornithine|Ornithine
C0941625|T201|COMP|25493-8|LNC|Penicillium brevicompactum Ab.IgE.RAST class|Penicillium brevicompactum Ab.IgE.RAST class
C0941626|T201|COMP|25495-3|LNC|Phenylalanine|Phenylalanine
C0941627|T201|COMP|25496-1|LNC|Triplochiton scleroxylon Ab.IgE.RAST class|Triplochiton scleroxylon Ab.IgE.RAST class
C0941628|T201|COMP|25498-7|LNC|Adenosine monophosphate.cyclic|Adenosine monophosphate.cyclic
C0941629|T201|COMP|25500-0|LNC|Phenylbutazone|Phenylbutazone
C0941630|T201|COMP|25501-8|LNC|Phosphate|Phosphate
C0941631|T201|COMP|25503-4|LNC|Phosphoserine|Phosphoserine
C0941632|T201|COMP|15942-6|LNC|Pinus radiata Ab.IgE.RAST class|Pinus radiata Ab.IgE.RAST class
C0941633|T201|COMP|25505-9|LNC|Pituitary glycoprotein hormone.alpha subunit|Pituitary glycoprotein hormone.alpha subunit
C0941634|T201|COMP|25506-7|LNC|Potassium|Potassium
C0941635|T201|COMP|25508-3|LNC|Progesterone^2nd specimen post XXX challenge|Progesterone^2nd specimen post XXX challenge
C0941636|T201|COMP|25509-1|LNC|Progesterone^3rd specimen post XXX challenge|Progesterone^3rd specimen post XXX challenge
C0941637|T201|COMP|25511-7|LNC|Propafenone|Propafenone
C0941638|T201|COMP|25512-5|LNC|Protoporphyrin|Protoporphyrin
C0941639|T201|COMP|25513-3|LNC|Renin^1st specimen post XXX challenge|Renin^1st specimen post XXX challenge
C0941640|T201|COMP|25517-4|LNC|Crocus sativus Ab.IgE.RAST class|Crocus sativus Ab.IgE.RAST class
C0941641|T201|COMP|25518-2|LNC|Sarcosine|Sarcosine
C0941642|T201|COMP|25520-8|LNC|Secobarbital|Secobarbital
C0941643|T201|COMP|25522-4|LNC|Seminal fluid Ab.IgE.RAST class|Seminal fluid Ab.IgE.RAST class
C0941644|T201|COMP|25523-2|LNC|Serine|Serine
C0941645|T201|COMP|25524-0|LNC|Serotonin|Serotonin
C0941646|T201|COMP|25526-5|LNC|Silicon|Silicon
C0941647|T201|COMP|25528-1|LNC|Insulin-like growth factor|Insulin-like growth factor
C0941648|T201|COMP|25529-9|LNC|Somatotropin|Somatotropin
C0941649|T201|COMP|25530-7|LNC|Specimen weight|Specimen weight
C0941650|T201|COMP|25531-5|LNC|Streptococcus pneumoniae Ab|Streptococcus pneumoniae Ab
C0941651|T201|COMP|25532-3|LNC|Swine serum albumin Ab.IgE.RAST class|Swine serum albumin Ab.IgE.RAST class
C0941652|T201|COMP|25533-1|LNC|Taurine|Taurine
C0941653|T201|COMP|25534-9|LNC|Teicoplanin^peak|Teicoplanin^peak
C0941654|T201|COMP|25535-6|LNC|Teicoplanin^trough|Teicoplanin^trough
C0941655|T201|COMP|25536-4|LNC|Clostridium tetani toxoid Ab.IgE.RAST class|Clostridium tetani toxoid Ab.IgE.RAST class
C0941656|T201|COMP|25537-2|LNC|Thallium|Thallium
C0941657|T201|COMP|25538-0|LNC|Thermoactinomyces vulgaris Ab.IgG|Thermoactinomyces vulgaris Ab.IgG
C0941658|T201|COMP|25539-8|LNC|Thermoactinomyces vulgaris Ab.IgG.RAST class|Thermoactinomyces vulgaris Ab.IgG.RAST class
C0941659|T201|COMP|25540-6|LNC|Threonine|Threonine
C0941660|T201|COMP|25541-4|LNC|Topiramate|Topiramate
C0941661|T201|COMP|25542-2|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0941662|T201|COMP|25543-0|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C0941663|T201|COMP|25546-3|LNC|Tryptophan|Tryptophan
C0941664|T201|COMP|25548-9|LNC|Urate|Urate
C0941665|T201|COMP|25549-7|LNC|Urea|Urea
C0941666|T201|COMP|25550-5|LNC|Urea|Urea
C0941667|T201|COMP|25551-3|LNC|Urobilinogen|Urobilinogen
C0941668|T201|COMP|25552-1|LNC|Uroporphyrin|Uroporphyrin
C0941669|T201|COMP|25553-9|LNC|Valine|Valine
C0941670|T201|COMP|25554-7|LNC|Tenebrio mollitor Ab.IgE.RAST class|Tenebrio mollitor Ab.IgE.RAST class
C0941671|T201|COMP|25555-4|LNC|Wuchereria bancrofti Ag|Wuchereria bancrofti Ag
C0941672|T201|COMP|25556-2|LNC|Xylose|Xylose
C0941673|T201|COMP|25557-0|LNC|Zinc|Zinc
C0941674|T201|COMP|25558-8|LNC|Zinc|Zinc
C0941675|T201|COMP|25559-6|LNC|Zolpidem|Zolpidem
C0941676|T201|COMP|25560-4|LNC|Allobarbital|Allobarbital
C0941677|T201|COMP|25561-2|LNC|11-Deoxycorticosterone|11-Deoxycorticosterone
C0941678|T201|COMP|25562-0|LNC|Angiotensin II^supine|Angiotensin II^supine
C0941679|T201|COMP|25563-8|LNC|Angiotensin II^upright|Angiotensin II^upright
C0941680|T201|COMP|25565-3|LNC|Bougainvillea Ab.IgE|Bougainvillea Ab.IgE
C0941681|T201|COMP|25566-1|LNC|Bougainvillea Ab.IgE.RAST class|Bougainvillea Ab.IgE.RAST class
C0941682|T201|COMP|25567-9|LNC|Budgerigar serum proteins Ab.IgE.RAST class|Budgerigar serum proteins Ab.IgE.RAST class
C0941683|T201|COMP|25568-7|LNC|C peptide^10th specimen post XXX challenge|C peptide^10th specimen post XXX challenge
C0941684|T201|COMP|25569-5|LNC|C peptide^11th specimen post XXX challenge|C peptide^11th specimen post XXX challenge
C0941685|T201|COMP|25570-3|LNC|C peptide^12th specimen post XXX challenge|C peptide^12th specimen post XXX challenge
C0941686|T201|COMP|25571-1|LNC|C peptide^13th specimen post XXX challenge|C peptide^13th specimen post XXX challenge
C0941687|T201|COMP|25572-9|LNC|C peptide^14th specimen post XXX challenge|C peptide^14th specimen post XXX challenge
C0941688|T201|COMP|25575-2|LNC|C peptide^2nd specimen post XXX challenge|C peptide^2nd specimen post XXX challenge
C0941689|T201|COMP|25576-0|LNC|C peptide^3rd specimen post XXX challenge|C peptide^3rd specimen post XXX challenge
C0941690|T201|COMP|25577-8|LNC|C peptide^4th specimen post XXX challenge|C peptide^4th specimen post XXX challenge
C0941691|T201|COMP|25578-6|LNC|C peptide^5th specimen post XXX challenge|C peptide^5th specimen post XXX challenge
C0941692|T201|COMP|25579-4|LNC|C peptide^6th specimen post XXX challenge|C peptide^6th specimen post XXX challenge
C0941693|T201|COMP|25580-2|LNC|C peptide^7th specimen post XXX challenge|C peptide^7th specimen post XXX challenge
C0941694|T201|COMP|25581-0|LNC|C peptide^8th specimen post XXX challenge|C peptide^8th specimen post XXX challenge
C0941695|T201|COMP|25582-8|LNC|C peptide^9th specimen post XXX challenge|C peptide^9th specimen post XXX challenge
C0941696|T201|COMP|25584-4|LNC|Calcium^5H post 500 mg calcium PO|Calcium^5H post 500 mg calcium PO
C0941697|T201|COMP|25585-1|LNC|Cat serum albumin Ab.IgE.RAST class|Cat serum albumin Ab.IgE.RAST class
C0941698|T201|COMP|25589-3|LNC|Citalopram|Citalopram
C0941699|T201|COMP|25593-5|LNC|Rotavirus Ab.IgG|Rotavirus Ab.IgG
C0941700|T201|COMP|25596-8|LNC|Fosfomycin|Fosfomycin
C0941701|T201|COMP|25597-6|LNC|Josamycine|Josamycine
C0941702|T201|COMP|25598-4|LNC|Cladosporium cladosporioides Ab.IgG|Cladosporium cladosporioides Ab.IgG
C0941703|T201|COMP|25599-2|LNC|Rotavirus Ab.IgG|Rotavirus Ab.IgG
C0941704|T201|COMP|25600-8|LNC|Rotavirus Ab.IgM|Rotavirus Ab.IgM
C0941705|T201|COMP|25601-6|LNC|Rotavirus Ab.IgM|Rotavirus Ab.IgM
C0941706|T201|COMP|25603-2|LNC|Rickettsia prowazekii Ab.IgG|Rickettsia prowazekii Ab.IgG
C0941707|T201|COMP|25604-0|LNC|Rickettsia prowazekii Ab.IgM|Rickettsia prowazekii Ab.IgM
C0941708|T201|COMP|25607-3|LNC|Miconazole|Miconazole
C0941710|T201|COMP|25609-9|LNC|Cochineal extract Ab.IgE|Cochineal extract Ab.IgE
C0941711|T201|COMP|25610-7|LNC|Cochineal extract Ab.IgE.RAST class|Cochineal extract Ab.IgE.RAST class
C0941712|T201|COMP|25611-5|LNC|Blatta orientalis Ab.IgE|Blatta orientalis Ab.IgE
C0941713|T201|COMP|25612-3|LNC|Blatta orientalis Ab.IgE.RAST class|Blatta orientalis Ab.IgE.RAST class
C0941714|T201|COMP|25614-9|LNC|Periplaneta fuliginosa Ab.IgE.RAST class|Periplaneta fuliginosa Ab.IgE.RAST class
C0941715|T201|COMP|25615-6|LNC|Conalbumin Ab.IgE|Conalbumin Ab.IgE
C0941716|T201|COMP|25616-4|LNC|Conalbumin Ab.IgE.RAST class|Conalbumin Ab.IgE.RAST class
C0941717|T201|COMP|25617-2|LNC|Cortisol^1H post 250 ug cortrosyn IM|Cortisol^1H post 250 ug cortrosyn IM
C0941718|T201|COMP|25618-0|LNC|Cortisol^1st specimen post XXX challenge|Cortisol^1st specimen post XXX challenge
C0941719|T201|COMP|25619-8|LNC|Cortisol^2nd specimen post XXX challenge|Cortisol^2nd specimen post XXX challenge
C0941720|T201|COMP|25620-6|LNC|Cortisol^30M post 250 ug cortrosyn IM|Cortisol^30M post 250 ug cortrosyn IM
C0941721|T201|COMP|25621-4|LNC|Cortisol^3rd specimen post XXX challenge|Cortisol^3rd specimen post XXX challenge
C0941722|T201|COMP|25622-2|LNC|Cortisol^4th specimen post XXX challenge|Cortisol^4th specimen post XXX challenge
C0941723|T201|COMP|25623-0|LNC|Cortisol^5th specimen post XXX challenge|Cortisol^5th specimen post XXX challenge
C0941724|T201|COMP|25624-8|LNC|Cortisol^6th specimen post XXX challenge|Cortisol^6th specimen post XXX challenge
C0941725|T201|COMP|25625-5|LNC|Cortisol^7th specimen post XXX challenge|Cortisol^7th specimen post XXX challenge
C0941726|T201|COMP|25627-1|LNC|Cortisol^8th specimen post XXX challenge|Cortisol^8th specimen post XXX challenge
C0941727|T201|COMP|25628-9|LNC|Cortisol^9th specimen post XXX challenge|Cortisol^9th specimen post XXX challenge
C0941728|T201|COMP|25629-7|LNC|Cortisol^pre 250 ug cortrosyn IM|Cortisol^pre 250 ug cortrosyn IM
C0941729|T201|COMP|25630-5|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0941730|T201|COMP|25631-3|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0941731|T201|COMP|25632-1|LNC|Plasmodium sp Ab|Plasmodium sp Ab
C0941732|T201|COMP|25634-7|LNC|Ribes sylvestre Ab.IgE.RAST class|Ribes sylvestre Ab.IgE.RAST class
C0941733|T201|COMP|25637-0|LNC|Econazole|Econazole
C0941734|T201|COMP|25638-8|LNC|Eosinophil cationic protein|Eosinophil cationic protein
C0941735|T201|COMP|25639-6|LNC|Follitropin|Follitropin
C0941738|T201|COMP|25642-0|LNC|Follitropin^1st specimen post XXX challenge|Follitropin^1st specimen post XXX challenge
C0941739|T201|COMP|25644-6|LNC|Follitropin^2nd specimen post XXX challenge|Follitropin^2nd specimen post XXX challenge
C0941741|T201|COMP|25646-1|LNC|Follitropin^3rd specimen post XXX challenge|Follitropin^3rd specimen post XXX challenge
C0941742|T201|COMP|25648-7|LNC|Follitropin^5th specimen post XXX challenge|Follitropin^5th specimen post XXX challenge
C0941743|T201|COMP|25649-5|LNC|Follitropin^6th specimen post XXX challenge|Follitropin^6th specimen post XXX challenge
C0941744|T201|COMP|25650-3|LNC|Follitropin^7th specimen post XXX challenge|Follitropin^7th specimen post XXX challenge
C0941745|T201|COMP|25651-1|LNC|Follitropin^8th specimen post XXX challenge|Follitropin^8th specimen post XXX challenge
C0941746|T201|COMP|25652-9|LNC|Follitropin^9th specimen post XXX challenge|Follitropin^9th specimen post XXX challenge
C0941747|T201|COMP|25653-7|LNC|Fosfomycin|Fosfomycin
C0941748|T201|COMP|25655-2|LNC|Gastrin^2nd specimen post XXX challenge|Gastrin^2nd specimen post XXX challenge
C0941749|T201|COMP|25656-0|LNC|Gastrin^3rd specimen post XXX challenge|Gastrin^3rd specimen post XXX challenge
C0941750|T201|COMP|25657-8|LNC|Gastrin^4th specimen post XXX challenge|Gastrin^4th specimen post XXX challenge
C0941751|T201|COMP|25658-6|LNC|Gastrin^5th specimen post XXX challenge|Gastrin^5th specimen post XXX challenge
C0941752|T201|COMP|25659-4|LNC|Gastrin^6th specimen post XXX challenge|Gastrin^6th specimen post XXX challenge
C0941753|T201|COMP|25660-2|LNC|Gastrin^7th specimen post XXX challenge|Gastrin^7th specimen post XXX challenge
C0941754|T201|COMP|25661-0|LNC|Gastrin^8th specimen post XXX challenge|Gastrin^8th specimen post XXX challenge
C0941755|T201|COMP|25662-8|LNC|Gastrin^9th specimen post XXX challenge|Gastrin^9th specimen post XXX challenge
C0941756|T201|COMP|25663-6|LNC|Glucose^15M post dose glucose|Glucose^15M post dose glucose
C0941757|T201|COMP|25664-4|LNC|Glucose^1H post dose glucose|Glucose^1H post dose glucose
C0941758|T201|COMP|25665-1|LNC|Glucose^1H post XXX challenge|Glucose^1H post XXX challenge
C0941759|T201|COMP|25667-7|LNC|Glucose^2H post dose glucose|Glucose^2H post dose glucose
C0941760|T201|COMP|25668-5|LNC|Glucose^2H post XXX challenge|Glucose^2H post XXX challenge
C0941761|T201|COMP|25669-3|LNC|Glucose^3.5H post dose glucose|Glucose^3.5H post dose glucose
C0941762|T201|COMP|25670-1|LNC|Glucose^30M post dose glucose|Glucose^30M post dose glucose
C0941763|T201|COMP|25671-9|LNC|Glucose^30M post XXX challenge|Glucose^30M post XXX challenge
C0941764|T201|COMP|25672-7|LNC|Glucose^4.5H post dose glucose|Glucose^4.5H post dose glucose
C0941765|T201|COMP|25673-5|LNC|Glucose^45M post dose glucose|Glucose^45M post dose glucose
C0941766|T201|COMP|25674-3|LNC|Glucose^45M post XXX challenge|Glucose^45M post XXX challenge
C0941767|T201|COMP|25675-0|LNC|Glucose^4H post dose glucose|Glucose^4H post dose glucose
C0941768|T201|COMP|25676-8|LNC|Glucose^5.5H post dose glucose|Glucose^5.5H post dose glucose
C0941769|T201|COMP|25677-6|LNC|Glucose^6H post dose glucose|Glucose^6H post dose glucose
C0941770|T201|COMP|25679-2|LNC|Glucose^1.5H post XXX challenge|Glucose^1.5H post XXX challenge
C0941771|T201|COMP|25680-0|LNC|Glucose^pre 50 g glucose PO|Glucose^pre 50 g glucose PO
C0941772|T201|COMP|25681-8|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C0941773|T201|COMP|25682-6|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C0941774|T201|COMP|25683-4|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C0941775|T201|COMP|25684-2|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C0941776|T201|COMP|25685-9|LNC|Insulin^10th specimen post XXX challenge|Insulin^10th specimen post XXX challenge
C0941777|T201|COMP|25686-7|LNC|Insulin^11th specimen post XXX challenge|Insulin^11th specimen post XXX challenge
C0941778|T201|COMP|25687-5|LNC|Insulin^12th specimen post XXX challenge|Insulin^12th specimen post XXX challenge
C0941779|T201|COMP|25688-3|LNC|Insulin^13th specimen post XXX challenge|Insulin^13th specimen post XXX challenge
C0941780|T201|COMP|25689-1|LNC|Insulin^14th specimen post XXX challenge|Insulin^14th specimen post XXX challenge
C0941781|T201|COMP|25691-7|LNC|Insulin^1st specimen post XXX challenge|Insulin^1st specimen post XXX challenge
C0941782|T201|COMP|25692-5|LNC|Insulin^2nd specimen post XXX challenge|Insulin^2nd specimen post XXX challenge
C0941783|T201|COMP|25693-3|LNC|Insulin^3rd specimen post XXX challenge|Insulin^3rd specimen post XXX challenge
C0941784|T201|COMP|25694-1|LNC|Insulin^4th specimen post XXX challenge|Insulin^4th specimen post XXX challenge
C0941785|T201|COMP|25695-8|LNC|Insulin^5th specimen post XXX challenge|Insulin^5th specimen post XXX challenge
C0941786|T201|COMP|25697-4|LNC|Insulin^7th specimen post XXX challenge|Insulin^7th specimen post XXX challenge
C0941787|T201|COMP|25698-2|LNC|Insulin^8th specimen post XXX challenge|Insulin^8th specimen post XXX challenge
C0941788|T201|COMP|25700-6|LNC|Interpretation|Interpretation
C0941789|T201|COMP|25701-4|LNC|Artocarpus heterophyllus Ab.IgE.RAST class|Artocarpus heterophyllus Ab.IgE.RAST class
C0941790|T201|COMP|25702-2|LNC|Josamycine|Josamycine
C0941791|T201|COMP|25703-0|LNC|Ziziphus jujuba Ab.IgE|Ziziphus jujuba Ab.IgE
C0941792|T201|COMP|25705-5|LNC|Ketones^1H post 50 g glucose PO|Ketones^1H post 50 g glucose PO
C0941793|T201|COMP|25706-3|LNC|Ketones^2H post dose glucose|Ketones^2H post dose glucose
C0941794|T201|COMP|25707-1|LNC|Ketones^4H post dose glucose|Ketones^4H post dose glucose
C0941795|T201|COMP|25708-9|LNC|Leishmania donovani Ab|Leishmania donovani Ab
C0941796|T201|COMP|25710-5|LNC|Leptospira interrogans serovar Grippotyphosa Ab|Leptospira interrogans serovar Grippotyphosa Ab
C0941799|T201|COMP|25714-7|LNC|Litchi chinensis Ab.IgE|Litchi chinensis Ab.IgE
C0941800|T201|COMP|25715-4|LNC|Litchi chinensis Ab.IgE.RAST class|Litchi chinensis Ab.IgE.RAST class
C0941801|T201|COMP|25716-2|LNC|Lutropin|Lutropin
C0941806|T201|COMP|25721-2|LNC|Mianserin|Mianserin
C0941807|T201|COMP|25722-0|LNC|Miconazole|Miconazole
C0941808|T201|COMP|25723-8|LNC|Nitroxoline|Nitroxoline
C0941809|T201|COMP|6897-3|LNC|Norsertraline|Norsertraline
C0941810|T201|COMP|25725-3|LNC|Ovary Ab|Ovary Ab
C0941811|T201|COMP|25726-1|LNC|OXcarbazepine|OXcarbazepine
C0941812|T201|COMP|25728-7|LNC|Parkinsonia florida Ab.IgE.RAST class|Parkinsonia florida Ab.IgE.RAST class
C0941813|T201|COMP|25729-5|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0941814|T201|COMP|25730-3|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0941815|T201|COMP|25731-1|LNC|Plasmodium sp Ab|Plasmodium sp Ab
C0941816|T201|COMP|25732-9|LNC|Pregnanetriolone|Pregnanetriolone
C0941817|T201|COMP|25733-7|LNC|Procollagen type III|Procollagen type III
C0941818|T201|COMP|25734-5|LNC|Prolactin^10M post 200 ug TRH IV|Prolactin^10M post 200 ug TRH IV
C0941819|T201|COMP|25736-0|LNC|Prolactin^1st specimen post XXX challenge|Prolactin^1st specimen post XXX challenge
C0941820|T201|COMP|25737-8|LNC|Prolactin^20M post 200 ug TRH IV|Prolactin^20M post 200 ug TRH IV
C0941821|T201|COMP|25738-6|LNC|Prolactin^2H post 200 ug TRH IV|Prolactin^2H post 200 ug TRH IV
C0941822|T201|COMP|25739-4|LNC|Prolactin^30M post 200 ug TRH IV|Prolactin^30M post 200 ug TRH IV
C0941823|T201|COMP|25740-2|LNC|Prolactin^40M post 200 ug TRH IV|Prolactin^40M post 200 ug TRH IV
C0941824|T201|COMP|25741-0|LNC|Prolactin^50M post 200 ug TRH IV|Prolactin^50M post 200 ug TRH IV
C0941825|T201|COMP|25742-8|LNC|Prothrombin fragment 1+2|Prothrombin fragment 1+2
C0941826|T201|COMP|25743-6|LNC|Chenopodium quinoa Ab.IgE|Chenopodium quinoa Ab.IgE
C0941827|T201|COMP|25744-4|LNC|Chenopodium quinoa Ab.IgE.RAST class|Chenopodium quinoa Ab.IgE.RAST class
C0941828|T201|COMP|25745-1|LNC|Rheumatoid factor|Rheumatoid factor
C0941829|T201|COMP|25747-7|LNC|Ribosomal Ab|Ribosomal Ab
C0941830|T201|COMP|25749-3|LNC|Rickettsia conorii Ab.IgG|Rickettsia conorii Ab.IgG
C0941831|T201|COMP|25751-9|LNC|Rickettsia prowazekii Ab.IgG|Rickettsia prowazekii Ab.IgG
C0941832|T201|COMP|25752-7|LNC|Rickettsia prowazekii Ab.IgM|Rickettsia prowazekii Ab.IgM
C0941833|T201|COMP|25753-5|LNC|Rotavirus Ab.IgG|Rotavirus Ab.IgG
C0941834|T201|COMP|25754-3|LNC|Rotavirus Ab.IgG|Rotavirus Ab.IgG
C0941835|T201|COMP|25756-8|LNC|Rotavirus Ab.IgM|Rotavirus Ab.IgM
C0941836|T201|COMP|25757-6|LNC|Schistosoma sp Ab.IgG|Schistosoma sp Ab.IgG
C0941849|T201|COMP|25772-5|LNC|Somatotropin^11th specimen post XXX challenge|Somatotropin^11th specimen post XXX challenge
C0941850|T201|COMP|25773-3|LNC|Somatotropin^12th specimen post XXX challenge|Somatotropin^12th specimen post XXX challenge
C0941851|T201|COMP|25774-1|LNC|Somatotropin^13th specimen post XXX challenge|Somatotropin^13th specimen post XXX challenge
C0941852|T201|COMP|25775-8|LNC|Somatotropin^14th specimen post XXX challenge|Somatotropin^14th specimen post XXX challenge
C0941853|T201|COMP|25776-6|LNC|Somatotropin^1st specimen post XXX challenge|Somatotropin^1st specimen post XXX challenge
C0941854|T201|COMP|25777-4|LNC|Somatotropin^40M post XXX challenge|Somatotropin^40M post XXX challenge
C0941855|T201|COMP|25778-2|LNC|Somatotropin^50M post XXX challenge|Somatotropin^50M post XXX challenge
C0941856|T201|COMP|25779-0|LNC|Stachybotrys chartarum Ab.IgG|Stachybotrys chartarum Ab.IgG
C0941857|T201|COMP|25780-8|LNC|Stachybotrys chartarum Ab.IgG.RAST class|Stachybotrys chartarum Ab.IgG.RAST class
C0941858|T201|COMP|25788-1|LNC|Streptolysin O Ab|Streptolysin O Ab
C0941859|T201|COMP|25789-9|LNC|Thyrotropin^1st specimen post XXX challenge|Thyrotropin^1st specimen post XXX challenge
C0941860|T201|COMP|25790-7|LNC|Thyroxine.free^1st specimen post XXX challenge|Thyroxine.free^1st specimen post XXX challenge
C0941861|T201|COMP|25791-5|LNC|Thyroxine.free^2nd specimen post XXX challenge|Thyroxine.free^2nd specimen post XXX challenge
C0941862|T201|COMP|25792-3|LNC|Thyroxine.free^3rd specimen post XXX challenge|Thyroxine.free^3rd specimen post XXX challenge
C0941863|T201|COMP|25794-9|LNC|Thyroxine.free^5th specimen post XXX challenge|Thyroxine.free^5th specimen post XXX challenge
C0941864|T201|COMP|25795-6|LNC|Thyroxine.free^6th specimen post XXX challenge|Thyroxine.free^6th specimen post XXX challenge
C0941865|T201|COMP|25796-4|LNC|Thyroxine.free^7th specimen post XXX challenge|Thyroxine.free^7th specimen post XXX challenge
C0941866|T201|COMP|25797-2|LNC|Thyroxine.free^8th specimen post XXX challenge|Thyroxine.free^8th specimen post XXX challenge
C0941867|T201|COMP|25798-0|LNC|Thyroxine.free^9th specimen post XXX challenge|Thyroxine.free^9th specimen post XXX challenge
C0941868|T201|COMP|25799-8|LNC|Tissue polypeptide specific Ag|Tissue polypeptide specific Ag
C0941869|T201|COMP|25800-4|LNC|Tobramycin|Tobramycin
C0941880|T201|COMP|25813-7|LNC|Trypanosoma cruzi Ab|Trypanosoma cruzi Ab
C0941881|T201|COMP|25815-2|LNC|Lathyrus sativus Ab.IgE.RAST class|Lathyrus sativus Ab.IgE.RAST class
C0941882|T201|COMP|25818-6|LNC|Xylose^1H post dose xylose PO|Xylose^1H post dose xylose PO
C0941883|T201|COMP|25819-4|LNC|Xylose^baseline|Xylose^baseline
C0941884|T201|COMP|25820-2|LNC|Cysteate|Cysteate
C0941885|T201|COMP|25821-0|LNC|Staphylococcus aureus enterotoxin A Ab.IgE|Staphylococcus aureus enterotoxin A Ab.IgE
C0941887|T201|COMP|25824-4|LNC|Staphylococcus aureus enterotoxin C Ab.IgE|Staphylococcus aureus enterotoxin C Ab.IgE
C0941889|T201|COMP|25826-9|LNC|Staphylococcus aureus enterotoxin D Ab.IgE|Staphylococcus aureus enterotoxin D Ab.IgE
C0941890|T201|COMP|25828-5|LNC|Parkinsonia florida Ab.IgE|Parkinsonia florida Ab.IgE
C0941891|T201|COMP|25829-3|LNC|Glucosylceramidase|Glucosylceramidase
C0941892|T201|COMP|25830-1|LNC|Beta glucosidase activator|Beta glucosidase activator
C0941893|T201|COMP|25831-9|LNC|Beta-N-acetylhexosaminidase.A|Beta-N-acetylhexosaminidase.A
C0941894|T201|COMP|25832-7|LNC|Beta-N-acetylhexosaminidase.A activator|Beta-N-acetylhexosaminidase.A activator
C0941895|T201|COMP|25834-3|LNC|Cancer associated retinopathy Ab|Cancer associated retinopathy Ab
C0941896|T201|COMP|25836-8|LNC|HIV 1 RNA|HIV 1 RNA
C0941897|T201|COMP|25837-6|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C0941898|T201|COMP|25838-4|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C0941899|T201|COMP|25839-2|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C0941900|T201|COMP|25840-0|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C0941901|T201|COMP|25841-8|LNC|HIV 2 proviral DNA|HIV 2 proviral DNA
C0941902|T201|COMP|25842-6|LNC|HIV 2 proviral DNA|HIV 2 proviral DNA
C0941903|T201|COMP|25843-4|LNC|Alanine|Alanine
C0941904|T201|COMP|25844-2|LNC|Alanine/Creatinine|Alanine/Creatinine
C0941905|T201|COMP|25845-9|LNC|Aldosterone|Aldosterone
C0941906|T201|COMP|25846-7|LNC|Alpha aminoadipate|Alpha aminoadipate
C0941907|T201|COMP|25847-5|LNC|Alpha aminoadipate/Creatinine|Alpha aminoadipate/Creatinine
C0941908|T201|COMP|25848-3|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0941909|T201|COMP|25849-1|LNC|Alpha aminobutyrate/Creatinine|Alpha aminobutyrate/Creatinine
C0941910|T201|COMP|25850-9|LNC|Ammonia|Ammonia
C0941911|T201|COMP|25851-7|LNC|Ammonia/Creatinine|Ammonia/Creatinine
C0941912|T201|COMP|25852-5|LNC|17-Hydroxycorticosteroids|17-Hydroxycorticosteroids
C0941913|T201|COMP|25853-3|LNC|1-Methylhistidine|1-Methylhistidine
C0941914|T201|COMP|25854-1|LNC|1-Methylhistidine/Creatinine|1-Methylhistidine/Creatinine
C0941915|T201|COMP|25855-8|LNC|3-Alpha-Androstanediol glucuronide|3-Alpha-Androstanediol glucuronide
C0941916|T201|COMP|25856-6|LNC|3-Methylhistidine|3-Methylhistidine
C0941917|T201|COMP|25857-4|LNC|3-Methylhistidine/Creatinine|3-Methylhistidine/Creatinine
C0941918|T201|COMP|25858-2|LNC|Anserine|Anserine
C0941919|T201|COMP|25859-0|LNC|Anserine/Creatinine|Anserine/Creatinine
C0941920|T201|COMP|25860-8|LNC|Arginine|Arginine
C0941921|T201|COMP|25861-6|LNC|Arginine/Creatinine|Arginine/Creatinine
C0941922|T201|COMP|25862-4|LNC|Asparagine|Asparagine
C0941923|T201|COMP|25864-0|LNC|Aspartate|Aspartate
C0941924|T201|COMP|25867-3|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0941925|T201|COMP|25869-9|LNC|Beta alanine/Creatinine|Beta alanine/Creatinine
C0941926|T201|COMP|25870-7|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0941927|T201|COMP|25871-5|LNC|Beta aminoisobutyrate/Creatinine|Beta aminoisobutyrate/Creatinine
C0941928|T201|COMP|25873-1|LNC|Calcium^pre 500 mg calcium PO|Calcium^pre 500 mg calcium PO
C0941929|T201|COMP|25874-9|LNC|Carnosine|Carnosine
C0941930|T201|COMP|25875-6|LNC|Carnosine/Creatinine|Carnosine/Creatinine
C0941931|T201|COMP|25877-2|LNC|Citrulline|Citrulline
C0941932|T201|COMP|25878-0|LNC|Citrulline/Creatinine|Citrulline/Creatinine
C0941933|T201|COMP|25879-8|LNC|Copper|Copper
C0941934|T201|COMP|25880-6|LNC|Copper/Creatinine|Copper/Creatinine
C0941935|T201|COMP|25881-4|LNC|Coproporphyrin|Coproporphyrin
C0941936|T201|COMP|25882-2|LNC|Cortisol.free|Cortisol.free
C0941937|T201|COMP|25883-0|LNC|Cortisol.free|Cortisol.free
C0941938|T201|COMP|25885-5|LNC|Cortisol.free|Cortisol.free
C0941939|T201|COMP|25886-3|LNC|Creatinine|Creatinine
C0941940|T201|COMP|25887-1|LNC|Cystathionine|Cystathionine
C0941941|T201|COMP|25888-9|LNC|Cystathionine/Creatinine|Cystathionine/Creatinine
C0941942|T201|COMP|25890-5|LNC|Cysteate/Creatinine|Cysteate/Creatinine
C0941943|T201|COMP|25891-3|LNC|Cysteine|Cysteine
C0941944|T201|COMP|25893-9|LNC|Cysteine/Creatinine|Cysteine/Creatinine
C0941945|T201|COMP|25894-7|LNC|Cystine/Creatinine|Cystine/Creatinine
C0941946|T201|COMP|25895-4|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C0941947|T201|COMP|25896-2|LNC|Delta aminolevulinate|Delta aminolevulinate
C0941948|T201|COMP|25897-0|LNC|Delta aminolevulinate/Creatinine|Delta aminolevulinate/Creatinine
C0941949|T201|COMP|25898-8|LNC|Deoxypyridinoline|Deoxypyridinoline
C0941950|T201|COMP|25899-6|LNC|D-Lactate^1st specimen post exercise|D-Lactate^1st specimen post exercise
C0941951|T201|COMP|25901-0|LNC|D-Lactate^3rd specimen post exercise|D-Lactate^3rd specimen post exercise
C0941952|T201|COMP|25902-8|LNC|D-Lactate^4th specimen post exercise|D-Lactate^4th specimen post exercise
C0941953|T201|COMP|25904-4|LNC|D-Lactate^6th specimen post exercise|D-Lactate^6th specimen post exercise
C0941954|T201|COMP|25905-1|LNC|D-lactate^pre exercise|D-lactate^pre exercise
C0941955|T201|COMP|25906-9|LNC|DOPamine|DOPamine
C0941956|T201|COMP|25907-7|LNC|Elastase.pancreatic|Elastase.pancreatic
C0941957|T201|COMP|25908-5|LNC|EPINEPHrine|EPINEPHrine
C0941958|T201|COMP|25909-3|LNC|EPINEPHrine/Creatinine|EPINEPHrine/Creatinine
C0941959|T201|COMP|25910-1|LNC|Ethanolamine|Ethanolamine
C0941960|T201|COMP|25911-9|LNC|Ethanolamine/Creatinine|Ethanolamine/Creatinine
C0941961|T201|COMP|25912-7|LNC|Fluoride|Fluoride
C0941962|T201|COMP|25913-5|LNC|Fluoride/Creatinine|Fluoride/Creatinine
C0941963|T201|COMP|25914-3|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0941964|T201|COMP|25915-0|LNC|Gamma aminobutyrate/Creatinine|Gamma aminobutyrate/Creatinine
C0941965|T201|COMP|25916-8|LNC|Glucose|Glucose
C0941966|T201|COMP|25917-6|LNC|Glutamate|Glutamate
C0941967|T201|COMP|25918-4|LNC|Glutamate/Creatinine|Glutamate/Creatinine
C0941968|T201|COMP|25919-2|LNC|Glutamine|Glutamine
C0941969|T201|COMP|25920-0|LNC|Glutamine/Creatinine|Glutamine/Creatinine
C0941970|T201|COMP|25921-8|LNC|Glycine|Glycine
C0941971|T201|COMP|25922-6|LNC|Glycine/Creatinine|Glycine/Creatinine
C0941972|T201|COMP|25923-4|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C0941973|T201|COMP|25924-2|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C0941974|T201|COMP|25926-7|LNC|Histidine|Histidine
C0941975|T201|COMP|25927-5|LNC|Histidine/Creatinine|Histidine/Creatinine
C0941976|T201|COMP|25928-3|LNC|Homocystine|Homocystine
C0941977|T201|COMP|25929-1|LNC|Homocystine/Creatinine|Homocystine/Creatinine
C0941978|T201|COMP|25930-9|LNC|Homovanillate|Homovanillate
C0941979|T201|COMP|25931-7|LNC|Homovanillate/Creatinine|Homovanillate/Creatinine
C0941980|T201|COMP|25932-5|LNC|Hydroxylysine|Hydroxylysine
C0941981|T201|COMP|25934-1|LNC|Hydroxyproline|Hydroxyproline
C0941982|T201|COMP|25939-0|LNC|Isoleucine/Creatinine|Isoleucine/Creatinine
C0941983|T201|COMP|25940-8|LNC|Leptospira borgpetersenii serovar Sejroe Ab|Leptospira borgpetersenii serovar Sejroe Ab
C0941984|T201|COMP|25941-6|LNC|Leucine|Leucine
C0941985|T201|COMP|25943-2|LNC|Lutropin^1st specimen post XXX challenge|Lutropin^1st specimen post XXX challenge
C0941986|T201|COMP|25944-0|LNC|Lutropin^2nd specimen post XXX challenge|Lutropin^2nd specimen post XXX challenge
C0941987|T201|COMP|25945-7|LNC|Lutropin^3rd specimen post XXX challenge|Lutropin^3rd specimen post XXX challenge
C0941988|T201|COMP|25947-3|LNC|Lutropin^5th specimen post XXX challenge|Lutropin^5th specimen post XXX challenge
C0941989|T201|COMP|25948-1|LNC|Lutropin^6th specimen post XXX challenge|Lutropin^6th specimen post XXX challenge
C0941990|T201|COMP|25949-9|LNC|Lutropin^7th specimen post XXX challenge|Lutropin^7th specimen post XXX challenge
C0941991|T201|COMP|25950-7|LNC|Lutropin^8th specimen post XXX challenge|Lutropin^8th specimen post XXX challenge
C0941992|T201|COMP|25951-5|LNC|Lutropin^9th specimen post XXX challenge|Lutropin^9th specimen post XXX challenge
C0941993|T201|COMP|25953-1|LNC|Lysine/Creatinine|Lysine/Creatinine
C0941994|T201|COMP|25954-9|LNC|Magnesium|Magnesium
C0941995|T201|COMP|25955-6|LNC|Metanephrine|Metanephrine
C0941996|T201|COMP|25957-2|LNC|Methionine sulfoxide|Methionine sulfoxide
C0941997|T201|COMP|25958-0|LNC|Methionine sulfoxide/Creatinine|Methionine sulfoxide/Creatinine
C0941998|T201|COMP|25959-8|LNC|Methionine/Creatinine|Methionine/Creatinine
C0942000|T201|COMP|25961-4|LNC|Nickel|Nickel
C0942001|T201|COMP|25962-2|LNC|Nickel/Creatinine|Nickel/Creatinine
C0942002|T201|COMP|25964-8|LNC|Normetanephrine|Normetanephrine
C0942003|T201|COMP|25965-5|LNC|Ornithine|Ornithine
C0942004|T201|COMP|25966-3|LNC|Ornithine/Creatinine|Ornithine/Creatinine
C0942005|T201|COMP|25967-1|LNC|Penicillium roqueforti Ab.IgE.RAST class|Penicillium roqueforti Ab.IgE.RAST class
C0942006|T201|COMP|25968-9|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C0942007|T201|COMP|25969-7|LNC|Phenylalanine|Phenylalanine
C0942008|T201|COMP|25970-5|LNC|Phenylalanine/Creatinine|Phenylalanine/Creatinine
C0942009|T201|COMP|25971-3|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C0942010|T201|COMP|25972-1|LNC|Adenosine monophosphate.cyclic/Creatinine|Adenosine monophosphate.cyclic/Creatinine
C0942011|T201|COMP|25973-9|LNC|Phosphate|Phosphate
C0942012|T201|COMP|25974-7|LNC|Phosphoserine/Creatinine|Phosphoserine/Creatinine
C0942013|T201|COMP|25975-4|LNC|Proline|Proline
C0942014|T201|COMP|25976-2|LNC|Proline/Creatinine|Proline/Creatinine
C0942015|T201|COMP|25977-0|LNC|Pyridinoline|Pyridinoline
C0942016|T201|COMP|25978-8|LNC|Sarcosine/Creatinine|Sarcosine/Creatinine
C0942017|T201|COMP|25979-6|LNC|Serine|Serine
C0942018|T201|COMP|25980-4|LNC|Serine/Creatinine|Serine/Creatinine
C0942019|T201|COMP|25981-2|LNC|Serotonin|Serotonin
C0942020|T201|COMP|25982-0|LNC|Sheep milk Ab.IgE.RAST class|Sheep milk Ab.IgE.RAST class
C0942021|T201|COMP|25983-8|LNC|Sheep whey Ab.IgE.RAST class|Sheep whey Ab.IgE.RAST class
C0942022|T201|COMP|25984-6|LNC|Somatotropin^30M post XXX challenge|Somatotropin^30M post XXX challenge
C0942023|T201|COMP|25985-3|LNC|Taurine/Creatinine|Taurine/Creatinine
C0942024|T201|COMP|25986-1|LNC|Testosterone|Testosterone
C0942025|T201|COMP|25987-9|LNC|Testosterone.free|Testosterone.free
C0942026|T201|COMP|25988-7|LNC|Threonine|Threonine
C0942027|T201|COMP|25989-5|LNC|Threonine/Creatinine|Threonine/Creatinine
C0942028|T201|COMP|25991-1|LNC|Thyrotropin^pre dose TRH IN|Thyrotropin^pre dose TRH IN
C0942029|T201|COMP|25993-7|LNC|Trichinella spiralis Ab|Trichinella spiralis Ab
C0942030|T201|COMP|25994-5|LNC|Tryptophan/Creatinine|Tryptophan/Creatinine
C0942031|T201|COMP|25995-2|LNC|Tyrosine|Tyrosine
C0942032|T201|COMP|25997-8|LNC|Urate|Urate
C0942033|T201|COMP|25998-6|LNC|Urea|Urea
C0942034|T201|COMP|25999-4|LNC|Urea/Creatinine|Urea/Creatinine
C0942035|T201|COMP|26000-0|LNC|Uroporphyrin|Uroporphyrin
C0942036|T201|COMP|26001-8|LNC|Valine|Valine
C0942037|T201|COMP|26003-4|LNC|Vanillylmandelate|Vanillylmandelate
C0942038|T201|COMP|26004-2|LNC|Vanillylmandelate/Creatinine|Vanillylmandelate/Creatinine
C0942039|T201|COMP|26005-9|LNC|Xylose^2H post dose xylose PO|Xylose^2H post dose xylose PO
C0942040|T201|COMP|26006-7|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0942041|T201|COMP|26008-3|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0942042|T201|COMP|26009-1|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C0942044|T201|COMP|26012-5|LNC|17-Hydroxycorticosteroids^1D post XXX challenge|17-Hydroxycorticosteroids^1D post XXX challenge
C0942045|T201|COMP|26013-3|LNC|17-Hydroxycorticosteroids^2D post XXX challenge|17-Hydroxycorticosteroids^2D post XXX challenge
C0942046|T201|COMP|26014-1|LNC|Arbovirus NOS Ab|Arbovirus NOS Ab
C0942047|T201|COMP|26015-8|LNC|Cholesterol.in HDL 2|Cholesterol.in HDL 2
C0942048|T201|COMP|26017-4|LNC|Cholesterol.in HDL 3|Cholesterol.in HDL 3
C0942051|T201|COMP|26021-6|LNC|Nordiazepam|Nordiazepam
C0942052|T201|COMP|26022-4|LNC|Enterovirus NOS Ab|Enterovirus NOS Ab
C0942053|T201|COMP|26023-2|LNC|Extractable nuclear Ab identified|Extractable nuclear Ab identified
C0942054|T201|COMP|26024-0|LNC|Gastrin^post meal|Gastrin^post meal
C0942055|T201|COMP|26026-5|LNC|Hexahydrophthalic anhydride Ab.IgE.RAST class|Hexahydrophthalic anhydride Ab.IgE.RAST class
C0942056|T201|COMP|26027-3|LNC|Histiocytes|Histiocytes
C0942057|T201|COMP|26028-1|LNC|HLA-B27|HLA-B27
C0942058|T201|COMP|26029-9|LNC|Lactoferrin bovine Ab.IgE|Lactoferrin bovine Ab.IgE
C0942059|T201|COMP|26030-7|LNC|Lactoferrin bovine Ab.IgE.RAST class|Lactoferrin bovine Ab.IgE.RAST class
C0942060|T201|COMP|26031-5|LNC|Sialate.lipid bound|Sialate.lipid bound
C0942061|T201|COMP|26032-3|LNC|Pepsin Ab.IgE.RAST class|Pepsin Ab.IgE.RAST class
C0942062|T201|COMP|26033-1|LNC|Pronormoblasts/100 cells|Pronormoblasts/100 cells
C0942063|T201|COMP|26034-9|LNC|Protein|Protein
C0942064|T201|COMP|26035-6|LNC|Serotonin|Serotonin
C0942066|T201|COMP|26037-2|LNC|Trichophyton mentagrophytes var goetzii Ab.IgE|Trichophyton mentagrophytes var goetzii Ab.IgE
C0942067|T201|COMP|26040-6|LNC|Norcitalopram|Norcitalopram
C0942068|T201|COMP|26041-4|LNC|Normephenytoin|Normephenytoin
C0942069|T201|COMP|26042-2|LNC|Didesmethylcitalopram|Didesmethylcitalopram
C0942070|T201|COMP|26043-0|LNC|HLA-B27|HLA-B27
C0942071|T201|COMP|26044-8|LNC|Pepsin Ab.IgE|Pepsin Ab.IgE
C0942072|T201|COMP|26045-5|LNC|Pheneturide|Pheneturide
C0942073|T201|COMP|26046-3|LNC|5-Hydroxypropafenone|5-Hydroxypropafenone
C0942074|T201|COMP|26047-1|LNC|Phytate|Phytate
C0942075|T201|COMP|26048-9|LNC|Canary serum proteins Ab.IgE.RAST class|Canary serum proteins Ab.IgE.RAST class
C0942076|T201|COMP|26049-7|LNC|Libocedrus decurrens Ab.IgE|Libocedrus decurrens Ab.IgE
C0942077|T201|COMP|26050-5|LNC|Libocedrus decurrens Ab.IgE.RAST class|Libocedrus decurrens Ab.IgE.RAST class
C0942078|T201|COMP|26051-3|LNC|Epithelial cells.extrarenal|Epithelial cells.extrarenal
C0942079|T201|COMP|26052-1|LNC|Epithelial cells.renal|Epithelial cells.renal
C0942080|T201|COMP|26054-7|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C0942081|T201|COMP|26055-4|LNC|Pyridoxine^pre 250 mg pyridoxine PO|Pyridoxine^pre 250 mg pyridoxine PO
C0942082|T201|COMP|26056-2|LNC|Pyridoxine^post 250 mg pyridoxine PO|Pyridoxine^post 250 mg pyridoxine PO
C0942083|T201|COMP|26058-8|LNC|European tick borne encephalitis virus Ab|European tick borne encephalitis virus Ab
C0942084|T201|COMP|26059-6|LNC|European tick borne encephalitis virus Ab.IgG|European tick borne encephalitis virus Ab.IgG
C0942085|T201|COMP|26060-4|LNC|European tick borne encephalitis virus Ab.IgM|European tick borne encephalitis virus Ab.IgM
C0942086|T201|COMP|26061-2|LNC|European tick borne encephalitis virus Ab|European tick borne encephalitis virus Ab
C0942087|T201|COMP|26063-8|LNC|European tick borne encephalitis virus Ab.IgM|European tick borne encephalitis virus Ab.IgM
C0942378|T201|COMP|26403-6|LNC|Alternaria alternata Ab.IgG4|Alternaria alternata Ab.IgG4
C0942379|T201|COMP|26404-4|LNC|Alternaria alternata Ab.IgG4.RAST class|Alternaria alternata Ab.IgG4.RAST class
C0942380|T201|COMP|26406-9|LNC|Aspergillus fumigatus Ab.IgG4.RAST class|Aspergillus fumigatus Ab.IgG4.RAST class
C0942381|T201|COMP|26407-7|LNC|Apis mellifera Ab.IgG4|Apis mellifera Ab.IgG4
C0942382|T201|COMP|26408-5|LNC|Apis mellifera Ab.IgG4.RAST class|Apis mellifera Ab.IgG4.RAST class
C0942383|T201|COMP|26409-3|LNC|Betula verrucosa Ab.IgG4|Betula verrucosa Ab.IgG4
C0942384|T201|COMP|26410-1|LNC|Betula verrucosa Ab.IgG4.RAST class|Betula verrucosa Ab.IgG4.RAST class
C0942385|T201|COMP|26411-9|LNC|Bran wheat Ab.IgG4|Bran wheat Ab.IgG4
C0942386|T201|COMP|26412-7|LNC|Bran wheat Ab.IgG4.RAST class|Bran wheat Ab.IgG4.RAST class
C0942387|T201|COMP|26413-5|LNC|Candida albicans Ab.IgG4|Candida albicans Ab.IgG4
C0942388|T201|COMP|26415-0|LNC|Casein Ab.IgG4|Casein Ab.IgG4
C0942389|T201|COMP|26416-8|LNC|Casein Ab.IgG4.RAST class|Casein Ab.IgG4.RAST class
C0942390|T201|COMP|26417-6|LNC|Cladosporium herbarum Ab.IgG4|Cladosporium herbarum Ab.IgG4
C0942391|T201|COMP|26418-4|LNC|Cladosporium herbarum Ab.IgG4.RAST class|Cladosporium herbarum Ab.IgG4.RAST class
C0942392|T201|COMP|26419-2|LNC|Dermatophagoides farinae Ab.IgG4|Dermatophagoides farinae Ab.IgG4
C0942393|T201|COMP|26420-0|LNC|Dermatophagoides farinae Ab.IgG4.RAST class|Dermatophagoides farinae Ab.IgG4.RAST class
C0942394|T201|COMP|26421-8|LNC|Dermatophagoides pteronyssinus Ab.IgG4|Dermatophagoides pteronyssinus Ab.IgG4
C0942395|T201|COMP|26422-6|LNC|Dermatophagoides pteronyssinus Ab.IgG4.RAST class|Dermatophagoides pteronyssinus Ab.IgG4.RAST class
C0942396|T201|COMP|26423-4|LNC|Egg white Ab.IgG4|Egg white Ab.IgG4
C0942397|T201|COMP|26424-2|LNC|Egg white Ab.IgG4.RAST class|Egg white Ab.IgG4.RAST class
C0942398|T201|COMP|26425-9|LNC|Lactalbumin alpha Ab.IgG4|Lactalbumin alpha Ab.IgG4
C0942399|T201|COMP|26427-5|LNC|Lactoglobulin Ab.IgG4|Lactoglobulin Ab.IgG4
C0942400|T201|COMP|26428-3|LNC|Oryza sativa Ab.IgG4|Oryza sativa Ab.IgG4
C0942401|T201|COMP|26430-9|LNC|Phleum pratense Ab.IgG4|Phleum pratense Ab.IgG4
C0942402|T201|COMP|26431-7|LNC|Phleum pratense Ab.IgG4.RAST class|Phleum pratense Ab.IgG4.RAST class
C0942403|T201|COMP|26432-5|LNC|Wasp venom Ab.IgG4|Wasp venom Ab.IgG4
C0942404|T201|COMP|26433-3|LNC|Wasp venom Ab.IgG4.RAST class|Wasp venom Ab.IgG4.RAST class
C0942405|T201|COMP|26434-1|LNC|Lactoglobulin Ab.IgG4.RAST class|Lactoglobulin Ab.IgG4.RAST class
C0942414|T201|COMP|26444-0|LNC|Basophils|Basophils
C0942415|T201|COMP|26445-7|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0942416|T201|COMP|26446-5|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C0942417|T201|COMP|26447-3|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C0942418|T201|COMP|26448-1|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C0942419|T201|COMP|26449-9|LNC|Eosinophils|Eosinophils
C0942420|T201|COMP|26451-5|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0942421|T201|COMP|26452-3|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0942422|T201|COMP|26453-1|LNC|Erythrocytes|Erythrocytes
C0942423|T201|COMP|26454-9|LNC|Erythrocytes|Erythrocytes
C0942424|T201|COMP|26456-4|LNC|Erythrocytes|Erythrocytes
C0942425|T201|COMP|26457-2|LNC|Erythrocytes|Erythrocytes
C0942426|T201|COMP|26458-0|LNC|Erythrocytes|Erythrocytes
C0942427|T201|COMP|26460-6|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C0942428|T201|COMP|26462-2|LNC|Large unstained cells|Large unstained cells
C0942429|T201|COMP|26463-0|LNC|Large unstained cells/100 leukocytes|Large unstained cells/100 leukocytes
C0942430|T201|COMP|26465-5|LNC|Leukocytes|Leukocytes
C0942431|T201|COMP|26466-3|LNC|Leukocytes|Leukocytes
C0942432|T201|COMP|26467-1|LNC|Leukocytes|Leukocytes
C0942433|T201|COMP|26469-7|LNC|Leukocytes|Leukocytes
C0942434|T201|COMP|26470-5|LNC|Leukocytes other|Leukocytes other
C0942435|T201|COMP|26472-1|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0942436|T201|COMP|26473-9|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0942437|T201|COMP|26474-7|LNC|Lymphocytes|Lymphocytes
C0942438|T201|COMP|26475-4|LNC|Lymphocytes|Lymphocytes
C0942439|T201|COMP|26476-2|LNC|Lymphocytes|Lymphocytes
C0942440|T201|COMP|26478-8|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0942441|T201|COMP|26479-6|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0942442|T201|COMP|26480-4|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0942443|T201|COMP|26481-2|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0942444|T201|COMP|26482-0|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0942445|T201|COMP|26483-8|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0942446|T201|COMP|26484-6|LNC|Monocytes|Monocytes
C0942447|T201|COMP|26485-3|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0942448|T201|COMP|26486-1|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0942449|T201|COMP|26487-9|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0942450|T201|COMP|26488-7|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0942451|T201|COMP|26489-5|LNC|Mononuclear cells|Mononuclear cells
C0942452|T201|COMP|26490-3|LNC|Mononuclear cells|Mononuclear cells
C0942453|T201|COMP|26491-1|LNC|Mononuclear cells|Mononuclear cells
C0942454|T201|COMP|26492-9|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0942455|T201|COMP|26493-7|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0942456|T201|COMP|26494-5|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0942457|T201|COMP|26495-2|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0942458|T201|COMP|26496-0|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0942459|T201|COMP|26497-8|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C0942460|T201|COMP|26498-6|LNC|Myelocytes/100 leukocytes|Myelocytes/100 leukocytes
C0942461|T201|COMP|26499-4|LNC|Neutrophils|Neutrophils
C0942462|T201|COMP|26500-9|LNC|Neutrophils|Neutrophils
C0942463|T201|COMP|26501-7|LNC|Neutrophils|Neutrophils
C0942464|T201|COMP|26502-5|LNC|Neutrophils|Neutrophils
C0942465|T201|COMP|26503-3|LNC|Neutrophils|Neutrophils
C0942466|T201|COMP|26505-8|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C0942467|T201|COMP|26506-6|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C0942468|T201|COMP|26508-2|LNC|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0942469|T201|COMP|26509-0|LNC|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0942470|T201|COMP|26510-8|LNC|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0942471|T201|COMP|26511-6|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0942472|T201|COMP|32709-8|LNC|Neutrophils|Neutrophils
C0942473|T201|COMP|26514-0|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0942474|T201|COMP|26515-7|LNC|Platelets|Platelets
C0942475|T201|COMP|26516-5|LNC|Platelets|Platelets
C0942476|T201|COMP|26518-1|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0942477|T201|COMP|26519-9|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0942478|T201|COMP|26520-7|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0942479|T201|COMP|26521-5|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0942480|T201|COMP|26523-1|LNC|Promyelocytes|Promyelocytes
C0942482|T201|COMP|26525-6|LNC|Cortisol.free^24H post dose corticotropin|Cortisol.free^24H post dose corticotropin
C0942483|T201|COMP|26526-4|LNC|Cortisol.free^48H post dose corticotropin|Cortisol.free^48H post dose corticotropin
C0942484|T201|COMP|26528-0|LNC|Cortisol^1H post dose corticotropin|Cortisol^1H post dose corticotropin
C0942485|T201|COMP|26529-8|LNC|Cortisol^24H post dose corticotropin|Cortisol^24H post dose corticotropin
C0942486|T201|COMP|26530-6|LNC|Cortisol^30M post dose corticotropin|Cortisol^30M post dose corticotropin
C0942487|T201|COMP|26531-4|LNC|Cortisol^32H post dose corticotropin|Cortisol^32H post dose corticotropin
C0942488|T201|COMP|26534-8|LNC|Cortisol^8H post dose corticotropin|Cortisol^8H post dose corticotropin
C0942489|T201|COMP|26535-5|LNC|Cortisol^30M post dose corticotropin|Cortisol^30M post dose corticotropin
C0942490|T201|COMP|26536-3|LNC|Cortisol^1H post dose corticotropin|Cortisol^1H post dose corticotropin
C0942491|T201|COMP|26537-1|LNC|Glucose^2.5H post dose glucose|Glucose^2.5H post dose glucose
C0942492|T201|COMP|26539-7|LNC|Glucose^45M post dose glucose|Glucose^45M post dose glucose
C0942493|T201|COMP|26540-5|LNC|Glucose^3H post dose glucose|Glucose^3H post dose glucose
C0942494|T201|COMP|26541-3|LNC|Glucose^4H post dose glucose|Glucose^4H post dose glucose
C0942495|T201|COMP|26542-1|LNC|Glucose^5H post dose glucose|Glucose^5H post dose glucose
C0942496|T201|COMP|26543-9|LNC|Glucose^5H post dose glucose|Glucose^5H post dose glucose
C0942497|T201|COMP|26544-7|LNC|Glucose^6H post dose glucose|Glucose^6H post dose glucose
C0942498|T201|COMP|26545-4|LNC|Glucose^6H post dose glucose|Glucose^6H post dose glucose
C0942499|T201|COMP|26546-2|LNC|Glucose^1H post dose glucose|Glucose^1H post dose glucose
C0942500|T201|COMP|26547-0|LNC|Glucose^2H post dose glucose|Glucose^2H post dose glucose
C0942501|T201|COMP|26548-8|LNC|Glucose^30M post dose glucose|Glucose^30M post dose glucose
C0942502|T201|COMP|26549-6|LNC|Glucose^3H post dose glucose|Glucose^3H post dose glucose
C0942503|T201|COMP|26550-4|LNC|Glucose^4H post dose glucose|Glucose^4H post dose glucose
C0942504|T201|COMP|26551-2|LNC|Glucose^5H post dose glucose|Glucose^5H post dose glucose
C0942505|T201|COMP|26552-0|LNC|Glucose^6H post dose glucose|Glucose^6H post dose glucose
C0942506|T201|COMP|26554-6|LNC|Glucose^2.5H post dose glucose|Glucose^2.5H post dose glucose
C0942507|T201|COMP|26555-3|LNC|Glucose^3.5H post dose glucose|Glucose^3.5H post dose glucose
C0942508|T201|COMP|26557-9|LNC|Cells.CD11b+CD56+/100 cells|Cells.CD11b+CD56+/100 cells
C0942509|T201|COMP|26558-7|LNC|Cells.CD11c+CD25+/100 cells|Cells.CD11c+CD25+/100 cells
C0942510|T201|COMP|26559-5|LNC|Cells.CD38+CD56+/100 cells|Cells.CD38+CD56+/100 cells
C0942511|T201|COMP|26560-3|LNC|Cells.CD16/100 cells|Cells.CD16/100 cells
C0942512|T201|COMP|26561-1|LNC|Cells.CD16+CD56+|Cells.CD16+CD56+
C0942513|T201|COMP|26562-9|LNC|Cells.CD19+CD38+/100 cells|Cells.CD19+CD38+/100 cells
C0942514|T201|COMP|26563-7|LNC|Cells.CD1a/100 cells|Cells.CD1a/100 cells
C0942515|T201|COMP|26564-5|LNC|Cells.CD30|Cells.CD30
C0942516|T201|COMP|26565-2|LNC|Cells.CD19+Kappa+/100 cells|Cells.CD19+Kappa+/100 cells
C0942517|T201|COMP|26566-0|LNC|Cells.CD19+Lambda+/100 cells|Cells.CD19+Lambda+/100 cells
C0942518|T201|COMP|26567-8|LNC|Lymphocytes.IgA/100 lymphocytes|Lymphocytes.IgA/100 lymphocytes
C0942519|T201|COMP|26568-6|LNC|Cells.CD3+HLA-DR+|Cells.CD3+HLA-DR+
C0942520|T201|COMP|26569-4|LNC|Cells.CD4+CD29+|Cells.CD4+CD29+
C0942521|T201|COMP|26570-2|LNC|Cells.CD4+CD45+|Cells.CD4+CD45+
C0942522|T201|COMP|33586-9|LNC|Cells.CD2+CD7+|Cells.CD2+CD7+
C0942523|T201|COMP|26573-6|LNC|Cells.CD4+CD45+/100 cells|Cells.CD4+CD45+/100 cells
C0942524|T201|COMP|26574-4|LNC|1-Methylhistidine/Creatinine|1-Methylhistidine/Creatinine
C0942525|T201|COMP|26575-1|LNC|3-Methylhistidine/Creatinine|3-Methylhistidine/Creatinine
C0942526|T201|COMP|26577-7|LNC|Asparagine/Creatinine|Asparagine/Creatinine
C0942527|T201|COMP|26578-5|LNC|Beta alanine/Creatinine|Beta alanine/Creatinine
C0942529|T201|COMP|26581-9|LNC|Gamma aminobutyrate/Creatinine|Gamma aminobutyrate/Creatinine
C0942530|T201|COMP|26582-7|LNC|Homocysteine/Creatinine|Homocysteine/Creatinine
C0942531|T201|COMP|26583-5|LNC|3-Hydroxy,3-Methylglutarate/Creatinine|3-Hydroxy,3-Methylglutarate/Creatinine
C0942532|T201|COMP|26585-0|LNC|3-Methylhistidine|3-Methylhistidine
C0942533|T201|COMP|26587-6|LNC|Alpha aminoadipate|Alpha aminoadipate
C0942534|T201|COMP|26588-4|LNC|Anserine|Anserine
C0942535|T201|COMP|26590-0|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0942536|T201|COMP|26591-8|LNC|Carnosine|Carnosine
C0942537|T201|COMP|26594-2|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0942538|T201|COMP|26595-9|LNC|Hydroxylysine|Hydroxylysine
C0942539|T201|COMP|26596-7|LNC|Hydroxyproline|Hydroxyproline
C0942540|T201|COMP|26598-3|LNC|Sarcosine|Sarcosine
C0942541|T201|COMP|26599-1|LNC|Anserine|Anserine
C0942542|T201|COMP|26600-7|LNC|Alpha aminoadipate|Alpha aminoadipate
C0942543|T201|COMP|26601-5|LNC|Alpha aminoadipate/Creatinine|Alpha aminoadipate/Creatinine
C0942544|T201|COMP|26602-3|LNC|Tryptophan|Tryptophan
C0942545|T201|COMP|26603-1|LNC|Asparagine|Asparagine
C0942546|T201|COMP|26604-9|LNC|Beta alanine|Beta alanine
C0942547|T201|COMP|26605-6|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0942548|T201|COMP|26606-4|LNC|Carnosine|Carnosine
C0942549|T201|COMP|26607-2|LNC|Cystathionine|Cystathionine
C0942550|T201|COMP|26608-0|LNC|Ethanolamine|Ethanolamine
C0942551|T201|COMP|26609-8|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0942552|T201|COMP|26610-6|LNC|Hydroxylysine|Hydroxylysine
C0942553|T201|COMP|26611-4|LNC|Phosphoethanolamine|Phosphoethanolamine
C0942554|T201|COMP|26612-2|LNC|Phosphoethanolamine|Phosphoethanolamine
C0942555|T201|COMP|26613-0|LNC|Sarcosine|Sarcosine
C0942556|T201|COMP|26614-8|LNC|Taurine|Taurine
C0942557|T201|COMP|26615-5|LNC|Erythrocytes.CD55|Erythrocytes.CD55
C0942558|T201|COMP|26616-3|LNC|Erythrocytes.CD59|Erythrocytes.CD59
C0942559|T201|COMP|26617-1|LNC|Trypanosoma brucei gambiense Ab|Trypanosoma brucei gambiense Ab
C0942560|T201|COMP|26619-7|LNC|Campylobacter sp Ab|Campylobacter sp Ab
C0942561|T201|COMP|26620-5|LNC|Hantavirus Ab.IgG|Hantavirus Ab.IgG
C0942562|T201|COMP|26622-1|LNC|Babesia duncani Ab|Babesia duncani Ab
C0942563|T201|COMP|26623-9|LNC|Chikungunya virus Ab|Chikungunya virus Ab
C0942564|T201|COMP|26624-7|LNC|Rickettsia conorii Ab|Rickettsia conorii Ab
C0942565|T201|COMP|26625-4|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C0942566|T201|COMP|26626-2|LNC|Chlamydia trachomatis L2 Ab|Chlamydia trachomatis L2 Ab
C0942567|T201|COMP|26627-0|LNC|Legionella polyvalent A Ab|Legionella polyvalent A Ab
C0942568|T201|COMP|26628-8|LNC|Legionella polyvalent B Ab|Legionella polyvalent B Ab
C0942569|T201|COMP|26629-6|LNC|Legionella polyvalent C Ab|Legionella polyvalent C Ab
C0942570|T201|COMP|26630-4|LNC|Corynebacterium diphtheriae toxin Ab|Corynebacterium diphtheriae toxin Ab
C0942571|T201|COMP|26631-2|LNC|Borrelia hermsii Ab|Borrelia hermsii Ab
C0942572|T201|COMP|26632-0|LNC|Legionella dumoffii Ab|Legionella dumoffii Ab
C0942573|T201|COMP|26633-8|LNC|Legionella bozemaniae Ab|Legionella bozemaniae Ab
C0942574|T201|COMP|26634-6|LNC|Legionella gormanii Ab|Legionella gormanii Ab
C0942575|T201|COMP|26636-1|LNC|Candida sp Ab|Candida sp Ab
C0942576|T201|COMP|26637-9|LNC|Leishmania braziliensis Ab|Leishmania braziliensis Ab
C0942577|T201|COMP|26638-7|LNC|Leishmania donovani Ab|Leishmania donovani Ab
C0942578|T201|COMP|26639-5|LNC|Leishmania tropica Ab|Leishmania tropica Ab
C0942579|T201|COMP|26640-3|LNC|Paracoccidioides brasiliensis Ab|Paracoccidioides brasiliensis Ab
C0942580|T201|COMP|26641-1|LNC|Histoplasma sp Ab|Histoplasma sp Ab
C0942581|T201|COMP|26642-9|LNC|Jamestown canyon virus Ab|Jamestown canyon virus Ab
C0942582|T201|COMP|26644-5|LNC|Getah virus Ab|Getah virus Ab
C0942583|T201|COMP|26645-2|LNC|BK virus Ab|BK virus Ab
C0942584|T201|COMP|26646-0|LNC|Powassan virus Ab|Powassan virus Ab
C0942585|T201|COMP|26647-8|LNC|Semliki forest virus Ab|Semliki forest virus Ab
C0942586|T201|COMP|26649-4|LNC|Snowshoe hare virus Ab|Snowshoe hare virus Ab
C0942587|T201|COMP|26650-2|LNC|Hantavirus sin nombre Ab.IgM|Hantavirus sin nombre Ab.IgM
C0942588|T201|COMP|26653-6|LNC|Colorado tick fever virus Ab|Colorado tick fever virus Ab
C0942589|T201|COMP|26654-4|LNC|Hantavirus sin nombre Ab.IgG|Hantavirus sin nombre Ab.IgG
C0942590|T201|COMP|26657-7|LNC|Schistosoma haematobium Ab|Schistosoma haematobium Ab
C0942591|T201|COMP|26658-5|LNC|Treponema sp Ab|Treponema sp Ab
C0942592|T201|COMP|26659-3|LNC|Leptospira autumnalis Ab|Leptospira autumnalis Ab
C0942593|T201|COMP|26661-9|LNC|Trichinella sp Ab|Trichinella sp Ab
C0942594|T201|COMP|26662-7|LNC|Bebaru virus Ab|Bebaru virus Ab
C0942595|T201|COMP|26663-5|LNC|Chlamydia trachomatis D Ab|Chlamydia trachomatis D Ab
C0942596|T201|COMP|26665-0|LNC|Chlamydia trachomatis F Ab|Chlamydia trachomatis F Ab
C0942597|T201|COMP|26666-8|LNC|Chlamydia trachomatis H Ab|Chlamydia trachomatis H Ab
C0942598|T201|COMP|26667-6|LNC|Chlamydia trachomatis I Ab|Chlamydia trachomatis I Ab
C0942599|T201|COMP|26668-4|LNC|Chlamydia trachomatis L1 Ab|Chlamydia trachomatis L1 Ab
C0942600|T201|COMP|26669-2|LNC|Absidia corymbifera Ab|Absidia corymbifera Ab
C0942601|T201|COMP|26670-0|LNC|Rhizomucor pusillus Ab|Rhizomucor pusillus Ab
C0942602|T201|COMP|26671-8|LNC|Ascaris sp Ab|Ascaris sp Ab
C0942603|T201|COMP|26672-6|LNC|Ross river virus Ab|Ross river virus Ab
C0942604|T201|COMP|26673-4|LNC|Echinococcus granulosus Ab|Echinococcus granulosus Ab
C0942605|T201|COMP|26674-2|LNC|Legionella longbeachae 1 Ab|Legionella longbeachae 1 Ab
C0942606|T201|COMP|26675-9|LNC|Legionella longbeachae 2 Ab|Legionella longbeachae 2 Ab
C0942607|T201|COMP|26676-7|LNC|Bartonella henselae Ab|Bartonella henselae Ab
C0942608|T201|COMP|26678-3|LNC|Bartonella elizabethae Ab|Bartonella elizabethae Ab
C0942609|T201|COMP|26679-1|LNC|Secobarbital|Secobarbital
C0942610|T201|COMP|26681-7|LNC|Streptococcus pneumoniae 23 Ab|Streptococcus pneumoniae 23 Ab
C0942611|T201|COMP|26682-5|LNC|Glycolate|Glycolate
C0942612|T201|COMP|26683-3|LNC|Estazolam|Estazolam
C0942613|T201|COMP|26684-1|LNC|Mycoplasma pneumoniae Ab.IgA|Mycoplasma pneumoniae Ab.IgA
C0942614|T201|COMP|26685-8|LNC|3-Hydroxyisovalerate|3-Hydroxyisovalerate
C0942615|T201|COMP|26686-6|LNC|Triazolam|Triazolam
C0942616|T201|COMP|26687-4|LNC|Amobarbital|Amobarbital
C0942617|T201|COMP|26688-2|LNC|Mercury/Creatinine|Mercury/Creatinine
C0942618|T201|COMP|26689-0|LNC|Butabarbital|Butabarbital
C0942619|T201|COMP|26690-8|LNC|Western equine encephalitis virus RNA|Western equine encephalitis virus RNA
C0942620|T201|COMP|26691-6|LNC|Uroporphyrin 1 isomer|Uroporphyrin 1 isomer
C0942621|T201|COMP|26692-4|LNC|Streptococcus pneumoniae 19 Ab|Streptococcus pneumoniae 19 Ab
C0942622|T201|COMP|26693-2|LNC|Streptococcus pneumoniae 12f Ab|Streptococcus pneumoniae 12f Ab
C0942623|T201|COMP|26694-0|LNC|Clostridioides difficile Ab.IgM|Clostridioides difficile Ab.IgM
C0942624|T201|COMP|26695-7|LNC|Glucose^7th specimen post XXX challenge|Glucose^7th specimen post XXX challenge
C0942625|T201|COMP|26696-5|LNC|Morphine.free|Morphine.free
C0942626|T201|COMP|26697-3|LNC|Clostridioides difficile Ab.IgA|Clostridioides difficile Ab.IgA
C0942627|T201|COMP|26698-1|LNC|Listeria monocytogenes Ab.IgG|Listeria monocytogenes Ab.IgG
C0942628|T201|COMP|26699-9|LNC|Indicans|Indicans
C0942631|T201|COMP|26704-7|LNC|Isospora belli|Isospora belli
C0942632|T201|COMP|26706-2|LNC|Vanillylmandelate|Vanillylmandelate
C0942633|T201|COMP|26708-8|LNC|Magnesium|Magnesium
C0942634|T201|COMP|26710-4|LNC|Leucine|Leucine
C0942635|T201|COMP|26712-0|LNC|Phenmetrazine|Phenmetrazine
C0942636|T201|COMP|26713-8|LNC|Phentermine|Phentermine
C0942637|T201|COMP|26714-6|LNC|Phenylpropanolamine|Phenylpropanolamine
C0942638|T201|COMP|26716-1|LNC|Chlorphentermine|Chlorphentermine
C0942639|T201|COMP|26717-9|LNC|Phosphoethanolamine|Phosphoethanolamine
C0942640|T201|COMP|26718-7|LNC|HYDROmorphone|HYDROmorphone
C0942641|T201|COMP|26719-5|LNC|HYDROcodone|HYDROcodone
C0942642|T201|COMP|26720-3|LNC|Codeine|Codeine
C0942643|T201|COMP|26721-1|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0942644|T201|COMP|26722-9|LNC|oxyCODONE|oxyCODONE
C0942645|T201|COMP|26723-7|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C0942646|T201|COMP|26725-2|LNC|Alpha aminoadipate|Alpha aminoadipate
C0942647|T201|COMP|26726-0|LNC|Proline|Proline
C0942648|T201|COMP|26727-8|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C0942649|T201|COMP|26729-4|LNC|Ovary Ab.IgG|Ovary Ab.IgG
C0942650|T201|COMP|26730-2|LNC|Isoleucine|Isoleucine
C0942651|T201|COMP|26731-0|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0942652|T201|COMP|26732-8|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0942653|T201|COMP|26733-6|LNC|Butabarbital|Butabarbital
C0942654|T201|COMP|26734-4|LNC|Methamphetamine|Methamphetamine
C0942655|T201|COMP|26735-1|LNC|Rhodococcus equi Ab|Rhodococcus equi Ab
C0942656|T201|COMP|26736-9|LNC|Promethazine|Promethazine
C0942657|T201|COMP|26737-7|LNC|Phosphoserine|Phosphoserine
C0942658|T201|COMP|26738-5|LNC|Phosphoserine|Phosphoserine
C0942659|T201|COMP|26739-3|LNC|Xylose^4th specimen post XXX challenge|Xylose^4th specimen post XXX challenge
C0942660|T201|COMP|26740-1|LNC|Hydroxyproline|Hydroxyproline
C0942661|T201|COMP|26741-9|LNC|Serine|Serine
C0942662|T201|COMP|26742-7|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0942663|T201|COMP|26743-5|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0942664|T201|COMP|26744-3|LNC|Opiates|Opiates
C0942665|T201|COMP|26745-0|LNC|Citrulline|Citrulline
C0942666|T201|COMP|26746-8|LNC|Magnesium|Magnesium
C0942667|T201|COMP|26747-6|LNC|Cannabinoids/Creatinine|Cannabinoids/Creatinine
C0942668|T201|COMP|26748-4|LNC|Osmium|Osmium
C0942669|T201|COMP|26750-0|LNC|Carnosine|Carnosine
C0942670|T201|COMP|26751-8|LNC|Adipate|Adipate
C0942671|T201|COMP|26752-6|LNC|Creatinine renal clearance|Creatinine renal clearance
C0942672|T201|COMP|26753-4|LNC|Carnitine esters|Carnitine esters
C0942673|T201|COMP|26754-2|LNC|Streptococcus pneumoniae Danish serotype 7F Ab|Streptococcus pneumoniae Danish serotype 7F Ab
C0942674|T201|COMP|26755-9|LNC|Streptococcus pneumoniae Danish serotype 18C Ab|Streptococcus pneumoniae Danish serotype 18C Ab
C0942675|T201|COMP|26756-7|LNC|Isoniazid|Isoniazid
C0942676|T201|COMP|26757-5|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C0942677|T201|COMP|26758-3|LNC|Cocaine|Cocaine
C0942678|T201|COMP|26759-1|LNC|Cells.CD4+CD45RA+|Cells.CD4+CD45RA+
C0942679|T201|COMP|26761-7|LNC|Sodium renal clearance|Sodium renal clearance
C0942680|T201|COMP|26762-5|LNC|Chloride|Chloride
C0942681|T201|COMP|26763-3|LNC|Sodium|Sodium
C0942682|T201|COMP|26764-1|LNC|Cannabinoids|Cannabinoids
C0942683|T201|COMP|26766-6|LNC|Bacteroides fragilis Ab.IgG|Bacteroides fragilis Ab.IgG
C0942684|T201|COMP|26767-4|LNC|Clostridium perfringens Ab.IgG|Clostridium perfringens Ab.IgG
C0942685|T201|COMP|26768-2|LNC|Clostridium perfringens Ab.IgM|Clostridium perfringens Ab.IgM
C0942686|T201|COMP|26770-8|LNC|Trichloroacetate/Creatinine|Trichloroacetate/Creatinine
C0942687|T201|COMP|26771-6|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C0942688|T201|COMP|26773-2|LNC|Benzfetamine|Benzfetamine
C0942689|T201|COMP|26774-0|LNC|Flurazepam|Flurazepam
C0942690|T201|COMP|26775-7|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C0942691|T201|COMP|26776-5|LNC|QUEtiapine|QUEtiapine
C0942692|T201|COMP|26778-1|LNC|Glucose^1H post dose lactose PO|Glucose^1H post dose lactose PO
C0942693|T201|COMP|26780-7|LNC|Glucose^2H post dose lactose PO|Glucose^2H post dose lactose PO
C0942694|T201|COMP|26783-1|LNC|Glucose^5H post dose lactose PO|Glucose^5H post dose lactose PO
C0942695|T201|COMP|26784-9|LNC|diazePAM|diazePAM
C0942696|T201|COMP|26785-6|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C0942697|T201|COMP|26787-2|LNC|Anserine|Anserine
C0942698|T201|COMP|26788-0|LNC|Carnitine|Carnitine
C0942699|T201|COMP|26789-8|LNC|Escherichia coli Ab.IgM|Escherichia coli Ab.IgM
C0942700|T201|COMP|26791-4|LNC|Amphetamine|Amphetamine
C0942701|T201|COMP|26792-2|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0942702|T201|COMP|26793-0|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0942703|T201|COMP|26795-5|LNC|Alanine|Alanine
C0942704|T201|COMP|26796-3|LNC|Oxalate|Oxalate
C0942705|T201|COMP|26797-1|LNC|Alpha hydroxybutyrate|Alpha hydroxybutyrate
C0942706|T201|COMP|26798-9|LNC|Succinate|Succinate
C0942707|T201|COMP|26799-7|LNC|Fumarate|Fumarate
C0942708|T201|COMP|26800-3|LNC|Escherichia coli Ab.IgG|Escherichia coli Ab.IgG
C0942709|T201|COMP|26801-1|LNC|Protein|Protein
C0942710|T201|COMP|26802-9|LNC|Midazolam|Midazolam
C0942711|T201|COMP|26803-7|LNC|Ethanolamine|Ethanolamine
C0942712|T201|COMP|26804-5|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0942713|T201|COMP|26805-2|LNC|Glutamate|Glutamate
C0942714|T201|COMP|26806-0|LNC|Glutamine|Glutamine
C0942715|T201|COMP|26807-8|LNC|Glycine|Glycine
C0942716|T201|COMP|26808-6|LNC|Histidine|Histidine
C0942717|T201|COMP|26809-4|LNC|Homocystine|Homocystine
C0942718|T201|COMP|26810-2|LNC|Hydroxyproline|Hydroxyproline
C0942719|T201|COMP|26811-0|LNC|2-Methylcitrate|2-Methylcitrate
C0942720|T201|COMP|26813-6|LNC|Acidity.titratable|Acidity.titratable
C0942721|T201|COMP|26814-4|LNC|IgG.monoclonal|IgG.monoclonal
C0942722|T201|COMP|26816-9|LNC|Nordiazepam|Nordiazepam
C0942723|T201|COMP|26817-7|LNC|Glucose^11H post XXX challenge|Glucose^11H post XXX challenge
C0942724|T201|COMP|26818-5|LNC|Campylobacter jejuni Ab|Campylobacter jejuni Ab
C0942725|T201|COMP|26819-3|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0942726|T201|COMP|26820-1|LNC|Stachybotrys chartarum Ab.IgA|Stachybotrys chartarum Ab.IgA
C0942727|T201|COMP|26821-9|LNC|Lipoprotein.beta|Lipoprotein.beta
C0942728|T201|COMP|26822-7|LNC|Lipoprotein.alpha|Lipoprotein.alpha
C0942729|T201|COMP|26823-5|LNC|Lutropin.beta subunit|Lutropin.beta subunit
C0942730|T201|COMP|26824-3|LNC|Phosphoserine|Phosphoserine
C0942731|T201|COMP|26825-0|LNC|Eastern equine encephalitis virus RNA|Eastern equine encephalitis virus RNA
C0942732|T201|COMP|26826-8|LNC|Testosterone|Testosterone
C0942733|T201|COMP|26827-6|LNC|Testosterone/Creatinine|Testosterone/Creatinine
C0942734|T201|COMP|26829-2|LNC|Phencyclidine|Phencyclidine
C0942735|T201|COMP|26830-0|LNC|Prochlorperazine|Prochlorperazine
C0942736|T201|COMP|26831-8|LNC|Suberate|Suberate
C0942737|T201|COMP|26833-4|LNC|Hippurate|Hippurate
C0942738|T201|COMP|26834-2|LNC|Temazepam|Temazepam
C0942739|T201|COMP|26835-9|LNC|Sebacate|Sebacate
C0942740|T201|COMP|26837-5|LNC|diazePAM|diazePAM
C0942741|T201|COMP|26838-3|LNC|LORazepam|LORazepam
C0942742|T201|COMP|26839-1|LNC|Oxazepam|Oxazepam
C0942743|T201|COMP|26841-7|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0942744|T201|COMP|26842-5|LNC|Iodine|Iodine
C0942745|T201|COMP|26843-3|LNC|Cystine|Cystine
C0942746|T201|COMP|26845-8|LNC|Sialate.lipid bound|Sialate.lipid bound
C0942747|T201|COMP|26847-4|LNC|Haloperidol|Haloperidol
C0942748|T201|COMP|26849-0|LNC|IgA.secretory|IgA.secretory
C0942749|T201|COMP|26850-8|LNC|Oxazepam|Oxazepam
C0942750|T201|COMP|26851-6|LNC|LORazepam|LORazepam
C0942751|T201|COMP|26853-2|LNC|Glucose^7th specimen post XXX challenge|Glucose^7th specimen post XXX challenge
C0942752|T201|COMP|26854-0|LNC|Glucose^8th specimen post XXX challenge|Glucose^8th specimen post XXX challenge
C0942753|T201|COMP|26855-7|LNC|Parainfluenza virus Ab|Parainfluenza virus Ab
C0942754|T201|COMP|26856-5|LNC|Cannabinoids|Cannabinoids
C0942755|T201|COMP|26858-1|LNC|Cells.CD3+CD56+|Cells.CD3+CD56+
C0942756|T201|COMP|26859-9|LNC|Phencyclidine|Phencyclidine
C0942757|T201|COMP|26861-5|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0942758|T201|COMP|26862-3|LNC|HYDROmorphone|HYDROmorphone
C0942759|T201|COMP|26863-1|LNC|HYDROcodone|HYDROcodone
C0942760|T201|COMP|26864-9|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C0942761|T201|COMP|26865-6|LNC|Codeine|Codeine
C0942762|T201|COMP|26866-4|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0942763|T201|COMP|26867-2|LNC|fentaNYL|fentaNYL
C0942764|T201|COMP|26868-0|LNC|Phenolphthalein|Phenolphthalein
C0942765|T201|COMP|26869-8|LNC|oxyCODONE|oxyCODONE
C0942766|T201|COMP|26870-6|LNC|Ganglioside GD1b Ab|Ganglioside GD1b Ab
C0942767|T201|COMP|26871-4|LNC|IgA|IgA
C0942768|T201|COMP|26872-2|LNC|Orotate|Orotate
C0942769|T201|COMP|26873-0|LNC|Valine|Valine
C0942770|T201|COMP|26874-8|LNC|Follitropin.beta subunit|Follitropin.beta subunit
C0942771|T201|COMP|26875-5|LNC|Streptococcus pneumoniae 4 Ab|Streptococcus pneumoniae 4 Ab
C0942772|T201|COMP|26876-3|LNC|Streptococcus pneumoniae 1 Ab|Streptococcus pneumoniae 1 Ab
C0942773|T201|COMP|26877-1|LNC|Hydroxytriazolam|Hydroxytriazolam
C0942774|T201|COMP|26878-9|LNC|ALPRAZolam|ALPRAZolam
C0942775|T201|COMP|26879-7|LNC|Triiodothyronine|Triiodothyronine
C0942776|T201|COMP|26881-3|LNC|Interleukin 6|Interleukin 6
C0942777|T201|COMP|26882-1|LNC|Homocystine|Homocystine
C0942778|T201|COMP|26700-5|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0942779|T201|COMP|26884-7|LNC|Ketones^3H post XXX challenge|Ketones^3H post XXX challenge
C0942780|T201|COMP|26885-4|LNC|Ova & parasites identified|Ova & parasites identified
C0942781|T201|COMP|26886-2|LNC|ALPRAZolam|ALPRAZolam
C0942782|T201|COMP|26887-0|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C0942783|T201|COMP|26888-8|LNC|Sulfate|Sulfate
C0942784|T201|COMP|26889-6|LNC|Sulfate|Sulfate
C0942785|T201|COMP|26890-4|LNC|Canine distemper virus Ab.IgM|Canine distemper virus Ab.IgM
C0942786|T201|COMP|26892-0|LNC|Intrinsic factor blocking Ab.IgG|Intrinsic factor blocking Ab.IgG
C0942787|T201|COMP|26893-8|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0942788|T201|COMP|26894-6|LNC|Glutamine|Glutamine
C0942789|T201|COMP|26896-1|LNC|Taurine|Taurine
C0942790|T201|COMP|26897-9|LNC|Threonine|Threonine
C0942791|T201|COMP|26898-7|LNC|Temazepam|Temazepam
C0942792|T201|COMP|26900-1|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0942793|T201|COMP|26902-7|LNC|Doxycycline|Doxycycline
C0942794|T201|COMP|26903-5|LNC|Canine distemper virus Ab.IgG|Canine distemper virus Ab.IgG
C0942795|T201|COMP|26904-3|LNC|2-Methylcitrate|2-Methylcitrate
C0942796|T201|COMP|26905-0|LNC|PHENobarbital|PHENobarbital
C0942797|T201|COMP|26907-6|LNC|Listeria sp Ab|Listeria sp Ab
C0942798|T201|COMP|26908-4|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C0942799|T201|COMP|26909-2|LNC|Alpha aminoadipate|Alpha aminoadipate
C0942800|T201|COMP|26910-0|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C0942801|T201|COMP|26911-8|LNC|ALPRAZolam|ALPRAZolam
C0942802|T201|COMP|26912-6|LNC|Hydroxytriazolam|Hydroxytriazolam
C0942803|T201|COMP|26913-4|LNC|Triazolam|Triazolam
C0942804|T201|COMP|26915-9|LNC|Pyridoxine|Pyridoxine
C0942805|T201|COMP|26916-7|LNC|Cobalamins|Cobalamins
C0942807|T201|COMP|26919-1|LNC|Alpha aminobutyrate/Creatinine|Alpha aminobutyrate/Creatinine
C0942808|T201|COMP|26920-9|LNC|Amobarbital|Amobarbital
C0942810|T201|COMP|26923-3|LNC|Butabarbital|Butabarbital
C0942811|T201|COMP|26925-8|LNC|Acetophenazine|Acetophenazine
C0942812|T201|COMP|26928-2|LNC|Vasopressin|Vasopressin
C0942813|T201|COMP|26929-0|LNC|Glycine|Glycine
C0942814|T201|COMP|26930-8|LNC|Secobarbital|Secobarbital
C0942815|T201|COMP|26931-6|LNC|Complement C4|Complement C4
C0942816|T201|COMP|26932-4|LNC|Sarcosine|Sarcosine
C0942817|T201|COMP|26933-2|LNC|Oxazepam|Oxazepam
C0942818|T201|COMP|26934-0|LNC|LORazepam|LORazepam
C0942819|T201|COMP|26935-7|LNC|diazePAM|diazePAM
C0942820|T201|COMP|26936-5|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C0942821|T201|COMP|26937-3|LNC|Temazepam|Temazepam
C0942822|T201|COMP|26938-1|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0942823|T201|COMP|26940-7|LNC|Myelin basic protein|Myelin basic protein
C0942824|T201|COMP|26701-3|LNC|Streptococcus pneumoniae 9 Ab|Streptococcus pneumoniae 9 Ab
C0942825|T201|COMP|26942-3|LNC|Mumps virus Ab|Mumps virus Ab
C0942826|T201|COMP|26944-9|LNC|11-Ketoandrosterone|11-Ketoandrosterone
C0942827|T201|COMP|26945-6|LNC|Triazolam|Triazolam
C0942828|T201|COMP|26946-4|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C0942829|T201|COMP|26947-2|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C0942830|T201|COMP|26948-0|LNC|Saccharopolyspora rectivirgula Ab.IgG|Saccharopolyspora rectivirgula Ab.IgG
C0942831|T201|COMP|26949-8|LNC|Thermoactinomyces sp Ab.IgG|Thermoactinomyces sp Ab.IgG
C0942832|T201|COMP|26950-6|LNC|11-Hydroxyetiocholanolone|11-Hydroxyetiocholanolone
C0942833|T201|COMP|26951-4|LNC|Alternaria alternata Ab.IgG|Alternaria alternata Ab.IgG
C0942834|T201|COMP|26952-2|LNC|Phoma herbarum Ab.IgG|Phoma herbarum Ab.IgG
C0942835|T201|COMP|26953-0|LNC|Dichlorodiphenyltrichloroethane|Dichlorodiphenyltrichloroethane
C0942836|T201|COMP|26954-8|LNC|Aspergillus fumigatus Ab.IgG|Aspergillus fumigatus Ab.IgG
C0942837|T201|COMP|26955-5|LNC|Aureobasidium pullulans Ab.IgG|Aureobasidium pullulans Ab.IgG
C0942838|T201|COMP|26956-3|LNC|Cocaine|Cocaine
C0942839|T201|COMP|26957-1|LNC|Penicillium notatum Ab.IgG|Penicillium notatum Ab.IgG
C0942840|T201|COMP|26958-9|LNC|IgM|IgM
C0942841|T201|COMP|26959-7|LNC|Amphetamine|Amphetamine
C0942842|T201|COMP|26960-5|LNC|Trypsin|Trypsin
C0942843|T201|COMP|26961-3|LNC|Valine|Valine
C0942844|T201|COMP|26962-1|LNC|Cystine|Cystine
C0942845|T201|COMP|26963-9|LNC|Methionine|Methionine
C0942846|T201|COMP|26965-4|LNC|Isoleucine|Isoleucine
C0942847|T201|COMP|26966-2|LNC|Tyrosine|Tyrosine
C0942848|T201|COMP|26967-0|LNC|Phenylalanine|Phenylalanine
C0942849|T201|COMP|26969-6|LNC|Parietal cell Ab|Parietal cell Ab
C0942850|T201|COMP|26970-4|LNC|Reticulin Ab.IgG|Reticulin Ab.IgG
C0942851|T201|COMP|26972-0|LNC|Herpes virus 7 Ab.IgG|Herpes virus 7 Ab.IgG
C0942852|T201|COMP|26975-3|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C0942853|T201|COMP|26977-9|LNC|Coproporphyrin 1|Coproporphyrin 1
C0942854|T201|COMP|26978-7|LNC|Protriptyline|Protriptyline
C0942855|T201|COMP|26979-5|LNC|Flurazepam|Flurazepam
C0942856|T201|COMP|26981-1|LNC|Phenylalanine|Phenylalanine
C0942857|T201|COMP|26982-9|LNC|Cells.CD4+CD25+|Cells.CD4+CD25+
C0942858|T201|COMP|26983-7|LNC|Cells.CD4+HLA-DR+|Cells.CD4+HLA-DR+
C0942859|T201|COMP|26984-5|LNC|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C0942860|T201|COMP|26986-0|LNC|Trichoderma viride Ab.IgG|Trichoderma viride Ab.IgG
C0942861|T201|COMP|26987-8|LNC|Pentachlorophenol/Creatinine|Pentachlorophenol/Creatinine
C0942862|T201|COMP|26988-6|LNC|18-Hydroxydeoxycorticosterone|18-Hydroxydeoxycorticosterone
C0942863|T201|COMP|26990-2|LNC|Phentermine|Phentermine
C0942864|T201|COMP|26991-0|LNC|Phenylpropanolamine|Phenylpropanolamine
C0942865|T201|COMP|26992-8|LNC|Mephentermine|Mephentermine
C0942866|T201|COMP|26994-4|LNC|Phencyclidine|Phencyclidine
C0942867|T201|COMP|26995-1|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0942868|T201|COMP|26996-9|LNC|Complement C7|Complement C7
C0942869|T201|COMP|26997-7|LNC|Cells.CD3+CD25+|Cells.CD3+CD25+
C0942870|T201|COMP|26998-5|LNC|Thyrotropin|Thyrotropin
C0942871|T201|COMP|26999-3|LNC|Homocystine|Homocystine
C0942872|T201|COMP|27000-9|LNC|Thyroxine|Thyroxine
C0942873|T201|COMP|27001-7|LNC|Diethyl ether|Diethyl ether
C0942874|T201|COMP|27002-5|LNC|Secobarbital|Secobarbital
C0942875|T201|COMP|27003-3|LNC|Mephobarbital|Mephobarbital
C0942876|T201|COMP|27005-8|LNC|Xylose^9th specimen post XXX challenge|Xylose^9th specimen post XXX challenge
C0942877|T201|COMP|27006-6|LNC|Xylose^8th specimen post XXX challenge|Xylose^8th specimen post XXX challenge
C0942878|T201|COMP|27007-4|LNC|acetoHEXAMIDE|acetoHEXAMIDE
C0942879|T201|COMP|27008-2|LNC|Xylose^6th specimen post XXX challenge|Xylose^6th specimen post XXX challenge
C0942880|T201|COMP|27009-0|LNC|Coccidioides sp Ab.IgG|Coccidioides sp Ab.IgG
C0942881|T201|COMP|27010-8|LNC|Mesoporphyrin|Mesoporphyrin
C0942882|T201|COMP|27011-6|LNC|Cells.CD14|Cells.CD14
C0942883|T201|COMP|27012-4|LNC|Benzaldehyde|Benzaldehyde
C0942884|T201|COMP|27013-2|LNC|Alanine|Alanine
C0942885|T201|COMP|27014-0|LNC|Inhibin A|Inhibin A
C0942886|T201|COMP|27015-7|LNC|Polychlorinated biphenyl|Polychlorinated biphenyl
C0942887|T201|COMP|27016-5|LNC|Xylose^7th specimen post XXX challenge|Xylose^7th specimen post XXX challenge
C0942888|T201|COMP|27018-1|LNC|IgG.monoclonal|IgG.monoclonal
C0942889|T201|COMP|27019-9|LNC|IgA.monoclonal|IgA.monoclonal
C0942890|T201|COMP|27020-7|LNC|IgM.monoclonal|IgM.monoclonal
C0942891|T201|COMP|27021-5|LNC|Neisseria gonorrhoeae Ab|Neisseria gonorrhoeae Ab
C0942892|T201|COMP|27023-1|LNC|Cells.CD8+CD11b+|Cells.CD8+CD11b+
C0942893|T201|COMP|27025-6|LNC|glipiZIDE|glipiZIDE
C0942894|T201|COMP|27026-4|LNC|Benzoylecgonine|Benzoylecgonine
C0942895|T201|COMP|27027-2|LNC|Cystine|Cystine
C0942896|T201|COMP|27029-8|LNC|Norpropoxyphene|Norpropoxyphene
C0942897|T201|COMP|27030-6|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C0942898|T201|COMP|27031-4|LNC|Oxyphenisatin|Oxyphenisatin
C0942899|T201|COMP|27032-2|LNC|Zirconium|Zirconium
C0942900|T201|COMP|27034-8|LNC|Drugs identified|Drugs identified
C0942901|T201|COMP|27035-5|LNC|Dihydrocodeine+Hydrocodeinone|Dihydrocodeine+Hydrocodeinone
C0942902|T201|COMP|27036-3|LNC|Norchlordiazepoxide|Norchlordiazepoxide
C0942903|T201|COMP|27038-9|LNC|Endomysium Ab.IgA|Endomysium Ab.IgA
C0942904|T201|COMP|27039-7|LNC|Ammonia|Ammonia
C0942905|T201|COMP|27040-5|LNC|Ketones^1H post XXX challenge|Ketones^1H post XXX challenge
C0942906|T201|COMP|27042-1|LNC|Methohexital|Methohexital
C0942907|T201|COMP|27043-9|LNC|Glutamine|Glutamine
C0942908|T201|COMP|27044-7|LNC|1-Methylhistidine|1-Methylhistidine
C0942909|T201|COMP|27046-2|LNC|3-Methylhistidine|3-Methylhistidine
C0942910|T201|COMP|27047-0|LNC|Anserine|Anserine
C0942912|T201|COMP|27049-6|LNC|Secobarbital|Secobarbital
C0942913|T201|COMP|27050-4|LNC|Mephobarbital|Mephobarbital
C0942914|T201|COMP|27052-0|LNC|Methadone|Methadone
C0942915|T201|COMP|27054-6|LNC|Morphine.free|Morphine.free
C0942916|T201|COMP|27055-3|LNC|Catecholamines.free|Catecholamines.free
C0942917|T201|COMP|27056-1|LNC|Citrulline|Citrulline
C0942918|T201|COMP|27058-7|LNC|Beta alanine|Beta alanine
C0942919|T201|COMP|27059-5|LNC|traZODone|traZODone
C0942920|T201|COMP|27060-3|LNC|Melatonin|Melatonin
C0942921|T201|COMP|27061-1|LNC|Butabarbital|Butabarbital
C0942922|T201|COMP|27062-9|LNC|Ketones^1H post XXX challenge|Ketones^1H post XXX challenge
C0942923|T201|COMP|27063-7|LNC|Benzodiazepines|Benzodiazepines
C0942924|T201|COMP|27064-5|LNC|Opiates|Opiates
C0942925|T201|COMP|27065-2|LNC|Ketones^2H post XXX challenge|Ketones^2H post XXX challenge
C0942926|T201|COMP|27066-0|LNC|Ketones^3H post XXX challenge|Ketones^3H post XXX challenge
C0942927|T201|COMP|27067-8|LNC|Propoxyphene|Propoxyphene
C0942928|T201|COMP|27068-6|LNC|Purkinje cells Ab|Purkinje cells Ab
C0942929|T201|COMP|27069-4|LNC|Cisapride|Cisapride
C0942930|T201|COMP|27070-2|LNC|Loratadine|Loratadine
C0942931|T201|COMP|27071-0|LNC|Cells.CD45|Cells.CD45
C0942932|T201|COMP|27072-8|LNC|14-3-3 Ag|14-3-3 Ag
C0942934|T201|COMP|27075-1|LNC|Lycopene|Lycopene
C0942935|T201|COMP|27076-9|LNC|Dextromethorphan+Levorphanol|Dextromethorphan+Levorphanol
C0942936|T201|COMP|27077-7|LNC|Enterococcus sp Ab.IgM|Enterococcus sp Ab.IgM
C0942937|T201|COMP|27078-5|LNC|Carotene.alpha|Carotene.alpha
C0942938|T201|COMP|27079-3|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C0942939|T201|COMP|27080-1|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C0942940|T201|COMP|27081-9|LNC|Itraconazole+Hydroxyitraconazole|Itraconazole+Hydroxyitraconazole
C0942941|T201|COMP|27082-7|LNC|Delavirdine|Delavirdine
C0942942|T201|COMP|27083-5|LNC|Norflunitrazepam|Norflunitrazepam
C0942943|T201|COMP|27084-3|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C0942944|T201|COMP|27085-0|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C0942945|T201|COMP|27086-8|LNC|Cannabinoids|Cannabinoids
C0942946|T201|COMP|27087-6|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C0942947|T201|COMP|27088-4|LNC|Folate|Folate
C0942948|T201|COMP|27089-2|LNC|Asparagine|Asparagine
C0942949|T201|COMP|27090-0|LNC|Entamoeba histolytica Ab.IgA|Entamoeba histolytica Ab.IgA
C0942950|T201|COMP|27091-8|LNC|Calcium|Calcium
C0942951|T201|COMP|27092-6|LNC|Streptococcus pneumoniae 1 Ab.IgG|Streptococcus pneumoniae 1 Ab.IgG
C0942952|T201|COMP|27094-2|LNC|Streptococcus pneumoniae 4 Ab.IgG|Streptococcus pneumoniae 4 Ab.IgG
C0942953|T201|COMP|27095-9|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0942954|T201|COMP|27096-7|LNC|Streptococcus pneumoniae 3 Ab.IgG|Streptococcus pneumoniae 3 Ab.IgG
C0942955|T201|COMP|27099-1|LNC|Riboflavin|Riboflavin
C0942956|T201|COMP|27100-7|LNC|Probenecid|Probenecid
C0942957|T201|COMP|27102-3|LNC|Phendimetrazine|Phendimetrazine
C0942958|T201|COMP|27103-1|LNC|Procyclidine|Procyclidine
C0942959|T201|COMP|27104-9|LNC|Glutamate|Glutamate
C0942960|T201|COMP|27106-4|LNC|Zinc|Zinc
C0942961|T201|COMP|27108-0|LNC|Oleate|Oleate
C0942962|T201|COMP|27109-8|LNC|PARoxetine|PARoxetine
C0942963|T201|COMP|27110-6|LNC|Androsterone|Androsterone
C0942964|T201|COMP|27111-4|LNC|Histidine|Histidine
C0942966|T201|COMP|27114-8|LNC|Cocaine|Cocaine
C0942967|T201|COMP|27115-5|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0942968|T201|COMP|27116-3|LNC|Methamphetamine|Methamphetamine
C0942969|T201|COMP|27117-1|LNC|Cadmium|Cadmium
C0942970|T201|COMP|27119-7|LNC|Streptococcus pneumoniae 23 Ab^2nd specimen|Streptococcus pneumoniae 23 Ab^2nd specimen
C0942973|T201|COMP|27122-1|LNC|Magnesium|Magnesium
C0942974|T201|COMP|27124-7|LNC|Copper|Copper
C0942975|T201|COMP|27125-4|LNC|Zinc|Zinc
C0942976|T201|COMP|27126-2|LNC|Streptococcus pneumoniae 14 Ab^2nd specimen|Streptococcus pneumoniae 14 Ab^2nd specimen
C0942977|T201|COMP|27127-0|LNC|Arsenic|Arsenic
C0942978|T201|COMP|27128-8|LNC|Streptococcus pneumoniae 12 Ab^2nd specimen|Streptococcus pneumoniae 12 Ab^2nd specimen
C0942979|T201|COMP|27129-6|LNC|Lead|Lead
C0942980|T201|COMP|27130-4|LNC|Mercury|Mercury
C0942981|T201|COMP|27131-2|LNC|Phencyclidine|Phencyclidine
C0942982|T201|COMP|27133-8|LNC|Citrate|Citrate
C0942983|T201|COMP|27135-3|LNC|Tryptophan|Tryptophan
C0942984|T201|COMP|27136-1|LNC|Opiates|Opiates
C0942985|T201|COMP|27137-9|LNC|Antimony|Antimony
C0942986|T201|COMP|27138-7|LNC|Streptococcus pneumoniae 23 Ab^1st specimen|Streptococcus pneumoniae 23 Ab^1st specimen
C0942987|T201|COMP|27139-5|LNC|Streptococcus pneumoniae 7f Ab.IgG|Streptococcus pneumoniae 7f Ab.IgG
C0942988|T201|COMP|27140-3|LNC|Follitropin.alpha subunit|Follitropin.alpha subunit
C0942989|T201|COMP|27141-1|LNC|Streptococcus pneumoniae 1 Ab^1st specimen|Streptococcus pneumoniae 1 Ab^1st specimen
C0942990|T201|COMP|27142-9|LNC|Streptococcus pneumoniae 3 Ab^1st specimen|Streptococcus pneumoniae 3 Ab^1st specimen
C0942991|T201|COMP|27143-7|LNC|Streptococcus pneumoniae 4 Ab^1st specimen|Streptococcus pneumoniae 4 Ab^1st specimen
C0942992|T201|COMP|27144-5|LNC|Streptococcus pneumoniae 8 Ab^1st specimen|Streptococcus pneumoniae 8 Ab^1st specimen
C0942993|T201|COMP|27145-2|LNC|Streptococcus pneumoniae 9 Ab^1st specimen|Streptococcus pneumoniae 9 Ab^1st specimen
C0942994|T201|COMP|27146-0|LNC|Streptococcus pneumoniae 12 Ab^1st specimen|Streptococcus pneumoniae 12 Ab^1st specimen
C0942995|T201|COMP|27147-8|LNC|Streptococcus pneumoniae 19 Ab^2nd specimen|Streptococcus pneumoniae 19 Ab^2nd specimen
C0942996|T201|COMP|27148-6|LNC|Streptococcus pneumoniae 19 Ab^1st specimen|Streptococcus pneumoniae 19 Ab^1st specimen
C0942997|T201|COMP|27149-4|LNC|Thiamine|Thiamine
C0943000|T201|COMP|27152-8|LNC|Streptococcus pneumoniae 1 Ab^2nd specimen|Streptococcus pneumoniae 1 Ab^2nd specimen
C0943001|T201|COMP|27153-6|LNC|Streptococcus pneumoniae 3 Ab^2nd specimen|Streptococcus pneumoniae 3 Ab^2nd specimen
C0943002|T201|COMP|27154-4|LNC|Streptococcus pneumoniae 4 Ab^2nd specimen|Streptococcus pneumoniae 4 Ab^2nd specimen
C0943003|T201|COMP|27156-9|LNC|Streptococcus pneumoniae 8 Ab^2nd specimen|Streptococcus pneumoniae 8 Ab^2nd specimen
C0943004|T201|COMP|27157-7|LNC|Streptococcus pneumoniae 9 Ab^2nd specimen|Streptococcus pneumoniae 9 Ab^2nd specimen
C0943005|T201|COMP|27159-3|LNC|Herpes virus 6 Ab.IgM|Herpes virus 6 Ab.IgM
C0943006|T201|COMP|27161-9|LNC|Interleukin 4|Interleukin 4
C0943007|T201|COMP|27162-7|LNC|1-Methylhistidine|1-Methylhistidine
C0943008|T201|COMP|27163-5|LNC|N-methylacetamide/Creatinine|N-methylacetamide/Creatinine
C0943009|T201|COMP|27166-8|LNC|TOLAZamide|TOLAZamide
C0943010|T201|COMP|27167-6|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C0943011|T201|COMP|27168-4|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C0943012|T201|COMP|27170-0|LNC|TOLBUTamide|TOLBUTamide
C0943013|T201|COMP|27171-8|LNC|Chlorphentermine|Chlorphentermine
C0943014|T201|COMP|27173-4|LNC|Propylthiouracil|Propylthiouracil
C0943015|T201|COMP|27174-2|LNC|Inhibin|Inhibin
C0943016|T201|COMP|27175-9|LNC|glyBURIDE|glyBURIDE
C0943017|T201|COMP|27176-7|LNC|3-Methylhistidine|3-Methylhistidine
C0943018|T201|COMP|27178-3|LNC|Phendimetrazine|Phendimetrazine
C0943019|T201|COMP|27179-1|LNC|Threonine|Threonine
C0943020|T201|COMP|27181-7|LNC|Hydroxyproline|Hydroxyproline
C0943021|T201|COMP|27182-5|LNC|Calcium|Calcium
C0943022|T201|COMP|27183-3|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C0943023|T201|COMP|27184-1|LNC|Alpha 1 globulin|Alpha 1 globulin
C0943024|T201|COMP|27186-6|LNC|Lysozyme|Lysozyme
C0943025|T201|COMP|27187-4|LNC|Methohexital|Methohexital
C0943026|T201|COMP|27188-2|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0943027|T201|COMP|27189-0|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0943028|T201|COMP|27191-6|LNC|PHENobarbital|PHENobarbital
C0943029|T201|COMP|27192-4|LNC|diazePAM|diazePAM
C0943030|T201|COMP|27193-2|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C0943031|T201|COMP|27194-0|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0943032|T201|COMP|27195-7|LNC|Hydroxylysine|Hydroxylysine
C0943033|T201|COMP|27196-5|LNC|HYDROmorphone.free|HYDROmorphone.free
C0943034|T201|COMP|27197-3|LNC|Benzodiazepines|Benzodiazepines
C0943035|T201|COMP|27198-1|LNC|Bilirubin|Bilirubin
C0943036|T201|COMP|27199-9|LNC|18-Hydroxycortisol/Creatinine|18-Hydroxycortisol/Creatinine
C0943037|T201|COMP|27200-5|LNC|Nuclear Ab|Nuclear Ab
C0943038|T201|COMP|27201-3|LNC|Zinc/Creatinine|Zinc/Creatinine
C0943039|T201|COMP|27202-1|LNC|Halothane|Halothane
C0943040|T201|COMP|27203-9|LNC|Follitropin|Follitropin
C0943041|T201|COMP|27204-7|LNC|Cocaine|Cocaine
C0943042|T201|COMP|27205-4|LNC|Amphetamines|Amphetamines
C0943043|T201|COMP|27206-2|LNC|Morphine.free|Morphine.free
C0943044|T201|COMP|27207-0|LNC|Methadone|Methadone
C0943045|T201|COMP|27208-8|LNC|Drugs identified|Drugs identified
C0943046|T201|COMP|27210-4|LNC|Magnesium|Magnesium
C0943047|T201|COMP|27211-2|LNC|Norpropoxyphene|Norpropoxyphene
C0943048|T201|COMP|27212-0|LNC|DOPamine|DOPamine
C0943049|T201|COMP|27213-8|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0943050|T201|COMP|27214-6|LNC|Purkinje cells Ab|Purkinje cells Ab
C0943051|T201|COMP|27216-1|LNC|sulfADIAZINE|sulfADIAZINE
C0943052|T201|COMP|27217-9|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0943053|T201|COMP|27218-7|LNC|quiNINE|quiNINE
C0943054|T201|COMP|27219-5|LNC|Ornithine|Ornithine
C0943055|T201|COMP|27220-3|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C0943056|T201|COMP|27222-9|LNC|Oxalate|Oxalate
C0943057|T201|COMP|27223-7|LNC|Serine|Serine
C0943058|T201|COMP|27224-5|LNC|Barbiturates|Barbiturates
C0943059|T201|COMP|27226-0|LNC|Cocaethylene|Cocaethylene
C0943060|T201|COMP|27227-8|LNC|Streptococcus pneumoniae 1 Ab.IgG|Streptococcus pneumoniae 1 Ab.IgG
C0943061|T201|COMP|27228-6|LNC|Streptococcus pneumoniae 3 Ab.IgG|Streptococcus pneumoniae 3 Ab.IgG
C0943062|T201|COMP|27230-2|LNC|Streptococcus pneumoniae 19 Ab.IgG|Streptococcus pneumoniae 19 Ab.IgG
C0943063|T201|COMP|27231-0|LNC|Streptococcus pneumoniae 23 Ab.IgG|Streptococcus pneumoniae 23 Ab.IgG
C0943064|T201|COMP|27232-8|LNC|Lead|Lead
C0943065|T201|COMP|27233-6|LNC|Lecithin|Lecithin
C0943066|T201|COMP|27235-1|LNC|PHENobarbital|PHENobarbital
C0943067|T201|COMP|27236-9|LNC|Azatadine|Azatadine
C0943068|T201|COMP|27237-7|LNC|LORazepam|LORazepam
C0943069|T201|COMP|27239-3|LNC|Nordiazepam|Nordiazepam
C0943070|T201|COMP|27240-1|LNC|PHENobarbital|PHENobarbital
C0943071|T201|COMP|27242-7|LNC|Secobarbital|Secobarbital
C0943072|T201|COMP|27243-5|LNC|PENTobarbital|PENTobarbital
C0943073|T201|COMP|27244-3|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0943074|T201|COMP|27245-0|LNC|Amobarbital|Amobarbital
C0943075|T201|COMP|27247-6|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C0943076|T201|COMP|27250-0|LNC|Phenmetrazine|Phenmetrazine
C0943077|T201|COMP|27251-8|LNC|Phenylpropanolamine|Phenylpropanolamine
C0943078|T201|COMP|27252-6|LNC|Choriogonadotropin.alpha subunit|Choriogonadotropin.alpha subunit
C0943079|T201|COMP|27253-4|LNC|Chlorphentermine|Chlorphentermine
C0943080|T201|COMP|27254-2|LNC|Amino beta guanidinopropionate/Creatinine|Amino beta guanidinopropionate/Creatinine
C0943081|T201|COMP|27255-9|LNC|Magnesium|Magnesium
C0943082|T201|COMP|27256-7|LNC|Aspartate|Aspartate
C0943083|T201|COMP|27257-5|LNC|Sodium|Sodium
C0943084|T201|COMP|27258-3|LNC|Protein|Protein
C0943085|T201|COMP|27259-1|LNC|Estriol.unconjugated|Estriol.unconjugated
C0943086|T201|COMP|27260-9|LNC|Schistosoma sp Ab.IgG|Schistosoma sp Ab.IgG
C0943087|T201|COMP|27261-7|LNC|Polio virus Ab|Polio virus Ab
C0943088|T201|COMP|27262-5|LNC|Methaqualone|Methaqualone
C0943089|T201|COMP|27263-3|LNC|Amphetamines|Amphetamines
C0943090|T201|COMP|27265-8|LNC|Giardia sp Ag|Giardia sp Ag
C0943091|T201|COMP|27266-6|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0943092|T201|COMP|27267-4|LNC|Homovanillate|Homovanillate
C0943093|T201|COMP|27268-2|LNC|Hydroxydecanedioate|Hydroxydecanedioate
C0943094|T201|COMP|27269-0|LNC|Isocitrate|Isocitrate
C0943095|T201|COMP|27270-8|LNC|4-Hydroxyphenylacetate|4-Hydroxyphenylacetate
C0943096|T201|COMP|27271-6|LNC|Alpha ketoglutarate|Alpha ketoglutarate
C0943097|T201|COMP|27272-4|LNC|3-Hydroxyisobutyrate|3-Hydroxyisobutyrate
C0943098|T201|COMP|27273-2|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C0943099|T201|COMP|27004-1|LNC|Benzfetamine|Benzfetamine
C0943100|T201|COMP|27275-7|LNC|diazePAM|diazePAM
C0943101|T201|COMP|27276-5|LNC|Azatadine|Azatadine
C0943102|T201|COMP|27277-3|LNC|Methamphetamine|Methamphetamine
C0943103|T201|COMP|27278-1|LNC|Phosphoethanolamine|Phosphoethanolamine
C0943104|T201|COMP|27279-9|LNC|Paraoxon|Paraoxon
C0943105|T201|COMP|27280-7|LNC|Tripelennamine|Tripelennamine
C0943106|T201|COMP|27281-5|LNC|Propoxyphene|Propoxyphene
C0943107|T201|COMP|27282-3|LNC|Carbinoxamine|Carbinoxamine
C0943108|T201|COMP|27283-1|LNC|Methadone|Methadone
C0943109|T201|COMP|27284-9|LNC|Brompheniramine|Brompheniramine
C0943110|T201|COMP|27286-4|LNC|Triazolam|Triazolam
C0943111|T201|COMP|27287-2|LNC|Flurazepam|Flurazepam
C0943112|T201|COMP|27288-0|LNC|Midazolam|Midazolam
C0943113|T201|COMP|27290-6|LNC|Phenmetrazine|Phenmetrazine
C0943114|T201|COMP|27291-4|LNC|Hydroxylysine|Hydroxylysine
C0943115|T201|COMP|27294-8|LNC|Carnosine|Carnosine
C0943116|T201|COMP|27295-5|LNC|Cocaethylene|Cocaethylene
C0943117|T201|COMP|27296-3|LNC|Arginine|Arginine
C0943118|T201|COMP|27298-9|LNC|Protein|Protein
C0943119|T201|COMP|27301-1|LNC|Glutarate|Glutarate
C0943120|T201|COMP|27302-9|LNC|Midazolam|Midazolam
C0943121|T201|COMP|27303-7|LNC|Phendimetrazine|Phendimetrazine
C0943122|T201|COMP|27305-2|LNC|Phentermine|Phentermine
C0943123|T201|COMP|27306-0|LNC|Testosterone|Testosterone
C0943124|T201|COMP|27307-8|LNC|Chlorphentermine|Chlorphentermine
C0943125|T201|COMP|27309-4|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C0943126|T201|COMP|27310-2|LNC|Taurine|Taurine
C0943127|T201|COMP|27311-0|LNC|Codeine.free|Codeine.free
C0943128|T201|COMP|27313-6|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C0943129|T201|COMP|27314-4|LNC|HYDROmorphone.free|HYDROmorphone.free
C0943130|T201|COMP|27315-1|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0943131|T201|COMP|27316-9|LNC|Dioxin|Dioxin
C0943132|T201|COMP|27318-5|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C0943133|T201|COMP|27319-3|LNC|Reducing substances|Reducing substances
C0943134|T201|COMP|27321-9|LNC|Opiates|Opiates
C0943135|T201|COMP|27322-7|LNC|Threonine|Threonine
C0943136|T201|COMP|27323-5|LNC|Leucine|Leucine
C0943137|T201|COMP|27324-3|LNC|Amobarbital|Amobarbital
C0943138|T201|COMP|27326-8|LNC|Alanine|Alanine
C0943140|T201|COMP|27328-4|LNC|Somatotropin^6th specimen post XXX challenge|Somatotropin^6th specimen post XXX challenge
C0943141|T201|COMP|27329-2|LNC|Feline panleukopenia virus Ab.IgM|Feline panleukopenia virus Ab.IgM
C0943142|T201|COMP|27330-0|LNC|Insulin^1.5H post XXX challenge|Insulin^1.5H post XXX challenge
C0943143|T201|COMP|27331-8|LNC|Imipenem|Imipenem
C0943144|T201|COMP|27332-6|LNC|Feline panleukopenia virus Ab.IgG|Feline panleukopenia virus Ab.IgG
C0943145|T201|COMP|27333-4|LNC|Lysine|Lysine
C0943146|T201|COMP|27334-2|LNC|Tryptophan|Tryptophan
C0943147|T201|COMP|27335-9|LNC|Ornithine|Ornithine
C0943148|T201|COMP|27336-7|LNC|Amino acids|Amino acids
C0943149|T201|COMP|27337-5|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0943150|T201|COMP|27338-3|LNC|2,4-Dichlorophenoxyacetate|2,4-Dichlorophenoxyacetate
C0943151|T201|COMP|27339-1|LNC|Nicotinamide|Nicotinamide
C0943152|T201|COMP|27340-9|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C0943153|T201|COMP|27341-7|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0943154|T201|COMP|27342-5|LNC|Fasciola hepatica Ab|Fasciola hepatica Ab
C0943155|T201|COMP|27343-3|LNC|Molybdenum|Molybdenum
C0943156|T201|COMP|27344-1|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C0943157|T201|COMP|27345-8|LNC|Hemoglobin A2|Hemoglobin A2
C0943158|T201|COMP|27346-6|LNC|Benzfetamine|Benzfetamine
C0943159|T201|COMP|27347-4|LNC|Methaqualone|Methaqualone
C0943160|T201|COMP|27348-2|LNC|DOPamine^2H post XXX challenge|DOPamine^2H post XXX challenge
C0943161|T201|COMP|27349-0|LNC|Cystathionine|Cystathionine
C0943162|T201|COMP|27350-8|LNC|Cystine|Cystine
C0943163|T201|COMP|27351-6|LNC|Pantothenate|Pantothenate
C0943164|T201|COMP|27352-4|LNC|Homocystine|Homocystine
C0943165|T201|COMP|27353-2|LNC|Estimated average glucose|Estimated average glucose
C0943166|T201|COMP|27356-5|LNC|Phencyclidine|Phencyclidine
C0943167|T201|COMP|27357-3|LNC|HYDROcodone.free|HYDROcodone.free
C0943168|T201|COMP|27358-1|LNC|Benzoylecgonine|Benzoylecgonine
C0943169|T201|COMP|27360-7|LNC|Myelin basic protein Ab|Myelin basic protein Ab
C0943170|T201|COMP|27361-5|LNC|Tyrosine|Tyrosine
C0943171|T201|COMP|27362-3|LNC|Phenylalanine|Phenylalanine
C0943172|T201|COMP|27363-1|LNC|DOPamine^3H post XXX challenge|DOPamine^3H post XXX challenge
C0943173|T201|COMP|27365-6|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C0943174|T201|COMP|27366-4|LNC|Somatotropin^22nd specimen post XXX challenge|Somatotropin^22nd specimen post XXX challenge
C0943175|T201|COMP|27367-2|LNC|Manganese/Creatinine|Manganese/Creatinine
C0943176|T201|COMP|27368-0|LNC|Chlamydia trachomatis B Ab|Chlamydia trachomatis B Ab
C0943177|T201|COMP|27370-6|LNC|Chlamydia trachomatis C Ab|Chlamydia trachomatis C Ab
C0943178|T201|COMP|27371-4|LNC|Chlamydia trachomatis G+F+K Ab|Chlamydia trachomatis G+F+K Ab
C0943179|T201|COMP|27372-2|LNC|Insulin^20M post XXX challenge|Insulin^20M post XXX challenge
C0943180|T201|COMP|27374-8|LNC|Streptococcus pneumoniae 12 Ab.IgG|Streptococcus pneumoniae 12 Ab.IgG
C0943181|T201|COMP|27375-5|LNC|Aspergillus fumigatus Ab|Aspergillus fumigatus Ab
C0943182|T201|COMP|27377-1|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C0943183|T201|COMP|27379-7|LNC|Insulin^1H post XXX challenge|Insulin^1H post XXX challenge
C0943184|T201|COMP|27380-5|LNC|DOPamine^4H post XXX challenge|DOPamine^4H post XXX challenge
C0943185|T201|COMP|27383-9|LNC|Feline herpesvirus 1 Ab|Feline herpesvirus 1 Ab
C0943186|T201|COMP|27384-7|LNC|Leptospira sp Ab.IgM|Leptospira sp Ab.IgM
C0943187|T201|COMP|27386-2|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0943188|T201|COMP|27387-0|LNC|Streptococcus pneumoniae 14 Ab.IgG|Streptococcus pneumoniae 14 Ab.IgG
C0943190|T201|COMP|27389-6|LNC|Streptococcus pneumoniae 23 Ab.IgG|Streptococcus pneumoniae 23 Ab.IgG
C0943191|T201|COMP|27390-4|LNC|Streptococcus pneumoniae 19 Ab.IgG|Streptococcus pneumoniae 19 Ab.IgG
C0943192|T201|COMP|27391-2|LNC|Candida sp Ab.IgM|Candida sp Ab.IgM
C0943193|T201|COMP|27392-0|LNC|Streptococcus pneumoniae 9 Ab.IgG|Streptococcus pneumoniae 9 Ab.IgG
C0943194|T201|COMP|27393-8|LNC|Streptococcus pneumoniae 23f Ab.IgG|Streptococcus pneumoniae 23f Ab.IgG
C0943195|T201|COMP|27394-6|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C0943197|T201|COMP|27396-1|LNC|Hemoglobin.gastrointestinal|Hemoglobin.gastrointestinal
C0943198|T201|COMP|27397-9|LNC|Streptococcus pneumoniae 12f Ab.IgG|Streptococcus pneumoniae 12f Ab.IgG
C0943199|T201|COMP|27398-7|LNC|Streptococcus pneumoniae 9n Ab.IgG|Streptococcus pneumoniae 9n Ab.IgG
C0943200|T201|COMP|27399-5|LNC|1-Methylhistidine|1-Methylhistidine
C0943201|T201|COMP|27400-1|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C0943202|T201|COMP|27401-9|LNC|Hemoglobin.gastrointestinal^6th specimen|Hemoglobin.gastrointestinal^6th specimen
C0943203|T201|COMP|27402-7|LNC|Norparamethadione|Norparamethadione
C0943204|T201|COMP|27404-3|LNC|Chlamydophila psittaci Ab.IgM|Chlamydophila psittaci Ab.IgM
C0943206|T201|COMP|27406-8|LNC|Streptococcus pneumoniae 19f Ab.IgG|Streptococcus pneumoniae 19f Ab.IgG
C0943207|T201|COMP|27407-6|LNC|Streptococcus pneumoniae 14 Ab.IgG^1st specimen|Streptococcus pneumoniae 14 Ab.IgG^1st specimen
C0943208|T201|COMP|27408-4|LNC|C peptide^20M post XXX challenge|C peptide^20M post XXX challenge
C0943209|T201|COMP|27409-2|LNC|Methylenedianiline|Methylenedianiline
C0943211|T201|COMP|27411-8|LNC|Iron/Creatinine|Iron/Creatinine
C0943212|T201|COMP|27413-4|LNC|Dextromethorphan|Dextromethorphan
C0943213|T201|COMP|27414-2|LNC|Fungus identified|Fungus identified
C0943214|T201|COMP|27415-9|LNC|Interferon.gamma|Interferon.gamma
C0943215|T201|COMP|27416-7|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C0943216|T201|COMP|27417-5|LNC|Candida sp Ab.IgA|Candida sp Ab.IgA
C0943217|T201|COMP|27418-3|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0943218|T201|COMP|27420-9|LNC|Phosphatidylglycerol|Phosphatidylglycerol
C0943219|T201|COMP|27421-7|LNC|C peptide^40M post XXX challenge|C peptide^40M post XXX challenge
C0943220|T201|COMP|27422-5|LNC|Streptococcus pneumoniae 3 Ab.IgG^2nd specimen|Streptococcus pneumoniae 3 Ab.IgG^2nd specimen
C0943221|T201|COMP|27424-1|LNC|Deoxypyridinoline|Deoxypyridinoline
C0943222|T201|COMP|27425-8|LNC|Streptococcus pneumoniae 14 Ab.IgG^2nd specimen|Streptococcus pneumoniae 14 Ab.IgG^2nd specimen
C0943223|T201|COMP|27426-6|LNC|Trichinella sp Ab.IgM|Trichinella sp Ab.IgM
C0943224|T201|COMP|27428-2|LNC|Streptococcus pneumoniae 1 Ab.IgG^1st specimen|Streptococcus pneumoniae 1 Ab.IgG^1st specimen
C0943225|T201|COMP|27429-0|LNC|Streptococcus pneumoniae 19 Ab.IgG^2nd specimen|Streptococcus pneumoniae 19 Ab.IgG^2nd specimen
C0943226|T201|COMP|27430-8|LNC|Streptococcus pneumoniae 3 Ab.IgG^1st specimen|Streptococcus pneumoniae 3 Ab.IgG^1st specimen
C0943227|T201|COMP|27431-6|LNC|Streptococcus pneumoniae 1 Ab.IgG^2nd specimen|Streptococcus pneumoniae 1 Ab.IgG^2nd specimen
C0943229|T201|COMP|27434-0|LNC|Streptococcus pneumoniae 23 Ab.IgG^1st specimen|Streptococcus pneumoniae 23 Ab.IgG^1st specimen
C0943230|T201|COMP|27436-5|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C0943231|T201|COMP|27437-3|LNC|Streptococcus pneumoniae 23 Ab.IgG^2nd specimen|Streptococcus pneumoniae 23 Ab.IgG^2nd specimen
C0943232|T201|COMP|27439-9|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C0943233|T201|COMP|27440-7|LNC|Candida sp Ag|Candida sp Ag
C0943234|T201|COMP|27441-5|LNC|Potassium|Potassium
C0943235|T201|COMP|27443-1|LNC|DOPamine^1H post XXX challenge|DOPamine^1H post XXX challenge
C0943236|T201|COMP|27444-9|LNC|Insulin^40M post XXX challenge|Insulin^40M post XXX challenge
C0943506|T201|COMP|27811-9|LNC|Antithrombin actual/Normal|Antithrombin actual/Normal
C0943507|T201|COMP|27812-7|LNC|Antithrombin Ag actual/Normal|Antithrombin Ag actual/Normal
C0943508|T201|COMP|27813-5|LNC|Prothrombin Ag actual/Normal|Prothrombin Ag actual/Normal
C0943510|T201|COMP|27815-0|LNC|Coagulation factor XIII activity actual/Normal|Coagulation factor XIII activity actual/Normal
C0943511|T201|COMP|27816-8|LNC|von Willebrand factor Ag actual/Normal|von Willebrand factor Ag actual/Normal
C0943512|T201|COMP|27817-6|LNC|Beta 2 glycoprotein 1 Ab|Beta 2 glycoprotein 1 Ab
C0943513|T201|COMP|27818-4|LNC|Protein C actual/Normal|Protein C actual/Normal
C0943514|T201|COMP|27819-2|LNC|Protein C actual/Normal|Protein C actual/Normal
C0943515|T201|COMP|27820-0|LNC|Protein C Ag actual/Normal|Protein C Ag actual/Normal
C0943516|T201|COMP|27821-8|LNC|Protein S.free Ag actual/Normal|Protein S.free Ag actual/Normal
C0943517|T201|COMP|27823-4|LNC|Protein S Ag actual/Normal|Protein S Ag actual/Normal
C0943518|T201|COMP|27824-2|LNC|Prothrombin fragment 1+2 Ag|Prothrombin fragment 1+2 Ag
C0943519|T201|COMP|27825-9|LNC|Platelet associated Ab|Platelet associated Ab
C0943520|T201|COMP|27826-7|LNC|Insulin^2H post XXX challenge|Insulin^2H post XXX challenge
C0943521|T201|COMP|27828-3|LNC|Insulin^3H post XXX challenge|Insulin^3H post XXX challenge
C0943522|T201|COMP|27830-9|LNC|Insulin^1H post 75 g glucose PO|Insulin^1H post 75 g glucose PO
C0943523|T201|COMP|27832-5|LNC|Insulin^4th specimen post XXX challenge|Insulin^4th specimen post XXX challenge
C0943524|T201|COMP|27833-3|LNC|Insulin^7H post 75 g glucose PO|Insulin^7H post 75 g glucose PO
C0943525|T201|COMP|27834-1|LNC|Insulin^1.5H post 75 g glucose PO|Insulin^1.5H post 75 g glucose PO
C0943526|T201|COMP|27835-8|LNC|Somatotropin^11th specimen post XXX challenge|Somatotropin^11th specimen post XXX challenge
C0943527|T201|COMP|27836-6|LNC|Somatotropin^12th specimen post XXX challenge|Somatotropin^12th specimen post XXX challenge
C0943528|T201|COMP|27838-2|LNC|Somatotropin^14th specimen post XXX challenge|Somatotropin^14th specimen post XXX challenge
C0943529|T201|COMP|27839-0|LNC|C peptide^4H post XXX challenge|C peptide^4H post XXX challenge
C0943530|T201|COMP|27840-8|LNC|Somatotropin^16th specimen post XXX challenge|Somatotropin^16th specimen post XXX challenge
C0943531|T201|COMP|27841-6|LNC|Somatotropin^17th specimen post XXX challenge|Somatotropin^17th specimen post XXX challenge
C0943532|T201|COMP|27842-4|LNC|Somatotropin^19th specimen post XXX challenge|Somatotropin^19th specimen post XXX challenge
C0943533|T201|COMP|27843-2|LNC|Somatotropin^20th specimen post XXX challenge|Somatotropin^20th specimen post XXX challenge
C0943534|T201|COMP|27844-0|LNC|Somatotropin^21st specimen post XXX challenge|Somatotropin^21st specimen post XXX challenge
C0943535|T201|COMP|27845-7|LNC|Somatotropin^23rd specimen post XXX challenge|Somatotropin^23rd specimen post XXX challenge
C0943536|T201|COMP|27846-5|LNC|Somatotropin^24th specimen post XXX challenge|Somatotropin^24th specimen post XXX challenge
C0943537|T201|COMP|27848-1|LNC|Lutropin^2nd specimen post XXX challenge|Lutropin^2nd specimen post XXX challenge
C0943538|T201|COMP|27849-9|LNC|Aldosterone^2nd specimen post XXX challenge|Aldosterone^2nd specimen post XXX challenge
C0943539|T201|COMP|27850-7|LNC|Somatotropin^10M post XXX challenge|Somatotropin^10M post XXX challenge
C0943540|T201|COMP|27851-5|LNC|Lutropin^3rd specimen post XXX challenge|Lutropin^3rd specimen post XXX challenge
C0943541|T201|COMP|27852-3|LNC|Insulin^5H post XXX challenge|Insulin^5H post XXX challenge
C0943542|T201|COMP|27853-1|LNC|Lutropin^4th specimen post XXX challenge|Lutropin^4th specimen post XXX challenge
C0943543|T201|COMP|27854-9|LNC|Lutropin^5th specimen post XXX challenge|Lutropin^5th specimen post XXX challenge
C0943544|T201|COMP|27855-6|LNC|Lutropin^6th specimen post XXX challenge|Lutropin^6th specimen post XXX challenge
C0943545|T201|COMP|27856-4|LNC|Proinsulin^2H post XXX challenge|Proinsulin^2H post XXX challenge
C0943546|T201|COMP|27857-2|LNC|Proinsulin^3H post XXX challenge|Proinsulin^3H post XXX challenge
C0943547|T201|COMP|27858-0|LNC|Lutropin^7th specimen post XXX challenge|Lutropin^7th specimen post XXX challenge
C0943548|T201|COMP|27859-8|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C0943549|T201|COMP|27860-6|LNC|Insulin^2H post 75 g glucose PO|Insulin^2H post 75 g glucose PO
C0943550|T201|COMP|27861-4|LNC|Insulin^3H post 75 g glucose PO|Insulin^3H post 75 g glucose PO
C0943551|T201|COMP|27862-2|LNC|Insulin^4H post 75 g glucose PO|Insulin^4H post 75 g glucose PO
C0943552|T201|COMP|27863-0|LNC|Insulin^2.5H post XXX challenge|Insulin^2.5H post XXX challenge
C0943553|T201|COMP|27865-5|LNC|Follitropin^3rd specimen post XXX challenge|Follitropin^3rd specimen post XXX challenge
C0943554|T201|COMP|27866-3|LNC|17-Ketogenic steroids|17-Ketogenic steroids
C0943555|T201|COMP|27867-1|LNC|Insulin^7th specimen post XXX challenge|Insulin^7th specimen post XXX challenge
C0943556|T201|COMP|27868-9|LNC|Follitropin^5th specimen post XXX challenge|Follitropin^5th specimen post XXX challenge
C0943557|T201|COMP|27869-7|LNC|Follitropin^8th specimen post XXX challenge|Follitropin^8th specimen post XXX challenge
C0943558|T201|COMP|27870-5|LNC|Follitropin^4th specimen post XXX challenge|Follitropin^4th specimen post XXX challenge
C0943559|T201|COMP|27871-3|LNC|Interferon.beta Ab.IgG|Interferon.beta Ab.IgG
C0943560|T201|COMP|27872-1|LNC|Insulin^6H post 75 g glucose PO|Insulin^6H post 75 g glucose PO
C0943561|T201|COMP|27873-9|LNC|Insulin^post CFst|Insulin^post CFst
C0943562|T201|COMP|27874-7|LNC|Insulin^5th specimen post XXX challenge|Insulin^5th specimen post XXX challenge
C0943563|T201|COMP|27876-2|LNC|Cells.CD14+CD11b+/100 cells|Cells.CD14+CD11b+/100 cells
C0943564|T201|COMP|27877-0|LNC|Cells.CD33+CD11b+/100 cells|Cells.CD33+CD11b+/100 cells
C0943565|T201|COMP|27878-8|LNC|Cells.CD14+HLA-DR+/100 cells|Cells.CD14+HLA-DR+/100 cells
C0943566|T201|COMP|27879-6|LNC|Cells.CD33+HLA-DR+/100 cells|Cells.CD33+HLA-DR+/100 cells
C0943567|T201|COMP|27881-2|LNC|Somatotropin^4th specimen post XXX challenge|Somatotropin^4th specimen post XXX challenge
C0943568|T201|COMP|27882-0|LNC|Proinsulin|Proinsulin
C0943569|T201|COMP|27883-8|LNC|Lutropin^15M post XXX challenge|Lutropin^15M post XXX challenge
C0943570|T201|COMP|27886-1|LNC|Follitropin^40M post XXX challenge|Follitropin^40M post XXX challenge
C0943571|T201|COMP|27887-9|LNC|Follitropin^15M post XXX challenge|Follitropin^15M post XXX challenge
C0943572|T201|COMP|27888-7|LNC|Somatotropin^2nd specimen post XXX challenge|Somatotropin^2nd specimen post XXX challenge
C0943573|T201|COMP|27889-5|LNC|Somatotropin^3rd specimen post XXX challenge|Somatotropin^3rd specimen post XXX challenge
C0943574|T201|COMP|27891-1|LNC|Thyroxine^baseline|Thyroxine^baseline
C0943575|T201|COMP|27892-9|LNC|Butyrylglycine/Creatinine|Butyrylglycine/Creatinine
C0943576|T201|COMP|27893-7|LNC|Cells.CD19+CD23+/100 cells|Cells.CD19+CD23+/100 cells
C0943577|T201|COMP|27894-5|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C0943582|T201|COMP|27900-0|LNC|Lactobacillus sp Ab.IgG|Lactobacillus sp Ab.IgG
C0943583|T201|COMP|27901-8|LNC|Lactobacillus sp Ab.IgM|Lactobacillus sp Ab.IgM
C0943584|T201|COMP|27902-6|LNC|Enterococcus sp Ab.IgG|Enterococcus sp Ab.IgG
C0943585|T201|COMP|27903-4|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C0943586|T201|COMP|27904-2|LNC|Histidine|Histidine
C0943587|T201|COMP|27905-9|LNC|Bacteroides fragilis Ab.IgM|Bacteroides fragilis Ab.IgM
C0943588|T201|COMP|27906-7|LNC|Lymphocytes.immature/100 leukocytes|Lymphocytes.immature/100 leukocytes
C0943589|T201|COMP|27907-5|LNC|Cryptosporidium sp|Cryptosporidium sp
C0943590|T201|COMP|27910-9|LNC|Calcium^6th specimen post XXX challenge|Calcium^6th specimen post XXX challenge
C0943591|T201|COMP|27911-7|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0943592|T201|COMP|27912-5|LNC|Butalbital|Butalbital
C0943593|T201|COMP|27913-3|LNC|Calcium^7th specimen post XXX challenge|Calcium^7th specimen post XXX challenge
C0943594|T201|COMP|27914-1|LNC|Gamma aminoadipate|Gamma aminoadipate
C0943595|T201|COMP|27915-8|LNC|Alpha-1-Antichymotrypsin|Alpha-1-Antichymotrypsin
C0943596|T201|COMP|27916-6|LNC|Calcium^2nd specimen post XXX challenge|Calcium^2nd specimen post XXX challenge
C0943597|T201|COMP|27917-4|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C0943598|T201|COMP|27918-2|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C0943599|T201|COMP|27919-0|LNC|Calcium^3rd specimen post XXX challenge|Calcium^3rd specimen post XXX challenge
C0943600|T201|COMP|27920-8|LNC|Normeperidine|Normeperidine
C0943601|T201|COMP|27921-6|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C0943602|T201|COMP|27922-4|LNC|Echovirus 4 RNA|Echovirus 4 RNA
C0943603|T201|COMP|27923-2|LNC|Ubiquinone 10|Ubiquinone 10
C0943604|T201|COMP|27924-0|LNC|Ascaris sp Ab|Ascaris sp Ab
C0943605|T201|COMP|27925-7|LNC|Hemoglobin.gastrointestinal^7th specimen|Hemoglobin.gastrointestinal^7th specimen
C0943606|T201|COMP|27926-5|LNC|Hemoglobin.gastrointestinal^8th specimen|Hemoglobin.gastrointestinal^8th specimen
C0943607|T201|COMP|27927-3|LNC|Butalbital|Butalbital
C0943608|T201|COMP|27928-1|LNC|Echovirus 30 RNA|Echovirus 30 RNA
C0943609|T201|COMP|27929-9|LNC|Mandelate|Mandelate
C0943610|T201|COMP|27931-5|LNC|Bile acid^2H post meal|Bile acid^2H post meal
C0943611|T201|COMP|27932-3|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0943612|T201|COMP|27933-1|LNC|Calcium^5th specimen post XXX challenge|Calcium^5th specimen post XXX challenge
C0943613|T201|COMP|27934-9|LNC|Echovirus 11 RNA|Echovirus 11 RNA
C0943614|T201|COMP|27936-4|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0943615|T201|COMP|27938-0|LNC|Salmonella paratyphi B O Ab|Salmonella paratyphi B O Ab
C0943616|T201|COMP|27939-8|LNC|Collagen crosslinked N-telopeptide|Collagen crosslinked N-telopeptide
C0943617|T201|COMP|27941-4|LNC|Lactate|Lactate
C0943618|T201|COMP|27942-2|LNC|Follitropin|Follitropin
C0943619|T201|COMP|27943-0|LNC|Interferon.omega|Interferon.omega
C0943620|T201|COMP|27944-8|LNC|C peptide|C peptide
C0943621|T201|COMP|27947-1|LNC|Coxsackievirus A7 RNA|Coxsackievirus A7 RNA
C0943622|T201|COMP|27948-9|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C0943623|T201|COMP|27949-7|LNC|Lactate^4H post XXX challenge|Lactate^4H post XXX challenge
C0943624|T201|COMP|27950-5|LNC|Saint Louis encephalitis virus RNA|Saint Louis encephalitis virus RNA
C0943625|T201|COMP|27951-3|LNC|Coxiella burnetii phase 1 Ab|Coxiella burnetii phase 1 Ab
C0943626|T201|COMP|27952-1|LNC|Enterovirus RNA|Enterovirus RNA
C0943627|T201|COMP|27953-9|LNC|Methionine|Methionine
C0943628|T201|COMP|27955-4|LNC|Lactate^2H post XXX challenge|Lactate^2H post XXX challenge
C0943629|T201|COMP|27956-2|LNC|Proinsulin^1H post XXX challenge|Proinsulin^1H post XXX challenge
C0943630|T201|COMP|27957-0|LNC|Pyruvate^4H post XXX challenge|Pyruvate^4H post XXX challenge
C0943631|T201|COMP|27958-8|LNC|Proinsulin^4H post XXX challenge|Proinsulin^4H post XXX challenge
C0943632|T201|COMP|27959-6|LNC|Pyruvate^baseline|Pyruvate^baseline
C0943633|T201|COMP|27960-4|LNC|Coxsackievirus B5 RNA|Coxsackievirus B5 RNA
C0943634|T201|COMP|27961-2|LNC|Lactate^3H post XXX challenge|Lactate^3H post XXX challenge
C0943635|T201|COMP|27962-0|LNC|Butalbital|Butalbital
C0943636|T201|COMP|27963-8|LNC|Pyruvate^1H post XXX challenge|Pyruvate^1H post XXX challenge
C0943637|T201|COMP|27964-6|LNC|Streptococcus pneumoniae 6+26 Ab|Streptococcus pneumoniae 6+26 Ab
C0943638|T201|COMP|27965-3|LNC|Babesia microti Ab.IgM|Babesia microti Ab.IgM
C0943639|T201|COMP|27966-1|LNC|Legionella pneumophila atypical Ab|Legionella pneumophila atypical Ab
C0943640|T201|COMP|27967-9|LNC|Progesterone^baseline|Progesterone^baseline
C0943641|T201|COMP|27968-7|LNC|Pyruvate^2H post XXX challenge|Pyruvate^2H post XXX challenge
C0943642|T201|COMP|27969-5|LNC|Coxsackievirus A9 RNA|Coxsackievirus A9 RNA
C0943643|T201|COMP|27970-3|LNC|Pyruvate^3H post XXX challenge|Pyruvate^3H post XXX challenge
C0943644|T201|COMP|27971-1|LNC|Catecholamines^4H post XXX challenge|Catecholamines^4H post XXX challenge
C0943645|T201|COMP|27972-9|LNC|Histidine|Histidine
C0943646|T201|COMP|27973-7|LNC|3-Methylhistidine|3-Methylhistidine
C0943647|T201|COMP|27974-5|LNC|Arginine|Arginine
C0943648|T201|COMP|27975-2|LNC|Thyrotropin|Thyrotropin
C0943649|T201|COMP|27976-0|LNC|Lactate^post CFst|Lactate^post CFst
C0943650|T201|COMP|27978-6|LNC|Metanephrines/Creatinine|Metanephrines/Creatinine
C0943651|T201|COMP|27979-4|LNC|17-Ketogenic steroids|17-Ketogenic steroids
C0943652|T201|COMP|27981-0|LNC|2-Hydroxyisobutyrate|2-Hydroxyisobutyrate
C0943653|T201|COMP|27982-8|LNC|Borrelia burgdorferi 66kD Ab|Borrelia burgdorferi 66kD Ab
C0943654|T201|COMP|27984-4|LNC|SCA8 gene.CAG repeats|SCA8 gene.CAG repeats
C0943655|T201|COMP|27985-1|LNC|Borrelia burgdorferi 18kD Ab|Borrelia burgdorferi 18kD Ab
C0943656|T201|COMP|27986-9|LNC|Borrelia burgdorferi 28kD Ab|Borrelia burgdorferi 28kD Ab
C0943657|T201|COMP|27987-7|LNC|Thyroxine.free^baseline|Thyroxine.free^baseline
C0943658|T201|COMP|27988-5|LNC|Aldosterone^baseline|Aldosterone^baseline
C0943659|T201|COMP|27989-3|LNC|Thyroxine.free^1H post XXX challenge|Thyroxine.free^1H post XXX challenge
C0943660|T201|COMP|27990-1|LNC|Fibrinogen fragments|Fibrinogen fragments
C0943661|T201|COMP|27991-9|LNC|Fibrinogen fragments|Fibrinogen fragments
C0943662|T201|COMP|27992-7|LNC|Borrelia burgdorferi 23kD Ab|Borrelia burgdorferi 23kD Ab
C0943663|T201|COMP|27993-5|LNC|Sympathomimetics|Sympathomimetics
C0943664|T201|COMP|27995-0|LNC|Asparagine|Asparagine
C0943665|T201|COMP|27996-8|LNC|17-Hydroxyprogesterone^baseline|17-Hydroxyprogesterone^baseline
C0943666|T201|COMP|27997-6|LNC|Beta aminoadipate/Creatinine|Beta aminoadipate/Creatinine
C0943667|T201|COMP|27998-4|LNC|Estrone|Estrone
C0943668|T201|COMP|28000-8|LNC|von Willebrand factor Ag|von Willebrand factor Ag
C0943669|T201|COMP|28002-4|LNC|Borrelia burgdorferi 39kD Ab|Borrelia burgdorferi 39kD Ab
C0943670|T201|COMP|28003-2|LNC|Sodium/Potassium|Sodium/Potassium
C0943671|T201|COMP|28004-0|LNC|HIV 1 Ab.IgG|HIV 1 Ab.IgG
C0943672|T201|COMP|28005-7|LNC|MTHFR gene.c.677C>T|MTHFR gene.c.677C>T
C0943673|T201|COMP|28006-5|LNC|Hemoglobin F|Hemoglobin F
C0943674|T201|COMP|28009-9|LNC|Specimen volume|Specimen volume
C0943695|T201|COMP|28035-4|LNC|Escherichia coli shiga-like toxin|Escherichia coli shiga-like toxin
C0943696|T201|COMP|28036-2|LNC|Borrelia burgdorferi 39kD Ab.IgG|Borrelia burgdorferi 39kD Ab.IgG
C0943697|T201|COMP|28037-0|LNC|Borrelia burgdorferi 39kD Ab.IgM|Borrelia burgdorferi 39kD Ab.IgM
C0943698|T201|COMP|28038-8|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C0943699|T201|COMP|28039-6|LNC|Borrelia burgdorferi 66kD Ab.IgG|Borrelia burgdorferi 66kD Ab.IgG
C0943700|T201|COMP|28040-4|LNC|Borrelia burgdorferi 41kD Ab.IgG|Borrelia burgdorferi 41kD Ab.IgG
C0943701|T201|COMP|28042-0|LNC|Organophosphate pesticides|Organophosphate pesticides
C0943702|T201|COMP|28043-8|LNC|Borrelia burgdorferi 41kD Ab.IgM|Borrelia burgdorferi 41kD Ab.IgM
C0943703|T201|COMP|28045-3|LNC|Cortisol^1st specimen|Cortisol^1st specimen
C0943704|T201|COMP|28046-1|LNC|Cortisol^2nd specimen|Cortisol^2nd specimen
C0943705|T201|COMP|28047-9|LNC|Carbamate pesticides|Carbamate pesticides
C0943706|T201|COMP|28048-7|LNC|Borrelia burgdorferi 58kD Ab.IgG|Borrelia burgdorferi 58kD Ab.IgG
C0943707|T201|COMP|28049-5|LNC|1,2,4-Trichlorobenzene|1,2,4-Trichlorobenzene
C0943708|T201|COMP|28050-3|LNC|1,2,3-Trichlorobenzene|1,2,3-Trichlorobenzene
C0943709|T201|COMP|28052-9|LNC|HIV 1 Ab.IgG band pattern|HIV 1 Ab.IgG band pattern
C0943710|T201|COMP|28053-7|LNC|Borrelia burgdorferi 30kD Ab.IgG|Borrelia burgdorferi 30kD Ab.IgG
C0943711|T201|COMP|28054-5|LNC|Borrelia burgdorferi 93kD Ab.IgG|Borrelia burgdorferi 93kD Ab.IgG
C0943712|T201|COMP|28055-2|LNC|Borrelia burgdorferi 45kD Ab.IgG|Borrelia burgdorferi 45kD Ab.IgG
C0943713|T201|COMP|28057-8|LNC|Borrelia burgdorferi 23kD Ab.IgG|Borrelia burgdorferi 23kD Ab.IgG
C0943714|T201|COMP|28058-6|LNC|Borrelia burgdorferi 21kD Ab.IgG|Borrelia burgdorferi 21kD Ab.IgG
C0943715|T201|COMP|28059-4|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C0943716|T201|COMP|28060-2|LNC|MTHFR gene.c.1298A>C|MTHFR gene.c.1298A>C
C0943717|T201|COMP|28062-8|LNC|Borrelia burgdorferi 23kD Ab.IgM|Borrelia burgdorferi 23kD Ab.IgM
C0943718|T201|COMP|28063-6|LNC|Mercury^2nd specimen|Mercury^2nd specimen
C0943719|T201|COMP|28064-4|LNC|amLODIPine|amLODIPine
C0943720|T201|COMP|28066-9|LNC|Celecoxib|Celecoxib
C0943721|T201|COMP|28067-7|LNC|Hemoglobin F|Hemoglobin F
C0943722|T201|COMP|28068-5|LNC|Beta aminobutyrate|Beta aminobutyrate
C0943723|T201|COMP|28069-3|LNC|Meat fibers|Meat fibers
C0943724|T201|COMP|28070-1|LNC|Vegetable fibers|Vegetable fibers
C0943725|T201|COMP|28071-9|LNC|E selectin|E selectin
C0943726|T201|COMP|28072-7|LNC|Dihydrocodeine+Hydrocodeinone|Dihydrocodeine+Hydrocodeinone
C0943727|T201|COMP|28074-3|LNC|Tritium|Tritium
C0943728|T201|COMP|28076-8|LNC|SUMAtriptan|SUMAtriptan
C0943729|T201|COMP|28077-6|LNC|Hexachlorobutadiene|Hexachlorobutadiene
C0944135|T201|COMP|28541-1|LNC|Metamyelocytes/100 leukocytes|Metamyelocytes/100 leukocytes
C0944136|T201|COMP|28542-9|LNC|Platelet mean volume|Platelet mean volume
C0944137|T201|COMP|28543-7|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C0944138|T201|COMP|28545-2|LNC|Mucus|Mucus
C0944139|T201|COMP|28546-0|LNC|Neisseria meningitidis serogroup A Ab.IgG|Neisseria meningitidis serogroup A Ab.IgG
C0944140|T201|COMP|28547-8|LNC|Neisseria meningitidis serogroup C Ab.IgG|Neisseria meningitidis serogroup C Ab.IgG
C0944141|T201|COMP|28548-6|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C0944142|T201|COMP|28550-2|LNC|Cortisol|Cortisol
C0944143|T201|COMP|28551-0|LNC|Bladder tumor Ag|Bladder tumor Ag
C0944144|T201|COMP|28552-8|LNC|Cladosporium herbarum Ab.IgM|Cladosporium herbarum Ab.IgM
C0944145|T201|COMP|28553-6|LNC|Streptococcus pneumoniae 6+26 Ab^1st specimen|Streptococcus pneumoniae 6+26 Ab^1st specimen
C0944146|T201|COMP|28555-1|LNC|Nicotine+Cotinine|Nicotine+Cotinine
C0944147|T201|COMP|28556-9|LNC|Chlamydia trachomatis D+K Ab.IgG|Chlamydia trachomatis D+K Ab.IgG
C0944148|T201|COMP|28557-7|LNC|Chlamydia trachomatis D+K Ab.IgA|Chlamydia trachomatis D+K Ab.IgA
C0944149|T201|COMP|28558-5|LNC|Chlamydia trachomatis D+K Ab.IgM|Chlamydia trachomatis D+K Ab.IgM
C0944150|T201|COMP|28559-3|LNC|Hemoglobin A2|Hemoglobin A2
C0944151|T201|COMP|28560-1|LNC|Neuronal thread protein|Neuronal thread protein
C0944173|T201|COMP|28584-1|LNC|2-Oxoadipate/Creatinine|2-Oxoadipate/Creatinine
C0944174|T201|COMP|28585-8|LNC|4-Hydroxyphenylacetate/Creatinine|4-Hydroxyphenylacetate/Creatinine
C0944175|T201|COMP|28586-6|LNC|4-Hydroxyphenyllactate/Creatinine|4-Hydroxyphenyllactate/Creatinine
C0944176|T201|COMP|28587-4|LNC|Benzoate/Creatinine|Benzoate/Creatinine
C0944177|T201|COMP|28588-2|LNC|Beta alanine/Creatinine|Beta alanine/Creatinine
C0944178|T201|COMP|28590-8|LNC|Alpha aminobutyrate/Creatinine|Alpha aminobutyrate/Creatinine
C0944180|T201|COMP|28592-4|LNC|Beta aminoadipate/Creatinine|Beta aminoadipate/Creatinine
C0944181|T201|COMP|28594-0|LNC|3-Methylhistidine/Creatinine|3-Methylhistidine/Creatinine
C0944182|T201|COMP|28595-7|LNC|Taurine/Creatinine|Taurine/Creatinine
C0944183|T201|COMP|28596-5|LNC|Anserine/Creatinine|Anserine/Creatinine
C0944184|T201|COMP|28597-3|LNC|Carnosine/Creatinine|Carnosine/Creatinine
C0944185|T201|COMP|28599-9|LNC|Cystathionine/Creatinine|Cystathionine/Creatinine
C0944186|T201|COMP|28600-5|LNC|Phosphoserine/Creatinine|Phosphoserine/Creatinine
C0944187|T201|COMP|28602-1|LNC|Beta aminoisobutyrate/Creatinine|Beta aminoisobutyrate/Creatinine
C0944188|T201|COMP|28603-9|LNC|Asparagine/Creatinine|Asparagine/Creatinine
C0944189|T201|COMP|28604-7|LNC|Phosphoethanolamine/Creatinine|Phosphoethanolamine/Creatinine
C0944190|T201|COMP|28605-4|LNC|Ethanolamine/Creatinine|Ethanolamine/Creatinine
C0944191|T201|COMP|28607-0|LNC|Canine parvovirus Ab|Canine parvovirus Ab
C0944192|T201|COMP|28608-8|LNC|Tryptophan/Creatinine|Tryptophan/Creatinine
C0944193|T201|COMP|28609-6|LNC|Alpha aminobutyrate/Creatinine|Alpha aminobutyrate/Creatinine
C0944194|T201|COMP|28591-6|LNC|Amino beta guanidinopropionate/Creatinine|Amino beta guanidinopropionate/Creatinine
C0944195|T201|COMP|28612-0|LNC|Legionella sp Ab.IgM|Legionella sp Ab.IgM
C0944218|T201|COMP|28637-7|LNC|Base deficit|Base deficit
C0944219|T201|COMP|28638-5|LNC|Base excess|Base excess
C0944220|T201|COMP|28639-3|LNC|Base excess|Base excess
C0944221|T201|COMP|28640-1|LNC|Bicarbonate|Bicarbonate
C0944222|T201|COMP|28641-9|LNC|Bicarbonate|Bicarbonate
C0944223|T201|COMP|28642-7|LNC|Oxygen saturation|Oxygen saturation
C0944224|T201|COMP|28644-3|LNC|Carbon dioxide|Carbon dioxide
C0944225|T201|COMP|28645-0|LNC|Carbon dioxide|Carbon dioxide
C0944227|T201|COMP|28648-4|LNC|Oxygen|Oxygen
C0944229|T201|COMP|28652-6|LNC|Heparinoid|Heparinoid
C0944233|T201|COMP|28657-5|LNC|Coagulation factor X activated actual/Normal|Coagulation factor X activated actual/Normal
C0944234|T201|COMP|28658-3|LNC|Plasmin inhibitor actual/Normal|Plasmin inhibitor actual/Normal
C0944235|T201|COMP|28659-1|LNC|Prekallikrein actual/Normal|Prekallikrein actual/Normal
C0944619|T201|COMP|29113-8|LNC|Abacavir|Abacavir
C0944620|T201|COMP|29114-6|LNC|Amprenavir|Amprenavir
C0944621|T201|COMP|29117-9|LNC|Efavirenz|Efavirenz
C0944622|T201|COMP|29119-5|LNC|lamiVUDine|lamiVUDine
C0944623|T201|COMP|29120-3|LNC|Nelfinavir|Nelfinavir
C0944624|T201|COMP|29121-1|LNC|Nevirapine|Nevirapine
C0944625|T201|COMP|29122-9|LNC|Ritonavir|Ritonavir
C0944626|T201|COMP|29124-5|LNC|Stavudine|Stavudine
C0944627|T201|COMP|29125-2|LNC|Zalcitabine|Zalcitabine
C0944628|T201|COMP|29126-0|LNC|Zidovudine|Zidovudine
C0944640|T201|COMP|29141-9|LNC|Metanephrine|Metanephrine
C0944641|T201|COMP|29142-7|LNC|Metanephrines|Metanephrines
C0944642|T201|COMP|29143-5|LNC|1,4-Dimethylbenzene|1,4-Dimethylbenzene
C0944643|T201|COMP|29144-3|LNC|1,2-Dimethylbenzene|1,2-Dimethylbenzene
C0944644|T201|COMP|29145-0|LNC|1,3-Dimethylbenzene|1,3-Dimethylbenzene
C0944645|T201|COMP|29146-8|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C0944646|T201|COMP|29147-6|LNC|carBAMazepine 10,11-Epoxide.bound|carBAMazepine 10,11-Epoxide.bound
C0944647|T201|COMP|29148-4|LNC|carBAMazepine.bound|carBAMazepine.bound
C0944648|T201|COMP|29149-2|LNC|Mefloquine|Mefloquine
C0944649|T201|COMP|29150-0|LNC|Mefloquine|Mefloquine
C0944650|T201|COMP|29152-6|LNC|Somatotropin^5H post XXX challenge|Somatotropin^5H post XXX challenge
C0944651|T201|COMP|29153-4|LNC|Cancer Ag 15-3|Cancer Ag 15-3
C0944652|T201|COMP|29154-2|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0944653|T201|COMP|29155-9|LNC|Follitropin/Creatinine|Follitropin/Creatinine
C0944654|T201|COMP|29156-7|LNC|Lutropin|Lutropin
C0944655|T201|COMP|29157-5|LNC|Lutropin/Creatinine|Lutropin/Creatinine
C0944656|T201|COMP|29158-3|LNC|Opiates|Opiates
C0944657|T201|COMP|29159-1|LNC|Methadone|Methadone
C0944658|T201|COMP|29160-9|LNC|Benzodiazepines|Benzodiazepines
C0944659|T201|COMP|29161-7|LNC|Barbiturates|Barbiturates
C0944696|T201|COMP|29207-8|LNC|Amiodarone|Amiodarone
C0944697|T201|COMP|29208-6|LNC|Streptolysin O Ab|Streptolysin O Ab
C0944698|T201|COMP|29209-4|LNC|Benzodiazepines|Benzodiazepines
C0944699|T201|COMP|29210-2|LNC|Bilirubin.non-glucuronidated|Bilirubin.non-glucuronidated
C0944700|T201|COMP|29211-0|LNC|Caffeine|Caffeine
C0944701|T201|COMP|29212-8|LNC|carBAMazepine|carBAMazepine
C0944702|T201|COMP|29213-6|LNC|Ceruloplasmin|Ceruloplasmin
C0944703|T201|COMP|29214-4|LNC|Chloramphenicol|Chloramphenicol
C0944704|T201|COMP|29215-1|LNC|Digitoxin|Digitoxin
C0944705|T201|COMP|29216-9|LNC|Digoxin|Digoxin
C0944706|T201|COMP|29217-7|LNC|Disopyramide|Disopyramide
C0944707|T201|COMP|29218-5|LNC|Ethosuximide|Ethosuximide
C0944708|T201|COMP|29219-3|LNC|FLUoxetine|FLUoxetine
C0944709|T201|COMP|29220-1|LNC|Haptoglobin|Haptoglobin
C0944710|T201|COMP|29221-9|LNC|Mercury|Mercury
C0944711|T201|COMP|29222-7|LNC|Mexiletine|Mexiletine
C0944712|T201|COMP|29223-5|LNC|PHENobarbital|PHENobarbital
C0944713|T201|COMP|29224-3|LNC|Phenytoin|Phenytoin
C0944714|T201|COMP|29225-0|LNC|Primidone|Primidone
C0944715|T201|COMP|29226-8|LNC|quiNIDine|quiNIDine
C0944716|T201|COMP|29227-6|LNC|Salicylates|Salicylates
C0944717|T201|COMP|29228-4|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C0944718|T201|COMP|29231-8|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C0944719|T201|COMP|29233-4|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C0944720|T201|COMP|29234-2|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C0944721|T201|COMP|29235-9|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C0944722|T201|COMP|29238-3|LNC|Insulin|Insulin
C0944723|T201|COMP|29239-1|LNC|Triiodothyronine.free|Triiodothyronine.free
C0944724|T201|COMP|29240-9|LNC|Hyaluronate|Hyaluronate
C0944725|T201|COMP|29242-5|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C0944726|T201|COMP|29243-3|LNC|Thiodiglycolate|Thiodiglycolate
C0944727|T201|COMP|29244-1|LNC|Thiodiglycolate/Creatinine|Thiodiglycolate/Creatinine
C0944728|T201|COMP|29245-8|LNC|Zinc|Zinc
C0944729|T201|COMP|29247-4|LNC|Sirolimus|Sirolimus
C0944730|T201|COMP|29248-2|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C0944731|T201|COMP|29249-0|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0944732|T201|COMP|29250-8|LNC|Brucella sp Ab^1st specimen|Brucella sp Ab^1st specimen
C0944733|T201|COMP|29251-6|LNC|Brucella sp Ab^2nd specimen|Brucella sp Ab^2nd specimen
C0944735|T201|COMP|29254-0|LNC|Linezolid|Linezolid
C0944736|T201|COMP|29255-7|LNC|Linezolid|Linezolid
C0944737|T201|COMP|29256-5|LNC|Fat.microscopic observation|Fat.microscopic observation
C0944738|T201|COMP|29257-3|LNC|Mycoplasma pneumoniae DNA|Mycoplasma pneumoniae DNA
C0944739|T201|COMP|29258-1|LNC|Linezolid|Linezolid
C0944740|T201|COMP|29259-9|LNC|Monocytes.abnormal/100 leukocytes|Monocytes.abnormal/100 leukocytes
C0944741|T201|COMP|29260-7|LNC|Monocytes.abnormal|Monocytes.abnormal
C0944742|T201|COMP|29261-5|LNC|Lymphocytes.abnormal/100 leukocytes|Lymphocytes.abnormal/100 leukocytes
C0944743|T201|COMP|29262-3|LNC|Lymphocytes.abnormal|Lymphocytes.abnormal
C0944744|T201|COMP|29263-1|LNC|Fibrin degradation products|Fibrin degradation products
C0944745|T201|COMP|29264-9|LNC|Collection time|Collection time
C0944746|T201|COMP|29265-6|LNC|Calcium^^corrected for albumin|Calcium^^corrected for albumin
C0944747|T201|COMP|29266-4|LNC|Coproporphyrin|Coproporphyrin
C0944748|T201|COMP|29267-2|LNC|Protoporphyrin|Protoporphyrin
C0944755|T201|COMP|29276-3|LNC|Calcium|Calcium
C0944756|T201|COMP|29277-1|LNC|Carbon disulfide|Carbon disulfide
C0944757|T201|COMP|29278-9|LNC|Codeine|Codeine
C0944758|T201|COMP|29279-7|LNC|Ethylene glycol|Ethylene glycol
C0944759|T201|COMP|29280-5|LNC|Fibrin D-dimer|Fibrin D-dimer
C0944760|T201|COMP|29281-3|LNC|Glutathione reductase|Glutathione reductase
C0944761|T201|COMP|29282-1|LNC|Glutethimide|Glutethimide
C0944762|T201|COMP|29283-9|LNC|Hydrogen sulfide|Hydrogen sulfide
C0944763|T201|COMP|29284-7|LNC|Leucine|Leucine
C0944764|T201|COMP|29285-4|LNC|Methadone|Methadone
C0944765|T201|COMP|29286-2|LNC|Methamphetamine|Methamphetamine
C0944766|T201|COMP|29287-0|LNC|Morphine|Morphine
C0944767|T201|COMP|29288-8|LNC|Orphenadrine|Orphenadrine
C0944768|T201|COMP|29289-6|LNC|Phenylethylmalonamide|Phenylethylmalonamide
C0944769|T201|COMP|29290-4|LNC|Carbon disulfide|Carbon disulfide
C0944770|T201|COMP|29291-2|LNC|Glutethimide|Glutethimide
C0944771|T201|COMP|29292-0|LNC|Hydrogen sulfide|Hydrogen sulfide
C0944772|T201|COMP|29293-8|LNC|Leucine|Leucine
C0944773|T201|COMP|29295-3|LNC|Phenylethylmalonamide|Phenylethylmalonamide
C0944774|T201|COMP|29296-1|LNC|Dimethylbenzene|Dimethylbenzene
C0944783|T201|COMP|29310-0|LNC|Treponema pallidum|Treponema pallidum
C0944784|T201|COMP|29314-2|LNC|Adenovirus Ab|Adenovirus Ab
C0944785|T201|COMP|29315-9|LNC|Isoniazid 0.4 ug/mL|Isoniazid 0.4 ug/mL
C0944786|T201|COMP|29316-7|LNC|Thyrotropin^30M post XXX challenge|Thyrotropin^30M post XXX challenge
C0944787|T201|COMP|29317-5|LNC|Thyrotropin^1H post XXX challenge|Thyrotropin^1H post XXX challenge
C0944788|T201|COMP|29319-1|LNC|Streptococcus pneumoniae group B Ag|Streptococcus pneumoniae group B Ag
C0944789|T201|COMP|29320-9|LNC|Streptococcus pneumoniae group B Ag|Streptococcus pneumoniae group B Ag
C0944790|T201|COMP|29321-7|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C0944791|T201|COMP|29322-5|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C0944792|T201|COMP|29324-1|LNC|Cocaethylene|Cocaethylene
C0944793|T201|COMP|29325-8|LNC|Cocaethylene|Cocaethylene
C0944794|T201|COMP|29326-6|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0944795|T201|COMP|29327-4|LNC|HIV 1 Ab|HIV 1 Ab
C0944796|T201|COMP|29330-8|LNC|Glucose^4H post XXX challenge|Glucose^4H post XXX challenge
C0944797|T201|COMP|29331-6|LNC|Glucose^5H post XXX challenge|Glucose^5H post XXX challenge
C0944798|T201|COMP|29332-4|LNC|Glucose^2.5H post XXX challenge|Glucose^2.5H post XXX challenge
C0944799|T201|COMP|22572-2|LNC|Saccharomonospora viridis Ab|Saccharomonospora viridis Ab
C0944800|T201|COMP|29334-0|LNC|Aspergillus fumigatus 2 Ab|Aspergillus fumigatus 2 Ab
C0944801|T201|COMP|29335-7|LNC|Mexiletine|Mexiletine
C0944802|T201|COMP|29336-5|LNC|Mexiletine|Mexiletine
C0944803|T201|COMP|29337-3|LNC|Morphine.free|Morphine.free
C0944804|T201|COMP|29338-1|LNC|Flecainide|Flecainide
C0944805|T201|COMP|29339-9|LNC|Flecainide|Flecainide
C0944806|T201|COMP|29340-7|LNC|Cells.CD71|Cells.CD71
C0944807|T201|COMP|29341-5|LNC|Cells.CD11b|Cells.CD11b
C0944808|T201|COMP|29342-3|LNC|Methylmalonate|Methylmalonate
C0944809|T201|COMP|29343-1|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0944810|T201|COMP|29344-9|LNC|LORazepam|LORazepam
C0944811|T201|COMP|29345-6|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C0944812|T201|COMP|29346-4|LNC|Chloramphenicol|Chloramphenicol
C0944813|T201|COMP|29347-2|LNC|Chloramphenicol|Chloramphenicol
C0944814|T201|COMP|29348-0|LNC|ALPRAZolam|ALPRAZolam
C0944815|T201|COMP|29349-8|LNC|Potassium^post dialysis|Potassium^post dialysis
C0944816|T201|COMP|29350-6|LNC|Cells.CD42|Cells.CD42
C0944817|T201|COMP|29351-4|LNC|Rheumatoid factor|Rheumatoid factor
C0944818|T201|COMP|29352-2|LNC|Salicylates|Salicylates
C0944819|T201|COMP|29353-0|LNC|17-Ketosteroids.total neutral|17-Ketosteroids.total neutral
C0944820|T201|COMP|29354-8|LNC|Reovirus Ab|Reovirus Ab
C0944821|T201|COMP|29355-5|LNC|Reovirus Ab|Reovirus Ab
C0944822|T201|COMP|29356-3|LNC|fentaNYL|fentaNYL
C0944823|T201|COMP|29359-7|LNC|Parainfluenza virus 2 Ab|Parainfluenza virus 2 Ab
C0944824|T201|COMP|29361-3|LNC|Streptococcus pneumoniae group B Ag|Streptococcus pneumoniae group B Ag
C0944825|T201|COMP|29363-9|LNC|Cortisol^1.5H post XXX challenge|Cortisol^1.5H post XXX challenge
C0944826|T201|COMP|29364-7|LNC|Magnesium|Magnesium
C0944827|T201|COMP|29365-4|LNC|Magnesium|Magnesium
C0944828|T201|COMP|29367-0|LNC|Parainfluenza virus 2 Ab|Parainfluenza virus 2 Ab
C0944829|T201|COMP|29368-8|LNC|Parainfluenza virus 3 Ab|Parainfluenza virus 3 Ab
C0944830|T201|COMP|29369-6|LNC|N-acetylprocainamide/Procainamide|N-acetylprocainamide/Procainamide
C0944831|T201|COMP|29371-2|LNC|cloZAPine^peak|cloZAPine^peak
C0944832|T201|COMP|29372-0|LNC|Codeine|Codeine
C0944833|T201|COMP|29373-8|LNC|Ethchlorvynol|Ethchlorvynol
C0944834|T201|COMP|29375-3|LNC|Methanol|Methanol
C0944835|T201|COMP|29376-1|LNC|Narcotics|Narcotics
C0944836|T201|COMP|29377-9|LNC|Narcotics|Narcotics
C0944837|T201|COMP|29378-7|LNC|Insulin^4H post XXX challenge|Insulin^4H post XXX challenge
C0944838|T201|COMP|29379-5|LNC|Insulin^6H post XXX challenge|Insulin^6H post XXX challenge
C0944839|T201|COMP|29380-3|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0944840|T201|COMP|29381-1|LNC|Meprobamate|Meprobamate
C0944841|T201|COMP|29382-9|LNC|Warfarin|Warfarin
C0944842|T201|COMP|29384-5|LNC|diazePAM|diazePAM
C0944843|T201|COMP|29385-2|LNC|Nordiazepam|Nordiazepam
C0944844|T201|COMP|29386-0|LNC|chlorproMAZINE|chlorproMAZINE
C0944845|T201|COMP|29388-6|LNC|Methaqualone|Methaqualone
C0944846|T201|COMP|29389-4|LNC|Acetaminophen|Acetaminophen
C0944847|T201|COMP|29390-2|LNC|Parathyrin.mid molecule|Parathyrin.mid molecule
C0944848|T201|COMP|29391-0|LNC|Gastrin^2H post XXX challenge|Gastrin^2H post XXX challenge
C0944849|T201|COMP|29393-6|LNC|Gastrin^3H post XXX challenge|Gastrin^3H post XXX challenge
C0944850|T201|COMP|29394-4|LNC|Gastrin^2.5H post XXX challenge|Gastrin^2.5H post XXX challenge
C0944851|T201|COMP|29395-1|LNC|Gastrin^post CFst|Gastrin^post CFst
C0944852|T201|COMP|29396-9|LNC|Gastrin^1.5H post XXX challenge|Gastrin^1.5H post XXX challenge
C0944853|T201|COMP|29397-7|LNC|Gastrin^30M pre XXX challenge|Gastrin^30M pre XXX challenge
C0944854|T201|COMP|29398-5|LNC|Gastrin^1M pre XXX challenge|Gastrin^1M pre XXX challenge
C0944855|T201|COMP|29399-3|LNC|clonazePAM|clonazePAM
C0944856|T201|COMP|29400-9|LNC|Meperidine|Meperidine
C0944857|T201|COMP|29401-7|LNC|Disopyramide|Disopyramide
C0944858|T201|COMP|29402-5|LNC|Trimipramine|Trimipramine
C0944859|T201|COMP|29403-3|LNC|Thiothixene|Thiothixene
C0944860|T201|COMP|29404-1|LNC|Thiothixene|Thiothixene
C0944861|T201|COMP|29405-8|LNC|Maprotiline|Maprotiline
C0944862|T201|COMP|29406-6|LNC|Amitriptyline|Amitriptyline
C0944863|T201|COMP|29407-4|LNC|Nortriptyline|Nortriptyline
C0944864|T201|COMP|29408-2|LNC|Imipramine|Imipramine
C0944865|T201|COMP|29409-0|LNC|Desipramine|Desipramine
C0944866|T201|COMP|29410-8|LNC|Doxepin|Doxepin
C0944867|T201|COMP|29411-6|LNC|Nordoxepin|Nordoxepin
C0944868|T201|COMP|29413-2|LNC|Reovirus Ab|Reovirus Ab
C0944869|T201|COMP|29414-0|LNC|Parainfluenza virus 3 Ab|Parainfluenza virus 3 Ab
C0944870|T201|COMP|29415-7|LNC|Reovirus Ab|Reovirus Ab
C0944871|T201|COMP|29416-5|LNC|Adenovirus Ab|Adenovirus Ab
C0944872|T201|COMP|29417-3|LNC|Parainfluenza virus 1 Ab|Parainfluenza virus 1 Ab
C0944936|T201|COMP|29492-6|LNC|Methicillin|Methicillin
C0944937|T201|COMP|29493-4|LNC|Colistin|Colistin
C0944938|T201|COMP|29495-9|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C0944939|T201|COMP|29496-7|LNC|Platelet associated Ab.IgA|Platelet associated Ab.IgA
C0944940|T201|COMP|29498-3|LNC|Platelet associated Ab.IgM|Platelet associated Ab.IgM
C0944941|T201|COMP|29499-1|LNC|Selenium|Selenium
C0944942|T201|COMP|29500-6|LNC|2-Hydroxyadipate/Creatinine|2-Hydroxyadipate/Creatinine
C0944943|T201|COMP|29501-4|LNC|2-Hydroxyisobutyrate/Creatinine|2-Hydroxyisobutyrate/Creatinine
C0944944|T201|COMP|29502-2|LNC|2-Hydroxyglutarate/Creatinine|2-Hydroxyglutarate/Creatinine
C0944945|T201|COMP|29503-0|LNC|2-Hydroxyisocaproate/Creatinine|2-Hydroxyisocaproate/Creatinine
C0944946|T201|COMP|29504-8|LNC|2-Hydroxyisovalerate/Creatinine|2-Hydroxyisovalerate/Creatinine
C0944947|T201|COMP|29505-5|LNC|2-Hydroxy-3-Methylvalerate/Creatinine|2-Hydroxy-3-Methylvalerate/Creatinine
C0944948|T201|COMP|29506-3|LNC|2-Oxoadipate/Creatinine|2-Oxoadipate/Creatinine
C0944949|T201|COMP|29507-1|LNC|Alpha ketoglutarate/Creatinine|Alpha ketoglutarate/Creatinine
C0944950|T201|COMP|29508-9|LNC|3-Hydroxyadipate/Creatinine|3-Hydroxyadipate/Creatinine
C0944951|T201|COMP|29509-7|LNC|Beta hydroxybutyrate/Creatinine|Beta hydroxybutyrate/Creatinine
C0944952|T201|COMP|29510-5|LNC|3-Hydroxyglutarate/Creatinine|3-Hydroxyglutarate/Creatinine
C0944953|T201|COMP|29511-3|LNC|3-Hydroxyisobutyrate/Creatinine|3-Hydroxyisobutyrate/Creatinine
C0944954|T201|COMP|29512-1|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C0944955|T201|COMP|16708-0|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C0944956|T201|COMP|29514-7|LNC|3-Hydroxyisovalerate/Creatinine|3-Hydroxyisovalerate/Creatinine
C0944957|T201|COMP|29515-4|LNC|3-Hydroxypropionate/Creatinine|3-Hydroxypropionate/Creatinine
C0944958|T201|COMP|29516-2|LNC|3-Hydroxyvalerate/Creatinine|3-Hydroxyvalerate/Creatinine
C0944959|T201|COMP|29517-0|LNC|Vanillylmandelate/Creatinine|Vanillylmandelate/Creatinine
C0944960|T201|COMP|29518-8|LNC|3-Methylglutarate/Creatinine|3-Methylglutarate/Creatinine
C0944961|T201|COMP|29519-6|LNC|4-Hydroxyphenylpyruvate/Creatinine|4-Hydroxyphenylpyruvate/Creatinine
C0944962|T201|COMP|29520-4|LNC|5-Hydroxyindoleacetate/Creatinine|5-Hydroxyindoleacetate/Creatinine
C0944963|T201|COMP|29521-2|LNC|5-Hydroxyhexanoate/Creatinine|5-Hydroxyhexanoate/Creatinine
C0944964|T201|COMP|29522-0|LNC|5-Oxoproline/Creatinine|5-Oxoproline/Creatinine
C0944965|T201|COMP|29523-8|LNC|2-Ethyl-3-Hydroxypropionate/Creatinine|2-Ethyl-3-Hydroxypropionate/Creatinine
C0944966|T201|COMP|29524-6|LNC|Acetoacetate/Creatinine|Acetoacetate/Creatinine
C0944967|T201|COMP|29526-1|LNC|Azelate/Creatinine|Azelate/Creatinine
C0944968|T201|COMP|29527-9|LNC|Citrate/Creatinine|Citrate/Creatinine
C0944969|T201|COMP|29529-5|LNC|Acetaminophen|Acetaminophen
C0944970|T201|COMP|29531-1|LNC|diphenhydrAMINE|diphenhydrAMINE
C0944971|T201|COMP|29532-9|LNC|Methadone|Methadone
C0944972|T201|COMP|29533-7|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C0944973|T201|COMP|29535-2|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C0944974|T201|COMP|29536-0|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C0944975|T201|COMP|29537-8|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C0944976|T201|COMP|29538-6|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C0944977|T201|COMP|29540-2|LNC|E-cadherin|E-cadherin
C0944978|T201|COMP|29541-0|LNC|HIV 1 RNA|HIV 1 RNA
C0944979|T201|COMP|29542-8|LNC|Beta-N-acetylhexosaminidase|Beta-N-acetylhexosaminidase
C0944988|T201|COMP|29553-5|LNC|Age|Age
C0944992|T201|COMP|29558-4|LNC|Enterovirus RNA|Enterovirus RNA
C0944993|T201|COMP|29559-2|LNC|Haemophilus ducreyi DNA|Haemophilus ducreyi DNA
C0944994|T201|COMP|29560-0|LNC|Anaplasma phagocytophilum DNA|Anaplasma phagocytophilum DNA
C0944995|T201|COMP|29561-8|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C0944996|T201|COMP|29562-6|LNC|Jamestown canyon virus Ab|Jamestown canyon virus Ab
C0944997|T201|COMP|29563-4|LNC|La Crosse virus Ab|La Crosse virus Ab
C0944998|T201|COMP|29564-2|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C0944999|T201|COMP|29565-9|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C0945000|T201|COMP|29566-7|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C0945001|T201|COMP|29567-5|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C0945002|T201|COMP|29568-3|LNC|West Nile virus Ab|West Nile virus Ab
C0945003|T201|COMP|29569-1|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C0945004|T201|COMP|29570-9|LNC|West Nile virus Ab|West Nile virus Ab
C0945005|T201|COMP|29571-7|LNC|Phenylalanine|Phenylalanine
C0945006|T201|COMP|29572-5|LNC|Phenylalanine|Phenylalanine
C0945007|T201|COMP|29573-3|LNC|Phenylalanine|Phenylalanine
C0945008|T201|COMP|29574-1|LNC|Thyrotropin|Thyrotropin
C0945009|T201|COMP|29575-8|LNC|Thyrotropin|Thyrotropin
C0945010|T201|COMP|29576-6|LNC|Bacterial susceptibility panel|Bacterial susceptibility panel
C0945011|T201|COMP|29577-4|LNC|Fungal susceptibility panel|Fungal susceptibility panel
C0945012|T201|COMP|29579-0|LNC|Mycobacterial susceptibility panel|Mycobacterial susceptibility panel
C0945013|T201|COMP|29580-8|LNC|Differential panel|Differential panel
C0945014|T201|COMP|29581-6|LNC|Differential panel|Differential panel
C0945015|T201|COMP|29582-4|LNC|Differential panel|Differential panel
C0945016|T201|COMP|29584-0|LNC|Differential panel|Differential panel
C0945017|T201|COMP|29585-7|LNC|Immunoelectrophoresis panel|Immunoelectrophoresis panel
C0945018|T201|COMP|29586-5|LNC|Immunoelectrophoresis panel|Immunoelectrophoresis panel
C0945019|T201|COMP|29587-3|LNC|Toxicology panel|Toxicology panel
C0945020|T201|COMP|29588-1|LNC|Heavy metals panel|Heavy metals panel
C0945021|T201|COMP|29589-9|LNC|Heavy metals panel|Heavy metals panel
C0945022|T201|COMP|29591-5|LNC|Enterovirus RNA|Enterovirus RNA
C0945023|T201|COMP|29592-3|LNC|Amphetamine|Amphetamine
C0945024|T201|COMP|29593-1|LNC|Cells.Ki-67 nuclear Ag/100 cells|Cells.Ki-67 nuclear Ag/100 cells
C0945025|T201|COMP|29594-9|LNC|CD45RO Ag|CD45RO Ag
C0945026|T201|COMP|29596-4|LNC|CD25 Ag|CD25 Ag
C0945027|T201|COMP|29597-2|LNC|Mephentermine|Mephentermine
C0945028|T201|COMP|29598-0|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C0945029|T201|COMP|29599-8|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C0945030|T201|COMP|29600-4|LNC|Benzfetamine|Benzfetamine
C0945031|T201|COMP|29601-2|LNC|Phenylpropanolamine|Phenylpropanolamine
C0945032|T201|COMP|29602-0|LNC|Chlorphentermine|Chlorphentermine
C0945033|T201|COMP|29604-6|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C0945034|T201|COMP|29605-3|LNC|Appearance|Appearance
C0945035|T201|COMP|29606-1|LNC|Appearance|Appearance
C0945036|T201|COMP|29607-9|LNC|Tropheryma whippelii DNA|Tropheryma whippelii DNA
C0945037|T201|COMP|29609-5|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C0945038|T201|COMP|29611-1|LNC|Ethchlorvynol|Ethchlorvynol
C0945039|T201|COMP|29613-7|LNC|Phendimetrazine|Phendimetrazine
C0945040|T201|COMP|29614-5|LNC|Phenmetrazine|Phenmetrazine
C0945041|T201|COMP|29615-2|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C0945042|T201|COMP|29618-6|LNC|Stachybotrys chartarum Ab.IgE.RAST class|Stachybotrys chartarum Ab.IgE.RAST class
C0945043|T201|COMP|29619-4|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C0945044|T201|COMP|29620-2|LNC|Zonisamide|Zonisamide
C0945045|T201|COMP|29621-0|LNC|3-Hydroxyadipate|3-Hydroxyadipate
C0945046|T201|COMP|29622-8|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C0945047|T201|COMP|29623-6|LNC|3-Hydroxydodecanoate|3-Hydroxydodecanoate
C0945048|T201|COMP|29624-4|LNC|3-Hydroxyglutarate|3-Hydroxyglutarate
C0945049|T201|COMP|29625-1|LNC|3-Hydroxypropionate|3-Hydroxypropionate
C0945051|T201|COMP|29627-7|LNC|3-Hydroxyvalerate|3-Hydroxyvalerate
C0945052|T201|COMP|29628-5|LNC|3-Methylcrotonylglycine|3-Methylcrotonylglycine
C0945053|T201|COMP|29629-3|LNC|3-Methylglutaconate|3-Methylglutaconate
C0945054|T201|COMP|29630-1|LNC|3-Methylglutarate|3-Methylglutarate
C0945055|T201|COMP|29631-9|LNC|N-acetylaspartate|N-acetylaspartate
C0945056|T201|COMP|29632-7|LNC|N-acetyltyrosine|N-acetyltyrosine
C0945057|T201|COMP|29633-5|LNC|CD122 Ag|CD122 Ag
C0945058|T201|COMP|29634-3|LNC|Terbutaline|Terbutaline
C0945059|T201|COMP|29636-8|LNC|Appearance|Appearance
C0945060|T201|COMP|29638-4|LNC|Specimen weight|Specimen weight
C0945061|T201|COMP|29639-2|LNC|Alkaline phosphatase|Alkaline phosphatase
C0945062|T201|COMP|29640-0|LNC|Isomaltase|Isomaltase
C0945063|T201|COMP|29641-8|LNC|Neutrophil cytoplasmic Ab.atypical|Neutrophil cytoplasmic Ab.atypical
C0945064|T201|COMP|29642-6|LNC|Neutrophil cytoplasmic Ab.classic.atypical|Neutrophil cytoplasmic Ab.classic.atypical
C0945065|T201|COMP|29643-4|LNC|Myeloperoxidase Ab|Myeloperoxidase Ab
C0945066|T201|COMP|29644-2|LNC|Proteinase 3|Proteinase 3
C0945067|T201|COMP|29645-9|LNC|Echovirus+Coxsackievirus Ab.IgA|Echovirus+Coxsackievirus Ab.IgA
C0945068|T201|COMP|29646-7|LNC|Parainfluenza virus 2 Ab.IgM|Parainfluenza virus 2 Ab.IgM
C0945069|T201|COMP|29647-5|LNC|Interferon.beta Ab|Interferon.beta Ab
C0945070|T201|COMP|29648-3|LNC|Rickettsia australis Ab|Rickettsia australis Ab
C0945071|T201|COMP|29649-1|LNC|Rickettsia australis Ab|Rickettsia australis Ab
C0945072|T201|COMP|29651-7|LNC|Rickettsia honei Ab|Rickettsia honei Ab
C0945073|T201|COMP|29652-5|LNC|Dothiepin|Dothiepin
C0945074|T201|COMP|29653-3|LNC|Dothiepin|Dothiepin
C0945075|T201|COMP|29654-1|LNC|Temazepam|Temazepam
C0945076|T201|COMP|29656-6|LNC|Sympathomimetics|Sympathomimetics
C0945077|T201|COMP|29657-4|LNC|Bordetella pertussis Ab.IgA|Bordetella pertussis Ab.IgA
C0945078|T201|COMP|29658-2|LNC|Bordetella pertussis Ab.IgM|Bordetella pertussis Ab.IgM
C0945079|T201|COMP|29660-8|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0945080|T201|COMP|29661-6|LNC|Dengue virus Ab.IgG|Dengue virus Ab.IgG
C0945081|T201|COMP|29662-4|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0945082|T201|COMP|29665-7|LNC|Rickettsia conorii Ab|Rickettsia conorii Ab
C0945083|T201|COMP|29667-3|LNC|Parainfluenza virus 2 Ab.IgM|Parainfluenza virus 2 Ab.IgM
C0945084|T201|COMP|29669-9|LNC|Rickettsia australis Ab|Rickettsia australis Ab
C0945085|T201|COMP|29670-7|LNC|Rickettsia honei Ab|Rickettsia honei Ab
C0945086|T201|COMP|29671-5|LNC|Rickettsia honei Ab|Rickettsia honei Ab
C0945087|T201|COMP|29673-1|LNC|Bordetella pertussis Ab.IgM|Bordetella pertussis Ab.IgM
C0945088|T201|COMP|29674-9|LNC|Bordetella pertussis Ab.IgG|Bordetella pertussis Ab.IgG
C0945089|T201|COMP|29675-6|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0945090|T201|COMP|29676-4|LNC|Dengue virus Ab.IgG|Dengue virus Ab.IgG
C0945091|T201|COMP|29678-0|LNC|Rickettsia conorii Ab|Rickettsia conorii Ab
C0945092|T201|COMP|29679-8|LNC|Rickettsia sibirica Ab|Rickettsia sibirica Ab
C0945093|T201|COMP|29680-6|LNC|Rickettsia akari Ab|Rickettsia akari Ab
C0945094|T201|COMP|29682-2|LNC|Rickettsia prowazekii Ab|Rickettsia prowazekii Ab
C0945095|T201|COMP|29683-0|LNC|Rickettsia prowazekii Ab|Rickettsia prowazekii Ab
C0945096|T201|COMP|29684-8|LNC|Rickettsia typhi Ab|Rickettsia typhi Ab
C0945097|T201|COMP|29685-5|LNC|Rickettsia typhi Ab|Rickettsia typhi Ab
C0945098|T201|COMP|29686-3|LNC|Orientia tsutsugamushi Gilliam Ab|Orientia tsutsugamushi Gilliam Ab
C0945099|T201|COMP|29687-1|LNC|Orientia tsutsugamushi Gilliam Ab|Orientia tsutsugamushi Gilliam Ab
C0945100|T201|COMP|29689-7|LNC|Orientia tsutsugamushi Karp Ab|Orientia tsutsugamushi Karp Ab
C0945101|T201|COMP|29690-5|LNC|Orientia tsutsugamushi Kato Ab|Orientia tsutsugamushi Kato Ab
C0945102|T201|COMP|29691-3|LNC|Orientia tsutsugamushi Kato Ab|Orientia tsutsugamushi Kato Ab
C0945103|T201|COMP|29692-1|LNC|Orientia tsutsugamushi Litchfield Ab|Orientia tsutsugamushi Litchfield Ab
C0945104|T201|COMP|29693-9|LNC|Orientia tsutsugamushi Litchfield Ab|Orientia tsutsugamushi Litchfield Ab
C0945105|T201|COMP|29694-7|LNC|Leptospira interrogans serovar Celledoni Ab|Leptospira interrogans serovar Celledoni Ab
C0945106|T201|COMP|29695-4|LNC|Leptospira interrogans serovar Bulgarica Ab|Leptospira interrogans serovar Bulgarica Ab
C0945107|T201|COMP|29696-2|LNC|Leptospira interrogans serovar Cynopteri Ab|Leptospira interrogans serovar Cynopteri Ab
C0945108|T201|COMP|29697-0|LNC|Leptospira interrogans serovar Djasiman Ab|Leptospira interrogans serovar Djasiman Ab
C0945109|T201|COMP|29698-8|LNC|Leptospira interrogans serovar Javanica Ab|Leptospira interrogans serovar Javanica Ab
C0945110|T201|COMP|29699-6|LNC|Leptospira interrogans serovar Panama Ab|Leptospira interrogans serovar Panama Ab
C0945111|T201|COMP|29700-2|LNC|Leptospira interrogans serovar Shermani Ab|Leptospira interrogans serovar Shermani Ab
C0945112|T201|COMP|29701-0|LNC|Leptospira interrogans serovar Zanoni Ab|Leptospira interrogans serovar Zanoni Ab
C0945113|T201|COMP|29702-8|LNC|Rickettsia conorii Ab|Rickettsia conorii Ab
C0945114|T201|COMP|29703-6|LNC|Rickettsia sibirica Ab|Rickettsia sibirica Ab
C0945115|T201|COMP|29704-4|LNC|Rickettsia sibirica Ab|Rickettsia sibirica Ab
C0945116|T201|COMP|29705-1|LNC|Rickettsia rickettsii Ab|Rickettsia rickettsii Ab
C0945117|T201|COMP|29706-9|LNC|Rickettsia rickettsii Ab|Rickettsia rickettsii Ab
C0945118|T201|COMP|29707-7|LNC|Rickettsia akari Ab|Rickettsia akari Ab
C0945119|T201|COMP|29708-5|LNC|Rickettsia akari Ab|Rickettsia akari Ab
C0945120|T201|COMP|29709-3|LNC|Rickettsia prowazekii Ab|Rickettsia prowazekii Ab
C0945121|T201|COMP|29711-9|LNC|Rickettsia typhi Ab|Rickettsia typhi Ab
C0945122|T201|COMP|29712-7|LNC|Rickettsia typhi Ab|Rickettsia typhi Ab
C0945123|T201|COMP|29714-3|LNC|Orientia tsutsugamushi Gilliam Ab|Orientia tsutsugamushi Gilliam Ab
C0945124|T201|COMP|29715-0|LNC|Orientia tsutsugamushi Karp Ab|Orientia tsutsugamushi Karp Ab
C0945125|T201|COMP|29716-8|LNC|Orientia tsutsugamushi Karp Ab|Orientia tsutsugamushi Karp Ab
C0945126|T201|COMP|29717-6|LNC|Orientia tsutsugamushi Kato Ab|Orientia tsutsugamushi Kato Ab
C0945127|T201|COMP|29718-4|LNC|Orientia tsutsugamushi Kato Ab|Orientia tsutsugamushi Kato Ab
C0945128|T201|COMP|29721-8|LNC|Influenza virus C Ag|Influenza virus C Ag
C0945129|T201|COMP|29722-6|LNC|Chlamydophila pneumoniae Ag|Chlamydophila pneumoniae Ag
C0945130|T201|COMP|29723-4|LNC|Bordetella parapertussis DNA|Bordetella parapertussis DNA
C0945131|T201|COMP|29725-9|LNC|Leptospira interrogans serovar Bulgarica Ab|Leptospira interrogans serovar Bulgarica Ab
C0945132|T201|COMP|29726-7|LNC|Leptospira interrogans serovar Cynopteri Ab|Leptospira interrogans serovar Cynopteri Ab
C0945133|T201|COMP|29727-5|LNC|Leptospira interrogans serovar Djasiman Ab|Leptospira interrogans serovar Djasiman Ab
C0945134|T201|COMP|29728-3|LNC|Leptospira interrogans serovar Javanica Ab|Leptospira interrogans serovar Javanica Ab
C0945135|T201|COMP|29729-1|LNC|Leptospira interrogans serovar Panama Ab|Leptospira interrogans serovar Panama Ab
C0945136|T201|COMP|29730-9|LNC|Leptospira interrogans serovar Shermani Ab|Leptospira interrogans serovar Shermani Ab
C0945137|T201|COMP|29731-7|LNC|Leptospira interrogans serovar Zanoni Ab|Leptospira interrogans serovar Zanoni Ab
C0945138|T201|COMP|29732-5|LNC|Leptospira interrogans serovar Robinsoni Ab|Leptospira interrogans serovar Robinsoni Ab
C0945139|T201|COMP|29734-1|LNC|Leptospira interrogans serovar Szwajizak Ab|Leptospira interrogans serovar Szwajizak Ab
C0945140|T201|COMP|29735-8|LNC|Leptospira interrogans serovar Medanensis Ab|Leptospira interrogans serovar Medanensis Ab
C0945141|T201|COMP|29736-6|LNC|Rickettsia sibirica Ab|Rickettsia sibirica Ab
C0945142|T201|COMP|29737-4|LNC|Rickettsia rickettsii Ab|Rickettsia rickettsii Ab
C0945143|T201|COMP|29738-2|LNC|Leptospira interrogans serovar Robinsoni Ab|Leptospira interrogans serovar Robinsoni Ab
C0945144|T201|COMP|29740-8|LNC|Leptospira interrogans serovar Szwajizak Ab|Leptospira interrogans serovar Szwajizak Ab
C0945145|T201|COMP|29741-6|LNC|Leptospira interrogans serovar Medanensis Ab|Leptospira interrogans serovar Medanensis Ab
C0945146|T201|COMP|29742-4|LNC|Date last dose|Date last dose
C0945147|T201|COMP|29743-2|LNC|Cryofibrinogen|Cryofibrinogen
C0945148|T201|COMP|29744-0|LNC|Cryofibrinogen|Cryofibrinogen
C0945149|T201|COMP|29745-7|LNC|Cryoglobulin|Cryoglobulin
C0945150|T201|COMP|29746-5|LNC|Cryoglobulin|Cryoglobulin
C0945151|T201|COMP|29748-1|LNC|Protein|Protein
C0945163|T201|COMP|29760-6|LNC|Bilirubin.glucuronidated|Bilirubin.glucuronidated
C0945166|T201|COMP|29763-0|LNC|Protoporphyrin.zinc|Protoporphyrin.zinc
C0945167|T201|COMP|29764-8|LNC|Iron|Iron
C0945168|T201|COMP|29765-5|LNC|Cholesterol|Cholesterol
C0945169|T201|COMP|29766-3|LNC|Triglyceride|Triglyceride
C0945170|T201|COMP|25088-6|LNC|4-Hydroxyphenylacetate/Creatinine|4-Hydroxyphenylacetate/Creatinine
C0945171|T201|COMP|25090-2|LNC|Benzoate/Creatinine|Benzoate/Creatinine
C0945172|T201|COMP|25112-4|LNC|Lactate/Creatinine|Lactate/Creatinine
C0945173|T201|COMP|25117-3|LNC|Methylsuccinate/Creatinine|Methylsuccinate/Creatinine
C0945174|T201|COMP|25119-9|LNC|N-acetyltyrosine/Creatinine|N-acetyltyrosine/Creatinine
C0945175|T201|COMP|25120-7|LNC|Octanoate/Creatinine|Octanoate/Creatinine
C0945176|T201|COMP|25121-5|LNC|Octenedioate/Creatinine|Octenedioate/Creatinine
C0945177|T201|COMP|25126-4|LNC|Phenylpyruvate/Creatinine|Phenylpyruvate/Creatinine
C0945178|T201|COMP|25130-6|LNC|Pyridinoline/Creatinine|Pyridinoline/Creatinine
C0945179|T201|COMP|25134-8|LNC|Sebacate/Creatinine|Sebacate/Creatinine
C0945180|T201|COMP|25139-7|LNC|Tryptophan/Creatinine|Tryptophan/Creatinine
C0945181|T201|COMP|25147-0|LNC|Calcium carbonate crystals|Calcium carbonate crystals
C0945182|T201|COMP|25156-1|LNC|Eosinophils|Eosinophils
C0945183|T201|COMP|25178-5|LNC|Amikacin 30.0 ug/mL|Amikacin 30.0 ug/mL
C0945184|T201|COMP|25182-7|LNC|Kanamycin 5.0 ug/mL|Kanamycin 5.0 ug/mL
C0945185|T201|COMP|25184-3|LNC|rifAMPin 14.0 ug/mL|rifAMPin 14.0 ug/mL
C0945186|T201|COMP|25187-6|LNC|Ethambutol 7.5 ug/mL|Ethambutol 7.5 ug/mL
C0945187|T201|COMP|25191-8|LNC|Clarithromycin 16.0 ug/mL|Clarithromycin 16.0 ug/mL
C0945188|T201|COMP|25199-1|LNC|Rifabutin 1.0 ug/mL|Rifabutin 1.0 ug/mL
C0945189|T201|COMP|25202-3|LNC|rifAMPin 1.0 ug/mL|rifAMPin 1.0 ug/mL
C0945190|T201|COMP|25223-9|LNC|Doxycycline 30.0 ug/mL|Doxycycline 30.0 ug/mL
C0945191|T201|COMP|25232-0|LNC|Nafcillin|Nafcillin
C0945192|T201|COMP|25237-9|LNC|Cefonicid|Cefonicid
C0945193|T201|COMP|25240-3|LNC|cefOXitin|cefOXitin
C0945194|T201|COMP|25244-5|LNC|cefTRIAXone|cefTRIAXone
C0945195|T201|COMP|25249-4|LNC|Clindamycin|Clindamycin
C0945196|T201|COMP|25252-8|LNC|Dicloxacillin|Dicloxacillin
C0945197|T201|COMP|25257-7|LNC|Imipenem|Imipenem
C0945198|T201|COMP|25261-9|LNC|Nalidixate|Nalidixate
C0945199|T201|COMP|25264-3|LNC|Ofloxacin|Ofloxacin
C0945200|T201|COMP|25265-0|LNC|Oxacillin|Oxacillin
C0945201|T201|COMP|25273-4|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0945203|T201|COMP|25308-8|LNC|Ammonia|Ammonia
C0945204|T201|COMP|25311-2|LNC|Amylase|Amylase
C0945205|T201|COMP|25315-3|LNC|11-Deoxycortisol|11-Deoxycortisol
C0945206|T201|COMP|25324-5|LNC|Arsenic/Creatinine|Arsenic/Creatinine
C0945207|T201|COMP|25325-2|LNC|Ascaris sp Ab.IgE|Ascaris sp Ab.IgE
C0945209|T201|COMP|25361-7|LNC|Caffeine|Caffeine
C0945210|T201|COMP|25362-5|LNC|Calcium|Calcium
C0945211|T201|COMP|25365-8|LNC|Carnosine|Carnosine
C0945212|T201|COMP|25370-8|LNC|Chocolate Ab.IgE.RAST class|Chocolate Ab.IgE.RAST class
C0945213|T201|COMP|25375-7|LNC|Chymotrypsin|Chymotrypsin
C0945214|T201|COMP|25379-9|LNC|Cobalt|Cobalt
C0945215|T201|COMP|25382-3|LNC|Cortisone|Cortisone
C0945216|T201|COMP|25387-2|LNC|Cyanide|Cyanide
C0945217|T201|COMP|25390-6|LNC|Cytokeratin 19|Cytokeratin 19
C0945218|T201|COMP|25398-9|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0945219|T201|COMP|25422-7|LNC|Schistosoma sp Ab|Schistosoma sp Ab
C0945220|T201|COMP|25424-3|LNC|Trypanosoma sp Ab|Trypanosoma sp Ab
C0945221|T201|COMP|25427-6|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C0945222|T201|COMP|25431-8|LNC|Glycine|Glycine
C0945223|T201|COMP|25435-9|LNC|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C0945224|T201|COMP|32690-0|LNC|Homocysteine|Homocysteine
C0945225|T201|COMP|25456-5|LNC|Lactoglobulin Ab.IgA.RAST class|Lactoglobulin Ab.IgA.RAST class
C0945226|T201|COMP|25466-4|LNC|Manganese|Manganese
C0945227|T201|COMP|25484-7|LNC|Nefazodone|Nefazodone
C0945228|T201|COMP|25492-0|LNC|Oxipurinol|Oxipurinol
C0945229|T201|COMP|25494-6|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C0945230|T201|COMP|25499-5|LNC|Adrenal cortex Ab|Adrenal cortex Ab
C0945231|T201|COMP|25502-6|LNC|Phosphoethanolamine|Phosphoethanolamine
C0945232|T201|COMP|25507-5|LNC|Pregnenolone|Pregnenolone
C0945233|T201|COMP|25510-9|LNC|Proline|Proline
C0945234|T201|COMP|25514-1|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0945235|T201|COMP|25521-6|LNC|Selenium|Selenium
C0945236|T201|COMP|25525-7|LNC|Serpula lacrymans Ab.IgE.RAST class|Serpula lacrymans Ab.IgE.RAST class
C0945237|T201|COMP|25527-3|LNC|Silver|Silver
C0945238|T201|COMP|25547-1|LNC|Tyrosine|Tyrosine
C0945239|T201|COMP|25564-6|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C0945240|T201|COMP|25573-7|LNC|C peptide^15th specimen post XXX challenge|C peptide^15th specimen post XXX challenge
C0945241|T201|COMP|25574-5|LNC|C peptide^1st specimen post XXX challenge|C peptide^1st specimen post XXX challenge
C0945242|T201|COMP|25583-6|LNC|Calcium|Calcium
C0945243|T201|COMP|25586-9|LNC|Chicken droppings Ab.IgE.RAST class|Chicken droppings Ab.IgE.RAST class
C0945244|T201|COMP|25587-7|LNC|Chromogranin A|Chromogranin A
C0945245|T201|COMP|25595-0|LNC|Econazole|Econazole
C0945246|T201|COMP|25613-1|LNC|Periplaneta fuliginosa Ab.IgE|Periplaneta fuliginosa Ab.IgE
C0945248|T201|COMP|25633-9|LNC|Leishmania donovani Ab|Leishmania donovani Ab
C0945250|T201|COMP|25647-9|LNC|Follitropin^4th specimen post XXX challenge|Follitropin^4th specimen post XXX challenge
C0945251|T201|COMP|25654-5|LNC|Gastrin^1st specimen post XXX challenge|Gastrin^1st specimen post XXX challenge
C0945252|T201|COMP|25666-9|LNC|Glucose^2.5H post dose glucose|Glucose^2.5H post dose glucose
C0945253|T201|COMP|25678-4|LNC|Glucose^1.5H post dose glucose|Glucose^1.5H post dose glucose
C0945254|T201|COMP|25696-6|LNC|Insulin^7.5H post XXX challenge|Insulin^7.5H post XXX challenge
C0945255|T201|COMP|25699-0|LNC|Insulin^9th specimen post XXX challenge|Insulin^9th specimen post XXX challenge
C0945256|T201|COMP|25704-8|LNC|Ziziphus jujuba Ab.IgE.RAST class|Ziziphus jujuba Ab.IgE.RAST class
C0945257|T201|COMP|25712-1|LNC|Leptospira interrogans serovar Pomona Ab|Leptospira interrogans serovar Pomona Ab
C0945258|T201|COMP|25735-2|LNC|Prolactin^1H post 200 ug TRH IV|Prolactin^1H post 200 ug TRH IV
C0945259|T201|COMP|25746-9|LNC|Rheumatoid factor|Rheumatoid factor
C0945260|T201|COMP|25750-1|LNC|Rickettsia conorii Ab.IgM|Rickettsia conorii Ab.IgM
C0945261|T201|COMP|25755-0|LNC|Rotavirus Ab.IgM|Rotavirus Ab.IgM
C0945264|T201|COMP|25793-1|LNC|Thyroxine.free^4th specimen post XXX challenge|Thyroxine.free^4th specimen post XXX challenge
C0945266|T201|COMP|25812-9|LNC|Trimipramine+Nortrimipramine|Trimipramine+Nortrimipramine
C0945267|T201|COMP|25816-0|LNC|Vigabatrin|Vigabatrin
C0945268|T201|COMP|25817-8|LNC|Xylose^1.5H post dose xylose PO|Xylose^1.5H post dose xylose PO
C0945269|T201|COMP|25822-8|LNC|Staphylococcus aureus enterotoxin B Ab.IgE|Staphylococcus aureus enterotoxin B Ab.IgE
C0945271|T201|COMP|25833-5|LNC|Cerebroside sulfatase activator|Cerebroside sulfatase activator
C0945272|T201|COMP|25835-0|LNC|HIV 1 RNA|HIV 1 RNA
C0945273|T201|COMP|25863-2|LNC|Asparagine/Creatinine|Asparagine/Creatinine
C0945274|T201|COMP|25865-7|LNC|Aspartate/Creatinine|Aspartate/Creatinine
C0945275|T201|COMP|25866-5|LNC|Leptospira borgpetersenii serovar Sejroe Ab|Leptospira borgpetersenii serovar Sejroe Ab
C0945276|T201|COMP|25868-1|LNC|Beta alanine|Beta alanine
C0945277|T201|COMP|25876-4|LNC|Citrate|Citrate
C0945278|T201|COMP|25884-8|LNC|Cortisol.free|Cortisol.free
C0945279|T201|COMP|25889-7|LNC|Cysteate|Cysteate
C0945280|T201|COMP|25892-1|LNC|Cysteine|Cysteine
C0945281|T201|COMP|25900-2|LNC|D-Lactate^2nd specimen post exercise|D-Lactate^2nd specimen post exercise
C0945282|T201|COMP|25903-6|LNC|D-Lactate^5th specimen post exercise|D-Lactate^5th specimen post exercise
C0945283|T201|COMP|25925-9|LNC|Histamine/Creatinine|Histamine/Creatinine
C0945284|T201|COMP|25933-3|LNC|Hydroxylysine/Creatinine|Hydroxylysine/Creatinine
C0945285|T201|COMP|25936-6|LNC|Iodine|Iodine
C0945286|T201|COMP|25937-4|LNC|Iron|Iron
C0945287|T201|COMP|25938-2|LNC|Isoleucine|Isoleucine
C0945288|T201|COMP|25942-4|LNC|Leucine/Creatinine|Leucine/Creatinine
C0945289|T201|COMP|25946-5|LNC|Lutropin^4th specimen post XXX challenge|Lutropin^4th specimen post XXX challenge
C0945290|T201|COMP|25952-3|LNC|Lysine|Lysine
C0945291|T201|COMP|25956-4|LNC|Methionine|Methionine
C0945292|T201|COMP|25963-0|LNC|Norepinephrine|Norepinephrine
C0945293|T201|COMP|25990-3|LNC|Thyrotropin^30M post dose TRH IN|Thyrotropin^30M post dose TRH IN
C0945294|T201|COMP|25992-9|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C0945295|T201|COMP|25996-0|LNC|Tyrosine/Creatinine|Tyrosine/Creatinine
C0945296|T201|COMP|26007-5|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C0945297|T201|COMP|26011-7|LNC|Macroamylase/Amylase.total|Macroamylase/Amylase.total
C0945298|T201|COMP|26016-6|LNC|Cholesterol.in HDL 2|Cholesterol.in HDL 2
C0945299|T201|COMP|26018-2|LNC|Cladosporium cladosporioides Ab.IgG.RAST class|Cladosporium cladosporioides Ab.IgG.RAST class
C0945301|T201|COMP|26039-8|LNC|Norflunitrazepam|Norflunitrazepam
C0945302|T201|COMP|26053-9|LNC|N-methylhistamine|N-methylhistamine
C0945303|T201|COMP|26057-0|LNC|Pyridoxine^post pyridoxine PO|Pyridoxine^post pyridoxine PO
C0945304|T201|COMP|26062-0|LNC|European tick borne encephalitis virus Ab.IgG|European tick borne encephalitis virus Ab.IgG
C0945350|T201|COMP|26405-1|LNC|Aspergillus fumigatus Ab.IgG4|Aspergillus fumigatus Ab.IgG4
C0945351|T201|COMP|26414-3|LNC|Candida albicans Ab.IgG4.RAST class|Candida albicans Ab.IgG4.RAST class
C0945352|T201|COMP|26426-7|LNC|Lactalbumin alpha Ab.IgG4.RAST class|Lactalbumin alpha Ab.IgG4.RAST class
C0945353|T201|COMP|26429-1|LNC|Oryza sativa Ab.IgG4.RAST class|Oryza sativa Ab.IgG4.RAST class
C0945354|T201|COMP|26450-7|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0945355|T201|COMP|26455-6|LNC|Erythrocytes|Erythrocytes
C0945356|T201|COMP|26461-4|LNC|Erythrocytes.nucleated/100 erythrocytes|Erythrocytes.nucleated/100 erythrocytes
C0945357|T201|COMP|26464-8|LNC|Leukocytes|Leukocytes
C0945358|T201|COMP|26468-9|LNC|Leukocytes|Leukocytes
C0945359|T201|COMP|26471-3|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0945360|T201|COMP|26477-0|LNC|Lymphocytes.variant|Lymphocytes.variant
C0945361|T201|COMP|26504-1|LNC|Neutrophils|Neutrophils
C0945362|T201|COMP|26507-4|LNC|Neutrophils.band form|Neutrophils.band form
C0945363|T201|COMP|26512-4|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0945364|T201|COMP|26517-3|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0945365|T201|COMP|26522-3|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0945366|T201|COMP|26527-2|LNC|Cortisol.free^72H post dose corticotropin|Cortisol.free^72H post dose corticotropin
C0945367|T201|COMP|26533-0|LNC|Cortisol^56H post dose corticotropin|Cortisol^56H post dose corticotropin
C0945368|T201|COMP|26538-9|LNC|Glucose^3.5H post dose glucose|Glucose^3.5H post dose glucose
C0945369|T201|COMP|26553-8|LNC|Glucose^1.5H post dose glucose|Glucose^1.5H post dose glucose
C0945370|T201|COMP|26556-1|LNC|Cells.CD103/100 cells|Cells.CD103/100 cells
C0945371|T201|COMP|26571-0|LNC|Cells.CD16|Cells.CD16
C0945372|T201|COMP|26580-1|LNC|Carnosine/Creatinine|Carnosine/Creatinine
C0945373|T201|COMP|26586-8|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0945374|T201|COMP|26589-2|LNC|Beta alanine|Beta alanine
C0945375|T201|COMP|26592-6|LNC|Cystathionine|Cystathionine
C0945376|T201|COMP|26593-4|LNC|Ethanolamine|Ethanolamine
C0945377|T201|COMP|26597-5|LNC|Phosphoethanolamine|Phosphoethanolamine
C0945378|T201|COMP|26618-9|LNC|Trypanosoma brucei rhodesiense Ab|Trypanosoma brucei rhodesiense Ab
C0945379|T201|COMP|26621-3|LNC|Legionella sp Ag|Legionella sp Ag
C0945380|T201|COMP|26635-3|LNC|Legionella micdadei Ab|Legionella micdadei Ab
C0945381|T201|COMP|26643-7|LNC|Clostridium tetani toxoid Ab|Clostridium tetani toxoid Ab
C0945382|T201|COMP|26648-6|LNC|Sindbis virus Ab|Sindbis virus Ab
C0945383|T201|COMP|26651-0|LNC|Rhizopus arrhizus Ab|Rhizopus arrhizus Ab
C0945384|T201|COMP|26652-8|LNC|Banzi virus Ab|Banzi virus Ab
C0945385|T201|COMP|26655-1|LNC|Entamoeba sp Ab|Entamoeba sp Ab
C0945386|T201|COMP|26656-9|LNC|HTLV II Ab|HTLV II Ab
C0945387|T201|COMP|26660-1|LNC|Toxocara sp Ab|Toxocara sp Ab
C0945388|T201|COMP|26664-3|LNC|Chlamydia trachomatis E Ab|Chlamydia trachomatis E Ab
C0945389|T201|COMP|26677-5|LNC|Bartonella quintana Ab|Bartonella quintana Ab
C0945390|T201|COMP|26680-9|LNC|Aspartate|Aspartate
C0945391|T201|COMP|26702-1|LNC|Clostridioides difficile Ab.IgG|Clostridioides difficile Ab.IgG
C0945392|T201|COMP|26705-4|LNC|Epstein Barr virus nuclear Ab.IgM|Epstein Barr virus nuclear Ab.IgM
C0945393|T201|COMP|26707-0|LNC|Aluminum|Aluminum
C0945394|T201|COMP|26709-6|LNC|Xylose^5th specimen post XXX challenge|Xylose^5th specimen post XXX challenge
C0945395|T201|COMP|26711-2|LNC|Phendimetrazine|Phendimetrazine
C0945396|T201|COMP|26715-3|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C0945397|T201|COMP|26724-5|LNC|Sarcosine|Sarcosine
C0945398|T201|COMP|26728-6|LNC|Cells.CD38|Cells.CD38
C0945399|T201|COMP|26749-2|LNC|Urea nitrogen^2nd specimen|Urea nitrogen^2nd specimen
C0945400|T201|COMP|26760-9|LNC|Cannabinoids|Cannabinoids
C0945401|T201|COMP|26769-0|LNC|Endothelin|Endothelin
C0945402|T201|COMP|26772-4|LNC|Mephentermine|Mephentermine
C0945403|T201|COMP|26779-9|LNC|Glucose^1.5H post dose lactose PO|Glucose^1.5H post dose lactose PO
C0945404|T201|COMP|26782-3|LNC|Glucose^4H post dose lactose PO|Glucose^4H post dose lactose PO
C0945405|T201|COMP|26786-4|LNC|Mephentermine|Mephentermine
C0945406|T201|COMP|26790-6|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C0945407|T201|COMP|26794-8|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C0945408|T201|COMP|26812-8|LNC|Xylose^3rd specimen post XXX challenge|Xylose^3rd specimen post XXX challenge
C0945409|T201|COMP|26815-1|LNC|Cocaethylene|Cocaethylene
C0945410|T201|COMP|26828-4|LNC|Cortisol|Cortisol
C0945411|T201|COMP|26832-6|LNC|Aconitate|Aconitate
C0945412|T201|COMP|26836-7|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C0945413|T201|COMP|26840-9|LNC|Nordiazepam|Nordiazepam
C0945414|T201|COMP|26844-1|LNC|Methionine|Methionine
C0945415|T201|COMP|26846-6|LNC|Perphenazine|Perphenazine
C0945416|T201|COMP|26848-2|LNC|Interleukin 10|Interleukin 10
C0945417|T201|COMP|26852-4|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C0945418|T201|COMP|26860-7|LNC|Morphine|Morphine
C0945420|T201|COMP|26891-2|LNC|Nordiazepam|Nordiazepam
C0945421|T201|COMP|26895-3|LNC|Amphetamines|Amphetamines
C0945422|T201|COMP|26899-5|LNC|Midazolam|Midazolam
C0945423|T201|COMP|26901-9|LNC|Flurazepam|Flurazepam
C0945424|T201|COMP|26906-8|LNC|Mephobarbital|Mephobarbital
C0945425|T201|COMP|26914-2|LNC|Estazolam|Estazolam
C0945426|T201|COMP|26918-3|LNC|PENTobarbital|PENTobarbital
C0945427|T201|COMP|26921-7|LNC|Cells.CD2+CD26+|Cells.CD2+CD26+
C0945428|T201|COMP|26924-1|LNC|Cancer Ag 19-9|Cancer Ag 19-9
C0945429|T201|COMP|26927-4|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C0945431|T201|COMP|26943-1|LNC|11-Ketoandrosterone|11-Ketoandrosterone
C0945432|T201|COMP|26964-7|LNC|Cystathionine|Cystathionine
C0945433|T201|COMP|26968-8|LNC|Beta alanine|Beta alanine
C0945434|T201|COMP|26971-2|LNC|Smooth muscle Ab|Smooth muscle Ab
C0945435|T201|COMP|26973-8|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C0945436|T201|COMP|26974-6|LNC|Delta aminolevulinate|Delta aminolevulinate
C0945437|T201|COMP|26976-1|LNC|Hydroxytriazolam|Hydroxytriazolam
C0945438|T201|COMP|26980-3|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C0945439|T201|COMP|26985-2|LNC|Arginine|Arginine
C0945440|T201|COMP|26989-4|LNC|Trypanosoma cruzi Ab.IgM|Trypanosoma cruzi Ab.IgM
C0945441|T201|COMP|27022-3|LNC|Para aminophenol/Creatinine|Para aminophenol/Creatinine
C0945442|T201|COMP|27024-9|LNC|Cannabinoids|Cannabinoids
C0945443|T201|COMP|27028-0|LNC|Ketones^2H post XXX challenge|Ketones^2H post XXX challenge
C0945444|T201|COMP|27037-1|LNC|Calcium/Creatinine|Calcium/Creatinine
C0945445|T201|COMP|27041-3|LNC|Norpropoxyphene|Norpropoxyphene
C0945446|T201|COMP|27045-4|LNC|Microscopic exam|Microscopic exam
C0945447|T201|COMP|27051-2|LNC|PHENobarbital|PHENobarbital
C0945448|T201|COMP|27053-8|LNC|Morphine|Morphine
C0945449|T201|COMP|27057-9|LNC|Serotonin|Serotonin
C0945450|T201|COMP|27074-4|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C0945451|T201|COMP|27093-4|LNC|Leptospira sp Ab.IgG|Leptospira sp Ab.IgG
C0945452|T201|COMP|27097-5|LNC|2-Methylbutyrylglycine/Creatinine|2-Methylbutyrylglycine/Creatinine
C0945453|T201|COMP|27098-3|LNC|Methionine|Methionine
C0945454|T201|COMP|27101-5|LNC|Phenmetrazine|Phenmetrazine
C0945455|T201|COMP|27105-6|LNC|Amphetamines|Amphetamines
C0945456|T201|COMP|27107-2|LNC|Lysine|Lysine
C0945457|T201|COMP|27113-0|LNC|Streptococcus pneumoniae 8 Ab.IgG|Streptococcus pneumoniae 8 Ab.IgG
C0945459|T201|COMP|27123-9|LNC|Phosphate|Phosphate
C0945460|T201|COMP|27132-0|LNC|Acetoacetate|Acetoacetate
C0945461|T201|COMP|27134-6|LNC|Argininosuccinate|Argininosuccinate
C0945462|T201|COMP|27155-1|LNC|Streptococcus pneumoniae 6 Ab^2nd specimen|Streptococcus pneumoniae 6 Ab^2nd specimen
C0945463|T201|COMP|27158-5|LNC|Streptococcus pneumoniae 14 Ab^1st specimen|Streptococcus pneumoniae 14 Ab^1st specimen
C0945464|T201|COMP|27160-1|LNC|Hydrastine|Hydrastine
C0945465|T201|COMP|27164-3|LNC|acetoHEXAMIDE|acetoHEXAMIDE
C0945466|T201|COMP|27165-0|LNC|Hexobarbital|Hexobarbital
C0945467|T201|COMP|27169-2|LNC|Butyrate|Butyrate
C0945468|T201|COMP|27172-6|LNC|Calcium|Calcium
C0945469|T201|COMP|27177-5|LNC|Herpes virus 7 Ab.IgM|Herpes virus 7 Ab.IgM
C0945470|T201|COMP|27180-9|LNC|Bisacodyl|Bisacodyl
C0945471|T201|COMP|27185-8|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C0945472|T201|COMP|27190-8|LNC|Propoxyphene|Propoxyphene
C0945473|T201|COMP|27209-6|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C0945474|T201|COMP|27221-1|LNC|Norepinephrine|Norepinephrine
C0945475|T201|COMP|27225-2|LNC|Estriol|Estriol
C0945476|T201|COMP|27229-4|LNC|Streptococcus pneumoniae 14 Ab.IgG|Streptococcus pneumoniae 14 Ab.IgG
C0945477|T201|COMP|27234-4|LNC|Phentermine|Phentermine
C0945478|T201|COMP|27238-5|LNC|Oxazepam|Oxazepam
C0945479|T201|COMP|27241-9|LNC|Mephobarbital|Mephobarbital
C0945480|T201|COMP|27246-8|LNC|Butalbital|Butalbital
C0945481|T201|COMP|27248-4|LNC|Benzoylecgonine|Benzoylecgonine
C0945482|T201|COMP|27249-2|LNC|Temazepam|Temazepam
C0945483|T201|COMP|27264-1|LNC|Aluminum|Aluminum
C0945484|T201|COMP|27285-6|LNC|Estazolam|Estazolam
C0945485|T201|COMP|27289-8|LNC|Methamphetamine|Methamphetamine
C0945486|T201|COMP|27292-2|LNC|Ornithine|Ornithine
C0945487|T201|COMP|27293-0|LNC|oxyCODONE.free|oxyCODONE.free
C0945488|T201|COMP|27297-1|LNC|Leukocyte esterase|Leukocyte esterase
C0945489|T201|COMP|27299-7|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C0945490|T201|COMP|27300-3|LNC|Mephentermine|Mephentermine
C0945491|T201|COMP|27308-6|LNC|PENTobarbital|PENTobarbital
C0945492|T201|COMP|27320-1|LNC|Parietal cell Ab|Parietal cell Ab
C0945493|T201|COMP|27325-0|LNC|Glycine|Glycine
C0945494|T201|COMP|27354-0|LNC|Toxoplasma gondii Ab.IgE|Toxoplasma gondii Ab.IgE
C0945495|T201|COMP|27359-9|LNC|Somatotropin^15th specimen post XXX challenge|Somatotropin^15th specimen post XXX challenge
C0945496|T201|COMP|27364-9|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C0945497|T201|COMP|27369-8|LNC|Somatotropin^2.5H post XXX challenge|Somatotropin^2.5H post XXX challenge
C0945499|T201|COMP|27381-3|LNC|Alloisoleucine|Alloisoleucine
C0945500|T201|COMP|27382-1|LNC|Porphobilinogen|Porphobilinogen
C0945501|T201|COMP|27385-4|LNC|Somatotropin^18th specimen post XXX challenge|Somatotropin^18th specimen post XXX challenge
C0945502|T201|COMP|27403-5|LNC|Gamma glutamyl transferase|Gamma glutamyl transferase
C0945503|T201|COMP|27412-6|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C0945504|T201|COMP|27419-1|LNC|Sodium|Sodium
C0945506|T201|COMP|27432-4|LNC|Glucose^8th specimen post XXX challenge|Glucose^8th specimen post XXX challenge
C0945507|T201|COMP|27435-7|LNC|Streptococcus pneumoniae 19 Ab.IgG^1st specimen|Streptococcus pneumoniae 19 Ab.IgG^1st specimen
C0945508|T201|COMP|27438-1|LNC|Protein C Ag/Coagulation factor VII Ag|Protein C Ag/Coagulation factor VII Ag
C0945509|T201|COMP|27442-3|LNC|Phenylpropanolamine|Phenylpropanolamine
C0945541|T201|COMP|27822-6|LNC|Protein S actual/Normal|Protein S actual/Normal
C0945542|T201|COMP|27827-5|LNC|Insulin^30M post XXX challenge|Insulin^30M post XXX challenge
C0945543|T201|COMP|27829-1|LNC|Somatotropin^8th specimen post XXX challenge|Somatotropin^8th specimen post XXX challenge
C0945544|T201|COMP|27831-7|LNC|Immune complex|Immune complex
C0945545|T201|COMP|27837-4|LNC|Somatotropin^13th specimen post XXX challenge|Somatotropin^13th specimen post XXX challenge
C0945546|T201|COMP|27847-3|LNC|Somatotropin^25th specimen post XXX challenge|Somatotropin^25th specimen post XXX challenge
C0945547|T201|COMP|27875-4|LNC|Insulin^6th specimen post XXX challenge|Insulin^6th specimen post XXX challenge
C0945548|T201|COMP|27880-4|LNC|Follitropin^6th specimen post XXX challenge|Follitropin^6th specimen post XXX challenge
C0945549|T201|COMP|27884-6|LNC|Lutropin^40M post XXX challenge|Lutropin^40M post XXX challenge
C0945550|T201|COMP|27890-3|LNC|Somatotropin^5th specimen post XXX challenge|Somatotropin^5th specimen post XXX challenge
C0945552|T201|COMP|27908-3|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C0945553|T201|COMP|27909-1|LNC|Calcium^1st specimen post XXX challenge|Calcium^1st specimen post XXX challenge
C0945554|T201|COMP|27935-6|LNC|Calcium^4th specimen post XXX challenge|Calcium^4th specimen post XXX challenge
C0945555|T201|COMP|27937-2|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C0945556|T201|COMP|27945-5|LNC|Coxiella burnetii phase 2 Ab|Coxiella burnetii phase 2 Ab
C0945557|T201|COMP|27946-3|LNC|Lactate^1H post XXX challenge|Lactate^1H post XXX challenge
C0945558|T201|COMP|27954-7|LNC|Coxsackievirus B6 RNA|Coxsackievirus B6 RNA
C0945559|T201|COMP|27977-8|LNC|Norepinephrine/Creatinine|Norepinephrine/Creatinine
C0945560|T201|COMP|27980-2|LNC|Thyroxine binding globulin|Thyroxine binding globulin
C0945561|T201|COMP|27994-3|LNC|Ehrlichia chaffeensis DNA|Ehrlichia chaffeensis DNA
C0945562|T201|COMP|27999-2|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C0945563|T201|COMP|28001-6|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C0945564|T201|COMP|28007-3|LNC|Urobilinogen|Urobilinogen
C0945568|T201|COMP|28041-2|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C0945569|T201|COMP|28044-6|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C0945570|T201|COMP|28051-1|LNC|1,3,5-Trichlorobenzene|1,3,5-Trichlorobenzene
C0945571|T201|COMP|28056-0|LNC|Borrelia burgdorferi 28kD Ab.IgG|Borrelia burgdorferi 28kD Ab.IgG
C0945572|T201|COMP|28061-0|LNC|Naloxone|Naloxone
C0945573|T201|COMP|28073-5|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C0945574|T201|COMP|28075-0|LNC|Sildenafil citrate|Sildenafil citrate
C0945575|T201|COMP|28078-4|LNC|Bladder tumor Ag|Bladder tumor Ag
C0945625|T201|COMP|28539-5|LNC|Erythrocyte mean corpuscular hemoglobin|Erythrocyte mean corpuscular hemoglobin
C0945626|T201|COMP|28544-5|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C0945627|T201|COMP|28554-4|LNC|Triglyceride|Triglyceride
C0945630|T201|COMP|28589-0|LNC|Carnitine esters/Creatinine|Carnitine esters/Creatinine
C0945631|T201|COMP|28598-1|LNC|Alpha aminoadipate/Creatinine|Alpha aminoadipate/Creatinine
C0945632|T201|COMP|28601-3|LNC|Hydroxyproline/Creatinine|Hydroxyproline/Creatinine
C0945633|T201|COMP|28606-2|LNC|1-Methylhistidine/Creatinine|1-Methylhistidine/Creatinine
C0945634|T201|COMP|28610-4|LNC|Sarcosine/Creatinine|Sarcosine/Creatinine
C0945637|T201|COMP|28643-5|LNC|Oxygen saturation|Oxygen saturation
C0945639|T201|COMP|28649-2|LNC|Oxygen|Oxygen
C0945642|T201|COMP|28660-9|LNC|Plasminogen actual/Normal|Plasminogen actual/Normal
C0945703|T201|COMP|29115-3|LNC|Delavirdine|Delavirdine
C0945704|T201|COMP|29116-1|LNC|Didanosine|Didanosine
C0945705|T201|COMP|29118-7|LNC|Indinavir|Indinavir
C0945706|T201|COMP|29123-7|LNC|Saquinavir|Saquinavir
C0945709|T201|COMP|29151-8|LNC|Somatotropin^4H post XXX challenge|Somatotropin^4H post XXX challenge
C0945718|T201|COMP|29229-2|LNC|Valproate|Valproate
C0945719|T201|COMP|29230-0|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C0945720|T201|COMP|29232-6|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C0945721|T201|COMP|29237-5|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C0945722|T201|COMP|29241-7|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0945723|T201|COMP|29253-2|LNC|Alpha-1-Fetoprotein^^adjusted|Alpha-1-Fetoprotein^^adjusted
C0945726|T201|COMP|29294-6|LNC|Methadone|Methadone
C0945732|T201|COMP|29311-8|LNC|Neisseria gonorrhoeae Ag|Neisseria gonorrhoeae Ag
C0945733|T201|COMP|29318-3|LNC|Streptococcus pneumoniae group B Ag|Streptococcus pneumoniae group B Ag
C0945734|T201|COMP|29323-3|LNC|Cocaine|Cocaine
C0945735|T201|COMP|29328-2|LNC|Xylose^2.5H post dose xylose PO|Xylose^2.5H post dose xylose PO
C0945736|T201|COMP|29357-1|LNC|Cyanide|Cyanide
C0945737|T201|COMP|29358-9|LNC|Cortisol^pre XXX challenge|Cortisol^pre XXX challenge
C0945738|T201|COMP|29360-5|LNC|Streptococcus pneumoniae group B Ag|Streptococcus pneumoniae group B Ag
C0945739|T201|COMP|29362-1|LNC|Streptococcus pneumoniae group B Ag|Streptococcus pneumoniae group B Ag
C0945740|T201|COMP|29366-2|LNC|Parainfluenza virus 1 Ab|Parainfluenza virus 1 Ab
C0945741|T201|COMP|29370-4|LNC|cloZAPine^trough|cloZAPine^trough
C0945742|T201|COMP|29374-6|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0945743|T201|COMP|29383-7|LNC|Warfarin|Warfarin
C0945744|T201|COMP|29387-8|LNC|Norpropoxyphene|Norpropoxyphene
C0945745|T201|COMP|29392-8|LNC|Gastrin^1H post XXX challenge|Gastrin^1H post XXX challenge
C0945746|T201|COMP|29412-4|LNC|Glucose^6H post XXX challenge|Glucose^6H post XXX challenge
C0945758|T201|COMP|29494-2|LNC|Demeclocycline|Demeclocycline
C0945759|T201|COMP|29525-3|LNC|Aconitate/Creatinine|Aconitate/Creatinine
C0945760|T201|COMP|29528-7|LNC|Hippurate/Creatinine|Hippurate/Creatinine
C0945761|T201|COMP|29530-3|LNC|Amphetamines|Amphetamines
C0945762|T201|COMP|29534-5|LNC|Anguilla anguilla Ab.IgE.RAST class|Anguilla anguilla Ab.IgE.RAST class
C0945763|T201|COMP|29539-4|LNC|HIV 1 RNA|HIV 1 RNA
C0945767|T201|COMP|29578-2|LNC|Viral susceptibility panel|Viral susceptibility panel
C0945768|T201|COMP|29583-2|LNC|Differential panel|Differential panel
C0945769|T201|COMP|29590-7|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C0945770|T201|COMP|29595-6|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0945771|T201|COMP|29603-8|LNC|CD5 Ag|CD5 Ag
C0945772|T201|COMP|29608-7|LNC|Phentermine|Phentermine
C0945773|T201|COMP|29610-3|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C0945774|T201|COMP|29612-9|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C0945775|T201|COMP|29616-0|LNC|Stachybotrys chartarum Ab.IgE|Stachybotrys chartarum Ab.IgE
C0945776|T201|COMP|29617-8|LNC|CD23 Ag|CD23 Ag
C0945777|T201|COMP|29635-0|LNC|Albuterol|Albuterol
C0945778|T201|COMP|29637-6|LNC|Time last dose|Time last dose
C0945779|T201|COMP|29650-9|LNC|Rickettsia honei Ab|Rickettsia honei Ab
C0945780|T201|COMP|29655-8|LNC|Oxazepam|Oxazepam
C0945781|T201|COMP|29659-0|LNC|Bordetella pertussis Ab.IgG|Bordetella pertussis Ab.IgG
C0945782|T201|COMP|29664-0|LNC|Chlamydia sp Ab.IgA|Chlamydia sp Ab.IgA
C0945783|T201|COMP|29666-5|LNC|Echovirus+Coxsackievirus Ab.IgA|Echovirus+Coxsackievirus Ab.IgA
C0945784|T201|COMP|29668-1|LNC|Rickettsia australis Ab|Rickettsia australis Ab
C0945785|T201|COMP|29672-3|LNC|Bordetella pertussis Ab.IgA|Bordetella pertussis Ab.IgA
C0945786|T201|COMP|29677-2|LNC|Chlamydia sp Ab.IgA|Chlamydia sp Ab.IgA
C0945787|T201|COMP|29681-4|LNC|Rickettsia akari Ab|Rickettsia akari Ab
C0945788|T201|COMP|29710-1|LNC|Rickettsia prowazekii Ab|Rickettsia prowazekii Ab
C0945789|T201|COMP|29713-5|LNC|Orientia tsutsugamushi Gilliam Ab|Orientia tsutsugamushi Gilliam Ab
C0945790|T201|COMP|29719-2|LNC|Orientia tsutsugamushi Litchfield Ab|Orientia tsutsugamushi Litchfield Ab
C0945791|T201|COMP|29720-0|LNC|Orientia tsutsugamushi Litchfield Ab|Orientia tsutsugamushi Litchfield Ab
C0945792|T201|COMP|29724-2|LNC|Leptospira interrogans serovar Celledoni Ab|Leptospira interrogans serovar Celledoni Ab
C0945793|T201|COMP|29733-3|LNC|Leptospira interrogans serovar Kremastos Ab|Leptospira interrogans serovar Kremastos Ab
C0945794|T201|COMP|29739-0|LNC|Leptospira interrogans serovar Kremastos Ab|Leptospira interrogans serovar Kremastos Ab
C0945795|T201|COMP|29747-3|LNC|Tocopherols|Tocopherols
C0947214|T201|COMP|25366-6|LNC|cefOXitin|cefOXitin
C0947215|T201|COMP|25446-6|LNC|IgM|IgM
C0947216|T201|COMP|25690-9|LNC|Insulin^15th specimen post XXX challenge|Insulin^15th specimen post XXX challenge
C0947217|T201|COMP|25709-7|LNC|Leptospira interrogans serovar Canicola Ab|Leptospira interrogans serovar Canicola Ab
C0947218|T201|COMP|25872-3|LNC|C peptide|C peptide
C0947219|T201|COMP|26002-6|LNC|Valine/Creatinine|Valine/Creatinine
C0947220|T201|COMP|26532-2|LNC|Cortisol^48H post dose corticotropin|Cortisol^48H post dose corticotropin
C0947221|T201|COMP|26576-9|LNC|Anserine/Creatinine|Anserine/Creatinine
C0947222|T201|COMP|26584-3|LNC|1-Methylhistidine|1-Methylhistidine
C0947223|T201|COMP|26765-8|LNC|Antimony|Antimony
C0947224|T201|COMP|26777-3|LNC|Glucose^30M post dose lactose PO|Glucose^30M post dose lactose PO
C0947225|T201|COMP|26781-5|LNC|Glucose^3H post dose lactose PO|Glucose^3H post dose lactose PO
C0947226|T201|COMP|26857-3|LNC|Mephentermine|Mephentermine
C0947227|T201|COMP|26926-6|LNC|Ganglioside GD1b Ab|Ganglioside GD1b Ab
C0947228|T201|COMP|26993-6|LNC|Benzfetamine|Benzfetamine
C0947229|T201|COMP|27033-0|LNC|Proline|Proline
C0947230|T201|COMP|27304-5|LNC|Lysine|Lysine
C0947231|T201|COMP|27312-8|LNC|HYDROcodone.free|HYDROcodone.free
C0947232|T201|COMP|27317-7|LNC|Asparagine|Asparagine
C0947233|T201|COMP|27373-0|LNC|Calcium|Calcium
C0947234|T201|COMP|27423-3|LNC|1,4-Dioxane|1,4-Dioxane
C0947235|T201|COMP|27885-3|LNC|Lutropin^1.5H post XXX challenge|Lutropin^1.5H post XXX challenge
C0947236|T201|COMP|27930-7|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0947240|T201|COMP|28549-4|LNC|Yersinia sp identified|Yersinia sp identified
C0947241|T201|COMP|28593-2|LNC|Gamma aminobutyrate/Creatinine|Gamma aminobutyrate/Creatinine
C0947249|T201|COMP|29246-6|LNC|Lactate|Lactate
C0947250|T201|COMP|29663-2|LNC|Dengue virus Ab.IgM|Dengue virus Ab.IgM
C0947251|T201|COMP|29767-1|LNC|Bilirubin|Bilirubin
C0947252|T201|COMP|25748-5|LNC|Ribosomal Ab|Ribosomal Ab
C0947257|T201|COMP|26459-8|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C0947258|T201|COMP|27355-7|LNC|Lipoprotein.pre-beta|Lipoprotein.pre-beta
C0947259|T201|COMP|27810-1|LNC|Plasmin inhibitor actual/Normal|Plasmin inhibitor actual/Normal
C0947260|T201|COMP|28008-1|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C0947265|T201|COMP|29236-7|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C0947266|T201|COMP|29329-0|LNC|Glucose^3.5H post XXX challenge|Glucose^3.5H post XXX challenge
C0947267|T201|COMP|29497-5|LNC|Platelet associated Ab.IgG|Platelet associated Ab.IgG
C0947495|T201|COMP|14251-3|LNC|Mitochondria M2 Ab.IgG|Mitochondria M2 Ab.IgG
C0947496|T201|COMP|27864-8|LNC|Follitropin^9th specimen post XXX challenge|Follitropin^9th specimen post XXX challenge
C0947498|T201|COMP|27017-3|LNC|Allyl alcohol|Allyl alcohol
C0947553|T201|COMP|29688-9|LNC|Orientia tsutsugamushi Karp Ab|Orientia tsutsugamushi Karp Ab
C1113710|T201|COMP|29770-5|LNC|Karyotype|Karyotype
C1113711|T201|COMP|29771-3|LNC|Hemoglobin.gastrointestinal.lower|Hemoglobin.gastrointestinal.lower
C1113712|T201|COMP|29772-1|LNC|Coxiella burnetii phase 2 Ab|Coxiella burnetii phase 2 Ab
C1113713|T201|COMP|29773-9|LNC|Coxiella burnetii phase 2 Ab.IgM|Coxiella burnetii phase 2 Ab.IgM
C1113714|T201|COMP|29774-7|LNC|Coxiella burnetii phase 1 Ab|Coxiella burnetii phase 1 Ab
C1113715|T201|COMP|29775-4|LNC|Insulin-like growth factor-I|Insulin-like growth factor-I
C1113717|T201|COMP|29777-0|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C1113718|T201|COMP|29778-8|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1113719|T201|COMP|29779-6|LNC|West Nile virus Ab|West Nile virus Ab
C1113720|T201|COMP|29780-4|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1113721|T201|COMP|29781-2|LNC|West Nile virus Ab|West Nile virus Ab
C1113722|T201|COMP|29783-8|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C1113723|T201|COMP|29785-3|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C1113724|T201|COMP|29786-1|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113725|T201|COMP|29787-9|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113726|T201|COMP|29789-5|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C1113727|T201|COMP|29790-3|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C1113728|T201|COMP|29791-1|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1113729|T201|COMP|29792-9|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1113730|T201|COMP|29794-5|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1113731|T201|COMP|29795-2|LNC|Trivittatus virus Ab|Trivittatus virus Ab
C1113732|T201|COMP|29796-0|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C1113733|T201|COMP|29797-8|LNC|Highlands J virus Ab|Highlands J virus Ab
C1113734|T201|COMP|29799-4|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113735|T201|COMP|29800-0|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113736|T201|COMP|29801-8|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C1113737|T201|COMP|29803-4|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C1113738|T201|COMP|29804-2|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1113739|T201|COMP|29805-9|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1113740|T201|COMP|29806-7|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1113741|T201|COMP|29807-5|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1113742|T201|COMP|29808-3|LNC|Trivittatus virus Ab|Trivittatus virus Ab
C1113743|T201|COMP|29809-1|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C1113744|T201|COMP|29810-9|LNC|Highlands J virus Ab|Highlands J virus Ab
C1113745|T201|COMP|29811-7|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C1113746|T201|COMP|29812-5|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113747|T201|COMP|29813-3|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113748|T201|COMP|29814-1|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C1113749|T201|COMP|29816-6|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C1113750|T201|COMP|29817-4|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1113751|T201|COMP|29818-2|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1113752|T201|COMP|29819-0|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1113753|T201|COMP|29820-8|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1113754|T201|COMP|29821-6|LNC|Trivittatus virus Ab|Trivittatus virus Ab
C1113755|T201|COMP|29822-4|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C1113756|T201|COMP|29823-2|LNC|Highlands J virus Ab|Highlands J virus Ab
C1113757|T201|COMP|29824-0|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C1113758|T201|COMP|29825-7|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113759|T201|COMP|29826-5|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113760|T201|COMP|29827-3|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C1113761|T201|COMP|29828-1|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C1113762|T201|COMP|29829-9|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C1113763|T201|COMP|29830-7|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1113764|T201|COMP|29831-5|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1113765|T201|COMP|29832-3|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1113766|T201|COMP|29833-1|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1113767|T201|COMP|29834-9|LNC|Trivittatus virus Ab|Trivittatus virus Ab
C1113768|T201|COMP|29835-6|LNC|Highlands J virus Ab|Highlands J virus Ab
C1113769|T201|COMP|29836-4|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C1113770|T201|COMP|29838-0|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113771|T201|COMP|29839-8|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C1113772|T201|COMP|29840-6|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C1113773|T201|COMP|29842-2|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1113774|T201|COMP|29843-0|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1113775|T201|COMP|29844-8|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1113776|T201|COMP|29847-1|LNC|Highlands J virus Ab|Highlands J virus Ab
C1113777|T201|COMP|29848-9|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C1113778|T201|COMP|29849-7|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1113779|T201|COMP|29851-3|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C1113780|T201|COMP|29852-1|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C1113781|T201|COMP|29853-9|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C1113782|T201|COMP|29854-7|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1113783|T201|COMP|29856-2|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1113784|T201|COMP|29857-0|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1113785|T201|COMP|29858-8|LNC|Alpha hydroxybutyrate/Creatinine|Alpha hydroxybutyrate/Creatinine
C1113786|T201|COMP|29859-6|LNC|Adipate/Creatinine|Adipate/Creatinine
C1113787|T201|COMP|29860-4|LNC|Cardiolipin Ab|Cardiolipin Ab
C1113788|T201|COMP|29861-2|LNC|Levisticum officinale Ab.IgE.RAST class|Levisticum officinale Ab.IgE.RAST class
C1113789|T201|COMP|29862-0|LNC|Diospyros kaki Ab.IgE.RAST class|Diospyros kaki Ab.IgE.RAST class
C1113790|T201|COMP|29864-6|LNC|2-Oxo,3-Methylvalerate|2-Oxo,3-Methylvalerate
C1113791|T201|COMP|29865-3|LNC|2-Oxoisocaproate|2-Oxoisocaproate
C1113792|T201|COMP|29866-1|LNC|2-Oxoisovalerate|2-Oxoisovalerate
C1113793|T201|COMP|29867-9|LNC|3-Hydroxy,3-Methylglutarate|3-Hydroxy,3-Methylglutarate
C1113794|T201|COMP|29868-7|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C1113795|T201|COMP|29869-5|LNC|4-Hydroxycyclohexylacetate|4-Hydroxycyclohexylacetate
C1113796|T201|COMP|29870-3|LNC|4-Hydroxyphenyllactate|4-Hydroxyphenyllactate
C1113797|T201|COMP|29871-1|LNC|4-Hydroxyphenylpyruvate|4-Hydroxyphenylpyruvate
C1113798|T201|COMP|29872-9|LNC|5-Oxoproline|5-Oxoproline
C1113799|T201|COMP|29873-7|LNC|Isobutyrylglycine|Isobutyrylglycine
C1113800|T201|COMP|29874-5|LNC|Isovalerylglycine|Isovalerylglycine
C1113801|T201|COMP|29875-2|LNC|Lactate|Lactate
C1113802|T201|COMP|29876-0|LNC|2-Methylcitrate|2-Methylcitrate
C1113803|T201|COMP|29877-8|LNC|Methylmalonate|Methylmalonate
C1113804|T201|COMP|29878-6|LNC|Argininosuccinate/Creatinine|Argininosuccinate/Creatinine
C1113805|T201|COMP|29879-4|LNC|Dehydroepiandrosterone/Creatinine|Dehydroepiandrosterone/Creatinine
C1113806|T201|COMP|29880-2|LNC|2-Hydroxy-3-Methylvalerate|2-Hydroxy-3-Methylvalerate
C1113807|T201|COMP|29881-0|LNC|2-Hydroxyglutarate|2-Hydroxyglutarate
C1113808|T201|COMP|29882-8|LNC|2-Hydroxyisovalerate|2-Hydroxyisovalerate
C1113809|T201|COMP|29883-6|LNC|2-Hydroxyphenylacetate|2-Hydroxyphenylacetate
C1113810|T201|COMP|29884-4|LNC|2-Methylbutyrylglycine|2-Methylbutyrylglycine
C1113811|T201|COMP|29885-1|LNC|Actinobacillus sp identified|Actinobacillus sp identified
C1113812|T201|COMP|29886-9|LNC|Encephalomyocarditis virus Ab|Encephalomyocarditis virus Ab
C1113813|T201|COMP|29887-7|LNC|Pasteurella multocida type|Pasteurella multocida type
C1113814|T201|COMP|29889-3|LNC|Encephalomyocarditis virus Ab|Encephalomyocarditis virus Ab
C1113815|T201|COMP|29890-1|LNC|Pseudorabies virus.G1 gene deletion Ab|Pseudorabies virus.G1 gene deletion Ab
C1113816|T201|COMP|29891-9|LNC|Carbon dioxide^post dose urea|Carbon dioxide^post dose urea
C1113817|T201|COMP|29892-7|LNC|Carbon dioxide^post dose urea|Carbon dioxide^post dose urea
C1113818|T201|COMP|29893-5|LNC|HIV 1 Ab|HIV 1 Ab
C1113819|T201|COMP|29894-3|LNC|Phosphorus|Phosphorus
C1113820|T201|COMP|29895-0|LNC|Phosphorus|Phosphorus
C1113821|T201|COMP|29896-8|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1113822|T201|COMP|29897-6|LNC|Styrene|Styrene
C1113823|T201|COMP|29898-4|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C1113824|T201|COMP|29899-2|LNC|Gamma globulin|Gamma globulin
C1113825|T201|COMP|29900-8|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1113826|T201|COMP|29901-6|LNC|HTLV I+II Ab|HTLV I+II Ab
C1113827|T201|COMP|29902-4|LNC|Chlorobenzene|Chlorobenzene
C1113828|T201|COMP|29904-0|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1113829|T201|COMP|29905-7|LNC|Entamoeba histolytica Ag|Entamoeba histolytica Ag
C1113830|T201|COMP|29906-5|LNC|Haemophilus influenzae A DNA|Haemophilus influenzae A DNA
C1113831|T201|COMP|29907-3|LNC|Haemophilus influenzae B DNA|Haemophilus influenzae B DNA
C1113832|T201|COMP|29909-9|LNC|Parainfluenza virus 2 RNA|Parainfluenza virus 2 RNA
C1113833|T201|COMP|29910-7|LNC|Parainfluenza virus 3 RNA|Parainfluenza virus 3 RNA
C1113834|T201|COMP|29911-5|LNC|Magnesium|Magnesium
C1113835|T201|COMP|29913-1|LNC|Xylose^2H post 5 g xylose PO|Xylose^2H post 5 g xylose PO
C1113836|T201|COMP|29914-9|LNC|Arsenic|Arsenic
C1113837|T201|COMP|29915-6|LNC|Tellurium|Tellurium
C1113838|T201|COMP|29916-4|LNC|Cobalt|Cobalt
C1113839|T201|COMP|29918-0|LNC|Bismuth|Bismuth
C1113840|T201|COMP|29919-8|LNC|Chromium/Creatinine|Chromium/Creatinine
C1113841|T201|COMP|29921-4|LNC|Boron|Boron
C1113842|T201|COMP|29922-2|LNC|Boron/Creatinine|Boron/Creatinine
C1113843|T201|COMP|29923-0|LNC|Scandium|Scandium
C1113844|T201|COMP|29926-3|LNC|Boron|Boron
C1113845|T201|COMP|29927-1|LNC|Beryllium|Beryllium
C1113846|T201|COMP|29928-9|LNC|Titanium|Titanium
C1113847|T201|COMP|29929-7|LNC|Titanium|Titanium
C1113848|T201|COMP|29930-5|LNC|Titanium/Creatinine|Titanium/Creatinine
C1113849|T201|COMP|29931-3|LNC|Vanadium|Vanadium
C1113850|T201|COMP|29932-1|LNC|Vanadium|Vanadium
C1113851|T201|COMP|29933-9|LNC|Vanadium/Creatinine|Vanadium/Creatinine
C1113852|T201|COMP|29934-7|LNC|Cobalt/Creatinine|Cobalt/Creatinine
C1113853|T201|COMP|29935-4|LNC|Manganese/Creatinine|Manganese/Creatinine
C1113854|T201|COMP|29936-2|LNC|Nickel|Nickel
C1113855|T201|COMP|29937-0|LNC|Aluminum/Creatinine|Aluminum/Creatinine
C1113856|T201|COMP|29938-8|LNC|Thallium/Creatinine|Thallium/Creatinine
C1113857|T201|COMP|29939-6|LNC|Tellurium/Creatinine|Tellurium/Creatinine
C1113858|T201|COMP|29940-4|LNC|Bismuth/Creatinine|Bismuth/Creatinine
C1113859|T201|COMP|29941-2|LNC|Antimony/Creatinine|Antimony/Creatinine
C1113860|T201|COMP|29942-0|LNC|Copper/Creatinine|Copper/Creatinine
C1113861|T201|COMP|29943-8|LNC|Lead/Creatinine|Lead/Creatinine
C1113862|T201|COMP|29944-6|LNC|Alpha-2-Macroglobulin|Alpha-2-Macroglobulin
C1113863|T201|COMP|29945-3|LNC|Alpha 1 globulin|Alpha 1 globulin
C1113864|T201|COMP|29946-1|LNC|Albumin|Albumin
C1113865|T201|COMP|29947-9|LNC|Alpha 2 globulin|Alpha 2 globulin
C1113866|T201|COMP|29948-7|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C1113867|T201|COMP|29949-5|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C1113868|T201|COMP|29950-3|LNC|Nuclear Ab.IgG|Nuclear Ab.IgG
C1113869|T201|COMP|29951-1|LNC|Beta globulin|Beta globulin
C1113870|T201|COMP|29952-9|LNC|Borrelia burgdorferi Ag|Borrelia burgdorferi Ag
C1113871|T201|COMP|29954-5|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C1113872|T201|COMP|29955-2|LNC|Legionella pneumophila Ab.IgG|Legionella pneumophila Ab.IgG
C1113873|T201|COMP|29956-0|LNC|Lysozyme|Lysozyme
C1113874|T201|COMP|29957-8|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1113875|T201|COMP|29958-6|LNC|Ribonucleoprotein extractable nuclear Ab.IgG|Ribonucleoprotein extractable nuclear Ab.IgG
C1113876|T201|COMP|29959-4|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C1113877|T201|COMP|29960-2|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C1113878|T201|COMP|29961-0|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C1113879|T201|COMP|29962-8|LNC|Asialoganglioside GM1 Ab.IgM|Asialoganglioside GM1 Ab.IgM
C1113880|T201|COMP|29963-6|LNC|Parietal cell Ab.IgG|Parietal cell Ab.IgG
C1113881|T201|COMP|29965-1|LNC|Sjogrens syndrome-B extractable nuclear Ab.IgG|Sjogrens syndrome-B extractable nuclear Ab.IgG
C1113882|T201|COMP|29966-9|LNC|Centromere Ab.IgG|Centromere Ab.IgG
C1113883|T201|COMP|29967-7|LNC|Neutrophil cytoplasmic Ab.IgG|Neutrophil cytoplasmic Ab.IgG
C1113884|T201|COMP|29968-5|LNC|Rubidium|Rubidium
C1113885|T201|COMP|29969-3|LNC|Rubidium|Rubidium
C1113886|T201|COMP|29970-1|LNC|Rubidium/Creatinine|Rubidium/Creatinine
C1113887|T201|COMP|29971-9|LNC|Strontium|Strontium
C1113888|T201|COMP|29972-7|LNC|Strontium|Strontium
C1113889|T201|COMP|29974-3|LNC|Molybdenum|Molybdenum
C1113890|T201|COMP|29975-0|LNC|Molybdenum|Molybdenum
C1113891|T201|COMP|29976-8|LNC|Molybdenum/Creatinine|Molybdenum/Creatinine
C1113892|T201|COMP|29977-6|LNC|Silver|Silver
C1113893|T201|COMP|29979-2|LNC|Tin|Tin
C1113894|T201|COMP|29980-0|LNC|Tin|Tin
C1113895|T201|COMP|29983-4|LNC|Cesium|Cesium
C1113896|T201|COMP|29984-2|LNC|Cesium/Creatinine|Cesium/Creatinine
C1113897|T201|COMP|29985-9|LNC|Barium|Barium
C1113898|T201|COMP|29987-5|LNC|Gold|Gold
C1113899|T201|COMP|29988-3|LNC|Gold/Creatinine|Gold/Creatinine
C1113900|T201|COMP|29989-1|LNC|Uranium/Creatinine|Uranium/Creatinine
C1113901|T201|COMP|29990-9|LNC|Spermatozoa^post vasectomy|Spermatozoa^post vasectomy
C1113902|T201|COMP|29991-7|LNC|Fibrin+Fibrinogen fragments|Fibrin+Fibrinogen fragments
C1113903|T201|COMP|29992-5|LNC|Eosinophils|Eosinophils
C1113904|T201|COMP|29993-3|LNC|Eosinophils|Eosinophils
C1113905|T201|COMP|29995-8|LNC|Basement membrane Ab.IgA|Basement membrane Ab.IgA
C1113906|T201|COMP|29996-6|LNC|Histone Ab.IgG|Histone Ab.IgG
C1113907|T201|COMP|29997-4|LNC|Basement membrane Ab.IgG|Basement membrane Ab.IgG
C1113908|T201|COMP|29998-2|LNC|Striated muscle Ab.IgG|Striated muscle Ab.IgG
C1113909|T201|COMP|29999-0|LNC|Xylose|Xylose
C1113910|T201|COMP|30000-4|LNC|Albumin/Creatinine|Albumin/Creatinine
C1113911|T201|COMP|30001-2|LNC|Albumin/Creatinine|Albumin/Creatinine
C1113912|T201|COMP|30002-0|LNC|Creatinine|Creatinine
C1113913|T201|COMP|30003-8|LNC|Albumin|Albumin
C1113914|T201|COMP|30004-6|LNC|Creatinine|Creatinine
C1113915|T201|COMP|30005-3|LNC|CYP21A2 gene targeted mutation analysis|CYP21A2 gene targeted mutation analysis
C1113916|T201|COMP|30006-1|LNC|Transfuse granulocytes|Transfuse granulocytes
C1113917|T201|COMP|30007-9|LNC|Transfuse cryoprecipitate poor plasma|Transfuse cryoprecipitate poor plasma
C1113918|T201|COMP|30008-7|LNC|Blood group antibody screen|Blood group antibody screen
C1113919|T201|COMP|30009-5|LNC|Fibrin+Fibrinogen fragments|Fibrin+Fibrinogen fragments
C1113920|T201|COMP|30010-3|LNC|Borrelia burgdorferi 93kD Ab.IgG|Borrelia burgdorferi 93kD Ab.IgG
C1113921|T201|COMP|30011-1|LNC|Borrelia burgdorferi 45kD Ab.IgG|Borrelia burgdorferi 45kD Ab.IgG
C1113922|T201|COMP|30012-9|LNC|Borrelia burgdorferi 28kD Ab.IgG|Borrelia burgdorferi 28kD Ab.IgG
C1113923|T201|COMP|30013-7|LNC|Borrelia burgdorferi 23kD Ab.IgG|Borrelia burgdorferi 23kD Ab.IgG
C1113924|T201|COMP|30014-5|LNC|Borrelia burgdorferi 21kD Ab.IgG|Borrelia burgdorferi 21kD Ab.IgG
C1113925|T201|COMP|30016-0|LNC|Borrelia burgdorferi 66kD Ab.IgG|Borrelia burgdorferi 66kD Ab.IgG
C1113926|T201|COMP|30017-8|LNC|Borrelia burgdorferi 58kD Ab.IgG|Borrelia burgdorferi 58kD Ab.IgG
C1113927|T201|COMP|30018-6|LNC|Borrelia burgdorferi 30kD Ab.IgG|Borrelia burgdorferi 30kD Ab.IgG
C1113928|T201|COMP|30019-4|LNC|Borrelia burgdorferi 41kD Ab.IgM|Borrelia burgdorferi 41kD Ab.IgM
C1113929|T201|COMP|30020-2|LNC|Borrelia burgdorferi 39kD Ab.IgM|Borrelia burgdorferi 39kD Ab.IgM
C1113930|T201|COMP|30021-0|LNC|Borrelia burgdorferi 23kD Ab.IgM|Borrelia burgdorferi 23kD Ab.IgM
C1113931|T201|COMP|30022-8|LNC|Botrytis cinerea Ab.IgG|Botrytis cinerea Ab.IgG
C1113932|T201|COMP|30024-4|LNC|Carbophenothion|Carbophenothion
C1113933|T201|COMP|30025-1|LNC|Coumaphos|Coumaphos
C1113934|T201|COMP|30026-9|LNC|Dichlorvos|Dichlorvos
C1113935|T201|COMP|30027-7|LNC|Dimethoate|Dimethoate
C1113936|T201|COMP|30029-3|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C1113937|T201|COMP|30030-1|LNC|Iron|Iron
C1113939|T201|COMP|30032-7|LNC|Phoma betae Ab.IgG|Phoma betae Ab.IgG
C1113940|T201|COMP|30034-3|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C1113941|T201|COMP|30035-0|LNC|Homocystine^post CFst|Homocystine^post CFst
C1113942|T201|COMP|30036-8|LNC|Aspergillus fumigatus 2 Ab|Aspergillus fumigatus 2 Ab
C1113944|T201|COMP|30038-4|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C1113945|T201|COMP|30040-0|LNC|Dirofilaria immitis Ab|Dirofilaria immitis Ab
C1113946|T201|COMP|30041-8|LNC|Curcuma longa Ab.IgE|Curcuma longa Ab.IgE
C1113947|T201|COMP|30042-6|LNC|Vigabatrin|Vigabatrin
C1113948|T201|COMP|30043-4|LNC|Rosmarinus officinalis Ab.IgE|Rosmarinus officinalis Ab.IgE
C1113949|T201|COMP|30045-9|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C1113950|T201|COMP|30046-7|LNC|Legionella pneumophila Ab|Legionella pneumophila Ab
C1113951|T201|COMP|30047-5|LNC|Histidine/Creatinine|Histidine/Creatinine
C1113952|T201|COMP|30049-1|LNC|Ornithine/Creatinine|Ornithine/Creatinine
C1113953|T201|COMP|30050-9|LNC|Hydroxylysine/Creatinine|Hydroxylysine/Creatinine
C1113954|T201|COMP|30053-3|LNC|Leucine/Creatinine|Leucine/Creatinine
C1113955|T201|COMP|30054-1|LNC|Tyrosine/Creatinine|Tyrosine/Creatinine
C1113956|T201|COMP|30055-8|LNC|Phenylalanine/Creatinine|Phenylalanine/Creatinine
C1113957|T201|COMP|30057-4|LNC|Threonine/Creatinine|Threonine/Creatinine
C1113958|T201|COMP|30058-2|LNC|Serine/Creatinine|Serine/Creatinine
C1113959|T201|COMP|30059-0|LNC|Glutamate/Creatinine|Glutamate/Creatinine
C1113960|T201|COMP|30060-8|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C1113961|T201|COMP|30061-6|LNC|Aspartate/Creatinine|Aspartate/Creatinine
C1113962|T201|COMP|30062-4|LNC|Arginine/Creatinine|Arginine/Creatinine
C1113963|T201|COMP|30063-2|LNC|Methionine/Creatinine|Methionine/Creatinine
C1113964|T201|COMP|30064-0|LNC|Valine/Creatinine|Valine/Creatinine
C1113965|T201|COMP|30065-7|LNC|Cystine/Creatinine|Cystine/Creatinine
C1113966|T201|COMP|30066-5|LNC|Glycine/Creatinine|Glycine/Creatinine
C1113967|T201|COMP|30067-3|LNC|Proline/Creatinine|Proline/Creatinine
C1113968|T201|COMP|30068-1|LNC|Alanine/Creatinine|Alanine/Creatinine
C1113969|T201|COMP|30069-9|LNC|Tyrosine|Tyrosine
C1113970|T201|COMP|30070-7|LNC|Cystathionine|Cystathionine
C1113971|T201|COMP|30071-5|LNC|Trichoderma viride Ab.IgG|Trichoderma viride Ab.IgG
C1113972|T201|COMP|30072-3|LNC|Cortisone|Cortisone
C1113973|T201|COMP|30073-1|LNC|Voltage-gated calcium channel Ab|Voltage-gated calcium channel Ab
C1113974|T201|COMP|30074-9|LNC|Hemoglobin F|Hemoglobin F
C1113975|T201|COMP|30075-6|LNC|Respiratory syncytial virus A RNA|Respiratory syncytial virus A RNA
C1113976|T201|COMP|30076-4|LNC|Respiratory syncytial virus B RNA|Respiratory syncytial virus B RNA
C1113977|T201|COMP|30077-2|LNC|Amylase/Creatinine renal clearance|Amylase/Creatinine renal clearance
C1113978|T201|COMP|30078-0|LNC|Specimen weight|Specimen weight
C1113979|T201|COMP|30079-8|LNC|Renal tubular casts|Renal tubular casts
C1113980|T201|COMP|30080-6|LNC|Cathepsin D|Cathepsin D
C1113981|T201|COMP|30081-4|LNC|IgD|IgD
C1113982|T201|COMP|30083-0|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C1113983|T201|COMP|30085-5|LNC|Legionella pneumophila Ab.IgG|Legionella pneumophila Ab.IgG
C1113984|T201|COMP|30086-3|LNC|Coagulation factor IX inhibitor|Coagulation factor IX inhibitor
C1113985|T201|COMP|30087-1|LNC|Cow hair+Cow dander Ab.IgE|Cow hair+Cow dander Ab.IgE
C1113986|T201|COMP|30088-9|LNC|Horse hair+Horse dander Ab.IgE|Horse hair+Horse dander Ab.IgE
C1113987|T201|COMP|30089-7|LNC|Transitional cells|Transitional cells
C1113988|T201|COMP|30090-5|LNC|Burkholderia pseudomallei Ab.IgG|Burkholderia pseudomallei Ab.IgG
C1113989|T201|COMP|30091-3|LNC|Burkholderia pseudomallei Ab.IgM|Burkholderia pseudomallei Ab.IgM
C1113990|T201|COMP|30092-1|LNC|Brucella canis Ab.IgG|Brucella canis Ab.IgG
C1113991|T201|COMP|30094-7|LNC|Neisseria meningitidis serogroup A Ag|Neisseria meningitidis serogroup A Ag
C1113992|T201|COMP|30095-4|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C1113993|T201|COMP|30096-2|LNC|Neisseria meningitidis serogroup C Ag|Neisseria meningitidis serogroup C Ag
C1113994|T201|COMP|30097-0|LNC|Neisseria meningitidis serogroup w135 Ag|Neisseria meningitidis serogroup w135 Ag
C1113995|T201|COMP|30099-6|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C1113996|T201|COMP|30100-2|LNC|Yersinia enterocolitica O:3 Ab|Yersinia enterocolitica O:3 Ab
C1113997|T201|COMP|30102-8|LNC|Yersinia enterocolitica O:8 Ab|Yersinia enterocolitica O:8 Ab
C1113998|T201|COMP|30103-6|LNC|Yersinia enterocolitica O:9 Ab|Yersinia enterocolitica O:9 Ab
C1113999|T201|COMP|30104-4|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C1114000|T201|COMP|30105-1|LNC|Trypanosoma cruzi Ab.IgM|Trypanosoma cruzi Ab.IgM
C1114001|T201|COMP|30107-7|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C1114002|T201|COMP|30108-5|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C1114003|T201|COMP|30109-3|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C1114004|T201|COMP|30111-9|LNC|Thermoactinomyces vulgaris 2 Ab|Thermoactinomyces vulgaris 2 Ab
C1114005|T201|COMP|30112-7|LNC|Amphetamine|Amphetamine
C1114006|T201|COMP|30113-5|LNC|Lymphocytes.IgG|Lymphocytes.IgG
C1114007|T201|COMP|30115-0|LNC|Lymphocytes.kappa|Lymphocytes.kappa
C1114010|T201|COMP|30118-4|LNC|Lymphocytes.IgA|Lymphocytes.IgA
C1114011|T201|COMP|30119-2|LNC|Lymphocytes.IgM|Lymphocytes.IgM
C1114012|T201|COMP|30120-0|LNC|Lymphocytes.IgD|Lymphocytes.IgD
C1114013|T201|COMP|30121-8|LNC|Colony count|Colony count
C1114014|T201|COMP|30122-6|LNC|Aeromonas sp|Aeromonas sp
C1114015|T201|COMP|30123-4|LNC|Testosterone.bound|Testosterone.bound
C1114016|T201|COMP|30124-2|LNC|Amylase|Amylase
C1114017|T201|COMP|30125-9|LNC|Gerbil hair Ab.IgE.RAST class|Gerbil hair Ab.IgE.RAST class
C1114018|T201|COMP|30126-7|LNC|Platanus acerifolia Ab.IgE.RAST class|Platanus acerifolia Ab.IgE.RAST class
C1114019|T201|COMP|30127-5|LNC|Gerbil hair Ab.IgE|Gerbil hair Ab.IgE
C1114020|T201|COMP|30128-3|LNC|Borrelia burgdorferi Ab^2nd specimen|Borrelia burgdorferi Ab^2nd specimen
C1114021|T201|COMP|30129-1|LNC|Brucella sp Ab^1st specimen|Brucella sp Ab^1st specimen
C1114022|T201|COMP|30130-9|LNC|Brucella sp Ab^2nd specimen|Brucella sp Ab^2nd specimen
C1114023|T201|COMP|30131-7|LNC|Complement total hemolytic CH50|Complement total hemolytic CH50
C1114024|T201|COMP|30132-5|LNC|Coxsackievirus Ab^1st specimen|Coxsackievirus Ab^1st specimen
C1114025|T201|COMP|30133-3|LNC|Coxsackievirus Ab^2nd specimen|Coxsackievirus Ab^2nd specimen
C1114026|T201|COMP|30134-1|LNC|Echovirus Ab^1st specimen|Echovirus Ab^1st specimen
C1114027|T201|COMP|30135-8|LNC|Echovirus Ab^2nd specimen|Echovirus Ab^2nd specimen
C1114028|T201|COMP|30136-6|LNC|Epstein Barr virus capsid Ab.IgG^2nd specimen|Epstein Barr virus capsid Ab.IgG^2nd specimen
C1114029|T201|COMP|30137-4|LNC|Epstein Barr virus capsid Ab.IgM^2nd specimen|Epstein Barr virus capsid Ab.IgM^2nd specimen
C1114030|T201|COMP|30139-0|LNC|Hydroxyproline.free|Hydroxyproline.free
C1114031|T201|COMP|30140-8|LNC|IgA|IgA
C1114032|T201|COMP|30141-6|LNC|IgG|IgG
C1114033|T201|COMP|30142-4|LNC|IgM|IgM
C1114034|T201|COMP|30143-2|LNC|Legionella sp Ab^1st specimen|Legionella sp Ab^1st specimen
C1114035|T201|COMP|30144-0|LNC|Legionella sp Ab^2nd specimen|Legionella sp Ab^2nd specimen
C1114036|T201|COMP|30145-7|LNC|Monocytes|Monocytes
C1114037|T201|COMP|30146-5|LNC|Mumps virus Ab^2nd specimen|Mumps virus Ab^2nd specimen
C1114038|T201|COMP|30147-3|LNC|Respiratory syncytial virus Ab^1st specimen|Respiratory syncytial virus Ab^1st specimen
C1114039|T201|COMP|30148-1|LNC|Respiratory syncytial virus Ab^2nd specimen|Respiratory syncytial virus Ab^2nd specimen
C1114040|T201|COMP|30150-7|LNC|Streptolysin O Ab^2nd specimen|Streptolysin O Ab^2nd specimen
C1114041|T201|COMP|30151-5|LNC|Thyrotropin.long acting|Thyrotropin.long acting
C1114042|T201|COMP|30152-3|LNC|Mannose-binding protein|Mannose-binding protein
C1114043|T201|COMP|30154-9|LNC|Protein/Creatinine|Protein/Creatinine
C1114044|T201|COMP|30155-6|LNC|Reticulocytes.punctate/100 erythrocytes|Reticulocytes.punctate/100 erythrocytes
C1114045|T201|COMP|30156-4|LNC|Reticulocytes.aggregate/100 erythrocytes|Reticulocytes.aggregate/100 erythrocytes
C1114046|T201|COMP|30157-2|LNC|Heterophils/100 leukocytes|Heterophils/100 leukocytes
C1114047|T201|COMP|30159-8|LNC|HTLV I+II DNA|HTLV I+II DNA
C1114048|T201|COMP|30160-6|LNC|Tau protein|Tau protein
C1114049|T201|COMP|30161-4|LNC|Citrulline/Creatinine|Citrulline/Creatinine
C1114050|T201|COMP|30163-0|LNC|Agapostemon texanus Ab.IgE|Agapostemon texanus Ab.IgE
C1114052|T201|COMP|30165-5|LNC|Phosphatidylcholine/Albumin|Phosphatidylcholine/Albumin
C1114053|T201|COMP|30166-3|LNC|Thyroid stimulating immunoglobulins actual/Normal|Thyroid stimulating immunoglobulins actual/Normal
C1114054|T201|COMP|30168-9|LNC|Juniperus monosperma Ab.IgE|Juniperus monosperma Ab.IgE
C1114055|T201|COMP|30169-7|LNC|Chromogranin A|Chromogranin A
C1114056|T201|COMP|30170-5|LNC|Periplaneta americana Ab.IgE|Periplaneta americana Ab.IgE
C1114057|T201|COMP|30171-3|LNC|Cortisol.free/Creatinine|Cortisol.free/Creatinine
C1114058|T201|COMP|30172-1|LNC|Cortisol.free/Creatinine|Cortisol.free/Creatinine
C1114059|T201|COMP|30174-7|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C1114060|T201|COMP|30175-4|LNC|Jamestown canyon virus Ab|Jamestown canyon virus Ab
C1114061|T201|COMP|30176-2|LNC|La Crosse virus Ab|La Crosse virus Ab
C1114062|T201|COMP|30177-0|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1114063|T201|COMP|30178-8|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C1114064|T201|COMP|30179-6|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1114065|T201|COMP|30180-4|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1114066|T201|COMP|30181-2|LNC|Lymphocytes.clefted|Lymphocytes.clefted
C1114075|T201|COMP|30190-3|LNC|3-Hydroxytetradecenoylcarnitine (C14:1-OH)|3-Hydroxytetradecenoylcarnitine (C14:1-OH)
C1114076|T201|COMP|30191-1|LNC|Acetylcarnitine (C2)|Acetylcarnitine (C2)
C1114078|T201|COMP|30193-7|LNC|Acylcarnitine/Carnitine.free (C0)|Acylcarnitine/Carnitine.free (C0)
C1114079|T201|COMP|30194-5|LNC|Fatty acids.very long chain.C22:0|Fatty acids.very long chain.C22:0
C1114080|T201|COMP|30195-2|LNC|Fatty acids.very long chain.C24:0|Fatty acids.very long chain.C24:0
C1114081|T201|COMP|30196-0|LNC|Fatty acids.very long chain.C24:0/C22:0|Fatty acids.very long chain.C24:0/C22:0
C1114082|T201|COMP|30197-8|LNC|Fatty acids.very long chain.C26:0|Fatty acids.very long chain.C26:0
C1114083|T201|COMP|30198-6|LNC|Fatty acids.very long chain.C26:0/C22:0|Fatty acids.very long chain.C26:0/C22:0
C1114084|T201|COMP|30199-4|LNC|Alpha subunit|Alpha subunit
C1114085|T201|COMP|30200-0|LNC|Asialoganglioside GM1 Ab.IgM|Asialoganglioside GM1 Ab.IgM
C1114086|T201|COMP|30201-8|LNC|B Ab|B Ab
C1114087|T201|COMP|30202-6|LNC|Brucella sp Ab|Brucella sp Ab
C1114088|T201|COMP|30204-2|LNC|Chlamydia trachomatis Ab|Chlamydia trachomatis Ab
C1114089|T201|COMP|30206-7|LNC|Choriogonadotropin.alpha subunit.free|Choriogonadotropin.alpha subunit.free
C1114090|T201|COMP|30207-5|LNC|Coccidioides immitis Ab.IgG|Coccidioides immitis Ab.IgG
C1114091|T201|COMP|30208-3|LNC|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C1114092|T201|COMP|30209-1|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C1114094|T201|COMP|30211-7|LNC|Collection duration|Collection duration
C1114095|T201|COMP|30212-5|LNC|Coxiella burnetii Ab.IgG|Coxiella burnetii Ab.IgG
C1114096|T201|COMP|30213-3|LNC|Coxiella burnetii Ab.IgM|Coxiella burnetii Ab.IgM
C1114097|T201|COMP|30215-8|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C1114098|T201|COMP|30216-6|LNC|Coxsackievirus A2 Ab|Coxsackievirus A2 Ab
C1114099|T201|COMP|30217-4|LNC|Coxsackievirus A4 Ab|Coxsackievirus A4 Ab
C1114100|T201|COMP|30218-2|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C1114101|T201|COMP|30220-8|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C1114102|T201|COMP|30221-6|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C1114103|T201|COMP|30223-2|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C1114104|T201|COMP|30224-0|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C1114105|T201|COMP|30225-7|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C1114106|T201|COMP|30226-5|LNC|Fibrin+Fibrinogen fragments|Fibrin+Fibrinogen fragments
C1114107|T201|COMP|30228-1|LNC|Mumps reaction wheal^2D post 0.1 mL mumps ID|Mumps reaction wheal^2D post 0.1 mL mumps ID
C1114108|T201|COMP|30229-9|LNC|Neutrophils.band form|Neutrophils.band form
C1114109|T201|COMP|30230-7|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C1114110|T201|COMP|30231-5|LNC|Rheumatoid factor|Rheumatoid factor
C1114112|T201|COMP|30233-1|LNC|3-Hydroxydodecanoylcarnitine (C12-OH)|3-Hydroxydodecanoylcarnitine (C12-OH)
C1114113|T201|COMP|30235-6|LNC|3-Hydroxypalmitoleylcarnitine (C16:1-OH)|3-Hydroxypalmitoleylcarnitine (C16:1-OH)
C1114114|T201|COMP|30236-4|LNC|3-Hydroxyhexanoylcarnitine (C6-OH)|3-Hydroxyhexanoylcarnitine (C6-OH)
C1114115|T201|COMP|30237-2|LNC|3-Hydroxylinoleoylcarnitine (C18:2-OH)|3-Hydroxylinoleoylcarnitine (C18:2-OH)
C1114116|T201|COMP|30238-0|LNC|3-Hydroxytetradecanoylcarnitine (C14-OH)|3-Hydroxytetradecanoylcarnitine (C14-OH)
C1114117|T201|COMP|30239-8|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C1114118|T201|COMP|30240-6|LNC|Fibrin D-dimer|Fibrin D-dimer
C1114119|T201|COMP|30241-4|LNC|Lactate|Lactate
C1114120|T201|COMP|30242-2|LNC|Lactate|Lactate
C1114121|T201|COMP|30243-0|LNC|Choriogonadotropin.intact|Choriogonadotropin.intact
C1114122|T201|COMP|30244-8|LNC|Acetylcholinesterase|Acetylcholinesterase
C1114123|T201|COMP|30245-5|LNC|HIV 1 DNA|HIV 1 DNA
C1114124|T201|COMP|30246-3|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1114125|T201|COMP|30247-1|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1114126|T201|COMP|30248-9|LNC|Transferrin receptor.soluble|Transferrin receptor.soluble
C1114127|T201|COMP|30249-7|LNC|Barbiturates|Barbiturates
C1114128|T201|COMP|30250-5|LNC|Benzodiazepines|Benzodiazepines
C1114129|T201|COMP|30251-3|LNC|Glucose^2.6H post dose glucose|Glucose^2.6H post dose glucose
C1114130|T201|COMP|30252-1|LNC|Glucose^3.3H post dose glucose|Glucose^3.3H post dose glucose
C1114131|T201|COMP|30253-9|LNC|Glucose^3.6H post dose glucose|Glucose^3.6H post dose glucose
C1114132|T201|COMP|30254-7|LNC|Insulin^15M post XXX challenge|Insulin^15M post XXX challenge
C1114133|T201|COMP|30255-4|LNC|Insulin^45M post XXX challenge|Insulin^45M post XXX challenge
C1114134|T201|COMP|30256-2|LNC|Insulin^1.3H post XXX challenge|Insulin^1.3H post XXX challenge
C1114135|T201|COMP|30257-0|LNC|Insulin^1.6H post XXX challenge|Insulin^1.6H post XXX challenge
C1114136|T201|COMP|30258-8|LNC|Insulin^2.3H post XXX challenge|Insulin^2.3H post XXX challenge
C1114137|T201|COMP|30259-6|LNC|Insulin^2.6H post XXX challenge|Insulin^2.6H post XXX challenge
C1114138|T201|COMP|30260-4|LNC|Insulin^3.3H post XXX challenge|Insulin^3.3H post XXX challenge
C1114139|T201|COMP|30262-0|LNC|Insulin^3.6H post XXX challenge|Insulin^3.6H post XXX challenge
C1114140|T201|COMP|30263-8|LNC|Glucose^20M post dose glucose|Glucose^20M post dose glucose
C1114141|T201|COMP|30265-3|LNC|Glucose^1.3H post dose glucose|Glucose^1.3H post dose glucose
C1114142|T201|COMP|30267-9|LNC|Glucose^2.3H post dose glucose|Glucose^2.3H post dose glucose
C1114143|T201|COMP|30268-7|LNC|Zidovudine|Zidovudine
C1114144|T201|COMP|30269-5|LNC|lamiVUDine|lamiVUDine
C1114145|T201|COMP|30270-3|LNC|Didanosine|Didanosine
C1114146|T201|COMP|30272-9|LNC|Stavudine|Stavudine
C1114147|T201|COMP|30273-7|LNC|Abacavir|Abacavir
C1114148|T201|COMP|30274-5|LNC|Adefovir|Adefovir
C1114149|T201|COMP|30275-2|LNC|Nevirapine|Nevirapine
C1114150|T201|COMP|30277-8|LNC|Efavirenz|Efavirenz
C1114151|T201|COMP|30278-6|LNC|Indinavir|Indinavir
C1114152|T201|COMP|30279-4|LNC|Ritonavir|Ritonavir
C1114153|T201|COMP|30281-0|LNC|Saquinavir|Saquinavir
C1114154|T201|COMP|30282-8|LNC|Zidovudine|Zidovudine
C1114155|T201|COMP|30283-6|LNC|lamiVUDine|lamiVUDine
C1114156|T201|COMP|30284-4|LNC|Didanosine|Didanosine
C1114157|T201|COMP|30286-9|LNC|Stavudine|Stavudine
C1114158|T201|COMP|30287-7|LNC|Abacavir|Abacavir
C1114159|T201|COMP|30288-5|LNC|Adefovir|Adefovir
C1114160|T201|COMP|30289-3|LNC|Nevirapine|Nevirapine
C1114161|T201|COMP|30290-1|LNC|Delavirdine|Delavirdine
C1114162|T201|COMP|30291-9|LNC|Efavirenz|Efavirenz
C1114163|T201|COMP|30292-7|LNC|Indinavir|Indinavir
C1114164|T201|COMP|30293-5|LNC|Ritonavir|Ritonavir
C1114165|T201|COMP|30294-3|LNC|Nelfinavir|Nelfinavir
C1114166|T201|COMP|30295-0|LNC|Saquinavir|Saquinavir
C1114167|T201|COMP|30296-8|LNC|Amprenavir|Amprenavir
C1114168|T201|COMP|30297-6|LNC|Amprenavir|Amprenavir
C1114169|T201|COMP|30298-4|LNC|lamiVUDine|lamiVUDine
C1114170|T201|COMP|30299-2|LNC|Amprenavir|Amprenavir
C1114171|T201|COMP|30300-8|LNC|Didanosine|Didanosine
C1114172|T201|COMP|30301-6|LNC|Zalcitabine|Zalcitabine
C1114173|T201|COMP|30302-4|LNC|Stavudine|Stavudine
C1114174|T201|COMP|30303-2|LNC|Abacavir|Abacavir
C1114175|T201|COMP|30304-0|LNC|Adefovir|Adefovir
C1114176|T201|COMP|30305-7|LNC|Delavirdine|Delavirdine
C1114177|T201|COMP|30306-5|LNC|Efavirenz|Efavirenz
C1114178|T201|COMP|30307-3|LNC|Indinavir|Indinavir
C1114179|T201|COMP|30308-1|LNC|Ritonavir|Ritonavir
C1114180|T201|COMP|30309-9|LNC|Nelfinavir|Nelfinavir
C1114181|T201|COMP|30310-7|LNC|Saquinavir|Saquinavir
C1114182|T201|COMP|30311-5|LNC|Nevirapine|Nevirapine
C1114183|T201|COMP|30312-3|LNC|3-Hydroxyoleoylcarnitine (C18:1-OH)|3-Hydroxyoleoylcarnitine (C18:1-OH)
C1114184|T201|COMP|30313-1|LNC|Hemoglobin|Hemoglobin
C1114185|T201|COMP|30314-9|LNC|A Ab|A Ab
C1114186|T201|COMP|30316-4|LNC|Alpha subunit.free|Alpha subunit.free
C1114187|T201|COMP|30317-2|LNC|Base deficit|Base deficit
C1114188|T201|COMP|30318-0|LNC|Base deficit|Base deficit
C1114189|T201|COMP|30319-8|LNC|Beta galactosidase|Beta galactosidase
C1114190|T201|COMP|30320-6|LNC|Cells.CD3+IL2R1+|Cells.CD3+IL2R1+
C1114194|T201|COMP|30325-5|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C1114195|T201|COMP|30326-3|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1114196|T201|COMP|30327-1|LNC|Decanoylcarnitine (C10)|Decanoylcarnitine (C10)
C1114197|T201|COMP|30328-9|LNC|Decenoylcarnitine (C10:1)|Decenoylcarnitine (C10:1)
C1114198|T201|COMP|30330-5|LNC|Disialylganglioside GD1b Ab.IgM|Disialylganglioside GD1b Ab.IgM
C1114199|T201|COMP|30331-3|LNC|Dodecanoylcarnitine (C12)|Dodecanoylcarnitine (C12)
C1114200|T201|COMP|30332-1|LNC|Dodecenoylcarnitine (C12:1)|Dodecenoylcarnitine (C12:1)
C1114201|T201|COMP|30334-7|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C1114202|T201|COMP|30335-4|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C1114203|T201|COMP|30336-2|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C1114204|T201|COMP|30338-8|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C1114205|T201|COMP|30339-6|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C1114206|T201|COMP|30340-4|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C1114207|T201|COMP|30342-0|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C1114208|T201|COMP|30343-8|LNC|Glomerular basement membrane Ab.IgG|Glomerular basement membrane Ab.IgG
C1114209|T201|COMP|30344-6|LNC|Glucose^1H post 1.2 g/kg lactose PO|Glucose^1H post 1.2 g/kg lactose PO
C1114210|T201|COMP|30345-3|LNC|Glucose^2H post 1.2 g/kg lactose PO|Glucose^2H post 1.2 g/kg lactose PO
C1114211|T201|COMP|30347-9|LNC|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C1114212|T201|COMP|30349-5|LNC|Glutarylcarnitine (C5-DC)|Glutarylcarnitine (C5-DC)
C1114213|T201|COMP|30350-3|LNC|Hemoglobin|Hemoglobin
C1114214|T201|COMP|30351-1|LNC|Hemoglobin|Hemoglobin
C1114215|T201|COMP|30352-9|LNC|Hemoglobin|Hemoglobin
C1114216|T201|COMP|30353-7|LNC|Hemoglobin|Hemoglobin
C1114217|T201|COMP|30355-2|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1114218|T201|COMP|30356-0|LNC|Palmitoylcarnitine (C16)|Palmitoylcarnitine (C16)
C1114219|T201|COMP|30357-8|LNC|Palmitoleylcarnitine (C16:1)|Palmitoleylcarnitine (C16:1)
C1114220|T201|COMP|30358-6|LNC|Hexanoylcarnitine (C6)|Hexanoylcarnitine (C6)
C1114221|T201|COMP|30359-4|LNC|Histone Ab|Histone Ab
C1114222|T201|COMP|30360-2|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C1114223|T201|COMP|30361-0|LNC|HIV 2 Ab|HIV 2 Ab
C1114224|T201|COMP|30362-8|LNC|Insulin^30M post 75 g glucose PO|Insulin^30M post 75 g glucose PO
C1114225|T201|COMP|30363-6|LNC|Insulin^post 12H CFst|Insulin^post 12H CFst
C1114226|T201|COMP|30364-4|LNC|Lymphocytes|Lymphocytes
C1114227|T201|COMP|30365-1|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C1114228|T201|COMP|30366-9|LNC|Metamyelocytes/100 leukocytes|Metamyelocytes/100 leukocytes
C1114229|T201|COMP|30367-7|LNC|Myeloblasts/100 leukocytes|Myeloblasts/100 leukocytes
C1114230|T201|COMP|30368-5|LNC|Myelocytes/100 leukocytes|Myelocytes/100 leukocytes
C1114231|T201|COMP|30369-3|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C1114232|T201|COMP|30370-1|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C1114233|T201|COMP|30371-9|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C1114234|T201|COMP|30372-7|LNC|Sucrase|Sucrase
C1114235|T201|COMP|30373-5|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1114236|T201|COMP|30374-3|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1114237|T201|COMP|30375-0|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1114238|T201|COMP|30376-8|LNC|Blasts|Blasts
C1114239|T201|COMP|30377-6|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1114240|T201|COMP|30378-4|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1114241|T201|COMP|30379-2|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1114242|T201|COMP|30380-0|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1114243|T201|COMP|30381-8|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1114244|T201|COMP|30383-4|LNC|Epithelial cells|Epithelial cells
C1114245|T201|COMP|30384-2|LNC|Erythrocyte distribution width|Erythrocyte distribution width
C1114246|T201|COMP|30385-9|LNC|Erythrocyte distribution width|Erythrocyte distribution width
C1114247|T201|COMP|30386-7|LNC|Erythrocyte mean corpuscular diameter|Erythrocyte mean corpuscular diameter
C1114248|T201|COMP|30388-3|LNC|Erythrocytes|Erythrocytes
C1114249|T201|COMP|30389-1|LNC|Erythrocytes|Erythrocytes
C1114250|T201|COMP|30391-7|LNC|Erythrocytes|Erythrocytes
C1114251|T201|COMP|30392-5|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C1114252|T201|COMP|19048-8|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C1114253|T201|COMP|30395-8|LNC|Granulocytes/100 leukocytes|Granulocytes/100 leukocytes
C1114254|T201|COMP|30396-6|LNC|Granulocytes/100 leukocytes|Granulocytes/100 leukocytes
C1114255|T201|COMP|30397-4|LNC|Hairy cells|Hairy cells
C1114256|T201|COMP|30398-2|LNC|Hematocrit|Hematocrit
C1114257|T201|COMP|30400-6|LNC|Hypochromia|Hypochromia
C1114258|T201|COMP|30401-4|LNC|Leukocytes|Leukocytes
C1114259|T201|COMP|30403-0|LNC|Leukocytes|Leukocytes
C1114260|T201|COMP|30404-8|LNC|Leukocytes|Leukocytes
C1114261|T201|COMP|30405-5|LNC|Leukocytes|Leukocytes
C1114262|T201|COMP|30407-1|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C1114263|T201|COMP|30408-9|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C1114264|T201|COMP|30411-3|LNC|Leukocytes.left shift|Leukocytes.left shift
C1114265|T201|COMP|30412-1|LNC|Lymphocytes.abnormal|Lymphocytes.abnormal
C1114266|T201|COMP|30413-9|LNC|Lymphocytes.abnormal/100 leukocytes|Lymphocytes.abnormal/100 leukocytes
C1114267|T201|COMP|30414-7|LNC|Lymphocytes.abnormal/100 leukocytes|Lymphocytes.abnormal/100 leukocytes
C1114268|T201|COMP|30415-4|LNC|Lymphocytes.abnormal/100 leukocytes|Lymphocytes.abnormal/100 leukocytes
C1114269|T201|COMP|30416-2|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C1114270|T201|COMP|30417-0|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C1114271|T201|COMP|30418-8|LNC|Lymphocytes.clefted|Lymphocytes.clefted
C1114272|T201|COMP|30419-6|LNC|Lymphocytes.clefted/100 leukocytes|Lymphocytes.clefted/100 leukocytes
C1114273|T201|COMP|30420-4|LNC|Lymphocytes.large granular/100 leukocytes|Lymphocytes.large granular/100 leukocytes
C1114274|T201|COMP|30421-2|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C1114275|T201|COMP|30422-0|LNC|Lymphoma cells|Lymphoma cells
C1114276|T201|COMP|30423-8|LNC|Lymphoma cells/100 leukocytes|Lymphoma cells/100 leukocytes
C1114277|T201|COMP|30424-6|LNC|Macrocytes|Macrocytes
C1114278|T201|COMP|30425-3|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C1114279|T201|COMP|30426-1|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C1114280|T201|COMP|30427-9|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C1114281|T201|COMP|30428-7|LNC|Erythrocyte mean corpuscular volume|Erythrocyte mean corpuscular volume
C1114282|T201|COMP|30429-5|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C1114283|T201|COMP|30430-3|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C1114284|T201|COMP|30431-1|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C1114285|T201|COMP|30432-9|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C1114286|T201|COMP|30433-7|LNC|Metamyelocytes|Metamyelocytes
C1114287|T201|COMP|30434-5|LNC|Microcytes|Microcytes
C1114288|T201|COMP|30435-2|LNC|Monocytes|Monocytes
C1114289|T201|COMP|30436-0|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1114290|T201|COMP|30437-8|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1114291|T201|COMP|30439-4|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1114292|T201|COMP|30440-2|LNC|Monocytes.abnormal|Monocytes.abnormal
C1114293|T201|COMP|30441-0|LNC|Monocytes.abnormal/100 leukocytes|Monocytes.abnormal/100 leukocytes
C1114294|T201|COMP|30442-8|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C1114295|T201|COMP|30443-6|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C1114296|T201|COMP|30444-4|LNC|Myeloblasts|Myeloblasts
C1114297|T201|COMP|30445-1|LNC|Myeloblasts/100 leukocytes|Myeloblasts/100 leukocytes
C1114298|T201|COMP|30447-7|LNC|Myelocytes/100 leukocytes|Myelocytes/100 leukocytes
C1114299|T201|COMP|30448-5|LNC|Neutrophils|Neutrophils
C1114300|T201|COMP|30449-3|LNC|Neutrophils.hypersegmented|Neutrophils.hypersegmented
C1114301|T201|COMP|30450-1|LNC|Neutrophils.hypersegmented/100 leukocytes|Neutrophils.hypersegmented/100 leukocytes
C1114302|T201|COMP|30451-9|LNC|Neutrophils.segmented|Neutrophils.segmented
C1114303|T201|COMP|30452-7|LNC|Neutrophils.segmented|Neutrophils.segmented
C1114304|T201|COMP|30453-5|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C1114305|T201|COMP|30455-0|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C1114306|T201|COMP|30456-8|LNC|Nonhematic cells/100 leukocytes|Nonhematic cells/100 leukocytes
C1114307|T201|COMP|30457-6|LNC|Nonhematic cells/100 leukocytes|Nonhematic cells/100 leukocytes
C1114308|T201|COMP|30458-4|LNC|Plasma cells|Plasma cells
C1114309|T201|COMP|30460-0|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C1114310|T201|COMP|30461-8|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C1114311|T201|COMP|30462-6|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C1114312|T201|COMP|30464-2|LNC|Prolymphocytes|Prolymphocytes
C1114313|T201|COMP|30465-9|LNC|Prolymphocytes/100 leukocytes|Prolymphocytes/100 leukocytes
C1114314|T201|COMP|30466-7|LNC|Promonocytes/100 leukocytes|Promonocytes/100 leukocytes
C1114315|T201|COMP|30467-5|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C1114316|T201|COMP|30468-3|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C1114317|T201|COMP|30470-9|LNC|Cardiolipin Ab.IgA|Cardiolipin Ab.IgA
C1114318|T201|COMP|30471-7|LNC|levETIRAcetam|levETIRAcetam
C1114319|T201|COMP|30472-5|LNC|Ethylmalonate|Ethylmalonate
C1114320|T201|COMP|30475-8|LNC|Glycerate|Glycerate
C1114321|T201|COMP|30476-6|LNC|Glyoxylate|Glyoxylate
C1114322|T201|COMP|30478-2|LNC|Malonate|Malonate
C1114323|T201|COMP|30479-0|LNC|Methylsuccinate|Methylsuccinate
C1114324|T201|COMP|30480-8|LNC|Orotate|Orotate
C1114325|T201|COMP|30481-6|LNC|Pyruvate|Pyruvate
C1114326|T201|COMP|30482-4|LNC|Suberylglycine|Suberylglycine
C1114327|T201|COMP|30483-2|LNC|Succinylacetone|Succinylacetone
C1114328|T201|COMP|30484-0|LNC|Tiglylglycine|Tiglylglycine
C1114329|T201|COMP|30485-7|LNC|Uracil|Uracil
C1114330|T201|COMP|30486-5|LNC|Catecholamines^baseline|Catecholamines^baseline
C1114331|T201|COMP|30487-3|LNC|Catecholamines^1H post XXX challenge|Catecholamines^1H post XXX challenge
C1114332|T201|COMP|30488-1|LNC|Streptococcus pneumoniae 12 Ab.IgG^1st specimen|Streptococcus pneumoniae 12 Ab.IgG^1st specimen
C1114333|T201|COMP|30489-9|LNC|Streptococcus pneumoniae 12 Ab.IgG^2nd specimen|Streptococcus pneumoniae 12 Ab.IgG^2nd specimen
C1114336|T201|COMP|30492-3|LNC|Streptococcus pneumoniae 19 Ab.IgG^1st specimen|Streptococcus pneumoniae 19 Ab.IgG^1st specimen
C1114337|T201|COMP|30493-1|LNC|Streptococcus pneumoniae 19 Ab.IgG^2nd specimen|Streptococcus pneumoniae 19 Ab.IgG^2nd specimen
C1114338|T201|COMP|30494-9|LNC|Streptococcus pneumoniae 23 Ab.IgG^1st specimen|Streptococcus pneumoniae 23 Ab.IgG^1st specimen
C1114339|T201|COMP|30495-6|LNC|Streptococcus pneumoniae 23 Ab.IgG^2nd specimen|Streptococcus pneumoniae 23 Ab.IgG^2nd specimen
C1114340|T201|COMP|30496-4|LNC|Streptococcus pneumoniae 4 Ab.IgG^1st specimen|Streptococcus pneumoniae 4 Ab.IgG^1st specimen
C1114341|T201|COMP|30497-2|LNC|Streptococcus pneumoniae 4 Ab.IgG^2nd specimen|Streptococcus pneumoniae 4 Ab.IgG^2nd specimen
C1114343|T201|COMP|30500-3|LNC|Phosphatidylserine Ab.IgA|Phosphatidylserine Ab.IgA
C1114346|T201|COMP|30503-7|LNC|Streptococcus pneumoniae 8 Ab.IgG^1st specimen|Streptococcus pneumoniae 8 Ab.IgG^1st specimen
C1114347|T201|COMP|30504-5|LNC|Streptococcus pneumoniae 8 Ab.IgG^2nd specimen|Streptococcus pneumoniae 8 Ab.IgG^2nd specimen
C1114348|T201|COMP|30505-2|LNC|Streptococcus pneumoniae 9 Ab.IgG^1st specimen|Streptococcus pneumoniae 9 Ab.IgG^1st specimen
C1114349|T201|COMP|30506-0|LNC|Streptococcus pneumoniae 9 Ab.IgG^2nd specimen|Streptococcus pneumoniae 9 Ab.IgG^2nd specimen
C1114350|T201|COMP|30507-8|LNC|Cumene|Cumene
C1114351|T201|COMP|30508-6|LNC|Etiocholanolone/Creatinine|Etiocholanolone/Creatinine
C1114352|T201|COMP|30509-4|LNC|Androsterone/Creatinine|Androsterone/Creatinine
C1114353|T201|COMP|30510-2|LNC|Estriol/Creatinine|Estriol/Creatinine
C1114354|T201|COMP|30511-0|LNC|Cortisone/Creatinine|Cortisone/Creatinine
C1114355|T201|COMP|30512-8|LNC|Pregnanetriol/Creatinine|Pregnanetriol/Creatinine
C1114356|T201|COMP|30513-6|LNC|Pregnanetriolone/Creatinine|Pregnanetriolone/Creatinine
C1114357|T201|COMP|30515-1|LNC|Tetrahydroaldosterone/Creatinine|Tetrahydroaldosterone/Creatinine
C1114358|T201|COMP|30516-9|LNC|Bromodiphenhydramine|Bromodiphenhydramine
C1114359|T201|COMP|30517-7|LNC|Carbinoxamine|Carbinoxamine
C1114360|T201|COMP|30518-5|LNC|Cholate|Cholate
C1114361|T201|COMP|30520-1|LNC|Deoxycholate|Deoxycholate
C1114362|T201|COMP|30521-9|LNC|Inhibin B|Inhibin B
C1114363|T201|COMP|30522-7|LNC|C reactive protein|C reactive protein
C1114364|T201|COMP|30524-3|LNC|Triglyceride^post 12H CFst|Triglyceride^post 12H CFst
C1114365|T201|COMP|30525-0|LNC|Age|Age
C1114366|T201|COMP|30526-8|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C1114367|T201|COMP|30527-6|LNC|Calcium|Calcium
C1114368|T201|COMP|30529-2|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C1114369|T201|COMP|30530-0|LNC|Intrinsic factor Ab|Intrinsic factor Ab
C1114370|T201|COMP|30532-6|LNC|levoFLOXacin^peak|levoFLOXacin^peak
C1114371|T201|COMP|30533-4|LNC|levoFLOXacin^trough|levoFLOXacin^trough
C1114372|T201|COMP|30534-2|LNC|Linoleoylcarnitine (C18:2)|Linoleoylcarnitine (C18:2)
C1114373|T201|COMP|30535-9|LNC|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C1114374|T201|COMP|30538-3|LNC|Neutrophil cytoplasmic Ab.classic|Neutrophil cytoplasmic Ab.classic
C1114375|T201|COMP|30539-1|LNC|Neutrophil cytoplasmic Ab.perinuclear|Neutrophil cytoplasmic Ab.perinuclear
C1114376|T201|COMP|30540-9|LNC|Octanoylcarnitine (C8)|Octanoylcarnitine (C8)
C1114377|T201|COMP|30541-7|LNC|Octenoylcarnitine (C8:1)|Octenoylcarnitine (C8:1)
C1114378|T201|COMP|30542-5|LNC|Oleoylcarnitine (C18:1)|Oleoylcarnitine (C18:1)
C1114379|T201|COMP|30543-3|LNC|Osmotic fragility^0.75% sodium chloride|Osmotic fragility^0.75% sodium chloride
C1114380|T201|COMP|30544-1|LNC|Phosphate|Phosphate
C1114381|T201|COMP|30545-8|LNC|Platelet Ab|Platelet Ab
C1114382|T201|COMP|30547-4|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C1114383|T201|COMP|30548-2|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C1114384|T201|COMP|30549-0|LNC|Potassium|Potassium
C1114385|T201|COMP|30550-8|LNC|Pristanate/Phytanate|Pristanate/Phytanate
C1114386|T201|COMP|30551-6|LNC|Propionylcarnitine (C3)|Propionylcarnitine (C3)
C1114387|T201|COMP|30552-4|LNC|Pyridoxal phosphate|Pyridoxal phosphate
C1114388|T201|COMP|30553-2|LNC|Rabies virus Ab|Rabies virus Ab
C1114389|T201|COMP|30554-0|LNC|HIV reverse transcriptase gene mutations detected|HIV reverse transcriptase gene mutations detected
C1114390|T201|COMP|30555-7|LNC|Rickettsia typhus group Ab.IgG|Rickettsia typhus group Ab.IgG
C1114392|T201|COMP|30557-3|LNC|Smooth muscle Ab.IgG|Smooth muscle Ab.IgG
C1114393|T201|COMP|30558-1|LNC|Sodium|Sodium
C1114394|T201|COMP|30559-9|LNC|Spermatozoa Ab|Spermatozoa Ab
C1114395|T201|COMP|30560-7|LNC|Stearoylcarnitine (C18)|Stearoylcarnitine (C18)
C1114396|T201|COMP|30561-5|LNC|Streptococcus pneumoniae 6 Ab.IgG|Streptococcus pneumoniae 6 Ab.IgG
C1114397|T201|COMP|30562-3|LNC|Surfactant/Albumin|Surfactant/Albumin
C1114398|T201|COMP|30563-1|LNC|Taurine|Taurine
C1114399|T201|COMP|30564-9|LNC|Tetradecadienoylcarnitine (C14:2)|Tetradecadienoylcarnitine (C14:2)
C1114400|T201|COMP|30565-6|LNC|Tetradecanoylcarnitine (C14)|Tetradecanoylcarnitine (C14)
C1114401|T201|COMP|30566-4|LNC|Tetradecenoylcarnitine (C14:1)|Tetradecenoylcarnitine (C14:1)
C1114402|T201|COMP|30567-2|LNC|Thyroid stimulating immunoglobulins|Thyroid stimulating immunoglobulins
C1114403|T201|COMP|30568-0|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C1114404|T201|COMP|30569-8|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C1114405|T201|COMP|30570-6|LNC|Triglyceride|Triglyceride
C1114406|T201|COMP|30571-4|LNC|Vanillylmandelate/Creatinine|Vanillylmandelate/Creatinine
C1114407|T201|COMP|30574-8|LNC|Acetoacetate+Acetone|Acetoacetate+Acetone
C1114408|T201|COMP|30575-5|LNC|Xylose^baseline|Xylose^baseline
C1114409|T201|COMP|30576-3|LNC|2-Ethyl-3-Hydroxypropionate|2-Ethyl-3-Hydroxypropionate
C1114410|T201|COMP|30577-1|LNC|2-Methyl-3-Hydroxybutyrate|2-Methyl-3-Hydroxybutyrate
C1114689|T201|COMP|30894-0|LNC|Aldosterone/Renin|Aldosterone/Renin
C1114690|T201|COMP|30895-7|LNC|Renin|Renin
C1114691|T201|COMP|30896-5|LNC|Reference lab test identifier|Reference lab test identifier
C1114692|T201|COMP|30897-3|LNC|Erythrocyte volume|Erythrocyte volume
C1114693|T201|COMP|30898-1|LNC|Plasma volume|Plasma volume
C1114694|T201|COMP|30899-9|LNC|Blood volume|Blood volume
C1114695|T201|COMP|30900-5|LNC|Cold agglutinin|Cold agglutinin
C1114696|T201|COMP|30901-3|LNC|Cold agglutinin|Cold agglutinin
C1114697|T201|COMP|30902-1|LNC|Fibrinogen|Fibrinogen
C1114698|T201|COMP|30903-9|LNC|Neutrophil oxidative burst|Neutrophil oxidative burst
C1114699|T201|COMP|30904-7|LNC|Cobalamins^post dose cyanocobalamin|Cobalamins^post dose cyanocobalamin
C1114703|T201|COMP|30910-4|LNC|Antimicrobials|Antimicrobials
C1114704|T201|COMP|30912-0|LNC|DNA index|DNA index
C1114705|T201|COMP|30913-8|LNC|Cells.S phase/100 cells|Cells.S phase/100 cells
C1114706|T201|COMP|30914-6|LNC|Cells.hyperdiploid/100 cells|Cells.hyperdiploid/100 cells
C1114707|T201|COMP|30915-3|LNC|Cells.aneuploid/100 cells|Cells.aneuploid/100 cells
C1114708|T201|COMP|30917-9|LNC|DNA ploidy|DNA ploidy
C1114709|T201|COMP|30918-7|LNC|Gold|Gold
C1114710|T201|COMP|30919-5|LNC|Iron|Iron
C1114711|T201|COMP|30921-1|LNC|Mercury|Mercury
C1114712|T201|COMP|30922-9|LNC|Magnesium|Magnesium
C1114713|T201|COMP|30923-7|LNC|Chromium|Chromium
C1114714|T201|COMP|30925-2|LNC|Cadmium|Cadmium
C1114715|T201|COMP|30926-0|LNC|Aluminum|Aluminum
C1114716|T201|COMP|30927-8|LNC|Selenium|Selenium
C1114717|T201|COMP|30928-6|LNC|Silver|Silver
C1114718|T201|COMP|30930-2|LNC|Zinc|Zinc
C1114719|T201|COMP|30931-0|LNC|Lead|Lead
C1114720|T201|COMP|30933-6|LNC|Nickel|Nickel
C1114721|T201|COMP|30934-4|LNC|Natriuretic peptide.B|Natriuretic peptide.B
C1114767|T201|COMP|30983-1|LNC|Aesculus hippocastanum Ab.IgE|Aesculus hippocastanum Ab.IgE
C1114768|T201|COMP|30985-6|LNC|Betula verrucosa recombinant (rBet v) 2 Ab.IgE|Betula verrucosa recombinant (rBet v) 2 Ab.IgE
C1114770|T201|COMP|30987-2|LNC|Chinchilla epithelium Ab.IgE|Chinchilla epithelium Ab.IgE
C1114772|T201|COMP|30989-8|LNC|Sardinops melanostictus Ab.IgE|Sardinops melanostictus Ab.IgE
C1114777|T201|COMP|30994-8|LNC|Phleum pratense recombinant (rPhl p) 1 Ab.IgE|Phleum pratense recombinant (rPhl p) 1 Ab.IgE
C1114778|T201|COMP|30995-5|LNC|Phleum pratense recombinant (rPhl p) 2 Ab.IgE|Phleum pratense recombinant (rPhl p) 2 Ab.IgE
C1114779|T201|COMP|30996-3|LNC|Phleum pratense recombinant (rPhl p) 5 Ab.IgE|Phleum pratense recombinant (rPhl p) 5 Ab.IgE
C1114780|T201|COMP|30997-1|LNC|Phleum pratense native (nPhl p) 4 Ab.IgE|Phleum pratense native (nPhl p) 4 Ab.IgE
C1114781|T201|COMP|30998-9|LNC|Phleum pratense recombinant (rPhl p) 6 Ab.IgE|Phleum pratense recombinant (rPhl p) 6 Ab.IgE
C1114782|T201|COMP|30999-7|LNC|Phleum pratense recombinant (rPhl p) 7 Ab.IgE|Phleum pratense recombinant (rPhl p) 7 Ab.IgE
C1114783|T201|COMP|31000-3|LNC|Phleum pratense recombinant (rPhl p) 11 Ab.IgE|Phleum pratense recombinant (rPhl p) 11 Ab.IgE
C1114784|T201|COMP|31001-1|LNC|Parietaria judaica Ab.IgE.RAST class|Parietaria judaica Ab.IgE.RAST class
C1114785|T201|COMP|31002-9|LNC|Phoenix dactylifera Ab.IgE|Phoenix dactylifera Ab.IgE
C1114789|T201|COMP|31007-8|LNC|(Beef+Chicken meat+Pork+Turkey meat) Ab.IgE|(Beef+Chicken meat+Pork+Turkey meat) Ab.IgE
C1114793|T201|COMP|31011-0|LNC|Sardinops melanostictus Ab.IgE.RAST class|Sardinops melanostictus Ab.IgE.RAST class
C1114794|T201|COMP|31012-8|LNC|Vancomycin|Vancomycin
C1114795|T201|COMP|31013-6|LNC|DehydrochlormethylTESTOSTERone|DehydrochlormethylTESTOSTERone
C1114796|T201|COMP|31014-4|LNC|Corynebacterium diphtheriae Ab^2nd specimen|Corynebacterium diphtheriae Ab^2nd specimen
C1114797|T201|COMP|31015-1|LNC|Ethylestrenol|Ethylestrenol
C1114798|T201|COMP|31016-9|LNC|Levoamphetamine/Amphetamines.total|Levoamphetamine/Amphetamines.total
C1114799|T201|COMP|31017-7|LNC|Tissue transglutaminase Ab.IgA|Tissue transglutaminase Ab.IgA
C1114800|T201|COMP|31018-5|LNC|Haemophilus influenzae B Ab.IgG^2nd specimen|Haemophilus influenzae B Ab.IgG^2nd specimen
C1114801|T201|COMP|31019-3|LNC|10-Hydroxycarbazepine|10-Hydroxycarbazepine
C1114802|T201|COMP|31021-9|LNC|Interferon.beta 1 Ab|Interferon.beta 1 Ab
C1114803|T201|COMP|31022-7|LNC|Filaria identified|Filaria identified
C1114804|T201|COMP|31023-5|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C1114805|T201|COMP|31024-3|LNC|Voltage-gated calcium channel Ab|Voltage-gated calcium channel Ab
C1114806|T201|COMP|31026-8|LNC|Dextromethamphetamine/Amphetamines.total|Dextromethamphetamine/Amphetamines.total
C1114807|T201|COMP|31027-6|LNC|Ritonavir|Ritonavir
C1114808|T201|COMP|31028-4|LNC|Amprenavir|Amprenavir
C1114809|T201|COMP|31029-2|LNC|Stenbolone|Stenbolone
C1114810|T201|COMP|31030-0|LNC|Testosterone/Epitestosterone|Testosterone/Epitestosterone
C1114811|T201|COMP|31031-8|LNC|Saccharomyces cerevisiae Ab.IgG|Saccharomyces cerevisiae Ab.IgG
C1114812|T201|COMP|31032-6|LNC|Saccharomyces cerevisiae Ab.IgA|Saccharomyces cerevisiae Ab.IgA
C1114813|T201|COMP|31033-4|LNC|Indinavir|Indinavir
C1114815|T201|COMP|31036-7|LNC|Gatifloxacin|Gatifloxacin
C1114816|T201|COMP|31037-5|LNC|Moxifloxacin|Moxifloxacin
C1114817|T201|COMP|31039-1|LNC|Moxifloxacin|Moxifloxacin
C1114818|T201|COMP|31040-9|LNC|Gatifloxacin|Gatifloxacin
C1114819|T201|COMP|31041-7|LNC|Moxifloxacin|Moxifloxacin
C1114820|T201|COMP|31043-3|LNC|Moxifloxacin|Moxifloxacin
C1114822|T201|COMP|29782-0|LNC|Trivittatus virus Ab|Trivittatus virus Ab
C1114823|T201|COMP|29784-6|LNC|Highlands J virus Ab|Highlands J virus Ab
C1114824|T201|COMP|29788-7|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C1114825|T201|COMP|29793-7|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1114826|T201|COMP|29798-6|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C1114827|T201|COMP|29802-6|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C1114828|T201|COMP|29815-8|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C1114829|T201|COMP|29837-2|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1114830|T201|COMP|29841-4|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C1114831|T201|COMP|29845-5|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1114832|T201|COMP|29846-3|LNC|Trivittatus virus Ab|Trivittatus virus Ab
C1114833|T201|COMP|29850-5|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1114834|T201|COMP|29855-4|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1114835|T201|COMP|29863-8|LNC|IgD Ag|IgD Ag
C1114836|T201|COMP|29888-5|LNC|Pseudorabies virus.G1 gene deletion Ab|Pseudorabies virus.G1 gene deletion Ab
C1114837|T201|COMP|29903-2|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1114838|T201|COMP|29908-1|LNC|Parainfluenza virus 1 RNA|Parainfluenza virus 1 RNA
C1114839|T201|COMP|29917-2|LNC|Selenium/Creatinine|Selenium/Creatinine
C1114840|T201|COMP|29920-6|LNC|Beryllium/Creatinine|Beryllium/Creatinine
C1114841|T201|COMP|29924-8|LNC|Scandium|Scandium
C1114842|T201|COMP|29925-5|LNC|Scandium/Creatinine|Scandium/Creatinine
C1114843|T201|COMP|29953-7|LNC|Nuclear Ab|Nuclear Ab
C1114844|T201|COMP|29964-4|LNC|Sjogrens syndrome-A extractable nuclear Ab.IgG|Sjogrens syndrome-A extractable nuclear Ab.IgG
C1114845|T201|COMP|29973-5|LNC|Strontium/Creatinine|Strontium/Creatinine
C1114846|T201|COMP|29978-4|LNC|Silver/Creatinine|Silver/Creatinine
C1114847|T201|COMP|29981-8|LNC|Tin/Creatinine|Tin/Creatinine
C1114848|T201|COMP|29982-6|LNC|Cesium|Cesium
C1114849|T201|COMP|29986-7|LNC|Barium/Creatinine|Barium/Creatinine
C1114850|T201|COMP|29994-1|LNC|Basement membrane Ab.IgG|Basement membrane Ab.IgG
C1114851|T201|COMP|30015-2|LNC|Borrelia burgdorferi 41kD Ab.IgG|Borrelia burgdorferi 41kD Ab.IgG
C1114852|T201|COMP|30023-6|LNC|Bacillus subtilis Ab.IgE|Bacillus subtilis Ab.IgE
C1114853|T201|COMP|30033-5|LNC|Homocystine^6H post dose methionine|Homocystine^6H post dose methionine
C1114854|T201|COMP|30039-2|LNC|Anaplasma phagocytophilum DNA|Anaplasma phagocytophilum DNA
C1114855|T201|COMP|30044-2|LNC|Dirofilaria immitis Ab|Dirofilaria immitis Ab
C1114856|T201|COMP|30048-3|LNC|Lysine/Creatinine|Lysine/Creatinine
C1114857|T201|COMP|30051-7|LNC|Homocystine/Creatinine|Homocystine/Creatinine
C1114858|T201|COMP|30052-5|LNC|Isoleucine/Creatinine|Isoleucine/Creatinine
C1114859|T201|COMP|30056-6|LNC|Glutamine/Creatinine|Glutamine/Creatinine
C1114860|T201|COMP|30084-8|LNC|Lupus erythematosus deoxynucleoproteins Ab.IgG|Lupus erythematosus deoxynucleoproteins Ab.IgG
C1114861|T201|COMP|30093-9|LNC|Brucella canis Ab.IgM|Brucella canis Ab.IgM
C1114862|T201|COMP|30098-8|LNC|Neisseria meningitidis serogroup Y Ag|Neisseria meningitidis serogroup Y Ag
C1114863|T201|COMP|30101-0|LNC|Yersinia enterocolitica O:5 Ab|Yersinia enterocolitica O:5 Ab
C1114864|T201|COMP|30106-9|LNC|Acetylcholinesterase|Acetylcholinesterase
C1114865|T201|COMP|30110-1|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C1114866|T201|COMP|30114-3|LNC|Lymphocytes.lambda|Lymphocytes.lambda
C1114867|T201|COMP|30138-2|LNC|Epstein Barr virus nuclear Ab^2nd specimen|Epstein Barr virus nuclear Ab^2nd specimen
C1114868|T201|COMP|30149-9|LNC|Streptolysin O Ab^1st specimen|Streptolysin O Ab^1st specimen
C1114870|T201|COMP|30158-0|LNC|Toxoplasma gondii|Toxoplasma gondii
C1114871|T201|COMP|30162-2|LNC|Cynara scolymus Ab.IgG|Cynara scolymus Ab.IgG
C1114872|T201|COMP|30173-9|LNC|Cortisol.free|Cortisol.free
C1114874|T201|COMP|30205-9|LNC|Chlamydophila pneumoniae Ab|Chlamydophila pneumoniae Ab
C1114875|T201|COMP|30214-1|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C1114876|T201|COMP|30219-0|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C1114877|T201|COMP|30222-4|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C1114879|T201|COMP|30234-9|LNC|3-Hydroxypalmitoylcarnitine (C16-OH)|3-Hydroxypalmitoylcarnitine (C16-OH)
C1114880|T201|COMP|30261-2|LNC|Insulin^3.5H post XXX challenge|Insulin^3.5H post XXX challenge
C1114881|T201|COMP|30264-6|LNC|Glucose^40M post dose glucose|Glucose^40M post dose glucose
C1114882|T201|COMP|30266-1|LNC|Glucose^1.6H post dose glucose|Glucose^1.6H post dose glucose
C1114883|T201|COMP|30271-1|LNC|Zalcitabine|Zalcitabine
C1114884|T201|COMP|30276-0|LNC|Delavirdine|Delavirdine
C1114885|T201|COMP|30285-1|LNC|Zalcitabine|Zalcitabine
C1114886|T201|COMP|30315-6|LNC|Acid alpha glucosidase|Acid alpha glucosidase
C1114887|T201|COMP|30324-8|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1114888|T201|COMP|30329-7|LNC|Disialylganglioside GD1b Ab.IgG|Disialylganglioside GD1b Ab.IgG
C1114889|T201|COMP|30333-9|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C1114890|T201|COMP|30337-0|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C1114891|T201|COMP|30341-2|LNC|Erythrocyte sedimentation rate|Erythrocyte sedimentation rate
C1114892|T201|COMP|30346-1|LNC|Glucose^3H post 1.2 g/kg lactose PO|Glucose^3H post 1.2 g/kg lactose PO
C1114893|T201|COMP|30354-5|LNC|Hemoglobin|Hemoglobin
C1114894|T201|COMP|30382-6|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1114895|T201|COMP|30387-5|LNC|Erythrocytes|Erythrocytes
C1114896|T201|COMP|30390-9|LNC|Erythrocytes|Erythrocytes
C1114897|T201|COMP|30394-1|LNC|Granulocytes|Granulocytes
C1114898|T201|COMP|30399-0|LNC|Hemoglobin distribution width|Hemoglobin distribution width
C1114899|T201|COMP|30402-2|LNC|Leukocytes|Leukocytes
C1114900|T201|COMP|30406-3|LNC|Leukocytes other|Leukocytes other
C1114901|T201|COMP|30409-7|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C1114902|T201|COMP|30438-6|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1114903|T201|COMP|30446-9|LNC|Myelocytes|Myelocytes
C1114904|T201|COMP|30454-3|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C1114905|T201|COMP|30459-2|LNC|Platelet mean diameter|Platelet mean diameter
C1114906|T201|COMP|26524-9|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C1114907|T201|COMP|30469-1|LNC|Unspecified cells/100 leukocytes|Unspecified cells/100 leukocytes
C1114908|T201|COMP|30473-3|LNC|Glutaconate|Glutaconate
C1114909|T201|COMP|30474-1|LNC|Glutarate|Glutarate
C1114910|T201|COMP|30477-4|LNC|Hexanoylglycine|Hexanoylglycine
C1114912|T201|COMP|30514-4|LNC|Tetrahydrocortisone/Creatinine|Tetrahydrocortisone/Creatinine
C1114913|T201|COMP|30519-3|LNC|Chenodeoxycholate|Chenodeoxycholate
C1114914|T201|COMP|30523-5|LNC|Mycobacterium sp DNA|Mycobacterium sp DNA
C1114915|T201|COMP|30528-4|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C1114916|T201|COMP|30531-8|LNC|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)
C1114917|T201|COMP|30536-7|LNC|Magnesium|Magnesium
C1114918|T201|COMP|30537-5|LNC|Myocardium Ab|Myocardium Ab
C1114919|T201|COMP|30546-6|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C1114920|T201|COMP|30572-2|LNC|Pyridoxal|Pyridoxal
C1114958|T201|COMP|30911-2|LNC|DNA ploidy|DNA ploidy
C1114959|T201|COMP|30916-1|LNC|Cells.euploid+Cells.aneuploid/100 cells|Cells.euploid+Cells.aneuploid/100 cells
C1114960|T201|COMP|30920-3|LNC|Copper|Copper
C1114961|T201|COMP|30924-5|LNC|Arsenic|Arsenic
C1114962|T201|COMP|30929-4|LNC|Thallium|Thallium
C1114963|T201|COMP|30932-8|LNC|Manganese|Manganese
C1114965|T201|COMP|30984-9|LNC|Betula verrucosa recombinant (rBet v) 1 Ab.IgE|Betula verrucosa recombinant (rBet v) 1 Ab.IgE
C1114967|T201|COMP|31020-1|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C1114968|T201|COMP|31025-0|LNC|Dextroamphetamine/Amphetamines.total|Dextroamphetamine/Amphetamines.total
C1114970|T201|COMP|31038-3|LNC|Gatifloxacin|Gatifloxacin
C1114971|T201|COMP|31042-5|LNC|Gatifloxacin|Gatifloxacin
C1116460|T201|COMP|29912-3|LNC|Magnesium|Magnesium
C1116461|T201|COMP|30028-5|LNC|O-Ethyl O-(p-nitrophenyl) phenylphosphonothionate|O-Ethyl O-(p-nitrophenyl) phenylphosphonothionate
C1116463|T201|COMP|30280-2|LNC|Nelfinavir|Nelfinavir
C1116464|T201|COMP|30410-5|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C1116470|T201|COMP|30082-2|LNC|IgE|IgE
C1116519|T201|COMP|30348-7|LNC|Glutamate|Glutamate
C1141680|T201|COMP|23515-0|LNC|Trypanosoma equiperdum Ab|Trypanosoma equiperdum Ab
C1145645|T201|COMP|2703-7|LNC|Oxygen|Oxygen
C1145646|T201|COMP|2704-5|LNC|Oxygen|Oxygen
C1145647|T201|COMP|2705-2|LNC|Oxygen|Oxygen
C1145648|T201|COMP|3394-4|LNC|Benzoylecgonine|Benzoylecgonine
C1145649|T201|COMP|6584-7|LNC|Virus identified|Virus identified
C1145650|T201|COMP|580-1|LNC|Fungus identified|Fungus identified
C1145651|T201|COMP|602-3|LNC|Bacteria identified|Bacteria identified
C1145652|T201|COMP|603-1|LNC|Bacteria identified|Bacteria identified
C1145653|T201|COMP|616-3|LNC|Bacteria identified|Bacteria identified
C1145654|T201|COMP|619-7|LNC|Bacteria identified|Bacteria identified
C1145655|T201|COMP|622-1|LNC|Bacteria identified|Bacteria identified
C1145656|T201|COMP|625-4|LNC|Bacteria identified|Bacteria identified
C1145657|T201|COMP|627-0|LNC|Bacteria identified|Bacteria identified
C1145658|T201|COMP|628-8|LNC|Bacteria identified|Bacteria identified
C1145704|T201|COMP|17876-4|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1145705|T201|COMP|17875-6|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1145706|T201|COMP|17874-9|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1145707|T201|COMP|17873-1|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1145708|T201|COMP|17940-8|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1145709|T201|COMP|17939-0|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1145710|T201|COMP|17938-2|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1145711|T201|COMP|17937-4|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1145712|T201|COMP|5074-0|LNC|Candida albicans Ab|Candida albicans Ab
C1145715|T201|COMP|13445-2|LNC|Creatinine renal clearance/1.73 sq M|Creatinine renal clearance/1.73 sq M
C1145716|T201|COMP|12195-4|LNC|Creatinine renal clearance/1.73 sq M|Creatinine renal clearance/1.73 sq M
C1145717|T201|COMP|17948-1|LNC|Fungus identified^^^3|Fungus identified^^^3
C1145718|T201|COMP|17947-3|LNC|Fungus identified^^^2|Fungus identified^^^2
C1145719|T201|COMP|17886-3|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1145720|T201|COMP|17885-5|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1145721|T201|COMP|17884-8|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1145722|T201|COMP|17883-0|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1145723|T201|COMP|10352-3|LNC|Bacteria identified|Bacteria identified
C1145724|T201|COMP|17891-3|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1145725|T201|COMP|17890-5|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1145726|T201|COMP|17889-7|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1145727|T201|COMP|17888-9|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1145728|T201|COMP|10353-1|LNC|Bacteria identified|Bacteria identified
C1145729|T201|COMP|17962-2|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1145730|T201|COMP|17961-4|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1145731|T201|COMP|17960-6|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1145732|T201|COMP|17959-8|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1145733|T201|COMP|17896-2|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1145734|T201|COMP|17895-4|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1145735|T201|COMP|17894-7|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1145736|T201|COMP|17893-9|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1146730|T201|COMP|31045-8|LNC|Creatinine/Urea nitrogen|Creatinine/Urea nitrogen
C1146731|T201|COMP|31046-6|LNC|Rheumatoid factor|Rheumatoid factor
C1146732|T201|COMP|31047-4|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C1146733|T201|COMP|31048-2|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C1146734|T201|COMP|31049-0|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C1146735|T201|COMP|31050-8|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C1146736|T201|COMP|31051-6|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C1146737|T201|COMP|31052-4|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C1146738|T201|COMP|31053-2|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C1146739|T201|COMP|31054-0|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C1146740|T201|COMP|31055-7|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C1146741|T201|COMP|31056-5|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C1146742|T201|COMP|31057-3|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C1146743|T201|COMP|31058-1|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C1146744|T201|COMP|31059-9|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C1146745|T201|COMP|31060-7|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C1146746|T201|COMP|31061-5|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C1146747|T201|COMP|31062-3|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C1146748|T201|COMP|31063-1|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C1146749|T201|COMP|31064-9|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C1146750|T201|COMP|31065-6|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C1146751|T201|COMP|31066-4|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C1146752|T201|COMP|31067-2|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C1146753|T201|COMP|31068-0|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C1146754|T201|COMP|31069-8|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C1146755|T201|COMP|31070-6|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C1146756|T201|COMP|31071-4|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C1146757|T201|COMP|31072-2|LNC|HIV 1 p41 Ab|HIV 1 p41 Ab
C1146758|T201|COMP|31073-0|LNC|HIV 2 Ab band pattern|HIV 2 Ab band pattern
C1146759|T201|COMP|31074-8|LNC|Cells.CD30|Cells.CD30
C1146760|T201|COMP|31075-5|LNC|Legionella pneumophila 1 Ab.IgM|Legionella pneumophila 1 Ab.IgM
C1146761|T201|COMP|31076-3|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C1146762|T201|COMP|31077-1|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C1146763|T201|COMP|31078-9|LNC|Casuarina equisetifolia Ab.IgE.RAST class|Casuarina equisetifolia Ab.IgE.RAST class
C1146764|T201|COMP|31079-7|LNC|Gerbil epithelium Ab.IgE.RAST class|Gerbil epithelium Ab.IgE.RAST class
C1146765|T201|COMP|31080-5|LNC|Cannabinoids|Cannabinoids
C1146766|T201|COMP|31081-3|LNC|Benzodiazepines|Benzodiazepines
C1146767|T201|COMP|31082-1|LNC|Ethylene glycol|Ethylene glycol
C1146768|T201|COMP|31083-9|LNC|Lead|Lead
C1146769|T201|COMP|31084-7|LNC|Methadone|Methadone
C1146770|T201|COMP|31085-4|LNC|Methaqualone|Methaqualone
C1146771|T201|COMP|31086-2|LNC|Morphine.free|Morphine.free
C1146772|T201|COMP|31087-0|LNC|Thioridazine|Thioridazine
C1146773|T201|COMP|31088-8|LNC|Narcotics|Narcotics
C1146774|T201|COMP|31089-6|LNC|Acetaminophen|Acetaminophen
C1146775|T201|COMP|31090-4|LNC|Ethchlorvynol|Ethchlorvynol
C1146776|T201|COMP|31091-2|LNC|Gentamicin^peak post extended interval dosing|Gentamicin^peak post extended interval dosing
C1146777|T201|COMP|31092-0|LNC|Gentamicin^trough post extended interval dosing|Gentamicin^trough post extended interval dosing
C1146778|T201|COMP|31093-8|LNC|Gentamicin^random post extended interval dosing|Gentamicin^random post extended interval dosing
C1146779|T201|COMP|31094-6|LNC|Tobramycin^peak post extended interval dosing|Tobramycin^peak post extended interval dosing
C1146780|T201|COMP|31095-3|LNC|Tobramycin^trough post extended interval dosing|Tobramycin^trough post extended interval dosing
C1146781|T201|COMP|31096-1|LNC|Tobramycin^random post extended interval dosing|Tobramycin^random post extended interval dosing
C1146782|T201|COMP|31097-9|LNC|Amikacin^peak post extended interval dosing|Amikacin^peak post extended interval dosing
C1146783|T201|COMP|31098-7|LNC|Amikacin^trough post extended interval dosing|Amikacin^trough post extended interval dosing
C1146784|T201|COMP|31099-5|LNC|Amikacin^random post extended interval dosing|Amikacin^random post extended interval dosing
C1146785|T201|COMP|31100-1|LNC|Hematocrit|Hematocrit
C1146786|T201|COMP|31101-9|LNC|Creatinine|Creatinine
C1146787|T201|COMP|31102-7|LNC|Protein S actual/Normal|Protein S actual/Normal
C1146797|T201|COMP|31112-6|LNC|Reticulocytes/100 erythrocytes|Reticulocytes/100 erythrocytes
C1146798|T201|COMP|33617-2|LNC|Cells.HLA-DR+|Cells.HLA-DR+
C1146799|T201|COMP|31114-2|LNC|Cells.aneuploid.population 1/100 cells|Cells.aneuploid.population 1/100 cells
C1146800|T201|COMP|31115-9|LNC|Cells.aneuploid.population 2/100 cells|Cells.aneuploid.population 2/100 cells
C1146803|T201|COMP|31118-3|LNC|Cells.G2+M phase/100 cells|Cells.G2+M phase/100 cells
C1146804|T201|COMP|31119-1|LNC|Cells.CD227/100 cells|Cells.CD227/100 cells
C1146805|T201|COMP|31120-9|LNC|Cells.CD227|Cells.CD227
C1146806|T201|COMP|17221-3|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C1146807|T201|COMP|31122-5|LNC|Cells.CD235a|Cells.CD235a
C1146808|T201|COMP|31123-3|LNC|Cells.CD25|Cells.CD25
C1146809|T201|COMP|31124-1|LNC|Cells.CD20+CD25+/100 cells|Cells.CD20+CD25+/100 cells
C1146810|T201|COMP|31125-8|LNC|Cells.CD20+CD25+|Cells.CD20+CD25+
C1146811|T201|COMP|31126-6|LNC|Cells.CD20+CD25-/100 cells|Cells.CD20+CD25-/100 cells
C1146812|T201|COMP|31127-4|LNC|Cells.CD20+CD25-|Cells.CD20+CD25-
C1146813|T201|COMP|31128-2|LNC|Cells.CD11c-CD20+/100 cells|Cells.CD11c-CD20+/100 cells
C1146814|T201|COMP|31129-0|LNC|Cells.CD11c-CD20+|Cells.CD11c-CD20+
C1146815|T201|COMP|31130-8|LNC|Mumps virus soluble Ab|Mumps virus soluble Ab
C1146816|T201|COMP|31131-6|LNC|Mumps virus particle-bound Ab|Mumps virus particle-bound Ab
C1146817|T201|COMP|31132-4|LNC|Mumps virus soluble Ab|Mumps virus soluble Ab
C1146818|T201|COMP|31133-2|LNC|Mumps virus particle-bound Ab|Mumps virus particle-bound Ab
C1146819|T201|COMP|31134-0|LNC|Nuclear matrix protein 22|Nuclear matrix protein 22
C1146820|T201|COMP|31135-7|LNC|Cocaethylene|Cocaethylene
C1146821|T201|COMP|31136-5|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C1146822|T201|COMP|31137-3|LNC|Cocaine|Cocaine
C1146823|T201|COMP|31138-1|LNC|Cefotaxime|Cefotaxime
C1146824|T201|COMP|31139-9|LNC|Cefotaxime|Cefotaxime
C1146825|T201|COMP|31140-7|LNC|cefTRIAXone|cefTRIAXone
C1146826|T201|COMP|31141-5|LNC|cefTRIAXone|cefTRIAXone
C1146827|T201|COMP|31142-3|LNC|Cefepime|Cefepime
C1146828|T201|COMP|31143-1|LNC|Cefepime|Cefepime
C1146829|T201|COMP|31144-9|LNC|Thyroxine|Thyroxine
C1146830|T201|COMP|31145-6|LNC|Thyroxine|Thyroxine
C1146831|T201|COMP|31146-4|LNC|Reagin Ab|Reagin Ab
C1146832|T201|COMP|31147-2|LNC|Reagin Ab|Reagin Ab
C1146833|T201|COMP|31148-0|LNC|Heavy metals|Heavy metals
C1146834|T201|COMP|31149-8|LNC|P53 protein Ag/100 cells|P53 protein Ag/100 cells
C1146835|T201|COMP|31150-6|LNC|HER2|HER2
C1146836|T201|COMP|31151-4|LNC|Alpha-2-Microglobulin|Alpha-2-Microglobulin
C1146837|T201|COMP|31152-2|LNC|Immunoglobulin light chains|Immunoglobulin light chains
C1146838|T201|COMP|31153-0|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1146839|T201|COMP|31154-8|LNC|Coccidioides sp Ab.IgG|Coccidioides sp Ab.IgG
C1146840|T201|COMP|31155-5|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C1146841|T201|COMP|31156-3|LNC|Hemoglobin Barts/Hemoglobin.total|Hemoglobin Barts/Hemoglobin.total
C1146842|T201|COMP|31157-1|LNC|Carboxyhemoglobin|Carboxyhemoglobin
C1146843|T201|COMP|31158-9|LNC|Fibrinogen Ag/Fibrinogen|Fibrinogen Ag/Fibrinogen
C1146844|T201|COMP|31159-7|LNC|Heparin anti Xa|Heparin anti Xa
C1146845|T201|COMP|31160-5|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C1146847|T201|COMP|31162-1|LNC|Sulfate-3-Glucuronyl paragloboside Ab|Sulfate-3-Glucuronyl paragloboside Ab
C1146848|T201|COMP|31163-9|LNC|Ganglioside GD1b Ab|Ganglioside GD1b Ab
C1146849|T201|COMP|31164-7|LNC|Ganglioside GQ1b Ab|Ganglioside GQ1b Ab
C1146850|T201|COMP|31165-4|LNC|Methyl butyl ketone|Methyl butyl ketone
C1146851|T201|COMP|31166-2|LNC|Methyl isoamyl ketone|Methyl isoamyl ketone
C1146852|T201|COMP|31167-0|LNC|Methyl propyl ketone|Methyl propyl ketone
C1146853|T201|COMP|31168-8|LNC|Mesityl oxide|Mesityl oxide
C1146854|T201|COMP|31169-6|LNC|Theobromine|Theobromine
C1146855|T201|COMP|31170-4|LNC|2,5-Hexanedione|2,5-Hexanedione
C1146856|T201|COMP|31171-2|LNC|2,5-Hexanedione/Creatinine|2,5-Hexanedione/Creatinine
C1146857|T201|COMP|31172-0|LNC|Fonofos|Fonofos
C1146858|T201|COMP|31173-8|LNC|Mevinphos|Mevinphos
C1146859|T201|COMP|31174-6|LNC|Terbufos|Terbufos
C1146860|T201|COMP|31175-3|LNC|Metasystox|Metasystox
C1146861|T201|COMP|31176-1|LNC|Estradiol|Estradiol
C1146862|T201|COMP|31177-9|LNC|Estrone|Estrone
C1146863|T201|COMP|31178-7|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C1146864|T201|COMP|31179-5|LNC|Lopinavir|Lopinavir
C1146865|T201|COMP|31180-3|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C1146866|T201|COMP|31181-1|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C1146867|T201|COMP|31182-9|LNC|7-Aminonitrazepam|7-Aminonitrazepam
C1146868|T201|COMP|31183-7|LNC|Streptococcus pneumoniae 5 Ab.IgG|Streptococcus pneumoniae 5 Ab.IgG
C1146869|T201|COMP|31184-5|LNC|Methyl amyl ketone|Methyl amyl ketone
C1146870|T201|COMP|31185-2|LNC|Platelet Ab.IgA|Platelet Ab.IgA
C1146871|T201|COMP|31186-0|LNC|Platelet Ab.IgM|Platelet Ab.IgM
C1146885|T201|COMP|31200-9|LNC|Histoplasma capsulatum Ab.IgG|Histoplasma capsulatum Ab.IgG
C1146886|T201|COMP|31201-7|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C1146887|T201|COMP|31202-5|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C1146888|T201|COMP|31203-3|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C1146889|T201|COMP|31204-1|LNC|Hepatitis B virus core Ab.IgM|Hepatitis B virus core Ab.IgM
C1146892|T201|COMP|31207-4|LNC|Progesterone receptor|Progesterone receptor
C1146893|T201|COMP|31208-2|LNC|Specimen source|Specimen source
C1146894|T201|COMP|31209-0|LNC|Islet cell 512 Ab|Islet cell 512 Ab
C1146897|T201|COMP|31212-4|LNC|Actinobacillus pleuropneumoniae serotype 1 Ab|Actinobacillus pleuropneumoniae serotype 1 Ab
C1146898|T201|COMP|31213-2|LNC|Actinobacillus pleuropneumoniae serotype 3 Ab|Actinobacillus pleuropneumoniae serotype 3 Ab
C1146899|T201|COMP|31214-0|LNC|Actinobacillus pleuropneumoniae serotype 5 Ab|Actinobacillus pleuropneumoniae serotype 5 Ab
C1146900|T201|COMP|31215-7|LNC|Actinobacillus pleuropneumoniae serotype 7 Ab|Actinobacillus pleuropneumoniae serotype 7 Ab
C1146901|T201|COMP|31216-5|LNC|Actinobacillus pleuropneumoniae Ab|Actinobacillus pleuropneumoniae Ab
C1146902|T201|COMP|31217-3|LNC|Adenovirus Ab|Adenovirus Ab
C1146903|T201|COMP|31218-1|LNC|Afipia felis Ab.IgG|Afipia felis Ab.IgG
C1146904|T201|COMP|31219-9|LNC|Afipia felis Ab.IgM|Afipia felis Ab.IgM
C1146905|T201|COMP|31220-7|LNC|African horse sickness virus Ab|African horse sickness virus Ab
C1146906|T201|COMP|31221-5|LNC|Alcelaphine herpesvirus 1 Ab|Alcelaphine herpesvirus 1 Ab
C1146907|T201|COMP|31222-3|LNC|Anaplasma marginale Ab|Anaplasma marginale Ab
C1146908|T201|COMP|31223-1|LNC|Arbovirus NOS Ab|Arbovirus NOS Ab
C1146909|T201|COMP|31224-9|LNC|Ascaris sp Ab|Ascaris sp Ab
C1146910|T201|COMP|31225-6|LNC|Asialoganglioside GM1 Ab|Asialoganglioside GM1 Ab
C1146911|T201|COMP|31226-4|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C1146912|T201|COMP|31227-2|LNC|Asialoganglioside GM1 Ab.IgM|Asialoganglioside GM1 Ab.IgM
C1146913|T201|COMP|31228-0|LNC|Aspergillus clavatus Ab|Aspergillus clavatus Ab
C1146914|T201|COMP|31229-8|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C1146915|T201|COMP|31230-6|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C1146916|T201|COMP|31231-4|LNC|Aspergillus nidulans Ab|Aspergillus nidulans Ab
C1146917|T201|COMP|31232-2|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C1146918|T201|COMP|31233-0|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C1146919|T201|COMP|31234-8|LNC|Aspergillus terreus Ab|Aspergillus terreus Ab
C1146920|T201|COMP|31235-5|LNC|Aureobasidium pullulans Ab.IgG|Aureobasidium pullulans Ab.IgG
C1146921|T201|COMP|31236-3|LNC|Infectious bronchitis virus Ab|Infectious bronchitis virus Ab
C1146922|T201|COMP|31237-1|LNC|Infectious bronchitis virus Ark-99 Ab|Infectious bronchitis virus Ark-99 Ab
C1146923|T201|COMP|31238-9|LNC|Infectious bronchitis virus Conn-42 Ab|Infectious bronchitis virus Conn-42 Ab
C1146924|T201|COMP|31239-7|LNC|Infectious bronchitis virus Mass-41 Ab|Infectious bronchitis virus Mass-41 Ab
C1146925|T201|COMP|31240-5|LNC|Avian infectious laryngotracheitis virus Ab|Avian infectious laryngotracheitis virus Ab
C1146926|T201|COMP|31241-3|LNC|Influenza virus A Ab|Influenza virus A Ab
C1146927|T201|COMP|31242-1|LNC|Avian paramyxovirus 1 Ab|Avian paramyxovirus 1 Ab
C1146928|T201|COMP|31243-9|LNC|Avian paramyxovirus 2 Ab|Avian paramyxovirus 2 Ab
C1146929|T201|COMP|31244-7|LNC|Babesia microti Ab.IgG|Babesia microti Ab.IgG
C1146930|T201|COMP|31245-4|LNC|Babesia microti Ab.IgM|Babesia microti Ab.IgM
C1146931|T201|COMP|31246-2|LNC|Babesia sp Ab.IgG|Babesia sp Ab.IgG
C1146932|T201|COMP|31247-0|LNC|Barmah forest virus Ab.IgG|Barmah forest virus Ab.IgG
C1146933|T201|COMP|31248-8|LNC|Barmah forest virus Ab.IgM|Barmah forest virus Ab.IgM
C1146934|T201|COMP|31249-6|LNC|Bartonella henselae Ab|Bartonella henselae Ab
C1146935|T201|COMP|31250-4|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C1146936|T201|COMP|31251-2|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C1146937|T201|COMP|31252-0|LNC|Basement membrane Ab|Basement membrane Ab
C1146938|T201|COMP|31253-8|LNC|Basement membrane Ab.IgA|Basement membrane Ab.IgA
C1146939|T201|COMP|31254-6|LNC|Basement membrane Ab.IgG|Basement membrane Ab.IgG
C1146940|T201|COMP|31255-3|LNC|Basement membrane Ab.IgG|Basement membrane Ab.IgG
C1146941|T201|COMP|31256-1|LNC|Beta 2 glycoprotein 1 Ab|Beta 2 glycoprotein 1 Ab
C1146942|T201|COMP|31257-9|LNC|Beta tubulin Ab.IgG|Beta tubulin Ab.IgG
C1146943|T201|COMP|31258-7|LNC|Beta tubulin Ab.IgM|Beta tubulin Ab.IgM
C1146944|T201|COMP|31259-5|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C1146945|T201|COMP|31260-3|LNC|Bluetongue virus 10 Ab|Bluetongue virus 10 Ab
C1146946|T201|COMP|31261-1|LNC|Bluetongue virus 11 Ab|Bluetongue virus 11 Ab
C1146947|T201|COMP|31262-9|LNC|Bluetongue virus 13 Ab|Bluetongue virus 13 Ab
C1146948|T201|COMP|31263-7|LNC|Bluetongue virus 17 Ab|Bluetongue virus 17 Ab
C1146949|T201|COMP|31264-5|LNC|Bluetongue virus 2 Ab|Bluetongue virus 2 Ab
C1146950|T201|COMP|31265-2|LNC|Bordetella avium Ab|Bordetella avium Ab
C1146951|T201|COMP|31266-0|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C1146952|T201|COMP|31267-8|LNC|Bordetella pertussis.secretory Ab.IgA|Bordetella pertussis.secretory Ab.IgA
C1146953|T201|COMP|31268-6|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C1146954|T201|COMP|31269-4|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C1146955|T201|COMP|31270-2|LNC|Bovine diarrhea virus 1 Ab|Bovine diarrhea virus 1 Ab
C1146956|T201|COMP|31271-0|LNC|Bovine diarrhea virus 2 Ab|Bovine diarrhea virus 2 Ab
C1146957|T201|COMP|31272-8|LNC|Bovine diarrhea virus Ab|Bovine diarrhea virus Ab
C1146958|T201|COMP|31273-6|LNC|Bovine herpesvirus 1 Ab|Bovine herpesvirus 1 Ab
C1146959|T201|COMP|31274-4|LNC|Bovine leukemia virus Ab|Bovine leukemia virus Ab
C1146960|T201|COMP|31275-1|LNC|Brush border Ab|Brush border Ab
C1146961|T201|COMP|31276-9|LNC|Burkholderia pseudomallei Ab.IgG|Burkholderia pseudomallei Ab.IgG
C1146962|T201|COMP|31277-7|LNC|Burkholderia pseudomallei Ab.IgM|Burkholderia pseudomallei Ab.IgM
C1146963|T201|COMP|31278-5|LNC|Campylobacter fetus Ab|Campylobacter fetus Ab
C1146964|T201|COMP|31279-3|LNC|Campylobacter jejuni Ab|Campylobacter jejuni Ab
C1146965|T201|COMP|31280-1|LNC|Canary serum proteins Ab|Canary serum proteins Ab
C1146966|T201|COMP|31281-9|LNC|Cancer associated retinopathy Ab|Cancer associated retinopathy Ab
C1146967|T201|COMP|31282-7|LNC|Canine adenovirus 1 Ab|Canine adenovirus 1 Ab
C1146968|T201|COMP|31283-5|LNC|Canine coronavirus Ab|Canine coronavirus Ab
C1146969|T201|COMP|31284-3|LNC|Canine distemper virus Ab|Canine distemper virus Ab
C1146970|T201|COMP|31285-0|LNC|Canine distemper virus Ab|Canine distemper virus Ab
C1146971|T201|COMP|31286-8|LNC|Canine parvovirus Ab|Canine parvovirus Ab
C1146972|T201|COMP|31287-6|LNC|Canine parvovirus Ab|Canine parvovirus Ab
C1146973|T201|COMP|31288-4|LNC|Canine parvovirus Ab.IgG|Canine parvovirus Ab.IgG
C1146974|T201|COMP|31289-2|LNC|Canine parvovirus Ab.IgM|Canine parvovirus Ab.IgM
C1146975|T201|COMP|31290-0|LNC|Centromere Ab.IgG|Centromere Ab.IgG
C1146976|T201|COMP|31291-8|LNC|Chicken serum Ab|Chicken serum Ab
C1146977|T201|COMP|31292-6|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C1146978|T201|COMP|31293-4|LNC|Chlamydia trachomatis Ab.IgA|Chlamydia trachomatis Ab.IgA
C1146979|T201|COMP|31294-2|LNC|Chlamydia trachomatis B Ab.IgA|Chlamydia trachomatis B Ab.IgA
C1146980|T201|COMP|31295-9|LNC|Chlamydia trachomatis B Ab.IgM|Chlamydia trachomatis B Ab.IgM
C1146981|T201|COMP|31296-7|LNC|Chlamydia trachomatis D+K Ab.IgA|Chlamydia trachomatis D+K Ab.IgA
C1146982|T201|COMP|31297-5|LNC|Chlamydia trachomatis D+K Ab.IgG|Chlamydia trachomatis D+K Ab.IgG
C1146983|T201|COMP|31298-3|LNC|Chlamydia trachomatis D+K Ab.IgM|Chlamydia trachomatis D+K Ab.IgM
C1146984|T201|COMP|31299-1|LNC|Chlamydophila pneumoniae Ab.IgA|Chlamydophila pneumoniae Ab.IgA
C1146985|T201|COMP|31300-7|LNC|Chlamydophila pneumoniae Ab.IgA|Chlamydophila pneumoniae Ab.IgA
C1146986|T201|COMP|31301-5|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C1146987|T201|COMP|31302-3|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C1146988|T201|COMP|31303-1|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C1146989|T201|COMP|31304-9|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C1146990|T201|COMP|31305-6|LNC|Chlamydophila psittaci Ab.IgA|Chlamydophila psittaci Ab.IgA
C1146991|T201|COMP|31306-4|LNC|Chlamydophila psittaci Ab.IgA|Chlamydophila psittaci Ab.IgA
C1146992|T201|COMP|31307-2|LNC|Chlamydophila psittaci Ab.IgG|Chlamydophila psittaci Ab.IgG
C1146993|T201|COMP|31308-0|LNC|Clostridioides difficile Ab|Clostridioides difficile Ab
C1146994|T201|COMP|31309-8|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C1146995|T201|COMP|31310-6|LNC|Cockatiel droppings Ab|Cockatiel droppings Ab
C1146996|T201|COMP|31311-4|LNC|Coxiella burnetii phase 1 Ab|Coxiella burnetii phase 1 Ab
C1146997|T201|COMP|31312-2|LNC|Coxiella burnetii phase 1 Ab.IgA|Coxiella burnetii phase 1 Ab.IgA
C1146998|T201|COMP|31313-0|LNC|Coxiella burnetii phase 2 Ab|Coxiella burnetii phase 2 Ab
C1146999|T201|COMP|31314-8|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C1147000|T201|COMP|31315-5|LNC|Coxiella burnetii phase 2 Ab.IgM|Coxiella burnetii phase 2 Ab.IgM
C1147001|T201|COMP|31316-3|LNC|Coxiella burnetii phase 2 Ab.IgA|Coxiella burnetii phase 2 Ab.IgA
C1147002|T201|COMP|31317-1|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C1147003|T201|COMP|31318-9|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C1147004|T201|COMP|31319-7|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C1147005|T201|COMP|31320-5|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C1147006|T201|COMP|31321-3|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C1147007|T201|COMP|31322-1|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C1147008|T201|COMP|31323-9|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C1147009|T201|COMP|31324-7|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C1147010|T201|COMP|31325-4|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C1147011|T201|COMP|31326-2|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C1147012|T201|COMP|31327-0|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C1147013|T201|COMP|31328-8|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C1147014|T201|COMP|31329-6|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C1147015|T201|COMP|31330-4|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C1147016|T201|COMP|31331-2|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C1147017|T201|COMP|31332-0|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C1147018|T201|COMP|31333-8|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C1147019|T201|COMP|31334-6|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C1147020|T201|COMP|31335-3|LNC|Cryptococcus sp Ab|Cryptococcus sp Ab
C1147021|T201|COMP|31336-1|LNC|Cryptostroma corticale Ab|Cryptostroma corticale Ab
C1147022|T201|COMP|31337-9|LNC|Cytotoxic percent reactive Ab|Cytotoxic percent reactive Ab
C1147023|T201|COMP|31338-7|LNC|Dengue virus 1 Ab|Dengue virus 1 Ab
C1147024|T201|COMP|31339-5|LNC|Dengue virus 2 Ab|Dengue virus 2 Ab
C1147025|T201|COMP|31340-3|LNC|Dengue virus 3 Ab|Dengue virus 3 Ab
C1147026|T201|COMP|31341-1|LNC|Dengue virus 4 Ab|Dengue virus 4 Ab
C1147027|T201|COMP|31342-9|LNC|Dengue virus Ab|Dengue virus Ab
C1147028|T201|COMP|31343-7|LNC|Dengue virus Ab|Dengue virus Ab
C1147029|T201|COMP|31344-5|LNC|Ganglioside GD1a Ab|Ganglioside GD1a Ab
C1147030|T201|COMP|31345-2|LNC|Ganglioside GD1b Ab|Ganglioside GD1b Ab
C1147031|T201|COMP|31346-0|LNC|Ganglioside GD1b Ab.IgG|Ganglioside GD1b Ab.IgG
C1147032|T201|COMP|31347-8|LNC|Ganglioside GD1b Ab.IgM|Ganglioside GD1b Ab.IgM
C1147033|T201|COMP|31348-6|LNC|DNA double strand Ab|DNA double strand Ab
C1147034|T201|COMP|31349-4|LNC|Eastern equine encephalomyelitis virus Ab|Eastern equine encephalomyelitis virus Ab
C1147035|T201|COMP|31350-2|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C1147036|T201|COMP|31351-0|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C1147037|T201|COMP|31352-8|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C1147038|T201|COMP|31353-6|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C1147039|T201|COMP|31354-4|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C1147040|T201|COMP|31355-1|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C1147041|T201|COMP|31356-9|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C1147042|T201|COMP|31357-7|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C1147043|T201|COMP|31358-5|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C1147044|T201|COMP|31359-3|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C1147045|T201|COMP|31360-1|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C1147046|T201|COMP|31361-9|LNC|Ehrlichia canis Ab|Ehrlichia canis Ab
C1147047|T201|COMP|31362-7|LNC|Ehrlichia chaffeensis Ab.IgM|Ehrlichia chaffeensis Ab.IgM
C1147048|T201|COMP|31363-5|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C1147049|T201|COMP|31364-3|LNC|Encephalomyocarditis virus Ab|Encephalomyocarditis virus Ab
C1147050|T201|COMP|31365-0|LNC|Endomysium Ab|Endomysium Ab
C1147051|T201|COMP|31366-8|LNC|Endomysium Ab.IgA|Endomysium Ab.IgA
C1147052|T201|COMP|31367-6|LNC|Enterovirus NOS Ab|Enterovirus NOS Ab
C1147053|T201|COMP|31368-4|LNC|Epidermis Ab|Epidermis Ab
C1147054|T201|COMP|31369-2|LNC|Epstein Barr virus capsid Ab.IgA|Epstein Barr virus capsid Ab.IgA
C1147055|T201|COMP|31370-0|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C1147056|T201|COMP|31371-8|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C1147057|T201|COMP|31372-6|LNC|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C1147058|T201|COMP|31373-4|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C1147059|T201|COMP|31374-2|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C1147060|T201|COMP|31375-9|LNC|Epstein Barr virus nuclear Ab.IgM|Epstein Barr virus nuclear Ab.IgM
C1147061|T201|COMP|31376-7|LNC|Equine arteritis virus Ab|Equine arteritis virus Ab
C1147062|T201|COMP|31377-5|LNC|Equine herpesvirus 1 Ab|Equine herpesvirus 1 Ab
C1147063|T201|COMP|31378-3|LNC|Equine herpesvirus 1+4 Ab|Equine herpesvirus 1+4 Ab
C1147064|T201|COMP|31379-1|LNC|Equine influenza virus A1 Ab|Equine influenza virus A1 Ab
C1147065|T201|COMP|31380-9|LNC|Equine influenza virus A2 Ab|Equine influenza virus A2 Ab
C1147066|T201|COMP|31381-7|LNC|Escherichia coli verotoxin 1 Ab|Escherichia coli verotoxin 1 Ab
C1147067|T201|COMP|31382-5|LNC|Escherichia coli verotoxin 2 Ab|Escherichia coli verotoxin 2 Ab
C1147068|T201|COMP|31383-3|LNC|European tick borne encephalitis virus Ab|European tick borne encephalitis virus Ab
C1147069|T201|COMP|31384-1|LNC|Feline calicivirus Ab|Feline calicivirus Ab
C1147070|T201|COMP|31385-8|LNC|Feline coronavirus Ab|Feline coronavirus Ab
C1147071|T201|COMP|31386-6|LNC|Feline herpesvirus 1 Ab|Feline herpesvirus 1 Ab
C1147072|T201|COMP|31387-4|LNC|Feline herpesvirus Ab|Feline herpesvirus Ab
C1147073|T201|COMP|31388-2|LNC|Feline immunodeficiency virus Ab|Feline immunodeficiency virus Ab
C1147074|T201|COMP|31389-0|LNC|Feline leukemia virus Ab|Feline leukemia virus Ab
C1147075|T201|COMP|31390-8|LNC|Feline panleukopenia virus Ab|Feline panleukopenia virus Ab
C1147076|T201|COMP|31391-6|LNC|Feline panleukopenia virus Ab.IgG|Feline panleukopenia virus Ab.IgG
C1147077|T201|COMP|31392-4|LNC|Feline panleukopenia virus Ab.IgM|Feline panleukopenia virus Ab.IgM
C1147078|T201|COMP|31393-2|LNC|Feline herpesvirus 1 Ab|Feline herpesvirus 1 Ab
C1147079|T201|COMP|31394-0|LNC|Feline syncytial virus Ab|Feline syncytial virus Ab
C1147080|T201|COMP|31395-7|LNC|Filovirus Ab|Filovirus Ab
C1147081|T201|COMP|31396-5|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C1147082|T201|COMP|31397-3|LNC|Ganglioside GD1a Ab.IgG|Ganglioside GD1a Ab.IgG
C1147083|T201|COMP|31398-1|LNC|Ganglioside GD1a Ab.IgM|Ganglioside GD1a Ab.IgM
C1147084|T201|COMP|31399-9|LNC|Ganglioside GD1a Ab.IgM|Ganglioside GD1a Ab.IgM
C1147085|T201|COMP|31400-5|LNC|Ganglioside GD1b Ab|Ganglioside GD1b Ab
C1147086|T201|COMP|31401-3|LNC|Ganglioside GD1b Ab.IgG|Ganglioside GD1b Ab.IgG
C1147087|T201|COMP|31402-1|LNC|Ganglioside GD1b Ab.IgG|Ganglioside GD1b Ab.IgG
C1147088|T201|COMP|31403-9|LNC|Ganglioside GD1b Ab.IgM|Ganglioside GD1b Ab.IgM
C1147089|T201|COMP|31404-7|LNC|Ganglioside GM1b Ab.IgG|Ganglioside GM1b Ab.IgG
C1147090|T201|COMP|31405-4|LNC|Ganglioside GM1b Ab.IgM|Ganglioside GM1b Ab.IgM
C1147091|T201|COMP|31406-2|LNC|Glomerular basement membrane Ab.IgG|Glomerular basement membrane Ab.IgG
C1147092|T201|COMP|31407-0|LNC|Haemophilus somnus Ab|Haemophilus somnus Ab
C1147093|T201|COMP|31408-8|LNC|Hantavirus sin nombre Ab.IgG|Hantavirus sin nombre Ab.IgG
C1147094|T201|COMP|31409-6|LNC|Hantavirus sin nombre Ab.IgM|Hantavirus sin nombre Ab.IgM
C1147095|T201|COMP|31410-4|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C1147096|T201|COMP|31411-2|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C1147097|T201|COMP|31412-0|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C1147098|T201|COMP|31413-8|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C1147099|T201|COMP|31414-6|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C1147100|T201|COMP|31415-3|LNC|Herpes virus 6 Ab.IgM|Herpes virus 6 Ab.IgM
C1147101|T201|COMP|31416-1|LNC|Herpes virus 7 Ab.IgG|Herpes virus 7 Ab.IgG
C1147102|T201|COMP|31417-9|LNC|Herpes virus 7 Ab.IgM|Herpes virus 7 Ab.IgM
C1147103|T201|COMP|31418-7|LNC|Heterophile Ab|Heterophile Ab
C1147104|T201|COMP|31419-5|LNC|Heterophile Ab|Heterophile Ab
C1147105|T201|COMP|31420-3|LNC|Highlands J virus Ab|Highlands J virus Ab
C1147106|T201|COMP|31421-1|LNC|Highlands J virus Ab|Highlands J virus Ab
C1147107|T201|COMP|31422-9|LNC|Highlands J virus Ab|Highlands J virus Ab
C1147108|T201|COMP|31423-7|LNC|Histone Ab.IgG|Histone Ab.IgG
C1147109|T201|COMP|31424-5|LNC|Histone H2a+H2b Ab|Histone H2a+H2b Ab
C1147110|T201|COMP|31425-2|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C1147111|T201|COMP|31426-0|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C1147112|T201|COMP|31427-8|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C1147113|T201|COMP|31428-6|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C1147114|T201|COMP|31429-4|LNC|Histoplasma sp Ab|Histoplasma sp Ab
C1147115|T201|COMP|31430-2|LNC|HIV 1 Ab.IgG|HIV 1 Ab.IgG
C1147116|T201|COMP|31431-0|LNC|HTLV I+II Ab.IgG|HTLV I+II Ab.IgG
C1147117|T201|COMP|31432-8|LNC|Human antimouse Ab|Human antimouse Ab
C1147118|T201|COMP|31433-6|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1147119|T201|COMP|31434-4|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1147120|T201|COMP|31435-1|LNC|Hyaluronidase Ab|Hyaluronidase Ab
C1147121|T201|COMP|31436-9|LNC|Infectious bursal disease virus Ab|Infectious bursal disease virus Ab
C1147122|T201|COMP|31437-7|LNC|Influenza virus A Ab.IgG|Influenza virus A Ab.IgG
C1147123|T201|COMP|31438-5|LNC|Influenza virus A Ab.IgM|Influenza virus A Ab.IgM
C1147124|T201|COMP|31439-3|LNC|Insulin receptor Ab|Insulin receptor Ab
C1147125|T201|COMP|31440-1|LNC|Intercalated disk Ab|Intercalated disk Ab
C1147126|T201|COMP|31441-9|LNC|Intercellular substance Ab|Intercellular substance Ab
C1147127|T201|COMP|31442-7|LNC|Interferon.beta 1 Ab|Interferon.beta 1 Ab
C1147128|T201|COMP|31443-5|LNC|Intrinsic factor blocking Ab|Intrinsic factor blocking Ab
C1147129|T201|COMP|31444-3|LNC|Intrinsic factor blocking Ab|Intrinsic factor blocking Ab
C1147130|T201|COMP|31445-0|LNC|Intrinsic factor blocking Ab.IgG|Intrinsic factor blocking Ab.IgG
C1147131|T201|COMP|31446-8|LNC|Jamestown canyon virus Ab|Jamestown canyon virus Ab
C1147132|T201|COMP|31448-4|LNC|La Crosse virus Ab|La Crosse virus Ab
C1147133|T201|COMP|31449-2|LNC|La Crosse virus Ab|La Crosse virus Ab
C1147134|T201|COMP|31450-0|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C1147135|T201|COMP|31451-8|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C1147136|T201|COMP|31452-6|LNC|Lassa virus Ab.IgG|Lassa virus Ab.IgG
C1147137|T201|COMP|31453-4|LNC|Lassa virus Ab.IgM|Lassa virus Ab.IgM
C1147138|T201|COMP|31454-2|LNC|Legionella pneumophila 1 Ab|Legionella pneumophila 1 Ab
C1147139|T201|COMP|31455-9|LNC|Legionella pneumophila 1 Ab.IgG|Legionella pneumophila 1 Ab.IgG
C1147140|T201|COMP|31456-7|LNC|Legionella pneumophila 1 Ab.IgM|Legionella pneumophila 1 Ab.IgM
C1147141|T201|COMP|31457-5|LNC|Legionella pneumophila 2 Ab|Legionella pneumophila 2 Ab
C1147142|T201|COMP|31458-3|LNC|Legionella pneumophila 2 Ab.IgG|Legionella pneumophila 2 Ab.IgG
C1147143|T201|COMP|31459-1|LNC|Legionella pneumophila 3 Ab|Legionella pneumophila 3 Ab
C1147144|T201|COMP|31460-9|LNC|Legionella pneumophila 3 Ab.IgG|Legionella pneumophila 3 Ab.IgG
C1147145|T201|COMP|31461-7|LNC|Legionella pneumophila 4 Ab|Legionella pneumophila 4 Ab
C1147146|T201|COMP|31462-5|LNC|Legionella pneumophila 4 Ab.IgG|Legionella pneumophila 4 Ab.IgG
C1147147|T201|COMP|31463-3|LNC|Legionella pneumophila 5 Ab|Legionella pneumophila 5 Ab
C1147148|T201|COMP|31464-1|LNC|Legionella pneumophila 5 Ab.IgG|Legionella pneumophila 5 Ab.IgG
C1147149|T201|COMP|31465-8|LNC|Legionella pneumophila 6 Ab|Legionella pneumophila 6 Ab
C1147150|T201|COMP|31466-6|LNC|Legionella pneumophila 6 Ab.IgG|Legionella pneumophila 6 Ab.IgG
C1147151|T201|COMP|31467-4|LNC|Legionella pneumophila 6 Ab.IgM|Legionella pneumophila 6 Ab.IgM
C1147152|T201|COMP|31468-2|LNC|Legionella pneumophila 7 Ab|Legionella pneumophila 7 Ab
C1147153|T201|COMP|31469-0|LNC|Legionella pneumophila 8 Ab|Legionella pneumophila 8 Ab
C1147154|T201|COMP|31470-8|LNC|Legionella pneumophila 9 Ab|Legionella pneumophila 9 Ab
C1147155|T201|COMP|31471-6|LNC|Legionella pneumophila Ab|Legionella pneumophila Ab
C1147156|T201|COMP|31472-4|LNC|Legionella pneumophila Ab.IgM|Legionella pneumophila Ab.IgM
C1147157|T201|COMP|31473-2|LNC|Legionella pneumophila atypical Ab|Legionella pneumophila atypical Ab
C1147158|T201|COMP|31474-0|LNC|Legionella sp Ab.IgM|Legionella sp Ab.IgM
C1147159|T201|COMP|31475-7|LNC|Leishmania donovani Ab|Leishmania donovani Ab
C1147160|T201|COMP|31476-5|LNC|Leptospira borgpetersenii serovar Sejroe Ab|Leptospira borgpetersenii serovar Sejroe Ab
C1147161|T201|COMP|31477-3|LNC|Leptospira interrogans serovar Bratislava Ab|Leptospira interrogans serovar Bratislava Ab
C1147162|T201|COMP|31478-1|LNC|Leptospira interrogans serovar Canicola Ab|Leptospira interrogans serovar Canicola Ab
C1147163|T201|COMP|31479-9|LNC|Leptospira interrogans serovar Grippotyphosa Ab|Leptospira interrogans serovar Grippotyphosa Ab
C1147164|T201|COMP|31480-7|LNC|Leptospira interrogans serovar Hardjo Ab|Leptospira interrogans serovar Hardjo Ab
C1147166|T201|COMP|31482-3|LNC|Leptospira interrogans serovar Pomona Ab|Leptospira interrogans serovar Pomona Ab
C1147167|T201|COMP|31483-1|LNC|Leptospira sp Ab|Leptospira sp Ab
C1147168|T201|COMP|31484-9|LNC|Leptospira sp Ab.IgG|Leptospira sp Ab.IgG
C1147169|T201|COMP|31485-6|LNC|Leptospira sp Ab.IgG|Leptospira sp Ab.IgG
C1147170|T201|COMP|31486-4|LNC|Leptospira sp Ab.IgM|Leptospira sp Ab.IgM
C1147171|T201|COMP|31487-2|LNC|Leptospira sp Ab.IgM|Leptospira sp Ab.IgM
C1147172|T201|COMP|31488-0|LNC|Listeria sp Ab|Listeria sp Ab
C1147173|T201|COMP|31489-8|LNC|Lumpy skin disease virus Ab|Lumpy skin disease virus Ab
C1147174|T201|COMP|31490-6|LNC|Lupus erythematosus deoxynucleoproteins Ab.IgG|Lupus erythematosus deoxynucleoproteins Ab.IgG
C1147175|T201|COMP|31491-4|LNC|Lymphocytic choriomeningitis virus Ab|Lymphocytic choriomeningitis virus Ab
C1147176|T201|COMP|31492-2|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C1147177|T201|COMP|31493-0|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C1147178|T201|COMP|31494-8|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C1147179|T201|COMP|31495-5|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C1147180|T201|COMP|31496-3|LNC|Ganglioside GM1 Ab|Ganglioside GM1 Ab
C1147181|T201|COMP|31497-1|LNC|Ganglioside GM1 Ab|Ganglioside GM1 Ab
C1147182|T201|COMP|31498-9|LNC|Ganglioside GM1 Ab.IgA|Ganglioside GM1 Ab.IgA
C1147183|T201|COMP|31499-7|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C1147184|T201|COMP|31500-2|LNC|Ganglioside GM1 Ab.IgG+IgM|Ganglioside GM1 Ab.IgG+IgM
C1147185|T201|COMP|31501-0|LNC|Ganglioside GM1 Ab.IgG+IgM|Ganglioside GM1 Ab.IgG+IgM
C1147186|T201|COMP|31502-8|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C1147187|T201|COMP|31503-6|LNC|Mumps virus Ab|Mumps virus Ab
C1147188|T201|COMP|31504-4|LNC|Mumps virus soluble Ab|Mumps virus soluble Ab
C1147189|T201|COMP|31505-1|LNC|Mumps virus soluble Ab|Mumps virus soluble Ab
C1147190|T201|COMP|31506-9|LNC|Mumps virus particle-bound Ab|Mumps virus particle-bound Ab
C1147191|T201|COMP|31507-7|LNC|Mumps virus particle-bound Ab|Mumps virus particle-bound Ab
C1147195|T201|COMP|31511-9|LNC|Mycoplasma gallisepticum Ab|Mycoplasma gallisepticum Ab
C1147196|T201|COMP|31512-7|LNC|Mycoplasma hominis Ab|Mycoplasma hominis Ab
C1147197|T201|COMP|31513-5|LNC|Mycoplasma hyopneumoniae Ab|Mycoplasma hyopneumoniae Ab
C1147199|T201|COMP|31515-0|LNC|Mycoplasma pneumoniae Ab.IgA|Mycoplasma pneumoniae Ab.IgA
C1147200|T201|COMP|31516-8|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C1147201|T201|COMP|31517-6|LNC|Mycoplasma sp Ab|Mycoplasma sp Ab
C1147202|T201|COMP|31518-4|LNC|Mycoplasma synoviae Ab|Mycoplasma synoviae Ab
C1147203|T201|COMP|31519-2|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C1147204|T201|COMP|31520-0|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C1147205|T201|COMP|31521-8|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C1147206|T201|COMP|31522-6|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C1147207|T201|COMP|31523-4|LNC|Myxoma virus Ab|Myxoma virus Ab
C1147208|T201|COMP|31524-2|LNC|Nairobi sheep disease virus Ab|Nairobi sheep disease virus Ab
C1147209|T201|COMP|31525-9|LNC|Neisseria gonorrhoeae Ab|Neisseria gonorrhoeae Ab
C1147210|T201|COMP|31526-7|LNC|Neisseria meningitidis serogroup A Ab.IgG|Neisseria meningitidis serogroup A Ab.IgG
C1147211|T201|COMP|31527-5|LNC|Neisseria meningitidis serogroup C Ab.IgG|Neisseria meningitidis serogroup C Ab.IgG
C1147212|T201|COMP|31528-3|LNC|Neisseria meningitidis serogroup Y Ab|Neisseria meningitidis serogroup Y Ab
C1147213|T201|COMP|31529-1|LNC|Neospora caninum Ab|Neospora caninum Ab
C1147214|T201|COMP|31530-9|LNC|Neuronal Ab|Neuronal Ab
C1147215|T201|COMP|31531-7|LNC|Neuronal Ab|Neuronal Ab
C1147216|T201|COMP|31532-5|LNC|Neuronal Ab|Neuronal Ab
C1147217|T201|COMP|31533-3|LNC|Neuronal Ab|Neuronal Ab
C1147218|T201|COMP|31534-1|LNC|Neuronal Ab.IgG|Neuronal Ab.IgG
C1147219|T201|COMP|31535-8|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C1147220|T201|COMP|31536-6|LNC|Neuronal nuclear Ab.IgG|Neuronal nuclear Ab.IgG
C1147221|T201|COMP|31537-4|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C1147222|T201|COMP|31538-2|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C1147223|T201|COMP|31539-0|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C1147224|T201|COMP|31540-8|LNC|Nuclear Ab|Nuclear Ab
C1147225|T201|COMP|31541-6|LNC|Nuclear Ab|Nuclear Ab
C1147226|T201|COMP|31542-4|LNC|Nuclear Ab|Nuclear Ab
C1147227|T201|COMP|31543-2|LNC|Nuclear Ab|Nuclear Ab
C1147228|T201|COMP|31544-0|LNC|Nuclear Ab|Nuclear Ab
C1147229|T201|COMP|31545-7|LNC|Nuclear Ab.IgG|Nuclear Ab.IgG
C1147230|T201|COMP|31546-5|LNC|Ovary Ab.IgG|Ovary Ab.IgG
C1147231|T201|COMP|31547-3|LNC|Pancreatic islet cell Ab|Pancreatic islet cell Ab
C1147232|T201|COMP|31548-1|LNC|Parainfluenza virus 1 Ab|Parainfluenza virus 1 Ab
C1147233|T201|COMP|31549-9|LNC|Parainfluenza virus 1 Ab.IgM|Parainfluenza virus 1 Ab.IgM
C1147234|T201|COMP|31550-7|LNC|Parainfluenza virus 2 Ab|Parainfluenza virus 2 Ab
C1147235|T201|COMP|31551-5|LNC|Parainfluenza virus 2 Ab.IgM|Parainfluenza virus 2 Ab.IgM
C1147236|T201|COMP|31552-3|LNC|Parainfluenza virus 3 Ab|Parainfluenza virus 3 Ab
C1147237|T201|COMP|31553-1|LNC|Parainfluenza virus 3 Ab.IgG|Parainfluenza virus 3 Ab.IgG
C1147238|T201|COMP|31554-9|LNC|Parainfluenza virus 3 Ab.IgM|Parainfluenza virus 3 Ab.IgM
C1147239|T201|COMP|31555-6|LNC|Parainfluenza virus Ab|Parainfluenza virus Ab
C1147240|T201|COMP|31556-4|LNC|Parietal cell Ab.IgG|Parietal cell Ab.IgG
C1147241|T201|COMP|31557-2|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C1147242|T201|COMP|31558-0|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C1147243|T201|COMP|31559-8|LNC|Pasteurella multocida Ab|Pasteurella multocida Ab
C1147244|T201|COMP|31560-6|LNC|Peste des petits ruminants virus Ab|Peste des petits ruminants virus Ab
C1147245|T201|COMP|31561-4|LNC|Phospholipid Ab.IgA|Phospholipid Ab.IgA
C1147246|T201|COMP|31562-2|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C1147247|T201|COMP|31563-0|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C1147248|T201|COMP|31564-8|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C1147249|T201|COMP|31565-5|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C1147250|T201|COMP|31566-3|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C1147251|T201|COMP|31567-1|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C1147252|T201|COMP|31568-9|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C1147253|T201|COMP|31569-7|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C1147254|T201|COMP|31570-5|LNC|Porcine influenza virus A Ab|Porcine influenza virus A Ab
C1147255|T201|COMP|31571-3|LNC|Porcine parvovirus Ab|Porcine parvovirus Ab
C1147257|T201|COMP|31573-9|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1147258|T201|COMP|31574-7|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1147259|T201|COMP|31575-4|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1147260|T201|COMP|31576-2|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1147261|T201|COMP|31577-0|LNC|Pseudorabies virus Ab|Pseudorabies virus Ab
C1147262|T201|COMP|31578-8|LNC|Pullularia sp Ab|Pullularia sp Ab
C1147263|T201|COMP|31579-6|LNC|Purkinje cells Ab|Purkinje cells Ab
C1147264|T201|COMP|31580-4|LNC|Purkinje cells Ab.IgG|Purkinje cells Ab.IgG
C1147265|T201|COMP|31581-2|LNC|Reovirus Ab|Reovirus Ab
C1147266|T201|COMP|31582-0|LNC|Reovirus Ab|Reovirus Ab
C1147267|T201|COMP|31583-8|LNC|Respiratory syncytial virus Ab.IgG|Respiratory syncytial virus Ab.IgG
C1147268|T201|COMP|31584-6|LNC|Reticulin Ab.IgG|Reticulin Ab.IgG
C1147269|T201|COMP|31585-3|LNC|Reticulin Ab.IgG|Reticulin Ab.IgG
C1147270|T201|COMP|31586-1|LNC|Rhodococcus equi Ab|Rhodococcus equi Ab
C1147271|T201|COMP|31587-9|LNC|Rhodococcus equi Ab|Rhodococcus equi Ab
C1147272|T201|COMP|31588-7|LNC|Ribonucleoprotein extractable nuclear Ab.IgG|Ribonucleoprotein extractable nuclear Ab.IgG
C1147273|T201|COMP|31589-5|LNC|Ribosomal Ab|Ribosomal Ab
C1147274|T201|COMP|31590-3|LNC|Ribosomal Ab|Ribosomal Ab
C1147275|T201|COMP|31591-1|LNC|Ribosomal P Ab|Ribosomal P Ab
C1147276|T201|COMP|31592-9|LNC|Ribosomal P Ab|Ribosomal P Ab
C1147277|T201|COMP|31593-7|LNC|Rickettsia (Proteus OX19) Ab|Rickettsia (Proteus OX19) Ab
C1147278|T201|COMP|31594-5|LNC|Rickettsia (Proteus OXK) Ab|Rickettsia (Proteus OXK) Ab
C1147279|T201|COMP|31595-2|LNC|Rickettsia akari Ab|Rickettsia akari Ab
C1147280|T201|COMP|31596-0|LNC|Rickettsia australis Ab|Rickettsia australis Ab
C1147281|T201|COMP|31597-8|LNC|Rickettsia conorii Ab|Rickettsia conorii Ab
C1147282|T201|COMP|31598-6|LNC|Rickettsia honei Ab|Rickettsia honei Ab
C1147283|T201|COMP|31599-4|LNC|Rickettsia prowazekii Ab.IgG|Rickettsia prowazekii Ab.IgG
C1147284|T201|COMP|31600-0|LNC|Rickettsia prowazekii Ab.IgM|Rickettsia prowazekii Ab.IgM
C1147285|T201|COMP|31601-8|LNC|Rickettsia spotted fever group Ab.IgM|Rickettsia spotted fever group Ab.IgM
C1147286|T201|COMP|31602-6|LNC|Rickettsia typhus group Ab.IgM|Rickettsia typhus group Ab.IgM
C1147287|T201|COMP|31603-4|LNC|Rickettsia rickettsii Ab|Rickettsia rickettsii Ab
C1147288|T201|COMP|31604-2|LNC|Rickettsia rickettsii Ab|Rickettsia rickettsii Ab
C1147289|T201|COMP|31605-9|LNC|Rickettsia sibirica Ab|Rickettsia sibirica Ab
C1147290|T201|COMP|31606-7|LNC|Orientia tsutsugamushi Ab.IgG|Orientia tsutsugamushi Ab.IgG
C1147291|T201|COMP|31607-5|LNC|Orientia tsutsugamushi Gilliam Ab|Orientia tsutsugamushi Gilliam Ab
C1147292|T201|COMP|31608-3|LNC|Orientia tsutsugamushi Karp Ab|Orientia tsutsugamushi Karp Ab
C1147293|T201|COMP|31609-1|LNC|Orientia tsutsugamushi Kato Ab|Orientia tsutsugamushi Kato Ab
C1147294|T201|COMP|31610-9|LNC|Orientia tsutsugamushi Litchfield Ab|Orientia tsutsugamushi Litchfield Ab
C1147295|T201|COMP|31611-7|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C1147296|T201|COMP|31612-5|LNC|Rift valley fever virus Ab|Rift valley fever virus Ab
C1147297|T201|COMP|31613-3|LNC|Rinderpest virus Ab|Rinderpest virus Ab
C1147298|T201|COMP|31614-1|LNC|Ross river virus Ab.IgG|Ross river virus Ab.IgG
C1147299|T201|COMP|31615-8|LNC|Ross river virus Ab.IgM|Ross river virus Ab.IgM
C1147300|T201|COMP|31616-6|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C1147301|T201|COMP|31617-4|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C1147302|T201|COMP|31618-2|LNC|Salmonella paratyphi B H Ab|Salmonella paratyphi B H Ab
C1147303|T201|COMP|31619-0|LNC|Salmonella paratyphi B O Ab|Salmonella paratyphi B O Ab
C1147304|T201|COMP|31620-8|LNC|Salmonella pullorum Ab|Salmonella pullorum Ab
C1147305|T201|COMP|31621-6|LNC|Salmonella typhi H D Ab|Salmonella typhi H D Ab
C1147306|T201|COMP|31622-4|LNC|Salmonella typhi O D Ab|Salmonella typhi O D Ab
C1147307|T201|COMP|31623-2|LNC|Salmonella typhimurium Ab|Salmonella typhimurium Ab
C1147308|T201|COMP|31624-0|LNC|Schistosoma sp Ab.IgG|Schistosoma sp Ab.IgG
C1147309|T201|COMP|31625-7|LNC|Sjogrens syndrome-A extractable nuclear Ab.IgG|Sjogrens syndrome-A extractable nuclear Ab.IgG
C1147310|T201|COMP|31626-5|LNC|Sjogrens syndrome-B extractable nuclear Ab.IgG|Sjogrens syndrome-B extractable nuclear Ab.IgG
C1147311|T201|COMP|31627-3|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C1147313|T201|COMP|31629-9|LNC|Smooth muscle Ab|Smooth muscle Ab
C1147314|T201|COMP|31630-7|LNC|Spermatozoa Ab|Spermatozoa Ab
C1147315|T201|COMP|31631-5|LNC|Spermatozoa Ab|Spermatozoa Ab
C1147316|T201|COMP|31632-3|LNC|Spermatozoa Ab|Spermatozoa Ab
C1147317|T201|COMP|31633-1|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C1147318|T201|COMP|31634-9|LNC|Stachybotrys chartarum Ab.IgA|Stachybotrys chartarum Ab.IgA
C1147319|T201|COMP|31635-6|LNC|Streptococcus pneumoniae 1 Ab.IgG^1st specimen|Streptococcus pneumoniae 1 Ab.IgG^1st specimen
C1147320|T201|COMP|31636-4|LNC|Streptococcus pneumoniae 14 Ab|Streptococcus pneumoniae 14 Ab
C1147321|T201|COMP|31637-2|LNC|Streptococcus pneumoniae 23 Ab.IgG^1st specimen|Streptococcus pneumoniae 23 Ab.IgG^1st specimen
C1147322|T201|COMP|31638-0|LNC|Streptococcus pneumoniae 23 Ab.IgG^2nd specimen|Streptococcus pneumoniae 23 Ab.IgG^2nd specimen
C1147324|T201|COMP|31640-6|LNC|Streptococcus pneumoniae 3 Ab|Streptococcus pneumoniae 3 Ab
C1147325|T201|COMP|31641-4|LNC|Streptococcus pneumoniae 3 Ab.IgG^1st specimen|Streptococcus pneumoniae 3 Ab.IgG^1st specimen
C1147326|T201|COMP|31642-2|LNC|Streptococcus pneumoniae 3 Ab.IgG^2nd specimen|Streptococcus pneumoniae 3 Ab.IgG^2nd specimen
C1147327|T201|COMP|31643-0|LNC|Streptococcus pneumoniae 4 Ab.IgG^1st specimen|Streptococcus pneumoniae 4 Ab.IgG^1st specimen
C1147328|T201|COMP|31644-8|LNC|Streptococcus pneumoniae 4 Ab.IgG^2nd specimen|Streptococcus pneumoniae 4 Ab.IgG^2nd specimen
C1147332|T201|COMP|31648-9|LNC|Streptococcus pneumoniae 6 Ab.IgG|Streptococcus pneumoniae 6 Ab.IgG
C1147333|T201|COMP|31649-7|LNC|Streptococcus pneumoniae 6 Ab^2nd specimen|Streptococcus pneumoniae 6 Ab^2nd specimen
C1147335|T201|COMP|31651-3|LNC|Streptococcus pneumoniae 6a+6b Ab|Streptococcus pneumoniae 6a+6b Ab
C1147336|T201|COMP|31652-1|LNC|Streptococcus pneumoniae 6+26 Ab^1st specimen|Streptococcus pneumoniae 6+26 Ab^1st specimen
C1147337|T201|COMP|31653-9|LNC|Streptococcus pneumoniae 8 Ab.IgG^1st specimen|Streptococcus pneumoniae 8 Ab.IgG^1st specimen
C1147338|T201|COMP|31654-7|LNC|Streptococcus pneumoniae 8 Ab.IgG^2nd specimen|Streptococcus pneumoniae 8 Ab.IgG^2nd specimen
C1147339|T201|COMP|31655-4|LNC|Streptococcus pneumoniae 9 Ab|Streptococcus pneumoniae 9 Ab
C1147340|T201|COMP|31656-2|LNC|Streptococcus pneumoniae 9 Ab.IgG^1st specimen|Streptococcus pneumoniae 9 Ab.IgG^1st specimen
C1147341|T201|COMP|31657-0|LNC|Streptococcus pneumoniae 9 Ab.IgG^2nd specimen|Streptococcus pneumoniae 9 Ab.IgG^2nd specimen
C1147342|T201|COMP|31658-8|LNC|Streptococcus pyogenes enzyme Ab|Streptococcus pyogenes enzyme Ab
C1147343|T201|COMP|31659-6|LNC|Striated muscle Ab|Striated muscle Ab
C1147344|T201|COMP|31660-4|LNC|Striated muscle Ab.IgG|Striated muscle Ab.IgG
C1147345|T201|COMP|31661-2|LNC|Sulfate-3-Glucuronyl paragloboside Ab|Sulfate-3-Glucuronyl paragloboside Ab
C1147346|T201|COMP|31662-0|LNC|Sulfate-3-Glucuronyl paragloboside Ab|Sulfate-3-Glucuronyl paragloboside Ab
C1147347|T201|COMP|31663-8|LNC|Sulfate-3-Glucuronyl paragloboside Ab.IgM|Sulfate-3-Glucuronyl paragloboside Ab.IgM
C1147348|T201|COMP|31664-6|LNC|Sulfate-3-Glucuronyl paragloboside Ab.IgM|Sulfate-3-Glucuronyl paragloboside Ab.IgM
C1147349|T201|COMP|31665-3|LNC|Sulfate-3-Glucuronyl paragloboside Ab.IgM|Sulfate-3-Glucuronyl paragloboside Ab.IgM
C1147350|T201|COMP|31666-1|LNC|Sulfate-3-Glucuronyl paragloboside Ab.IgM|Sulfate-3-Glucuronyl paragloboside Ab.IgM
C1147351|T201|COMP|31667-9|LNC|Sulfatide Ab|Sulfatide Ab
C1147352|T201|COMP|31668-7|LNC|Sulfatide Ab|Sulfatide Ab
C1147353|T201|COMP|31669-5|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C1147354|T201|COMP|31670-3|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C1147355|T201|COMP|31671-1|LNC|Sulfatide Ab.IgM|Sulfatide Ab.IgM
C1147356|T201|COMP|31672-9|LNC|Taylorella equigenitalis Ab|Taylorella equigenitalis Ab
C1147357|T201|COMP|31673-7|LNC|Teichoate Ab|Teichoate Ab
C1147358|T201|COMP|31674-5|LNC|Ganglioside GQ1b Ab|Ganglioside GQ1b Ab
C1147358|T201|COMP|48397-4|LNC|Ganglioside GQ1b Ab|Ganglioside GQ1b Ab
C1147359|T201|COMP|31675-2|LNC|Tetrasialylganglioside GQ1b Ab|Tetrasialylganglioside GQ1b Ab
C1147360|T201|COMP|31676-0|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C1147361|T201|COMP|31677-8|LNC|Tetrasialylganglioside GQ1b Ab.IgG|Tetrasialylganglioside GQ1b Ab.IgG
C1147362|T201|COMP|31678-6|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C1147363|T201|COMP|31679-4|LNC|Tetrasialylganglioside GQ1b Ab.IgG|Tetrasialylganglioside GQ1b Ab.IgG
C1147364|T201|COMP|31680-2|LNC|Theileria annulata Ab|Theileria annulata Ab
C1147365|T201|COMP|31681-0|LNC|Theileria mutans Ab|Theileria mutans Ab
C1147366|T201|COMP|31682-8|LNC|Theileria parva Ab|Theileria parva Ab
C1147367|T201|COMP|31683-6|LNC|Thermoactinomyces sp Ab.IgG|Thermoactinomyces sp Ab.IgG
C1147368|T201|COMP|31684-4|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C1147369|T201|COMP|31685-1|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C1147370|T201|COMP|31686-9|LNC|Transmissible gastroenteritis virus Ab|Transmissible gastroenteritis virus Ab
C1147371|T201|COMP|31687-7|LNC|Trichinella sp Ab.IgM|Trichinella sp Ab.IgM
C1147372|T201|COMP|31688-5|LNC|Trivittatus virus Ab|Trivittatus virus Ab
C1147373|T201|COMP|31689-3|LNC|Trivittatus virus Ab|Trivittatus virus Ab
C1147374|T201|COMP|31690-1|LNC|Trivittatus virus Ab|Trivittatus virus Ab
C1147375|T201|COMP|31691-9|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C1147376|T201|COMP|31692-7|LNC|Trypanosoma equiperdum Ab|Trypanosoma equiperdum Ab
C1147377|T201|COMP|31693-5|LNC|Unidentified extractable nuclear Ab|Unidentified extractable nuclear Ab
C1147378|T201|COMP|31694-3|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C1147379|T201|COMP|31695-0|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C1147380|T201|COMP|31696-8|LNC|Vesicular stomatitis Indiana virus Ab|Vesicular stomatitis Indiana virus Ab
C1147381|T201|COMP|31697-6|LNC|Vesicular stomatitis New Jersey virus Ab|Vesicular stomatitis New Jersey virus Ab
C1147382|T201|COMP|31698-4|LNC|Vibrio cholerae Ab|Vibrio cholerae Ab
C1147383|T201|COMP|31699-2|LNC|Viral hemorrhagic disease virus Ab|Viral hemorrhagic disease virus Ab
C1147384|T201|COMP|31700-8|LNC|West Nile virus Ab|West Nile virus Ab
C1147385|T201|COMP|31701-6|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C1147386|T201|COMP|31702-4|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C1147387|T201|COMP|31703-2|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1147388|T201|COMP|31704-0|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1147389|T201|COMP|31705-7|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C1147390|T201|COMP|31706-5|LNC|Western equine encephalitis virus Ab.IgG|Western equine encephalitis virus Ab.IgG
C1147391|T201|COMP|31707-3|LNC|Yersinia enterocolitica O:5 Ab|Yersinia enterocolitica O:5 Ab
C1147392|T201|COMP|31708-1|LNC|Yersinia enterocolitica Ab|Yersinia enterocolitica Ab
C1147393|T201|COMP|31709-9|LNC|Adenovirus 40+41 Ag|Adenovirus 40+41 Ag
C1147394|T201|COMP|31710-7|LNC|Adenovirus Ag|Adenovirus Ag
C1147395|T201|COMP|31711-5|LNC|Adenovirus Ag|Adenovirus Ag
C1147396|T201|COMP|31712-3|LNC|Adenovirus Ag|Adenovirus Ag
C1147397|T201|COMP|31713-1|LNC|Adenovirus Ag|Adenovirus Ag
C1147398|T201|COMP|31714-9|LNC|Adenovirus Ag|Adenovirus Ag
C1147399|T201|COMP|31715-6|LNC|African horse sickness virus Ag|African horse sickness virus Ag
C1147400|T201|COMP|31716-4|LNC|African swine fever virus Ag|African swine fever virus Ag
C1147401|T201|COMP|31717-2|LNC|Alcelaphine herpesvirus 1 Ag|Alcelaphine herpesvirus 1 Ag
C1147402|T201|COMP|31718-0|LNC|Astrovirus Ag|Astrovirus Ag
C1147403|T201|COMP|31719-8|LNC|Infectious bronchitis virus Ag|Infectious bronchitis virus Ag
C1147404|T201|COMP|31720-6|LNC|Avian infectious laryngotracheitis virus Ag|Avian infectious laryngotracheitis virus Ag
C1147405|T201|COMP|31721-4|LNC|Avian infectious laryngotracheitis virus Ag|Avian infectious laryngotracheitis virus Ag
C1147406|T201|COMP|31722-2|LNC|Avian infectious laryngotracheitis virus Ag|Avian infectious laryngotracheitis virus Ag
C1147407|T201|COMP|31723-0|LNC|Avian leukosis virus Ag|Avian leukosis virus Ag
C1147408|T201|COMP|31724-8|LNC|Avian leukosis virus Ag|Avian leukosis virus Ag
C1147409|T201|COMP|31725-5|LNC|Avian paramyxovirus 1 Ag|Avian paramyxovirus 1 Ag
C1147410|T201|COMP|31726-3|LNC|Bacillus anthracis Ag|Bacillus anthracis Ag
C1147411|T201|COMP|31727-1|LNC|Bacteroides fragilis Ag|Bacteroides fragilis Ag
C1147412|T201|COMP|31728-9|LNC|Bacteroides melaninogenicus Ag|Bacteroides melaninogenicus Ag
C1147413|T201|COMP|31729-7|LNC|Bladder tumor Ag|Bladder tumor Ag
C1147414|T201|COMP|31730-5|LNC|Bladder tumor Ag|Bladder tumor Ag
C1147415|T201|COMP|31731-3|LNC|Blastomyces dermatitidis Ag|Blastomyces dermatitidis Ag
C1147416|T201|COMP|31732-1|LNC|Bluetongue virus Ag|Bluetongue virus Ag
C1147417|T201|COMP|31733-9|LNC|Border disease virus Ag|Border disease virus Ag
C1147418|T201|COMP|31734-7|LNC|Border disease virus Ag|Border disease virus Ag
C1147419|T201|COMP|31735-4|LNC|Bordetella bronchiseptica Ag|Bordetella bronchiseptica Ag
C1147420|T201|COMP|31736-2|LNC|Bordetella parapertussis Ag|Bordetella parapertussis Ag
C1147421|T201|COMP|31737-0|LNC|Bordetella pertussis Ag|Bordetella pertussis Ag
C1147422|T201|COMP|31738-8|LNC|Borrelia burgdorferi Ag|Borrelia burgdorferi Ag
C1147423|T201|COMP|31739-6|LNC|Borrelia sp Ag|Borrelia sp Ag
C1147424|T201|COMP|31740-4|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C1147425|T201|COMP|31741-2|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C1147426|T201|COMP|31742-0|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C1147427|T201|COMP|31743-8|LNC|Bovine diarrhea virus Ag|Bovine diarrhea virus Ag
C1147428|T201|COMP|31744-6|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C1147429|T201|COMP|31745-3|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C1147430|T201|COMP|31746-1|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C1147431|T201|COMP|31747-9|LNC|Bovine herpesvirus 1 Ag|Bovine herpesvirus 1 Ag
C1147432|T201|COMP|31748-7|LNC|Bovine herpesvirus 2 Ag|Bovine herpesvirus 2 Ag
C1147433|T201|COMP|31749-5|LNC|Bovine herpesvirus 4 Ag|Bovine herpesvirus 4 Ag
C1147434|T201|COMP|31750-3|LNC|Bovine inner ear Ag|Bovine inner ear Ag
C1147435|T201|COMP|31751-1|LNC|Bovine respiratory syncytial virus Ag|Bovine respiratory syncytial virus Ag
C1147436|T201|COMP|31752-9|LNC|Bovine virus diarrhea virus Ag|Bovine virus diarrhea virus Ag
C1147437|T201|COMP|31753-7|LNC|Brucella sp Ag|Brucella sp Ag
C1147438|T201|COMP|31754-5|LNC|Brucella sp Ag|Brucella sp Ag
C1147439|T201|COMP|31755-2|LNC|Campylobacter fetus Ag|Campylobacter fetus Ag
C1147440|T201|COMP|31756-0|LNC|Campylobacter fetus Ag|Campylobacter fetus Ag
C1147441|T201|COMP|31757-8|LNC|Canarypox virus Ag|Canarypox virus Ag
C1147442|T201|COMP|31758-6|LNC|Candida albicans Ag|Candida albicans Ag
C1147443|T201|COMP|31759-4|LNC|Candida albicans Ag|Candida albicans Ag
C1147444|T201|COMP|31760-2|LNC|Candida sp Ag|Candida sp Ag
C1147445|T201|COMP|31761-0|LNC|Canine parvovirus Ag|Canine parvovirus Ag
C1147446|T201|COMP|31762-8|LNC|Capripox virus Ag|Capripox virus Ag
C1147447|T201|COMP|31763-6|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1147448|T201|COMP|31764-4|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1147449|T201|COMP|31765-1|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1147450|T201|COMP|31766-9|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1147451|T201|COMP|31767-7|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1147452|T201|COMP|31768-5|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147453|T201|COMP|31769-3|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147454|T201|COMP|31770-1|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147455|T201|COMP|31771-9|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147456|T201|COMP|31772-7|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147457|T201|COMP|31773-5|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147458|T201|COMP|31774-3|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147459|T201|COMP|31775-0|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147460|T201|COMP|31776-8|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147461|T201|COMP|31777-6|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1147462|T201|COMP|31778-4|LNC|Chlamydophila pneumoniae Ag|Chlamydophila pneumoniae Ag
C1147463|T201|COMP|31779-2|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C1147464|T201|COMP|31780-0|LNC|Chlamydophila psittaci Ag|Chlamydophila psittaci Ag
C1147465|T201|COMP|31781-8|LNC|Classical swine fever virus Ag|Classical swine fever virus Ag
C1147466|T201|COMP|31782-6|LNC|Coccidioides immitis Ag|Coccidioides immitis Ag
C1147467|T201|COMP|31783-4|LNC|Coxiella burnetii Ag|Coxiella burnetii Ag
C1147468|T201|COMP|31784-2|LNC|Coxiella burnetii Ag|Coxiella burnetii Ag
C1147469|T201|COMP|31785-9|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C1147470|T201|COMP|31786-7|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C1147471|T201|COMP|31787-5|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C1147472|T201|COMP|31788-3|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1147473|T201|COMP|31789-1|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1147474|T201|COMP|31790-9|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1147475|T201|COMP|31791-7|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1147476|T201|COMP|31792-5|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1147477|T201|COMP|31793-3|LNC|Cryptosporidium sp Ag|Cryptosporidium sp Ag
C1147478|T201|COMP|31794-1|LNC|Cryptosporidium sp Ag|Cryptosporidium sp Ag
C1147479|T201|COMP|31795-8|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C1147480|T201|COMP|31796-6|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C1147481|T201|COMP|31797-4|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C1147482|T201|COMP|31798-2|LNC|Dengue virus Ag|Dengue virus Ag
C1147483|T201|COMP|31799-0|LNC|Dengue virus Ag|Dengue virus Ag
C1147484|T201|COMP|31800-6|LNC|Dermatophilus congolensis Ag|Dermatophilus congolensis Ag
C1147485|T201|COMP|31801-4|LNC|Dirofilaria immitis Ag|Dirofilaria immitis Ag
C1147486|T201|COMP|31802-2|LNC|Duck enteritis virus Ag|Duck enteritis virus Ag
C1147487|T201|COMP|31803-0|LNC|Duck hepatitis virus 1 Ag|Duck hepatitis virus 1 Ag
C1147488|T201|COMP|31804-8|LNC|Duck hepatitis virus 2 Ag|Duck hepatitis virus 2 Ag
C1147489|T201|COMP|31805-5|LNC|Duck hepatitis virus 3 Ag|Duck hepatitis virus 3 Ag
C1147490|T201|COMP|31806-3|LNC|Eastern equine encephalitis virus Ag|Eastern equine encephalitis virus Ag
C1147491|T201|COMP|31807-1|LNC|Eastern equine encephalitis virus Ag|Eastern equine encephalitis virus Ag
C1147492|T201|COMP|31808-9|LNC|Eastern equine encephalitis virus Ag|Eastern equine encephalitis virus Ag
C1147493|T201|COMP|31809-7|LNC|Echinococcus sp Ag|Echinococcus sp Ag
C1147494|T201|COMP|31810-5|LNC|Entamoeba histolytica Ag|Entamoeba histolytica Ag
C1147495|T201|COMP|31811-3|LNC|Entamoeba histolytica Ag|Entamoeba histolytica Ag
C1147496|T201|COMP|31812-1|LNC|Entamoeba histolytica Ag|Entamoeba histolytica Ag
C1147497|T201|COMP|31813-9|LNC|Epizootic hemorrhagic disease virus Ag|Epizootic hemorrhagic disease virus Ag
C1147498|T201|COMP|31814-7|LNC|Equine adenovirus Ag|Equine adenovirus Ag
C1147499|T201|COMP|31815-4|LNC|Equine arteritis virus Ag|Equine arteritis virus Ag
C1147500|T201|COMP|31816-2|LNC|Equine herpesvirus 1 Ag|Equine herpesvirus 1 Ag
C1147501|T201|COMP|31817-0|LNC|Equine herpesvirus 1 Ag|Equine herpesvirus 1 Ag
C1147502|T201|COMP|31818-8|LNC|Equine herpesvirus 1+4 Ag|Equine herpesvirus 1+4 Ag
C1147503|T201|COMP|31819-6|LNC|Equine herpesvirus 4 Ag|Equine herpesvirus 4 Ag
C1147504|T201|COMP|31820-4|LNC|Equine infectious anemia virus Ag|Equine infectious anemia virus Ag
C1147505|T201|COMP|31821-2|LNC|Equine influenza virus A1 Ag|Equine influenza virus A1 Ag
C1147506|T201|COMP|31822-0|LNC|Equine influenza virus A2 Ag|Equine influenza virus A2 Ag
C1147507|T201|COMP|31823-8|LNC|Equine influenza virus Ag|Equine influenza virus Ag
C1147508|T201|COMP|31824-6|LNC|Escherichia coli K1 Ag|Escherichia coli K1 Ag
C1147509|T201|COMP|31825-3|LNC|Escherichia coli K1 Ag|Escherichia coli K1 Ag
C1147510|T201|COMP|31826-1|LNC|Feline infectious peritonitis virus Ag|Feline infectious peritonitis virus Ag
C1147511|T201|COMP|31827-9|LNC|Foot and mouth disease virus Ag|Foot and mouth disease virus Ag
C1147512|T201|COMP|31828-7|LNC|Francisella tularensis Ag|Francisella tularensis Ag
C1147513|T201|COMP|31829-5|LNC|Francisella tularensis Ag|Francisella tularensis Ag
C1147514|T201|COMP|31830-3|LNC|Giardia lamblia Ag|Giardia lamblia Ag
C1147515|T201|COMP|31831-1|LNC|Giardia lamblia Ag^2nd specimen|Giardia lamblia Ag^2nd specimen
C1147516|T201|COMP|31832-9|LNC|Giardia lamblia Ag^3rd specimen|Giardia lamblia Ag^3rd specimen
C1147517|T201|COMP|31833-7|LNC|Haemophilus influenzae A Ag|Haemophilus influenzae A Ag
C1147518|T201|COMP|31834-5|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C1147519|T201|COMP|31835-2|LNC|Haemophilus influenzae C Ag|Haemophilus influenzae C Ag
C1147520|T201|COMP|31836-0|LNC|Haemophilus influenzae C Ag|Haemophilus influenzae C Ag
C1147521|T201|COMP|31837-8|LNC|Haemophilus influenzae D Ag|Haemophilus influenzae D Ag
C1147522|T201|COMP|31838-6|LNC|Haemophilus influenzae D Ag|Haemophilus influenzae D Ag
C1147523|T201|COMP|31839-4|LNC|Haemophilus influenzae E Ag|Haemophilus influenzae E Ag
C1147524|T201|COMP|31840-2|LNC|Haemophilus influenzae E Ag|Haemophilus influenzae E Ag
C1147525|T201|COMP|31841-0|LNC|Haemophilus influenzae F Ag|Haemophilus influenzae F Ag
C1147526|T201|COMP|31842-8|LNC|Haemophilus influenzae F Ag|Haemophilus influenzae F Ag
C1147527|T201|COMP|31843-6|LNC|Helicobacter pylori Ag|Helicobacter pylori Ag
C1147528|T201|COMP|31844-4|LNC|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C1147529|T201|COMP|31845-1|LNC|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C1147530|T201|COMP|31846-9|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1147531|T201|COMP|31847-7|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1147532|T201|COMP|31848-5|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1147533|T201|COMP|31849-3|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1147534|T201|COMP|31850-1|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1147535|T201|COMP|31851-9|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1147536|T201|COMP|31852-7|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1147537|T201|COMP|31853-5|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1147538|T201|COMP|31854-3|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1147539|T201|COMP|31855-0|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1147540|T201|COMP|31856-8|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1147541|T201|COMP|31857-6|LNC|Infectious bursal disease virus Ag|Infectious bursal disease virus Ag
C1147542|T201|COMP|31858-4|LNC|Influenza virus A Ag|Influenza virus A Ag
C1147543|T201|COMP|31859-2|LNC|Influenza virus A Ag|Influenza virus A Ag
C1147544|T201|COMP|31860-0|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C1147545|T201|COMP|31861-8|LNC|Influenza virus A+B+C Ag|Influenza virus A+B+C Ag
C1147546|T201|COMP|31862-6|LNC|Influenza virus A+B+C Ag|Influenza virus A+B+C Ag
C1147547|T201|COMP|31863-4|LNC|Influenza virus B Ag|Influenza virus B Ag
C1147548|T201|COMP|31864-2|LNC|Influenza virus B Ag|Influenza virus B Ag
C1147549|T201|COMP|31865-9|LNC|Influenza virus C Ag|Influenza virus C Ag
C1147550|T201|COMP|31866-7|LNC|Japanese encephalitis virus Ag|Japanese encephalitis virus Ag
C1147551|T201|COMP|31867-5|LNC|Lassa virus Ag|Lassa virus Ag
C1147552|T201|COMP|31868-3|LNC|Legionella pneumophila 1 Ag|Legionella pneumophila 1 Ag
C1147553|T201|COMP|31869-1|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C1147554|T201|COMP|31870-9|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C1147555|T201|COMP|31871-7|LNC|Leptospira interrogans Ag|Leptospira interrogans Ag
C1147556|T201|COMP|31872-5|LNC|Leptospira sp Ag|Leptospira sp Ag
C1147557|T201|COMP|31873-3|LNC|Mareks disease virus Ag|Mareks disease virus Ag
C1147558|T201|COMP|31874-1|LNC|Mareks disease virus Ag|Mareks disease virus Ag
C1147559|T201|COMP|31875-8|LNC|Measles virus Ag|Measles virus Ag
C1147560|T201|COMP|31876-6|LNC|Measles virus Ag|Measles virus Ag
C1147561|T201|COMP|31877-4|LNC|Measles virus Ag|Measles virus Ag
C1147562|T201|COMP|31878-2|LNC|Measles virus Ag|Measles virus Ag
C1147563|T201|COMP|31879-0|LNC|Measles virus Ag|Measles virus Ag
C1147564|T201|COMP|31880-8|LNC|Measles virus Ag|Measles virus Ag
C1147565|T201|COMP|31881-6|LNC|Measles virus Ag|Measles virus Ag
C1147566|T201|COMP|31882-4|LNC|Measles virus Ag|Measles virus Ag
C1147567|T201|COMP|31883-2|LNC|Measles virus Ag|Measles virus Ag
C1147568|T201|COMP|31884-0|LNC|Measles virus Ag|Measles virus Ag
C1147569|T201|COMP|31885-7|LNC|Measles virus Ag|Measles virus Ag
C1147570|T201|COMP|31886-5|LNC|Measles virus Ag|Measles virus Ag
C1147571|T201|COMP|31887-3|LNC|Measles virus Ag|Measles virus Ag
C1147572|T201|COMP|31888-1|LNC|Mumps virus Ag|Mumps virus Ag
C1147573|T201|COMP|31889-9|LNC|Mumps virus Ag|Mumps virus Ag
C1147574|T201|COMP|31890-7|LNC|Mumps virus Ag|Mumps virus Ag
C1147575|T201|COMP|31891-5|LNC|Mumps virus Ag|Mumps virus Ag
C1147576|T201|COMP|31892-3|LNC|Mumps virus Ag|Mumps virus Ag
C1147577|T201|COMP|31893-1|LNC|Mumps virus Ag|Mumps virus Ag
C1147578|T201|COMP|31894-9|LNC|Mumps virus Ag|Mumps virus Ag
C1147579|T201|COMP|31895-6|LNC|Mumps virus Ag|Mumps virus Ag
C1147580|T201|COMP|31896-4|LNC|Mumps virus Ag|Mumps virus Ag
C1147581|T201|COMP|31897-2|LNC|Mumps virus Ag|Mumps virus Ag
C1147582|T201|COMP|31898-0|LNC|Mumps virus Ag|Mumps virus Ag
C1147583|T201|COMP|31899-8|LNC|Mumps virus Ag|Mumps virus Ag
C1147584|T201|COMP|31900-4|LNC|Mumps virus Ag|Mumps virus Ag
C1147585|T201|COMP|31901-2|LNC|Mycoplasma gallisepticum Ag|Mycoplasma gallisepticum Ag
C1147587|T201|COMP|31903-8|LNC|Myxoma virus Ag|Myxoma virus Ag
C1147588|T201|COMP|31904-6|LNC|Nairobi sheep disease virus Ag|Nairobi sheep disease virus Ag
C1147589|T201|COMP|31905-3|LNC|Neisseria gonorrhoeae Ag|Neisseria gonorrhoeae Ag
C1147590|T201|COMP|31906-1|LNC|Neisseria gonorrhoeae Ag|Neisseria gonorrhoeae Ag
C1147591|T201|COMP|31907-9|LNC|Neisseria meningitidis serogroup A Ag|Neisseria meningitidis serogroup A Ag
C1147592|T201|COMP|31908-7|LNC|Neisseria meningitidis serogroup A Ag|Neisseria meningitidis serogroup A Ag
C1147593|T201|COMP|31909-5|LNC|Neisseria meningitidis serogroups A+C+w135+Y Ag|Neisseria meningitidis serogroups A+C+w135+Y Ag
C1147594|T201|COMP|31910-3|LNC|Neisseria meningitidis serogroups A+C+w135+Y Ag|Neisseria meningitidis serogroups A+C+w135+Y Ag
C1147595|T201|COMP|31911-1|LNC|Neisseria meningitidis Ag|Neisseria meningitidis Ag
C1147596|T201|COMP|31912-9|LNC|Neisseria meningitidis Ag|Neisseria meningitidis Ag
C1147597|T201|COMP|31913-7|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C1147600|T201|COMP|31916-0|LNC|Neisseria meningitidis serogroup C Ag|Neisseria meningitidis serogroup C Ag
C1147601|T201|COMP|31917-8|LNC|Neisseria meningitidis serogroup C Ag|Neisseria meningitidis serogroup C Ag
C1147602|T201|COMP|31918-6|LNC|Neisseria meningitidis serogroup w135 Ag|Neisseria meningitidis serogroup w135 Ag
C1147603|T201|COMP|31919-4|LNC|Neisseria meningitidis serogroup w135 Ag|Neisseria meningitidis serogroup w135 Ag
C1147604|T201|COMP|31920-2|LNC|Neisseria meningitidis serogroup w135 Ag|Neisseria meningitidis serogroup w135 Ag
C1147605|T201|COMP|31921-0|LNC|Neisseria meningitidis serogroup Y Ag|Neisseria meningitidis serogroup Y Ag
C1147606|T201|COMP|31922-8|LNC|Ovine progressive pneumonia virus Ag|Ovine progressive pneumonia virus Ag
C1147607|T201|COMP|31923-6|LNC|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C1147608|T201|COMP|31924-4|LNC|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C1147609|T201|COMP|31925-1|LNC|Parainfluenza virus 2 Ag|Parainfluenza virus 2 Ag
C1147610|T201|COMP|31926-9|LNC|Parainfluenza virus 2 Ag|Parainfluenza virus 2 Ag
C1147611|T201|COMP|31927-7|LNC|Parainfluenza virus 3 Ag|Parainfluenza virus 3 Ag
C1147612|T201|COMP|31928-5|LNC|Parainfluenza virus 3 Ag|Parainfluenza virus 3 Ag
C1147613|T201|COMP|31929-3|LNC|Parainfluenza virus Ag|Parainfluenza virus Ag
C1147614|T201|COMP|31930-1|LNC|Pasteurella multocida Ag|Pasteurella multocida Ag
C1147615|T201|COMP|31931-9|LNC|Plasmodium vivax Ag|Plasmodium vivax Ag
C1147616|T201|COMP|31932-7|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147617|T201|COMP|31933-5|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147618|T201|COMP|31934-3|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147619|T201|COMP|31935-0|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147620|T201|COMP|31936-8|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147621|T201|COMP|31937-6|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147622|T201|COMP|31938-4|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147623|T201|COMP|31939-2|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147624|T201|COMP|31940-0|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147625|T201|COMP|31941-8|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147626|T201|COMP|31942-6|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147627|T201|COMP|31943-4|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C1147628|T201|COMP|31944-2|LNC|Porcine enterovirus Ag|Porcine enterovirus Ag
C1147629|T201|COMP|31945-9|LNC|Pseudorabies virus Ag|Pseudorabies virus Ag
C1147630|T201|COMP|31946-7|LNC|Rabies virus Ag|Rabies virus Ag
C1147631|T201|COMP|31947-5|LNC|Rabies virus Ag|Rabies virus Ag
C1147632|T201|COMP|31948-3|LNC|Rabies virus Ag|Rabies virus Ag
C1147633|T201|COMP|31949-1|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C1147634|T201|COMP|31950-9|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C1147635|T201|COMP|31951-7|LNC|Rift valley fever virus Ag|Rift valley fever virus Ag
C1147636|T201|COMP|31952-5|LNC|Rinderpest virus Ag|Rinderpest virus Ag
C1147637|T201|COMP|31953-3|LNC|Rinderpest virus Ag|Rinderpest virus Ag
C1147638|T201|COMP|31954-1|LNC|Rinderpest virus Ag|Rinderpest virus Ag
C1147639|T201|COMP|31955-8|LNC|Rubella virus Ag|Rubella virus Ag
C1147640|T201|COMP|31956-6|LNC|Rubella virus Ag|Rubella virus Ag
C1147641|T201|COMP|31957-4|LNC|Rubella virus Ag|Rubella virus Ag
C1147642|T201|COMP|31958-2|LNC|Rubella virus Ag|Rubella virus Ag
C1147643|T201|COMP|31959-0|LNC|Rubella virus Ag|Rubella virus Ag
C1147644|T201|COMP|31960-8|LNC|Rubella virus Ag|Rubella virus Ag
C1147645|T201|COMP|31961-6|LNC|Rubella virus Ag|Rubella virus Ag
C1147646|T201|COMP|31962-4|LNC|Rubella virus Ag|Rubella virus Ag
C1147647|T201|COMP|31963-2|LNC|Rubella virus Ag|Rubella virus Ag
C1147648|T201|COMP|31964-0|LNC|Rubella virus Ag|Rubella virus Ag
C1147649|T201|COMP|31965-7|LNC|Rubella virus Ag|Rubella virus Ag
C1147650|T201|COMP|31966-5|LNC|Rubella virus Ag|Rubella virus Ag
C1147651|T201|COMP|31967-3|LNC|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C1147652|T201|COMP|31968-1|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C1147653|T201|COMP|31969-9|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C1147654|T201|COMP|31970-7|LNC|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C1147655|T201|COMP|31971-5|LNC|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C1147656|T201|COMP|31972-3|LNC|Swine vesicular disease virus Ag|Swine vesicular disease virus Ag
C1147657|T201|COMP|31973-1|LNC|Swine vesicular disease virus Ag|Swine vesicular disease virus Ag
C1147658|T201|COMP|31974-9|LNC|Taenia hydatigena Ag|Taenia hydatigena Ag
C1147659|T201|COMP|31975-6|LNC|Taenia sp Ag|Taenia sp Ag
C1147660|T201|COMP|31976-4|LNC|Taylorella equigenitalis Ag|Taylorella equigenitalis Ag
C1147661|T201|COMP|31977-2|LNC|Transmissible gastroenteritis virus Ag|Transmissible gastroenteritis virus Ag
C1147662|T201|COMP|31978-0|LNC|Trichomonas vaginalis Ag|Trichomonas vaginalis Ag
C1147663|T201|COMP|31979-8|LNC|Trypanosoma evansi Ag|Trypanosoma evansi Ag
C1147664|T201|COMP|31980-6|LNC|Trypanosoma sp Ag|Trypanosoma sp Ag
C1147665|T201|COMP|31981-4|LNC|Varicella zoster virus Ag|Varicella zoster virus Ag
C1147666|T201|COMP|31982-2|LNC|Varicella zoster virus Ag|Varicella zoster virus Ag
C1147667|T201|COMP|31983-0|LNC|Venezuelan equine encephalitis virus Ag|Venezuelan equine encephalitis virus Ag
C1147668|T201|COMP|31984-8|LNC|Venezuelan equine encephalitis virus Ag|Venezuelan equine encephalitis virus Ag
C1147669|T201|COMP|31985-5|LNC|Vesicular stomatitis virus Ag|Vesicular stomatitis virus Ag
C1147670|T201|COMP|31986-3|LNC|Vesicular stomatitis virus Ag|Vesicular stomatitis virus Ag
C1147671|T201|COMP|31987-1|LNC|Western equine encephalitis virus Ag|Western equine encephalitis virus Ag
C1147672|T201|COMP|31988-9|LNC|Western equine encephalitis virus Ag|Western equine encephalitis virus Ag
C1147673|T201|COMP|31989-7|LNC|14-3-3 Ag|14-3-3 Ag
C1147674|T201|COMP|31990-5|LNC|14-3-3 Ag|14-3-3 Ag
C1147675|T201|COMP|31991-3|LNC|Acylcarnitine|Acylcarnitine
C1147676|T201|COMP|31992-1|LNC|Aldosterone|Aldosterone
C1147677|T201|COMP|31993-9|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C1147678|T201|COMP|31994-7|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1147679|T201|COMP|31995-4|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1147680|T201|COMP|31996-2|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1147681|T201|COMP|31997-0|LNC|Biotin|Biotin
C1147682|T201|COMP|31998-8|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C1147683|T201|COMP|31999-6|LNC|Broad casts|Broad casts
C1147684|T201|COMP|32000-2|LNC|Catecholamines|Catecholamines
C1147685|T201|COMP|32001-0|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1147686|T201|COMP|32002-8|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1147687|T201|COMP|32003-6|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1147688|T201|COMP|32004-4|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1147689|T201|COMP|32005-1|LNC|Chlamydia trachomatis B Ab|Chlamydia trachomatis B Ab
C1147690|T201|COMP|32006-9|LNC|Chlamydia trachomatis C Ab|Chlamydia trachomatis C Ab
C1147691|T201|COMP|32007-7|LNC|Chlamydia trachomatis G+F+K Ab|Chlamydia trachomatis G+F+K Ab
C1147692|T201|COMP|32008-5|LNC|Coproporphyrin/Creatinine|Coproporphyrin/Creatinine
C1147693|T201|COMP|32009-3|LNC|Cortisol.free/Creatinine|Cortisol.free/Creatinine
C1147694|T201|COMP|32010-1|LNC|Diuretics|Diuretics
C1147695|T201|COMP|32011-9|LNC|Ehrlichia sp Ab.IgG|Ehrlichia sp Ab.IgG
C1147696|T201|COMP|32012-7|LNC|Ehrlichia sp Ab.IgM|Ehrlichia sp Ab.IgM
C1147697|T201|COMP|32013-5|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1147698|T201|COMP|32014-3|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1147699|T201|COMP|32015-0|LNC|EPINEPHrine|EPINEPHrine
C1147700|T201|COMP|32016-8|LNC|Glucose|Glucose
C1147701|T201|COMP|32017-6|LNC|Hemoglobin.other/Hemoglobin.total|Hemoglobin.other/Hemoglobin.total
C1147702|T201|COMP|32018-4|LNC|Hepatitis A virus Ab.IgG|Hepatitis A virus Ab.IgG
C1147703|T201|COMP|32019-2|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C1147704|T201|COMP|32020-0|LNC|Homocysteine|Homocysteine
C1147705|T201|COMP|32021-8|LNC|HTLV I DNA|HTLV I DNA
C1147706|T201|COMP|32022-6|LNC|Hydroxyproline.free|Hydroxyproline.free
C1147707|T201|COMP|32023-4|LNC|Insulin-like growth factor-I|Insulin-like growth factor-I
C1147708|T201|COMP|32024-2|LNC|Magnesium|Magnesium
C1147709|T201|COMP|32025-9|LNC|Malignin Ab|Malignin Ab
C1147711|T201|COMP|32027-5|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1147712|T201|COMP|32028-3|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1147713|T201|COMP|32029-1|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1147714|T201|COMP|32030-9|LNC|Nitrate|Nitrate
C1147715|T201|COMP|32031-7|LNC|Phosphatidylserine Ab.IgA|Phosphatidylserine Ab.IgA
C1147716|T201|COMP|32032-5|LNC|Phosphatidylserine Ab.IgG|Phosphatidylserine Ab.IgG
C1147717|T201|COMP|32033-3|LNC|Phosphatidylserine Ab.IgM|Phosphatidylserine Ab.IgM
C1147718|T201|COMP|32034-1|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1147719|T201|COMP|32035-8|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1147720|T201|COMP|32036-6|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1147721|T201|COMP|32037-4|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1147722|T201|COMP|32038-2|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1147723|T201|COMP|32039-0|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1147724|T201|COMP|32040-8|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C1147726|T201|COMP|32042-4|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C1147727|T201|COMP|32043-2|LNC|Uroporphyrin/Creatinine|Uroporphyrin/Creatinine
C1147728|T201|COMP|32044-0|LNC|Volatiles|Volatiles
C1147729|T201|COMP|32045-7|LNC|Parathyrin.biointact|Parathyrin.biointact
C1147730|T201|COMP|32046-5|LNC|Pregnancy associated plasma protein A|Pregnancy associated plasma protein A
C1147732|T201|COMP|32048-1|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C1147733|T201|COMP|32049-9|LNC|Amobarbital|Amobarbital
C1147734|T201|COMP|32050-7|LNC|Barbital|Barbital
C1147735|T201|COMP|32051-5|LNC|Barbital|Barbital
C1147736|T201|COMP|32052-3|LNC|Benzodiazepines|Benzodiazepines
C1147737|T201|COMP|32053-1|LNC|Bupivacaine|Bupivacaine
C1147738|T201|COMP|32054-9|LNC|Butabarbital|Butabarbital
C1147739|T201|COMP|32055-6|LNC|Butalbital|Butalbital
C1147740|T201|COMP|32056-4|LNC|Butalbital|Butalbital
C1147741|T201|COMP|32057-2|LNC|Butalbital|Butalbital
C1147742|T201|COMP|32058-0|LNC|carBAMazepine.free|carBAMazepine.free
C1147743|T201|COMP|32059-8|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C1147744|T201|COMP|32060-6|LNC|Chloroquine|Chloroquine
C1147745|T201|COMP|32061-4|LNC|chlorproMAZINE|chlorproMAZINE
C1147746|T201|COMP|32062-2|LNC|chlorproPAMIDE|chlorproPAMIDE
C1147747|T201|COMP|32063-0|LNC|Cimetidine|Cimetidine
C1147748|T201|COMP|32064-8|LNC|Clorazepate|Clorazepate
C1147749|T201|COMP|32065-5|LNC|cloZAPine|cloZAPine
C1147750|T201|COMP|32066-3|LNC|cloZAPine|cloZAPine
C1147751|T201|COMP|32067-1|LNC|Digoxin.free|Digoxin.free
C1147752|T201|COMP|32068-9|LNC|diphenhydrAMINE+Dimenhydrinate|diphenhydrAMINE+Dimenhydrinate
C1147753|T201|COMP|32069-7|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C1147754|T201|COMP|32070-5|LNC|Ethanol|Ethanol
C1147755|T201|COMP|32071-3|LNC|Ethchlorvynol|Ethchlorvynol
C1147756|T201|COMP|32072-1|LNC|FLUoxetine|FLUoxetine
C1147757|T201|COMP|32073-9|LNC|fluvoxaMINE|fluvoxaMINE
C1147758|T201|COMP|32074-7|LNC|fluvoxaMINE|fluvoxaMINE
C1147759|T201|COMP|32075-4|LNC|fluvoxaMINE|fluvoxaMINE
C1147760|T201|COMP|32076-2|LNC|Glutethimide|Glutethimide
C1147761|T201|COMP|32077-0|LNC|Glutethimide|Glutethimide
C1147762|T201|COMP|32078-8|LNC|glyBURIDE|glyBURIDE
C1147763|T201|COMP|32079-6|LNC|Gold|Gold
C1147764|T201|COMP|32080-4|LNC|HYDROcodone|HYDROcodone
C1147765|T201|COMP|32081-2|LNC|HYDROmorphone|HYDROmorphone
C1147766|T201|COMP|32082-0|LNC|Ibuprofen|Ibuprofen
C1147767|T201|COMP|32083-8|LNC|Imipramine+Desipramine|Imipramine+Desipramine
C1147768|T201|COMP|32084-6|LNC|Isopropanol|Isopropanol
C1147769|T201|COMP|32085-3|LNC|Isopropanol|Isopropanol
C1147770|T201|COMP|32086-1|LNC|Lidocaine|Lidocaine
C1147771|T201|COMP|32087-9|LNC|Loxapine|Loxapine
C1147772|T201|COMP|32088-7|LNC|Meperidine|Meperidine
C1147773|T201|COMP|32089-5|LNC|Mephobarbital|Mephobarbital
C1147774|T201|COMP|32090-3|LNC|Mepivacaine|Mepivacaine
C1147775|T201|COMP|32091-1|LNC|Meprobamate|Meprobamate
C1147776|T201|COMP|32092-9|LNC|Meprobamate|Meprobamate
C1147777|T201|COMP|32093-7|LNC|Methadone|Methadone
C1147778|T201|COMP|32094-5|LNC|Methanol|Methanol
C1147779|T201|COMP|32095-2|LNC|Methanol|Methanol
C1147780|T201|COMP|32096-0|LNC|Methaqualone|Methaqualone
C1147781|T201|COMP|32097-8|LNC|Methyprylon|Methyprylon
C1147782|T201|COMP|32098-6|LNC|Mexiletine|Mexiletine
C1147783|T201|COMP|32099-4|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C1147784|T201|COMP|32100-0|LNC|Morphine|Morphine
C1147785|T201|COMP|32101-8|LNC|oxyCODONE|oxyCODONE
C1147786|T201|COMP|32102-6|LNC|PARoxetine|PARoxetine
C1147787|T201|COMP|32103-4|LNC|PENTobarbital|PENTobarbital
C1147788|T201|COMP|32104-2|LNC|PENTobarbital|PENTobarbital
C1147789|T201|COMP|32105-9|LNC|Perphenazine|Perphenazine
C1147790|T201|COMP|32106-7|LNC|Perphenazine|Perphenazine
C1147791|T201|COMP|32107-5|LNC|Phencyclidine|Phencyclidine
C1147792|T201|COMP|32108-3|LNC|PHENobarbital|PHENobarbital
C1147793|T201|COMP|32109-1|LNC|Phenytoin.free|Phenytoin.free
C1147794|T201|COMP|32110-9|LNC|Procyclidine|Procyclidine
C1147795|T201|COMP|32111-7|LNC|Secobarbital|Secobarbital
C1147796|T201|COMP|32112-5|LNC|Sertraline|Sertraline
C1147797|T201|COMP|32113-3|LNC|Sertraline|Sertraline
C1147798|T201|COMP|32114-1|LNC|Thallium|Thallium
C1147799|T201|COMP|32115-8|LNC|Theophylline^peak|Theophylline^peak
C1147800|T201|COMP|32116-6|LNC|Theophylline^trough|Theophylline^trough
C1147801|T201|COMP|32117-4|LNC|Thiopental|Thiopental
C1147802|T201|COMP|32118-2|LNC|TOLBUTamide|TOLBUTamide
C1147803|T201|COMP|32119-0|LNC|Valproate.free|Valproate.free
C1147804|T201|COMP|32120-8|LNC|Venlafaxine|Venlafaxine
C1147805|T201|COMP|32121-6|LNC|Venlafaxine|Venlafaxine
C1147806|T201|COMP|32122-4|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C1147807|T201|COMP|32123-2|LNC|Pregnancy associated plasma protein A|Pregnancy associated plasma protein A
C1147808|T201|COMP|32124-0|LNC|Bromazepam|Bromazepam
C1147809|T201|COMP|32125-7|LNC|Propoxyphene|Propoxyphene
C1147810|T201|COMP|32126-5|LNC|Propylene glycol|Propylene glycol
C1147811|T201|COMP|32127-3|LNC|raNITIdine|raNITIdine
C1147812|T201|COMP|32128-1|LNC|risperiDONE|risperiDONE
C1147813|T201|COMP|32129-9|LNC|risperiDONE|risperiDONE
C1147814|T201|COMP|32130-7|LNC|risperiDONE|risperiDONE
C1147815|T201|COMP|32131-5|LNC|Hantavirus Ab.IgM|Hantavirus Ab.IgM
C1147816|T201|COMP|32132-3|LNC|Lactate|Lactate
C1147817|T201|COMP|32133-1|LNC|Lactate|Lactate
C1147818|T201|COMP|32134-9|LNC|Adenovirus+Rotavirus|Adenovirus+Rotavirus
C1147819|T201|COMP|32135-6|LNC|Alkaline phosphatase.liver|Alkaline phosphatase.liver
C1147820|T201|COMP|32136-4|LNC|Antidepressants|Antidepressants
C1147821|T201|COMP|32137-2|LNC|Calcium phosphate/Total|Calcium phosphate/Total
C1147822|T201|COMP|32138-0|LNC|Cystine/Total|Cystine/Total
C1147823|T201|COMP|32139-8|LNC|Haemophilus influenzae Ag|Haemophilus influenzae Ag
C1147824|T201|COMP|32140-6|LNC|Hemoglobin F|Hemoglobin F
C1147825|T201|COMP|32141-4|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1147826|T201|COMP|32142-2|LNC|Leukocytes|Leukocytes
C1147827|T201|COMP|32143-0|LNC|Triple phosphate/Total|Triple phosphate/Total
C1147828|T201|COMP|32144-8|LNC|Pathologist review|Pathologist review
C1147829|T201|COMP|32145-5|LNC|Phosphate crystals.amorphous|Phosphate crystals.amorphous
C1147830|T201|COMP|32146-3|LNC|Platelets.large|Platelets.large
C1147831|T201|COMP|32147-1|LNC|Reducing substances|Reducing substances
C1147832|T201|COMP|32148-9|LNC|Substance.toxic identified|Substance.toxic identified
C1147833|T201|COMP|32149-7|LNC|Urate/Total|Urate/Total
C1147834|T201|COMP|32150-5|LNC|Urate crystals.amorphous|Urate crystals.amorphous
C1147836|T201|COMP|32152-1|LNC|17-Hydroxyketosteroids|17-Hydroxyketosteroids
C1147837|T201|COMP|32153-9|LNC|Alpha-Phenyl-2-Piperidine acetate|Alpha-Phenyl-2-Piperidine acetate
C1147838|T201|COMP|32154-7|LNC|Basophils+Eosinophils+Monocytes|Basophils+Eosinophils+Monocytes
C1147839|T201|COMP|32155-4|LNC|Basophils+Eosinophils+Monocytes/100 leukocytes|Basophils+Eosinophils+Monocytes/100 leukocytes
C1147840|T201|COMP|32156-2|LNC|Calcium carbonate/Total|Calcium carbonate/Total
C1147841|T201|COMP|32157-0|LNC|Calcium oxalate/Total|Calcium oxalate/Total
C1147842|T201|COMP|32158-8|LNC|Klebsiella granulomatis|Klebsiella granulomatis
C1147843|T201|COMP|32159-6|LNC|Carbonated calcium phosphate/Total|Carbonated calcium phosphate/Total
C1147844|T201|COMP|32160-4|LNC|Carboxyhemoglobin|Carboxyhemoglobin
C1147845|T201|COMP|32161-2|LNC|Catecholamines|Catecholamines
C1147846|T201|COMP|32162-0|LNC|Cells|Cells
C1147847|T201|COMP|32163-8|LNC|Cells|Cells
C1147848|T201|COMP|32164-6|LNC|Cells|Cells
C1147849|T201|COMP|32165-3|LNC|Cells counted.total|Cells counted.total
C1147850|T201|COMP|32166-1|LNC|Choriogonadotropin^^adjusted|Choriogonadotropin^^adjusted
C1147851|T201|COMP|32167-9|LNC|Clarity|Clarity
C1147852|T201|COMP|32168-7|LNC|Color|Color
C1147853|T201|COMP|32169-5|LNC|Cystine|Cystine
C1147854|T201|COMP|32170-3|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C1147855|T201|COMP|32171-1|LNC|Echinococcus sp Ab.IgG|Echinococcus sp Ab.IgG
C1147856|T201|COMP|32172-9|LNC|Ehrlichia chaffeensis Ab|Ehrlichia chaffeensis Ab
C1147857|T201|COMP|32173-7|LNC|Eosinophils|Eosinophils
C1147858|T201|COMP|32174-5|LNC|Glucose|Glucose
C1147859|T201|COMP|32175-2|LNC|Granular casts.coarse|Granular casts.coarse
C1147860|T201|COMP|32176-0|LNC|Granular casts.fine|Granular casts.fine
C1147861|T201|COMP|32177-8|LNC|Granulocytes/100 leukocytes|Granulocytes/100 leukocytes
C1147862|T201|COMP|32178-6|LNC|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C1147863|T201|COMP|32179-4|LNC|Heptacarboxylporphyrin/Creatinine|Heptacarboxylporphyrin/Creatinine
C1147864|T201|COMP|32180-2|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C1147865|T201|COMP|32181-0|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C1147866|T201|COMP|32182-8|LNC|Herpes virus 6 Ab.IgM|Herpes virus 6 Ab.IgM
C1147867|T201|COMP|32183-6|LNC|Hydroxyproline.free|Hydroxyproline.free
C1147868|T201|COMP|32184-4|LNC|Itraconazole^peak|Itraconazole^peak
C1147869|T201|COMP|32185-1|LNC|Itraconazole^trough|Itraconazole^trough
C1147875|T201|COMP|32191-9|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1147876|T201|COMP|32192-7|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1147877|T201|COMP|32193-5|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1147878|T201|COMP|32194-3|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1147879|T201|COMP|32195-0|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1147880|T201|COMP|32196-8|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1147881|T201|COMP|32197-6|LNC|Myoglobin|Myoglobin
C1147882|T201|COMP|32198-4|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1147883|T201|COMP|32199-2|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1147884|T201|COMP|32200-8|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C1147885|T201|COMP|32201-6|LNC|Unidentified cells|Unidentified cells
C1147886|T201|COMP|32202-4|LNC|Unidentified cells|Unidentified cells
C1147887|T201|COMP|32203-2|LNC|Unidentified cells|Unidentified cells
C1147888|T201|COMP|32204-0|LNC|Unidentified cells|Unidentified cells
C1147889|T201|COMP|32205-7|LNC|Unidentified cells|Unidentified cells
C1147890|T201|COMP|32206-5|LNC|Plasmodium sp identified|Plasmodium sp identified
C1147891|T201|COMP|32207-3|LNC|Platelet distribution width|Platelet distribution width
C1147892|T201|COMP|32208-1|LNC|Platelets.small|Platelets.small
C1147893|T201|COMP|32209-9|LNC|Protein|Protein
C1147894|T201|COMP|32210-7|LNC|Protein pattern|Protein pattern
C1147895|T201|COMP|32211-5|LNC|Reducing substances|Reducing substances
C1147896|T201|COMP|32212-3|LNC|Salmonella paratyphi A Ab|Salmonella paratyphi A Ab
C1147897|T201|COMP|32213-1|LNC|Salmonella paratyphi B Ab|Salmonella paratyphi B Ab
C1147898|T201|COMP|32214-9|LNC|Thyroid stimulating immunoglobulins|Thyroid stimulating immunoglobulins
C1147899|T201|COMP|32215-6|LNC|Thyroxine free index|Thyroxine free index
C1147900|T201|COMP|32216-4|LNC|Uroporphyrin|Uroporphyrin
C1147901|T201|COMP|32217-2|LNC|von Willebrand factor multimers|von Willebrand factor multimers
C1147902|T201|COMP|32218-0|LNC|Cyclic citrullinated peptide Ab|Cyclic citrullinated peptide Ab
C1147903|T201|COMP|32219-8|LNC|Soluble liver Ab|Soluble liver Ab
C1147904|T201|COMP|32220-6|LNC|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C1147905|T201|COMP|32221-4|LNC|Alanine|Alanine
C1147906|T201|COMP|32222-2|LNC|Alanine|Alanine
C1147907|T201|COMP|32223-0|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C1147908|T201|COMP|32224-8|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C1147909|T201|COMP|32225-5|LNC|Arginine|Arginine
C1147910|T201|COMP|32226-3|LNC|Arginine|Arginine
C1147911|T201|COMP|32227-1|LNC|Argininosuccinate|Argininosuccinate
C1147912|T201|COMP|32228-9|LNC|Argininosuccinate|Argininosuccinate
C1147913|T201|COMP|32229-7|LNC|Argininosuccinate/Creatinine|Argininosuccinate/Creatinine
C1147914|T201|COMP|32230-5|LNC|Asparagine|Asparagine
C1147915|T201|COMP|32231-3|LNC|Aspartate|Aspartate
C1147916|T201|COMP|32232-1|LNC|Aspartate|Aspartate
C1147917|T201|COMP|32233-9|LNC|Carbamoyl phosphate synthetase|Carbamoyl phosphate synthetase
C1147918|T201|COMP|32234-7|LNC|Citrulline|Citrulline
C1147919|T201|COMP|32235-4|LNC|Citrulline|Citrulline
C1147920|T201|COMP|32236-2|LNC|Cystathionine|Cystathionine
C1147921|T201|COMP|32237-0|LNC|Cystine|Cystine
C1147922|T201|COMP|32238-8|LNC|Cystine|Cystine
C1147923|T201|COMP|32239-6|LNC|Ethanolamine|Ethanolamine
C1147924|T201|COMP|32240-4|LNC|Fructose|Fructose
C1147925|T201|COMP|32241-2|LNC|Glutamate|Glutamate
C1147926|T201|COMP|32242-0|LNC|Glutamine|Glutamine
C1147927|T201|COMP|32243-8|LNC|Glutamine|Glutamine
C1147928|T201|COMP|32244-6|LNC|Glycine|Glycine
C1147929|T201|COMP|32245-3|LNC|Glycine|Glycine
C1147930|T201|COMP|32246-1|LNC|Histidine|Histidine
C1147931|T201|COMP|32247-9|LNC|Histidine|Histidine
C1147932|T201|COMP|32248-7|LNC|Homocitrulline/Creatinine|Homocitrulline/Creatinine
C1147933|T201|COMP|32249-5|LNC|Hydroxyproline|Hydroxyproline
C1147934|T201|COMP|32250-3|LNC|Hydroxyproline|Hydroxyproline
C1147935|T201|COMP|32251-1|LNC|Isoleucine|Isoleucine
C1147936|T201|COMP|32252-9|LNC|Isoleucine|Isoleucine
C1147937|T201|COMP|32253-7|LNC|Leucine|Leucine
C1147938|T201|COMP|32254-5|LNC|Leucine|Leucine
C1147939|T201|COMP|32255-2|LNC|Lysine|Lysine
C1147940|T201|COMP|32256-0|LNC|Lysine|Lysine
C1147941|T201|COMP|32257-8|LNC|Methionine|Methionine
C1147942|T201|COMP|32258-6|LNC|Methionine|Methionine
C1147943|T201|COMP|32259-4|LNC|Methylmalonate|Methylmalonate
C1147944|T201|COMP|32260-2|LNC|Ornithine|Ornithine
C1147945|T201|COMP|32261-0|LNC|Ornithine|Ornithine
C1147946|T201|COMP|32262-8|LNC|Orotate/Creatinine|Orotate/Creatinine
C1147947|T201|COMP|32263-6|LNC|Phenylalanine|Phenylalanine
C1147948|T201|COMP|32264-4|LNC|Phenylalanine|Phenylalanine
C1147949|T201|COMP|32265-1|LNC|Phenylalanine/Tyrosine|Phenylalanine/Tyrosine
C1147950|T201|COMP|32266-9|LNC|Proline|Proline
C1147951|T201|COMP|32267-7|LNC|Proline|Proline
C1147952|T201|COMP|32268-5|LNC|Ribose|Ribose
C1147953|T201|COMP|32269-3|LNC|Serine|Serine
C1147954|T201|COMP|32270-1|LNC|Serine|Serine
C1147955|T201|COMP|32271-9|LNC|Taurine|Taurine
C1147956|T201|COMP|32272-7|LNC|Threonine|Threonine
C1147957|T201|COMP|32273-5|LNC|Threonine|Threonine
C1147958|T201|COMP|32274-3|LNC|Thiosulfate/Creatinine|Thiosulfate/Creatinine
C1147959|T201|COMP|32275-0|LNC|Tryptophan|Tryptophan
C1147960|T201|COMP|32276-8|LNC|Tyrosine|Tyrosine
C1147961|T201|COMP|32277-6|LNC|Tyrosine|Tyrosine
C1147962|T201|COMP|32278-4|LNC|Valine|Valine
C1147963|T201|COMP|32279-2|LNC|Valine|Valine
C1147964|T201|COMP|32280-0|LNC|Acylglycines|Acylglycines
C1147965|T201|COMP|32281-8|LNC|Carnitine.free (C0)/Carnitine.total|Carnitine.free (C0)/Carnitine.total
C1147966|T201|COMP|32282-6|LNC|Succinylpurines|Succinylpurines
C1147967|T201|COMP|32283-4|LNC|Valproate.free/Valproate.total|Valproate.free/Valproate.total
C1147968|T201|COMP|32284-2|LNC|BK virus DNA|BK virus DNA
C1147969|T201|COMP|32285-9|LNC|BK virus DNA|BK virus DNA
C1147970|T201|COMP|32286-7|LNC|Hepatitis C virus genotype|Hepatitis C virus genotype
C1147971|T201|COMP|32287-5|LNC|Methylmalonate|Methylmalonate
C1147972|T201|COMP|32288-3|LNC|17-Hydroxyprogesterone^baseline|17-Hydroxyprogesterone^baseline
C1147973|T201|COMP|32289-1|LNC|7-Dehydrocholesterol|7-Dehydrocholesterol
C1147974|T201|COMP|32290-9|LNC|Acetone|Acetone
C1147975|T201|COMP|32291-7|LNC|Acetone|Acetone
C1147976|T201|COMP|32292-5|LNC|Acetone|Acetone
C1147977|T201|COMP|32293-3|LNC|Albumin|Albumin
C1147978|T201|COMP|32294-1|LNC|Albumin/Creatinine|Albumin/Creatinine
C1147979|T201|COMP|32295-8|LNC|Aluminum|Aluminum
C1147980|T201|COMP|32296-6|LNC|Amino acid pattern|Amino acid pattern
C1147981|T201|COMP|32297-4|LNC|Amino acids|Amino acids
C1147982|T201|COMP|32298-2|LNC|Amylase|Amylase
C1147983|T201|COMP|32299-0|LNC|Androstenedione^baseline|Androstenedione^baseline
C1147984|T201|COMP|32300-6|LNC|Base excess|Base excess
C1147985|T201|COMP|32301-4|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C1147986|T201|COMP|32302-2|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C1147987|T201|COMP|32303-0|LNC|Bilirubin|Bilirubin
C1147988|T201|COMP|32304-8|LNC|Cadmium|Cadmium
C1147989|T201|COMP|32305-5|LNC|Calcium|Calcium
C1147990|T201|COMP|32306-3|LNC|Carbon dioxide|Carbon dioxide
C1147991|T201|COMP|32307-1|LNC|Chloride|Chloride
C1147992|T201|COMP|32308-9|LNC|Cholesterol|Cholesterol
C1147993|T201|COMP|32309-7|LNC|Cholesterol.total/Cholesterol.in HDL|Cholesterol.total/Cholesterol.in HDL
C1147994|T201|COMP|32310-5|LNC|Cortisol|Cortisol
C1147995|T201|COMP|32311-3|LNC|Cortisol^1H post XXX challenge|Cortisol^1H post XXX challenge
C1147996|T201|COMP|32312-1|LNC|Cortisol^2H post XXX challenge|Cortisol^2H post XXX challenge
C1147997|T201|COMP|32313-9|LNC|Cortisol^30M post XXX challenge|Cortisol^30M post XXX challenge
C1147998|T201|COMP|32314-7|LNC|Cortisol^1.5H post XXX challenge|Cortisol^1.5H post XXX challenge
C1147999|T201|COMP|32315-4|LNC|Cortisol^baseline|Cortisol^baseline
C1148000|T201|COMP|32316-2|LNC|Follitropin^30M post XXX challenge|Follitropin^30M post XXX challenge
C1148001|T201|COMP|32317-0|LNC|Follitropin^baseline|Follitropin^baseline
C1148002|T201|COMP|32318-8|LNC|Glucose|Glucose
C1148003|T201|COMP|32319-6|LNC|Glucose^30M post 75 g glucose PO|Glucose^30M post 75 g glucose PO
C1148004|T201|COMP|32320-4|LNC|Glucose^3H post 75 g glucose PO|Glucose^3H post 75 g glucose PO
C1148005|T201|COMP|32321-2|LNC|Glucose^4H post 75 g glucose PO|Glucose^4H post 75 g glucose PO
C1148006|T201|COMP|32322-0|LNC|Glucose^5H post 75 g glucose PO|Glucose^5H post 75 g glucose PO
C1148007|T201|COMP|32323-8|LNC|Ketones|Ketones
C1148008|T201|COMP|32324-6|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C1148009|T201|COMP|32325-3|LNC|Lead|Lead
C1148010|T201|COMP|32326-1|LNC|Lutropin^30M post XXX challenge|Lutropin^30M post XXX challenge
C1148011|T201|COMP|32327-9|LNC|Lutropin^1H post XXX challenge|Lutropin^1H post XXX challenge
C1148012|T201|COMP|32328-7|LNC|Lutropin^baseline|Lutropin^baseline
C1148013|T201|COMP|32329-5|LNC|Magnesium|Magnesium
C1148014|T201|COMP|32330-3|LNC|Mercury|Mercury
C1148015|T201|COMP|32331-1|LNC|Myoglobin|Myoglobin
C1148016|T201|COMP|32332-9|LNC|Neopterin/Biopterin|Neopterin/Biopterin
C1148017|T201|COMP|32333-7|LNC|Phenylpropanolamine|Phenylpropanolamine
C1148018|T201|COMP|32334-5|LNC|Pipecolate|Pipecolate
C1148019|T201|COMP|32335-2|LNC|Pipecolate|Pipecolate
C1148020|T201|COMP|32336-0|LNC|Potassium|Potassium
C1148021|T201|COMP|32337-8|LNC|Protein|Protein
C1148022|T201|COMP|32338-6|LNC|Pyruvate|Pyruvate
C1148023|T201|COMP|32339-4|LNC|Serotonin|Serotonin
C1148024|T201|COMP|32340-2|LNC|Sodium|Sodium
C1148025|T201|COMP|32341-0|LNC|Transcobalamin II|Transcobalamin II
C1148026|T201|COMP|32342-8|LNC|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C1148027|T201|COMP|32343-6|LNC|Urate|Urate
C1148028|T201|COMP|32344-4|LNC|Urobilin|Urobilin
C1148029|T201|COMP|32345-1|LNC|Uroporphyrin|Uroporphyrin
C1148030|T201|COMP|32346-9|LNC|Uroporphyrin|Uroporphyrin
C1148031|T201|COMP|32347-7|LNC|Xylose|Xylose
C1148032|T201|COMP|32348-5|LNC|Zinc|Zinc
C1148033|T201|COMP|32349-3|LNC|Basophils+Eosinophils+Monocytes|Basophils+Eosinophils+Monocytes
C1148034|T201|COMP|32350-1|LNC|Basophils+Eosinophils+Monocytes/100 leukocytes|Basophils+Eosinophils+Monocytes/100 leukocytes
C1148035|T201|COMP|32351-9|LNC|Alkaline phosphatase.heat labile|Alkaline phosphatase.heat labile
C1148036|T201|COMP|32352-7|LNC|Alkaline phosphatase.heat stable|Alkaline phosphatase.heat stable
C1148037|T201|COMP|32353-5|LNC|Estriol|Estriol
C1148038|T201|COMP|32354-3|LNC|Hematocrit|Hematocrit
C1148039|T201|COMP|32355-0|LNC|Bacteria identified|Bacteria identified
C1148040|T201|COMP|32356-8|LNC|Yeast|Yeast
C1148041|T201|COMP|32357-6|LNC|Ova+Parasites identified|Ova+Parasites identified
C1148042|T201|COMP|32358-4|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C1148043|T201|COMP|32359-2|LNC|Glucose^10M post dose glucose|Glucose^10M post dose glucose
C1148044|T201|COMP|32360-0|LNC|Insulin^10M post XXX challenge|Insulin^10M post XXX challenge
C1148045|T201|COMP|32361-8|LNC|West Nile virus RNA|West Nile virus RNA
C1148046|T201|COMP|32362-6|LNC|BK virus DNA|BK virus DNA
C1148047|T201|COMP|32363-4|LNC|JC virus DNA|JC virus DNA
C1148048|T201|COMP|32364-2|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1148049|T201|COMP|32365-9|LNC|Torque teno virus DNA|Torque teno virus DNA
C1148050|T201|COMP|32366-7|LNC|Hepatitis B virus genotype|Hepatitis B virus genotype
C1148051|T201|COMP|32367-5|LNC|Bacteria identified|Bacteria identified
C1148052|T201|COMP|32368-3|LNC|Ureaplasma sp identified|Ureaplasma sp identified
C1148053|T201|COMP|32369-1|LNC|Clostridium perfringens enterotoxin|Clostridium perfringens enterotoxin
C1148054|T201|COMP|32370-9|LNC|West Nile virus RNA|West Nile virus RNA
C1148055|T201|COMP|32371-7|LNC|West Nile virus Ag|West Nile virus Ag
C1148056|T201|COMP|32372-5|LNC|Fleroxacin|Fleroxacin
C1148057|T201|COMP|32373-3|LNC|Arbekacin|Arbekacin
C1148058|T201|COMP|32374-1|LNC|Cefotiam|Cefotiam
C1148059|T201|COMP|32375-8|LNC|Cefmenoxime|Cefmenoxime
C1148061|T201|COMP|32377-4|LNC|Cefetamet|Cefetamet
C1148062|T201|COMP|32378-2|LNC|Caspofungin|Caspofungin
C1148063|T201|COMP|32379-0|LNC|Voriconazole|Voriconazole
C1148064|T201|COMP|18916-7|LNC|Dicloxacillin|Dicloxacillin
C1148065|T201|COMP|32381-6|LNC|Isepamicin|Isepamicin
C1148066|T201|COMP|25608-1|LNC|Nitroxoline|Nitroxoline
C1148067|T201|COMP|32383-2|LNC|Pristinamycin|Pristinamycin
C1148068|T201|COMP|32384-0|LNC|Thiacetazone|Thiacetazone
C1148177|T201|COMP|32493-9|LNC|Cells.CD25/100 cells|Cells.CD25/100 cells
C1148178|T201|COMP|32494-7|LNC|Cells.CD25/100 cells|Cells.CD25/100 cells
C1148179|T201|COMP|32495-4|LNC|Cells.CD25/100 cells|Cells.CD25/100 cells
C1148180|T201|COMP|32496-2|LNC|Cells.CD57/100 cells|Cells.CD57/100 cells
C1148181|T201|COMP|32497-0|LNC|Cells.CD57/100 cells|Cells.CD57/100 cells
C1148182|T201|COMP|32498-8|LNC|Cells.CD57/100 cells|Cells.CD57/100 cells
C1148183|T201|COMP|32499-6|LNC|Cells.CD7-CD13+CD33+/100 cells|Cells.CD7-CD13+CD33+/100 cells
C1148184|T201|COMP|32500-1|LNC|Cells.CD10+CD19+/100 cells|Cells.CD10+CD19+/100 cells
C1148185|T201|COMP|32501-9|LNC|Cells.CD10+CD19+/100 cells|Cells.CD10+CD19+/100 cells
C1148186|T201|COMP|32502-7|LNC|Cells.CD10+CD19+/100 cells|Cells.CD10+CD19+/100 cells
C1148187|T201|COMP|33582-8|LNC|Cells.CD13+CD33+|Cells.CD13+CD33+
C1148188|T201|COMP|32504-3|LNC|Cells.CD13+CD33+/100 cells|Cells.CD13+CD33+/100 cells
C1148189|T201|COMP|32505-0|LNC|Cells.CD13+CD33+/100 cells|Cells.CD13+CD33+/100 cells
C1148190|T201|COMP|32506-8|LNC|Cells.CD14/100 cells|Cells.CD14/100 cells
C1148191|T201|COMP|32507-6|LNC|Cells.CD14/100 cells|Cells.CD14/100 cells
C1148192|T201|COMP|32508-4|LNC|Cells.CD3-CD16+CD56+/100 cells|Cells.CD3-CD16+CD56+/100 cells
C1148193|T201|COMP|32509-2|LNC|Cells.CD3-CD16+CD56+/100 cells|Cells.CD3-CD16+CD56+/100 cells
C1148194|T201|COMP|32510-0|LNC|Cells.CD5+CD19+/100 cells|Cells.CD5+CD19+/100 cells
C1148195|T201|COMP|32511-8|LNC|Cells.CD5+CD19+/100 cells|Cells.CD5+CD19+/100 cells
C1148196|T201|COMP|32512-6|LNC|Cells.CD2|Cells.CD2
C1148197|T201|COMP|32513-4|LNC|Cells.CD3+CD25+|Cells.CD3+CD25+
C1148198|T201|COMP|32514-2|LNC|Cells.CD3+CD25+/100 cells|Cells.CD3+CD25+/100 cells
C1148199|T201|COMP|32515-9|LNC|Cells.CD3+CD4+|Cells.CD3+CD4+
C1148200|T201|COMP|32516-7|LNC|Cells.CD3+CD4+/100 cells|Cells.CD3+CD4+/100 cells
C1148201|T201|COMP|32517-5|LNC|Cells.CD3+CD8+|Cells.CD3+CD8+
C1148202|T201|COMP|32518-3|LNC|Cells.CD3+CD8+/100 cells|Cells.CD3+CD8+/100 cells
C1148203|T201|COMP|32519-1|LNC|Cells.CD3-CD16+CD56+/100 cells|Cells.CD3-CD16+CD56+/100 cells
C1148204|T201|COMP|32520-9|LNC|Cells.CD7-CD13+CD33+/100 cells|Cells.CD7-CD13+CD33+/100 cells
C1148205|T201|COMP|32521-7|LNC|Cells.CD10+CD19+/100 cells|Cells.CD10+CD19+/100 cells
C1148206|T201|COMP|32522-5|LNC|Cells.CD13+CD33+/100 cells|Cells.CD13+CD33+/100 cells
C1148207|T201|COMP|32523-3|LNC|Cells.CD5+CD19+/100 cells|Cells.CD5+CD19+/100 cells
C1148208|T201|COMP|32524-1|LNC|Cells.CD19|Cells.CD19
C1148209|T201|COMP|32525-8|LNC|Cells.CD19/100 cells|Cells.CD19/100 cells
C1148210|T201|COMP|32526-6|LNC|Cells.CD2|Cells.CD2
C1148211|T201|COMP|32527-4|LNC|Cells.CD2/100 cells|Cells.CD2/100 cells
C1148212|T201|COMP|32528-2|LNC|Cells.CD3|Cells.CD3
C1148213|T201|COMP|32529-0|LNC|Cells.CD3/100 cells|Cells.CD3/100 cells
C1148214|T201|COMP|32530-8|LNC|Cells.CD3+CD25+|Cells.CD3+CD25+
C1148215|T201|COMP|32531-6|LNC|Cells.CD3+CD25+/100 cells|Cells.CD3+CD25+/100 cells
C1148216|T201|COMP|32532-4|LNC|Cells.CD3+CD4+|Cells.CD3+CD4+
C1148217|T201|COMP|32533-2|LNC|Cells.CD3+CD4+/100 cells|Cells.CD3+CD4+/100 cells
C1148218|T201|COMP|32534-0|LNC|Cells.CD3+CD8+|Cells.CD3+CD8+
C1148219|T201|COMP|32535-7|LNC|Cells.CD3+CD8+/100 cells|Cells.CD3+CD8+/100 cells
C1148220|T201|COMP|32536-5|LNC|Cells.CD3-CD16+CD56+|Cells.CD3-CD16+CD56+
C1148221|T201|COMP|32537-3|LNC|Cells.CD3+CD4+/Cells.CD3+CD8+|Cells.CD3+CD4+/Cells.CD3+CD8+
C1148222|T201|COMP|32538-1|LNC|17-Hydroxyprogesterone^2H post XXX challenge|17-Hydroxyprogesterone^2H post XXX challenge
C1148223|T201|COMP|32539-9|LNC|17-Hydroxyprogesterone^1H post XXX challenge|17-Hydroxyprogesterone^1H post XXX challenge
C1148224|T201|COMP|32540-7|LNC|Glucosylceramidase|Glucosylceramidase
C1148225|T201|COMP|32541-5|LNC|Calcium|Calcium
C1148226|T201|COMP|32542-3|LNC|Chloride|Chloride
C1148227|T201|COMP|32543-1|LNC|Creatinine|Creatinine
C1148230|T201|COMP|32546-4|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C1148231|T201|COMP|32547-2|LNC|Ketones|Ketones
C1148232|T201|COMP|32548-0|LNC|Nitroprusside reacting substances|Nitroprusside reacting substances
C1148233|T201|COMP|32549-8|LNC|Norepinephrine/Creatinine|Norepinephrine/Creatinine
C1148234|T201|COMP|32550-6|LNC|Potassium|Potassium
C1148235|T201|COMP|32551-4|LNC|Protein|Protein
C1148236|T201|COMP|32552-2|LNC|Pyruvate kinase|Pyruvate kinase
C1148237|T201|COMP|32553-0|LNC|Sodium|Sodium
C1148238|T201|COMP|32554-8|LNC|Thiamine|Thiamine
C1148239|T201|COMP|32555-5|LNC|Urate|Urate
C1148240|T201|COMP|32556-3|LNC|Urea|Urea
C1148242|T201|COMP|32558-9|LNC|Mumps reaction wheal^1D post 0.1 mL mumps ID|Mumps reaction wheal^1D post 0.1 mL mumps ID
C1148243|T201|COMP|32559-7|LNC|Tau protein|Tau protein
C1148246|T201|COMP|32562-1|LNC|Lymphocytes.IgG/100 lymphocytes|Lymphocytes.IgG/100 lymphocytes
C1148247|T201|COMP|32563-9|LNC|Lymphocytes.IgG/100 lymphocytes|Lymphocytes.IgG/100 lymphocytes
C1148248|T201|COMP|32564-7|LNC|Cells.CD3+CD7+/100 cells|Cells.CD3+CD7+/100 cells
C1148249|T201|COMP|32565-4|LNC|SCA3 gene.CAG repeats|SCA3 gene.CAG repeats
C1148250|T201|COMP|32566-2|LNC|Coxiella burnetii Ab|Coxiella burnetii Ab
C1148253|T201|COMP|32569-6|LNC|Corynebacterium diphtheriae Ab^1st specimen|Corynebacterium diphtheriae Ab^1st specimen
C1148254|T201|COMP|32570-4|LNC|Tetrahydroaldosterone/Creatinine|Tetrahydroaldosterone/Creatinine
C1148255|T201|COMP|32571-2|LNC|HIV 1 Ab|HIV 1 Ab
C1148256|T201|COMP|32572-0|LNC|Tilapia Ab.IgE|Tilapia Ab.IgE
C1148257|T201|COMP|32573-8|LNC|Tilapia Ab.IgE.RAST class|Tilapia Ab.IgE.RAST class
C1148258|T201|COMP|32574-6|LNC|Zaleplon|Zaleplon
C1148259|T201|COMP|32575-3|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C1148260|T201|COMP|32576-1|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C1148261|T201|COMP|32577-9|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C1148262|T201|COMP|32578-7|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C1148263|T201|COMP|32579-5|LNC|Phentermine|Phentermine
C1148264|T201|COMP|32580-3|LNC|Chromatin Ab.IgG|Chromatin Ab.IgG
C1148265|T201|COMP|32581-1|LNC|Epidermal growth factor receptor Ag|Epidermal growth factor receptor Ag
C1148266|T201|COMP|32582-9|LNC|Phenylpropionylglycine|Phenylpropionylglycine
C1148267|T201|COMP|32583-7|LNC|Phenyllactate|Phenyllactate
C1148268|T201|COMP|32584-5|LNC|Propionylglycine|Propionylglycine
C1148269|T201|COMP|32585-2|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1148270|T201|COMP|32586-0|LNC|Follitropin^20M post XXX challenge|Follitropin^20M post XXX challenge
C1148271|T201|COMP|32587-8|LNC|Androstenedione^2H post XXX challenge|Androstenedione^2H post XXX challenge
C1148272|T201|COMP|32588-6|LNC|Androstenedione^1H post XXX challenge|Androstenedione^1H post XXX challenge
C1148274|T201|COMP|32590-2|LNC|Granulocytes units available|Granulocytes units available
C1148275|T201|COMP|32591-0|LNC|Heavy metals|Heavy metals
C1148276|T201|COMP|32592-8|LNC|Cryoprecipitate poor plasma units available|Cryoprecipitate poor plasma units available
C1148277|T201|COMP|32593-6|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1148278|T201|COMP|32594-4|LNC|Tacrolimus|Tacrolimus
C1148279|T201|COMP|32595-1|LNC|Topiramate|Topiramate
C1148280|T201|COMP|32596-9|LNC|Trifluoperazine|Trifluoperazine
C1148281|T201|COMP|32597-7|LNC|Natamycin|Natamycin
C1148282|T201|COMP|32598-5|LNC|Sertraline|Sertraline
C1148283|T201|COMP|32599-3|LNC|Lutropin^30M post XXX challenge|Lutropin^30M post XXX challenge
C1148284|T201|COMP|32600-9|LNC|Felbamate|Felbamate
C1148285|T201|COMP|32601-7|LNC|Cells.CD59/100 cells|Cells.CD59/100 cells
C1148286|T201|COMP|32602-5|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C1148287|T201|COMP|32603-3|LNC|Itraconazole|Itraconazole
C1148288|T201|COMP|32604-1|LNC|Leptospira sp Ab^1st specimen|Leptospira sp Ab^1st specimen
C1148289|T201|COMP|32605-8|LNC|Leptospira sp Ab^2nd specimen|Leptospira sp Ab^2nd specimen
C1148290|T201|COMP|32606-6|LNC|Lutropin^1H post XXX challenge|Lutropin^1H post XXX challenge
C1148292|T201|COMP|32608-2|LNC|cloZAPine|cloZAPine
C1148460|T201|COMP|20942-9|LNC|Plant identified|Plant identified
C1148462|T201|COMP|17942-4|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1148463|T201|COMP|17943-2|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1148464|T201|COMP|17944-0|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1148465|T201|COMP|17945-7|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1153739|T201|COMP|19049-6|LNC|Metanephrine|Metanephrine
C1153740|T201|COMP|17967-1|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1153741|T201|COMP|17966-3|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1153742|T201|COMP|17965-5|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1153743|T201|COMP|17964-8|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1153744|T201|COMP|17907-7|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1153745|T201|COMP|17906-9|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1153746|T201|COMP|17905-1|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1153747|T201|COMP|17904-4|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1153748|T201|COMP|17923-4|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1153749|T201|COMP|19214-6|LNC|Oxygen^^saturation adjusted to 0.5|Oxygen^^saturation adjusted to 0.5
C1153750|T201|COMP|19215-3|LNC|Oxygen^^saturation adjusted to 0.5|Oxygen^^saturation adjusted to 0.5
C1153751|T201|COMP|19216-1|LNC|Oxygen^^saturation adjusted to 0.5|Oxygen^^saturation adjusted to 0.5
C1153752|T201|COMP|17975-4|LNC|Virus identified^^^2|Virus identified^^^2
C1315083|T201|COMP|32609-0|LNC|Amino acids|Amino acids
C1315084|T201|COMP|32610-8|LNC|Amino acids|Amino acids
C1315085|T201|COMP|32611-6|LNC|Amino acids|Amino acids
C1315086|T201|COMP|32612-4|LNC|Amino acids|Amino acids
C1315087|T201|COMP|32613-2|LNC|Carnitine.free (C0)/Carnitine.total|Carnitine.free (C0)/Carnitine.total
C1315088|T201|COMP|32614-0|LNC|Glutamate|Glutamate
C1315089|T201|COMP|32615-7|LNC|Homocysteine cysteine disulfide|Homocysteine cysteine disulfide
C1315090|T201|COMP|32616-5|LNC|Homocysteine cysteine disulfide/Creatinine|Homocysteine cysteine disulfide/Creatinine
C1315091|T201|COMP|32617-3|LNC|Ornithine carbamoyltransferase|Ornithine carbamoyltransferase
C1315092|T201|COMP|32618-1|LNC|3-Methoxytyramine|3-Methoxytyramine
C1315093|T201|COMP|32619-9|LNC|Biotinidase|Biotinidase
C1315094|T201|COMP|32620-7|LNC|Corynebacterium diphtheriae Ab|Corynebacterium diphtheriae Ab
C1315095|T201|COMP|32621-5|LNC|HLA-DR|HLA-DR
C1315096|T201|COMP|32622-3|LNC|Hyaluronidase Ab|Hyaluronidase Ab
C1315099|T201|COMP|32625-6|LNC|Spermatozoa Ab.IgA|Spermatozoa Ab.IgA
C1315100|T201|COMP|32626-4|LNC|Spermatozoa Ab.IgG|Spermatozoa Ab.IgG
C1315101|T201|COMP|32627-2|LNC|Argininosuccinate lyase|Argininosuccinate lyase
C1315102|T201|COMP|32628-0|LNC|ACADM gene.c.985A>G|ACADM gene.c.985A>G
C1315103|T201|COMP|32629-8|LNC|Protein.monoclonal/Protein.total|Protein.monoclonal/Protein.total
C1315104|T201|COMP|32630-6|LNC|MSH2 gene+MLH1 gene targeted mutation analysis|MSH2 gene+MLH1 gene targeted mutation analysis
C1315105|T201|COMP|32631-4|LNC|Nitroblue tetrazolium test|Nitroblue tetrazolium test
C1315106|T201|COMP|32632-2|LNC|HEXA gene targeted mutation analysis|HEXA gene targeted mutation analysis
C1315107|T201|COMP|32633-0|LNC|Susceptibility organism^^^4|Susceptibility organism^^^4
C1315108|T201|COMP|32634-8|LNC|Metanephrine.free|Metanephrine.free
C1315109|T201|COMP|32635-5|LNC|Coagulation factor II inhibitor|Coagulation factor II inhibitor
C1315110|T201|COMP|32636-3|LNC|Islet cell 512 Ab|Islet cell 512 Ab
C1315111|T201|COMP|32637-1|LNC|Urease|Urease
C1315112|T201|COMP|32638-9|LNC|Blood group antibody screen|Blood group antibody screen
C1315113|T201|COMP|32639-7|LNC|FANCC gene targeted mutation analysis|FANCC gene targeted mutation analysis
C1315114|T201|COMP|32640-5|LNC|BLM gene targeted mutation analysis|BLM gene targeted mutation analysis
C1315115|T201|COMP|32641-3|LNC|SMPD1 gene targeted mutation analysis|SMPD1 gene targeted mutation analysis
C1315116|T201|COMP|32642-1|LNC|Dextroamphetamine/Levoamphetamine|Dextroamphetamine/Levoamphetamine
C1315117|T201|COMP|32643-9|LNC|Dextromethamphetamine/Levomethamphetamine|Dextromethamphetamine/Levomethamphetamine
C1315118|T201|COMP|32644-7|LNC|Coxiella burnetii phase 1 Ab.IgG|Coxiella burnetii phase 1 Ab.IgG
C1315119|T201|COMP|32645-4|LNC|Coxiella burnetii phase 1 Ab.IgM|Coxiella burnetii phase 1 Ab.IgM
C1315120|T201|COMP|32646-2|LNC|Nevirapine|Nevirapine
C1315121|T201|COMP|32647-0|LNC|Nelfinavir|Nelfinavir
C1315122|T201|COMP|32648-8|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C1315123|T201|COMP|32649-6|LNC|Hydroxytriazolam|Hydroxytriazolam
C1315124|T201|COMP|32650-4|LNC|Norflunitrazepam|Norflunitrazepam
C1315125|T201|COMP|32651-2|LNC|Ethion|Ethion
C1315126|T201|COMP|32652-0|LNC|Fenthion|Fenthion
C1315127|T201|COMP|32653-8|LNC|DYS gene targeted mutation analysis|DYS gene targeted mutation analysis
C1315128|T201|COMP|32654-6|LNC|6-Methylmercaptopurine|6-Methylmercaptopurine
C1315129|T201|COMP|35644-4|LNC|Metanephrine/Creatinine|Metanephrine/Creatinine
C1315130|T201|COMP|32656-1|LNC|Aflatoxin Ab.IgG|Aflatoxin Ab.IgG
C1315131|T201|COMP|32657-9|LNC|Aflatoxin Ab.IgA|Aflatoxin Ab.IgA
C1315132|T201|COMP|32658-7|LNC|Aflatoxin Ab.IgM|Aflatoxin Ab.IgM
C1315133|T201|COMP|32659-5|LNC|Aflatoxin Ab.IgE|Aflatoxin Ab.IgE
C1315134|T201|COMP|32660-3|LNC|6-Thioguanine|6-Thioguanine
C1315135|T201|COMP|32661-1|LNC|Adrenal Ab|Adrenal Ab
C1315136|T201|COMP|32662-9|LNC|Afipia felis Ab.IgG|Afipia felis Ab.IgG
C1315137|T201|COMP|32663-7|LNC|Afipia felis Ab.IgM|Afipia felis Ab.IgM
C1315138|T201|COMP|32664-5|LNC|Ammonia|Ammonia
C1315139|T201|COMP|32665-2|LNC|Anticonvulsants|Anticonvulsants
C1315140|T201|COMP|32666-0|LNC|Borrelia burgdorferi 25kD Ab.IgM|Borrelia burgdorferi 25kD Ab.IgM
C1315141|T201|COMP|32667-8|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C1315142|T201|COMP|32668-6|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C1315143|T201|COMP|32669-4|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C1315144|T201|COMP|32670-2|LNC|Cells counted.total|Cells counted.total
C1315145|T201|COMP|32671-0|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1315146|T201|COMP|32672-8|LNC|Cold agglutinin|Cold agglutinin
C1315147|T201|COMP|32673-6|LNC|Creatine kinase.MB|Creatine kinase.MB
C1315148|T201|COMP|32674-4|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1315149|T201|COMP|32675-1|LNC|Cytomegalovirus|Cytomegalovirus
C1315150|T201|COMP|32676-9|LNC|Diuretics|Diuretics
C1315151|T201|COMP|32677-7|LNC|DNA double strand Ab|DNA double strand Ab
C1315152|T201|COMP|32678-5|LNC|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C1315153|T201|COMP|32679-3|LNC|Ehrlichia chaffeensis Ab.IgM|Ehrlichia chaffeensis Ab.IgM
C1315154|T201|COMP|32680-1|LNC|Granular casts.fine|Granular casts.fine
C1315155|T201|COMP|32681-9|LNC|Hemoglobin C/Hemoglobin.total|Hemoglobin C/Hemoglobin.total
C1315156|T201|COMP|32682-7|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C1315157|T201|COMP|32683-5|LNC|Hemoglobin S/Hemoglobin.total|Hemoglobin S/Hemoglobin.total
C1315158|T201|COMP|32684-3|LNC|Heparin.low molecular weight|Heparin.low molecular weight
C1315159|T201|COMP|32685-0|LNC|Hepatitis B virus core Ab.IgG|Hepatitis B virus core Ab.IgG
C1315160|T201|COMP|32686-8|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1315161|T201|COMP|32687-6|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C1315162|T201|COMP|32688-4|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C1315163|T201|COMP|32689-2|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1315164|T201|COMP|32691-8|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1315165|T201|COMP|32692-6|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1315166|T201|COMP|32693-4|LNC|Lactate|Lactate
C1315167|T201|COMP|32694-2|LNC|Legionella longbeachae 1+2 Ab|Legionella longbeachae 1+2 Ab
C1315168|T201|COMP|32695-9|LNC|Legionella pneumophila atypical Ab|Legionella pneumophila atypical Ab
C1315169|T201|COMP|32696-7|LNC|Legionella pneumophila 1+2+3+4+5+6 Ab|Legionella pneumophila 1+2+3+4+5+6 Ab
C1315170|T201|COMP|32698-3|LNC|Magnesium.ionized|Magnesium.ionized
C1315173|T201|COMP|32701-5|LNC|Microsporidia identified|Microsporidia identified
C1315174|T201|COMP|32702-3|LNC|Muscle sarcolemma Ab|Muscle sarcolemma Ab
C1315175|T201|COMP|32703-1|LNC|Cytochrome b5 reductase|Cytochrome b5 reductase
C1315176|T201|COMP|32704-9|LNC|Neisseria gonorrhoeae Ab|Neisseria gonorrhoeae Ab
C1315177|T201|COMP|32705-6|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C1315178|T201|COMP|32706-4|LNC|Neisseria meningitidis serogroups A+C+w135+Y Ag|Neisseria meningitidis serogroups A+C+w135+Y Ag
C1315180|T201|COMP|32708-0|LNC|Neutrophil cytoplasmic Ab.classic|Neutrophil cytoplasmic Ab.classic
C1315181|T201|COMP|32710-6|LNC|Nitrite|Nitrite
C1315182|T201|COMP|32623-1|LNC|Platelet mean volume|Platelet mean volume
C1315183|T201|COMP|32712-2|LNC|Platelets.giant/100 leukocytes|Platelets.giant/100 leukocytes
C1315184|T201|COMP|32713-0|LNC|Potassium|Potassium
C1315185|T201|COMP|32714-8|LNC|Rickettsia typhus group Ab.IgM|Rickettsia typhus group Ab.IgM
C1315186|T201|COMP|32715-5|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C1315187|T201|COMP|32716-3|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C1315188|T201|COMP|32717-1|LNC|Sodium|Sodium
C1315189|T201|COMP|32718-9|LNC|Spermatozoa Ab.IgA|Spermatozoa Ab.IgA
C1315190|T201|COMP|32719-7|LNC|Spermatozoa Ab.IgG|Spermatozoa Ab.IgG
C1315191|T201|COMP|32720-5|LNC|Spermatozoa Ab.IgM|Spermatozoa Ab.IgM
C1315192|T201|COMP|32721-3|LNC|Tacrolimus|Tacrolimus
C1315193|T201|COMP|32722-1|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C1315194|T201|COMP|32723-9|LNC|Trichinella sp Ab.IgG|Trichinella sp Ab.IgG
C1315195|T201|COMP|32724-7|LNC|Trichomonas sp|Trichomonas sp
C1315196|T201|COMP|32725-4|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C1315197|T201|COMP|32726-2|LNC|Trypanosoma cruzi Ab.IgM|Trypanosoma cruzi Ab.IgM
C1315198|T201|COMP|32727-0|LNC|Urobilinogen|Urobilinogen
C1315199|T201|COMP|32728-8|LNC|Beta 1 globulin/Protein.total|Beta 1 globulin/Protein.total
C1315200|T201|COMP|32729-6|LNC|Beta 2 globulin/Protein.total|Beta 2 globulin/Protein.total
C1315201|T201|COMP|32730-4|LNC|Beta 1 globulin|Beta 1 globulin
C1315202|T201|COMP|32731-2|LNC|Beta 2 globulin|Beta 2 globulin
C1315203|T201|COMP|32732-0|LNC|Beta 1 globulin/Protein.total|Beta 1 globulin/Protein.total
C1315204|T201|COMP|32733-8|LNC|Beta 2 globulin/Protein.total|Beta 2 globulin/Protein.total
C1315205|T201|COMP|32734-6|LNC|Beta 1 globulin|Beta 1 globulin
C1315206|T201|COMP|32735-3|LNC|Beta 2 globulin|Beta 2 globulin
C1315207|T201|COMP|32736-1|LNC|Beta 1 globulin/Protein.total|Beta 1 globulin/Protein.total
C1315208|T201|COMP|32737-9|LNC|Beta 2 globulin/Protein.total|Beta 2 globulin/Protein.total
C1315209|T201|COMP|32738-7|LNC|Beta 1 globulin|Beta 1 globulin
C1315210|T201|COMP|32739-5|LNC|Beta 2 globulin|Beta 2 globulin
C1315211|T201|COMP|32740-3|LNC|Beta 1 globulin/Protein.total|Beta 1 globulin/Protein.total
C1315212|T201|COMP|32741-1|LNC|Beta 2 globulin/Protein.total|Beta 2 globulin/Protein.total
C1315213|T201|COMP|32742-9|LNC|Cells.CD117/100 cells|Cells.CD117/100 cells
C1315214|T201|COMP|32743-7|LNC|Cells.CD138/100 cells|Cells.CD138/100 cells
C1315215|T201|COMP|32744-5|LNC|Cells.CD55/100 cells|Cells.CD55/100 cells
C1315216|T201|COMP|32745-2|LNC|Cells.CD62E/100 cells|Cells.CD62E/100 cells
C1315217|T201|COMP|32746-0|LNC|Cells.CD62P/100 cells|Cells.CD62P/100 cells
C1315218|T201|COMP|32747-8|LNC|Cells.CD64/100 cells|Cells.CD64/100 cells
C1315219|T201|COMP|32748-6|LNC|Cells.CD90/100 cells|Cells.CD90/100 cells
C1315220|T201|COMP|32749-4|LNC|Cells.cyclin D1/100 cells|Cells.cyclin D1/100 cells
C1315222|T201|COMP|32751-0|LNC|Cells.HLA-DR+/100 cells|Cells.HLA-DR+/100 cells
C1315223|T201|COMP|32752-8|LNC|Cells.CD3/100 cells|Cells.CD3/100 cells
C1315224|T201|COMP|32753-6|LNC|Cells.CD4/100 cells|Cells.CD4/100 cells
C1315225|T201|COMP|32754-4|LNC|Cells.CD8/100 cells|Cells.CD8/100 cells
C1315226|T201|COMP|32755-1|LNC|Cells.CD19/100 cells|Cells.CD19/100 cells
C1315227|T201|COMP|32756-9|LNC|Cells.CD3+CD4+/Cells.CD3+CD8+|Cells.CD3+CD4+/Cells.CD3+CD8+
C1315228|T201|COMP|32757-7|LNC|Cells.BCL2/100 cells|Cells.BCL2/100 cells
C1315229|T201|COMP|32758-5|LNC|Cells.CD11b/100 cells|Cells.CD11b/100 cells
C1315230|T201|COMP|32759-3|LNC|Cells.myeloperoxidase/100 cells|Cells.myeloperoxidase/100 cells
C1315231|T201|COMP|32760-1|LNC|Cell type|Cell type
C1315232|T201|COMP|32761-9|LNC|Leukocytes|Leukocytes
C1315233|T201|COMP|32762-7|LNC|Epithelial cells|Epithelial cells
C1315234|T201|COMP|32763-5|LNC|Bacteria|Bacteria
C1315235|T201|COMP|32764-3|LNC|Clue cells|Clue cells
C1315236|T201|COMP|32765-0|LNC|Yeast|Yeast
C1315237|T201|COMP|32766-8|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C1315238|T201|COMP|32767-6|LNC|Borrelia burgdorferi 25kD Ab.IgM|Borrelia burgdorferi 25kD Ab.IgM
C1315239|T201|COMP|32768-4|LNC|Trichinella sp Ab.IgG|Trichinella sp Ab.IgG
C1315240|T201|COMP|32769-2|LNC|Alpha 1 antitrypsin phenotyping|Alpha 1 antitrypsin phenotyping
C1315241|T201|COMP|32770-0|LNC|Transfusion band number|Transfusion band number
C1315243|T201|COMP|32772-6|LNC|Cells.CD14|Cells.CD14
C1315244|T201|COMP|32773-4|LNC|Cells.CD24|Cells.CD24
C1315245|T201|COMP|32774-2|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1315246|T201|COMP|32775-9|LNC|Clostridium tetani toxoid Ab|Clostridium tetani toxoid Ab
C1315247|T201|COMP|32776-7|LNC|Erythrocytes|Erythrocytes
C1315248|T201|COMP|32777-5|LNC|Escherichia coli O157:H7 Ag|Escherichia coli O157:H7 Ag
C1315249|T201|COMP|32778-3|LNC|Fibrin strands|Fibrin strands
C1315250|T201|COMP|32779-1|LNC|Glucose-6-Phosphatase|Glucose-6-Phosphatase
C1315251|T201|COMP|32780-9|LNC|Histoplasma sp Ag|Histoplasma sp Ag
C1315252|T201|COMP|32781-7|LNC|Legionella sp Ag|Legionella sp Ag
C1315253|T201|COMP|32782-5|LNC|Leukocyte esterase+Nitrite|Leukocyte esterase+Nitrite
C1315254|T201|COMP|32783-3|LNC|Leucine+Isoleucine+Valine|Leucine+Isoleucine+Valine
C1315255|T201|COMP|32784-1|LNC|Mean peroxidase activity index|Mean peroxidase activity index
C1315257|T201|COMP|32786-6|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C1315258|T201|COMP|32787-4|LNC|Neutrophil cytoplasmic Ab.perinuclear|Neutrophil cytoplasmic Ab.perinuclear
C1315259|T201|COMP|32788-2|LNC|Polymorphonuclear cells/Monocytes|Polymorphonuclear cells/Monocytes
C1315260|T201|COMP|32789-0|LNC|Viscosity|Viscosity
C1315262|T201|COMP|32791-6|LNC|Cytomegalovirus Ab.IgG^1st specimen/2nd specimen|Cytomegalovirus Ab.IgG^1st specimen/2nd specimen
C1315263|T201|COMP|32792-4|LNC|Parvovirus B19 Ab.IgG^2nd specimen|Parvovirus B19 Ab.IgG^2nd specimen
C1315264|T201|COMP|32793-2|LNC|Parvovirus B19 Ab.IgG^1st specimen/2nd specimen|Parvovirus B19 Ab.IgG^1st specimen/2nd specimen
C1315265|T201|COMP|32794-0|LNC|Parvovirus B19 Ab.IgM^1st specimen|Parvovirus B19 Ab.IgM^1st specimen
C1315266|T201|COMP|32795-7|LNC|Parvovirus B19 Ab.IgM^2nd specimen|Parvovirus B19 Ab.IgM^2nd specimen
C1315267|T201|COMP|32796-5|LNC|Parvovirus B19 Ab.IgM^1st specimen/2nd specimen|Parvovirus B19 Ab.IgM^1st specimen/2nd specimen
C1315268|T201|COMP|32797-3|LNC|Drugs identified|Drugs identified
C1315270|T201|COMP|32799-9|LNC|Glycosaminoglycans/Creatinine|Glycosaminoglycans/Creatinine
C1315271|T201|COMP|32800-5|LNC|Neisseria meningitidis serogroups C+w135 Ag|Neisseria meningitidis serogroups C+w135 Ag
C1315272|T201|COMP|32801-3|LNC|Specimen volume|Specimen volume
C1315273|T201|COMP|32802-1|LNC|Color|Color
C1315274|T201|COMP|32803-9|LNC|Appearance|Appearance
C1315275|T201|COMP|32804-7|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C1315276|T201|COMP|32805-4|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C1315277|T201|COMP|32806-2|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1315278|T201|COMP|32807-0|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C1315279|T201|COMP|32808-8|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C1315280|T201|COMP|32809-6|LNC|Fungus identified|Fungus identified
C1315281|T201|COMP|32810-4|LNC|Bacteria identified|Bacteria identified
C1315284|T201|COMP|32813-8|LNC|Pathologist interpretation|Pathologist interpretation
C1315290|T201|COMP|32819-5|LNC|Microsporidia identified|Microsporidia identified
C1315291|T201|COMP|32820-3|LNC|Glucose^45M post dose lactose PO|Glucose^45M post dose lactose PO
C1315292|T201|COMP|32821-1|LNC|Interpretation|Interpretation
C1315293|T201|COMP|32822-9|LNC|Epithelial cells.squamous/100 cells|Epithelial cells.squamous/100 cells
C1315294|T201|COMP|32823-7|LNC|Columnar cells/100 cells|Columnar cells/100 cells
C1315296|T201|COMP|32825-2|LNC|Leukocytes|Leukocytes
C1315297|T201|COMP|32826-0|LNC|Parvovirus B19 Ab.IgG^1st specimen|Parvovirus B19 Ab.IgG^1st specimen
C1315298|T201|COMP|32827-8|LNC|HIV 1 p17+p18 Ab|HIV 1 p17+p18 Ab
C1315299|T201|COMP|32828-6|LNC|Epstein Barr virus capsid Ab.IgG^1st specimen|Epstein Barr virus capsid Ab.IgG^1st specimen
C1315300|T201|COMP|32829-4|LNC|Epstein Barr virus capsid Ab.IgG^2nd specimen|Epstein Barr virus capsid Ab.IgG^2nd specimen
C1315303|T201|COMP|32832-8|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C1315304|T201|COMP|32833-6|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1315306|T201|COMP|32835-1|LNC|Cytomegalovirus Ab.IgG^1st specimen/2nd specimen|Cytomegalovirus Ab.IgG^1st specimen/2nd specimen
C1315307|T201|COMP|32836-9|LNC|Parvovirus B19 Ab.IgG^1st specimen|Parvovirus B19 Ab.IgG^1st specimen
C1315308|T201|COMP|32837-7|LNC|Parvovirus B19 Ab.IgG^2nd specimen|Parvovirus B19 Ab.IgG^2nd specimen
C1315309|T201|COMP|32838-5|LNC|Parvovirus B19 Ab.IgG^1st specimen/2nd specimen|Parvovirus B19 Ab.IgG^1st specimen/2nd specimen
C1315310|T201|COMP|32839-3|LNC|Parvovirus B19 Ab.IgM^2nd specimen|Parvovirus B19 Ab.IgM^2nd specimen
C1315311|T201|COMP|32840-1|LNC|Parvovirus B19 Ab.IgM^1st specimen/2nd specimen|Parvovirus B19 Ab.IgM^1st specimen/2nd specimen
C1315312|T201|COMP|32841-9|LNC|Neisseria meningitidis serogroups C+w135 Ag|Neisseria meningitidis serogroups C+w135 Ag
C1315313|T201|COMP|32842-7|LNC|HIV 1 p17+p18 Ab|HIV 1 p17+p18 Ab
C1315314|T201|COMP|32843-5|LNC|Epstein Barr virus capsid Ab.IgG^1st specimen|Epstein Barr virus capsid Ab.IgG^1st specimen
C1315315|T201|COMP|32844-3|LNC|Epstein Barr virus capsid Ab.IgG^2nd specimen|Epstein Barr virus capsid Ab.IgG^2nd specimen
C1315318|T201|COMP|32847-6|LNC|Streptococcus pneumoniae 18 Ab.IgG|Streptococcus pneumoniae 18 Ab.IgG
C1315319|T201|COMP|32848-4|LNC|Neisseria meningitidis serogroups A+Y Ag|Neisseria meningitidis serogroups A+Y Ag
C1315320|T201|COMP|32849-2|LNC|Streptococcus pneumoniae 18 Ab.IgG|Streptococcus pneumoniae 18 Ab.IgG
C1315321|T201|COMP|32850-0|LNC|Streptococcus pneumoniae 5 Ab.IgG|Streptococcus pneumoniae 5 Ab.IgG
C1315322|T201|COMP|32851-8|LNC|Neisseria meningitidis serogroups A+Y Ag|Neisseria meningitidis serogroups A+Y Ag
C1315323|T201|COMP|32852-6|LNC|carBAMazepine.free/carBAMazepine.total|carBAMazepine.free/carBAMazepine.total
C1315324|T201|COMP|32853-4|LNC|Neuronal Ab|Neuronal Ab
C1315325|T201|COMP|32854-2|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C1315326|T201|COMP|32855-9|LNC|Cells.CD62/100 cells|Cells.CD62/100 cells
C1315327|T201|COMP|32856-7|LNC|Cells.cytoplasmic CD22/100 cells|Cells.cytoplasmic CD22/100 cells
C1315328|T201|COMP|32857-5|LNC|Cells.cytoplasmic CD3/100 cells|Cells.cytoplasmic CD3/100 cells
C1315329|T201|COMP|32858-3|LNC|Cells.IgG/100 cells|Cells.IgG/100 cells
C1315330|T201|COMP|32859-1|LNC|Cells.multiple drug resistance/100 cells|Cells.multiple drug resistance/100 cells
C1315331|T201|COMP|32860-9|LNC|Cells.TCR alpha beta/100 cells|Cells.TCR alpha beta/100 cells
C1315332|T201|COMP|32861-7|LNC|Cells.TCR gamma delta/100 cells|Cells.TCR gamma delta/100 cells
C1315333|T201|COMP|32862-5|LNC|Osmotic fragility^incubated|Osmotic fragility^incubated
C1315334|T201|COMP|32863-3|LNC|Osmotic fragility^fresh|Osmotic fragility^fresh
C1315466|T201|COMP|32995-3|LNC|Lutropin^20M post XXX challenge|Lutropin^20M post XXX challenge
C1315467|T201|COMP|32996-1|LNC|HER2|HER2
C1315468|T201|COMP|32997-9|LNC|cycloSPORINE^2H post dose|cycloSPORINE^2H post dose
C1315469|T201|COMP|32998-7|LNC|Tissue transglutaminase Ab.IgG|Tissue transglutaminase Ab.IgG
C1315470|T201|COMP|32999-5|LNC|Rickettsia spotted fever group Ab.IgG|Rickettsia spotted fever group Ab.IgG
C1315471|T201|COMP|33000-1|LNC|Rickettsia spotted fever group Ab.IgM|Rickettsia spotted fever group Ab.IgM
C1315472|T201|COMP|33001-9|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C1315473|T201|COMP|33002-7|LNC|Triticum spelta Ab.IgE|Triticum spelta Ab.IgE
C1315474|T201|COMP|33003-5|LNC|Triticum spelta Ab.IgE.RAST class|Triticum spelta Ab.IgE.RAST class
C1315475|T201|COMP|33004-3|LNC|Kelp Ab.IgE|Kelp Ab.IgE
C1315476|T201|COMP|33005-0|LNC|Kelp Ab.IgE.RAST class|Kelp Ab.IgE.RAST class
C1315477|T201|COMP|33006-8|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1315478|T201|COMP|33007-6|LNC|Protoporphyrin.zinc|Protoporphyrin.zinc
C1315479|T201|COMP|33008-4|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C1315480|T201|COMP|33009-2|LNC|Chylomicrons|Chylomicrons
C1315481|T201|COMP|33010-0|LNC|Cheese colby Ab.IgE|Cheese colby Ab.IgE
C1315482|T201|COMP|33011-8|LNC|Cheese colby Ab.IgE.RAST class|Cheese colby Ab.IgE.RAST class
C1315483|T201|COMP|33012-6|LNC|Cheese provolone Ab.IgE|Cheese provolone Ab.IgE
C1315484|T201|COMP|33013-4|LNC|Cheese provolone Ab.IgE.RAST class|Cheese provolone Ab.IgE.RAST class
C1315485|T201|COMP|33014-2|LNC|Cheese romano Ab.IgE|Cheese romano Ab.IgE
C1315486|T201|COMP|33015-9|LNC|Cheese romano Ab.IgE.RAST class|Cheese romano Ab.IgE.RAST class
C1315487|T201|COMP|33016-7|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C1315488|T201|COMP|33017-5|LNC|Parasites|Parasites
C1315489|T201|COMP|33018-3|LNC|Protein.monoclonal|Protein.monoclonal
C1315490|T201|COMP|33019-1|LNC|Pseudocasts|Pseudocasts
C1315491|T201|COMP|33020-9|LNC|Triple phosphate crystals|Triple phosphate crystals
C1315492|T201|COMP|33021-7|LNC|Tyrosine crystals|Tyrosine crystals
C1315494|T201|COMP|33023-3|LNC|Cells.CD34/100 cells|Cells.CD34/100 cells
C1315495|T201|COMP|33024-1|LNC|Glucose^30M post 1.2 g/kg lactose PO|Glucose^30M post 1.2 g/kg lactose PO
C1315496|T201|COMP|33025-8|LNC|Hemoglobin|Hemoglobin
C1315497|T201|COMP|33026-6|LNC|Hemoglobin|Hemoglobin
C1315498|T201|COMP|33027-4|LNC|Herpes simplex virus+Varicella zoster virus DNA|Herpes simplex virus+Varicella zoster virus DNA
C1315499|T201|COMP|33028-2|LNC|Leukocytes|Leukocytes
C1315500|T201|COMP|33029-0|LNC|Cells.CD3+TCR/100 cells|Cells.CD3+TCR/100 cells
C1315501|T201|COMP|33030-8|LNC|Cells.CD34|Cells.CD34
C1315502|T201|COMP|33031-6|LNC|Sodium urate crystals|Sodium urate crystals
C1315503|T201|COMP|33032-4|LNC|Spermatozoa.progressive|Spermatozoa.progressive
C1315504|T201|COMP|33033-2|LNC|CD45 positive events|CD45 positive events
C1315505|T201|COMP|33034-0|LNC|CD45 negative events|CD45 negative events
C1315506|T201|COMP|33035-7|LNC|Reason for lab test|Reason for lab test
C1315507|T201|COMP|33036-5|LNC|Fatty acids.very long chain.C26:1|Fatty acids.very long chain.C26:1
C1315508|T201|COMP|33037-3|LNC|Anion gap|Anion gap
C1315509|T201|COMP|33038-1|LNC|Candida sp identified|Candida sp identified
C1315510|T201|COMP|33039-9|LNC|Fungus identified|Fungus identified
C1315511|T201|COMP|33040-7|LNC|Hypnotics|Hypnotics
C1315512|T201|COMP|33041-5|LNC|Hypnotics|Hypnotics
C1315513|T201|COMP|33042-3|LNC|Interpretation|Interpretation
C1315514|T201|COMP|33043-1|LNC|Ketones|Ketones
C1315515|T201|COMP|33044-9|LNC|Pyknosis|Pyknosis
C1315516|T201|COMP|33045-6|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C1315517|T201|COMP|33046-4|LNC|Tranquilizers|Tranquilizers
C1315518|T201|COMP|33047-2|LNC|Tranquilizers|Tranquilizers
C1315519|T201|COMP|33048-0|LNC|Eosin-5-Maleimide binding|Eosin-5-Maleimide binding
C1315520|T201|COMP|33049-8|LNC|Hypertonic cryohemolysis|Hypertonic cryohemolysis
C1315521|T201|COMP|33050-6|LNC|Pseudocholinesterase phenotype|Pseudocholinesterase phenotype
C1315522|T201|COMP|33051-4|LNC|Erythrocytes|Erythrocytes
C1315523|T201|COMP|33052-2|LNC|Leukocytes|Leukocytes
C1315524|T201|COMP|33053-0|LNC|Protoporphyrin|Protoporphyrin
C1315525|T201|COMP|33054-8|LNC|BCL2 Ag|BCL2 Ag
C1315526|T201|COMP|33055-5|LNC|Ki-67 nuclear Ag|Ki-67 nuclear Ag
C1315527|T201|COMP|33056-3|LNC|Sezary cells|Sezary cells
C1315528|T201|COMP|33057-1|LNC|Heinz bodies/100 erythrocytes|Heinz bodies/100 erythrocytes
C1315529|T201|COMP|33058-9|LNC|Ketones|Ketones
C1315530|T201|COMP|33059-7|LNC|Fluorescence polarization|Fluorescence polarization
C1315531|T201|COMP|33060-5|LNC|chlordiazePOXIDE+Metabolites|chlordiazePOXIDE+Metabolites
C1315532|T201|COMP|33061-3|LNC|Homocystine^6H post dose methionine - post CFst|Homocystine^6H post dose methionine - post CFst
C1315533|T201|COMP|33062-1|LNC|Blood group antigens tested for|Blood group antigens tested for
C1315534|T201|COMP|33063-9|LNC|Alkaline phosphatase isoenzymes|Alkaline phosphatase isoenzymes
C1315535|T201|COMP|33064-7|LNC|Chromate|Chromate
C1315664|T201|COMP|33193-4|LNC|Viable cells/100 cells|Viable cells/100 cells
C1315665|T201|COMP|33194-2|LNC|Viable cells/100 cells|Viable cells/100 cells
C1315666|T201|COMP|33195-9|LNC|Viable cells/100 cells|Viable cells/100 cells
C1315671|T201|COMP|33200-7|LNC|Amyloid beta 42 peptide|Amyloid beta 42 peptide
C1315672|T201|COMP|33201-5|LNC|Cells.CD11c/100 cells|Cells.CD11c/100 cells
C1315673|T201|COMP|33202-3|LNC|Cells.CD11c/100 cells|Cells.CD11c/100 cells
C1315674|T201|COMP|33203-1|LNC|Amyloid beta 42 peptide|Amyloid beta 42 peptide
C1315675|T201|COMP|33204-9|LNC|Troponin T.cardiac|Troponin T.cardiac
C1315676|T201|COMP|33205-6|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C1315677|T201|COMP|33206-4|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C1315678|T201|COMP|33207-2|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C1315679|T201|COMP|33208-0|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C1315680|T201|COMP|33209-8|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C1315681|T201|COMP|33210-6|LNC|Transferrin receptor.soluble|Transferrin receptor.soluble
C1315682|T201|COMP|33211-4|LNC|Interleukin 8|Interleukin 8
C1315683|T201|COMP|33212-2|LNC|N-acetyl-L-aspartate|N-acetyl-L-aspartate
C1315684|T201|COMP|33213-0|LNC|Glycine plas/Glycine CSF|Glycine plas/Glycine CSF
C1315685|T201|COMP|33214-8|LNC|Taurine|Taurine
C1315686|T201|COMP|33215-5|LNC|Neutrophils.agranular|Neutrophils.agranular
C1315687|T201|COMP|33216-3|LNC|Platelets.agranular|Platelets.agranular
C1315688|T201|COMP|33217-1|LNC|Spermatozoa.agglutinated|Spermatozoa.agglutinated
C1315689|T201|COMP|33218-9|LNC|Bacteria|Bacteria
C1315690|T201|COMP|33219-7|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C1315691|T201|COMP|33220-5|LNC|Transitional cells|Transitional cells
C1315692|T201|COMP|33221-3|LNC|Epithelial cells.renal|Epithelial cells.renal
C1315693|T201|COMP|33222-1|LNC|Oval fat bodies (globules)|Oval fat bodies (globules)
C1315694|T201|COMP|33223-9|LNC|Hyaline casts|Hyaline casts
C1315695|T201|COMP|33224-7|LNC|Granular casts.fine|Granular casts.fine
C1315696|T201|COMP|33225-4|LNC|Granular casts.fine|Granular casts.fine
C1315697|T201|COMP|33226-2|LNC|Granular casts.coarse|Granular casts.coarse
C1315698|T201|COMP|33227-0|LNC|Granular casts.coarse|Granular casts.coarse
C1315699|T201|COMP|33228-8|LNC|Leukocyte casts|Leukocyte casts
C1315700|T201|COMP|33229-6|LNC|Erythrocyte casts|Erythrocyte casts
C1315701|T201|COMP|33230-4|LNC|Waxy casts|Waxy casts
C1315702|T201|COMP|33231-2|LNC|Fatty casts|Fatty casts
C1315703|T201|COMP|33232-0|LNC|Spermatozoa|Spermatozoa
C1315704|T201|COMP|33233-8|LNC|Urate crystals|Urate crystals
C1315705|T201|COMP|33234-6|LNC|Calcium oxalate crystals|Calcium oxalate crystals
C1315706|T201|COMP|33235-3|LNC|Calcium phosphate crystals|Calcium phosphate crystals
C1315707|T201|COMP|33236-1|LNC|Bilirubin crystals|Bilirubin crystals
C1315708|T201|COMP|33237-9|LNC|Sulfonamide crystals|Sulfonamide crystals
C1315709|T201|COMP|33238-7|LNC|Triple phosphate crystals|Triple phosphate crystals
C1315710|T201|COMP|33239-5|LNC|Ammonium urate crystals|Ammonium urate crystals
C1315711|T201|COMP|33240-3|LNC|Cystine crystals|Cystine crystals
C1315712|T201|COMP|33241-1|LNC|Calcium carbonate crystals|Calcium carbonate crystals
C1315713|T201|COMP|33242-9|LNC|Fungi.filamentous|Fungi.filamentous
C1315714|T201|COMP|33243-7|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C1315715|T201|COMP|33244-5|LNC|Guanidinoacetate|Guanidinoacetate
C1315716|T201|COMP|33245-2|LNC|Amylase|Amylase
C1315717|T201|COMP|33246-0|LNC|Ovary Ab|Ovary Ab
C1315718|T201|COMP|33247-8|LNC|Specimen weight|Specimen weight
C1315719|T201|COMP|33248-6|LNC|Diabetes status|Diabetes status
C1315720|T201|COMP|33249-4|LNC|Hyperchromia|Hyperchromia
C1315721|T201|COMP|33250-2|LNC|Cells.CD55|Cells.CD55
C1315722|T201|COMP|33253-6|LNC|Nuclear Ab|Nuclear Ab
C1315723|T201|COMP|33254-4|LNC|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1315724|T201|COMP|33255-1|LNC|Cell fractions|Cell fractions
C1315725|T201|COMP|33256-9|LNC|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C1315726|T201|COMP|33257-7|LNC|Cortisol|Cortisol
C1315727|T201|COMP|33258-5|LNC|Thyrotropin^30M post dose TRH|Thyrotropin^30M post dose TRH
C1315728|T201|COMP|33259-3|LNC|Thyrotropin^1H post dose TRH|Thyrotropin^1H post dose TRH
C1315729|T201|COMP|33260-1|LNC|Thyrotropin^1.5H post dose TRH|Thyrotropin^1.5H post dose TRH
C1315730|T201|COMP|33261-9|LNC|Thyrotropin^2H post dose TRH|Thyrotropin^2H post dose TRH
C1315731|T201|COMP|33262-7|LNC|Metamyelocytes/100 leukocytes|Metamyelocytes/100 leukocytes
C1315732|T201|COMP|33263-5|LNC|Metamyelocytes/100 leukocytes|Metamyelocytes/100 leukocytes
C1315733|T201|COMP|33264-3|LNC|Osmol gap|Osmol gap
C1315734|T201|COMP|33265-0|LNC|Toxoplasma gondii Ab.IgA|Toxoplasma gondii Ab.IgA
C1315735|T201|COMP|33266-8|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C1315736|T201|COMP|33267-6|LNC|Aspergillus sp Ab.IgG|Aspergillus sp Ab.IgG
C1315737|T201|COMP|33268-4|LNC|Bordetella pertussis.pertussis toxin Ab.IgG|Bordetella pertussis.pertussis toxin Ab.IgG
C1315738|T201|COMP|33269-2|LNC|Thyrotropin^pre dose TRH|Thyrotropin^pre dose TRH
C1315741|T201|COMP|33272-6|LNC|Cryoglobulin|Cryoglobulin
C1315742|T201|COMP|33273-4|LNC|3-Methylglutaconate|3-Methylglutaconate
C1315743|T201|COMP|33274-2|LNC|5-Methyltetrahydrofolate|5-Methyltetrahydrofolate
C1315744|T201|COMP|33275-9|LNC|7-Dehydrocholesterol|7-Dehydrocholesterol
C1315745|T201|COMP|33276-7|LNC|Aureobasidium pullulans Ab.IgG.RAST class|Aureobasidium pullulans Ab.IgG.RAST class
C1315746|T201|COMP|33277-5|LNC|Acetaminophen+Phenacetin|Acetaminophen+Phenacetin
C1315747|T201|COMP|33278-3|LNC|Acetylcholine receptor blocking Ab|Acetylcholine receptor blocking Ab
C1315748|T201|COMP|33279-1|LNC|Acetylcholine receptor modulation Ab|Acetylcholine receptor modulation Ab
C1315749|T201|COMP|33280-9|LNC|Amphetamine+Methamphetamine|Amphetamine+Methamphetamine
C1315750|T201|COMP|33281-7|LNC|Curvularia specifera Ab.IgG.RAST class|Curvularia specifera Ab.IgG.RAST class
C1315751|T201|COMP|33282-5|LNC|Cannabinoids|Cannabinoids
C1315752|T201|COMP|33283-3|LNC|Ictalurus punctatus Ab.IgG.RAST class|Ictalurus punctatus Ab.IgG.RAST class
C1315753|T201|COMP|32376-6|LNC|Clinafloxacin|Clinafloxacin
C1315754|T201|COMP|33285-8|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C1315755|T201|COMP|33286-6|LNC|Fusarium moniliforme Ab.IgG.RAST class|Fusarium moniliforme Ab.IgG.RAST class
C1315756|T201|COMP|33287-4|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C1315757|T201|COMP|33288-2|LNC|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C1315758|T201|COMP|33289-0|LNC|Helminthosporium sp Ab.IgG.RAST class|Helminthosporium sp Ab.IgG.RAST class
C1315759|T201|COMP|33290-8|LNC|Histamine|Histamine
C1315760|T201|COMP|33291-6|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C1315761|T201|COMP|33292-4|LNC|Herpes simplex virus 1+2 Ab|Herpes simplex virus 1+2 Ab
C1315762|T201|COMP|33293-2|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C1315763|T201|COMP|33294-0|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1315764|T201|COMP|33295-7|LNC|JC virus DNA|JC virus DNA
C1315765|T201|COMP|33296-5|LNC|Actinidia chinensis Ab.IgG.RAST class|Actinidia chinensis Ab.IgG.RAST class
C1315766|T201|COMP|33297-3|LNC|Mucor racemosus Ab.IgG.RAST class|Mucor racemosus Ab.IgG.RAST class
C1315767|T201|COMP|18859-9|LNC|Amdinocillin|Amdinocillin
C1315768|T201|COMP|33299-9|LNC|N-acetyl-L-aspartate|N-acetyl-L-aspartate
C1315769|T201|COMP|33300-5|LNC|Naproxen|Naproxen
C1315770|T201|COMP|33301-3|LNC|Norchlordiazepoxide|Norchlordiazepoxide
C1315771|T201|COMP|33302-1|LNC|Phthalic anhydride Ab.IgG.RAST class|Phthalic anhydride Ab.IgG.RAST class
C1315772|T201|COMP|33303-9|LNC|Phoma betae Ab.IgG.RAST class|Phoma betae Ab.IgG.RAST class
C1315773|T201|COMP|33304-7|LNC|Penicillium notatum Ab.IgG.RAST class|Penicillium notatum Ab.IgG.RAST class
C1315774|T201|COMP|33305-4|LNC|Perca spp Ab.IgG.RAST class|Perca spp Ab.IgG.RAST class
C1315775|T201|COMP|33306-2|LNC|Phosphatidate Ab|Phosphatidate Ab
C1315776|T201|COMP|33307-0|LNC|Phosphatidylcholine Ab|Phosphatidylcholine Ab
C1315777|T201|COMP|33308-8|LNC|Phosphatidylethanolamine Ab|Phosphatidylethanolamine Ab
C1315778|T201|COMP|33309-6|LNC|Phosphatidylinositol Ab|Phosphatidylinositol Ab
C1315779|T201|COMP|33310-4|LNC|Phosphatidylserine Ab|Phosphatidylserine Ab
C1315780|T201|COMP|33311-2|LNC|Porphyrins|Porphyrins
C1315781|T201|COMP|33312-0|LNC|Rhizopus nigricans Ab.IgG.RAST class|Rhizopus nigricans Ab.IgG.RAST class
C1315782|T201|COMP|33313-8|LNC|Rheumatoid factor.IgA|Rheumatoid factor.IgA
C1315783|T201|COMP|33314-6|LNC|Rheumatoid factor.IgG|Rheumatoid factor.IgG
C1315784|T201|COMP|33315-3|LNC|Stemphylium botryosum Ab.IgG.RAST class|Stemphylium botryosum Ab.IgG.RAST class
C1315785|T201|COMP|33316-1|LNC|Salmonella paratyphi A O Ab|Salmonella paratyphi A O Ab
C1315786|T201|COMP|33317-9|LNC|Schistosoma sp Ab.IgG|Schistosoma sp Ab.IgG
C1315787|T201|COMP|33318-7|LNC|Spermatozoa Ab.IgM|Spermatozoa Ab.IgM
C1315788|T201|COMP|33319-5|LNC|Toxoplasma gondii Ab.IgE|Toxoplasma gondii Ab.IgE
C1315789|T201|COMP|33320-3|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C1315790|T201|COMP|33321-1|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C1315791|T201|COMP|33322-9|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1315792|T201|COMP|33323-7|LNC|Theophylline|Theophylline
C1315793|T201|COMP|33324-5|LNC|Trichophyton Ab.IgG.RAST class|Trichophyton Ab.IgG.RAST class
C1315794|T201|COMP|33325-2|LNC|Trypsin|Trypsin
C1315795|T201|COMP|33326-0|LNC|Turbidity|Turbidity
C1315796|T201|COMP|33327-8|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C1315797|T201|COMP|33328-6|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C1315798|T201|COMP|33329-4|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C1315799|T201|COMP|33330-2|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1315800|T201|COMP|33331-0|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1315801|T201|COMP|33332-8|LNC|Linezolid|Linezolid
C1315802|T201|COMP|33333-6|LNC|Colistin|Colistin
C1315803|T201|COMP|33334-4|LNC|Quinupristin+Dalfopristin|Quinupristin+Dalfopristin
C1315804|T201|COMP|33335-1|LNC|Diphenylmethoxyacetate|Diphenylmethoxyacetate
C1315805|T201|COMP|33336-9|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C1315806|T201|COMP|33337-7|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C1315807|T201|COMP|33338-5|LNC|Zolpidem|Zolpidem
C1315808|T201|COMP|33339-3|LNC|Zolpidem|Zolpidem
C1315809|T201|COMP|33340-1|LNC|Zolpidem|Zolpidem
C1315810|T201|COMP|33341-9|LNC|Granular casts|Granular casts
C1315811|T201|COMP|33342-7|LNC|Epithelial cells|Epithelial cells
C1315812|T201|COMP|33343-5|LNC|Leukotriene E4/Creatinine|Leukotriene E4/Creatinine
C1315813|T201|COMP|33344-3|LNC|Leukotriene E4|Leukotriene E4
C1315814|T201|COMP|33345-0|LNC|Histrelin|Histrelin
C1315815|T201|COMP|33346-8|LNC|Cortisol.free|Cortisol.free
C1315816|T201|COMP|33347-6|LNC|17-Ketosteroids/Creatinine|17-Ketosteroids/Creatinine
C1315817|T201|COMP|33348-4|LNC|Pemoline|Pemoline
C1315818|T201|COMP|33349-2|LNC|Pemoline|Pemoline
C1315819|T201|COMP|33350-0|LNC|Lysergate diethylamide|Lysergate diethylamide
C1315820|T201|COMP|33351-8|LNC|11-Dehydro thromboxane beta 2|11-Dehydro thromboxane beta 2
C1315821|T201|COMP|33352-6|LNC|Glucose/Creatinine|Glucose/Creatinine
C1315822|T201|COMP|33353-4|LNC|Alanine aminopeptidase|Alanine aminopeptidase
C1315823|T201|COMP|33354-2|LNC|N-acetyl-beta-glucosaminidase|N-acetyl-beta-glucosaminidase
C1315824|T201|COMP|33355-9|LNC|Urea nitrogen|Urea nitrogen
C1315827|T201|COMP|33358-3|LNC|Protein.monoclonal|Protein.monoclonal
C1315828|T201|COMP|33359-1|LNC|Branched chain keto-acid dehydrogenase complex|Branched chain keto-acid dehydrogenase complex
C1315829|T201|COMP|33360-9|LNC|Galactose 1 phosphate|Galactose 1 phosphate
C1315830|T201|COMP|33361-7|LNC|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C1315831|T201|COMP|33362-5|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C1315832|T201|COMP|33363-3|LNC|Normocytic|Normocytic
C1315833|T201|COMP|33364-1|LNC|Normochromic|Normochromic
C1315834|T201|COMP|33365-8|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C1315835|T201|COMP|33366-6|LNC|Chloride|Chloride
C1315836|T201|COMP|33367-4|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C1315837|T201|COMP|33368-2|LNC|Amylase|Amylase
C1315838|T201|COMP|33369-0|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C1315839|T201|COMP|33370-8|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C1315840|T201|COMP|33371-6|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C1315841|T201|COMP|33372-4|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C1315842|T201|COMP|33373-2|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C1315843|T201|COMP|33374-0|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C1315844|T201|COMP|33375-7|LNC|Chylomicrons|Chylomicrons
C1315845|T201|COMP|33376-5|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C1315846|T201|COMP|33377-3|LNC|Blastomyces sp Ab|Blastomyces sp Ab
C1315847|T201|COMP|33378-1|LNC|Blastomyces sp Ab|Blastomyces sp Ab
C1315848|T201|COMP|33379-9|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1315849|T201|COMP|33380-7|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1315850|T201|COMP|33381-5|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1315851|T201|COMP|33382-3|LNC|Respiratory syncytial virus Ab|Respiratory syncytial virus Ab
C1315852|T201|COMP|33383-1|LNC|Influenza virus A Bangkok Ab|Influenza virus A Bangkok Ab
C1315853|T201|COMP|33384-9|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C1315854|T201|COMP|33385-6|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C1315855|T201|COMP|33386-4|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C1315856|T201|COMP|33387-2|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C1315857|T201|COMP|33388-0|LNC|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C1315858|T201|COMP|33389-8|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C1315859|T201|COMP|33390-6|LNC|Respiratory syncytial virus Ab|Respiratory syncytial virus Ab
C1315860|T201|COMP|33391-4|LNC|Coxsackievirus A8 Ab|Coxsackievirus A8 Ab
C1315861|T201|COMP|33392-2|LNC|Coxsackievirus A8 Ab|Coxsackievirus A8 Ab
C1315862|T201|COMP|33393-0|LNC|Granular casts.coarse|Granular casts.coarse
C1315863|T201|COMP|33394-8|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C1315864|T201|COMP|33395-5|LNC|Epstein Barr virus capsid Ab|Epstein Barr virus capsid Ab
C1315865|T201|COMP|33396-3|LNC|Neisseria meningitidis serogroups A+C+w135+Y Ag|Neisseria meningitidis serogroups A+C+w135+Y Ag
C1315866|T201|COMP|33397-1|LNC|Neisseria meningitidis serogroups A+C+w135+Y Ag|Neisseria meningitidis serogroups A+C+w135+Y Ag
C1315867|T201|COMP|33398-9|LNC|Neisseria meningitidis serogroups A+C+w135+Y Ag|Neisseria meningitidis serogroups A+C+w135+Y Ag
C1315871|T201|COMP|33402-9|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1315872|T201|COMP|33403-7|LNC|Fatty acids.very long chain.C26:0|Fatty acids.very long chain.C26:0
C1315874|T201|COMP|33405-2|LNC|Glucose|Glucose
C1315875|T201|COMP|33406-0|LNC|Candida albicans Ab|Candida albicans Ab
C1315876|T201|COMP|33407-8|LNC|Protein|Protein
C1315877|T201|COMP|33408-6|LNC|Complement C2|Complement C2
C1315878|T201|COMP|33409-4|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C1315879|T201|COMP|33410-2|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C1315880|T201|COMP|33411-0|LNC|Hemoglobin.free|Hemoglobin.free
C1315881|T201|COMP|33412-8|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C1315882|T201|COMP|33413-6|LNC|Lipoprotein.beta/Lipoprotein.total|Lipoprotein.beta/Lipoprotein.total
C1315883|T201|COMP|33414-4|LNC|Lipoprotein.pre-beta/Lipoprotein.total|Lipoprotein.pre-beta/Lipoprotein.total
C1315884|T201|COMP|33415-1|LNC|IgG|IgG
C1315885|T201|COMP|33416-9|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1315887|T201|COMP|33418-5|LNC|Neuronal Ab.IgG|Neuronal Ab.IgG
C1315888|T201|COMP|33419-3|LNC|Histoplasma sp Ag|Histoplasma sp Ag
C1315889|T201|COMP|33420-1|LNC|Histoplasma sp Ag|Histoplasma sp Ag
C1315890|T201|COMP|33421-9|LNC|Alkaline phosphatase.other fractions|Alkaline phosphatase.other fractions
C1315891|T201|COMP|33422-7|LNC|Amphiphysin Ab|Amphiphysin Ab
C1315892|T201|COMP|33423-5|LNC|Amphiphysin Ab|Amphiphysin Ab
C1315924|T201|COMP|33455-7|LNC|Appearance|Appearance
C1315927|T201|COMP|33458-1|LNC|Bilirubin.glucuronidated|Bilirubin.glucuronidated
C1315928|T201|COMP|33459-9|LNC|Toxoplasma gondii Ab.IgA|Toxoplasma gondii Ab.IgA
C1315930|T201|COMP|33461-5|LNC|Candida albicans Ab|Candida albicans Ab
C1315931|T201|COMP|33462-3|LNC|Hepatitis C virus Ab.IgG|Hepatitis C virus Ab.IgG
C1315932|T201|COMP|33463-1|LNC|Hepatitis B virus little e Ab.IgG|Hepatitis B virus little e Ab.IgG
C1315933|T201|COMP|33464-9|LNC|Hepatitis D virus Ag|Hepatitis D virus Ag
C1315934|T201|COMP|33465-6|LNC|Francisella tularensis Ab.IgG|Francisella tularensis Ab.IgG
C1315935|T201|COMP|33466-4|LNC|Francisella tularensis Ab.IgM|Francisella tularensis Ab.IgM
C1315936|T201|COMP|33467-2|LNC|Prealbumin|Prealbumin
C1315937|T201|COMP|33468-0|LNC|West Nile virus Ab|West Nile virus Ab
C1315938|T201|COMP|33469-8|LNC|Clostridium tetani Ab.IgG|Clostridium tetani Ab.IgG
C1315939|T201|COMP|33470-6|LNC|Salmonella paratyphi A O Ab|Salmonella paratyphi A O Ab
C1315940|T201|COMP|33471-4|LNC|Hydrogen/Expired gas^post XXX challenge|Hydrogen/Expired gas^post XXX challenge
C1315941|T201|COMP|33472-2|LNC|Acylcarnitine pattern|Acylcarnitine pattern
C1315942|T201|COMP|33473-0|LNC|Bile acid pattern|Bile acid pattern
C1315943|T201|COMP|33474-8|LNC|Glycosaminoglycans pattern|Glycosaminoglycans pattern
C1315944|T201|COMP|33475-5|LNC|Organic acids pattern|Organic acids pattern
C1315945|T201|COMP|33476-3|LNC|Organic acids pattern|Organic acids pattern
C1315946|T201|COMP|33477-1|LNC|Organic acids pattern|Organic acids pattern
C1315947|T201|COMP|33478-9|LNC|Fatty acids.very long chain pattern|Fatty acids.very long chain pattern
C1315948|T201|COMP|33479-7|LNC|Epstein Barr virus early restricted Ab|Epstein Barr virus early restricted Ab
C1315949|T201|COMP|33480-5|LNC|Methane/Expired gas^2H post dose lactose PO|Methane/Expired gas^2H post dose lactose PO
C1315950|T201|COMP|33481-3|LNC|Methane/Expired gas^2.5H post dose lactose PO|Methane/Expired gas^2.5H post dose lactose PO
C1315951|T201|COMP|33482-1|LNC|Methane/Expired gas^3H post dose lactose PO|Methane/Expired gas^3H post dose lactose PO
C1315952|T201|COMP|33483-9|LNC|Patient symptoms^pre dose lactose PO|Patient symptoms^pre dose lactose PO
C1315953|T201|COMP|33484-7|LNC|Patient symptoms^30M post dose lactose PO|Patient symptoms^30M post dose lactose PO
C1315954|T201|COMP|33485-4|LNC|Patient symptoms^1H post dose lactose PO|Patient symptoms^1H post dose lactose PO
C1315955|T201|COMP|33486-2|LNC|Patient symptoms^1.5H post dose lactose PO|Patient symptoms^1.5H post dose lactose PO
C1315956|T201|COMP|33487-0|LNC|Patient symptoms^2H post dose lactose PO|Patient symptoms^2H post dose lactose PO
C1315957|T201|COMP|33488-8|LNC|Patient symptoms^2.5H post dose lactose PO|Patient symptoms^2.5H post dose lactose PO
C1315959|T201|COMP|33490-4|LNC|Hydrogen/Expired gas^pre dose lactose PO|Hydrogen/Expired gas^pre dose lactose PO
C1315960|T201|COMP|33491-2|LNC|Hydrogen/Expired gas^30M post dose lactose PO|Hydrogen/Expired gas^30M post dose lactose PO
C1315961|T201|COMP|33492-0|LNC|Hydrogen/Expired gas^1H post dose lactose PO|Hydrogen/Expired gas^1H post dose lactose PO
C1315962|T201|COMP|33493-8|LNC|Hydrogen/Expired gas^1.5H post dose lactose PO|Hydrogen/Expired gas^1.5H post dose lactose PO
C1315963|T201|COMP|33494-6|LNC|Hydrogen/Expired gas^2H post dose lactose PO|Hydrogen/Expired gas^2H post dose lactose PO
C1315964|T201|COMP|33495-3|LNC|Hydrogen/Expired gas^2.5H post dose lactose PO|Hydrogen/Expired gas^2.5H post dose lactose PO
C1315965|T201|COMP|33496-1|LNC|Hydrogen/Expired gas^3H post dose lactose PO|Hydrogen/Expired gas^3H post dose lactose PO
C1315966|T201|COMP|33497-9|LNC|Methane/Expired gas^pre dose lactose PO|Methane/Expired gas^pre dose lactose PO
C1315967|T201|COMP|33498-7|LNC|Methane/Expired gas^30M post dose lactose PO|Methane/Expired gas^30M post dose lactose PO
C1315968|T201|COMP|33499-5|LNC|Methane/Expired gas^1H post dose lactose PO|Methane/Expired gas^1H post dose lactose PO
C1315969|T201|COMP|33500-0|LNC|Methane/Expired gas^1.5H post dose lactose PO|Methane/Expired gas^1.5H post dose lactose PO
C1315973|T201|COMP|33504-2|LNC|Hydrogen+Methane/Expired gas^pre dose lactose PO|Hydrogen+Methane/Expired gas^pre dose lactose PO
C1315976|T201|COMP|33507-5|LNC|Alpha-Phenyl-2-Piperidine acetate|Alpha-Phenyl-2-Piperidine acetate
C1315977|T201|COMP|33508-3|LNC|HIV 1 p65+p66 Ab|HIV 1 p65+p66 Ab
C1315978|T201|COMP|33509-1|LNC|Hemoglobin|Hemoglobin
C1315979|T201|COMP|33510-9|LNC|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C1315980|T201|COMP|33511-7|LNC|Appearance|Appearance
C1315981|T201|COMP|33512-5|LNC|Color|Color
C1315982|T201|COMP|33513-3|LNC|Specific gravity|Specific gravity
C1315983|T201|COMP|33514-1|LNC|Specimen volume|Specimen volume
C1315984|T201|COMP|33515-8|LNC|Clarity|Clarity
C1315985|T201|COMP|33516-6|LNC|Reticulocytes.immature/Reticulocytes.total|Reticulocytes.immature/Reticulocytes.total
C1315986|T201|COMP|33517-4|LNC|Hemoglobin|Hemoglobin
C1315989|T201|COMP|33520-8|LNC|Platelet aggregation.collagen induced^high dose|Platelet aggregation.collagen induced^high dose
C1315990|T201|COMP|33521-6|LNC|Platelet aggregation.collagen induced^low dose|Platelet aggregation.collagen induced^low dose
C1315991|T201|COMP|33522-4|LNC|Platelet aggregation.ristocetin induced^high dose|Platelet aggregation.ristocetin induced^high dose
C1315992|T201|COMP|33523-2|LNC|Platelet aggregation.ristocetin induced^low dose|Platelet aggregation.ristocetin induced^low dose
C1315993|T201|COMP|33524-0|LNC|Coagulum lysis|Coagulum lysis
C1315996|T201|COMP|33527-3|LNC|Methadone.long acting metabolite|Methadone.long acting metabolite
C1315999|T201|COMP|33530-7|LNC|Platelet aggregation.EPINEPHrine induced|Platelet aggregation.EPINEPHrine induced
C1316000|T201|COMP|33531-5|LNC|Platelet aggregation.arachidonate induced|Platelet aggregation.arachidonate induced
C1316001|T201|COMP|33532-3|LNC|Platelet aggregation.ristocetin induced^high dose|Platelet aggregation.ristocetin induced^high dose
C1316002|T201|COMP|33533-1|LNC|Platelet aggregation.ristocetin induced^low dose|Platelet aggregation.ristocetin induced^low dose
C1316003|T201|COMP|33534-9|LNC|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C1316004|T201|COMP|33535-6|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C1316005|T201|COMP|33536-4|LNC|Allergen.miscellaneous Ab.IgE.RAST class|Allergen.miscellaneous Ab.IgE.RAST class
C1316017|T201|COMP|33548-9|LNC|Lymphocytes.abnormal/100 leukocytes|Lymphocytes.abnormal/100 leukocytes
C1316018|T201|COMP|33549-7|LNC|Hantavirus sin nombre Ab|Hantavirus sin nombre Ab
C1316021|T201|COMP|33552-1|LNC|Platelet aggregation.ristocetin induced^900 ug/mL|Platelet aggregation.ristocetin induced^900 ug/mL
C1316022|T201|COMP|33553-9|LNC|Platelet aggregation.ristocetin induced^600 ug/mL|Platelet aggregation.ristocetin induced^600 ug/mL
C1316023|T201|COMP|33554-7|LNC|Platelet aggregation.ristocetin induced^300 ug/mL|Platelet aggregation.ristocetin induced^300 ug/mL
C1316027|T201|COMP|33558-8|LNC|Creatinine renal clearance|Creatinine renal clearance
C1316029|T201|COMP|33560-4|LNC|Benzodiazepines|Benzodiazepines
C1316030|T201|COMP|33561-2|LNC|Cannabinoids|Cannabinoids
C1316031|T201|COMP|33562-0|LNC|Ampicillin^peak|Ampicillin^peak
C1316032|T201|COMP|33563-8|LNC|Pancreatic islet cell Ab.IgG|Pancreatic islet cell Ab.IgG
C1316033|T201|COMP|33564-6|LNC|Smith extractable nuclear Ab.IgG|Smith extractable nuclear Ab.IgG
C1316034|T201|COMP|33565-3|LNC|Smith extractable nuclear Ab.IgG|Smith extractable nuclear Ab.IgG
C1316035|T201|COMP|33566-1|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C1316038|T201|COMP|33569-5|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C1316039|T201|COMP|33570-3|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C1316040|T201|COMP|33571-1|LNC|Jo-1 extractable nuclear Ab.IgG|Jo-1 extractable nuclear Ab.IgG
C1316041|T201|COMP|33572-9|LNC|Aureobasidium pullulans Ab.IgG|Aureobasidium pullulans Ab.IgG
C1316043|T201|COMP|33574-5|LNC|Chlamydia trachomatis I Ab.IgM|Chlamydia trachomatis I Ab.IgM
C1316044|T201|COMP|33575-2|LNC|Chlamydia trachomatis I Ab|Chlamydia trachomatis I Ab
C1316045|T201|COMP|33576-0|LNC|Francisella tularensis Ab.IgA|Francisella tularensis Ab.IgA
C1316046|T201|COMP|33577-8|LNC|Rheumatoid factor.IgM|Rheumatoid factor.IgM
C1316047|T201|COMP|33578-6|LNC|Dengue virus Ab|Dengue virus Ab
C1316048|T201|COMP|33579-4|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1316049|T201|COMP|33580-2|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1316050|T201|COMP|33581-0|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C1316051|T201|COMP|33583-6|LNC|Sjogrens syndrome-A extractable nuclear Ab.IgG|Sjogrens syndrome-A extractable nuclear Ab.IgG
C1316052|T201|COMP|33584-4|LNC|Gastrin^10M pre XXX challenge|Gastrin^10M pre XXX challenge
C1316053|T201|COMP|33585-1|LNC|Uroporphyrin 3 isomer|Uroporphyrin 3 isomer
C1316054|T201|COMP|33587-7|LNC|Trichinella sp Ab.IgA|Trichinella sp Ab.IgA
C1316055|T201|COMP|33588-5|LNC|Phosphatidylethanolamine Ab|Phosphatidylethanolamine Ab
C1316056|T201|COMP|33589-3|LNC|Phosphatidylinositol Ab|Phosphatidylinositol Ab
C1316057|T201|COMP|33590-1|LNC|Neuronal nuclear Ab.IgG|Neuronal nuclear Ab.IgG
C1316058|T201|COMP|33591-9|LNC|Neuronal nuclear Ab.IgG|Neuronal nuclear Ab.IgG
C1316059|T201|COMP|33592-7|LNC|Cells.CD10+HLA-DR+|Cells.CD10+HLA-DR+
C1316060|T201|COMP|33593-5|LNC|Hemoglobin G-Coushatta/Hemoglobin.total|Hemoglobin G-Coushatta/Hemoglobin.total
C1316061|T201|COMP|33594-3|LNC|Platelet factor 4|Platelet factor 4
C1316062|T201|COMP|33597-6|LNC|Borrelia burgdorferi 34kD Ab.IgM|Borrelia burgdorferi 34kD Ab.IgM
C1316063|T201|COMP|33598-4|LNC|Sjogrens syndrome-B extractable nuclear Ab.IgG|Sjogrens syndrome-B extractable nuclear Ab.IgG
C1316064|T201|COMP|33599-2|LNC|Amylase|Amylase
C1316065|T201|COMP|33600-8|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C1316066|T201|COMP|33601-6|LNC|Cells.CD23+CD38+|Cells.CD23+CD38+
C1316067|T201|COMP|33602-4|LNC|Myelin associated glycoprotein Ab.IgG|Myelin associated glycoprotein Ab.IgG
C1316069|T201|COMP|33604-0|LNC|Chlamydia trachomatis I Ab.IgM|Chlamydia trachomatis I Ab.IgM
C1316070|T201|COMP|33605-7|LNC|Chlamydia trachomatis I Ab|Chlamydia trachomatis I Ab
C1316071|T201|COMP|33606-5|LNC|Dengue virus Ab|Dengue virus Ab
C1316072|T201|COMP|33607-3|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1316073|T201|COMP|33608-1|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1316074|T201|COMP|33609-9|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C1316075|T201|COMP|33610-7|LNC|Sjogrens syndrome-A extractable nuclear Ab.IgG|Sjogrens syndrome-A extractable nuclear Ab.IgG
C1316076|T201|COMP|33611-5|LNC|Phosphatidylethanolamine Ab|Phosphatidylethanolamine Ab
C1316077|T201|COMP|33612-3|LNC|Phosphatidylinositol Ab|Phosphatidylinositol Ab
C1316078|T201|COMP|33613-1|LNC|Sjogrens syndrome-B extractable nuclear Ab.IgG|Sjogrens syndrome-B extractable nuclear Ab.IgG
C1316080|T201|COMP|33615-6|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C1316081|T201|COMP|33616-4|LNC|Cytomegalovirus early Ag|Cytomegalovirus early Ag
C1316082|T201|COMP|33618-0|LNC|Coproporphyrin 3/Coproporphyrin 1|Coproporphyrin 3/Coproporphyrin 1
C1316083|T201|COMP|33619-8|LNC|Deuteroporphyrin.semi-proto|Deuteroporphyrin.semi-proto
C1316084|T201|COMP|33620-6|LNC|Tricarboxylporphyrin 1|Tricarboxylporphyrin 1
C1316085|T201|COMP|33621-4|LNC|Tricarboxylporphyrin 3|Tricarboxylporphyrin 3
C1316086|T201|COMP|33622-2|LNC|Isotricarboxylporphyrin|Isotricarboxylporphyrin
C1316087|T201|COMP|33623-0|LNC|Pentacarboxylporphyrin I|Pentacarboxylporphyrin I
C1316088|T201|COMP|33624-8|LNC|Pentacarboxylporphyrin III|Pentacarboxylporphyrin III
C1316089|T201|COMP|33625-5|LNC|Isocoproporphyrin|Isocoproporphyrin
C1316090|T201|COMP|33626-3|LNC|Hematoporphyrin|Hematoporphyrin
C1316091|T201|COMP|33627-1|LNC|Tenofovir|Tenofovir
C1316092|T201|COMP|33628-9|LNC|Cidofovir|Cidofovir
C1316093|T201|COMP|33629-7|LNC|Hepatitis B virus sequencing|Hepatitis B virus sequencing
C1316094|T201|COMP|33630-5|LNC|HIV protease gene mutations detected|HIV protease gene mutations detected
C1316095|T201|COMP|33631-3|LNC|Cytomegalovirus UL54 gene mutations detected|Cytomegalovirus UL54 gene mutations detected
C1316096|T201|COMP|33632-1|LNC|Cytomegalovirus UL54+UL97 gene mutations detected|Cytomegalovirus UL54+UL97 gene mutations detected
C1316097|T201|COMP|33633-9|LNC|Hepatitis B virus precore TAG mutation|Hepatitis B virus precore TAG mutation
C1316099|T201|COMP|33635-4|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C1316100|T201|COMP|33636-2|LNC|IgA.secretory|IgA.secretory
C1316101|T201|COMP|33637-0|LNC|Phagocytic index|Phagocytic index
C1316105|T201|COMP|33641-2|LNC|Lymphocyte proliferation.tuberculin stimulation|Lymphocyte proliferation.tuberculin stimulation
C1316106|T201|COMP|33642-0|LNC|Lymphocyte Ab|Lymphocyte Ab
C1316107|T201|COMP|33643-8|LNC|Limulus amebocyte lysate test|Limulus amebocyte lysate test
C1316108|T201|COMP|33644-6|LNC|A1 Ab|A1 Ab
C1316109|T201|COMP|33645-3|LNC|A2 Ab|A2 Ab
C1316110|T201|COMP|33646-1|LNC|Methylenedianiline|Methylenedianiline
C1316111|T201|COMP|33647-9|LNC|Protein.monoclonal/Protein.total|Protein.monoclonal/Protein.total
C1316112|T201|COMP|33648-7|LNC|Cryoglobulin.rheumatoid factor|Cryoglobulin.rheumatoid factor
C1316113|T201|COMP|33649-5|LNC|Cryoglobulin.IgG|Cryoglobulin.IgG
C1316114|T201|COMP|33650-3|LNC|Cryoglobulin.IgA|Cryoglobulin.IgA
C1316115|T201|COMP|33651-1|LNC|Cryoglobulin.IgM|Cryoglobulin.IgM
C1316116|T201|COMP|33652-9|LNC|Cells.CD56/Cells.CD38|Cells.CD56/Cells.CD38
C1316117|T201|COMP|33653-7|LNC|Beta galactosidase|Beta galactosidase
C1316119|T201|COMP|33655-2|LNC|Beta-N-acetylhexosaminidase|Beta-N-acetylhexosaminidase
C1316120|T201|COMP|33656-0|LNC|Beta-N-acetylhexosaminidase.B|Beta-N-acetylhexosaminidase.B
C1316121|T201|COMP|33657-8|LNC|Beta-N-acetylhexosaminidase.A|Beta-N-acetylhexosaminidase.A
C1316123|T201|COMP|33659-4|LNC|Pipecolate/Creatinine|Pipecolate/Creatinine
C1316124|T201|COMP|33660-2|LNC|HIV 1 p24 Ag|HIV 1 p24 Ag
C1316125|T201|COMP|33661-0|LNC|Glucosylceramidase|Glucosylceramidase
C1316126|T201|COMP|33662-8|LNC|Erythrocytes.CD59 deficient/100 Cells.235a|Erythrocytes.CD59 deficient/100 Cells.235a
C1316127|T201|COMP|33663-6|LNC|Cells.CD59 deficient/100 cells|Cells.CD59 deficient/100 cells
C1316128|T201|COMP|33664-4|LNC|Cells.CD59|Cells.CD59
C1316129|T201|COMP|33665-1|LNC|HTLV I+II Ab band pattern|HTLV I+II Ab band pattern
C1316130|T201|COMP|33666-9|LNC|Erythrocytes.dysmorphic|Erythrocytes.dysmorphic
C1316131|T201|COMP|33667-7|LNC|Prostate specific Ag.protein bound|Prostate specific Ag.protein bound
C1316132|T201|COMP|33668-5|LNC|Erythrocytes|Erythrocytes
C1316133|T201|COMP|33669-3|LNC|Trypsin|Trypsin
C1316140|T201|COMP|33676-8|LNC|Francisella tularensis|Francisella tularensis
C1316141|T201|COMP|33677-6|LNC|Francisella tularensis|Francisella tularensis
C1316142|T201|COMP|33678-4|LNC|Francisella tularensis Ag|Francisella tularensis Ag
C1316143|T201|COMP|33679-2|LNC|Francisella tularensis DNA|Francisella tularensis DNA
C1316144|T201|COMP|33680-0|LNC|Francisella tularensis DNA|Francisella tularensis DNA
C1316145|T201|COMP|33681-8|LNC|Francisella tularensis|Francisella tularensis
C1316146|T201|COMP|33682-6|LNC|Francisella tularensis|Francisella tularensis
C1316147|T201|COMP|33683-4|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C1316148|T201|COMP|33684-2|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C1316149|T201|COMP|33685-9|LNC|Yersinia pestis|Yersinia pestis
C1316150|T201|COMP|33686-7|LNC|Yersinia pestis|Yersinia pestis
C1316151|T201|COMP|33687-5|LNC|Yersinia pestis Ag|Yersinia pestis Ag
C1316152|T201|COMP|33688-3|LNC|Yersinia pestis Ag|Yersinia pestis Ag
C1316153|T201|COMP|33689-1|LNC|Yersinia pestis Ab|Yersinia pestis Ab
C1316154|T201|COMP|33690-9|LNC|Yersinia pestis Ab|Yersinia pestis Ab
C1316155|T201|COMP|33691-7|LNC|Yersinia pestis DNA|Yersinia pestis DNA
C1316156|T201|COMP|33692-5|LNC|Yersinia pestis DNA|Yersinia pestis DNA
C1316157|T201|COMP|33693-3|LNC|Yersinia pestis|Yersinia pestis
C1316158|T201|COMP|33694-1|LNC|Clostridium botulinum|Clostridium botulinum
C1316159|T201|COMP|33695-8|LNC|Clostridium botulinum|Clostridium botulinum
C1316160|T201|COMP|33696-6|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C1316161|T201|COMP|33697-4|LNC|Bacillus anthracis Ag|Bacillus anthracis Ag
C1316162|T201|COMP|33698-2|LNC|Bacillus anthracis|Bacillus anthracis
C1316164|T201|COMP|33700-6|LNC|Spore identification|Spore identification
C1316165|T201|COMP|33701-4|LNC|Clostridium botulinum toxin A|Clostridium botulinum toxin A
C1316166|T201|COMP|33702-2|LNC|Clostridium botulinum toxin E|Clostridium botulinum toxin E
C1316167|T201|COMP|33703-0|LNC|Clostridium botulinum toxin F|Clostridium botulinum toxin F
C1316168|T201|COMP|33704-8|LNC|Clostridium botulinum toxin A+B+E|Clostridium botulinum toxin A+B+E
C1316169|T201|COMP|33705-5|LNC|Clostridium botulinum toxin B|Clostridium botulinum toxin B
C1316170|T201|COMP|33706-3|LNC|Yersinia pestis Ab|Yersinia pestis Ab
C1316171|T201|COMP|33707-1|LNC|Yersinia pestis Ab|Yersinia pestis Ab
C1316172|T201|COMP|33708-9|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C1316173|T201|COMP|33709-7|LNC|Clostridium botulinum toxin A|Clostridium botulinum toxin A
C1316174|T201|COMP|33710-5|LNC|Clostridium botulinum toxin E|Clostridium botulinum toxin E
C1316175|T201|COMP|33711-3|LNC|Clostridium botulinum toxin F|Clostridium botulinum toxin F
C1316176|T201|COMP|33712-1|LNC|Clostridium botulinum toxin A+B+E|Clostridium botulinum toxin A+B+E
C1316177|T201|COMP|33713-9|LNC|Clostridium botulinum toxin B|Clostridium botulinum toxin B
C1316178|T201|COMP|33714-7|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C1316179|T201|COMP|33715-4|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C1316182|T201|COMP|33718-8|LNC|Cytology report|Cytology report
C1316185|T201|COMP|33721-2|LNC|Pathology biopsy report|Pathology biopsy report
C1316186|T201|COMP|33722-0|LNC|Collection method|Collection method
C1316187|T201|COMP|33723-8|LNC|Specimen length|Specimen length
C1316188|T201|COMP|33724-6|LNC|Collection method|Collection method
C1316189|T201|COMP|33725-3|LNC|Tumor site|Tumor site
C1316190|T201|COMP|33726-1|LNC|Macroscopic tumor configuration|Macroscopic tumor configuration
C1316191|T201|COMP|33727-9|LNC|Macroscopic tumor configuration|Macroscopic tumor configuration
C1316192|T201|COMP|33728-7|LNC|Size.max.dimension|Size.max.dimension
C1316193|T201|COMP|33729-5|LNC|Size.additional dimension|Size.additional dimension
C1316194|T201|COMP|33730-3|LNC|Resection completeness|Resection completeness
C1316195|T201|COMP|33731-1|LNC|Histology type|Histology type
C1316196|T201|COMP|33732-9|LNC|Histology grade|Histology grade
C1316197|T201|COMP|33733-7|LNC|Sites of distant metastasis|Sites of distant metastasis
C1316198|T201|COMP|33734-5|LNC|Surgical margin tumor involvement.proximal|Surgical margin tumor involvement.proximal
C1316199|T201|COMP|33735-2|LNC|Surgical margin tumor involvement.distant|Surgical margin tumor involvement.distant
C1316200|T201|COMP|33736-0|LNC|Surgical margin tumor involvement.circumferential|Surgical margin tumor involvement.circumferential
C1316201|T201|COMP|33737-8|LNC|Distance of tumor from closest margin|Distance of tumor from closest margin
C1316202|T201|COMP|33738-6|LNC|Closest margin|Closest margin
C1316203|T201|COMP|33739-4|LNC|Lymphatic.small vessel.invasion|Lymphatic.small vessel.invasion
C1316204|T201|COMP|33740-2|LNC|Venous.large vessel.invasion|Venous.large vessel.invasion
C1316205|T201|COMP|33741-0|LNC|Perineural invasion|Perineural invasion
C1316206|T201|COMP|33742-8|LNC|Tumor border configuration|Tumor border configuration
C1316207|T201|COMP|33743-6|LNC|Intratumoral + Peritumoral lymphocytic response|Intratumoral + Peritumoral lymphocytic response
C1316208|T201|COMP|33744-4|LNC|Additional pathological findings|Additional pathological findings
C1316209|T201|COMP|33745-1|LNC|Polyps|Polyps
C1316210|T201|COMP|33746-9|LNC|Pathologic findings|Pathologic findings
C1316211|T201|COMP|33747-7|LNC|Number of fragmented pieces|Number of fragmented pieces
C1316212|T201|COMP|33748-5|LNC|Distance from anal verge|Distance from anal verge
C1316213|T201|COMP|33749-3|LNC|Distance from anal verge unknown|Distance from anal verge unknown
C1316214|T201|COMP|33750-1|LNC|Margins cannot be assessed|Margins cannot be assessed
C1316215|T201|COMP|33751-9|LNC|Surgical margin tumor involvement.lateral|Surgical margin tumor involvement.lateral
C1316216|T201|COMP|33752-7|LNC|Distance of carcinoma from closest lateral margin|Distance of carcinoma from closest lateral margin
C1316217|T201|COMP|33753-5|LNC|Lateral margin location|Lateral margin location
C1316218|T201|COMP|33754-3|LNC|Surgical margin tumor involvement.deep|Surgical margin tumor involvement.deep
C1316219|T201|COMP|33755-0|LNC|Distance of carcinoma from deep margin|Distance of carcinoma from deep margin
C1316220|T201|COMP|33756-8|LNC|Polyp size greatest dimension|Polyp size greatest dimension
C1316221|T201|COMP|33757-6|LNC|Polyp size additional dimensions|Polyp size additional dimensions
C1316222|T201|COMP|33758-4|LNC|Polyp stalk length|Polyp stalk length
C1316223|T201|COMP|33759-2|LNC|Extent of invasion deepest|Extent of invasion deepest
C1316224|T201|COMP|33760-0|LNC|Surgical margin tumor involvement.mucosal|Surgical margin tumor involvement.mucosal
C1316225|T201|COMP|33761-8|LNC|Venous + Lymphatic small vessel invasion|Venous + Lymphatic small vessel invasion
C1316226|T201|COMP|33762-6|LNC|Natriuretic peptide.B prohormone N-Terminal|Natriuretic peptide.B prohormone N-Terminal
C1316227|T201|COMP|33763-4|LNC|Natriuretic peptide.B prohormone N-Terminal|Natriuretic peptide.B prohormone N-Terminal
C1316228|T201|COMP|33764-2|LNC|Shiga toxin stx gene|Shiga toxin stx gene
C1316229|T201|COMP|33765-9|LNC|Leukocytes|Leukocytes
C1316230|T201|COMP|33766-7|LNC|Radioactivity^pre dose radioactive cyanocobalamin|Radioactivity^pre dose radioactive cyanocobalamin
C1316231|T201|COMP|33767-5|LNC|Acidity.total|Acidity.total
C1316232|T201|COMP|33768-3|LNC|Leukocyte clumps|Leukocyte clumps
C1316233|T201|COMP|33769-1|LNC|Mucin clot^15M post incubation|Mucin clot^15M post incubation
C1316234|T201|COMP|33770-9|LNC|Mucin clot^30M post incubation|Mucin clot^30M post incubation
C1316235|T201|COMP|33771-7|LNC|Pl-12 Ab|Pl-12 Ab
C1316236|T201|COMP|33772-5|LNC|Pl-7 Ab|Pl-7 Ab
C1316237|T201|COMP|33773-3|LNC|Karyotype|Karyotype
C1316238|T201|COMP|33774-1|LNC|Karyotype|Karyotype
C1316239|T201|COMP|33775-8|LNC|Cells.CD41a/100 cells|Cells.CD41a/100 cells
C1316240|T201|COMP|32750-2|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C1316241|T201|COMP|33777-4|LNC|Cells.SmIg/100 cells|Cells.SmIg/100 cells
C1316242|T201|COMP|33778-2|LNC|SmIg Ag|SmIg Ag
C1316243|T201|COMP|33779-0|LNC|IgG+IgM+IgA heavy chain Ag|IgG+IgM+IgA heavy chain Ag
C1316245|T201|COMP|33781-6|LNC|Alpha-1-Acid glycoprotein|Alpha-1-Acid glycoprotein
C1316246|T201|COMP|33782-4|LNC|Alpha-2-Retinol binding protein|Alpha-2-Retinol binding protein
C1316247|T201|COMP|33783-2|LNC|Atrial natriuretic factor|Atrial natriuretic factor
C1316248|T201|COMP|33784-0|LNC|Bacterial casts|Bacterial casts
C1316249|T201|COMP|33785-7|LNC|Basophils.immature|Basophils.immature
C1316250|T201|COMP|33786-5|LNC|Basophils.immature/100 leukocytes|Basophils.immature/100 leukocytes
C1316251|T201|COMP|33787-3|LNC|Calcitonin^10th specimen post XXX challenge|Calcitonin^10th specimen post XXX challenge
C1316252|T201|COMP|33788-1|LNC|Calcitonin^1st specimen post XXX challenge|Calcitonin^1st specimen post XXX challenge
C1316253|T201|COMP|33789-9|LNC|Calcium^10th specimen post XXX challenge|Calcium^10th specimen post XXX challenge
C1316254|T201|COMP|33790-7|LNC|Calcium^1st specimen post XXX challenge|Calcium^1st specimen post XXX challenge
C1316255|T201|COMP|33791-5|LNC|Calcium^5th specimen post XXX challenge|Calcium^5th specimen post XXX challenge
C1316256|T201|COMP|33792-3|LNC|Calcium^6th specimen post XXX challenge|Calcium^6th specimen post XXX challenge
C1316257|T201|COMP|33793-1|LNC|Calcium^7th specimen post XXX challenge|Calcium^7th specimen post XXX challenge
C1316258|T201|COMP|33794-9|LNC|Calcium^8th specimen post XXX challenge|Calcium^8th specimen post XXX challenge
C1316259|T201|COMP|33795-6|LNC|Calcium^9th specimen post XXX challenge|Calcium^9th specimen post XXX challenge
C1316260|T201|COMP|33796-4|LNC|Cotinine|Cotinine
C1316261|T201|COMP|33797-2|LNC|Creatine|Creatine
C1316262|T201|COMP|33798-0|LNC|Creatinine|Creatinine
C1316263|T201|COMP|33799-8|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C1316264|T201|COMP|33800-4|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C1316265|T201|COMP|33801-2|LNC|E selectin|E selectin
C1316266|T201|COMP|33802-0|LNC|Eosinophils.immature|Eosinophils.immature
C1316267|T201|COMP|33803-8|LNC|Eosinophils.immature/100 leukocytes|Eosinophils.immature/100 leukocytes
C1316268|T201|COMP|33804-6|LNC|Erythrocyte casts|Erythrocyte casts
C1316269|T201|COMP|33805-3|LNC|Fructosamine|Fructosamine
C1316270|T201|COMP|33806-1|LNC|HIV 2 Ab.IgG|HIV 2 Ab.IgG
C1316271|T201|COMP|33807-9|LNC|HIV 2 Ab.IgG|HIV 2 Ab.IgG
C1316272|T201|COMP|33808-7|LNC|Insulin-like growth factor binding protein 3|Insulin-like growth factor binding protein 3
C1316273|T201|COMP|33809-5|LNC|Insulin^10th specimen post XXX challenge|Insulin^10th specimen post XXX challenge
C1316274|T201|COMP|33810-3|LNC|Insulin^11th specimen post XXX challenge|Insulin^11th specimen post XXX challenge
C1316275|T201|COMP|33811-1|LNC|Insulin^12th specimen post XXX challenge|Insulin^12th specimen post XXX challenge
C1316276|T201|COMP|33812-9|LNC|Insulin^13th specimen post XXX challenge|Insulin^13th specimen post XXX challenge
C1316277|T201|COMP|33813-7|LNC|Insulin^14th specimen post XXX challenge|Insulin^14th specimen post XXX challenge
C1316278|T201|COMP|33814-5|LNC|Insulin^15th specimen post XXX challenge|Insulin^15th specimen post XXX challenge
C1316279|T201|COMP|33815-2|LNC|Insulin^1st specimen post XXX challenge|Insulin^1st specimen post XXX challenge
C1316280|T201|COMP|33816-0|LNC|Insulin^2nd specimen post XXX challenge|Insulin^2nd specimen post XXX challenge
C1316281|T201|COMP|33817-8|LNC|Insulin^3rd specimen post XXX challenge|Insulin^3rd specimen post XXX challenge
C1316282|T201|COMP|33818-6|LNC|Insulin^8th specimen post XXX challenge|Insulin^8th specimen post XXX challenge
C1316283|T201|COMP|33819-4|LNC|Insulin^9th specimen post XXX challenge|Insulin^9th specimen post XXX challenge
C1316284|T201|COMP|33820-2|LNC|Interferon.alpha|Interferon.alpha
C1316285|T201|COMP|33821-0|LNC|Interleukin 1 alpha|Interleukin 1 alpha
C1316286|T201|COMP|33822-8|LNC|Interleukin 13|Interleukin 13
C1316287|T201|COMP|33823-6|LNC|Interleukin 18|Interleukin 18
C1316288|T201|COMP|33824-4|LNC|Iron|Iron
C1316289|T201|COMP|33825-1|LNC|Leukocyte casts|Leukocyte casts
C1316290|T201|COMP|33826-9|LNC|Lutropin^10th specimen post XXX challenge|Lutropin^10th specimen post XXX challenge
C1316291|T201|COMP|33827-7|LNC|Lutropin^1st specimen post XXX challenge|Lutropin^1st specimen post XXX challenge
C1316292|T201|COMP|33828-5|LNC|Lutropin^8th specimen post XXX challenge|Lutropin^8th specimen post XXX challenge
C1316293|T201|COMP|33829-3|LNC|Lutropin^9th specimen post XXX challenge|Lutropin^9th specimen post XXX challenge
C1316294|T201|COMP|33830-1|LNC|Lymphoblasts|Lymphoblasts
C1316295|T201|COMP|33831-9|LNC|Lymphoblasts/100 leukocytes|Lymphoblasts/100 leukocytes
C1316296|T201|COMP|33832-7|LNC|Lymphocytes.immunoblastic|Lymphocytes.immunoblastic
C1316297|T201|COMP|33833-5|LNC|Lymphocytes.immunoblastic/100 leukocytes|Lymphocytes.immunoblastic/100 leukocytes
C1316298|T201|COMP|33834-3|LNC|Lymphocytes.plasmacytoid|Lymphocytes.plasmacytoid
C1316299|T201|COMP|33835-0|LNC|Lymphocytes.plasmacytoid/100 leukocytes|Lymphocytes.plasmacytoid/100 leukocytes
C1316300|T201|COMP|33836-8|LNC|Malignant cells|Malignant cells
C1316301|T201|COMP|33837-6|LNC|Malignant cells/100 leukocytes|Malignant cells/100 leukocytes
C1316302|T201|COMP|33838-4|LNC|Mannitol|Mannitol
C1316303|T201|COMP|33839-2|LNC|Monoblasts|Monoblasts
C1316304|T201|COMP|33840-0|LNC|Monoblasts/100 leukocytes|Monoblasts/100 leukocytes
C1316305|T201|COMP|33841-8|LNC|Monocytes.immature|Monocytes.immature
C1316306|T201|COMP|33842-6|LNC|Monocytes.immature/100 leukocytes|Monocytes.immature/100 leukocytes
C1316307|T201|COMP|33843-4|LNC|Norepinephrine^standing|Norepinephrine^standing
C1316308|T201|COMP|33844-2|LNC|Norepinephrine^supine|Norepinephrine^supine
C1316309|T201|COMP|33845-9|LNC|Parathyrin.intact^1H post XXX challenge|Parathyrin.intact^1H post XXX challenge
C1316310|T201|COMP|33846-7|LNC|Parathyrin.intact^2H post XXX challenge|Parathyrin.intact^2H post XXX challenge
C1316311|T201|COMP|33847-5|LNC|Parathyrin.intact^30M post XXX challenge|Parathyrin.intact^30M post XXX challenge
C1316312|T201|COMP|33848-3|LNC|Plasma cell precursor|Plasma cell precursor
C1316313|T201|COMP|33849-1|LNC|Plasma cell precursor/100 leukocytes|Plasma cell precursor/100 leukocytes
C1316314|T201|COMP|33850-9|LNC|Plasma cells.immature|Plasma cells.immature
C1316315|T201|COMP|33851-7|LNC|Progesterone^10th specimen post XXX challenge|Progesterone^10th specimen post XXX challenge
C1316316|T201|COMP|33852-5|LNC|Progesterone^1st specimen post XXX challenge|Progesterone^1st specimen post XXX challenge
C1316317|T201|COMP|33853-3|LNC|Progesterone^1st specimen post XXX challenge|Progesterone^1st specimen post XXX challenge
C1316318|T201|COMP|33854-1|LNC|Progesterone^4th specimen post XXX challenge|Progesterone^4th specimen post XXX challenge
C1316319|T201|COMP|33856-6|LNC|Sezary cells|Sezary cells
C1316320|T201|COMP|33857-4|LNC|Sezary cells/100 leukocytes|Sezary cells/100 leukocytes
C1316321|T201|COMP|33858-2|LNC|Somatotropin|Somatotropin
C1316322|T201|COMP|33859-0|LNC|Somatotropin/Creatinine|Somatotropin/Creatinine
C1316323|T201|COMP|33860-8|LNC|Somatotropin/Creatinine|Somatotropin/Creatinine
C1316324|T201|COMP|33861-6|LNC|Starch granules|Starch granules
C1316325|T201|COMP|33862-4|LNC|Waxy casts|Waxy casts
C1316326|T201|COMP|33863-2|LNC|Cystatin C|Cystatin C
C1316327|T201|COMP|33864-0|LNC|Elastase.leukocyte|Elastase.leukocyte
C1316328|T201|COMP|33865-7|LNC|Staphylococcus aureus enterotoxin|Staphylococcus aureus enterotoxin
C1316329|T201|COMP|33866-5|LNC|HIV 1 Ab|HIV 1 Ab
C1316333|T201|COMP|33870-7|LNC|Bilirubin|Bilirubin
C1316334|T201|COMP|33871-5|LNC|Xylose^1H post 5 g xylose PO|Xylose^1H post 5 g xylose PO
C1316335|T201|COMP|33872-3|LNC|Cystine|Cystine
C1316336|T201|COMP|33873-1|LNC|DOPamine/Creatinine|DOPamine/Creatinine
C1316337|T201|COMP|33874-9|LNC|EPINEPHrine/Creatinine|EPINEPHrine/Creatinine
C1316338|T201|COMP|33875-6|LNC|Oligosaccharides pattern|Oligosaccharides pattern
C1316339|T201|COMP|33876-4|LNC|Sulfocysteine/Creatinine|Sulfocysteine/Creatinine
C1316340|T201|COMP|33877-2|LNC|Tetrahydrobiopterin/Biopterin|Tetrahydrobiopterin/Biopterin
C1316342|T201|COMP|33879-8|LNC|Protein.monoclonal|Protein.monoclonal
C1316345|T201|COMP|33882-2|LNC|Collection date|Collection date
C1316356|T201|COMP|33893-9|LNC|Karyotype|Karyotype
C1316359|T201|COMP|33896-2|LNC|Orientia tsutsugamushi Ab.IgM|Orientia tsutsugamushi Ab.IgM
C1316360|T201|COMP|33897-0|LNC|Orientia tsutsugamushi Ab.IgM|Orientia tsutsugamushi Ab.IgM
C1316363|T201|COMP|33900-2|LNC|Fetal cell screen|Fetal cell screen
C1316364|T201|COMP|33901-0|LNC|Gestational age|Gestational age
C1316365|T201|COMP|33902-8|LNC|Immune complex|Immune complex
C1316366|T201|COMP|33903-6|LNC|Ketones|Ketones
C1316367|T201|COMP|33904-4|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1316368|T201|COMP|33905-1|LNC|Trichomonas sp|Trichomonas sp
C1316369|T201|COMP|33906-9|LNC|Prolactin^30M post 200 ug TRH IV|Prolactin^30M post 200 ug TRH IV
C1316370|T201|COMP|33907-7|LNC|Prolactin^1H post 200 ug TRH IV|Prolactin^1H post 200 ug TRH IV
C1316371|T201|COMP|33908-5|LNC|Prolactin^1.5H post 200 ug TRH IV|Prolactin^1.5H post 200 ug TRH IV
C1316372|T201|COMP|33909-3|LNC|Prolactin^2H post 200 ug TRH IV|Prolactin^2H post 200 ug TRH IV
C1316373|T201|COMP|33910-1|LNC|Rheumatoid factor|Rheumatoid factor
C1316374|T201|COMP|33911-9|LNC|Complement C1r actual/Normal|Complement C1r actual/Normal
C1316375|T201|COMP|33912-7|LNC|Complement C1s actual/Normal|Complement C1s actual/Normal
C1316377|T201|COMP|33914-3|LNC|Glomerular filtration rate/1.73 sq M.predicted|Glomerular filtration rate/1.73 sq M.predicted
C1316378|T201|COMP|33915-0|LNC|Anabasine|Anabasine
C1316379|T201|COMP|33916-8|LNC|Trans-3-Hydroxycotinine|Trans-3-Hydroxycotinine
C1316380|T201|COMP|33917-6|LNC|Nornicotine|Nornicotine
C1316381|T201|COMP|33918-4|LNC|Acetoacetate|Acetoacetate
C1316382|T201|COMP|33919-2|LNC|Ampicillin^trough|Ampicillin^trough
C1316383|T201|COMP|33920-0|LNC|S Ab|S Ab
C1316384|T201|COMP|33921-8|LNC|Signal recognition particle Ab|Signal recognition particle Ab
C1316385|T201|COMP|33922-6|LNC|Wasp venom Ab.IgE.RAST class|Wasp venom Ab.IgE.RAST class
C1316386|T201|COMP|33923-4|LNC|Hemosiderin|Hemosiderin
C1316387|T201|COMP|33924-2|LNC|Neuronal nuclear type 3 Ab|Neuronal nuclear type 3 Ab
C1316388|T201|COMP|33925-9|LNC|Purkinje cell cytoplasmic type 2 Ab|Purkinje cell cytoplasmic type 2 Ab
C1316389|T201|COMP|33926-7|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C1316390|T201|COMP|33927-5|LNC|Amphiphysin Ab|Amphiphysin Ab
C1316391|T201|COMP|33928-3|LNC|Efavirenz|Efavirenz
C1316392|T201|COMP|33929-1|LNC|Tacrolimus^trough|Tacrolimus^trough
C1316395|T201|COMP|33932-5|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C1316396|T201|COMP|33933-3|LNC|Glutaraldehyde Ab.IgE|Glutaraldehyde Ab.IgE
C1316397|T201|COMP|33934-1|LNC|Methylmethacrylate Ab.IgE|Methylmethacrylate Ab.IgE
C1316398|T201|COMP|33935-8|LNC|Cyclic citrullinated peptide Ab.IgG|Cyclic citrullinated peptide Ab.IgG
C1316399|T201|COMP|33936-6|LNC|Homocystine.free|Homocystine.free
C1316400|T201|COMP|33937-4|LNC|Homocystine.free|Homocystine.free
C1316401|T201|COMP|33938-2|LNC|Interleukin 5|Interleukin 5
C1316402|T201|COMP|33939-0|LNC|Interleukin 2|Interleukin 2
C1316403|T201|COMP|33940-8|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1316404|T201|COMP|33941-6|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1316405|T201|COMP|33942-4|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1316407|T201|COMP|33944-0|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C1316408|T201|COMP|33945-7|LNC|Brucella abortus Ab|Brucella abortus Ab
C1316409|T201|COMP|33946-5|LNC|Ziprasidone|Ziprasidone
C1316410|T201|COMP|33947-3|LNC|Clostridioides difficile toxin Ab|Clostridioides difficile toxin Ab
C1316411|T201|COMP|33948-1|LNC|IgG/Creatinine|IgG/Creatinine
C1316412|T201|COMP|33949-9|LNC|Potassium/Creatinine|Potassium/Creatinine
C1316413|T201|COMP|33950-7|LNC|Magnesium/Creatinine|Magnesium/Creatinine
C1316414|T201|COMP|33951-5|LNC|Sodium/Creatinine|Sodium/Creatinine
C1316415|T201|COMP|33952-3|LNC|Immune complex.IgM|Immune complex.IgM
C1316416|T201|COMP|33953-1|LNC|Immune complex.IgA|Immune complex.IgA
C1316417|T201|COMP|33954-9|LNC|Immune complex.IgG|Immune complex.IgG
C1316418|T201|COMP|33955-6|LNC|cycloSPORINE.monoclonal|cycloSPORINE.monoclonal
C1316419|T201|COMP|33956-4|LNC|cycloSPORINE.polyclonal|cycloSPORINE.polyclonal
C1316420|T201|COMP|33957-2|LNC|Normoblasts/100 blasts|Normoblasts/100 blasts
C1316421|T201|COMP|33958-0|LNC|Cholecalciferol|Cholecalciferol
C1316422|T201|COMP|33959-8|LNC|Procalcitonin|Procalcitonin
C1316423|T201|COMP|33960-6|LNC|Immune complex.IgE|Immune complex.IgE
C1316424|T201|COMP|33961-4|LNC|Sulthiame|Sulthiame
C1316425|T201|COMP|33962-2|LNC|Melanoma inhibitory activity protein|Melanoma inhibitory activity protein
C1316426|T201|COMP|33963-0|LNC|Granulocytes/100 leukocytes|Granulocytes/100 leukocytes
C1316427|T201|COMP|33964-8|LNC|SARS coronavirus Urbani RNA|SARS coronavirus Urbani RNA
C1316428|T201|COMP|33965-5|LNC|SARS coronavirus Urbani RNA|SARS coronavirus Urbani RNA
C1316429|T201|COMP|33966-3|LNC|SARS coronavirus Urbani RNA|SARS coronavirus Urbani RNA
C1316430|T201|COMP|33967-1|LNC|SARS coronavirus Urbani RNA|SARS coronavirus Urbani RNA
C1316431|T201|COMP|33968-9|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1316432|T201|COMP|33969-7|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1316433|T201|COMP|33970-5|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1316434|T201|COMP|33971-3|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1316435|T201|COMP|33972-1|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1316436|T201|COMP|33973-9|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1316437|T201|COMP|33974-7|LNC|SARS coronavirus Urbani Ab|SARS coronavirus Urbani Ab
C1316438|T201|COMP|33975-4|LNC|SARS coronavirus Urbani RNA|SARS coronavirus Urbani RNA
C1316439|T201|COMP|33976-2|LNC|Plasminogen activator inhibitor 1 Ag|Plasminogen activator inhibitor 1 Ag
C1316440|T201|COMP|33977-0|LNC|F little y super little a Ab|F little y super little a Ab
C1316441|T201|COMP|33978-8|LNC|BK virus DNA|BK virus DNA
C1316442|T201|COMP|33979-6|LNC|Voltage-gated calcium channel N type binding Ab|Voltage-gated calcium channel N type binding Ab
C1316443|T201|COMP|33980-4|LNC|Voltage-gated calcium channel PQ type binding Ab|Voltage-gated calcium channel PQ type binding Ab
C1316444|T201|COMP|33981-2|LNC|TBP gene.CAG repeats|TBP gene.CAG repeats
C1316445|T201|COMP|33982-0|LNC|Juglans california pollen Ab.IgE|Juglans california pollen Ab.IgE
C1316446|T201|COMP|33983-8|LNC|U1 small nuclear ribonucleoprotein Ab.IgG|U1 small nuclear ribonucleoprotein Ab.IgG
C1316447|T201|COMP|33984-6|LNC|Coagulation factor X activity actual/Normal|Coagulation factor X activity actual/Normal
C1316448|T201|COMP|33985-3|LNC|Bartonella henselae DNA|Bartonella henselae DNA
C1316449|T201|COMP|33986-1|LNC|Bartonella henselae DNA|Bartonella henselae DNA
C1316450|T201|COMP|33987-9|LNC|Heparin cofactor II actual/Normal|Heparin cofactor II actual/Normal
C1316451|T201|COMP|33988-7|LNC|Thymidine phosphorylase|Thymidine phosphorylase
C1316452|T201|COMP|33989-5|LNC|quiNINE induced platelet Ab|quiNINE induced platelet Ab
C1316453|T201|COMP|33990-3|LNC|Normoblasts/100 leukocytes|Normoblasts/100 leukocytes
C1316454|T201|COMP|33991-1|LNC|Cells.CD79b/100 cells|Cells.CD79b/100 cells
C1316516|T201|COMP|34053-9|LNC|Xylose^2H post 5 g xylose PO|Xylose^2H post 5 g xylose PO
C1316517|T201|COMP|34054-7|LNC|Thyrotropin^pre or post dose TRH|Thyrotropin^pre or post dose TRH
C1316518|T201|COMP|34055-4|LNC|Lutropin^pre or post XXX challenge|Lutropin^pre or post XXX challenge
C1316519|T201|COMP|34056-2|LNC|Glucose^pre or post dose arginine|Glucose^pre or post dose arginine
C1316520|T201|COMP|34057-0|LNC|Glucose^pre or post dose cloNIDine|Glucose^pre or post dose cloNIDine
C1316521|T201|COMP|34058-8|LNC|Glucose^pre or post dose glucagon|Glucose^pre or post dose glucagon
C1316522|T201|COMP|34059-6|LNC|Glucose^pre or post dose glucose|Glucose^pre or post dose glucose
C1316523|T201|COMP|34060-4|LNC|Glucose^pre or post dose insulin|Glucose^pre or post dose insulin
C1316524|T201|COMP|34061-2|LNC|Somatotropin^pre or post dose arginine|Somatotropin^pre or post dose arginine
C1316525|T201|COMP|34062-0|LNC|Somatotropin^pre or post dose cloNIDine|Somatotropin^pre or post dose cloNIDine
C1316526|T201|COMP|34063-8|LNC|Somatotropin^pre or post dose glucagon|Somatotropin^pre or post dose glucagon
C1316527|T201|COMP|34064-6|LNC|Somatotropin^pre or post dose insulin|Somatotropin^pre or post dose insulin
C1316528|T201|COMP|34065-3|LNC|Cortisol^pre or post dose corticotropin|Cortisol^pre or post dose corticotropin
C1316585|T201|COMP|34122-2|LNC|Pathology procedure note|Pathology procedure note
C1316605|T201|COMP|34142-0|LNC|Paraneoplastic Ab|Paraneoplastic Ab
C1316606|T201|COMP|34143-8|LNC|HLA-DQ locus 2|HLA-DQ locus 2
C1316607|T201|COMP|34144-6|LNC|HLA-DR W locus 2|HLA-DR W locus 2
C1316608|T201|COMP|34145-3|LNC|Human antichimeric Ab|Human antichimeric Ab
C1316609|T201|COMP|34146-1|LNC|Neopterin|Neopterin
C1316610|T201|COMP|34147-9|LNC|Treponema pallidum Ab.IgG+IgM|Treponema pallidum Ab.IgG+IgM
C1316611|T201|COMP|34148-7|LNC|Borrelia burgdorferi Ab.IgG+IgM|Borrelia burgdorferi Ab.IgG+IgM
C1316612|T201|COMP|34149-5|LNC|N-acetyl-L-aspartate|N-acetyl-L-aspartate
C1316613|T201|COMP|34150-3|LNC|Mycoplasma fermentans DNA|Mycoplasma fermentans DNA
C1316614|T201|COMP|34151-1|LNC|Cells.CD10+CD25+|Cells.CD10+CD25+
C1316615|T201|COMP|34152-9|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1316616|T201|COMP|34153-7|LNC|Influenza virus A Ab|Influenza virus A Ab
C1316617|T201|COMP|34154-5|LNC|Influenza virus B Ab|Influenza virus B Ab
C1316618|T201|COMP|34155-2|LNC|Guanidinoacetate/Creatinine|Guanidinoacetate/Creatinine
C1316619|T201|COMP|34156-0|LNC|Insulin.bound|Insulin.bound
C1316620|T201|COMP|34157-8|LNC|little e Ab|little e Ab
C1316621|T201|COMP|34158-6|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1316622|T201|COMP|34159-4|LNC|Tau protein|Tau protein
C1316623|T201|COMP|34160-2|LNC|Creatine kinase|Creatine kinase
C1316624|T201|COMP|34161-0|LNC|Cancer Ag 72-4|Cancer Ag 72-4
C1316625|T201|COMP|34162-8|LNC|Hepatitis C virus Ab.IgG band pattern|Hepatitis C virus Ab.IgG band pattern
C1316626|T201|COMP|34163-6|LNC|Oxygen content|Oxygen content
C1316627|T201|COMP|34164-4|LNC|N-Acetylglucosamine-6-Sulfatase|N-Acetylglucosamine-6-Sulfatase
C1316628|T201|COMP|34165-1|LNC|Granulocytes.immature|Granulocytes.immature
C1316630|T201|COMP|34167-7|LNC|Platelets.large|Platelets.large
C1316631|T201|COMP|34168-5|LNC|Sulfocysteine/Creatinine|Sulfocysteine/Creatinine
C1316632|T201|COMP|34169-3|LNC|Fatty acids.very long chain|Fatty acids.very long chain
C1316633|T201|COMP|34170-1|LNC|Biopterin|Biopterin
C1316634|T201|COMP|34171-9|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1316635|T201|COMP|34172-7|LNC|Streptococcus pneumoniae Danish serotype 6B Ab|Streptococcus pneumoniae Danish serotype 6B Ab
C1316636|T201|COMP|34173-5|LNC|Mixed cellular casts|Mixed cellular casts
C1316637|T201|COMP|34174-3|LNC|Hemoglobin casts|Hemoglobin casts
C1316638|T201|COMP|34175-0|LNC|Analgesics|Analgesics
C1316639|T201|COMP|34176-8|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C1316640|T201|COMP|34177-6|LNC|Opiates|Opiates
C1316641|T201|COMP|34178-4|LNC|Phenothiazines|Phenothiazines
C1316642|T201|COMP|34179-2|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C1316643|T201|COMP|34180-0|LNC|Ethanol|Ethanol
C1316644|T201|COMP|34181-8|LNC|Methanol|Methanol
C1316645|T201|COMP|34182-6|LNC|Methaqualone metabolite|Methaqualone metabolite
C1316646|T201|COMP|34183-4|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C1316647|T201|COMP|34184-2|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C1316648|T201|COMP|34185-9|LNC|methIMAzole|methIMAzole
C1316649|T201|COMP|34186-7|LNC|Para aminobenzoate|Para aminobenzoate
C1316650|T201|COMP|34187-5|LNC|DNA double strand Ab|DNA double strand Ab
C1316651|T201|COMP|34188-3|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C1316653|T201|COMP|34190-9|LNC|Thermoactinomyces vulgaris Ab.IgG|Thermoactinomyces vulgaris Ab.IgG
C1316654|T201|COMP|34191-7|LNC|Beta glucuronidase|Beta glucuronidase
C1316655|T201|COMP|34192-5|LNC|Beta galactosidase|Beta galactosidase
C1316656|T201|COMP|34193-3|LNC|SMPD1 gene mutations tested for|SMPD1 gene mutations tested for
C1316657|T201|COMP|34194-1|LNC|Fructose|Fructose
C1316658|T201|COMP|34195-8|LNC|little e Ab|little e Ab
C1316659|T201|COMP|34196-6|LNC|C Ab|C Ab
C1316660|T201|COMP|34197-4|LNC|Salicylamide^trough|Salicylamide^trough
C1316661|T201|COMP|34198-2|LNC|Salicylamide^peak|Salicylamide^peak
C1316662|T201|COMP|34199-0|LNC|Neutrophils.hypersegmented|Neutrophils.hypersegmented
C1316663|T201|COMP|34200-6|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C1316664|T201|COMP|34201-4|LNC|Cytomegalovirus|Cytomegalovirus
C1316665|T201|COMP|34202-2|LNC|Linezolid|Linezolid
C1316666|T201|COMP|34203-0|LNC|SCA12 gene.CAG repeats|SCA12 gene.CAG repeats
C1316667|T201|COMP|34204-8|LNC|11-Deoxycortisol|11-Deoxycortisol
C1316668|T201|COMP|34205-5|LNC|11-Deoxycortisol|11-Deoxycortisol
C1316669|T201|COMP|34206-3|LNC|11-Deoxycortisol/Creatinine|11-Deoxycortisol/Creatinine
C1316670|T201|COMP|34207-1|LNC|11-Hydroxyandrosterone|11-Hydroxyandrosterone
C1316671|T201|COMP|34208-9|LNC|11-Hydroxyandrosterone|11-Hydroxyandrosterone
C1316672|T201|COMP|34209-7|LNC|11-Hydroxyandrosterone/Creatinine|11-Hydroxyandrosterone/Creatinine
C1316673|T201|COMP|34210-5|LNC|11-Hydroxyetiocholanolone|11-Hydroxyetiocholanolone
C1316674|T201|COMP|34211-3|LNC|11-Hydroxyetiocholanolone|11-Hydroxyetiocholanolone
C1316675|T201|COMP|34212-1|LNC|11-Hydroxyetiocholanolone/Creatinine|11-Hydroxyetiocholanolone/Creatinine
C1316676|T201|COMP|34213-9|LNC|11-Ketoandrosterone|11-Ketoandrosterone
C1316677|T201|COMP|34214-7|LNC|11-Ketoandrosterone|11-Ketoandrosterone
C1316678|T201|COMP|34215-4|LNC|11-Ketoandrosterone/Creatinine|11-Ketoandrosterone/Creatinine
C1316679|T201|COMP|34216-2|LNC|11-Ketoetiocholanolone|11-Ketoetiocholanolone
C1316680|T201|COMP|34217-0|LNC|11-Ketoetiocholanolone|11-Ketoetiocholanolone
C1316681|T201|COMP|34218-8|LNC|17-Hydroxycorticosteroids|17-Hydroxycorticosteroids
C1316682|T201|COMP|34219-6|LNC|17-Hydroxycorticosteroids/Creatinine|17-Hydroxycorticosteroids/Creatinine
C1316683|T201|COMP|34220-4|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C1316684|T201|COMP|34221-2|LNC|17-Hydroxyprogesterone/Creatinine|17-Hydroxyprogesterone/Creatinine
C1316685|T201|COMP|34222-0|LNC|17-Ketosteroids|17-Ketosteroids
C1316686|T201|COMP|34223-8|LNC|17-Ketosteroids/Creatinine|17-Ketosteroids/Creatinine
C1316687|T201|COMP|34224-6|LNC|3-Alpha-Androstanediol glucuronide|3-Alpha-Androstanediol glucuronide
C1316688|T201|COMP|34225-3|LNC|3-Alpha-Androstanediol glucuronide|3-Alpha-Androstanediol glucuronide
C1316689|T201|COMP|34226-1|LNC|3-Alpha-Androstanediol glucuronide/Creatinine|3-Alpha-Androstanediol glucuronide/Creatinine
C1316690|T201|COMP|34227-9|LNC|Acylcarnitine|Acylcarnitine
C1316691|T201|COMP|34228-7|LNC|Acylcarnitine|Acylcarnitine
C1316692|T201|COMP|34229-5|LNC|Acylcarnitine/Creatinine|Acylcarnitine/Creatinine
C1316693|T201|COMP|34230-3|LNC|Adenosine monophosphate.cyclic|Adenosine monophosphate.cyclic
C1316694|T201|COMP|34231-1|LNC|Aldosterone/Creatinine|Aldosterone/Creatinine
C1316695|T201|COMP|34232-9|LNC|Pseudallescheria boydii Ab.IgG|Pseudallescheria boydii Ab.IgG
C1316696|T201|COMP|34233-7|LNC|Alternaria sp Ab.IgG|Alternaria sp Ab.IgG
C1316697|T201|COMP|34234-5|LNC|Ampicillin Ab.IgG|Ampicillin Ab.IgG
C1316698|T201|COMP|34235-2|LNC|Amylase/Creatinine|Amylase/Creatinine
C1316699|T201|COMP|34236-0|LNC|Androstenediol|Androstenediol
C1316700|T201|COMP|34237-8|LNC|Androstenediol|Androstenediol
C1316701|T201|COMP|34238-6|LNC|Androstenediol/Creatinine|Androstenediol/Creatinine
C1316702|T201|COMP|34239-4|LNC|Androstenedione|Androstenedione
C1316703|T201|COMP|34240-2|LNC|Androstenedione/Creatinine|Androstenedione/Creatinine
C1316704|T201|COMP|34241-0|LNC|Androsterone|Androsterone
C1316705|T201|COMP|34242-8|LNC|Androsterone|Androsterone
C1316706|T201|COMP|34243-6|LNC|Androsterone/Creatinine|Androsterone/Creatinine
C1316707|T201|COMP|34244-4|LNC|Arsenic|Arsenic
C1316708|T201|COMP|34245-1|LNC|Arsenic|Arsenic
C1316709|T201|COMP|34246-9|LNC|Ascorbate|Ascorbate
C1316710|T201|COMP|34247-7|LNC|Ascorbate|Ascorbate
C1316711|T201|COMP|34248-5|LNC|Ascorbate/Creatinine|Ascorbate/Creatinine
C1316712|T201|COMP|34249-3|LNC|Asialoganglioside GM2 Ab|Asialoganglioside GM2 Ab
C1316713|T201|COMP|34250-1|LNC|Betula verrucosa recombinant (rBet v) 4 Ab.IgE|Betula verrucosa recombinant (rBet v) 4 Ab.IgE
C1316714|T201|COMP|34251-9|LNC|Borrelia garinii Ab.IgG|Borrelia garinii Ab.IgG
C1316715|T201|COMP|34252-7|LNC|Borrelia garinii Ab.IgM|Borrelia garinii Ab.IgM
C1316716|T201|COMP|34253-5|LNC|C peptide|C peptide
C1316717|T201|COMP|34254-3|LNC|Cadmium|Cadmium
C1316718|T201|COMP|34255-0|LNC|Cadmium|Cadmium
C1316719|T201|COMP|34256-8|LNC|Cancer Ag 50|Cancer Ag 50
C1316720|T201|COMP|34257-6|LNC|Carnitine|Carnitine
C1316721|T201|COMP|34258-4|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C1316722|T201|COMP|34259-2|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C1316723|T201|COMP|34260-0|LNC|Catecholamines|Catecholamines
C1316724|T201|COMP|34261-8|LNC|Catecholamines|Catecholamines
C1316725|T201|COMP|34262-6|LNC|Catecholamines/Creatinine|Catecholamines/Creatinine
C1316726|T201|COMP|34263-4|LNC|Cefaclor Ab.IgG|Cefaclor Ab.IgG
C1316727|T201|COMP|34264-2|LNC|Chlamydia sp Ab.IgA|Chlamydia sp Ab.IgA
C1316728|T201|COMP|34265-9|LNC|Chloride/Creatinine|Chloride/Creatinine
C1316729|T201|COMP|34266-7|LNC|Citrate|Citrate
C1316730|T201|COMP|34267-5|LNC|Cladosporium sp Ab.IgG|Cladosporium sp Ab.IgG
C1316731|T201|COMP|34268-3|LNC|Cobalt|Cobalt
C1316732|T201|COMP|34269-1|LNC|Cobalt|Cobalt
C1316733|T201|COMP|34270-9|LNC|Cobalt/Creatinine|Cobalt/Creatinine
C1316734|T201|COMP|34271-7|LNC|Collagen crosslinked N-telopeptide|Collagen crosslinked N-telopeptide
C1316735|T201|COMP|34272-5|LNC|Collagen crosslinked N-telopeptide/Creatinine|Collagen crosslinked N-telopeptide/Creatinine
C1316736|T201|COMP|34273-3|LNC|Copper|Copper
C1316737|T201|COMP|34274-1|LNC|Creatine|Creatine
C1316738|T201|COMP|34275-8|LNC|Creatine/Creatinine|Creatine/Creatinine
C1316739|T201|COMP|34276-6|LNC|Cysteate|Cysteate
C1316740|T201|COMP|34277-4|LNC|Cysteine|Cysteine
C1316741|T201|COMP|34278-2|LNC|Cystine|Cystine
C1316742|T201|COMP|34279-0|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C1316743|T201|COMP|34280-8|LNC|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C1316744|T201|COMP|34281-6|LNC|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C1316745|T201|COMP|34282-4|LNC|Dehydroepiandrosterone sulfate/Creatinine|Dehydroepiandrosterone sulfate/Creatinine
C1316746|T201|COMP|34283-2|LNC|Dehydroepiandrosterone/Creatinine|Dehydroepiandrosterone/Creatinine
C1316747|T201|COMP|34284-0|LNC|Delta aminolevulinate|Delta aminolevulinate
C1316748|T201|COMP|34285-7|LNC|Ehrlichia sp Ab|Ehrlichia sp Ab
C1316749|T201|COMP|34286-5|LNC|Estradiol|Estradiol
C1316750|T201|COMP|34287-3|LNC|Estradiol|Estradiol
C1316751|T201|COMP|34288-1|LNC|Estradiol.unconjugated|Estradiol.unconjugated
C1316752|T201|COMP|34289-9|LNC|Estradiol.unconjugated|Estradiol.unconjugated
C1316753|T201|COMP|34290-7|LNC|Estradiol.unconjugated/Creatinine|Estradiol.unconjugated/Creatinine
C1316754|T201|COMP|34291-5|LNC|Estradiol/Creatinine|Estradiol/Creatinine
C1316755|T201|COMP|34292-3|LNC|Estriol|Estriol
C1316756|T201|COMP|34293-1|LNC|Estriol/Creatinine|Estriol/Creatinine
C1316757|T201|COMP|34294-9|LNC|Estrogen|Estrogen
C1316758|T201|COMP|34295-6|LNC|Estrogen|Estrogen
C1316759|T201|COMP|34296-4|LNC|Estrogen/Creatinine|Estrogen/Creatinine
C1316760|T201|COMP|34297-2|LNC|Estrone|Estrone
C1316761|T201|COMP|34298-0|LNC|Estrone|Estrone
C1316762|T201|COMP|34299-8|LNC|Estrone/Creatinine|Estrone/Creatinine
C1316763|T201|COMP|34300-4|LNC|Ethanolamine|Ethanolamine
C1316764|T201|COMP|34301-2|LNC|Etiocholanolone|Etiocholanolone
C1316765|T201|COMP|34302-0|LNC|Etiocholanolone|Etiocholanolone
C1316766|T201|COMP|34303-8|LNC|Etiocholanolone/Creatinine|Etiocholanolone/Creatinine
C1316767|T201|COMP|34304-6|LNC|Fluoride|Fluoride
C1316768|T201|COMP|34305-3|LNC|Flupenthixol|Flupenthixol
C1316769|T201|COMP|34306-1|LNC|Follitropin|Follitropin
C1316770|T201|COMP|34307-9|LNC|Fructose|Fructose
C1316771|T201|COMP|34308-7|LNC|Fructose|Fructose
C1316772|T201|COMP|34309-5|LNC|Fructose/Creatinine|Fructose/Creatinine
C1316773|T201|COMP|34310-3|LNC|Galactose|Galactose
C1316774|T201|COMP|34311-1|LNC|Galactose|Galactose
C1316775|T201|COMP|34312-9|LNC|Glucose/Creatinine|Glucose/Creatinine
C1316776|T201|COMP|34313-7|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C1316777|T201|COMP|34314-5|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C1316778|T201|COMP|34315-2|LNC|Hexacarboxylporphyrins|Hexacarboxylporphyrins
C1316779|T201|COMP|34316-0|LNC|Histamine|Histamine
C1316780|T201|COMP|34317-8|LNC|Histamine|Histamine
C1316781|T201|COMP|34318-6|LNC|HTLV I+II Ab|HTLV I+II Ab
C1316782|T201|COMP|34319-4|LNC|Inhibin B|Inhibin B
C1316783|T201|COMP|34320-2|LNC|Iodine|Iodine
C1316784|T201|COMP|34321-0|LNC|Iodine/Creatinine|Iodine/Creatinine
C1316785|T201|COMP|34322-8|LNC|Iron/Creatinine|Iron/Creatinine
C1316786|T201|COMP|34323-6|LNC|Lactate|Lactate
C1316787|T201|COMP|34324-4|LNC|Lactate|Lactate
C1316788|T201|COMP|34325-1|LNC|Lead|Lead
C1316789|T201|COMP|34326-9|LNC|Lead/Creatinine|Lead/Creatinine
C1316790|T201|COMP|34327-7|LNC|Lead/Creatinine|Lead/Creatinine
C1316791|T201|COMP|34328-5|LNC|Levodopa|Levodopa
C1316793|T201|COMP|34330-1|LNC|Lithium|Lithium
C1316794|T201|COMP|34331-9|LNC|Lithium/Creatinine|Lithium/Creatinine
C1316795|T201|COMP|34332-7|LNC|Lormetazepam|Lormetazepam
C1316796|T201|COMP|34333-5|LNC|Lutropin|Lutropin
C1316797|T201|COMP|34334-3|LNC|Lutropin/Creatinine|Lutropin/Creatinine
C1316798|T201|COMP|34335-0|LNC|Lysozyme|Lysozyme
C1316799|T201|COMP|34336-8|LNC|Lysozyme/Creatinine|Lysozyme/Creatinine
C1316800|T201|COMP|34337-6|LNC|Mercury|Mercury
C1316801|T201|COMP|34338-4|LNC|Mercury|Mercury
C1316802|T201|COMP|34340-0|LNC|Methionine sulfoxide|Methionine sulfoxide
C1316803|T201|COMP|34341-8|LNC|Mianserin+Normianserin|Mianserin+Normianserin
C1316804|T201|COMP|34342-6|LNC|Niacin|Niacin
C1316805|T201|COMP|34343-4|LNC|Nickel|Nickel
C1316806|T201|COMP|34344-2|LNC|N-methylhistamine|N-methylhistamine
C1316807|T201|COMP|34345-9|LNC|N-methylhistamine|N-methylhistamine
C1316808|T201|COMP|34346-7|LNC|N-methylhistamine/Creatinine|N-methylhistamine/Creatinine
C1316809|T201|COMP|34347-5|LNC|Normetanephrine|Normetanephrine
C1316810|T201|COMP|34348-3|LNC|Normetanephrine/Creatinine|Normetanephrine/Creatinine
C1316811|T201|COMP|34349-1|LNC|Oxalate|Oxalate
C1316812|T201|COMP|34350-9|LNC|Oxalate/Creatinine|Oxalate/Creatinine
C1316813|T201|COMP|34351-7|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C1316814|T201|COMP|34352-5|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C1316815|T201|COMP|34353-3|LNC|Pentacarboxylporphyrins/Creatinine|Pentacarboxylporphyrins/Creatinine
C1316816|T201|COMP|34354-1|LNC|Phosphate/Creatinine|Phosphate/Creatinine
C1316817|T201|COMP|34355-8|LNC|Phosphoethanolamine|Phosphoethanolamine
C1316818|T201|COMP|34356-6|LNC|Porphobilinogen|Porphobilinogen
C1316819|T201|COMP|34357-4|LNC|Porphobilinogen/Creatinine|Porphobilinogen/Creatinine
C1316820|T201|COMP|34358-2|LNC|Pregnanediol|Pregnanediol
C1316821|T201|COMP|34359-0|LNC|Pregnanediol/Creatinine|Pregnanediol/Creatinine
C1316822|T201|COMP|34360-8|LNC|Pregnanetriol|Pregnanetriol
C1316823|T201|COMP|34361-6|LNC|Pregnanetriol/Creatinine|Pregnanetriol/Creatinine
C1316824|T201|COMP|34362-4|LNC|Pregnanetriolone|Pregnanetriolone
C1316825|T201|COMP|34363-2|LNC|Pregnanetriolone|Pregnanetriolone
C1316826|T201|COMP|34364-0|LNC|Pregnanetriolone/Creatinine|Pregnanetriolone/Creatinine
C1316827|T201|COMP|34365-7|LNC|Primidone+PHENobarbital|Primidone+PHENobarbital
C1316828|T201|COMP|34366-5|LNC|Protein/Creatinine|Protein/Creatinine
C1316829|T201|COMP|34367-3|LNC|Pyridinoline|Pyridinoline
C1316830|T201|COMP|34368-1|LNC|Pyridinoline|Pyridinoline
C1316831|T201|COMP|34369-9|LNC|Salmonella paratyphi C H Ab|Salmonella paratyphi C H Ab
C1316832|T201|COMP|34370-7|LNC|Salmonella paratyphi C O Ab|Salmonella paratyphi C O Ab
C1316833|T201|COMP|34371-5|LNC|Salmonella typhi H Ab|Salmonella typhi H Ab
C1316834|T201|COMP|34372-3|LNC|Salmonella typhi O Ab|Salmonella typhi O Ab
C1316835|T201|COMP|34373-1|LNC|Serotonin|Serotonin
C1316836|T201|COMP|34374-9|LNC|Serotonin/Creatinine|Serotonin/Creatinine
C1316837|T201|COMP|34375-6|LNC|Streptokinase Ab|Streptokinase Ab
C1316838|T201|COMP|34376-4|LNC|Strongyloides sp Ab.IgG|Strongyloides sp Ab.IgG
C1316839|T201|COMP|34377-2|LNC|Sulthiame|Sulthiame
C1316840|T201|COMP|34378-0|LNC|Teicoplanin^peak|Teicoplanin^peak
C1316841|T201|COMP|34379-8|LNC|Teicoplanin^trough|Teicoplanin^trough
C1316842|T201|COMP|34380-6|LNC|Testosterone/Creatinine|Testosterone/Creatinine
C1316843|T201|COMP|34381-4|LNC|Thioguanine|Thioguanine
C1316844|T201|COMP|34382-2|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1316845|T201|COMP|34383-0|LNC|Trypanosoma brucei Ab|Trypanosoma brucei Ab
C1316846|T201|COMP|34384-8|LNC|Tryptophan|Tryptophan
C1316847|T201|COMP|34385-5|LNC|Urate/Creatinine|Urate/Creatinine
C1316848|T201|COMP|34386-3|LNC|Venlafaxine|Venlafaxine
C1316849|T201|COMP|34387-1|LNC|Zinc|Zinc
C1316850|T201|COMP|34388-9|LNC|Zinc|Zinc
C1316851|T201|COMP|34389-7|LNC|Zinc/Creatinine|Zinc/Creatinine
C1316858|T201|COMP|34396-2|LNC|11-Ketoetiocholanolone/Creatinine|11-Ketoetiocholanolone/Creatinine
C1316859|T201|COMP|34397-0|LNC|Amilsulpride|Amilsulpride
C1316860|T201|COMP|34398-8|LNC|Biotin|Biotin
C1316861|T201|COMP|34399-6|LNC|Buccal mucosa Ab|Buccal mucosa Ab
C1316862|T201|COMP|34400-2|LNC|Colon Ab|Colon Ab
C1316863|T201|COMP|34401-0|LNC|Complement C3d|Complement C3d
C1316864|T201|COMP|34402-8|LNC|Coproporphyrin/Hemoglobin|Coproporphyrin/Hemoglobin
C1316865|T201|COMP|34403-6|LNC|Cytomegalovirus Ab avidity|Cytomegalovirus Ab avidity
C1316866|T201|COMP|34404-4|LNC|Cytoskeleton Ab|Cytoskeleton Ab
C1316867|T201|COMP|34405-1|LNC|Escitalopram|Escitalopram
C1316868|T201|COMP|34406-9|LNC|Exocrine pancreas Ab|Exocrine pancreas Ab
C1316869|T201|COMP|34407-7|LNC|Interleukin 1|Interleukin 1
C1316870|T201|COMP|34408-5|LNC|Interleukin 2 receptor.soluble|Interleukin 2 receptor.soluble
C1316871|T201|COMP|34409-3|LNC|Keratin Ab|Keratin Ab
C1316872|T201|COMP|34410-1|LNC|Saccharopolyspora rectivirgula Ab.IgG|Saccharopolyspora rectivirgula Ab.IgG
C1316873|T201|COMP|34411-9|LNC|Mitochondria M4 Ab|Mitochondria M4 Ab
C1316874|T201|COMP|34412-7|LNC|Mitochondria M9 Ab|Mitochondria M9 Ab
C1316875|T201|COMP|34413-5|LNC|Moclobemide|Moclobemide
C1316876|T201|COMP|34414-3|LNC|Normianserin|Normianserin
C1316877|T201|COMP|34415-0|LNC|Normirtazapine|Normirtazapine
C1316878|T201|COMP|34416-8|LNC|Nucleosome Ab|Nucleosome Ab
C1316879|T201|COMP|34417-6|LNC|Protoporphyrin.zinc|Protoporphyrin.zinc
C1316880|T201|COMP|34418-4|LNC|Protoporphyrin|Protoporphyrin
C1316881|T201|COMP|34419-2|LNC|Reticulocytes.mature/Reticulocytes.total|Reticulocytes.mature/Reticulocytes.total
C1316882|T201|COMP|34420-0|LNC|Reticulocytes.mid/Reticulocytes.total|Reticulocytes.mid/Reticulocytes.total
C1316883|T201|COMP|34421-8|LNC|Rubella virus Ab.IgG avidity|Rubella virus Ab.IgG avidity
C1316884|T201|COMP|34422-6|LNC|Toxoplasma gondii Ab.IgG avidity|Toxoplasma gondii Ab.IgG avidity
C1316885|T201|COMP|34423-4|LNC|Salmonella enteritidis H Ab|Salmonella enteritidis H Ab
C1316886|T201|COMP|34424-2|LNC|Salmonella typhimurium H Ab|Salmonella typhimurium H Ab
C1316887|T201|COMP|34425-9|LNC|Betula verrucosa recombinant (rBet v) 1+2 Ab.IgE|Betula verrucosa recombinant (rBet v) 1+2 Ab.IgE
C1316888|T201|COMP|34426-7|LNC|cycloSPORINE.monoclonal|cycloSPORINE.monoclonal
C1316889|T201|COMP|34427-5|LNC|Methadone.R|Methadone.R
C1316890|T201|COMP|34428-3|LNC|Phleum pratense recombinant (rPhl p) 12 Ab.IgE|Phleum pratense recombinant (rPhl p) 12 Ab.IgE
C1316891|T201|COMP|34429-1|LNC|Phleum pratense recombinant (rPhl p) 1+5b Ab.IgE|Phleum pratense recombinant (rPhl p) 1+5b Ab.IgE
C1316892|T201|COMP|34430-9|LNC|Phleum pratense recombinant (rPhl p) 7+12 Ab.IgE|Phleum pratense recombinant (rPhl p) 7+12 Ab.IgE
C1316893|T201|COMP|34431-7|LNC|Salmonella enteritidis H Ab|Salmonella enteritidis H Ab
C1316894|T201|COMP|34432-5|LNC|Salmonella typhimurium H Ab|Salmonella typhimurium H Ab
C1316895|T201|COMP|34433-3|LNC|Bartonella henselae Ab|Bartonella henselae Ab
C1316896|T201|COMP|34434-1|LNC|Lutropin/Follitropin|Lutropin/Follitropin
C1316897|T201|COMP|34435-8|LNC|Protein pattern|Protein pattern
C1316898|T201|COMP|34436-6|LNC|Diethylene glycol|Diethylene glycol
C1316899|T201|COMP|34437-4|LNC|Coxsackievirus B Ab|Coxsackievirus B Ab
C1316900|T201|COMP|34438-2|LNC|Apolipoprotein E phenotyping|Apolipoprotein E phenotyping
C1316901|T201|COMP|34439-0|LNC|Natural killer cell function|Natural killer cell function
C1316902|T201|COMP|34440-8|LNC|Interpretation|Interpretation
C1316903|T201|COMP|34441-6|LNC|Spermatozoa|Spermatozoa
C1316904|T201|COMP|34442-4|LNC|Bilirubin.glucuronidated/Bilirubin.total|Bilirubin.glucuronidated/Bilirubin.total
C1316905|T201|COMP|34443-2|LNC|ZOLMitriptan|ZOLMitriptan
C1316906|T201|COMP|34444-0|LNC|Acarboxyprothrombin|Acarboxyprothrombin
C1316907|T201|COMP|34445-7|LNC|Leukocytes|Leukocytes
C1316908|T201|COMP|34446-5|LNC|Erythrocytes|Erythrocytes
C1316909|T201|COMP|34447-3|LNC|Cache valley virus RNA|Cache valley virus RNA
C1316910|T201|COMP|34448-1|LNC|Cache valley virus RNA|Cache valley virus RNA
C1316911|T201|COMP|34449-9|LNC|Eastern equine encephalitis virus RNA|Eastern equine encephalitis virus RNA
C1316912|T201|COMP|34450-7|LNC|Eastern equine encephalitis virus RNA|Eastern equine encephalitis virus RNA
C1316913|T201|COMP|34451-5|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C1316914|T201|COMP|34452-3|LNC|Jamestown canyon virus RNA|Jamestown canyon virus RNA
C1316915|T201|COMP|34453-1|LNC|Jamestown canyon virus RNA|Jamestown canyon virus RNA
C1316916|T201|COMP|34454-9|LNC|La Crosse virus RNA|La Crosse virus RNA
C1316917|T201|COMP|34455-6|LNC|La Crosse virus RNA|La Crosse virus RNA
C1316918|T201|COMP|34456-4|LNC|Powassan virus RNA|Powassan virus RNA
C1316919|T201|COMP|34457-2|LNC|Powassan virus RNA|Powassan virus RNA
C1316920|T201|COMP|34458-0|LNC|Saint Louis encephalitis virus RNA|Saint Louis encephalitis virus RNA
C1316921|T201|COMP|34459-8|LNC|Saint Louis encephalitis virus RNA|Saint Louis encephalitis virus RNA
C1316922|T201|COMP|34460-6|LNC|West Nile virus RNA|West Nile virus RNA
C1316923|T201|COMP|34461-4|LNC|West Nile virus RNA|West Nile virus RNA
C1316924|T201|COMP|34462-2|LNC|California serogroup virus RNA|California serogroup virus RNA
C1316925|T201|COMP|34463-0|LNC|California serogroup virus RNA|California serogroup virus RNA
C1316926|T201|COMP|34464-8|LNC|B Ab|B Ab
C1316927|T201|COMP|34465-5|LNC|B Ab|B Ab
C1316928|T201|COMP|34466-3|LNC|Carbohydrates|Carbohydrates
C1316929|T201|COMP|34467-1|LNC|Cholesterol.in chylomicrons|Cholesterol.in chylomicrons
C1316930|T201|COMP|34468-9|LNC|Clostridioides difficile toxin A+B|Clostridioides difficile toxin A+B
C1316931|T201|COMP|34469-7|LNC|Leukocytes|Leukocytes
C1316932|T201|COMP|34470-5|LNC|Giardia lamblia Ag|Giardia lamblia Ag
C1316933|T201|COMP|34471-3|LNC|Calcium bilirubinate crystals|Calcium bilirubinate crystals
C1316934|T201|COMP|34472-1|LNC|Cholesterol crystals|Cholesterol crystals
C1316935|T201|COMP|34473-9|LNC|Neutrophils.vacuolated+Segmented|Neutrophils.vacuolated+Segmented
C1316936|T201|COMP|34474-7|LNC|ABO & Rh group|ABO & Rh group
C1316937|T201|COMP|34475-4|LNC|Cells.CD4+CD45RO+|Cells.CD4+CD45RO+
C1316938|T201|COMP|34476-2|LNC|Cortisol^1H post 250 ug corticotropin|Cortisol^1H post 250 ug corticotropin
C1316939|T201|COMP|34477-0|LNC|Blood group antibodies identified|Blood group antibodies identified
C1316940|T201|COMP|34478-8|LNC|Blood group antibodies identified|Blood group antibodies identified
C1316941|T201|COMP|34479-6|LNC|Blood group antibodies identified|Blood group antibodies identified
C1316942|T201|COMP|34480-4|LNC|Blood group antibodies identified|Blood group antibodies identified
C1316943|T201|COMP|34481-2|LNC|Blood group antibodies identified|Blood group antibodies identified
C1316944|T201|COMP|34482-0|LNC|Blood group antibodies identified|Blood group antibodies identified
C1316947|T201|COMP|34485-3|LNC|Avian paramyxovirus 1.exotic RNA|Avian paramyxovirus 1.exotic RNA
C1316948|T201|COMP|34486-1|LNC|Avian paramyxovirus 1 RNA|Avian paramyxovirus 1 RNA
C1316949|T201|COMP|34487-9|LNC|Influenza virus A RNA|Influenza virus A RNA
C1316950|T201|COMP|34488-7|LNC|Avian paramyxovirus 1 subtype|Avian paramyxovirus 1 subtype
C1316951|T201|COMP|34489-5|LNC|TOR1A gene deletion|TOR1A gene deletion
C1316952|T201|COMP|34490-3|LNC|MT-TK gene targeted mutation analysis|MT-TK gene targeted mutation analysis
C1316953|T201|COMP|34491-1|LNC|PRF1 gene targeted mutation analysis|PRF1 gene targeted mutation analysis
C1316954|T201|COMP|34492-9|LNC|NOTCH3 gene targeted mutation analysis|NOTCH3 gene targeted mutation analysis
C1316955|T201|COMP|34493-7|LNC|PRF1 gene targeted mutation analysis|PRF1 gene targeted mutation analysis
C1316956|T201|COMP|34494-5|LNC|SCA10 gene.ATTCT repeats|SCA10 gene.ATTCT repeats
C1316957|T201|COMP|34495-2|LNC|TOR1A gene targeted mutation analysis|TOR1A gene targeted mutation analysis
C1316958|T201|COMP|34496-0|LNC|Chromosome 7 uniparental disomy|Chromosome 7 uniparental disomy
C1316959|T201|COMP|34497-8|LNC|SPINK1 gene targeted mutation analysis|SPINK1 gene targeted mutation analysis
C1316960|T201|COMP|34498-6|LNC|ACADS gene targeted mutation analysis|ACADS gene targeted mutation analysis
C1316961|T201|COMP|34499-4|LNC|GPC3 gene targeted mutation analysis|GPC3 gene targeted mutation analysis
C1316962|T201|COMP|34500-9|LNC|SHOX gene targeted mutation analysis|SHOX gene targeted mutation analysis
C1316963|T201|COMP|34501-7|LNC|HADHA gene.c.1528G>C|HADHA gene.c.1528G>C
C1316964|T201|COMP|34502-5|LNC|VHL gene targeted mutation analysis|VHL gene targeted mutation analysis
C1316965|T201|COMP|34503-3|LNC|Chromosome 15 uniparental disomy|Chromosome 15 uniparental disomy
C1316966|T201|COMP|34504-1|LNC|GJB6 gene targeted mutation analysis|GJB6 gene targeted mutation analysis
C1316967|T201|COMP|34505-8|LNC|NPDC gene targeted mutation analysis|NPDC gene targeted mutation analysis
C1316969|T201|COMP|34507-4|LNC|PRX gene targeted mutation analysis|PRX gene targeted mutation analysis
C1316970|T201|COMP|34508-2|LNC|PANK2 gene targeted mutation analysis|PANK2 gene targeted mutation analysis
C1316971|T201|COMP|34509-0|LNC|UGT1A1 gene targeted mutation analysis|UGT1A1 gene targeted mutation analysis
C1316972|T201|COMP|34510-8|LNC|SDHB gene targeted mutation analysis|SDHB gene targeted mutation analysis
C1316973|T201|COMP|34511-6|LNC|SDHD gene targeted mutation analysis|SDHD gene targeted mutation analysis
C1316974|T201|COMP|34512-4|LNC|NPHS1 gene targeted mutation analysis|NPHS1 gene targeted mutation analysis
C1316975|T201|COMP|34513-2|LNC|NPHS1 gene targeted mutation analysis|NPHS1 gene targeted mutation analysis
C1316976|T201|COMP|34514-0|LNC|SLC22A18 gene targeted mutation analysis|SLC22A18 gene targeted mutation analysis
C1316977|T201|COMP|34515-7|LNC|GLA gene targeted mutation analysis|GLA gene targeted mutation analysis
C1316978|T201|COMP|34516-5|LNC|SPAST gene targeted mutation analysis|SPAST gene targeted mutation analysis
C1316979|T201|COMP|34517-3|LNC|CATCH22 syndrome gene targeted mutation analysis|CATCH22 syndrome gene targeted mutation analysis
C1316980|T201|COMP|34518-1|LNC|SMPD1 gene targeted mutation analysis|SMPD1 gene targeted mutation analysis
C1316981|T201|COMP|34519-9|LNC|HFE gene targeted mutation analysis|HFE gene targeted mutation analysis
C1316982|T201|COMP|34520-7|LNC|Carbon dioxide|Carbon dioxide
C1316983|T201|COMP|34521-5|LNC|Carnitine acyltransferase|Carnitine acyltransferase
C1316984|T201|COMP|34522-3|LNC|Phosphorylase kinase|Phosphorylase kinase
C1316985|T201|COMP|34523-1|LNC|Succinate semialdehyde dehydrogenase|Succinate semialdehyde dehydrogenase
C1316986|T201|COMP|34524-9|LNC|Neutrophils.band form|Neutrophils.band form
C1316987|T201|COMP|34525-6|LNC|Erythrocytes.lytic resistant|Erythrocytes.lytic resistant
C1316988|T201|COMP|34526-4|LNC|Sialooligosaccharides/Creatinine|Sialooligosaccharides/Creatinine
C1316990|T201|COMP|34528-0|LNC|PT panel|PT panel
C1316991|T201|COMP|34529-8|LNC|PT & aPTT panel|PT & aPTT panel
C1316992|T201|COMP|34530-6|LNC|ABO & Rh group panel|ABO & Rh group panel
C1316993|T201|COMP|34531-4|LNC|Blood type & Crossmatch panel|Blood type & Crossmatch panel
C1316994|T201|COMP|34532-2|LNC|Blood type & Indirect antibody screen panel|Blood type & Indirect antibody screen panel
C1316997|T201|COMP|34535-5|LNC|Microalbumin/Creatinine ratio panel|Microalbumin/Creatinine ratio panel
C1317001|T201|COMP|34539-7|LNC|Protein fractions panel|Protein fractions panel
C1317002|T201|COMP|34541-3|LNC|ACTH stimulation test using IM corticosteroids|ACTH stimulation test using IM corticosteroids
C1317003|T201|COMP|34542-1|LNC|ACTH stimulation test using IV corticosteroids|ACTH stimulation test using IV corticosteroids
C1317004|T201|COMP|34543-9|LNC|Bilirubin direct & total panel|Bilirubin direct & total panel
C1317005|T201|COMP|34544-7|LNC|Complement C3 & C4 panel|Complement C3 & C4 panel
C1317006|T201|COMP|34545-4|LNC|carBAMazepine free & total panel|carBAMazepine free & total panel
C1317007|T201|COMP|34546-2|LNC|Protein & Glucose panel|Protein & Glucose panel
C1317008|T201|COMP|34547-0|LNC|Complement profile panel|Complement profile panel
C1317009|T201|COMP|34548-8|LNC|Sodium & Potassium panel|Sodium & Potassium panel
C1317010|T201|COMP|34549-6|LNC|Follitropin & Lutropin panel|Follitropin & Lutropin panel
C1317011|T201|COMP|34550-4|LNC|Immunoglobulin panel|Immunoglobulin panel
C1317012|T201|COMP|34551-2|LNC|Catecholamines 3 panel|Catecholamines 3 panel
C1317015|T201|COMP|34554-6|LNC|Electrolytes 1998 & Venous pH panel|Electrolytes 1998 & Venous pH panel
C1317016|T201|COMP|34555-3|LNC|Creatinine renal clearance panel|Creatinine renal clearance panel
C1317017|T201|COMP|34556-1|LNC|Cell count panel|Cell count panel
C1317018|T201|COMP|34557-9|LNC|Cell count & Differential panel|Cell count & Differential panel
C1317019|T201|COMP|34558-7|LNC|Cell count panel|Cell count panel
C1317020|T201|COMP|34559-5|LNC|Cell count panel|Cell count panel
C1317021|T201|COMP|34560-3|LNC|Cell count & Differential panel|Cell count & Differential panel
C1317022|T201|COMP|34561-1|LNC|Cell count panel|Cell count panel
C1317023|T201|COMP|34562-9|LNC|Cell count & Differential panel|Cell count & Differential panel
C1317024|T201|COMP|34563-7|LNC|Cell count panel|Cell count panel
C1317025|T201|COMP|34564-5|LNC|Cell count & Differential panel|Cell count & Differential panel
C1317028|T201|COMP|34567-8|LNC|Cell count & Differential panel|Cell count & Differential panel
C1317029|T201|COMP|34568-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C1317032|T201|COMP|34571-0|LNC|Coagulation surface induced.lupus sensitive|Coagulation surface induced.lupus sensitive
C1317033|T201|COMP|34572-8|LNC|Coagulation surface induced.lupus sensitive|Coagulation surface induced.lupus sensitive
C1317036|T201|COMP|34575-1|LNC|8-Hydroxyloxapine|8-Hydroxyloxapine
C1317037|T201|COMP|34576-9|LNC|Adenovirus Ab|Adenovirus Ab
C1317038|T201|COMP|34577-7|LNC|Apheresis.therapeutic|Apheresis.therapeutic
C1317039|T201|COMP|34578-5|LNC|Barbiturates|Barbiturates
C1317040|T201|COMP|34579-3|LNC|Basophils|Basophils
C1317041|T201|COMP|34580-1|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C1317042|T201|COMP|34581-9|LNC|Calcium.ionized|Calcium.ionized
C1317043|T201|COMP|34582-7|LNC|Candida sp Ab.IgA|Candida sp Ab.IgA
C1317044|T201|COMP|34583-5|LNC|Candida sp Ab.IgG|Candida sp Ab.IgG
C1317045|T201|COMP|34584-3|LNC|Candida sp Ab.IgM|Candida sp Ab.IgM
C1317046|T201|COMP|34585-0|LNC|Inner Ear 68kD Ab|Inner Ear 68kD Ab
C1317047|T201|COMP|34586-8|LNC|JC virus DNA|JC virus DNA
C1317048|T201|COMP|34587-6|LNC|Palmitoyl protein thioesterase|Palmitoyl protein thioesterase
C1317049|T201|COMP|34588-4|LNC|Feeding duration|Feeding duration
C1317050|T201|COMP|34589-2|LNC|von Willebrand factor cleaving protease|von Willebrand factor cleaving protease
C1317051|T201|COMP|34590-0|LNC|von Willebrand factor cleaving protease inhibitor|von Willebrand factor cleaving protease inhibitor
C1318451|T201|COMP|10573-4|LNC|Ferning|Ferning
C1369461|T201|COMP|34591-8|LNC|HIV 1 Ab|HIV 1 Ab
C1369462|T201|COMP|34592-6|LNC|HIV 1 Ab|HIV 1 Ab
C1369463|T201|COMP|34593-4|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1369464|T201|COMP|34594-2|LNC|Schistosoma sp Ab|Schistosoma sp Ab
C1369465|T201|COMP|34595-9|LNC|Collection time|Collection time
C1369466|T201|COMP|34596-7|LNC|3-O-Methyldopa|3-O-Methyldopa
C1369467|T201|COMP|34597-5|LNC|Hepatitis D virus Ab.IgM|Hepatitis D virus Ab.IgM
C1369468|T201|COMP|34598-3|LNC|Sialate|Sialate
C1369469|T201|COMP|34599-1|LNC|Methotrexate|Methotrexate
C1369470|T201|COMP|34600-7|LNC|Immunoglobulin heavy chain gene rearrangements|Immunoglobulin heavy chain gene rearrangements
C1369471|T201|COMP|34601-5|LNC|Drugs identified|Drugs identified
C1369472|T201|COMP|34604-9|LNC|M Ab|M Ab
C1369473|T201|COMP|34605-6|LNC|Collagen type 2 Ab|Collagen type 2 Ab
C1369474|T201|COMP|34606-4|LNC|Minocycline|Minocycline
C1369475|T201|COMP|34607-2|LNC|Interferon.beta Ab|Interferon.beta Ab
C1369476|T201|COMP|34608-0|LNC|Leishmania sp Ab.IgG|Leishmania sp Ab.IgG
C1369477|T201|COMP|34609-8|LNC|Transketolase|Transketolase
C1369478|T201|COMP|34610-6|LNC|N-acetylaspartate/Creatinine|N-acetylaspartate/Creatinine
C1369479|T201|COMP|34611-4|LNC|Prostate specific Ag|Prostate specific Ag
C1369480|T201|COMP|34612-2|LNC|Iron|Iron
C1369481|T201|COMP|34613-0|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C1369482|T201|COMP|34614-8|LNC|Spermatozoa Ab.IgM|Spermatozoa Ab.IgM
C1369483|T201|COMP|34615-5|LNC|Iron.microscopic observation|Iron.microscopic observation
C1369484|T201|COMP|34616-3|LNC|Amino acids|Amino acids
C1369485|T201|COMP|34617-1|LNC|Antibiotic XXX|Antibiotic XXX
C1369486|T201|COMP|34618-9|LNC|Hemoglobin|Hemoglobin
C1369487|T201|COMP|34619-7|LNC|Complement C1 esterase inhibitor.functional|Complement C1 esterase inhibitor.functional
C1369488|T201|COMP|34620-5|LNC|Camphor|Camphor
C1369489|T201|COMP|34621-3|LNC|Liver cytosol Ab|Liver cytosol Ab
C1369490|T201|COMP|34622-1|LNC|Cells.CD4+CD25+/100 cells|Cells.CD4+CD25+/100 cells
C1369491|T201|COMP|34623-9|LNC|Colorado tick fever virus Ab|Colorado tick fever virus Ab
C1369492|T201|COMP|34624-7|LNC|Cystine.free|Cystine.free
C1369493|T201|COMP|34625-4|LNC|Corynebacterium diphtheriae toxin Ab|Corynebacterium diphtheriae toxin Ab
C1369494|T201|COMP|34626-2|LNC|2-Methylcitrate|2-Methylcitrate
C1369495|T201|COMP|34627-0|LNC|Methylmalonate|Methylmalonate
C1369496|T201|COMP|34628-8|LNC|Methotrexate|Methotrexate
C1369497|T201|COMP|34629-6|LNC|CISplatin|CISplatin
C1369498|T201|COMP|34630-4|LNC|Substance P|Substance P
C1369499|T201|COMP|34631-2|LNC|Cyproheptadine|Cyproheptadine
C1369500|T201|COMP|34632-0|LNC|hydrALAZINE|hydrALAZINE
C1369501|T201|COMP|34633-8|LNC|Hypoglycemics.sulfonyluric|Hypoglycemics.sulfonyluric
C1369502|T201|COMP|34634-6|LNC|Cells.CD11+CD18+|Cells.CD11+CD18+
C1369503|T201|COMP|34635-3|LNC|Citalopram|Citalopram
C1369504|T201|COMP|34636-1|LNC|Ciprofloxacin|Ciprofloxacin
C1369505|T201|COMP|34637-9|LNC|5-Methyltetrahydrofolate|5-Methyltetrahydrofolate
C1369506|T201|COMP|34638-7|LNC|Clarithromycin|Clarithromycin
C1369507|T201|COMP|34639-5|LNC|Epstein Barr virus capsid Ab.IgA|Epstein Barr virus capsid Ab.IgA
C1369508|T201|COMP|34640-3|LNC|Bile acid|Bile acid
C1369509|T201|COMP|34641-1|LNC|Protein pattern|Protein pattern
C1369510|T201|COMP|34642-9|LNC|Thyroid colloidal Ab|Thyroid colloidal Ab
C1369511|T201|COMP|34643-7|LNC|Lopinavir|Lopinavir
C1369512|T201|COMP|34644-5|LNC|Tenofovir|Tenofovir
C1369513|T201|COMP|34645-2|LNC|Chlamydophila pneumoniae DNA|Chlamydophila pneumoniae DNA
C1369514|T201|COMP|34646-0|LNC|Sulfatides|Sulfatides
C1369515|T201|COMP|34647-8|LNC|PPT1 gene targeted mutation analysis|PPT1 gene targeted mutation analysis
C1369516|T201|COMP|34648-6|LNC|Specimen weight|Specimen weight
C1369517|T201|COMP|34649-4|LNC|MERRF gene targeted mutation analysis|MERRF gene targeted mutation analysis
C1369518|T201|COMP|34650-2|LNC|TSC gene targeted mutation analysis|TSC gene targeted mutation analysis
C1369519|T201|COMP|34652-8|LNC|Pancreatic islet cell Ab|Pancreatic islet cell Ab
C1369520|T201|COMP|34653-6|LNC|GJB1 gene targeted mutation analysis|GJB1 gene targeted mutation analysis
C1369521|T201|COMP|34654-4|LNC|MPZ gene targeted mutation analysis|MPZ gene targeted mutation analysis
C1369522|T201|COMP|34655-1|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1369523|T201|COMP|34656-9|LNC|KEL gene targeted mutation analysis|KEL gene targeted mutation analysis
C1369524|T201|COMP|34658-5|LNC|MCOLN1 gene targeted mutation analysis|MCOLN1 gene targeted mutation analysis
C1369525|T201|COMP|34659-3|LNC|ATP7A gene targeted mutation analysis|ATP7A gene targeted mutation analysis
C1369526|T201|COMP|34660-1|LNC|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C1369527|T201|COMP|34661-9|LNC|Actin Ab.IgG|Actin Ab.IgG
C1369528|T201|COMP|34662-7|LNC|Mephenytoin+Normephenytoin|Mephenytoin+Normephenytoin
C1369529|T201|COMP|34663-5|LNC|Hemoglobin S|Hemoglobin S
C1369530|T201|COMP|34664-3|LNC|Clostridium botulinum toxin A Ab|Clostridium botulinum toxin A Ab
C1369531|T201|COMP|34665-0|LNC|TORCH panel|TORCH panel
C1369532|T201|COMP|34666-8|LNC|Carisoprodol+Meprobamate|Carisoprodol+Meprobamate
C1369533|T201|COMP|34667-6|LNC|Heavy metals panel|Heavy metals panel
C1369534|T201|COMP|34668-4|LNC|Prilocaine|Prilocaine
C1369535|T201|COMP|34669-2|LNC|Pyrimethamine|Pyrimethamine
C1369536|T201|COMP|34670-0|LNC|Choriogonadotropin|Choriogonadotropin
C1369537|T201|COMP|34671-8|LNC|8-Dehydrocholesterol|8-Dehydrocholesterol
C1369538|T201|COMP|34672-6|LNC|Immunoelectrophoresis panel|Immunoelectrophoresis panel
C1369539|T201|COMP|34673-4|LNC|Propofol|Propofol
C1369540|T201|COMP|34674-2|LNC|Tripeptide aminopeptidase|Tripeptide aminopeptidase
C1369541|T201|COMP|34675-9|LNC|Mitochondria DNA targeted mutation analysis|Mitochondria DNA targeted mutation analysis
C1369542|T201|COMP|34676-7|LNC|SMA@ gene mutation analysis|SMA@ gene mutation analysis
C1369543|T201|COMP|34677-5|LNC|Mitotic spindle apparatus Ab|Mitotic spindle apparatus Ab
C1369544|T201|COMP|34678-3|LNC|MT-RNR1 gene.m.1555A>G|MT-RNR1 gene.m.1555A>G
C1369545|T201|COMP|34679-1|LNC|PTPN11 gene targeted mutation analysis|PTPN11 gene targeted mutation analysis
C1369546|T201|COMP|34680-9|LNC|Ceramide trihexoside|Ceramide trihexoside
C1369547|T201|COMP|34681-7|LNC|Biopsy|Biopsy
C1369555|T201|COMP|34689-0|LNC|Sulfatidase|Sulfatidase
C1369556|T201|COMP|34690-8|LNC|CV2 Ab|CV2 Ab
C1369557|T201|COMP|34691-6|LNC|Erythroamino alcohol|Erythroamino alcohol
C1369558|T201|COMP|34692-4|LNC|Threoamino alcohol|Threoamino alcohol
C1369559|T201|COMP|34693-2|LNC|GALOP Ab|GALOP Ab
C1369560|T201|COMP|34694-0|LNC|Vascular endothelial growth factor|Vascular endothelial growth factor
C1369561|T201|COMP|34695-7|LNC|Cholesterol.in VLDL/Triglyceride|Cholesterol.in VLDL/Triglyceride
C1369562|T201|COMP|34696-5|LNC|Collection method|Collection method
C1369563|T201|COMP|34697-3|LNC|Alpha 1 antitrypsin actual/Normal|Alpha 1 antitrypsin actual/Normal
C1369564|T201|COMP|34698-1|LNC|CSTB gene targeted mutation analysis|CSTB gene targeted mutation analysis
C1369565|T201|COMP|34699-9|LNC|HIV 2 proviral DNA|HIV 2 proviral DNA
C1369567|T201|COMP|34701-3|LNC|Platelet factor 4 heparin complex induced Ab|Platelet factor 4 heparin complex induced Ab
C1369568|T201|COMP|34702-1|LNC|Mycoplasma sp|Mycoplasma sp
C1369569|T201|COMP|34703-9|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1369570|T201|COMP|34704-7|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1369572|T201|COMP|34706-2|LNC|CFTR gene.c.3199del6|CFTR gene.c.3199del6
C1369573|T201|COMP|34707-0|LNC|Chlamydophila pneumoniae rRNA|Chlamydophila pneumoniae rRNA
C1369574|T201|COMP|34708-8|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1369575|T201|COMP|34709-6|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1369576|T201|COMP|34710-4|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1369577|T201|COMP|34711-2|LNC|Cholinesterase|Cholinesterase
C1369578|T201|COMP|34712-0|LNC|Clostridioides difficile|Clostridioides difficile
C1369579|T201|COMP|34713-8|LNC|Clostridioides difficile toxin A+B|Clostridioides difficile toxin A+B
C1369580|T201|COMP|34714-6|LNC|Coagulation tissue factor induced.INR|Coagulation tissue factor induced.INR
C1369581|T201|COMP|34715-3|LNC|Cocaine|Cocaine
C1369582|T201|COMP|34716-1|LNC|Coxiella burnetii phase 1 Ab.IgG|Coxiella burnetii phase 1 Ab.IgG
C1369583|T201|COMP|34717-9|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C1369584|T201|COMP|34718-7|LNC|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C1369585|T201|COMP|34719-5|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1369586|T201|COMP|34720-3|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1369587|T201|COMP|34721-1|LNC|Dengue virus Ab.IgM|Dengue virus Ab.IgM
C1369588|T201|COMP|34506-6|LNC|EGR2 gene targeted mutation analysis|EGR2 gene targeted mutation analysis
C1369589|T201|COMP|34723-7|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C1369590|T201|COMP|34724-5|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C1369591|T201|COMP|34725-2|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C1369592|T201|COMP|34726-0|LNC|Eosinophils|Eosinophils
C1369593|T201|COMP|34727-8|LNC|DMPK gene targeted mutation analysis|DMPK gene targeted mutation analysis
C1369594|T201|COMP|34728-6|LNC|Carbon dioxide|Carbon dioxide
C1369595|T201|COMP|34729-4|LNC|CFTR gene.p.Arg117His+5T variant|CFTR gene.p.Arg117His+5T variant
C1369596|T201|COMP|34730-2|LNC|Chromosome breakage|Chromosome breakage
C1369597|T201|COMP|34731-0|LNC|APOE gene allele 1|APOE gene allele 1
C1369598|T201|COMP|34732-8|LNC|APOE gene allele 2|APOE gene allele 2
C1369599|T201|COMP|34733-6|LNC|APOE gene allele 3|APOE gene allele 3
C1369600|T201|COMP|34734-4|LNC|APOE gene gentoype|APOE gene gentoype
C1369601|T201|COMP|34735-1|LNC|APOE gene allele 4|APOE gene allele 4
C1369602|T201|COMP|34736-9|LNC|Calcium oxalate index|Calcium oxalate index
C1369603|T201|COMP|34737-7|LNC|Nuclear mitotic apparatus Ab|Nuclear mitotic apparatus Ab
C1369604|T201|COMP|34738-5|LNC|K Ab|K Ab
C1369605|T201|COMP|34739-3|LNC|NR0B1 gene targeted mutation analysis|NR0B1 gene targeted mutation analysis
C1369606|T201|COMP|34740-1|LNC|NEFL gene targeted mutation analysis|NEFL gene targeted mutation analysis
C1369607|T201|COMP|34741-9|LNC|RHCE gene targeted mutation analysis|RHCE gene targeted mutation analysis
C1369608|T201|COMP|34742-7|LNC|Chromosome breakage|Chromosome breakage
C1369609|T201|COMP|34743-5|LNC|Hemoglobin.stable|Hemoglobin.stable
C1369685|T201|COMP|34819-3|LNC|Note|Note
C1369748|T201|COMP|34882-1|LNC|Ethanol|Ethanol
C1369749|T201|COMP|34883-9|LNC|Mycoplasma sp Ag|Mycoplasma sp Ag
C1369750|T201|COMP|34884-7|LNC|Haemophilus paragallinarum Ab|Haemophilus paragallinarum Ab
C1369751|T201|COMP|34885-4|LNC|African horse sickness virus Ab|African horse sickness virus Ab
C1369752|T201|COMP|34886-2|LNC|Viral hemorrhagic disease virus Ab|Viral hemorrhagic disease virus Ab
C1369753|T201|COMP|34887-0|LNC|Peste des petits ruminants virus Ag|Peste des petits ruminants virus Ag
C1369754|T201|COMP|34888-8|LNC|Aino virus Ab|Aino virus Ab
C1369755|T201|COMP|34889-6|LNC|Akabane virus Ab|Akabane virus Ab
C1369756|T201|COMP|34890-4|LNC|Coliform bacteria|Coliform bacteria
C1369757|T201|COMP|34891-2|LNC|Salmonella enteritidis|Salmonella enteritidis
C1369758|T201|COMP|34892-0|LNC|West Nile virus RNA|West Nile virus RNA
C1369759|T201|COMP|34893-8|LNC|Aino virus Ab|Aino virus Ab
C1369760|T201|COMP|34894-6|LNC|Akabane virus Ab|Akabane virus Ab
C1369773|T201|COMP|34907-6|LNC|Calcium^^corrected for total protein|Calcium^^corrected for total protein
C1369774|T201|COMP|34908-4|LNC|Neopterin|Neopterin
C1369775|T201|COMP|34909-2|LNC|Cortisol.free|Cortisol.free
C1369776|T201|COMP|34910-0|LNC|Basophils.immature|Basophils.immature
C1369777|T201|COMP|34911-8|LNC|Basophils.immature/100 leukocytes|Basophils.immature/100 leukocytes
C1369778|T201|COMP|34912-6|LNC|Eosinophils.immature|Eosinophils.immature
C1369779|T201|COMP|34913-4|LNC|Eosinophils.immature/100 leukocytes|Eosinophils.immature/100 leukocytes
C1369780|T201|COMP|34914-2|LNC|Malignant cells|Malignant cells
C1369781|T201|COMP|34915-9|LNC|Malignant cells/100 leukocytes|Malignant cells/100 leukocytes
C1369782|T201|COMP|34916-7|LNC|Plasma cell precursor|Plasma cell precursor
C1369783|T201|COMP|34917-5|LNC|Plasma cell precursor/100 leukocytes|Plasma cell precursor/100 leukocytes
C1369784|T201|COMP|34918-3|LNC|Sezary cells|Sezary cells
C1369785|T201|COMP|34919-1|LNC|Sezary cells/100 leukocytes|Sezary cells/100 leukocytes
C1369786|T201|COMP|34920-9|LNC|Lymphocytes.immunoblastic/100 leukocytes|Lymphocytes.immunoblastic/100 leukocytes
C1369787|T201|COMP|34921-7|LNC|Lymphocytes.plasmacytoid/100 leukocytes|Lymphocytes.plasmacytoid/100 leukocytes
C1369788|T201|COMP|34922-5|LNC|Lymphoblasts/100 leukocytes|Lymphoblasts/100 leukocytes
C1369789|T201|COMP|34923-3|LNC|Monoblasts/100 leukocytes|Monoblasts/100 leukocytes
C1369790|T201|COMP|34924-1|LNC|Monocytes.immature|Monocytes.immature
C1369791|T201|COMP|34925-8|LNC|Monocytes.immature/100 leukocytes|Monocytes.immature/100 leukocytes
C1369792|T201|COMP|34927-4|LNC|Urobilinogen|Urobilinogen
C1369793|T201|COMP|34928-2|LNC|Urobilinogen|Urobilinogen
C1369794|T201|COMP|34929-0|LNC|Cells.CD3+CD4+CD45RO+CD45RA-/100 cells|Cells.CD3+CD4+CD45RO+CD45RA-/100 cells
C1369795|T201|COMP|34930-8|LNC|Cells.CD3+CD4+CD45RO+CD45RA+/100 cells|Cells.CD3+CD4+CD45RO+CD45RA+/100 cells
C1369796|T201|COMP|34931-6|LNC|Cells.CD3+CD4+CD45RO-CD45RA-/100 cells|Cells.CD3+CD4+CD45RO-CD45RA-/100 cells
C1369797|T201|COMP|34932-4|LNC|Cells.CD3+CD4+CD45RO-CD45RA+/100 cells|Cells.CD3+CD4+CD45RO-CD45RA+/100 cells
C1369798|T201|COMP|34933-2|LNC|Cells.CD3+CD8+CD45RO+CD45RA-/100 cells|Cells.CD3+CD8+CD45RO+CD45RA-/100 cells
C1369799|T201|COMP|34934-0|LNC|Cells.CD3+CD8+CD45RO+CD45RA+/100 cells|Cells.CD3+CD8+CD45RO+CD45RA+/100 cells
C1369800|T201|COMP|34935-7|LNC|Cells.CD3+CD8+CD45RO-CD45RA-/100 cells|Cells.CD3+CD8+CD45RO-CD45RA-/100 cells
C1369801|T201|COMP|34936-5|LNC|Cells.CD3+CD8+CD45RO-CD45RA+/100 cells|Cells.CD3+CD8+CD45RO-CD45RA+/100 cells
C1369802|T201|COMP|34937-3|LNC|Fibrinopeptide A|Fibrinopeptide A
C1369803|T201|COMP|34938-1|LNC|Phosphate|Phosphate
C1369804|T201|COMP|34939-9|LNC|Tumor necrosis factor.alpha|Tumor necrosis factor.alpha
C1369805|T201|COMP|34940-7|LNC|Babesia microti Ab.IgG & IgM panel|Babesia microti Ab.IgG & IgM panel
C1369806|T201|COMP|34941-5|LNC|Bordetella pertussis Ab.IgG & IgM panel|Bordetella pertussis Ab.IgG & IgM panel
C1369807|T201|COMP|34942-3|LNC|Borrelia burgdorferi Ab.IgG & IgM panel|Borrelia burgdorferi Ab.IgG & IgM panel
C1369808|T201|COMP|34943-1|LNC|Borrelia burgdorferi Ab.IgG & IgM panel|Borrelia burgdorferi Ab.IgG & IgM panel
C1369809|T201|COMP|34944-9|LNC|Cytomegalovirus Ab.IgG & IgM panel|Cytomegalovirus Ab.IgG & IgM panel
C1369810|T201|COMP|34945-6|LNC|Herpes virus 6 Ab.IgG & IgM panel|Herpes virus 6 Ab.IgG & IgM panel
C1369811|T201|COMP|34946-4|LNC|Herpes virus 6 Ab.IgG & IgM panel|Herpes virus 6 Ab.IgG & IgM panel
C1369812|T201|COMP|34947-2|LNC|Herpes virus 7 Ab.IgG & IgM panel|Herpes virus 7 Ab.IgG & IgM panel
C1369813|T201|COMP|34948-0|LNC|Measles virus Ab.IgG & IgM panel|Measles virus Ab.IgG & IgM panel
C1369814|T201|COMP|34949-8|LNC|Measles virus Ab.IgG & IgM panel|Measles virus Ab.IgG & IgM panel
C1369815|T201|COMP|34950-6|LNC|Parvovirus B19 Ab.IgG & IgM panel|Parvovirus B19 Ab.IgG & IgM panel
C1369816|T201|COMP|34951-4|LNC|Phosphatidylserine Ab.IgG & IgM panel|Phosphatidylserine Ab.IgG & IgM panel
C1369817|T201|COMP|34952-2|LNC|Rubella virus Ab.IgG & IgM panel|Rubella virus Ab.IgG & IgM panel
C1369818|T201|COMP|34953-0|LNC|Rubella virus Ab.IgG & IgM panel|Rubella virus Ab.IgG & IgM panel
C1369819|T201|COMP|34954-8|LNC|Treponema pallidum Ab.IgG & IgM panel|Treponema pallidum Ab.IgG & IgM panel
C1369821|T201|COMP|34956-3|LNC|Western equine encephalitis virus Ab.IgM|Western equine encephalitis virus Ab.IgM
C1369823|T201|COMP|34960-5|LNC|HLA Ab|HLA Ab
C1369824|T201|COMP|34961-3|LNC|Rh|Rh
C1369825|T201|COMP|34962-1|LNC|Cells.CD3+TCR alpha beta+/100 cells|Cells.CD3+TCR alpha beta+/100 cells
C1369826|T201|COMP|34963-9|LNC|Cells.CD3+TCR alpha beta+|Cells.CD3+TCR alpha beta+
C1369827|T201|COMP|34964-7|LNC|Osmotic fragility|Osmotic fragility
C1369829|T201|COMP|34966-2|LNC|Osmotic fragility^0.10% sodium chloride|Osmotic fragility^0.10% sodium chloride
C1369831|T201|COMP|34968-8|LNC|Osmotic fragility^0.20% sodium chloride|Osmotic fragility^0.20% sodium chloride
C1369832|T201|COMP|34969-6|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C1369833|T201|COMP|34970-4|LNC|Date ultrasound|Date ultrasound
C1369834|T201|COMP|34971-2|LNC|Neutrophil associated Ab|Neutrophil associated Ab
C1369835|T201|COMP|34972-0|LNC|DNA index 3|DNA index 3
C1369836|T201|COMP|34973-8|LNC|DNA index 2|DNA index 2
C1369837|T201|COMP|34974-6|LNC|DNA index 3|DNA index 3
C1369838|T201|COMP|34976-1|LNC|DNA index 2|DNA index 2
C1369839|T201|COMP|34977-9|LNC|Platelet genotype|Platelet genotype
C1369840|T201|COMP|34978-7|LNC|Specimen volume|Specimen volume
C1369841|T201|COMP|34979-5|LNC|Specimen volume|Specimen volume
C1369842|T201|COMP|34980-3|LNC|Specimen volume|Specimen volume
C1369843|T201|COMP|34981-1|LNC|Specimen volume|Specimen volume
C1369844|T201|COMP|34982-9|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C1369845|T201|COMP|34983-7|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C1369846|T201|COMP|34984-5|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C1369847|T201|COMP|34985-2|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C1369848|T201|COMP|34986-0|LNC|Unidentified cells|Unidentified cells
C1369849|T201|COMP|34988-6|LNC|Unidentified cells|Unidentified cells
C1369850|T201|COMP|34989-4|LNC|Unidentified cells|Unidentified cells
C1369851|T201|COMP|34990-2|LNC|Unidentified cells|Unidentified cells
C1369852|T201|COMP|34991-0|LNC|Unidentified cells|Unidentified cells
C1369853|T201|COMP|34992-8|LNC|Smudge cells/100 leukocytes|Smudge cells/100 leukocytes
C1369854|T201|COMP|34993-6|LNC|Smudge cells|Smudge cells
C1369855|T201|COMP|34994-4|LNC|Smear morphology panel|Smear morphology panel
C1369856|T201|COMP|34999-3|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C1369857|T201|COMP|35003-3|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1369858|T201|COMP|35019-9|LNC|Monocytes+Macrophages/100 lymphocytes|Monocytes+Macrophages/100 lymphocytes
C1369859|T201|COMP|35020-7|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1369860|T201|COMP|35021-5|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1369861|T201|COMP|35022-3|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1369862|T201|COMP|35023-1|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1369863|T201|COMP|35029-8|LNC|Monoblasts|Monoblasts
C1369864|T201|COMP|35039-7|LNC|Lymphocytes.plasmacytoid|Lymphocytes.plasmacytoid
C1369865|T201|COMP|35040-5|LNC|Lymphocytes.immunoblastic|Lymphocytes.immunoblastic
C1369866|T201|COMP|35046-2|LNC|Lymphocytes.abnormal|Lymphocytes.abnormal
C1369867|T201|COMP|35050-4|LNC|Lymphoblasts|Lymphoblasts
C1369868|T201|COMP|35055-3|LNC|Histiocytes/100 leukocytes|Histiocytes/100 leukocytes
C1369869|T201|COMP|35057-9|LNC|Histiocytes|Histiocytes
C1369870|T201|COMP|35069-4|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1369871|T201|COMP|35070-2|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1369872|T201|COMP|35073-6|LNC|Basophils|Basophils
C1369873|T201|COMP|35075-1|LNC|Basophils|Basophils
C1369874|T201|COMP|35077-7|LNC|Lymphocytes.abnormal/100 leukocytes|Lymphocytes.abnormal/100 leukocytes
C1369875|T201|COMP|35083-5|LNC|Amino acids panel|Amino acids panel
C1369876|T201|COMP|35084-3|LNC|Fetal lung maturity|Fetal lung maturity
C1369877|T201|COMP|35085-0|LNC|Newborn screening panel|Newborn screening panel
C1369878|T201|COMP|35086-8|LNC|Second trimester triple maternal screen panel|Second trimester triple maternal screen panel
C1369879|T201|COMP|35087-6|LNC|Amino acids panel|Amino acids panel
C1369889|T201|COMP|35100-7|LNC|Enterovirus Ab.IgM|Enterovirus Ab.IgM
C1369890|T201|COMP|35101-5|LNC|Intrathecal pressure|Intrathecal pressure
C1369891|T201|COMP|35102-3|LNC|Acenocoumarol|Acenocoumarol
C1369892|T201|COMP|35103-1|LNC|Acyclovir^trough|Acyclovir^trough
C1369893|T201|COMP|35104-9|LNC|Acyclovir^peak|Acyclovir^peak
C1369894|T201|COMP|35105-6|LNC|Bromperidol|Bromperidol
C1369895|T201|COMP|35106-4|LNC|Norcitalopram|Norcitalopram
C1369896|T201|COMP|35107-2|LNC|Norclobazam|Norclobazam
C1369897|T201|COMP|35108-0|LNC|Normaprotiline|Normaprotiline
C1369898|T201|COMP|35109-8|LNC|Phenprocoumon|Phenprocoumon
C1369899|T201|COMP|35110-6|LNC|Flecainide^trough|Flecainide^trough
C1369900|T201|COMP|35111-4|LNC|Flecainide^peak|Flecainide^peak
C1369901|T201|COMP|35112-2|LNC|Floxacillin|Floxacillin
C1369902|T201|COMP|35113-0|LNC|Nelfinavir M8|Nelfinavir M8
C1369903|T201|COMP|35114-8|LNC|Nordothiepin|Nordothiepin
C1369904|T201|COMP|35115-5|LNC|Pipamperone|Pipamperone
C1369905|T201|COMP|35116-3|LNC|Sulforidazine|Sulforidazine
C1369906|T201|COMP|35117-1|LNC|Sulpiride|Sulpiride
C1369907|T201|COMP|35118-9|LNC|Acetaldehyde|Acetaldehyde
C1369908|T201|COMP|35119-7|LNC|Chloral hydrate|Chloral hydrate
C1369909|T201|COMP|35120-5|LNC|Dothiepin sulfoxide|Dothiepin sulfoxide
C1369910|T201|COMP|35121-3|LNC|E-10-Hydroxynortriptyline|E-10-Hydroxynortriptyline
C1369911|T201|COMP|35122-1|LNC|MTM1 gene targeted mutation analysis|MTM1 gene targeted mutation analysis
C1369912|T201|COMP|35123-9|LNC|Chromosome 14 uniparental disomy|Chromosome 14 uniparental disomy
C1369913|T201|COMP|35124-7|LNC|Dysferlin|Dysferlin
C1369914|T201|COMP|35125-4|LNC|Hemoglobin Lepore/Hemoglobin.total|Hemoglobin Lepore/Hemoglobin.total
C1369915|T201|COMP|35126-2|LNC|Hemoglobin O-Arab/Hemoglobin.total|Hemoglobin O-Arab/Hemoglobin.total
C1369916|T201|COMP|35127-0|LNC|Hemoglobin A2.prime/Hemoglobin.total|Hemoglobin A2.prime/Hemoglobin.total
C1369917|T201|COMP|35128-8|LNC|Perforin|Perforin
C1369918|T201|COMP|35129-6|LNC|Karyotype|Karyotype
C1369919|T201|COMP|35130-4|LNC|Salicylates|Salicylates
C1369920|T201|COMP|35131-2|LNC|L-dopa decarboxylase|L-dopa decarboxylase
C1369921|T201|COMP|35132-0|LNC|MELAS gene targeted mutation analysis|MELAS gene targeted mutation analysis
C1369922|T201|COMP|35133-8|LNC|Glutarate|Glutarate
C1369923|T201|COMP|35134-6|LNC|Thyrotropin Ab|Thyrotropin Ab
C1369924|T201|COMP|35135-3|LNC|Adenosine triphosphate/Adenosine diphosphate|Adenosine triphosphate/Adenosine diphosphate
C1369925|T201|COMP|35136-1|LNC|Patient symptoms^3H post dose lactose PO|Patient symptoms^3H post dose lactose PO
C1369926|T201|COMP|35137-9|LNC|MECP2 gene targeted mutation analysis|MECP2 gene targeted mutation analysis
C1369927|T201|COMP|35138-7|LNC|MEFV gene mutations tested for|MEFV gene mutations tested for
C1369928|T201|COMP|35139-5|LNC|Interferon.beta Ab|Interferon.beta Ab
C1369929|T201|COMP|35140-3|LNC|Trans-3-Hydroxycotinine|Trans-3-Hydroxycotinine
C1369930|T201|COMP|35141-1|LNC|Purine nucleoside phosphorylase|Purine nucleoside phosphorylase
C1369931|T201|COMP|35142-9|LNC|Amphiphysin Ab|Amphiphysin Ab
C1369932|T201|COMP|35143-7|LNC|Purkinje cell cytoplasmic type 2 Ab|Purkinje cell cytoplasmic type 2 Ab
C1369933|T201|COMP|35144-5|LNC|Neuronal nuclear type 3 Ab|Neuronal nuclear type 3 Ab
C1369934|T201|COMP|35145-2|LNC|Octanoate|Octanoate
C1369935|T201|COMP|35146-0|LNC|Decanoate|Decanoate
C1369936|T201|COMP|35147-8|LNC|Decenoate|Decenoate
C1369937|T201|COMP|35148-6|LNC|Tetradecadienoate|Tetradecadienoate
C1369938|T201|COMP|35149-4|LNC|Octadecanoate|Octadecanoate
C1369939|T201|COMP|35150-2|LNC|Laurate|Laurate
C1369940|T201|COMP|35151-0|LNC|Lauroleate|Lauroleate
C1369941|T201|COMP|35152-8|LNC|Fatty acids.very long chain.C26:0|Fatty acids.very long chain.C26:0
C1369942|T201|COMP|35153-6|LNC|Fatty acids.very long chain.C26:1|Fatty acids.very long chain.C26:1
C1369943|T201|COMP|35154-4|LNC|Hexadecadienoate|Hexadecadienoate
C1369944|T201|COMP|35155-1|LNC|Hexadecenoate|Hexadecenoate
C1369945|T201|COMP|35156-9|LNC|Fatty acids.very long chain.C24:0|Fatty acids.very long chain.C24:0
C1369946|T201|COMP|35157-7|LNC|Myristate|Myristate
C1369947|T201|COMP|35158-5|LNC|Myristoleate|Myristoleate
C1369948|T201|COMP|35159-3|LNC|Fatty acids.very long chain.C22:0|Fatty acids.very long chain.C22:0
C1369949|T201|COMP|35160-1|LNC|Docosenoate|Docosenoate
C1369950|T201|COMP|35161-9|LNC|Palmitate|Palmitate
C1369951|T201|COMP|35162-7|LNC|Palmitoleate|Palmitoleate
C1369952|T201|COMP|35163-5|LNC|Gamma linolenate|Gamma linolenate
C1369953|T201|COMP|35164-3|LNC|Alpha linolenate|Alpha linolenate
C1369954|T201|COMP|35165-0|LNC|Linoleate|Linoleate
C1369955|T201|COMP|35166-8|LNC|Oleate|Oleate
C1369956|T201|COMP|35167-6|LNC|Vaccenate|Vaccenate
C1369957|T201|COMP|35168-4|LNC|Arachidonate|Arachidonate
C1369958|T201|COMP|35169-2|LNC|Arachidate|Arachidate
C1369959|T201|COMP|35170-0|LNC|Nervonate|Nervonate
C1369960|T201|COMP|35171-8|LNC|Homo-gamma linolenate|Homo-gamma linolenate
C1369961|T201|COMP|35172-6|LNC|Mead acid|Mead acid
C1369962|T201|COMP|35173-4|LNC|Eicosapentaenoate|Eicosapentaenoate
C1369963|T201|COMP|35174-2|LNC|Docosahexaenoate|Docosahexaenoate
C1369964|T201|COMP|35175-9|LNC|Fatty acids.saturated|Fatty acids.saturated
C1369965|T201|COMP|35176-7|LNC|Fatty acids.monounsaturated|Fatty acids.monounsaturated
C1369966|T201|COMP|35177-5|LNC|Fatty acids.polyunsaturated|Fatty acids.polyunsaturated
C1369967|T201|COMP|35178-3|LNC|Fatty acids.omega 3|Fatty acids.omega 3
C1369968|T201|COMP|35179-1|LNC|Fatty acids.omega 6|Fatty acids.omega 6
C1369969|T201|COMP|35180-9|LNC|Docosapentaenate w3|Docosapentaenate w3
C1369970|T201|COMP|35181-7|LNC|Docosapentaenate w6|Docosapentaenate w6
C1369971|T201|COMP|35182-5|LNC|Docosatetraenoate|Docosatetraenoate
C1369972|T201|COMP|35183-3|LNC|Hemoglobin|Hemoglobin
C1369982|T201|COMP|1974-5|LNC|Bilirubin|Bilirubin
C1370010|T201|COMP|2777-1|LNC|Phosphate|Phosphate
C1370054|T201|COMP|35265-8|LNC|Path report.addendum|Path report.addendum
C1370055|T201|COMP|35266-6|LNC|Gleason score|Gleason score
C1370056|T201|COMP|35267-4|LNC|Age at pathology Dx|Age at pathology Dx
C1370058|T201|COMP|35269-0|LNC|Bartonella henselae Ab|Bartonella henselae Ab
C1370059|T201|COMP|35270-8|LNC|Candida sp Ab|Candida sp Ab
C1370060|T201|COMP|35271-6|LNC|Candida sp Ag|Candida sp Ag
C1370061|T201|COMP|35272-4|LNC|Centromere Ab.IgG|Centromere Ab.IgG
C1370062|T201|COMP|35273-2|LNC|Hepatitis D virus Ab.IgG|Hepatitis D virus Ab.IgG
C1370063|T201|COMP|35274-0|LNC|Histone Ab.IgG|Histone Ab.IgG
C1370064|T201|COMP|35275-7|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C1370065|T201|COMP|35276-5|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C1370066|T201|COMP|35277-3|LNC|Myocardium Ab.IgG|Myocardium Ab.IgG
C1370067|T201|COMP|35278-1|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C1370068|T201|COMP|35279-9|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C1370069|T201|COMP|35280-7|LNC|Tissue transglutaminase Ab.IgA|Tissue transglutaminase Ab.IgA
C1370070|T201|COMP|35281-5|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C1370071|T201|COMP|35282-3|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C1370072|T201|COMP|35283-1|LNC|Hepatitis D virus Ab.IgG|Hepatitis D virus Ab.IgG
C1370073|T201|COMP|35284-9|LNC|Histone Ab.IgG|Histone Ab.IgG
C1370074|T201|COMP|35285-6|LNC|Tissue transglutaminase Ab.IgA|Tissue transglutaminase Ab.IgA
C1378206|T201|COMP|35047-0|LNC|Lymphocytes.abnormal|Lymphocytes.abnormal
C1378210|T201|COMP|35048-8|LNC|Lymphocytes.abnormal|Lymphocytes.abnormal
C1378214|T201|COMP|35043-9|LNC|Lymphocytes.variant|Lymphocytes.variant
C1378215|T201|COMP|35045-4|LNC|Lymphocytes.variant|Lymphocytes.variant
C1378216|T201|COMP|35042-1|LNC|Lymphocytes.variant|Lymphocytes.variant
C1378217|T201|COMP|35041-3|LNC|Lymphocytes.variant|Lymphocytes.variant
C1378218|T201|COMP|35044-7|LNC|Lymphocytes.variant|Lymphocytes.variant
C1378223|T201|COMP|35072-8|LNC|Basophils|Basophils
C1378224|T201|COMP|35071-0|LNC|Basophils|Basophils
C1378225|T201|COMP|35074-4|LNC|Basophils|Basophils
C1378226|T201|COMP|35068-6|LNC|Blasts|Blasts
C1378227|T201|COMP|34958-9|LNC|Eosinophils|Eosinophils
C1378230|T201|COMP|35067-8|LNC|Blasts|Blasts
C1378231|T201|COMP|35066-0|LNC|Blasts|Blasts
C1378232|T201|COMP|34957-1|LNC|Eosinophils|Eosinophils
C1378233|T201|COMP|35065-2|LNC|Blasts|Blasts
C1378236|T201|COMP|35064-5|LNC|Blasts|Blasts
C1378237|T201|COMP|35063-7|LNC|Eosinophils|Eosinophils
C1378239|T201|COMP|35062-9|LNC|Eosinophils|Eosinophils
C1378240|T201|COMP|35061-1|LNC|Eosinophils|Eosinophils
C1378241|T201|COMP|35060-3|LNC|Eosinophils|Eosinophils
C1378250|T201|COMP|34651-0|LNC|CYP21A2 gene targeted mutation analysis|CYP21A2 gene targeted mutation analysis
C1378253|T201|COMP|34603-1|LNC|I Ab|I Ab
C1378254|T201|COMP|34975-3|LNC|DNA index|DNA index
C1378258|T201|COMP|35059-5|LNC|Granulocytes|Granulocytes
C1378264|T201|COMP|35058-7|LNC|Hairy cells/100 leukocytes|Hairy cells/100 leukocytes
C1378269|T201|COMP|34602-3|LNC|E Ab|E Ab
C1378279|T201|COMP|35056-1|LNC|Histiocytes|Histiocytes
C1378285|T201|COMP|35051-2|LNC|Leukocytes other|Leukocytes other
C1378287|T201|COMP|35052-0|LNC|Leukocytes other|Leukocytes other
C1378288|T201|COMP|35054-6|LNC|Leukocytes other|Leukocytes other
C1378289|T201|COMP|35053-8|LNC|Leukocytes other|Leukocytes other
C1378290|T201|COMP|35082-7|LNC|Lymphocytes.large granular|Lymphocytes.large granular
C1378297|T201|COMP|35098-3|LNC|Lymphocytes|Lymphocytes
C1378304|T201|COMP|35006-6|LNC|Plasma cells|Plasma cells
C1378305|T201|COMP|35097-5|LNC|Lymphocytes|Lymphocytes
C1378306|T201|COMP|35049-6|LNC|Lymphocytes|Lymphocytes
C1378307|T201|COMP|35081-9|LNC|Lymphocytes+Monocytes|Lymphocytes+Monocytes
C1378311|T201|COMP|35038-9|LNC|Macrophages|Macrophages
C1378313|T201|COMP|35036-3|LNC|Macrophages|Macrophages
C1378314|T201|COMP|35037-1|LNC|Macrophages|Macrophages
C1378316|T201|COMP|35001-7|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1378317|T201|COMP|35002-5|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1378318|T201|COMP|35000-9|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1378319|T201|COMP|35005-8|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1378321|T201|COMP|35004-1|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C1378324|T201|COMP|35034-8|LNC|Mesothelial cells|Mesothelial cells
C1378325|T201|COMP|35079-3|LNC|Mesothelial cells|Mesothelial cells
C1378327|T201|COMP|35033-0|LNC|Mesothelial cells|Mesothelial cells
C1378329|T201|COMP|35032-2|LNC|Mesothelial cells|Mesothelial cells
C1378330|T201|COMP|35035-5|LNC|Mesothelial cells|Mesothelial cells
C1378331|T201|COMP|34998-5|LNC|Prolymphocytes|Prolymphocytes
C1378332|T201|COMP|35030-6|LNC|Metamyelocytes|Metamyelocytes
C1378333|T201|COMP|34926-6|LNC|Promonocytes|Promonocytes
C1378334|T201|COMP|34997-7|LNC|Promonocytes|Promonocytes
C1378335|T201|COMP|35031-4|LNC|Metamyelocytes|Metamyelocytes
C1378336|T201|COMP|34995-1|LNC|Promyelocytes|Promyelocytes
C1378337|T201|COMP|35026-4|LNC|Monocytes|Monocytes
C1378338|T201|COMP|35076-9|LNC|Monocytes|Monocytes
C1378339|T201|COMP|34996-9|LNC|Promyelocytes|Promyelocytes
C1378341|T201|COMP|35028-0|LNC|Monocytes|Monocytes
C1378342|T201|COMP|35027-2|LNC|Monocytes|Monocytes
C1378343|T201|COMP|35099-1|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1378344|T201|COMP|35025-6|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1378361|T201|COMP|35024-9|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C1378363|T201|COMP|35018-1|LNC|Mononuclear cells|Mononuclear cells
C1378364|T201|COMP|35080-1|LNC|Mononuclear cells|Mononuclear cells
C1378397|T201|COMP|34657-7|LNC|Spermatozoa.immotile|Spermatozoa.immotile
C1378400|T201|COMP|35017-3|LNC|Myelocytes|Myelocytes
C1378401|T201|COMP|35016-5|LNC|Myelocytes|Myelocytes
C1378407|T201|COMP|35015-7|LNC|Neutrophils.band form|Neutrophils.band form
C1378408|T201|COMP|35014-0|LNC|Neutrophils.band form|Neutrophils.band form
C1378409|T201|COMP|35013-2|LNC|Neutrophils.band form|Neutrophils.band form
C1378410|T201|COMP|35011-6|LNC|Neutrophils.segmented|Neutrophils.segmented
C1378412|T201|COMP|35012-4|LNC|Neutrophils.segmented|Neutrophils.segmented
C1378413|T201|COMP|35010-8|LNC|Neutrophils.segmented|Neutrophils.segmented
C1378414|T201|COMP|35009-0|LNC|Neutrophils.segmented|Neutrophils.segmented
C1378415|T201|COMP|35007-4|LNC|Nonhematic cells|Nonhematic cells
C1378416|T201|COMP|35008-2|LNC|Nonhematic cells|Nonhematic cells
C1382693|T201|COMP|35078-5|LNC|Unspecified cells|Unspecified cells
C1382694|T201|COMP|34987-8|LNC|Unidentified cells|Unidentified cells
C1507396|T201|COMP|35618-8|LNC|Methadone|Methadone
C1507397|T201|COMP|35619-6|LNC|Methaqualone|Methaqualone
C1507398|T201|COMP|35620-4|LNC|Metoprolol|Metoprolol
C1507399|T201|COMP|35621-2|LNC|Norclomipramine|Norclomipramine
C1507400|T201|COMP|35622-0|LNC|Nordiazepam|Nordiazepam
C1507401|T201|COMP|35623-8|LNC|Nordoxepin|Nordoxepin
C1507402|T201|COMP|35624-6|LNC|Norfluoxetine|Norfluoxetine
C1507403|T201|COMP|35625-3|LNC|Normeperidine|Normeperidine
C1507404|T201|COMP|35812-7|LNC|Garenoxacin|Garenoxacin
C1507405|T201|COMP|35813-5|LNC|Garenoxacin|Garenoxacin
C1507406|T201|COMP|35814-3|LNC|Gemifloxacin|Gemifloxacin
C1507407|T201|COMP|35815-0|LNC|Gemifloxacin|Gemifloxacin
C1507408|T201|COMP|35816-8|LNC|Gemifloxacin|Gemifloxacin
C1507409|T201|COMP|35817-6|LNC|Gentamicin.high potency|Gentamicin.high potency
C1507410|T201|COMP|35818-4|LNC|Grepafloxacin|Grepafloxacin
C1507411|T201|COMP|35819-2|LNC|Imipenem+EDTA|Imipenem+EDTA
C1507412|T201|COMP|35865-5|LNC|Lipoprotein.intermediate density|Lipoprotein.intermediate density
C1507413|T201|COMP|35866-3|LNC|Organic acids panel|Organic acids panel
C1507414|T201|COMP|35867-1|LNC|Acetoacetate|Acetoacetate
C1507415|T201|COMP|35305-2|LNC|Toxoplasma gondii AC Ab|Toxoplasma gondii AC Ab
C1507416|T201|COMP|35306-0|LNC|TTR gene allele 2|TTR gene allele 2
C1507417|T201|COMP|35307-8|LNC|TTR gene allele 1|TTR gene allele 1
C1507418|T201|COMP|35308-6|LNC|Trypsin^5th specimen post dose sincalide|Trypsin^5th specimen post dose sincalide
C1507419|T201|COMP|35309-4|LNC|Trypsin^4th specimen post dose sincalide|Trypsin^4th specimen post dose sincalide
C1507420|T201|COMP|35310-2|LNC|Trypsin^3rd specimen post dose sincalide|Trypsin^3rd specimen post dose sincalide
C1507421|T201|COMP|35311-0|LNC|Trypsin^2nd specimen post dose sincalide|Trypsin^2nd specimen post dose sincalide
C1507422|T201|COMP|35312-8|LNC|Trypsin^1st specimen post dose sincalide|Trypsin^1st specimen post dose sincalide
C1507424|T201|COMP|35859-8|LNC|Virginiamycin|Virginiamycin
C1507425|T201|COMP|35860-6|LNC|Virginiamycin|Virginiamycin
C1507426|T201|COMP|35861-4|LNC|Virginiamycin|Virginiamycin
C1507427|T201|COMP|35862-2|LNC|Voriconazole|Voriconazole
C1507428|T201|COMP|35863-0|LNC|Voriconazole|Voriconazole
C1507430|T201|COMP|35287-2|LNC|Toxoplasma gondii HS Ab|Toxoplasma gondii HS Ab
C1507431|T201|COMP|35288-0|LNC|MEN1 gene targeted mutation analysis|MEN1 gene targeted mutation analysis
C1507432|T201|COMP|35289-8|LNC|Peroxide hemolysis|Peroxide hemolysis
C1507433|T201|COMP|35290-6|LNC|RPS6KA3 gene targeted mutation analysis|RPS6KA3 gene targeted mutation analysis
C1507434|T201|COMP|35291-4|LNC|UBE3A gene targeted mutation analysis|UBE3A gene targeted mutation analysis
C1507435|T201|COMP|35292-2|LNC|Chromosome 11 uniparental disomy|Chromosome 11 uniparental disomy
C1507436|T201|COMP|35293-0|LNC|TYR gene targeted mutation analysis|TYR gene targeted mutation analysis
C1507437|T201|COMP|35294-8|LNC|PYGM gene targeted mutation analysis|PYGM gene targeted mutation analysis
C1507438|T201|COMP|35295-5|LNC|BTK gene targeted mutation analysis|BTK gene targeted mutation analysis
C1507439|T201|COMP|35296-3|LNC|PAX3 gene targeted mutation analysis|PAX3 gene targeted mutation analysis
C1507440|T201|COMP|35297-1|LNC|LMNA gene targeted mutation analysis|LMNA gene targeted mutation analysis
C1507441|T201|COMP|35298-9|LNC|FXN gene targeted mutation analysis|FXN gene targeted mutation analysis
C1507442|T201|COMP|35299-7|LNC|PSEN1 gene targeted mutation analysis|PSEN1 gene targeted mutation analysis
C1507443|T201|COMP|35300-3|LNC|GJB2 gene targeted mutation analysis|GJB2 gene targeted mutation analysis
C1507444|T201|COMP|35301-1|LNC|Transferrin.carbohydrate deficient.asialo|Transferrin.carbohydrate deficient.asialo
C1507445|T201|COMP|35302-9|LNC|HYAL1 gene targeted mutation analysis|HYAL1 gene targeted mutation analysis
C1507446|T201|COMP|35303-7|LNC|Glucosylceramidase|Glucosylceramidase
C1507447|T201|COMP|35304-5|LNC|CLA2 gene targeted mutation analysis|CLA2 gene targeted mutation analysis
C1507451|T201|COMP|35317-7|LNC|Thermoactinomyces vulgaris 1 Ab|Thermoactinomyces vulgaris 1 Ab
C1507452|T201|COMP|35318-5|LNC|Thermoactinomyces sacchari Ab|Thermoactinomyces sacchari Ab
C1507453|T201|COMP|35319-3|LNC|Protein^5th specimen post dose sincalide|Protein^5th specimen post dose sincalide
C1507454|T201|COMP|35320-1|LNC|Protein^4th specimen post dose sincalide|Protein^4th specimen post dose sincalide
C1507455|T201|COMP|35321-9|LNC|Protein^3rd specimen post dose sincalide|Protein^3rd specimen post dose sincalide
C1507456|T201|COMP|35322-7|LNC|Protein^2nd specimen post dose sincalide|Protein^2nd specimen post dose sincalide
C1507457|T201|COMP|35323-5|LNC|Protein^1st specimen post dose sincalide|Protein^1st specimen post dose sincalide
C1507458|T201|COMP|35324-3|LNC|PMP22 gene allele 1|PMP22 gene allele 1
C1507459|T201|COMP|35325-0|LNC|PMP22 gene allele 2|PMP22 gene allele 2
C1507460|T201|COMP|35326-8|LNC|pH^5th specimen post dose sincalide|pH^5th specimen post dose sincalide
C1507461|T201|COMP|35327-6|LNC|pH^4th specimen post dose sincalide|pH^4th specimen post dose sincalide
C1507462|T201|COMP|35328-4|LNC|pH^3rd specimen post dose sincalide|pH^3rd specimen post dose sincalide
C1507463|T201|COMP|35329-2|LNC|pH^2nd specimen post dose sincalide|pH^2nd specimen post dose sincalide
C1507464|T201|COMP|35330-0|LNC|pH^1st specimen post dose sincalide|pH^1st specimen post dose sincalide
C1507465|T201|COMP|35331-8|LNC|OXcarbazepine|OXcarbazepine
C1507466|T201|COMP|35332-6|LNC|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C1507467|T201|COMP|35333-4|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C1507468|T201|COMP|35334-2|LNC|Collagen crosslinked N-telopeptide|Collagen crosslinked N-telopeptide
C1507469|T201|COMP|35335-9|LNC|Chymotrypsin^5th specimen post dose sincalide|Chymotrypsin^5th specimen post dose sincalide
C1507470|T201|COMP|35336-7|LNC|Chymotrypsin^4th specimen post dose sincalide|Chymotrypsin^4th specimen post dose sincalide
C1507471|T201|COMP|35337-5|LNC|Chymotrypsin^3rd specimen post dose sincalide|Chymotrypsin^3rd specimen post dose sincalide
C1507472|T201|COMP|35338-3|LNC|Chymotrypsin^2nd specimen post dose sincalide|Chymotrypsin^2nd specimen post dose sincalide
C1507473|T201|COMP|35339-1|LNC|Chymotrypsin^1st specimen post dose sincalide|Chymotrypsin^1st specimen post dose sincalide
C1507474|T201|COMP|35340-9|LNC|ASPA gene.p.Tyr231Ter|ASPA gene.p.Tyr231Ter
C1507475|T201|COMP|35341-7|LNC|ASPA gene.p.Ala305Glu|ASPA gene.p.Ala305Glu
C1507476|T201|COMP|35342-5|LNC|Amylase^5th specimen post dose sincalide|Amylase^5th specimen post dose sincalide
C1507477|T201|COMP|35343-3|LNC|Amylase^4th specimen post dose sincalide|Amylase^4th specimen post dose sincalide
C1507478|T201|COMP|35344-1|LNC|Amylase^3rd specimen post dose sincalide|Amylase^3rd specimen post dose sincalide
C1507479|T201|COMP|35345-8|LNC|Amylase^2nd specimen post dose sincalide|Amylase^2nd specimen post dose sincalide
C1507480|T201|COMP|35346-6|LNC|Amylase^1st specimen post dose sincalide|Amylase^1st specimen post dose sincalide
C1507482|T201|COMP|35348-2|LNC|Corynebacterium diphtheriae Ab|Corynebacterium diphtheriae Ab
C1507483|T201|COMP|35349-0|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C1507486|T201|COMP|35352-4|LNC|Mycobacterium tuberculosis genotype|Mycobacterium tuberculosis genotype
C1507487|T201|COMP|35353-2|LNC|FSHD gene targeted mutation analysis|FSHD gene targeted mutation analysis
C1507488|T201|COMP|35354-0|LNC|COL1A1+COL1A2 gene targeted mutation analysis|COL1A1+COL1A2 gene targeted mutation analysis
C1507489|T201|COMP|38406-5|LNC|PABPN1 gene targeted mutation analysis|PABPN1 gene targeted mutation analysis
C1507490|T201|COMP|35356-5|LNC|TWIST1 gene targeted mutation analysis|TWIST1 gene targeted mutation analysis
C1507491|T201|COMP|35357-3|LNC|PEO gene targeted mutation analysis|PEO gene targeted mutation analysis
C1507492|T201|COMP|35358-1|LNC|LHON syndrome gene targeted mutation analysis|LHON syndrome gene targeted mutation analysis
C1507493|T201|COMP|35359-9|LNC|AR gene targeted mutation analysis|AR gene targeted mutation analysis
C1507494|T201|COMP|35360-7|LNC|Triglyceride.in lipoprotein (little a)|Triglyceride.in lipoprotein (little a)
C1507495|T201|COMP|35361-5|LNC|Triglyceride.in lipoprotein (little a)|Triglyceride.in lipoprotein (little a)
C1507496|T201|COMP|35362-3|LNC|Triglyceride.in chylomicrons|Triglyceride.in chylomicrons
C1507497|T201|COMP|35363-1|LNC|Triglyceride.in chylomicrons|Triglyceride.in chylomicrons
C1507499|T201|COMP|35365-6|LNC|Vitamin D+Metabolites|Vitamin D+Metabolites
C1507500|T201|COMP|35366-4|LNC|SCA2 gene allele 2.CAG repeats|SCA2 gene allele 2.CAG repeats
C1507501|T201|COMP|35367-2|LNC|SCA2 gene allele 1.CAG repeats|SCA2 gene allele 1.CAG repeats
C1507502|T201|COMP|35368-0|LNC|SCA1 gene allele 2.CAG repeats|SCA1 gene allele 2.CAG repeats
C1507503|T201|COMP|35369-8|LNC|SCA1 gene allele 1.CAG repeats|SCA1 gene allele 1.CAG repeats
C1507504|T201|COMP|35370-6|LNC|GBA gene.g.S84GG|GBA gene.g.S84GG
C1507505|T201|COMP|35371-4|LNC|GBA gene.g.N370S|GBA gene.g.N370S
C1507506|T201|COMP|35372-2|LNC|GBA gene.p.Leu444Pro|GBA gene.p.Leu444Pro
C1507507|T201|COMP|35373-0|LNC|Platelet aggregation.XXX induced|Platelet aggregation.XXX induced
C1507508|T201|COMP|35374-8|LNC|DMPK gene allele 2.CTG repeats|DMPK gene allele 2.CTG repeats
C1507509|T201|COMP|35375-5|LNC|DMPK gene allele 1.CTG repeats|DMPK gene allele 1.CTG repeats
C1507510|T201|COMP|35376-3|LNC|MJD gene allele 2.CAG repeats|MJD gene allele 2.CAG repeats
C1507511|T201|COMP|35377-1|LNC|MJD gene allele 1.CAG repeats|MJD gene allele 1.CAG repeats
C1507512|T201|COMP|35378-9|LNC|HNPCC genes mutations tested for|HNPCC genes mutations tested for
C1507513|T201|COMP|35379-7|LNC|HNPCC genes targeted mutation analysis|HNPCC genes targeted mutation analysis
C1507514|T201|COMP|35380-5|LNC|HEXA gene.c.IVS7+1G>A|HEXA gene.c.IVS7+1G>A
C1507515|T201|COMP|35381-3|LNC|HEXA gene.c.IVS12+1G>C|HEXA gene.c.IVS12+1G>C
C1507516|T201|COMP|35382-1|LNC|HEXA gene.p.Gly269Ser|HEXA gene.p.Gly269Ser
C1507517|T201|COMP|35383-9|LNC|Galactomannan Ag|Galactomannan Ag
C1507518|T201|COMP|35384-7|LNC|Estradiol|Estradiol
C1507519|T201|COMP|35385-4|LNC|CV2 Ab.IgG|CV2 Ab.IgG
C1507520|T201|COMP|35386-2|LNC|CV2 Ab.IgG|CV2 Ab.IgG
C1507521|T201|COMP|35387-0|LNC|Cholesterol.in lipoprotein (little a)|Cholesterol.in lipoprotein (little a)
C1507522|T201|COMP|35388-8|LNC|Cholesterol.in lipoprotein (little a)|Cholesterol.in lipoprotein (little a)
C1507523|T201|COMP|35389-6|LNC|Cholesterol.in chylomicrons|Cholesterol.in chylomicrons
C1507524|T201|COMP|35390-4|LNC|Vaccinia virus DNA|Vaccinia virus DNA
C1507525|T201|COMP|35391-2|LNC|Taenia solium larva Ab.IgG|Taenia solium larva Ab.IgG
C1507526|T201|COMP|35392-0|LNC|Hantavirus Ab.IgG|Hantavirus Ab.IgG
C1507527|T201|COMP|35393-8|LNC|Hantavirus Ab.IgM|Hantavirus Ab.IgM
C1507528|T201|COMP|35394-6|LNC|Legionella pneumophila 1 Ab.IgG|Legionella pneumophila 1 Ab.IgG
C1507529|T201|COMP|35395-3|LNC|Legionella pneumophila 1 Ab.IgM|Legionella pneumophila 1 Ab.IgM
C1507530|T201|COMP|35396-1|LNC|Enterovirus RNA|Enterovirus RNA
C1507531|T201|COMP|35397-9|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1507532|T201|COMP|35398-7|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1507533|T201|COMP|35399-5|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1507534|T201|COMP|35400-1|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1507535|T201|COMP|35401-9|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1507536|T201|COMP|35402-7|LNC|Leishmania donovani Ab.IgG|Leishmania donovani Ab.IgG
C1507537|T201|COMP|35403-5|LNC|Leishmania donovani Ab.IgM|Leishmania donovani Ab.IgM
C1507538|T201|COMP|35404-3|LNC|Leishmania braziliensis Ab.IgG|Leishmania braziliensis Ab.IgG
C1507539|T201|COMP|35405-0|LNC|Leishmania braziliensis Ab.IgM|Leishmania braziliensis Ab.IgM
C1507540|T201|COMP|35406-8|LNC|Leishmania mexicana Ab.IgG|Leishmania mexicana Ab.IgG
C1507541|T201|COMP|35407-6|LNC|Leishmania mexicana Ab.IgM|Leishmania mexicana Ab.IgM
C1507542|T201|COMP|35408-4|LNC|Leishmania tropica Ab.IgG|Leishmania tropica Ab.IgG
C1507543|T201|COMP|35409-2|LNC|Leishmania tropica Ab.IgM|Leishmania tropica Ab.IgM
C1507545|T201|COMP|35411-8|LNC|Trienoate/Arachidonate|Trienoate/Arachidonate
C1507546|T201|COMP|35412-6|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507547|T201|COMP|35413-4|LNC|Coxsackievirus A4+A16 Ab|Coxsackievirus A4+A16 Ab
C1507548|T201|COMP|35414-2|LNC|Specific gravity|Specific gravity
C1507549|T201|COMP|35415-9|LNC|Oxytocin|Oxytocin
C1507550|T201|COMP|35416-7|LNC|Echinococcus granulosus Ab|Echinococcus granulosus Ab
C1507551|T201|COMP|35417-5|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507552|T201|COMP|35418-3|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507553|T201|COMP|35419-1|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507554|T201|COMP|35420-9|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507555|T201|COMP|35421-7|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507556|T201|COMP|35422-5|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507557|T201|COMP|35423-3|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507558|T201|COMP|35424-1|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507559|T201|COMP|35425-8|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507560|T201|COMP|35426-6|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507561|T201|COMP|35427-4|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507562|T201|COMP|35428-2|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507563|T201|COMP|35429-0|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507564|T201|COMP|35430-8|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507565|T201|COMP|35431-6|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507566|T201|COMP|35432-4|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507567|T201|COMP|35433-2|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507568|T201|COMP|35434-0|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507569|T201|COMP|35435-7|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C1507570|T201|COMP|35436-5|LNC|Spermatozoa^post reanastomosis|Spermatozoa^post reanastomosis
C1507571|T201|COMP|35437-3|LNC|HIV 1 Ab|HIV 1 Ab
C1507572|T201|COMP|35438-1|LNC|HIV 1 Ab|HIV 1 Ab
C1507573|T201|COMP|35439-9|LNC|HIV 1 Ab|HIV 1 Ab
C1507574|T201|COMP|35440-7|LNC|HIV 1 gp160 Ab|HIV 1 gp160 Ab
C1507575|T201|COMP|35441-5|LNC|HIV 1 gp120 Ab|HIV 1 gp120 Ab
C1507576|T201|COMP|35442-3|LNC|HIV 1 p66 Ab|HIV 1 p66 Ab
C1507577|T201|COMP|35443-1|LNC|HIV 1 p65 Ab|HIV 1 p65 Ab
C1507578|T201|COMP|35444-9|LNC|HIV 1 p55 Ab|HIV 1 p55 Ab
C1507579|T201|COMP|35445-6|LNC|HIV 1 p51 Ab|HIV 1 p51 Ab
C1507580|T201|COMP|35446-4|LNC|HIV 1 gp41 Ab|HIV 1 gp41 Ab
C1507581|T201|COMP|35447-2|LNC|HIV 1 p31 Ab|HIV 1 p31 Ab
C1507582|T201|COMP|35448-0|LNC|HIV 1 p24 Ab|HIV 1 p24 Ab
C1507583|T201|COMP|35449-8|LNC|HIV 1 p17 Ab|HIV 1 p17 Ab
C1507584|T201|COMP|35450-6|LNC|HIV 1 p18 Ab|HIV 1 p18 Ab
C1507585|T201|COMP|35451-4|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1507586|T201|COMP|35452-2|LNC|HIV 1 gp40 Ab|HIV 1 gp40 Ab
C1507587|T201|COMP|35453-0|LNC|ARSA gene PD allele|ARSA gene PD allele
C1507588|T201|COMP|35454-8|LNC|MLL gene rearrangements|MLL gene rearrangements
C1507589|T201|COMP|35455-5|LNC|X chromosome inactivation|X chromosome inactivation
C1507590|T201|COMP|35456-3|LNC|Y chromosome deletion|Y chromosome deletion
C1507591|T201|COMP|35457-1|LNC|Maternal cell contamination|Maternal cell contamination
C1507592|T201|COMP|35458-9|LNC|Ma+Ta Ab|Ma+Ta Ab
C1507593|T201|COMP|35459-7|LNC|T cell crossmatch|T cell crossmatch
C1507594|T201|COMP|35460-5|LNC|Platelet genotype|Platelet genotype
C1507595|T201|COMP|35461-3|LNC|ELN gene targeted mutation analysis|ELN gene targeted mutation analysis
C1507596|T201|COMP|35462-1|LNC|SMN1 gene targeted mutation analysis|SMN1 gene targeted mutation analysis
C1507597|T201|COMP|35463-9|LNC|Telomere analysis|Telomere analysis
C1507598|T201|COMP|35464-7|LNC|CMT axonal gene targeted mutation analysis|CMT axonal gene targeted mutation analysis
C1507599|T201|COMP|35465-4|LNC|RHD gene targeted mutation analysis|RHD gene targeted mutation analysis
C1507600|T201|COMP|35466-2|LNC|AS+PWS gene targeted mutation analysis|AS+PWS gene targeted mutation analysis
C1507601|T201|COMP|35467-0|LNC|M-chlorophenylpiperazine|M-chlorophenylpiperazine
C1507602|T201|COMP|35468-8|LNC|Cells.FLAER|Cells.FLAER
C1507604|T201|COMP|35470-4|LNC|Mitochondria DNA deletion|Mitochondria DNA deletion
C1507605|T201|COMP|35471-2|LNC|HLA Ab|HLA Ab
C1507606|T201|COMP|35472-0|LNC|HEXA gene.c.1277insTATC|HEXA gene.c.1277insTATC
C1507607|T201|COMP|35473-8|LNC|HEXA gene 7.6kb deletion|HEXA gene 7.6kb deletion
C1507608|T201|COMP|35474-6|LNC|Gene XXX targeted mutation analysis|Gene XXX targeted mutation analysis
C1507610|T201|COMP|35476-1|LNC|OKT3 blocking Ab|OKT3 blocking Ab
C1507611|T201|COMP|35477-9|LNC|Ciliated columnar lining cells/100 leukocytes|Ciliated columnar lining cells/100 leukocytes
C1507612|T201|COMP|35478-7|LNC|Cytosol aminopeptidase|Cytosol aminopeptidase
C1507613|T201|COMP|35479-5|LNC|Diazinon|Diazinon
C1507614|T201|COMP|35480-3|LNC|1-Naphthol|1-Naphthol
C1507615|T201|COMP|35481-1|LNC|Terbufos|Terbufos
C1507616|T201|COMP|35482-9|LNC|Para nitrophenol|Para nitrophenol
C1507617|T201|COMP|35483-7|LNC|Mevinphos|Mevinphos
C1507618|T201|COMP|35484-5|LNC|Methyl parathion|Methyl parathion
C1507619|T201|COMP|35485-2|LNC|Metasystox|Metasystox
C1507620|T201|COMP|35486-0|LNC|Fonofos|Fonofos
C1507621|T201|COMP|35487-8|LNC|Fenchlorphos|Fenchlorphos
C1507622|T201|COMP|35488-6|LNC|Diazinon|Diazinon
C1507623|T201|COMP|35489-4|LNC|Chlorpyrifos|Chlorpyrifos
C1507624|T201|COMP|35490-2|LNC|Azinphos-methyl|Azinphos-methyl
C1507625|T201|COMP|35491-0|LNC|Leptospira sp DNA|Leptospira sp DNA
C1507626|T201|COMP|35492-8|LNC|Staphylococcus aureus.methicillin resistant DNA|Staphylococcus aureus.methicillin resistant DNA
C1507627|T201|COMP|35493-6|LNC|Ricin|Ricin
C1507628|T201|COMP|35494-4|LNC|Succinate dehydrogenase|Succinate dehydrogenase
C1507629|T201|COMP|35495-1|LNC|Citrate synthase|Citrate synthase
C1507630|T201|COMP|35496-9|LNC|NADH dehydrogenase|NADH dehydrogenase
C1507631|T201|COMP|35497-7|LNC|NADH cytochrome C reductase|NADH cytochrome C reductase
C1507632|T201|COMP|35498-5|LNC|Succinate cytochrome C reductase|Succinate cytochrome C reductase
C1507633|T201|COMP|35499-3|LNC|Pesticide & Insecticide panel|Pesticide & Insecticide panel
C1507634|T201|COMP|35500-8|LNC|Pesticide & Insecticide panel|Pesticide & Insecticide panel
C1507635|T201|COMP|35501-6|LNC|Pesticide & Insecticide panel|Pesticide & Insecticide panel
C1507636|T201|COMP|35502-4|LNC|Mitochondrial myopathy enzyme panel|Mitochondrial myopathy enzyme panel
C1507638|T201|COMP|35504-0|LNC|Para aminobenzoate^6H post XXX bentiromide PO|Para aminobenzoate^6H post XXX bentiromide PO
C1507639|T201|COMP|35505-7|LNC|Lipoprotein.beta.subparticle|Lipoprotein.beta.subparticle
C1507641|T201|COMP|35507-3|LNC|Amino acids panel|Amino acids panel
C1507642|T201|COMP|35508-1|LNC|Amino acids panel|Amino acids panel
C1507643|T201|COMP|35509-9|LNC|Amino acids panel|Amino acids panel
C1507663|T201|COMP|35529-7|LNC|Beef Ab.IgG|Beef Ab.IgG
C1507664|T201|COMP|35530-5|LNC|Candida albicans Ab.IgG|Candida albicans Ab.IgG
C1507665|T201|COMP|35531-3|LNC|Saccharum officinarum Ab.IgG|Saccharum officinarum Ab.IgG
C1507666|T201|COMP|35532-1|LNC|Chicken Ab.IgG|Chicken Ab.IgG
C1507667|T201|COMP|35533-9|LNC|Coffea spp Ab.IgG|Coffea spp Ab.IgG
C1507668|T201|COMP|35534-7|LNC|Zea mays Ab.IgG|Zea mays Ab.IgG
C1507674|T201|COMP|38230-9|LNC|Calcium.ionized|Calcium.ionized
C1507675|T201|COMP|38231-7|LNC|Cells.CD11b+HLA-DR+/100 cells|Cells.CD11b+HLA-DR+/100 cells
C1507676|T201|COMP|38232-5|LNC|Cells.CD13+CD16+/100 cells|Cells.CD13+CD16+/100 cells
C1507677|T201|COMP|38233-3|LNC|Cells.CD3+CD62L+|Cells.CD3+CD62L+
C1507678|T201|COMP|38234-1|LNC|Cells.CD3+CD62L+/100 cells|Cells.CD3+CD62L+/100 cells
C1507679|T201|COMP|38235-8|LNC|Cells.CD3+TCR gamma delta+|Cells.CD3+TCR gamma delta+
C1507680|T201|COMP|38236-6|LNC|Cells.CD3+TCR gamma delta+/100 cells|Cells.CD3+TCR gamma delta+/100 cells
C1507681|T201|COMP|38237-4|LNC|Cells.CD4+CD28+|Cells.CD4+CD28+
C1507682|T201|COMP|38238-2|LNC|Cells.CD4+CD28+/100 cells|Cells.CD4+CD28+/100 cells
C1507683|T201|COMP|38239-0|LNC|Cells.CD4+CD95+|Cells.CD4+CD95+
C1507684|T201|COMP|38240-8|LNC|Cells.CD4+CD95+/100 cells|Cells.CD4+CD95+/100 cells
C1507685|T201|COMP|38241-6|LNC|Cells.CD8+CD95+|Cells.CD8+CD95+
C1507686|T201|COMP|38242-4|LNC|Cells.CD8+CD95+/100 cells|Cells.CD8+CD95+/100 cells
C1507687|T201|COMP|38243-2|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C1507688|T201|COMP|38244-0|LNC|Brucella abortus Ab.IgM|Brucella abortus Ab.IgM
C1507689|T201|COMP|38245-7|LNC|Brucella canis Ab.IgG|Brucella canis Ab.IgG
C1507690|T201|COMP|38246-5|LNC|Brucella canis Ab.IgM|Brucella canis Ab.IgM
C1507691|T201|COMP|38247-3|LNC|Brucella sp Ab.IgG|Brucella sp Ab.IgG
C1507692|T201|COMP|38248-1|LNC|Brucella sp Ab.IgM|Brucella sp Ab.IgM
C1507693|T201|COMP|38249-9|LNC|C peptide^15M post XXX challenge|C peptide^15M post XXX challenge
C1507694|T201|COMP|38250-7|LNC|Calcium|Calcium
C1507695|T201|COMP|35535-4|LNC|Egg white Ab.IgG|Egg white Ab.IgG
C1507696|T201|COMP|35536-2|LNC|Egg yolk Ab.IgG|Egg yolk Ab.IgG
C1507697|T201|COMP|35537-0|LNC|Triticum aestivum Ab.IgG|Triticum aestivum Ab.IgG
C1507698|T201|COMP|35538-8|LNC|Saccharomyces cerevisiae Ab.IgG|Saccharomyces cerevisiae Ab.IgG
C1507699|T201|COMP|35539-6|LNC|Cow milk Ab.IgG|Cow milk Ab.IgG
C1507700|T201|COMP|35540-4|LNC|Agaricus hortensis Ab.IgG|Agaricus hortensis Ab.IgG
C1507701|T201|COMP|35541-2|LNC|Allium cepa Ab.IgG|Allium cepa Ab.IgG
C1507702|T201|COMP|35542-0|LNC|Arachis hypogaea Ab.IgG|Arachis hypogaea Ab.IgG
C1507703|T201|COMP|35543-8|LNC|Pork Ab.IgG|Pork Ab.IgG
C1507704|T201|COMP|35544-6|LNC|Solanum tuberosum Ab.IgG|Solanum tuberosum Ab.IgG
C1507705|T201|COMP|35545-3|LNC|Oryza sativa Ab.IgG|Oryza sativa Ab.IgG
C1507706|T201|COMP|35546-1|LNC|Glycine max Ab.IgG|Glycine max Ab.IgG
C1507707|T201|COMP|35547-9|LNC|Lycopersicon lycopersicum Ab.IgG|Lycopersicon lycopersicum Ab.IgG
C1507708|T201|COMP|35548-7|LNC|Fusarium moniliforme Ab.IgG|Fusarium moniliforme Ab.IgG
C1507709|T201|COMP|35549-5|LNC|Mucor racemosus Ab.IgG|Mucor racemosus Ab.IgG
C1507710|T201|COMP|35550-3|LNC|Phthalic anhydride Ab.IgG|Phthalic anhydride Ab.IgG
C1507711|T201|COMP|35551-1|LNC|Phoma betae Ab.IgG|Phoma betae Ab.IgG
C1507712|T201|COMP|35552-9|LNC|Rhizopus nigricans Ab.IgG|Rhizopus nigricans Ab.IgG
C1507713|T201|COMP|35553-7|LNC|Stemphylium botryosum Ab.IgG|Stemphylium botryosum Ab.IgG
C1507714|T201|COMP|35554-5|LNC|Chocolate Ab.IgG|Chocolate Ab.IgG
C1507715|T201|COMP|35555-2|LNC|Setomelanomma rostrata Ab.IgG|Setomelanomma rostrata Ab.IgG
C1507716|T201|COMP|35556-0|LNC|Trichophyton rubrum Ab.IgG|Trichophyton rubrum Ab.IgG
C1507717|T201|COMP|35557-8|LNC|Cladosporium cladosporioides Ab.IgG|Cladosporium cladosporioides Ab.IgG
C1507718|T201|COMP|35558-6|LNC|Cholinesterase panel|Cholinesterase panel
C1507719|T201|COMP|35559-4|LNC|Protein.monoclonal band 2|Protein.monoclonal band 2
C1507720|T201|COMP|35560-2|LNC|Protein.monoclonal|Protein.monoclonal
C1507721|T201|COMP|35561-0|LNC|Protein.monoclonal band 2|Protein.monoclonal band 2
C1507722|T201|COMP|35562-8|LNC|Bile acid^post CFst|Bile acid^post CFst
C1507723|T201|COMP|35563-6|LNC|Rickettsia rickettsii Ab.IgG & IgM panel|Rickettsia rickettsii Ab.IgG & IgM panel
C1507724|T201|COMP|35564-4|LNC|HIV 1 p31+p32 Ab|HIV 1 p31+p32 Ab
C1507725|T201|COMP|35565-1|LNC|HIV 1 p40 Ab|HIV 1 p40 Ab
C1507726|T201|COMP|35566-9|LNC|Parathyrin^baseline|Parathyrin^baseline
C1507727|T201|COMP|35567-7|LNC|Parathyrin^10M post excision|Parathyrin^10M post excision
C1507728|T201|COMP|35568-5|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C1507729|T201|COMP|35569-3|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C1507730|T201|COMP|35570-1|LNC|Renin|Renin
C1507731|T201|COMP|35571-9|LNC|Tyrosine|Tyrosine
C1507732|T201|COMP|35572-7|LNC|Phenylalanine/Tyrosine|Phenylalanine/Tyrosine
C1507733|T201|COMP|35573-5|LNC|Procollagen+Collagen|Procollagen+Collagen
C1507734|T201|COMP|35574-3|LNC|Fatty acid oxidation|Fatty acid oxidation
C1507735|T201|COMP|35575-0|LNC|Pigeon antibody panel|Pigeon antibody panel
C1507736|T201|COMP|35576-8|LNC|Hydrocarbon and oxygenated volatiles panel|Hydrocarbon and oxygenated volatiles panel
C1507737|T201|COMP|35577-6|LNC|Hypersensitivity pneumonitis panel|Hypersensitivity pneumonitis panel
C1507738|T201|COMP|35578-4|LNC|1,2-Glyceryl dinitrate|1,2-Glyceryl dinitrate
C1507739|T201|COMP|35579-2|LNC|Tetrahydrofuran|Tetrahydrofuran
C1507740|T201|COMP|35580-0|LNC|N-methyl valine|N-methyl valine
C1507741|T201|COMP|35581-8|LNC|Hydroxyethyl valine|Hydroxyethyl valine
C1507742|T201|COMP|35582-6|LNC|Hydrazine|Hydrazine
C1507743|T201|COMP|35583-4|LNC|Hydrazine/Creatinine|Hydrazine/Creatinine
C1507744|T201|COMP|35584-2|LNC|Aniline|Aniline
C1507745|T201|COMP|35585-9|LNC|2-Butoxyacetate|2-Butoxyacetate
C1507746|T201|COMP|35586-7|LNC|4-Tert-Butylphenol|4-Tert-Butylphenol
C1507747|T201|COMP|35587-5|LNC|2-Ethoxyacetate|2-Ethoxyacetate
C1507748|T201|COMP|35588-3|LNC|Ethylene glycol dinitrate|Ethylene glycol dinitrate
C1507749|T201|COMP|35589-1|LNC|Furoate/Creatinine|Furoate/Creatinine
C1507750|T201|COMP|35590-9|LNC|Aniline|Aniline
C1507751|T201|COMP|35591-7|LNC|Creatinine renal clearance.predicted|Creatinine renal clearance.predicted
C1507752|T201|COMP|35592-5|LNC|Creatinine renal clearance/1.73 sq M.predicted|Creatinine renal clearance/1.73 sq M.predicted
C1507753|T201|COMP|35593-3|LNC|Creatinine renal clearance/1.73 sq M|Creatinine renal clearance/1.73 sq M
C1507754|T201|COMP|35594-1|LNC|Creatinine renal clearance/1.73 sq M|Creatinine renal clearance/1.73 sq M
C1507755|T201|COMP|35595-8|LNC|Acetaminophen|Acetaminophen
C1507756|T201|COMP|35596-6|LNC|Theophylline|Theophylline
C1507757|T201|COMP|35597-4|LNC|Salicylates|Salicylates
C1507758|T201|COMP|35598-2|LNC|Butalbital|Butalbital
C1507759|T201|COMP|35599-0|LNC|carBAMazepine|carBAMazepine
C1507760|T201|COMP|35600-6|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C1507761|T201|COMP|35601-4|LNC|chlorproMAZINE|chlorproMAZINE
C1507762|T201|COMP|35602-2|LNC|clomiPRAMINE|clomiPRAMINE
C1507763|T201|COMP|35603-0|LNC|clonazePAM|clonazePAM
C1507764|T201|COMP|35604-8|LNC|Cyclobenzaprine|Cyclobenzaprine
C1507765|T201|COMP|35605-5|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C1507766|T201|COMP|35606-3|LNC|Desipramine|Desipramine
C1507767|T201|COMP|35607-1|LNC|diazePAM|diazePAM
C1507768|T201|COMP|35608-9|LNC|diphenhydrAMINE|diphenhydrAMINE
C1507769|T201|COMP|35609-7|LNC|Doxepin|Doxepin
C1507770|T201|COMP|35610-5|LNC|FLUoxetine|FLUoxetine
C1507771|T201|COMP|35611-3|LNC|Flurazepam|Flurazepam
C1507772|T201|COMP|35612-1|LNC|fluvoxaMINE|fluvoxaMINE
C1507773|T201|COMP|35613-9|LNC|Glutethimide|Glutethimide
C1507774|T201|COMP|35614-7|LNC|Ibuprofen|Ibuprofen
C1507775|T201|COMP|35615-4|LNC|Lidocaine|Lidocaine
C1507776|T201|COMP|35616-2|LNC|LORazepam|LORazepam
C1507777|T201|COMP|35617-0|LNC|Meperidine|Meperidine
C1507778|T201|COMP|35626-1|LNC|Norpropoxyphene|Norpropoxyphene
C1507779|T201|COMP|35627-9|LNC|Nortriptyline|Nortriptyline
C1507780|T201|COMP|35628-7|LNC|Norverapamil|Norverapamil
C1507781|T201|COMP|35629-5|LNC|Oxazepam|Oxazepam
C1507782|T201|COMP|35630-3|LNC|PENTobarbital|PENTobarbital
C1507783|T201|COMP|35631-1|LNC|PHENobarbital|PHENobarbital
C1507784|T201|COMP|35632-9|LNC|Phenytoin|Phenytoin
C1507785|T201|COMP|35633-7|LNC|Propranolol|Propranolol
C1507786|T201|COMP|35634-5|LNC|Secobarbital|Secobarbital
C1507787|T201|COMP|35635-2|LNC|traZODone|traZODone
C1507788|T201|COMP|35636-0|LNC|Amitriptyline|Amitriptyline
C1507789|T201|COMP|35637-8|LNC|4-Hydroxyglutethimide|4-Hydroxyglutethimide
C1507790|T201|COMP|35638-6|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C1507792|T201|COMP|35640-2|LNC|Cells.CD5/100 cells|Cells.CD5/100 cells
C1507793|T201|COMP|35641-0|LNC|Cells.CD7/100 cells|Cells.CD7/100 cells
C1507794|T201|COMP|35642-8|LNC|Cotinine|Cotinine
C1507795|T201|COMP|35643-6|LNC|Collagen type 2 Ab|Collagen type 2 Ab
C1507796|T201|COMP|35645-1|LNC|NSD1 gene deletion|NSD1 gene deletion
C1507797|T201|COMP|35646-9|LNC|Deoxypyridinoline/Creatinine|Deoxypyridinoline/Creatinine
C1507798|T201|COMP|35647-7|LNC|Pyridinoline+Deoxypyridinoline/Creatinine|Pyridinoline+Deoxypyridinoline/Creatinine
C1507799|T201|COMP|35648-5|LNC|C reactive protein|C reactive protein
C1507800|T201|COMP|35649-3|LNC|Propoxyphene|Propoxyphene
C1507802|T201|COMP|35651-9|LNC|Synovial lining cells/100 cells|Synovial lining cells/100 cells
C1507803|T201|COMP|35652-7|LNC|Epithelial cells/100 cells|Epithelial cells/100 cells
C1507804|T201|COMP|35653-5|LNC|Cells.CD158|Cells.CD158
C1507805|T201|COMP|35654-3|LNC|Creatinine/body weight|Creatinine/body weight
C1507806|T201|COMP|35655-0|LNC|Butyrylcarnitine (C4)|Butyrylcarnitine (C4)
C1507807|T201|COMP|35656-8|LNC|3-Hydroxystearoylcarnitine (C18-OH)|3-Hydroxystearoylcarnitine (C18-OH)
C1507808|T201|COMP|35657-6|LNC|Urea nitrogen/body weight|Urea nitrogen/body weight
C1507812|T201|COMP|35661-8|LNC|JC virus DNA|JC virus DNA
C1507813|T201|COMP|35662-6|LNC|Glucose|Glucose
C1507814|T201|COMP|35663-4|LNC|Protein|Protein
C1507815|T201|COMP|35664-2|LNC|Ethanol|Ethanol
C1507816|T201|COMP|35665-9|LNC|Acetone|Acetone
C1507818|T201|COMP|35667-5|LNC|Atomoxetine|Atomoxetine
C1507819|T201|COMP|35668-3|LNC|Gentamicin|Gentamicin
C1507820|T201|COMP|35669-1|LNC|Amikacin|Amikacin
C1507821|T201|COMP|35670-9|LNC|Tobramycin|Tobramycin
C1507822|T201|COMP|35671-7|LNC|Galactomannan Ag|Galactomannan Ag
C1507824|T201|COMP|35673-3|LNC|Phosphate|Phosphate
C1507825|T201|COMP|35674-1|LNC|Creatinine|Creatinine
C1507826|T201|COMP|35675-8|LNC|Calcium|Calcium
C1507827|T201|COMP|35676-6|LNC|Chloride|Chloride
C1507828|T201|COMP|35677-4|LNC|Potassium|Potassium
C1507829|T201|COMP|35678-2|LNC|Sodium|Sodium
C1507830|T201|COMP|35679-0|LNC|Varicella zoster virus Ab.IgG & IgM panel|Varicella zoster virus Ab.IgG & IgM panel
C1507831|T201|COMP|35680-8|LNC|Hepatitis E virus Ab.IgG & IgM panel|Hepatitis E virus Ab.IgG & IgM panel
C1507832|T201|COMP|35681-6|LNC|Tissue transglutaminase Ab panel|Tissue transglutaminase Ab panel
C1507833|T201|COMP|35682-4|LNC|Trypanosoma cruzi Ab.IgG & IgM panel|Trypanosoma cruzi Ab.IgG & IgM panel
C1507834|T201|COMP|35683-2|LNC|Burkholderia pseudomallei Ab.IgG & IgM panel|Burkholderia pseudomallei Ab.IgG & IgM panel
C1507835|T201|COMP|35684-0|LNC|Colorado tick fever virus Ab.IgG & IgM panel|Colorado tick fever virus Ab.IgG & IgM panel
C1507836|T201|COMP|35685-7|LNC|Carbon dioxide|Carbon dioxide
C1507837|T201|COMP|35686-5|LNC|GBA gene.c.1226A>G|GBA gene.c.1226A>G
C1507838|T201|COMP|35687-3|LNC|GBA gene.c.1297G>T|GBA gene.c.1297G>T
C1507839|T201|COMP|35688-1|LNC|GBA gene.c.1448T>G & 1448T>C|GBA gene.c.1448T>G & 1448T>C
C1507840|T201|COMP|35689-9|LNC|GBA gene.c.84insG|GBA gene.c.84insG
C1507841|T201|COMP|35690-7|LNC|GBA gene.c.IVS2(+1)G>A & IVS2(+1)G>T|GBA gene.c.IVS2(+1)G>A & IVS2(+1)G>T
C1507842|T201|COMP|35691-5|LNC|XXX microorganism DNA|XXX microorganism DNA
C1507843|T201|COMP|35692-3|LNC|Cells.G0+G1 phase/100 cells|Cells.G0+G1 phase/100 cells
C1507844|T201|COMP|35693-1|LNC|GBA gene targeted mutation analysis|GBA gene targeted mutation analysis
C1507845|T201|COMP|35694-9|LNC|California encephalitis virus Ab.IgG|California encephalitis virus Ab.IgG
C1507846|T201|COMP|35695-6|LNC|California encephalitis virus Ab.IgM|California encephalitis virus Ab.IgM
C1507847|T201|COMP|35696-4|LNC|California encephalitis virus Ab|California encephalitis virus Ab
C1507848|T201|COMP|35697-2|LNC|La Crosse virus Ab|La Crosse virus Ab
C1507849|T201|COMP|35698-0|LNC|metFORMIN|metFORMIN
C1507850|T201|COMP|35699-8|LNC|Anti-hyperglycemics|Anti-hyperglycemics
C1507851|T201|COMP|35700-4|LNC|Acetaminophen|Acetaminophen
C1507852|T201|COMP|35701-2|LNC|Acetylcholinesterase|Acetylcholinesterase
C1507853|T201|COMP|35702-0|LNC|Acid hemolysis|Acid hemolysis
C1507854|T201|COMP|35703-8|LNC|Adenosine deaminase|Adenosine deaminase
C1507855|T201|COMP|35704-6|LNC|Adenosine deaminase|Adenosine deaminase
C1507856|T201|COMP|35705-3|LNC|Adenovirus Ag|Adenovirus Ag
C1507857|T201|COMP|35706-1|LNC|Albumin/Protein.total|Albumin/Protein.total
C1507859|T201|COMP|35708-7|LNC|Alpha 1 globulin|Alpha 1 globulin
C1507860|T201|COMP|35709-5|LNC|La Crosse virus Ab|La Crosse virus Ab
C1507861|T201|COMP|35710-3|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507862|T201|COMP|35711-1|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507863|T201|COMP|35712-9|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507864|T201|COMP|35713-7|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507865|T201|COMP|35714-5|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507866|T201|COMP|35715-2|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507867|T201|COMP|35716-0|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507868|T201|COMP|35717-8|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507869|T201|COMP|35718-6|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507870|T201|COMP|35719-4|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507871|T201|COMP|35720-2|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507872|T201|COMP|35721-0|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507873|T201|COMP|35722-8|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507874|T201|COMP|35723-6|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507875|T201|COMP|35724-4|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507876|T201|COMP|35725-1|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507877|T201|COMP|35726-9|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507878|T201|COMP|35727-7|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507879|T201|COMP|35728-5|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507880|T201|COMP|35729-3|LNC|Chlamydia sp DNA|Chlamydia sp DNA
C1507881|T201|COMP|35730-1|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507882|T201|COMP|35731-9|LNC|Corylus avellana Ab.IgG.RAST class|Corylus avellana Ab.IgG.RAST class
C1507883|T201|COMP|35732-7|LNC|Histoplasma capsulatum H Ab|Histoplasma capsulatum H Ab
C1507884|T201|COMP|35733-5|LNC|Histoplasma capsulatum M Ab|Histoplasma capsulatum M Ab
C1507885|T201|COMP|35734-3|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1507886|T201|COMP|35735-0|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C1507887|T201|COMP|35736-8|LNC|Chlamydia sp rRNA|Chlamydia sp rRNA
C1507889|T201|COMP|35738-4|LNC|Inhibin A|Inhibin A
C1507890|T201|COMP|35739-2|LNC|Brucella sp Ab.IgG & IgM panel|Brucella sp Ab.IgG & IgM panel
C1507891|T201|COMP|35740-0|LNC|Rickettsia sp Ab.IgG & IgM panel|Rickettsia sp Ab.IgG & IgM panel
C1507892|T201|COMP|35741-8|LNC|Prostate specific Ag|Prostate specific Ag
C1507893|T201|COMP|35742-6|LNC|SH2D1A gene targeted mutation analysis|SH2D1A gene targeted mutation analysis
C1507895|T201|COMP|35744-2|LNC|TP73L gene targeted mutation analysis|TP73L gene targeted mutation analysis
C1507896|T201|COMP|35745-9|LNC|Fat/Solids.total|Fat/Solids.total
C1507897|T201|COMP|35746-7|LNC|Hyperchromia|Hyperchromia
C1507898|T201|COMP|35747-5|LNC|Hydrogen ion|Hydrogen ion
C1507900|T201|COMP|35749-1|LNC|DMPK phenotype|DMPK phenotype
C1507901|T201|COMP|35750-9|LNC|DMPK gene allele 2.CTG repeats|DMPK gene allele 2.CTG repeats
C1507902|T201|COMP|35751-7|LNC|DMPK gene allele 1.CTG repeats|DMPK gene allele 1.CTG repeats
C1507903|T201|COMP|35752-5|LNC|Escherichia coli O157:H7 Ab.IgG & IgM panel|Escherichia coli O157:H7 Ab.IgG & IgM panel
C1507905|T201|COMP|35754-1|LNC|Avilamycin|Avilamycin
C1507906|T201|COMP|35755-8|LNC|Avilamycin|Avilamycin
C1507907|T201|COMP|35756-6|LNC|Avilamycin|Avilamycin
C1507908|T201|COMP|35757-4|LNC|Cefdinir|Cefdinir
C1507909|T201|COMP|35758-2|LNC|Cefdinir|Cefdinir
C1507910|T201|COMP|35759-0|LNC|Cefditoren|Cefditoren
C1507911|T201|COMP|35760-8|LNC|Cefditoren|Cefditoren
C1507912|T201|COMP|35761-6|LNC|Cefditoren|Cefditoren
C1507913|T201|COMP|35762-4|LNC|Cefditoren|Cefditoren
C1507914|T201|COMP|35763-2|LNC|Cefepime+Clavulanate|Cefepime+Clavulanate
C1507915|T201|COMP|35764-0|LNC|Cefetamet|Cefetamet
C1507916|T201|COMP|35765-7|LNC|Cefetamet|Cefetamet
C1507917|T201|COMP|35766-5|LNC|Cefixime|Cefixime
C1507918|T201|COMP|35767-3|LNC|Cefoperazone|Cefoperazone
C1507919|T201|COMP|35768-1|LNC|Cefoperazone+Sulbactam|Cefoperazone+Sulbactam
C1507920|T201|COMP|35769-9|LNC|Cefotaxime+Clavulanate|Cefotaxime+Clavulanate
C1507921|T201|COMP|35770-7|LNC|Cefotaxime+Clavulanate|Cefotaxime+Clavulanate
C1507922|T201|COMP|35771-5|LNC|Cefotaxime+Clavulanate|Cefotaxime+Clavulanate
C1507923|T201|COMP|35772-3|LNC|Cefotiam|Cefotiam
C1507924|T201|COMP|35773-1|LNC|Cefotiam|Cefotiam
C1507925|T201|COMP|35774-9|LNC|cefTAZidime+Clavulanate|cefTAZidime+Clavulanate
C1507926|T201|COMP|35775-6|LNC|cefTAZidime+Clavulanate|cefTAZidime+Clavulanate
C1507927|T201|COMP|35776-4|LNC|cefTAZidime+Clavulanate|cefTAZidime+Clavulanate
C1507928|T201|COMP|35777-2|LNC|Ceftibuten|Ceftibuten
C1507929|T201|COMP|35778-0|LNC|Ceftibuten|Ceftibuten
C1507930|T201|COMP|35779-8|LNC|Ceftibuten|Ceftibuten
C1507931|T201|COMP|35780-6|LNC|Ceftiofur|Ceftiofur
C1507932|T201|COMP|35781-4|LNC|Ceftiofur|Ceftiofur
C1507933|T201|COMP|35782-2|LNC|Cefuroxime.oral|Cefuroxime.oral
C1507934|T201|COMP|35783-0|LNC|Cefuroxime.oral|Cefuroxime.oral
C1507935|T201|COMP|35784-8|LNC|Cephalexin|Cephalexin
C1507936|T201|COMP|35785-5|LNC|Clinafloxacin|Clinafloxacin
C1507937|T201|COMP|35786-3|LNC|Clinafloxacin|Clinafloxacin
C1507938|T201|COMP|35787-1|LNC|DAPTOmycin|DAPTOmycin
C1507939|T201|COMP|35788-9|LNC|DAPTOmycin|DAPTOmycin
C1507940|T201|COMP|35789-7|LNC|DAPTOmycin|DAPTOmycin
C1507941|T201|COMP|35790-5|LNC|Difloxacin|Difloxacin
C1507942|T201|COMP|35791-3|LNC|Difloxacin|Difloxacin
C1507943|T201|COMP|35792-1|LNC|Difloxacin|Difloxacin
C1507944|T201|COMP|35793-9|LNC|Dirithromycin|Dirithromycin
C1507945|T201|COMP|35794-7|LNC|Dirithromycin|Dirithromycin
C1507946|T201|COMP|35795-4|LNC|Dirithromycin|Dirithromycin
C1507947|T201|COMP|35796-2|LNC|Enrofloxacin|Enrofloxacin
C1507948|T201|COMP|35797-0|LNC|Enrofloxacin|Enrofloxacin
C1507949|T201|COMP|35798-8|LNC|Enrofloxacin|Enrofloxacin
C1507950|T201|COMP|35799-6|LNC|Ertapenem|Ertapenem
C1507951|T201|COMP|35800-2|LNC|Ertapenem|Ertapenem
C1507952|T201|COMP|35801-0|LNC|Ertapenem|Ertapenem
C1507953|T201|COMP|35802-8|LNC|Ertapenem|Ertapenem
C1507954|T201|COMP|35803-6|LNC|Bambermycins|Bambermycins
C1507955|T201|COMP|35804-4|LNC|Bambermycins|Bambermycins
C1507956|T201|COMP|35805-1|LNC|Bambermycins|Bambermycins
C1507957|T201|COMP|35806-9|LNC|Fleroxacin|Fleroxacin
C1507958|T201|COMP|35807-7|LNC|Florfenicol|Florfenicol
C1507959|T201|COMP|35808-5|LNC|Florfenicol|Florfenicol
C1507960|T201|COMP|35809-3|LNC|Fosfomycin|Fosfomycin
C1507961|T201|COMP|35810-1|LNC|Fosfomycin|Fosfomycin
C1507962|T201|COMP|35811-9|LNC|Garenoxacin|Garenoxacin
C1507963|T201|COMP|35820-0|LNC|Isepamicin|Isepamicin
C1507964|T201|COMP|35821-8|LNC|Isepamicin|Isepamicin
C1507965|T201|COMP|35822-6|LNC|Mupirocin|Mupirocin
C1507966|T201|COMP|35823-4|LNC|Mupirocin|Mupirocin
C1507967|T201|COMP|35824-2|LNC|Nystatin|Nystatin
C1507968|T201|COMP|35825-9|LNC|Orbifloxacin|Orbifloxacin
C1507969|T201|COMP|35826-7|LNC|Orbifloxacin|Orbifloxacin
C1507970|T201|COMP|35827-5|LNC|Orbifloxacin|Orbifloxacin
C1507971|T201|COMP|35828-3|LNC|Pefloxacin|Pefloxacin
C1507972|T201|COMP|35829-1|LNC|Pirlimycin|Pirlimycin
C1507973|T201|COMP|35830-9|LNC|Pirlimycin|Pirlimycin
C1507974|T201|COMP|35831-7|LNC|Pirlimycin|Pirlimycin
C1507975|T201|COMP|35832-5|LNC|Polymyxin B|Polymyxin B
C1507976|T201|COMP|35833-3|LNC|Pristinamycin|Pristinamycin
C1507977|T201|COMP|35834-1|LNC|Pristinamycin|Pristinamycin
C1507978|T201|COMP|35835-8|LNC|Quinupristin+Dalfopristin|Quinupristin+Dalfopristin
C1507979|T201|COMP|35836-6|LNC|Salinomycin|Salinomycin
C1507980|T201|COMP|35837-4|LNC|Salinomycin|Salinomycin
C1507981|T201|COMP|35838-2|LNC|Salinomycin|Salinomycin
C1507982|T201|COMP|35839-0|LNC|Sparfloxacin|Sparfloxacin
C1507983|T201|COMP|35840-8|LNC|Spectinomycin|Spectinomycin
C1507984|T201|COMP|35841-6|LNC|Streptomycin.high potency|Streptomycin.high potency
C1507985|T201|COMP|35842-4|LNC|Sulfonamide|Sulfonamide
C1507986|T201|COMP|35843-2|LNC|Telithromycin|Telithromycin
C1507987|T201|COMP|35844-0|LNC|Telithromycin|Telithromycin
C1507988|T201|COMP|35845-7|LNC|Telithromycin|Telithromycin
C1507989|T201|COMP|35846-5|LNC|Tiamulin|Tiamulin
C1507990|T201|COMP|35847-3|LNC|Tiamulin|Tiamulin
C1507991|T201|COMP|35848-1|LNC|Tiamulin|Tiamulin
C1507992|T201|COMP|35849-9|LNC|Tilmicosin|Tilmicosin
C1507993|T201|COMP|35850-7|LNC|Tilmicosin|Tilmicosin
C1507994|T201|COMP|35851-5|LNC|Tilmicosin|Tilmicosin
C1507995|T201|COMP|35852-3|LNC|Trospectinomycin|Trospectinomycin
C1507996|T201|COMP|35853-1|LNC|Trospectinomycin|Trospectinomycin
C1507997|T201|COMP|35854-9|LNC|Trospectinomycin|Trospectinomycin
C1507998|T201|COMP|35855-6|LNC|Trovafloxacin|Trovafloxacin
C1507999|T201|COMP|35856-4|LNC|Tylosin|Tylosin
C1508000|T201|COMP|35857-2|LNC|Tylosin|Tylosin
C1508001|T201|COMP|35858-0|LNC|Tylosin|Tylosin
C1508002|T201|COMP|35868-9|LNC|2-Oxoisovalerate|2-Oxoisovalerate
C1508003|T201|COMP|35869-7|LNC|2-Oxo,3-Methylvalerate|2-Oxo,3-Methylvalerate
C1508004|T201|COMP|35870-5|LNC|2-Oxoisocaproate|2-Oxoisocaproate
C1508005|T201|COMP|35871-3|LNC|Succinate|Succinate
C1508006|T201|COMP|35872-1|LNC|Penicillin+Novobiocin|Penicillin+Novobiocin
C1508007|T201|COMP|35873-9|LNC|Penicillin+Novobiocin|Penicillin+Novobiocin
C1508008|T201|COMP|35874-7|LNC|Penicillin+Novobiocin|Penicillin+Novobiocin
C1508009|T201|COMP|35875-4|LNC|Herpes simplex virus 1+2 Ab|Herpes simplex virus 1+2 Ab
C1508010|T201|COMP|35876-2|LNC|Rickettsia sp Ab.IgM|Rickettsia sp Ab.IgM
C1508011|T201|COMP|35877-0|LNC|Rickettsia sp Ab.IgG|Rickettsia sp Ab.IgG
C1508012|T201|COMP|35878-8|LNC|Escherichia coli O157:H7 Ab.IgM|Escherichia coli O157:H7 Ab.IgM
C1508013|T201|COMP|35879-6|LNC|Escherichia coli O157:H7 Ab.IgG|Escherichia coli O157:H7 Ab.IgG
C1508014|T201|COMP|35880-4|LNC|Tissue transglutaminase Ab.IgM|Tissue transglutaminase Ab.IgM
C1508015|T201|COMP|36895-1|LNC|Arbovirus Ab|Arbovirus Ab
C1508016|T201|COMP|36896-9|LNC|West Nile virus polyvalent E Ab|West Nile virus polyvalent E Ab
C1508037|T201|COMP|36897-7|LNC|West Nile virus Ab|West Nile virus Ab
C1508038|T201|COMP|36898-5|LNC|West Nile virus NS5 Ab|West Nile virus NS5 Ab
C1508039|T201|COMP|36899-3|LNC|Arbovirus Ab|Arbovirus Ab
C1508040|T201|COMP|36900-9|LNC|West Nile virus polyvalent E Ab|West Nile virus polyvalent E Ab
C1508041|T201|COMP|36901-7|LNC|West Nile virus NS5 Ab|West Nile virus NS5 Ab
C1508042|T201|COMP|36902-5|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae DNA|Chlamydia trachomatis+Neisseria gonorrhoeae DNA
C1508043|T201|COMP|36903-3|LNC|Chlamydia trachomatis & Neisseria gonorrhoeae DNA|Chlamydia trachomatis & Neisseria gonorrhoeae DNA
C1508044|T201|COMP|36904-1|LNC|Inhibin A^^adjusted|Inhibin A^^adjusted
C1508045|T201|COMP|36905-8|LNC|Inhibin A^^unadjusted|Inhibin A^^unadjusted
C1508046|T201|COMP|36906-6|LNC|Complement C1 esterase inhibitor|Complement C1 esterase inhibitor
C1508047|T201|COMP|36907-4|LNC|Chromosome 8 trisomy|Chromosome 8 trisomy
C1508048|T201|COMP|36908-2|LNC|Gene mutations tested for|Gene mutations tested for
C1508049|T201|COMP|36909-0|LNC|Cells.G0+G1 phase/100 cells|Cells.G0+G1 phase/100 cells
C1508050|T201|COMP|36910-8|LNC|Cells.S phase/100 cells|Cells.S phase/100 cells
C1508052|T201|COMP|36912-4|LNC|CATCH22 syndrome gene mutations tested for|CATCH22 syndrome gene mutations tested for
C1508053|T201|COMP|36913-2|LNC|FMR1 gene targeted mutation analysis|FMR1 gene targeted mutation analysis
C1508054|T201|COMP|36914-0|LNC|FMR1 gene mutations tested for|FMR1 gene mutations tested for
C1508055|T201|COMP|36915-7|LNC|AS+PWS gene mutations tested for|AS+PWS gene mutations tested for
C1508056|T201|COMP|36916-5|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C1508057|T201|COMP|36917-3|LNC|Chromosome uniparental disomy|Chromosome uniparental disomy
C1508058|T201|COMP|36918-1|LNC|ALDOB gene targeted mutation analysis|ALDOB gene targeted mutation analysis
C1508059|T201|COMP|36919-9|LNC|ELN gene mutations tested for|ELN gene mutations tested for
C1508060|T201|COMP|36920-7|LNC|PROP1 gene targeted mutation analysis|PROP1 gene targeted mutation analysis
C1508061|T201|COMP|36921-5|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C1508062|T201|COMP|36922-3|LNC|TPMT gene targeted mutation analysis|TPMT gene targeted mutation analysis
C1508063|T201|COMP|36923-1|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1508064|T201|COMP|36924-9|LNC|14-3-3 Ag|14-3-3 Ag
C1508065|T201|COMP|36925-6|LNC|MEFV gene targeted mutation analysis|MEFV gene targeted mutation analysis
C1508066|T201|COMP|37424-9|LNC|Perchlorate|Perchlorate
C1508067|T201|COMP|37425-6|LNC|Prion protein.abnormal|Prion protein.abnormal
C1508068|T201|COMP|37982-6|LNC|Avian paramyxovirus|Avian paramyxovirus
C1508069|T201|COMP|37983-4|LNC|Eastern equine encephalitis virus RNA|Eastern equine encephalitis virus RNA
C1508070|T201|COMP|37984-2|LNC|Saint Louis encephalitis virus RNA|Saint Louis encephalitis virus RNA
C1508071|T201|COMP|37985-9|LNC|West Nile virus RNA|West Nile virus RNA
C1508072|T201|COMP|37986-7|LNC|California serogroup virus RNA|California serogroup virus RNA
C1508076|T201|COMP|37990-9|LNC|Corticotropin releasing hormone|Corticotropin releasing hormone
C1508077|T201|COMP|37991-7|LNC|Neutrophil cytoplasmic Ab.perinuclear|Neutrophil cytoplasmic Ab.perinuclear
C1508078|T201|COMP|37992-5|LNC|Neutrophil cytoplasmic Ab.classic|Neutrophil cytoplasmic Ab.classic
C1508079|T201|COMP|37993-3|LNC|DNA double strand Ab|DNA double strand Ab
C1508089|T201|COMP|38157-4|LNC|Parathyrin.intact^5M post excision|Parathyrin.intact^5M post excision
C1508090|T201|COMP|38158-2|LNC|Parathyrin.intact^baseline|Parathyrin.intact^baseline
C1508091|T201|COMP|38159-0|LNC|levETIRAcetam|levETIRAcetam
C1508092|T201|COMP|38160-8|LNC|Porphyrins/Creatinine|Porphyrins/Creatinine
C1508093|T201|COMP|38161-6|LNC|Pentacarboxylporphyrins/Creatinine|Pentacarboxylporphyrins/Creatinine
C1508094|T201|COMP|38162-4|LNC|Coproporphyrin/Creatinine|Coproporphyrin/Creatinine
C1508095|T201|COMP|38163-2|LNC|Heptacarboxylporphyrin/Creatinine|Heptacarboxylporphyrin/Creatinine
C1508096|T201|COMP|38164-0|LNC|Hexacarboxylporphyrin/Creatinine|Hexacarboxylporphyrin/Creatinine
C1508097|T201|COMP|38165-7|LNC|Uroporphyrin/Creatinine|Uroporphyrin/Creatinine
C1508098|T201|COMP|38166-5|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1508099|T201|COMP|38167-3|LNC|Major crossmatch|Major crossmatch
C1508100|T201|COMP|38168-1|LNC|Major crossmatch|Major crossmatch
C1508101|T201|COMP|38169-9|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C1508102|T201|COMP|38170-7|LNC|Cells.CD18/100 cells|Cells.CD18/100 cells
C1508103|T201|COMP|38171-5|LNC|Cells.CD3-CD19+/100 cells|Cells.CD3-CD19+/100 cells
C1508104|T201|COMP|38172-3|LNC|Organic acids|Organic acids
C1508105|T201|COMP|38173-1|LNC|Borrelia burgdorferi C6 Ab|Borrelia burgdorferi C6 Ab
C1508106|T201|COMP|38174-9|LNC|Borrelia burgdorferi C6 Ab|Borrelia burgdorferi C6 Ab
C1508107|T201|COMP|38175-6|LNC|Heptacarboxylate/Creatinine|Heptacarboxylate/Creatinine
C1508108|T201|COMP|38176-4|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C1508109|T201|COMP|38177-2|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C1508110|T201|COMP|38178-0|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C1508112|T201|COMP|38180-6|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1508113|T201|COMP|38182-2|LNC|Parainfluenza virus 1 Ab.IgG|Parainfluenza virus 1 Ab.IgG
C1508114|T201|COMP|38183-0|LNC|Parainfluenza virus 2 Ab.IgG|Parainfluenza virus 2 Ab.IgG
C1508115|T201|COMP|38184-8|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1508116|T201|COMP|38185-5|LNC|Beta galactosidase|Beta galactosidase
C1508117|T201|COMP|38186-3|LNC|Beta globulin|Beta globulin
C1508118|T201|COMP|38187-1|LNC|Bile acid.dihydroxy|Bile acid.dihydroxy
C1508119|T201|COMP|38188-9|LNC|Bile acid.trihydroxy|Bile acid.trihydroxy
C1508120|T201|COMP|38189-7|LNC|Alpha 2 globulin|Alpha 2 globulin
C1508121|T201|COMP|38190-5|LNC|Alpha 2 globulin|Alpha 2 globulin
C1508122|T201|COMP|38191-3|LNC|Ammonium urate/Total|Ammonium urate/Total
C1508123|T201|COMP|38192-1|LNC|Amylase|Amylase
C1508124|T201|COMP|38193-9|LNC|Amylase|Amylase
C1508125|T201|COMP|38194-7|LNC|Antidepressants|Antidepressants
C1508126|T201|COMP|38195-4|LNC|Antihistamines|Antihistamines
C1508127|T201|COMP|38196-2|LNC|Appearance|Appearance
C1508128|T201|COMP|38197-0|LNC|Bordetella parapertussis Ag|Bordetella parapertussis Ag
C1508129|T201|COMP|38198-8|LNC|Bordetella pertussis Ag|Bordetella pertussis Ag
C1508131|T201|COMP|38200-2|LNC|Specimen volume|Specimen volume
C1508136|T201|COMP|38251-5|LNC|Calcium oxalate|Calcium oxalate
C1508137|T201|COMP|38252-3|LNC|Calcium oxalate monohydrate/Total|Calcium oxalate monohydrate/Total
C1508138|T201|COMP|38253-1|LNC|Carbon dioxide|Carbon dioxide
C1508139|T201|COMP|38254-9|LNC|Carbonated calcium phosphate|Carbonated calcium phosphate
C1508140|T201|COMP|38255-6|LNC|Cat dander Ab.IgE/IgE.total|Cat dander Ab.IgE/IgE.total
C1508141|T201|COMP|38256-4|LNC|Cells counted.total|Cells counted.total
C1508142|T201|COMP|38257-2|LNC|Cells counted.total|Cells counted.total
C1508143|T201|COMP|38258-0|LNC|Cells counted.total|Cells counted.total
C1508144|T201|COMP|38259-8|LNC|Cells counted.total|Cells counted.total
C1508145|T201|COMP|38260-6|LNC|Cells counted.total|Cells counted.total
C1508146|T201|COMP|38270-5|LNC|Influenza virus A H7 RNA|Influenza virus A H7 RNA
C1508147|T201|COMP|38271-3|LNC|Influenza virus A H6 RNA|Influenza virus A H6 RNA
C1508148|T201|COMP|38272-1|LNC|Influenza virus A H5 RNA|Influenza virus A H5 RNA
C1508149|T201|COMP|38273-9|LNC|Influenza virus A Ab|Influenza virus A Ab
C1508150|T201|COMP|38274-7|LNC|Columbid circovirus DNA|Columbid circovirus DNA
C1508151|T201|COMP|38275-4|LNC|Transmissible spongiform encephalopathy|Transmissible spongiform encephalopathy
C1508152|T201|COMP|38276-2|LNC|Coagulation surface induced^1H post incubation|Coagulation surface induced^1H post incubation
C1508161|T201|COMP|38285-3|LNC|Erythrocytes|Erythrocytes
C1508162|T201|COMP|38286-1|LNC|2,4-Dichlorophenoxyacetate|2,4-Dichlorophenoxyacetate
C1508163|T201|COMP|38287-9|LNC|2,2-Dichloropropionate|2,2-Dichloropropionate
C1508164|T201|COMP|38288-7|LNC|1,2-Dibromo-3-Chloropropane|1,2-Dibromo-3-Chloropropane
C1508165|T201|COMP|38289-5|LNC|1,2-Dichlorobenzene|1,2-Dichlorobenzene
C1508166|T201|COMP|38290-3|LNC|1,4-Dichlorobenzene|1,4-Dichlorobenzene
C1508167|T201|COMP|38291-1|LNC|1,2-Dichloroethane|1,2-Dichloroethane
C1508168|T201|COMP|38292-9|LNC|1,1-Dichloroethylene|1,1-Dichloroethylene
C1508169|T201|COMP|38293-7|LNC|cis-1,2-Dichloroethylene|cis-1,2-Dichloroethylene
C1508170|T201|COMP|38294-5|LNC|Trans-1,2-Dichloroethylene|Trans-1,2-Dichloroethylene
C1508171|T201|COMP|38295-2|LNC|Methylene chloride|Methylene chloride
C1508172|T201|COMP|38296-0|LNC|1,2-Dichloropropane|1,2-Dichloropropane
C1508173|T201|COMP|38297-8|LNC|Di(2-Ethylhexyl) phthalate|Di(2-Ethylhexyl) phthalate
C1508174|T201|COMP|38298-6|LNC|Dinoseb|Dinoseb
C1508175|T201|COMP|38299-4|LNC|Dioxin|Dioxin
C1508176|T201|COMP|38300-0|LNC|Diquat|Diquat
C1508177|T201|COMP|38301-8|LNC|Endothall|Endothall
C1508178|T201|COMP|38302-6|LNC|Endrin|Endrin
C1508179|T201|COMP|38303-4|LNC|Epichlorohydrin|Epichlorohydrin
C1508180|T201|COMP|38304-2|LNC|Ethylene dibromide|Ethylene dibromide
C1508181|T201|COMP|38305-9|LNC|Glyphosate|Glyphosate
C1508182|T201|COMP|38306-7|LNC|Heptachlor|Heptachlor
C1508183|T201|COMP|38307-5|LNC|Heptachlorepoxide|Heptachlorepoxide
C1508184|T201|COMP|38308-3|LNC|Antimony|Antimony
C1508185|T201|COMP|38309-1|LNC|Asbestos|Asbestos
C1508186|T201|COMP|38310-9|LNC|Beryllium|Beryllium
C1508187|T201|COMP|38311-7|LNC|Thallium|Thallium
C1508188|T201|COMP|38312-5|LNC|Tetrachloroethylene|Tetrachloroethylene
C1508189|T201|COMP|38313-3|LNC|Toluene|Toluene
C1508190|T201|COMP|38314-1|LNC|Cyclohexanone|Cyclohexanone
C1508191|T201|COMP|38315-8|LNC|Dichlorobenzene|Dichlorobenzene
C1508192|T201|COMP|38316-6|LNC|Dichloroethane|Dichloroethane
C1508193|T201|COMP|38317-4|LNC|Hexane|Hexane
C1508194|T201|COMP|38318-2|LNC|Acrylamide|Acrylamide
C1508195|T201|COMP|38319-0|LNC|Alachlor|Alachlor
C1508196|T201|COMP|38320-8|LNC|Benzo alpha pyrene|Benzo alpha pyrene
C1508197|T201|COMP|38321-6|LNC|Carbofuran|Carbofuran
C1508198|T201|COMP|38322-4|LNC|Carbon tetrachloride|Carbon tetrachloride
C1508199|T201|COMP|38323-2|LNC|Lindane|Lindane
C1508200|T201|COMP|38324-0|LNC|Methoxychlor|Methoxychlor
C1508201|T201|COMP|38325-7|LNC|Oxamyl|Oxamyl
C1508202|T201|COMP|38326-5|LNC|Pentachlorophenol|Pentachlorophenol
C1508203|T201|COMP|38327-3|LNC|Picloram|Picloram
C1508204|T201|COMP|38328-1|LNC|Simazine|Simazine
C1508205|T201|COMP|38329-9|LNC|Styrene|Styrene
C1508206|T201|COMP|38330-7|LNC|Toxaphene|Toxaphene
C1508207|T201|COMP|38331-5|LNC|2,4,5-Trichlorophenoxyacetate|2,4,5-Trichlorophenoxyacetate
C1508208|T201|COMP|38332-3|LNC|1,2,4-Trichlorobenzene|1,2,4-Trichlorobenzene
C1508209|T201|COMP|38333-1|LNC|Trichloroethane|Trichloroethane
C1508210|T201|COMP|38334-9|LNC|1,1,2-Trichloroethane|1,1,2-Trichloroethane
C1508211|T201|COMP|38335-6|LNC|Vinyl chloride|Vinyl chloride
C1508212|T201|COMP|38336-4|LNC|Ethyl benzene|Ethyl benzene
C1508213|T201|COMP|38337-2|LNC|Hexachlorocyclopentadiene|Hexachlorocyclopentadiene
C1508214|T201|COMP|38338-0|LNC|Cyanide|Cyanide
C1508215|T201|COMP|38339-8|LNC|Benzene|Benzene
C1508216|T201|COMP|38340-6|LNC|Dichlorodiphenyltrichloroethane|Dichlorodiphenyltrichloroethane
C1508217|T201|COMP|38341-4|LNC|Chlordane|Chlordane
C1508218|T201|COMP|38342-2|LNC|Hexachlorobenzene|Hexachlorobenzene
C1508219|T201|COMP|38343-0|LNC|Chlorobenzene|Chlorobenzene
C1508220|T201|COMP|38344-8|LNC|Trichloroethylene|Trichloroethylene
C1508221|T201|COMP|38345-5|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C1508222|T201|COMP|38346-3|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C1508764|T201|COMP|13446-0|LNC|Creatinine renal clearance/1.73 sq M|Creatinine renal clearance/1.73 sq M
C1508765|T201|COMP|13447-8|LNC|Creatinine renal clearance/1.73 sq M|Creatinine renal clearance/1.73 sq M
C1508766|T201|COMP|13449-4|LNC|Creatinine renal clearance/1.73 sq M|Creatinine renal clearance/1.73 sq M
C1510482|T201|COMP|14822-1|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C1524719|T201|COMP|38391-9|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C1524720|T201|COMP|38392-7|LNC|Legionella sp Ab|Legionella sp Ab
C1524721|T201|COMP|38393-5|LNC|Legionella sp identified|Legionella sp identified
C1524722|T201|COMP|38394-3|LNC|Legionella sp identified|Legionella sp identified
C1524723|T201|COMP|38395-0|LNC|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C1524724|T201|COMP|38396-8|LNC|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C1524725|T201|COMP|38397-6|LNC|Crystals|Crystals
C1524726|T201|COMP|38398-4|LNC|Crystals|Crystals
C1524727|T201|COMP|38399-2|LNC|Crystals|Crystals
C1524728|T201|COMP|38400-8|LNC|Parainfluenza virus 1+2+3 Ab|Parainfluenza virus 1+2+3 Ab
C1525151|T201|COMP|38654-0|LNC|Chloroacetate|Chloroacetate
C1525152|T201|COMP|38655-7|LNC|2-Chloroacetophenone|2-Chloroacetophenone
C1525153|T201|COMP|38656-5|LNC|Chlorobenzilate|Chlorobenzilate
C1525154|T201|COMP|38657-3|LNC|Diazomethane|Diazomethane
C1525155|T201|COMP|38658-1|LNC|Acetate|Acetate
C1525156|T201|COMP|38659-9|LNC|Acetophenone|Acetophenone
C1525157|T201|COMP|38660-7|LNC|Acetylene|Acetylene
C1525158|T201|COMP|38661-5|LNC|Aldrin|Aldrin
C1525159|T201|COMP|38662-3|LNC|Aluminum oxide|Aluminum oxide
C1525160|T201|COMP|38764-7|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C1525921|T201|COMP|38757-1|LNC|1,3-Dimethylbenzene|1,3-Dimethylbenzene
C1525922|T201|COMP|38758-9|LNC|1,4-Dimethylbenzene|1,4-Dimethylbenzene
C1525923|T201|COMP|38759-7|LNC|Aluminum|Aluminum
C1525924|T201|COMP|38760-5|LNC|Dibenzofuran|Dibenzofuran
C1525925|T201|COMP|38761-3|LNC|Asphalt|Asphalt
C1525926|T201|COMP|38762-1|LNC|Isooctane|Isooctane
C1525927|T201|COMP|38763-9|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C1526359|T201|COMP|38347-1|LNC|XXX microorganism DNA|XXX microorganism DNA
C1526360|T201|COMP|38348-9|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1526361|T201|COMP|38349-7|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1526362|T201|COMP|38350-5|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1526363|T201|COMP|38351-3|LNC|Herpes virus 6 DNA panel|Herpes virus 6 DNA panel
C1526364|T201|COMP|38352-1|LNC|Interleukin 2 receptor|Interleukin 2 receptor
C1526365|T201|COMP|38353-9|LNC|Streptococcus sp identified|Streptococcus sp identified
C1526366|T201|COMP|38354-7|LNC|Bartonella sp identified|Bartonella sp identified
C1526367|T201|COMP|38355-4|LNC|Chitotriosidase|Chitotriosidase
C1526368|T201|COMP|38356-2|LNC|Thyroxine Ab|Thyroxine Ab
C1526369|T201|COMP|38357-0|LNC|B cell crossmatch|B cell crossmatch
C1526370|T201|COMP|38358-8|LNC|A Ab|A Ab
C1526371|T201|COMP|38359-6|LNC|A Ab|A Ab
C1526372|T201|COMP|38360-4|LNC|Isobutyrylglycine/Creatinine|Isobutyrylglycine/Creatinine
C1526374|T201|COMP|38362-0|LNC|Muscle specific receptor tyrosine kinase Ab|Muscle specific receptor tyrosine kinase Ab
C1526375|T201|COMP|38363-8|LNC|Cefepime|Cefepime
C1526376|T201|COMP|38364-6|LNC|Haloperidol.reduced|Haloperidol.reduced
C1526377|T201|COMP|38365-3|LNC|Hexadecadienoate/Creatinine|Hexadecadienoate/Creatinine
C1526378|T201|COMP|38366-1|LNC|Hypoxanthine/Creatinine|Hypoxanthine/Creatinine
C1526379|T201|COMP|38367-9|LNC|N-octanoylglycine/Creatinine|N-octanoylglycine/Creatinine
C1526380|T201|COMP|38368-7|LNC|Pigeon droppings Ab.IgG|Pigeon droppings Ab.IgG
C1526381|T201|COMP|38369-5|LNC|U1 small nuclear ribonucleoprotein Ab.IgG|U1 small nuclear ribonucleoprotein Ab.IgG
C1526382|T201|COMP|38370-3|LNC|Voriconazole|Voriconazole
C1526383|T201|COMP|38371-1|LNC|Xanthine/Creatinine|Xanthine/Creatinine
C1526385|T201|COMP|38373-7|LNC|Buprenorphine+Norbuprenorphine|Buprenorphine+Norbuprenorphine
C1526386|T201|COMP|38374-5|LNC|Tenofovir|Tenofovir
C1526387|T201|COMP|38375-2|LNC|Adenovirus DNA|Adenovirus DNA
C1526388|T201|COMP|38376-0|LNC|Cryptococcus sp identified|Cryptococcus sp identified
C1526389|T201|COMP|38377-8|LNC|Cryptococcus neoformans|Cryptococcus neoformans
C1526390|T201|COMP|38378-6|LNC|Mycobacterium tuberculosis complex rRNA|Mycobacterium tuberculosis complex rRNA
C1526391|T201|COMP|38379-4|LNC|Mycobacterium tuberculosis complex DNA|Mycobacterium tuberculosis complex DNA
C1526392|T201|COMP|38380-2|LNC|HFE gene.p.Ser65Cys|HFE gene.p.Ser65Cys
C1526393|T201|COMP|38381-0|LNC|Influenza virus A cDNA|Influenza virus A cDNA
C1526394|T201|COMP|38382-8|LNC|Influenza virus B|Influenza virus B
C1526395|T201|COMP|38383-6|LNC|Enterococcus sp rRNA|Enterococcus sp rRNA
C1526396|T201|COMP|38384-4|LNC|Cocaine|Cocaine
C1526397|T201|COMP|38385-1|LNC|Coccidioides immitis Ag|Coccidioides immitis Ag
C1526398|T201|COMP|38386-9|LNC|Color|Color
C1526399|T201|COMP|38387-7|LNC|C3 nephritic factor|C3 nephritic factor
C1526400|T201|COMP|38388-5|LNC|Complement C3|Complement C3
C1526401|T201|COMP|38389-3|LNC|Coxiella burnetii phase 2 Ab|Coxiella burnetii phase 2 Ab
C1526402|T201|COMP|38390-1|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C1526403|T201|COMP|38401-6|LNC|Protozoa identified|Protozoa identified
C1526404|T201|COMP|38402-4|LNC|Parasite identified|Parasite identified
C1526405|T201|COMP|38403-2|LNC|Cyclospora sp Ag|Cyclospora sp Ag
C1526406|T201|COMP|38404-0|LNC|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C1526407|T201|COMP|38405-7|LNC|MT-ATP6 gene targeted mutation analysis|MT-ATP6 gene targeted mutation analysis
C1526408|T201|COMP|38407-3|LNC|PAX3 gene targeted mutation analysis|PAX3 gene targeted mutation analysis
C1526409|T201|COMP|38408-1|LNC|PEO gene targeted mutation analysis|PEO gene targeted mutation analysis
C1526410|T201|COMP|38409-9|LNC|SERPINA1 gene targeted mutation analysis|SERPINA1 gene targeted mutation analysis
C1526411|T201|COMP|38410-7|LNC|Basement membrane zone Ab|Basement membrane zone Ab
C1526412|T201|COMP|38411-5|LNC|TOR1A gene targeted mutation analysis|TOR1A gene targeted mutation analysis
C1526413|T201|COMP|38412-3|LNC|FGFR2 gene targeted mutation analysis|FGFR2 gene targeted mutation analysis
C1526414|T201|COMP|38413-1|LNC|FGFR3 gene targeted mutation analysis|FGFR3 gene targeted mutation analysis
C1526415|T201|COMP|38414-9|LNC|Iron|Iron
C1526416|T201|COMP|38415-6|LNC|MTHFR gene targeted mutation analysis|MTHFR gene targeted mutation analysis
C1526417|T201|COMP|38416-4|LNC|Parasite identified|Parasite identified
C1526418|T201|COMP|38417-2|LNC|Trans-cinnamoylglycine/Creatinine|Trans-cinnamoylglycine/Creatinine
C1526419|T201|COMP|38418-0|LNC|Pigeon droppings Ab.IgG|Pigeon droppings Ab.IgG
C1526420|T201|COMP|38419-8|LNC|Cells.CD21/100 cells|Cells.CD21/100 cells
C1526421|T201|COMP|38420-6|LNC|Soluble liver Ab.IgG|Soluble liver Ab.IgG
C1526422|T201|COMP|38421-4|LNC|C peptide^30M post XXX challenge|C peptide^30M post XXX challenge
C1526423|T201|COMP|38422-2|LNC|C peptide^1H post XXX challenge|C peptide^1H post XXX challenge
C1526424|T201|COMP|38423-0|LNC|C peptide^1.5H post XXX challenge|C peptide^1.5H post XXX challenge
C1526425|T201|COMP|38424-8|LNC|C peptide^2H post XXX challenge|C peptide^2H post XXX challenge
C1526426|T201|COMP|38425-5|LNC|C peptide^2.5H post XXX challenge|C peptide^2.5H post XXX challenge
C1526427|T201|COMP|38426-3|LNC|C peptide^3H post XXX challenge|C peptide^3H post XXX challenge
C1526428|T201|COMP|38427-1|LNC|Thiocyanate|Thiocyanate
C1526429|T201|COMP|38428-9|LNC|Ibuprofen^pre dose|Ibuprofen^pre dose
C1526430|T201|COMP|38429-7|LNC|Ibuprofen^30M post dose|Ibuprofen^30M post dose
C1526431|T201|COMP|38430-5|LNC|Ibuprofen^1H post dose|Ibuprofen^1H post dose
C1526432|T201|COMP|38431-3|LNC|Ibuprofen^1.5H post dose|Ibuprofen^1.5H post dose
C1526433|T201|COMP|38432-1|LNC|Ibuprofen^2H post dose|Ibuprofen^2H post dose
C1526434|T201|COMP|38433-9|LNC|Ibuprofen^2.5H post dose|Ibuprofen^2.5H post dose
C1526435|T201|COMP|38434-7|LNC|Ibuprofen^3H post dose|Ibuprofen^3H post dose
C1526437|T201|COMP|38436-2|LNC|Colony count|Colony count
C1526438|T201|COMP|38437-0|LNC|Anacardium occidentale Ab.IgE/IgE.total|Anacardium occidentale Ab.IgE/IgE.total
C1526439|T201|COMP|38438-8|LNC|Aspergillus fumigatus Ab.IgE/IgE.total|Aspergillus fumigatus Ab.IgE/IgE.total
C1526440|T201|COMP|38439-6|LNC|Barbiturates|Barbiturates
C1526441|T201|COMP|38440-4|LNC|Basement membrane zone Ab|Basement membrane zone Ab
C1526442|T201|COMP|38441-2|LNC|Benzodiazepines|Benzodiazepines
C1526443|T201|COMP|38442-0|LNC|Bilirubin crystals|Bilirubin crystals
C1526444|T201|COMP|38443-8|LNC|Blastomyces dermatitidis Ab.IgM|Blastomyces dermatitidis Ab.IgM
C1526445|T201|COMP|38444-6|LNC|Bromide|Bromide
C1526446|T201|COMP|38445-3|LNC|Calprotectin|Calprotectin
C1526447|T201|COMP|38446-1|LNC|Catecholamines|Catecholamines
C1526448|T201|COMP|38447-9|LNC|CFTR gene.c.711+1G>T|CFTR gene.c.711+1G>T
C1526449|T201|COMP|38448-7|LNC|CFTR gene.p.Ala455Glu|CFTR gene.p.Ala455Glu
C1526450|T201|COMP|38449-5|LNC|CFTR gene.c.1078delT|CFTR gene.c.1078delT
C1526451|T201|COMP|38450-3|LNC|CFTR gene.c.2184delA|CFTR gene.c.2184delA
C1526452|T201|COMP|38451-1|LNC|CFTR gene.c.2789+5G>A|CFTR gene.c.2789+5G>A
C1526453|T201|COMP|38452-9|LNC|CFTR gene.c.3120+1G>A|CFTR gene.c.3120+1G>A
C1526454|T201|COMP|38453-7|LNC|CFTR gene.c.3659delC|CFTR gene.c.3659delC
C1526455|T201|COMP|38454-5|LNC|CFTR gene.p.Gly85Glu|CFTR gene.p.Gly85Glu
C1526456|T201|COMP|38455-2|LNC|CFTR gene.c.621+1G>T|CFTR gene.c.621+1G>T
C1526457|T201|COMP|38456-0|LNC|CFTR gene.c.3849+10kbC>T|CFTR gene.c.3849+10kbC>T
C1526458|T201|COMP|38457-8|LNC|Immune complex.C3d+IgG|Immune complex.C3d+IgG
C1526459|T201|COMP|38458-6|LNC|Crystals|Crystals
C1526460|T201|COMP|38459-4|LNC|Crystals|Crystals
C1526461|T201|COMP|38460-2|LNC|Legionella sp Ag|Legionella sp Ag
C1526462|T201|COMP|38461-0|LNC|Legionella sp Ag|Legionella sp Ag
C1526463|T201|COMP|38462-8|LNC|Legionella sp Ag|Legionella sp Ag
C1526464|T201|COMP|38463-6|LNC|Legionella sp Ag|Legionella sp Ag
C1526465|T201|COMP|38464-4|LNC|Juniperus sabinoides Ab.IgE/IgE.total|Juniperus sabinoides Ab.IgE/IgE.total
C1526466|T201|COMP|38465-1|LNC|Chicken Ab.IgE/IgE.total|Chicken Ab.IgE/IgE.total
C1526467|T201|COMP|38466-9|LNC|Chicken serum proteins Ab.IgG|Chicken serum proteins Ab.IgG
C1526468|T201|COMP|38467-7|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C1526469|T201|COMP|38468-5|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C1526470|T201|COMP|38469-3|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1526471|T201|COMP|38470-1|LNC|chlorproPAMIDE|chlorproPAMIDE
C1526472|T201|COMP|38471-9|LNC|Karyotype|Karyotype
C1526473|T201|COMP|38472-7|LNC|17-Hydroxycorticosteroids/Creatinine|17-Hydroxycorticosteroids/Creatinine
C1526474|T201|COMP|38473-5|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C1526475|T201|COMP|38474-3|LNC|Acylcarnitine|Acylcarnitine
C1526476|T201|COMP|38475-0|LNC|Acid alpha glucosidase|Acid alpha glucosidase
C1526477|T201|COMP|38476-8|LNC|Mullerian inhibiting substance|Mullerian inhibiting substance
C1526478|T201|COMP|38477-6|LNC|Glucosylceramidase|Glucosylceramidase
C1526479|T201|COMP|38478-4|LNC|Biotinidase|Biotinidase
C1526480|T201|COMP|38479-2|LNC|Branched chain keto-acid dehydrogenase complex|Branched chain keto-acid dehydrogenase complex
C1526481|T201|COMP|38480-0|LNC|Carnitine|Carnitine
C1526482|T201|COMP|38481-8|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C1526483|T201|COMP|38482-6|LNC|Creatine kinase.MB|Creatine kinase.MB
C1526484|T201|COMP|38483-4|LNC|Creatinine|Creatinine
C1526485|T201|COMP|38484-2|LNC|Cysteine|Cysteine
C1526486|T201|COMP|38485-9|LNC|Galactose 1 phosphate|Galactose 1 phosphate
C1526487|T201|COMP|38486-7|LNC|Homocystine|Homocystine
C1526488|T201|COMP|38487-5|LNC|IgA|IgA
C1526489|T201|COMP|38488-3|LNC|IgG|IgG
C1526490|T201|COMP|38489-1|LNC|Insulin bovine Ab|Insulin bovine Ab
C1526491|T201|COMP|38490-9|LNC|Insulin porcine Ab|Insulin porcine Ab
C1526493|T201|COMP|38492-5|LNC|Insulin-like growth factor-I|Insulin-like growth factor-I
C1526494|T201|COMP|38493-3|LNC|Ketones|Ketones
C1526495|T201|COMP|38494-1|LNC|Metanephrine.free|Metanephrine.free
C1526496|T201|COMP|38495-8|LNC|Phenylalanine+Tyrosine|Phenylalanine+Tyrosine
C1526497|T201|COMP|38496-6|LNC|Retinyl palmitate|Retinyl palmitate
C1526498|T201|COMP|38497-4|LNC|Spermatozoa.amorphous head|Spermatozoa.amorphous head
C1526499|T201|COMP|38498-2|LNC|Spermatozoa.nonviable/100 spermatozoa|Spermatozoa.nonviable/100 spermatozoa
C1526500|T201|COMP|38499-0|LNC|Spermatozoa.progressive^4H post ejaculation|Spermatozoa.progressive^4H post ejaculation
C1526501|T201|COMP|38500-5|LNC|Spermatozoa.progressive.grade 1/100 spermatozoa|Spermatozoa.progressive.grade 1/100 spermatozoa
C1526502|T201|COMP|38501-3|LNC|Spermatozoa.progressive.grade 2/100 spermatozoa|Spermatozoa.progressive.grade 2/100 spermatozoa
C1526503|T201|COMP|38502-1|LNC|Spermatozoa.progressive.grade 4/100 spermatozoa|Spermatozoa.progressive.grade 4/100 spermatozoa
C1526504|T201|COMP|38503-9|LNC|Spermatozoa.progressive.grade 3/100 spermatozoa|Spermatozoa.progressive.grade 3/100 spermatozoa
C1526505|T201|COMP|38504-7|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C1526506|T201|COMP|38505-4|LNC|Thyroglobulin recovery|Thyroglobulin recovery
C1526507|T201|COMP|38506-2|LNC|Thyroxine|Thyroxine
C1526508|T201|COMP|38507-0|LNC|Urobilinogen|Urobilinogen
C1526509|T201|COMP|38508-8|LNC|Uroporphyrin/Creatinine|Uroporphyrin/Creatinine
C1526510|T201|COMP|38509-6|LNC|Viscosity^30M post collection|Viscosity^30M post collection
C1526511|T201|COMP|38510-4|LNC|Cells.CD11b+CD11c+/100 cells|Cells.CD11b+CD11c+/100 cells
C1526512|T201|COMP|38511-2|LNC|Cells.CD19+CD33+/100 cells|Cells.CD19+CD33+/100 cells
C1526513|T201|COMP|38512-0|LNC|Cells.CD2+CD3+/100 cells|Cells.CD2+CD3+/100 cells
C1526514|T201|COMP|38513-8|LNC|Cells.CD2+CD3+|Cells.CD2+CD3+
C1526515|T201|COMP|38514-6|LNC|Cells.CD33+CD34+/100 cells|Cells.CD33+CD34+/100 cells
C1526516|T201|COMP|38515-3|LNC|Cells.cytoplasmic Ig mu|Cells.cytoplasmic Ig mu
C1526519|T201|COMP|38518-7|LNC|Granulocytes.immature/100 leukocytes|Granulocytes.immature/100 leukocytes
C1526521|T201|COMP|38520-3|LNC|Capillary fragility|Capillary fragility
C1526522|T201|COMP|38521-1|LNC|Coagulation factor VIII Ag actual/Normal|Coagulation factor VIII Ag actual/Normal
C1526523|T201|COMP|38522-9|LNC|Complement C4b binding protein actual/Normal|Complement C4b binding protein actual/Normal
C1526524|T201|COMP|38523-7|LNC|Fibrinopeptide A|Fibrinopeptide A
C1526525|T201|COMP|38524-5|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C1526526|T201|COMP|38525-2|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C1526527|T201|COMP|38526-0|LNC|Number of specimens tested|Number of specimens tested
C1526528|T201|COMP|38527-8|LNC|Number of specimens received|Number of specimens received
C1526529|T201|COMP|38528-6|LNC|Protein.abnormal band|Protein.abnormal band
C1526530|T201|COMP|38529-4|LNC|CMTX2 gene targeted mutation analysis|CMTX2 gene targeted mutation analysis
C1526531|T201|COMP|38530-2|LNC|BRCA2 gene targeted mutation analysis|BRCA2 gene targeted mutation analysis
C1526532|T201|COMP|38531-0|LNC|BRCA2 gene mutations tested for|BRCA2 gene mutations tested for
C1526533|T201|COMP|38532-8|LNC|SPG3A gene targeted mutation analysis|SPG3A gene targeted mutation analysis
C1526534|T201|COMP|38533-6|LNC|TCOF1 gene targeted mutation analysis|TCOF1 gene targeted mutation analysis
C1526535|T201|COMP|38534-4|LNC|COL5A1 gene targeted mutation analysis|COL5A1 gene targeted mutation analysis
C1526536|T201|COMP|38535-1|LNC|LAMA2 gene targeted mutation analysis|LAMA2 gene targeted mutation analysis
C1526537|T201|COMP|38536-9|LNC|MLH1 gene targeted mutation analysis|MLH1 gene targeted mutation analysis
C1526538|T201|COMP|38537-7|LNC|ARX gene targeted mutation analysis|ARX gene targeted mutation analysis
C1526539|T201|COMP|38538-5|LNC|Fatty acids.very long chain.C26:1/C22:0|Fatty acids.very long chain.C26:1/C22:0
C1526540|T201|COMP|38539-3|LNC|Spermatozoa.motile/100 spermatozoa^post washing|Spermatozoa.motile/100 spermatozoa^post washing
C1526541|T201|COMP|38540-1|LNC|Spermatozoa.motile/100 spermatozoa^pre washing|Spermatozoa.motile/100 spermatozoa^pre washing
C1526542|T201|COMP|38541-9|LNC|Spermatozoa.motile^pre washing|Spermatozoa.motile^pre washing
C1526543|T201|COMP|38542-7|LNC|Repaglinide|Repaglinide
C1526544|T201|COMP|38543-5|LNC|Spermatozoa^post washing|Spermatozoa^post washing
C1526545|T201|COMP|38544-3|LNC|Spermatozoa^pre washing|Spermatozoa^pre washing
C1526546|T201|COMP|38545-0|LNC|Methylmercury|Methylmercury
C1526547|T201|COMP|38546-8|LNC|HLA-B locus|HLA-B locus
C1526548|T201|COMP|38547-6|LNC|HLA-C locus|HLA-C locus
C1526549|T201|COMP|38548-4|LNC|HLA-A locus|HLA-A locus
C1526550|T201|COMP|38549-2|LNC|HLA-B W locus|HLA-B W locus
C1526551|T201|COMP|38550-0|LNC|MSH2 gene targeted mutation analysis|MSH2 gene targeted mutation analysis
C1526552|T201|COMP|38551-8|LNC|Cortisol^pre or post dose dexamethasone|Cortisol^pre or post dose dexamethasone
C1526553|T201|COMP|38552-6|LNC|Acylcarnitine.short chain|Acylcarnitine.short chain
C1526554|T201|COMP|38553-4|LNC|Narcolepsy associated Ag|Narcolepsy associated Ag
C1526555|T201|COMP|38554-2|LNC|Spermatozoa.head.motile with IgA/100 spermatozoa|Spermatozoa.head.motile with IgA/100 spermatozoa
C1526556|T201|COMP|38555-9|LNC|Spermatozoa.head.motile with IgG/100 spermatozoa|Spermatozoa.head.motile with IgG/100 spermatozoa
C1526557|T201|COMP|38556-7|LNC|Spermatozoa.head.motile with IgM/100 spermatozoa|Spermatozoa.head.motile with IgM/100 spermatozoa
C1526561|T201|COMP|38560-9|LNC|Spermatozoa.tail.motile with IgA/100 spermatozoa|Spermatozoa.tail.motile with IgA/100 spermatozoa
C1526562|T201|COMP|38561-7|LNC|Spermatozoa.tail.motile with IgG/100 spermatozoa|Spermatozoa.tail.motile with IgG/100 spermatozoa
C1526563|T201|COMP|38562-5|LNC|Spermatozoa.tail.motile with IgM/100 spermatozoa|Spermatozoa.tail.motile with IgM/100 spermatozoa
C1526567|T201|COMP|38566-6|LNC|Spermatozoa.motile^post washing|Spermatozoa.motile^post washing
C1526568|T201|COMP|38567-4|LNC|Aniline|Aniline
C1526569|T201|COMP|38568-2|LNC|Asbestos|Asbestos
C1526570|T201|COMP|38569-0|LNC|Arsenic|Arsenic
C1526571|T201|COMP|38570-8|LNC|Azinphos-methyl|Azinphos-methyl
C1526572|T201|COMP|38571-6|LNC|Barium|Barium
C1526573|T201|COMP|38572-4|LNC|Benzidine|Benzidine
C1526574|T201|COMP|38573-2|LNC|Acrylamide|Acrylamide
C1526575|T201|COMP|38574-0|LNC|Beryllium|Beryllium
C1526576|T201|COMP|38575-7|LNC|Bromoform|Bromoform
C1526577|T201|COMP|38576-5|LNC|Butane|Butane
C1526578|T201|COMP|38577-3|LNC|Carbon disulfide|Carbon disulfide
C1526579|T201|COMP|38578-1|LNC|Carbon tetrachloride|Carbon tetrachloride
C1526580|T201|COMP|38579-9|LNC|Chlordane|Chlordane
C1526581|T201|COMP|38580-7|LNC|Cresols|Cresols
C1526582|T201|COMP|38581-5|LNC|Cumene|Cumene
C1526583|T201|COMP|38582-3|LNC|2,4-Dichlorophenoxyacetate|2,4-Dichlorophenoxyacetate
C1526584|T201|COMP|38583-1|LNC|1,2-Dibromo-3-Chloropropane|1,2-Dibromo-3-Chloropropane
C1526585|T201|COMP|38584-9|LNC|Acetaldehyde|Acetaldehyde
C1526586|T201|COMP|38585-6|LNC|Acetone|Acetone
C1526587|T201|COMP|38586-4|LNC|Acetonitrile|Acetonitrile
C1526588|T201|COMP|38587-2|LNC|Acrylaldehyde|Acrylaldehyde
C1526589|T201|COMP|38588-0|LNC|Acrylonitrile|Acrylonitrile
C1526590|T201|COMP|38589-8|LNC|Ammonia|Ammonia
C1526591|T201|COMP|38590-6|LNC|1,4-Dichlorobenzene|1,4-Dichlorobenzene
C1526592|T201|COMP|38591-4|LNC|Dichlorvos|Dichlorvos
C1526593|T201|COMP|38592-2|LNC|Dimethylformamide|Dimethylformamide
C1526594|T201|COMP|38593-0|LNC|1,4-Dioxane|1,4-Dioxane
C1526595|T201|COMP|38594-8|LNC|Epichlorohydrin|Epichlorohydrin
C1526596|T201|COMP|38595-5|LNC|Ethylene dibromide|Ethylene dibromide
C1526597|T201|COMP|38596-3|LNC|Ethylene glycol|Ethylene glycol
C1526598|T201|COMP|38597-1|LNC|Heptachlor|Heptachlor
C1526599|T201|COMP|38598-9|LNC|Hexachlorobenzene|Hexachlorobenzene
C1526600|T201|COMP|38599-7|LNC|Hexachlorobutadiene|Hexachlorobutadiene
C1526601|T201|COMP|38600-3|LNC|Hexachloroethane|Hexachloroethane
C1526602|T201|COMP|38601-1|LNC|Hexane|Hexane
C1526603|T201|COMP|38602-9|LNC|Hydrazine|Hydrazine
C1526604|T201|COMP|38603-7|LNC|Hydrogen sulfide|Hydrogen sulfide
C1526605|T201|COMP|38604-5|LNC|Hydroquinone|Hydroquinone
C1526606|T201|COMP|38605-2|LNC|Lindane|Lindane
C1526607|T201|COMP|38606-0|LNC|Maleic anhydride|Maleic anhydride
C1526608|T201|COMP|38607-8|LNC|Methoxychlor|Methoxychlor
C1526609|T201|COMP|38608-6|LNC|Methyl bromide|Methyl bromide
C1526610|T201|COMP|38609-4|LNC|Methyl tert-butyl ether|Methyl tert-butyl ether
C1526611|T201|COMP|38610-2|LNC|Methylene chloride|Methylene chloride
C1526612|T201|COMP|38611-0|LNC|Methyl isobutyl ketone|Methyl isobutyl ketone
C1526613|T201|COMP|38612-8|LNC|Naphthalene|Naphthalene
C1526614|T201|COMP|38613-6|LNC|Parathion|Parathion
C1526615|T201|COMP|38614-4|LNC|Pentachlorophenol|Pentachlorophenol
C1526616|T201|COMP|38615-1|LNC|Phenol|Phenol
C1526617|T201|COMP|38616-9|LNC|Propoxur|Propoxur
C1526618|T201|COMP|38617-7|LNC|1,2-Dichloropropane|1,2-Dichloropropane
C1526619|T201|COMP|38618-5|LNC|Styrene|Styrene
C1526620|T201|COMP|38619-3|LNC|Dioxin|Dioxin
C1526621|T201|COMP|38620-1|LNC|Tetrachloroethylene|Tetrachloroethylene
C1526622|T201|COMP|38621-9|LNC|Toluene|Toluene
C1526623|T201|COMP|38622-7|LNC|Toxaphene|Toxaphene
C1526624|T201|COMP|38623-5|LNC|1,2,4-Trichlorobenzene|1,2,4-Trichlorobenzene
C1526625|T201|COMP|38624-3|LNC|1,1,2-Trichloroethane|1,1,2-Trichloroethane
C1526626|T201|COMP|38625-0|LNC|Trichloroethylene|Trichloroethylene
C1526627|T201|COMP|38626-8|LNC|Vinyl chloride|Vinyl chloride
C1526628|T201|COMP|38627-6|LNC|Benzene|Benzene
C1526629|T201|COMP|38628-4|LNC|Benzo alpha pyrene|Benzo alpha pyrene
C1526630|T201|COMP|38629-2|LNC|Acetamide|Acetamide
C1526631|T201|COMP|38630-0|LNC|Acrylate|Acrylate
C1526632|T201|COMP|38631-8|LNC|Allyl chloride|Allyl chloride
C1526633|T201|COMP|38632-6|LNC|4-Biphenylamine|4-Biphenylamine
C1526634|T201|COMP|38633-4|LNC|Benzotrichloride|Benzotrichloride
C1526635|T201|COMP|38634-2|LNC|Benzyl chloride|Benzyl chloride
C1526636|T201|COMP|38635-9|LNC|Biphenyl|Biphenyl
C1526637|T201|COMP|38636-7|LNC|Di(2-Ethylhexyl) phthalate|Di(2-Ethylhexyl) phthalate
C1526638|T201|COMP|38637-5|LNC|Bis(chloromethyl)ether|Bis(chloromethyl)ether
C1526639|T201|COMP|38638-3|LNC|Boron oxide|Boron oxide
C1526640|T201|COMP|38639-1|LNC|Boron trifluoride|Boron trifluoride
C1526641|T201|COMP|38640-9|LNC|Bromine|Bromine
C1526642|T201|COMP|38641-7|LNC|Ethyl bromide|Ethyl bromide
C1526643|T201|COMP|38642-5|LNC|1,3-Butadiene|1,3-Butadiene
C1526644|T201|COMP|38643-3|LNC|Calcium cyanamide|Calcium cyanamide
C1526645|T201|COMP|38644-1|LNC|Caprolactam|Caprolactam
C1526646|T201|COMP|38645-8|LNC|Captan|Captan
C1526647|T201|COMP|38646-6|LNC|Catechol|Catechol
C1526648|T201|COMP|38647-4|LNC|Chlorine|Chlorine
C1526649|T201|COMP|38648-2|LNC|Chlorobenzene|Chlorobenzene
C1526650|T201|COMP|38649-0|LNC|Chloroform|Chloroform
C1526651|T201|COMP|38650-8|LNC|Chloromethyl methyl ether|Chloromethyl methyl ether
C1526652|T201|COMP|38651-6|LNC|2-Chloro-1,3-Butadiene|2-Chloro-1,3-Butadiene
C1526653|T201|COMP|38652-4|LNC|Carbonyl sulfide|Carbonyl sulfide
C1526654|T201|COMP|38653-2|LNC|Amiben|Amiben
C1526655|T201|COMP|38663-1|LNC|Dichlorobenzidine|Dichlorobenzidine
C1526656|T201|COMP|38664-9|LNC|Bis(2-Chloroethyl) ether|Bis(2-Chloroethyl) ether
C1526657|T201|COMP|38665-6|LNC|Diethanolamine|Diethanolamine
C1526658|T201|COMP|38666-4|LNC|Diethylsulfate|Diethylsulfate
C1526659|T201|COMP|38667-2|LNC|3,3'-Dimethoxybenzidine|3,3'-Dimethoxybenzidine
C1526660|T201|COMP|38668-0|LNC|Dimethylaniline|Dimethylaniline
C1526661|T201|COMP|38669-8|LNC|Dichlorodiphenyldichloroethylene|Dichlorodiphenyldichloroethylene
C1526662|T201|COMP|38670-6|LNC|Orthocresol|Orthocresol
C1526663|T201|COMP|38671-4|LNC|M-cresol|M-cresol
C1526664|T201|COMP|38672-2|LNC|P-cresol|P-cresol
C1526665|T201|COMP|38673-0|LNC|Dimethylphthalate|Dimethylphthalate
C1526666|T201|COMP|38674-8|LNC|Spermatozoa.head Ab.IgA/100 spermatozoa|Spermatozoa.head Ab.IgA/100 spermatozoa
C1526667|T201|COMP|38675-5|LNC|Spermatozoa.midpiece Ab.IgA/100 spermatozoa|Spermatozoa.midpiece Ab.IgA/100 spermatozoa
C1526668|T201|COMP|38676-3|LNC|Spermatozoa.tail tip Ab.IgA/100 spermatozoa|Spermatozoa.tail tip Ab.IgA/100 spermatozoa
C1526669|T201|COMP|38677-1|LNC|Spermatozoa.tail Ab.IgA/100 spermatozoa|Spermatozoa.tail Ab.IgA/100 spermatozoa
C1526670|T201|COMP|38678-9|LNC|Spermatozoa.head Ab.IgG/100 spermatozoa|Spermatozoa.head Ab.IgG/100 spermatozoa
C1526671|T201|COMP|38679-7|LNC|Spermatozoa.midpiece Ab.IgG/100 spermatozoa|Spermatozoa.midpiece Ab.IgG/100 spermatozoa
C1526672|T201|COMP|38680-5|LNC|Spermatozoa.tail tip Ab.IgG/100 spermatozoa|Spermatozoa.tail tip Ab.IgG/100 spermatozoa
C1526673|T201|COMP|38681-3|LNC|Spermatozoa.tail Ab.IgG/100 spermatozoa|Spermatozoa.tail Ab.IgG/100 spermatozoa
C1526674|T201|COMP|38682-1|LNC|Spermatozoa.head Ab.IgM/100 spermatozoa|Spermatozoa.head Ab.IgM/100 spermatozoa
C1526675|T201|COMP|38683-9|LNC|Spermatozoa.midpiece Ab.IgM/100 spermatozoa|Spermatozoa.midpiece Ab.IgM/100 spermatozoa
C1526676|T201|COMP|38684-7|LNC|Spermatozoa.tail tip Ab.IgM/100 spermatozoa|Spermatozoa.tail tip Ab.IgM/100 spermatozoa
C1526677|T201|COMP|38685-4|LNC|Spermatozoa.tail Ab.IgM/100 spermatozoa|Spermatozoa.tail Ab.IgM/100 spermatozoa
C1526678|T201|COMP|38686-2|LNC|Spermatozoa Ab.IgA+IgG/100 spermatozoa|Spermatozoa Ab.IgA+IgG/100 spermatozoa
C1526679|T201|COMP|38687-0|LNC|2-Acetylaminofluorene|2-Acetylaminofluorene
C1526680|T201|COMP|38688-8|LNC|1,1-Dimethylhydrazine|1,1-Dimethylhydrazine
C1526681|T201|COMP|38689-6|LNC|Dimethyl sulfate|Dimethyl sulfate
C1526682|T201|COMP|38690-4|LNC|4,6-Dinitro-O-Cresol|4,6-Dinitro-O-Cresol
C1526683|T201|COMP|38691-2|LNC|1,2-Diphenylhydrazine|1,2-Diphenylhydrazine
C1526684|T201|COMP|38692-0|LNC|1-Butene oxide|1-Butene oxide
C1526685|T201|COMP|38693-8|LNC|Ethyl acrylate|Ethyl acrylate
C1526686|T201|COMP|38694-6|LNC|Chloroethane|Chloroethane
C1526687|T201|COMP|38695-3|LNC|1,2-Dichloroethane|1,2-Dichloroethane
C1526688|T201|COMP|38696-1|LNC|Ethylene oxide|Ethylene oxide
C1526689|T201|COMP|38697-9|LNC|Ethylene thiourea|Ethylene thiourea
C1526690|T201|COMP|38698-7|LNC|Ethyleneimine|Ethyleneimine
C1526691|T201|COMP|38699-5|LNC|1,1-Dichloroethane|1,1-Dichloroethane
C1526692|T201|COMP|38700-1|LNC|Formaldehyde|Formaldehyde
C1526693|T201|COMP|38701-9|LNC|Hexachlorocyclopentadiene|Hexachlorocyclopentadiene
C1526694|T201|COMP|38702-7|LNC|Hexamethylene diisocyanate|Hexamethylene diisocyanate
C1526695|T201|COMP|38703-5|LNC|Hexamethylphosphoramide|Hexamethylphosphoramide
C1526696|T201|COMP|38704-3|LNC|Isophorone|Isophorone
C1526697|T201|COMP|38705-0|LNC|Methanol|Methanol
C1526698|T201|COMP|38706-8|LNC|Chloromethane|Chloromethane
C1526699|T201|COMP|38707-6|LNC|Trichloroethane|Trichloroethane
C1526700|T201|COMP|38708-4|LNC|Methyl hydrazine|Methyl hydrazine
C1526701|T201|COMP|38709-2|LNC|Methyl iodide|Methyl iodide
C1526702|T201|COMP|38710-0|LNC|Nitrobenzene|Nitrobenzene
C1526703|T201|COMP|38711-8|LNC|2-Nitropropane|2-Nitropropane
C1526704|T201|COMP|38712-6|LNC|N-nitrosodimethylamine|N-nitrosodimethylamine
C1526705|T201|COMP|38713-4|LNC|N-nitrosomorpholine|N-nitrosomorpholine
C1526706|T201|COMP|38714-2|LNC|Pentachloronitrobenzene|Pentachloronitrobenzene
C1526707|T201|COMP|38715-9|LNC|Phosgene|Phosgene
C1526708|T201|COMP|38716-7|LNC|Phosphine|Phosphine
C1526709|T201|COMP|38717-5|LNC|Phosphate|Phosphate
C1526710|T201|COMP|38718-3|LNC|Phthalic anhydride|Phthalic anhydride
C1526711|T201|COMP|38719-1|LNC|1,3-Propane sultone|1,3-Propane sultone
C1526712|T201|COMP|38720-9|LNC|Beta-propiolactone|Beta-propiolactone
C1526713|T201|COMP|38721-7|LNC|Propionaldehyde|Propionaldehyde
C1526714|T201|COMP|38722-5|LNC|Propyleneimine|Propyleneimine
C1526715|T201|COMP|38723-3|LNC|1,4-Benzoquinone|1,4-Benzoquinone
C1526716|T201|COMP|38724-1|LNC|Quinoline|Quinoline
C1526717|T201|COMP|38725-8|LNC|Styrene-7,8-Oxide|Styrene-7,8-Oxide
C1526718|T201|COMP|38726-6|LNC|Titanium tetrachloride|Titanium tetrachloride
C1526719|T201|COMP|38727-4|LNC|2,4 toluenediamine|2,4 toluenediamine
C1526720|T201|COMP|38728-2|LNC|2-Aminotoluene|2-Aminotoluene
C1526721|T201|COMP|38729-0|LNC|2,4,5-Trichlorophenol|2,4,5-Trichlorophenol
C1526722|T201|COMP|38730-8|LNC|2,4,6-Trichlorophenol|2,4,6-Trichlorophenol
C1526723|T201|COMP|38731-6|LNC|Triethylamine|Triethylamine
C1526724|T201|COMP|38732-4|LNC|Trifluralin|Trifluralin
C1526725|T201|COMP|38733-2|LNC|Vinyl acetate|Vinyl acetate
C1526726|T201|COMP|38734-0|LNC|Vinyl bromide|Vinyl bromide
C1526727|T201|COMP|38735-7|LNC|1,1-Dichloroethylene|1,1-Dichloroethylene
C1526728|T201|COMP|38736-5|LNC|Animal hair+Epithelium|Animal hair+Epithelium
C1526729|T201|COMP|38737-3|LNC|O-anisidine|O-anisidine
C1526730|T201|COMP|38738-1|LNC|Carbaryl|Carbaryl
C1526731|T201|COMP|38739-9|LNC|1,3-Dichloropropene|1,3-Dichloropropene
C1526732|T201|COMP|38740-7|LNC|Dimethylcarbamoyl chloride|Dimethylcarbamoyl chloride
C1526733|T201|COMP|38741-5|LNC|2,4-Dinitrophenol|2,4-Dinitrophenol
C1526734|T201|COMP|38742-3|LNC|2,4-Dinitrotoluene|2,4-Dinitrotoluene
C1526735|T201|COMP|38743-1|LNC|Hydrogen chloride|Hydrogen chloride
C1526736|T201|COMP|38744-9|LNC|Hydrogen fluoride|Hydrogen fluoride
C1526737|T201|COMP|38745-6|LNC|Diphenylmethane diisocyanate (MDI)|Diphenylmethane diisocyanate (MDI)
C1526738|T201|COMP|38746-4|LNC|4,4'-Methylene bis(2-Chloroaniline)|4,4'-Methylene bis(2-Chloroaniline)
C1526739|T201|COMP|38747-2|LNC|Methyl isocyanate|Methyl isocyanate
C1526740|T201|COMP|38748-0|LNC|Methylenedianiline|Methylenedianiline
C1526741|T201|COMP|38749-8|LNC|P-nitrobiphenyl|P-nitrobiphenyl
C1526742|T201|COMP|38750-6|LNC|Para nitrophenol|Para nitrophenol
C1526743|T201|COMP|38751-4|LNC|1,4-Benzenediamine|1,4-Benzenediamine
C1526744|T201|COMP|38752-2|LNC|Polychlorinated biphenyl|Polychlorinated biphenyl
C1526745|T201|COMP|38753-0|LNC|Tetrachloroethane|Tetrachloroethane
C1526746|T201|COMP|38754-8|LNC|2,4-Toluene diisocyanate|2,4-Toluene diisocyanate
C1526747|T201|COMP|38755-5|LNC|Dimethylbenzene|Dimethylbenzene
C1526748|T201|COMP|38756-3|LNC|1,2-Dimethylbenzene|1,2-Dimethylbenzene
C1527419|T201|COMP|11553-5|LNC|Microscopic exam|Microscopic exam
C1542883|T201|COMP|39595-4|LNC|Hippoglossus hippoglossus Ab.IgE/IgE.total|Hippoglossus hippoglossus Ab.IgE/IgE.total
C1542884|T201|COMP|39596-2|LNC|Mytilus edulis Ab.IgE/IgE.total|Mytilus edulis Ab.IgE/IgE.total
C1542885|T201|COMP|39597-0|LNC|Cucurbita pepo Ab.IgE/IgE.total|Cucurbita pepo Ab.IgE/IgE.total
C1542886|T201|COMP|39598-8|LNC|Curvularia lunata Ab.IgE/IgE.total|Curvularia lunata Ab.IgE/IgE.total
C1542887|T201|COMP|39599-6|LNC|Epicoccum purpurascens Ab.IgE/IgE.total|Epicoccum purpurascens Ab.IgE/IgE.total
C1542888|T201|COMP|39600-2|LNC|Fusarium moniliforme Ab.IgE/IgE.total|Fusarium moniliforme Ab.IgE/IgE.total
C1542889|T201|COMP|39601-0|LNC|Stemphylium botryosum Ab.IgE/IgE.total|Stemphylium botryosum Ab.IgE/IgE.total
C1542890|T201|COMP|39602-8|LNC|Hamster epithelium Ab.IgE/IgE.total|Hamster epithelium Ab.IgE/IgE.total
C1542891|T201|COMP|39603-6|LNC|Guinea pig epithelium Ab.IgE/IgE.total|Guinea pig epithelium Ab.IgE/IgE.total
C1542892|T201|COMP|39604-4|LNC|Artemisia vulgaris Ab.IgE/IgE.total|Artemisia vulgaris Ab.IgE/IgE.total
C1542893|T201|COMP|39605-1|LNC|Goose feather Ab.IgE/IgE.total|Goose feather Ab.IgE/IgE.total
C1542894|T201|COMP|39606-9|LNC|Rabbit epithelium Ab.IgE/IgE.total|Rabbit epithelium Ab.IgE/IgE.total
C1542895|T201|COMP|39607-7|LNC|Spermatozoa.motile|Spermatozoa.motile
C1542928|T201|COMP|40039-0|LNC|Glucose^27H post XXX challenge|Glucose^27H post XXX challenge
C1542929|T201|COMP|40040-8|LNC|Glucose^28H post XXX challenge|Glucose^28H post XXX challenge
C1542930|T201|COMP|40041-6|LNC|Glucose^29H post XXX challenge|Glucose^29H post XXX challenge
C1542931|T201|COMP|40042-4|LNC|Glucose^30H post XXX challenge|Glucose^30H post XXX challenge
C1542932|T201|COMP|40043-2|LNC|Glucose^31H post XXX challenge|Glucose^31H post XXX challenge
C1542933|T201|COMP|40044-0|LNC|Glucose^36H post XXX challenge|Glucose^36H post XXX challenge
C1542934|T201|COMP|40045-7|LNC|Glucose^2D post XXX challenge|Glucose^2D post XXX challenge
C1542935|T201|COMP|40046-5|LNC|Albumin^pre XXX challenge|Albumin^pre XXX challenge
C1542936|T201|COMP|40047-3|LNC|Albumin^45M pre XXX challenge|Albumin^45M pre XXX challenge
C1542938|T201|COMP|40112-5|LNC|Creatinine^pre XXX challenge|Creatinine^pre XXX challenge
C1542939|T201|COMP|40113-3|LNC|Creatinine^1.5H pre XXX challenge|Creatinine^1.5H pre XXX challenge
C1542940|T201|COMP|40114-1|LNC|Creatinine^1H pre XXX challenge|Creatinine^1H pre XXX challenge
C1542941|T201|COMP|40115-8|LNC|Creatinine^45M pre XXX challenge|Creatinine^45M pre XXX challenge
C1542942|T201|COMP|40116-6|LNC|Creatinine^30M pre XXX challenge|Creatinine^30M pre XXX challenge
C1542943|T201|COMP|40117-4|LNC|Creatinine^45M post XXX challenge|Creatinine^45M post XXX challenge
C1542944|T201|COMP|40118-2|LNC|Creatinine^3.5H post XXX challenge|Creatinine^3.5H post XXX challenge
C1542945|T201|COMP|40119-0|LNC|Creatinine^4H post XXX challenge|Creatinine^4H post XXX challenge
C1542946|T201|COMP|40202-4|LNC|Glucose^8M post XXX challenge|Glucose^8M post XXX challenge
C1542947|T201|COMP|40203-2|LNC|Glucose^9M post XXX challenge|Glucose^9M post XXX challenge
C1542948|T201|COMP|40204-0|LNC|Glucose^12M post XXX challenge|Glucose^12M post XXX challenge
C1542949|T201|COMP|40205-7|LNC|Glucose^14M post XXX challenge|Glucose^14M post XXX challenge
C1542950|T201|COMP|40206-5|LNC|Glucose^16M post XXX challenge|Glucose^16M post XXX challenge
C1542951|T201|COMP|40207-3|LNC|Glucose^19M post XXX challenge|Glucose^19M post XXX challenge
C1542952|T201|COMP|40208-1|LNC|Glucose^22M post XXX challenge|Glucose^22M post XXX challenge
C1542953|T201|COMP|40209-9|LNC|Glucose^25M post XXX challenge|Glucose^25M post XXX challenge
C1542954|T201|COMP|40210-7|LNC|Glucose^27M post XXX challenge|Glucose^27M post XXX challenge
C1542955|T201|COMP|38894-2|LNC|Cells.CD158|Cells.CD158
C1542956|T201|COMP|38895-9|LNC|ELA2 gene targeted mutation analysis|ELA2 gene targeted mutation analysis
C1542957|T201|COMP|38896-7|LNC|F9 gene targeted mutation analysis|F9 gene targeted mutation analysis
C1542958|T201|COMP|38897-5|LNC|Fibers|Fibers
C1542959|T201|COMP|38898-3|LNC|Fibrin D-dimer|Fibrin D-dimer
C1542960|T201|COMP|38899-1|LNC|fluPHENAZine|fluPHENAZine
C1542961|T201|COMP|38900-7|LNC|HEXA gene mutations tested for|HEXA gene mutations tested for
C1542962|T201|COMP|38901-5|LNC|Leflunomide|Leflunomide
C1542963|T201|COMP|38902-3|LNC|LITAF gene targeted mutation analysis|LITAF gene targeted mutation analysis
C1542964|T201|COMP|38903-1|LNC|Lymphocytes|Lymphocytes
C1542980|T201|COMP|40163-8|LNC|Glucose^4H post XXX challenge|Glucose^4H post XXX challenge
C1542981|T201|COMP|40164-6|LNC|Glucose^5H post XXX challenge|Glucose^5H post XXX challenge
C1542982|T201|COMP|40165-3|LNC|Glucose^6H post XXX challenge|Glucose^6H post XXX challenge
C1542983|T201|COMP|40166-1|LNC|Glucose^6.5H post XXX challenge|Glucose^6.5H post XXX challenge
C1542984|T201|COMP|40167-9|LNC|Glucose^7H post XXX challenge|Glucose^7H post XXX challenge
C1542985|T201|COMP|40168-7|LNC|Glucose^7.5H post XXX challenge|Glucose^7.5H post XXX challenge
C1542986|T201|COMP|40169-5|LNC|Glucose^8H post XXX challenge|Glucose^8H post XXX challenge
C1542987|T201|COMP|40170-3|LNC|Glucose^8.5H post XXX challenge|Glucose^8.5H post XXX challenge
C1542988|T201|COMP|40171-1|LNC|Glucose^9H post XXX challenge|Glucose^9H post XXX challenge
C1542989|T201|COMP|40524-1|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C1542990|T201|COMP|40525-8|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C1542991|T201|COMP|40526-6|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C1542992|T201|COMP|40527-4|LNC|Cocaine|Cocaine
C1542993|T201|COMP|40528-2|LNC|Opiates|Opiates
C1542994|T201|COMP|40529-0|LNC|Amphetamines|Amphetamines
C1542995|T201|COMP|40530-8|LNC|Ethanol|Ethanol
C1542996|T201|COMP|40531-6|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C1542997|T201|COMP|40532-4|LNC|Methanol|Methanol
C1542998|T201|COMP|40533-2|LNC|Leukocytes|Leukocytes
C1542999|T201|COMP|40909-4|LNC|Streptococcus pneumoniae 4 Ab.IgG^1st specimen|Streptococcus pneumoniae 4 Ab.IgG^1st specimen
C1543000|T201|COMP|40910-2|LNC|Streptococcus pneumoniae 4 Ab.IgG^2nd specimen|Streptococcus pneumoniae 4 Ab.IgG^2nd specimen
C1543007|T201|COMP|38875-1|LNC|Coagulation tissue factor induced.INR|Coagulation tissue factor induced.INR
C1543023|T201|COMP|38891-8|LNC|ABCC8 gene targeted mutation analysis|ABCC8 gene targeted mutation analysis
C1543024|T201|COMP|38892-6|LNC|Anisocytosis|Anisocytosis
C1543025|T201|COMP|38893-4|LNC|ARIPiprazole|ARIPiprazole
C1543026|T201|COMP|38904-9|LNC|MFN2 gene targeted mutation analysis|MFN2 gene targeted mutation analysis
C1543027|T201|COMP|38905-6|LNC|MLL gene mutations tested for|MLL gene mutations tested for
C1543028|T201|COMP|38906-4|LNC|MSH6 gene targeted mutation analysis|MSH6 gene targeted mutation analysis
C1543029|T201|COMP|38907-2|LNC|NIPA1 gene targeted mutation analysis|NIPA1 gene targeted mutation analysis
C1543030|T201|COMP|38908-0|LNC|Poikilocytosis|Poikilocytosis
C1543031|T201|COMP|38909-8|LNC|PTCH gene targeted mutation analysis|PTCH gene targeted mutation analysis
C1543032|T201|COMP|38910-6|LNC|Schistocytes|Schistocytes
C1543033|T201|COMP|38911-4|LNC|SDHC gene targeted mutation analysis|SDHC gene targeted mutation analysis
C1543034|T201|COMP|38912-2|LNC|Succinylacetone|Succinylacetone
C1543035|T201|COMP|38913-0|LNC|TBX5 gene targeted mutation analysis|TBX5 gene targeted mutation analysis
C1543036|T201|COMP|38914-8|LNC|RS1 gene targeted mutation analysis|RS1 gene targeted mutation analysis
C1543037|T201|COMP|38915-5|LNC|Zinc finger protein of the cerebellum 4 Ab|Zinc finger protein of the cerebellum 4 Ab
C1543038|T201|COMP|38916-3|LNC|Calicivirus RNA|Calicivirus RNA
C1543039|T201|COMP|38917-1|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C1543040|T201|COMP|38918-9|LNC|ABCC8 gene targeted mutation analysis|ABCC8 gene targeted mutation analysis
C1543041|T201|COMP|38919-7|LNC|LITAF gene targeted mutation analysis|LITAF gene targeted mutation analysis
C1543042|T201|COMP|38920-5|LNC|MFN2 gene targeted mutation analysis|MFN2 gene targeted mutation analysis
C1543043|T201|COMP|38921-3|LNC|MSH6 gene targeted mutation analysis|MSH6 gene targeted mutation analysis
C1543044|T201|COMP|38922-1|LNC|PTCH gene targeted mutation analysis|PTCH gene targeted mutation analysis
C1543045|T201|COMP|38923-9|LNC|SDHC gene targeted mutation analysis|SDHC gene targeted mutation analysis
C1543046|T201|COMP|38924-7|LNC|TBX5 gene targeted mutation analysis|TBX5 gene targeted mutation analysis
C1543047|T201|COMP|38925-4|LNC|RS1 gene targeted mutation analysis|RS1 gene targeted mutation analysis
C1543048|T201|COMP|38926-2|LNC|Macroprolactin|Macroprolactin
C1543049|T201|COMP|38927-0|LNC|TRPS1 gene targeted mutation analysis|TRPS1 gene targeted mutation analysis
C1543050|T201|COMP|38928-8|LNC|FAH gene targeted mutation analysis|FAH gene targeted mutation analysis
C1543051|T201|COMP|38929-6|LNC|FAH gene targeted mutation analysis|FAH gene targeted mutation analysis
C1543052|T201|COMP|38930-4|LNC|EXT1 gene targeted mutation analysis|EXT1 gene targeted mutation analysis
C1543053|T201|COMP|38931-2|LNC|TRPS1 gene targeted mutation analysis|TRPS1 gene targeted mutation analysis
C1543111|T201|COMP|38989-0|LNC|Clostridium botulinum toxin A+B+E+F+G|Clostridium botulinum toxin A+B+E+F+G
C1543112|T201|COMP|38990-8|LNC|Escherichia coli O157:H7 DNA|Escherichia coli O157:H7 DNA
C1543113|T201|COMP|38991-6|LNC|Amylase|Amylase
C1543114|T201|COMP|38992-4|LNC|Amylase|Amylase
C1543115|T201|COMP|38993-2|LNC|Calcium oxalate dihydrate crystals|Calcium oxalate dihydrate crystals
C1543116|T201|COMP|38994-0|LNC|Histiocytes|Histiocytes
C1543117|T201|COMP|38995-7|LNC|Mixed cellular casts|Mixed cellular casts
C1543118|T201|COMP|38996-5|LNC|Neutrophils|Neutrophils
C1543119|T201|COMP|38997-3|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C1543120|T201|COMP|38998-1|LNC|HIV 1+Hepatitis C virus RNA|HIV 1+Hepatitis C virus RNA
C1543122|T201|COMP|39000-5|LNC|3-Hydroxybutyrylcarnitine (C4-OH)|3-Hydroxybutyrylcarnitine (C4-OH)
C1543123|T201|COMP|39001-3|LNC|3-Hydroxyisovalerylcarnitine (C5-OH)|3-Hydroxyisovalerylcarnitine (C5-OH)
C1543124|T201|COMP|39002-1|LNC|Adipoylcarnitine (C6-DC)|Adipoylcarnitine (C6-DC)
C1543125|T201|COMP|39003-9|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1543126|T201|COMP|39004-7|LNC|Epidermal growth factor receptor Ag|Epidermal growth factor receptor Ag
C1543127|T201|COMP|39005-4|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C1543128|T201|COMP|39006-2|LNC|Hepatitis B virus little e Ab|Hepatitis B virus little e Ab
C1543129|T201|COMP|39007-0|LNC|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C1543130|T201|COMP|39008-8|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C1543131|T201|COMP|39009-6|LNC|Isovalerylcarnitine (C5)|Isovalerylcarnitine (C5)
C1543132|T201|COMP|39010-4|LNC|Methylmalonylcarnitine (C4-DC)|Methylmalonylcarnitine (C4-DC)
C1543133|T201|COMP|39011-2|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C1543134|T201|COMP|39012-0|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C1543135|T201|COMP|39013-8|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C1543136|T201|COMP|39014-6|LNC|Suberylcarnitine (C8-DC)|Suberylcarnitine (C8-DC)
C1543137|T201|COMP|39015-3|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1543138|T201|COMP|39016-1|LNC|Age at death|Age at death
C1543140|T201|COMP|39019-5|LNC|Escherichia coli O157:H7 Ag|Escherichia coli O157:H7 Ag
C1543141|T201|COMP|39020-3|LNC|Prion protein.abnormal|Prion protein.abnormal
C1543142|T201|COMP|39021-1|LNC|Prion protein.abnormal|Prion protein.abnormal
C1543143|T201|COMP|39022-9|LNC|Sarcocystis neurona Ab|Sarcocystis neurona Ab
C1543144|T201|COMP|39023-7|LNC|Vesicular stomatitis Indiana virus RNA|Vesicular stomatitis Indiana virus RNA
C1543145|T201|COMP|39024-5|LNC|Vesicular stomatitis New Jersey virus RNA|Vesicular stomatitis New Jersey virus RNA
C1543146|T201|COMP|39025-2|LNC|Influenza virus A hemagglutinin cDNA|Influenza virus A hemagglutinin cDNA
C1543201|T201|COMP|39080-7|LNC|EPM2A gene targeted mutation analysis|EPM2A gene targeted mutation analysis
C1543202|T201|COMP|39081-5|LNC|Gadus morhua Ab.IgE/IgE.total|Gadus morhua Ab.IgE/IgE.total
C1543203|T201|COMP|39082-3|LNC|Gentamicin^peak|Gentamicin^peak
C1543204|T201|COMP|39083-1|LNC|Herpes virus 8 Ab|Herpes virus 8 Ab
C1543205|T201|COMP|39084-9|LNC|Iva ciliata Ab.IgE/IgE.total|Iva ciliata Ab.IgE/IgE.total
C1543206|T201|COMP|39085-6|LNC|Juglans california pollen Ab.IgE/IgE.total|Juglans california pollen Ab.IgE/IgE.total
C1543208|T201|COMP|39087-2|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C1543209|T201|COMP|39088-0|LNC|Pecten spp Ab.IgE/IgE.total|Pecten spp Ab.IgE/IgE.total
C1543210|T201|COMP|39089-8|LNC|PLP1 gene targeted mutation analysis|PLP1 gene targeted mutation analysis
C1543211|T201|COMP|39090-6|LNC|Ruditapes spp Ab.IgE/IgE.total|Ruditapes spp Ab.IgE/IgE.total
C1543212|T201|COMP|39091-4|LNC|Sorghum halepense Ab.IgE/IgE.total|Sorghum halepense Ab.IgE/IgE.total
C1543213|T201|COMP|39092-2|LNC|Vancomycin^peak|Vancomycin^peak
C1543223|T201|COMP|39102-9|LNC|Influenza virus A hemagglutinin cDNA|Influenza virus A hemagglutinin cDNA
C1543224|T201|COMP|39103-7|LNC|Influenza virus A neuraminidase cDNA|Influenza virus A neuraminidase cDNA
C1543381|T201|COMP|39295-1|LNC|Influenza virus A Ab|Influenza virus A Ab
C1543382|T201|COMP|39296-9|LNC|Influenza virus A H1 Ab|Influenza virus A H1 Ab
C1543383|T201|COMP|39297-7|LNC|Influenza virus A H10 Ab|Influenza virus A H10 Ab
C1543384|T201|COMP|39298-5|LNC|Influenza virus A H11 Ab|Influenza virus A H11 Ab
C1543385|T201|COMP|39299-3|LNC|Influenza virus A H12 Ab|Influenza virus A H12 Ab
C1543386|T201|COMP|39300-9|LNC|Influenza virus A H13 Ab|Influenza virus A H13 Ab
C1543387|T201|COMP|39301-7|LNC|Influenza virus A H14 Ab|Influenza virus A H14 Ab
C1543388|T201|COMP|39302-5|LNC|Influenza virus A H15 Ab|Influenza virus A H15 Ab
C1543389|T201|COMP|39303-3|LNC|Influenza virus A H2 Ab|Influenza virus A H2 Ab
C1543390|T201|COMP|39304-1|LNC|Influenza virus A H3 Ab|Influenza virus A H3 Ab
C1543391|T201|COMP|39305-8|LNC|Influenza virus A H4 Ab|Influenza virus A H4 Ab
C1543392|T201|COMP|39306-6|LNC|Influenza virus A H5 Ab|Influenza virus A H5 Ab
C1543393|T201|COMP|39307-4|LNC|Influenza virus A H6 Ab|Influenza virus A H6 Ab
C1543394|T201|COMP|39308-2|LNC|Influenza virus A H7 Ab|Influenza virus A H7 Ab
C1543395|T201|COMP|39309-0|LNC|Influenza virus A H8 Ab|Influenza virus A H8 Ab
C1543396|T201|COMP|39310-8|LNC|Influenza virus A H9 Ab|Influenza virus A H9 Ab
C1543397|T201|COMP|39311-6|LNC|Influenza virus A N1 Ab|Influenza virus A N1 Ab
C1543398|T201|COMP|39312-4|LNC|Influenza virus A N2 Ab|Influenza virus A N2 Ab
C1543399|T201|COMP|39313-2|LNC|Influenza virus A N3 Ab|Influenza virus A N3 Ab
C1543400|T201|COMP|39314-0|LNC|Influenza virus A N4 Ab|Influenza virus A N4 Ab
C1543401|T201|COMP|39315-7|LNC|Influenza virus A N5 Ab|Influenza virus A N5 Ab
C1543402|T201|COMP|39316-5|LNC|Influenza virus A N6 Ab|Influenza virus A N6 Ab
C1543403|T201|COMP|39317-3|LNC|Influenza virus A N7 Ab|Influenza virus A N7 Ab
C1543404|T201|COMP|39318-1|LNC|Influenza virus A N8 Ab|Influenza virus A N8 Ab
C1543405|T201|COMP|39319-9|LNC|Influenza virus A N9 Ab|Influenza virus A N9 Ab
C1543406|T201|COMP|39320-7|LNC|Prion protein.abnormal|Prion protein.abnormal
C1543439|T201|COMP|39354-6|LNC|Cholinesterase^dibucaine/Cholinesterase|Cholinesterase^dibucaine/Cholinesterase
C1543440|T201|COMP|39355-3|LNC|Cholinesterase.fluoride inhibited/Cholinesterase|Cholinesterase.fluoride inhibited/Cholinesterase
C1543441|T201|COMP|39356-1|LNC|Cholinesterase.scoline inhibited/Cholinesterase|Cholinesterase.scoline inhibited/Cholinesterase
C1543442|T201|COMP|39357-9|LNC|Cholinesterase.chloride inhibited/Cholinesterase|Cholinesterase.chloride inhibited/Cholinesterase
C1543443|T201|COMP|39358-7|LNC|Cholinesterase.RO 020683 inhibited/Cholinesterase|Cholinesterase.RO 020683 inhibited/Cholinesterase
C1543531|T201|COMP|39455-1|LNC|9-Hydroxyrisperidone|9-Hydroxyrisperidone
C1543532|T201|COMP|39456-9|LNC|Acetaminophen|Acetaminophen
C1543533|T201|COMP|39457-7|LNC|Beta aminobutyrate|Beta aminobutyrate
C1543534|T201|COMP|39458-5|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C1543535|T201|COMP|39459-3|LNC|Bicarbonate^^standard|Bicarbonate^^standard
C1543536|T201|COMP|39460-1|LNC|Bicarbonate^^standard|Bicarbonate^^standard
C1543537|T201|COMP|39461-9|LNC|Bilirubin|Bilirubin
C1543538|T201|COMP|39462-7|LNC|Bilirubin.glucuronidated|Bilirubin.glucuronidated
C1543539|T201|COMP|39463-5|LNC|Bilirubin.non-glucuronidated|Bilirubin.non-glucuronidated
C1543540|T201|COMP|39464-3|LNC|Carbon dioxide|Carbon dioxide
C1543541|T201|COMP|39465-0|LNC|Carbon dioxide|Carbon dioxide
C1543542|T201|COMP|39466-8|LNC|Carbon dioxide|Carbon dioxide
C1543543|T201|COMP|39467-6|LNC|Chloride|Chloride
C1543544|T201|COMP|39468-4|LNC|Cholesterol|Cholesterol
C1543545|T201|COMP|39469-2|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C1543546|T201|COMP|39470-0|LNC|Prochlorperazine|Prochlorperazine
C1543547|T201|COMP|39471-8|LNC|Creatinine|Creatinine
C1543548|T201|COMP|39472-6|LNC|Creatinine|Creatinine
C1543549|T201|COMP|39473-4|LNC|Creatinine|Creatinine
C1543550|T201|COMP|39474-2|LNC|Creatinine|Creatinine
C1543551|T201|COMP|39475-9|LNC|dimenhyDRINATE|dimenhyDRINATE
C1543552|T201|COMP|39476-7|LNC|diphenhydrAMINE|diphenhydrAMINE
C1543553|T201|COMP|39477-5|LNC|fluPHENAZine|fluPHENAZine
C1543554|T201|COMP|39478-3|LNC|Glucose|Glucose
C1543555|T201|COMP|39479-1|LNC|Glucose|Glucose
C1543556|T201|COMP|39480-9|LNC|Glucose|Glucose
C1543557|T201|COMP|39481-7|LNC|Glucose|Glucose
C1543558|T201|COMP|39482-5|LNC|Trimeprazine|Trimeprazine
C1543559|T201|COMP|39483-3|LNC|Normethsuximide|Normethsuximide
C1543560|T201|COMP|39484-1|LNC|OLANZapine|OLANZapine
C1543561|T201|COMP|39485-8|LNC|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1543562|T201|COMP|39486-6|LNC|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1543563|T201|COMP|39487-4|LNC|PHENobarbital|PHENobarbital
C1543564|T201|COMP|39488-2|LNC|Phensuximide|Phensuximide
C1543603|T201|COMP|39528-5|LNC|Adenovirus DNA|Adenovirus DNA
C1543604|T201|COMP|39529-3|LNC|Acetone|Acetone
C1543605|T201|COMP|39530-1|LNC|Isopropanol|Isopropanol
C1543606|T201|COMP|39531-9|LNC|Acetaldehyde|Acetaldehyde
C1543607|T201|COMP|39532-7|LNC|Inhibin B|Inhibin B
C1543608|T201|COMP|39533-5|LNC|Deoxyhemoglobin|Deoxyhemoglobin
C1543609|T201|COMP|39534-3|LNC|Cryptosporidium sp Ag|Cryptosporidium sp Ag
C1543610|T201|COMP|39535-0|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C1543611|T201|COMP|39536-8|LNC|Influenza virus A Ab|Influenza virus A Ab
C1543612|T201|COMP|39537-6|LNC|Influenza virus B Ab|Influenza virus B Ab
C1543613|T201|COMP|39538-4|LNC|Finch droppings Ab.IgG|Finch droppings Ab.IgG
C1543614|T201|COMP|39539-2|LNC|Cockatiel droppings Ab.IgG|Cockatiel droppings Ab.IgG
C1543615|T201|COMP|39540-0|LNC|Uranium/Creatinine|Uranium/Creatinine
C1543616|T201|COMP|39541-8|LNC|Legionella sp Ag|Legionella sp Ag
C1543617|T201|COMP|39542-6|LNC|Prunus dulcis Ab.IgE/IgE.total|Prunus dulcis Ab.IgE/IgE.total
C1543618|T201|COMP|39543-4|LNC|Corylus avellana Ab.IgE/IgE.total|Corylus avellana Ab.IgE/IgE.total
C1543619|T201|COMP|39544-2|LNC|Dolichovespula arenaria Ab.IgE/IgE.total|Dolichovespula arenaria Ab.IgE/IgE.total
C1543620|T201|COMP|39545-9|LNC|Cancer pagurus Ab.IgE/IgE.total|Cancer pagurus Ab.IgE/IgE.total
C1543621|T201|COMP|39546-7|LNC|Homarus gammarus Ab.IgE/IgE.total|Homarus gammarus Ab.IgE/IgE.total
C1543622|T201|COMP|39547-5|LNC|Thunnus albacares Ab.IgE/IgE.total|Thunnus albacares Ab.IgE/IgE.total
C1543623|T201|COMP|39548-3|LNC|Salmo salar Ab.IgE/IgE.total|Salmo salar Ab.IgE/IgE.total
C1543624|T201|COMP|39549-1|LNC|Helix aspersa Ab.IgE/IgE.total|Helix aspersa Ab.IgE/IgE.total
C1543625|T201|COMP|39550-9|LNC|Horse dander Ab.IgE/IgE.total|Horse dander Ab.IgE/IgE.total
C1543626|T201|COMP|39551-7|LNC|Cow dander Ab.IgE/IgE.total|Cow dander Ab.IgE/IgE.total
C1543627|T201|COMP|39552-5|LNC|Lamb Ab.IgE/IgE.total|Lamb Ab.IgE/IgE.total
C1543628|T201|COMP|39553-3|LNC|Penicillin V Ab.IgE/IgE.total|Penicillin V Ab.IgE/IgE.total
C1543629|T201|COMP|39554-1|LNC|Endomysium Ab.IgG|Endomysium Ab.IgG
C1543630|T201|COMP|39555-8|LNC|West Nile virus Ab|West Nile virus Ab
C1543631|T201|COMP|39556-6|LNC|Coagulation factor X inhibitor|Coagulation factor X inhibitor
C1543632|T201|COMP|39557-4|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1543633|T201|COMP|39558-2|LNC|West Nile virus Ab|West Nile virus Ab
C1543634|T201|COMP|39559-0|LNC|Legionella sp Ab.IgM|Legionella sp Ab.IgM
C1543635|T201|COMP|39560-8|LNC|Sulfate.inorganic|Sulfate.inorganic
C1543636|T201|COMP|39561-6|LNC|Glucose^1st specimen post dose lactose|Glucose^1st specimen post dose lactose
C1543637|T201|COMP|39562-4|LNC|Glucose^2nd specimen post dose lactose|Glucose^2nd specimen post dose lactose
C1543638|T201|COMP|39563-2|LNC|Glucose^3rd specimen post dose lactose|Glucose^3rd specimen post dose lactose
C1543639|T201|COMP|39564-0|LNC|Corticotropin^1st specimen post XXX challenge|Corticotropin^1st specimen post XXX challenge
C1543640|T201|COMP|39565-7|LNC|Complement C4d|Complement C4d
C1543641|T201|COMP|39566-5|LNC|Pregnanetriol/Creatinine|Pregnanetriol/Creatinine
C1543642|T201|COMP|39567-3|LNC|TOLAZamide|TOLAZamide
C1543643|T201|COMP|39568-1|LNC|TOLBUTamide|TOLBUTamide
C1543644|T201|COMP|39569-9|LNC|Trichoderma viride Ab|Trichoderma viride Ab
C1543645|T201|COMP|39570-7|LNC|Alternaria sp Ab.IgG|Alternaria sp Ab.IgG
C1543646|T201|COMP|39571-5|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1543647|T201|COMP|39572-3|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C1543648|T201|COMP|39573-1|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1543649|T201|COMP|39574-9|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C1543650|T201|COMP|39575-6|LNC|Fungus.microscopic observation|Fungus.microscopic observation
C1543651|T201|COMP|39576-4|LNC|Sulfate|Sulfate
C1543652|T201|COMP|39577-2|LNC|Leishmania sp Ab.IgM|Leishmania sp Ab.IgM
C1543653|T201|COMP|39578-0|LNC|Alternaria alternata Ab|Alternaria alternata Ab
C1543654|T201|COMP|39579-8|LNC|Penicillium notatum Ab|Penicillium notatum Ab
C1543655|T201|COMP|39580-6|LNC|Phoma herbarum Ab|Phoma herbarum Ab
C1543656|T201|COMP|39581-4|LNC|Rubella virus Ab|Rubella virus Ab
C1543657|T201|COMP|39582-2|LNC|Amino beta guanidinopropionate/Creatinine|Amino beta guanidinopropionate/Creatinine
C1543658|T201|COMP|39583-0|LNC|Mercury|Mercury
C1543659|T201|COMP|39584-8|LNC|Mercury|Mercury
C1543660|T201|COMP|39585-5|LNC|Tritium|Tritium
C1543661|T201|COMP|39586-3|LNC|Disialylganglioside GD1b Ab|Disialylganglioside GD1b Ab
C1543662|T201|COMP|39587-1|LNC|Neutrophil Ab|Neutrophil Ab
C1543663|T201|COMP|39588-9|LNC|Histoplasma capsulatum Ab.IgG|Histoplasma capsulatum Ab.IgG
C1543664|T201|COMP|39589-7|LNC|HTLV I p19 Ab|HTLV I p19 Ab
C1543665|T201|COMP|39590-5|LNC|HTLV I+II p19 Ab|HTLV I+II p19 Ab
C1543666|T201|COMP|39591-3|LNC|PARoxetine|PARoxetine
C1543667|T201|COMP|39592-1|LNC|Bertholletia excelsa Ab.IgE/IgE.total|Bertholletia excelsa Ab.IgE/IgE.total
C1543668|T201|COMP|39593-9|LNC|Cocos nucifera Ab.IgE/IgE.total|Cocos nucifera Ab.IgE/IgE.total
C1543669|T201|COMP|39594-7|LNC|Carya illinoinensis nut Ab.IgE/IgE.total|Carya illinoinensis nut Ab.IgE/IgE.total
C1543670|T201|COMP|39608-5|LNC|Spermatozoa.immotile|Spermatozoa.immotile
C1543671|T201|COMP|39609-3|LNC|Vaccinium myrtillus Ab.IgE/IgE.total|Vaccinium myrtillus Ab.IgE/IgE.total
C1543672|T201|COMP|39610-1|LNC|Neisseria meningitidis serogroup w135 Ab|Neisseria meningitidis serogroup w135 Ab
C1543673|T201|COMP|39611-9|LNC|Silicone Ab.IgG|Silicone Ab.IgG
C1543674|T201|COMP|39612-7|LNC|Silicone Ab.IgA|Silicone Ab.IgA
C1543675|T201|COMP|39613-5|LNC|Silicone Ab.IgM|Silicone Ab.IgM
C1543676|T201|COMP|39614-3|LNC|Silicone Ab.IgE|Silicone Ab.IgE
C1543677|T201|COMP|39615-0|LNC|Benzoylcarnitine (BzCn)|Benzoylcarnitine (BzCn)
C1543678|T201|COMP|39616-8|LNC|Palmitoylcarnitine|Palmitoylcarnitine
C1543679|T201|COMP|39617-6|LNC|3-Hydroxypalmitoylcarnitine|3-Hydroxypalmitoylcarnitine
C1543680|T201|COMP|39618-4|LNC|Neisseria meningitidis serogroup Y Ab|Neisseria meningitidis serogroup Y Ab
C1543813|T201|COMP|39771-1|LNC|Porphyrins|Porphyrins
C1543814|T201|COMP|39772-9|LNC|Sulfamethoxazole|Sulfamethoxazole
C1543815|T201|COMP|39773-7|LNC|Beta-2-Microglobulin/Creatinine|Beta-2-Microglobulin/Creatinine
C1543816|T201|COMP|39774-5|LNC|Porphyrins|Porphyrins
C1543817|T201|COMP|39775-2|LNC|Protoporphyrin.free|Protoporphyrin.free
C1543818|T201|COMP|39776-0|LNC|Urea^post dialysis|Urea^post dialysis
C1543819|T201|COMP|39777-8|LNC|Urea^pre dialysis|Urea^pre dialysis
C1543820|T201|COMP|39778-6|LNC|Iron/Iron binding capacity.total|Iron/Iron binding capacity.total
C1543821|T201|COMP|39779-4|LNC|Urea|Urea
C1543822|T201|COMP|39780-2|LNC|Urea|Urea
C1543823|T201|COMP|39781-0|LNC|Urea|Urea
C1543824|T201|COMP|39782-8|LNC|Delta aminolevulinate/Creatinine|Delta aminolevulinate/Creatinine
C1543825|T201|COMP|39783-6|LNC|Urea/Creatinine|Urea/Creatinine
C1543826|T201|COMP|39784-4|LNC|Porphyrins|Porphyrins
C1543827|T201|COMP|39785-1|LNC|Potassium|Potassium
C1543828|T201|COMP|39786-9|LNC|Pyridoxine|Pyridoxine
C1543829|T201|COMP|39787-7|LNC|Sodium|Sodium
C1543830|T201|COMP|39788-5|LNC|Urate|Urate
C1543831|T201|COMP|39789-3|LNC|Potassium|Potassium
C1543832|T201|COMP|39790-1|LNC|Potassium|Potassium
C1543833|T201|COMP|39791-9|LNC|Sodium|Sodium
C1543834|T201|COMP|39792-7|LNC|Sodium|Sodium
C1543835|T201|COMP|39793-5|LNC|Coproporphyrin 3/Coproporphyrin 1|Coproporphyrin 3/Coproporphyrin 1
C1543836|T201|COMP|39794-3|LNC|Tocainide|Tocainide
C1543837|T201|COMP|39795-0|LNC|Trifluoperazine|Trifluoperazine
C1543838|T201|COMP|39796-8|LNC|Vancomycin^peak|Vancomycin^peak
C1543839|T201|COMP|39797-6|LNC|Vancomycin^trough|Vancomycin^trough
C1543840|T201|COMP|39798-4|LNC|Warfarin|Warfarin
C1543841|T201|COMP|39799-2|LNC|risperiDONE|risperiDONE
C1543842|T201|COMP|39800-8|LNC|Risperidone+9-Hydroxyrisperidone|Risperidone+9-Hydroxyrisperidone
C1543843|T201|COMP|39801-6|LNC|Triglyceride|Triglyceride
C1543844|T201|COMP|39802-4|LNC|Creatinine dial fld/Creatinine ser_plas|Creatinine dial fld/Creatinine ser_plas
C1543845|T201|COMP|39803-2|LNC|inFLIXimab|inFLIXimab
C1543846|T201|COMP|39804-0|LNC|Lipoprotein associated phospholipase A2|Lipoprotein associated phospholipase A2
C1543847|T201|COMP|39805-7|LNC|Rabbit hair Ab.IgE|Rabbit hair Ab.IgE
C1543968|T201|COMP|39955-0|LNC|Creatinine^pre XXX challenge|Creatinine^pre XXX challenge
C1543969|T201|COMP|39956-8|LNC|Creatinine^1.5H pre XXX challenge|Creatinine^1.5H pre XXX challenge
C1543970|T201|COMP|39957-6|LNC|Creatinine^1H pre XXX challenge|Creatinine^1H pre XXX challenge
C1543971|T201|COMP|39958-4|LNC|Creatinine^45M pre XXX challenge|Creatinine^45M pre XXX challenge
C1543972|T201|COMP|39959-2|LNC|Creatinine^30M pre XXX challenge|Creatinine^30M pre XXX challenge
C1543973|T201|COMP|39960-0|LNC|Creatinine^45M post XXX challenge|Creatinine^45M post XXX challenge
C1543974|T201|COMP|39961-8|LNC|Creatinine^3.5H post XXX challenge|Creatinine^3.5H post XXX challenge
C1543975|T201|COMP|39962-6|LNC|Creatinine^3.75H post XXX challenge|Creatinine^3.75H post XXX challenge
C1543976|T201|COMP|39963-4|LNC|Creatinine^4H post XXX challenge|Creatinine^4H post XXX challenge
C1543977|T201|COMP|39964-2|LNC|Creatinine^4.5H post XXX challenge|Creatinine^4.5H post XXX challenge
C1543978|T201|COMP|39965-9|LNC|Creatinine^5.25H post XXX challenge|Creatinine^5.25H post XXX challenge
C1543979|T201|COMP|39966-7|LNC|Creatinine^5.5H post XXX challenge|Creatinine^5.5H post XXX challenge
C1543980|T201|COMP|39967-5|LNC|Creatinine^6.5H post XXX challenge|Creatinine^6.5H post XXX challenge
C1543981|T201|COMP|39968-3|LNC|Creatinine^8H post XXX challenge|Creatinine^8H post XXX challenge
C1543982|T201|COMP|39969-1|LNC|Creatinine^9H post XXX challenge|Creatinine^9H post XXX challenge
C1543983|T201|COMP|39970-9|LNC|Creatinine^10H post XXX challenge|Creatinine^10H post XXX challenge
C1543984|T201|COMP|39971-7|LNC|Creatinine^12H post XXX challenge|Creatinine^12H post XXX challenge
C1543985|T201|COMP|39972-5|LNC|Creatinine^16H post XXX challenge|Creatinine^16H post XXX challenge
C1543986|T201|COMP|39973-3|LNC|Creatinine^18H post XXX challenge|Creatinine^18H post XXX challenge
C1543987|T201|COMP|39974-1|LNC|Creatinine^2D post XXX challenge|Creatinine^2D post XXX challenge
C1543988|T201|COMP|39975-8|LNC|Creatinine^4D post XXX challenge|Creatinine^4D post XXX challenge
C1543989|T201|COMP|39976-6|LNC|Creatinine^7D post XXX challenge|Creatinine^7D post XXX challenge
C1543990|T201|COMP|39977-4|LNC|Creatinine^pre XXX challenge|Creatinine^pre XXX challenge
C1543991|T201|COMP|39978-2|LNC|Creatinine^2.25H pre XXX challenge|Creatinine^2.25H pre XXX challenge
C1543992|T201|COMP|39979-0|LNC|Creatinine^1.5H pre XXX challenge|Creatinine^1.5H pre XXX challenge
C1543993|T201|COMP|39980-8|LNC|Creatinine^1H pre XXX challenge|Creatinine^1H pre XXX challenge
C1543994|T201|COMP|39981-6|LNC|Creatinine^30M pre XXX challenge|Creatinine^30M pre XXX challenge
C1543995|T201|COMP|39982-4|LNC|Creatinine^baseline|Creatinine^baseline
C1543996|T201|COMP|39983-2|LNC|Creatinine^30M post XXX challenge|Creatinine^30M post XXX challenge
C1543997|T201|COMP|39984-0|LNC|Creatinine^1H post XXX challenge|Creatinine^1H post XXX challenge
C1543998|T201|COMP|39985-7|LNC|Creatinine^1.5H post XXX challenge|Creatinine^1.5H post XXX challenge
C1543999|T201|COMP|39986-5|LNC|Creatinine^2H post XXX challenge|Creatinine^2H post XXX challenge
C1544000|T201|COMP|39987-3|LNC|Creatinine^2.5H post XXX challenge|Creatinine^2.5H post XXX challenge
C1544001|T201|COMP|39988-1|LNC|Creatinine^3H post XXX challenge|Creatinine^3H post XXX challenge
C1544002|T201|COMP|39989-9|LNC|Creatinine^3.5H post XXX challenge|Creatinine^3.5H post XXX challenge
C1544003|T201|COMP|39990-7|LNC|Creatinine^4H post XXX challenge|Creatinine^4H post XXX challenge
C1544004|T201|COMP|39991-5|LNC|Creatinine^4.5H post XXX challenge|Creatinine^4.5H post XXX challenge
C1544005|T201|COMP|39992-3|LNC|Creatinine^5H post XXX challenge|Creatinine^5H post XXX challenge
C1544006|T201|COMP|39993-1|LNC|Creatinine^5.5H post XXX challenge|Creatinine^5.5H post XXX challenge
C1544007|T201|COMP|39994-9|LNC|Creatinine^6H post XXX challenge|Creatinine^6H post XXX challenge
C1544008|T201|COMP|39995-6|LNC|Creatinine^8H post XXX challenge|Creatinine^8H post XXX challenge
C1544009|T201|COMP|39996-4|LNC|Creatinine^1D post XXX challenge|Creatinine^1D post XXX challenge
C1544010|T201|COMP|39997-2|LNC|Glucose^pre XXX challenge|Glucose^pre XXX challenge
C1544011|T201|COMP|39998-0|LNC|Glucose^30M pre XXX challenge|Glucose^30M pre XXX challenge
C1544012|T201|COMP|39999-8|LNC|Glucose^15M pre XXX challenge|Glucose^15M pre XXX challenge
C1544013|T201|COMP|40000-2|LNC|Glucose^5M pre XXX challenge|Glucose^5M pre XXX challenge
C1544014|T201|COMP|40001-0|LNC|Glucose^5M post XXX challenge|Glucose^5M post XXX challenge
C1544015|T201|COMP|40002-8|LNC|Glucose^80M post XXX challenge|Glucose^80M post XXX challenge
C1544016|T201|COMP|40003-6|LNC|Glucose^1.5H post XXX challenge|Glucose^1.5H post XXX challenge
C1544017|T201|COMP|40004-4|LNC|Glucose^100M post XXX challenge|Glucose^100M post XXX challenge
C1544018|T201|COMP|40005-1|LNC|Glucose^110M post XXX challenge|Glucose^110M post XXX challenge
C1544019|T201|COMP|40006-9|LNC|Glucose^8.5H post XXX challenge|Glucose^8.5H post XXX challenge
C1544020|T201|COMP|40007-7|LNC|Glucose^9.5H post XXX challenge|Glucose^9.5H post XXX challenge
C1544021|T201|COMP|40008-5|LNC|Glucose^11.5H post XXX challenge|Glucose^11.5H post XXX challenge
C1544022|T201|COMP|40009-3|LNC|Glucose^12.5H post XXX challenge|Glucose^12.5H post XXX challenge
C1544023|T201|COMP|40010-1|LNC|Glucose^13H post XXX challenge|Glucose^13H post XXX challenge
C1544024|T201|COMP|40011-9|LNC|Glucose^13.5H post XXX challenge|Glucose^13.5H post XXX challenge
C1544025|T201|COMP|40012-7|LNC|Glucose^14H post XXX challenge|Glucose^14H post XXX challenge
C1544026|T201|COMP|40013-5|LNC|Glucose^15.5H post XXX challenge|Glucose^15.5H post XXX challenge
C1544027|T201|COMP|40014-3|LNC|Glucose^16H post XXX challenge|Glucose^16H post XXX challenge
C1544028|T201|COMP|40015-0|LNC|Glucose^17.5H post XXX challenge|Glucose^17.5H post XXX challenge
C1544029|T201|COMP|40016-8|LNC|Glucose^18H post XXX challenge|Glucose^18H post XXX challenge
C1544030|T201|COMP|40017-6|LNC|Glucose^18.5H post XXX challenge|Glucose^18.5H post XXX challenge
C1544031|T201|COMP|40018-4|LNC|Glucose^19.5H post XXX challenge|Glucose^19.5H post XXX challenge
C1544032|T201|COMP|40019-2|LNC|Glucose^20H post XXX challenge|Glucose^20H post XXX challenge
C1544033|T201|COMP|40020-0|LNC|Glucose^20.5H post XXX challenge|Glucose^20.5H post XXX challenge
C1544034|T201|COMP|40021-8|LNC|Glucose^21.5H post XXX challenge|Glucose^21.5H post XXX challenge
C1544035|T201|COMP|40022-6|LNC|Glucose^22H post XXX challenge|Glucose^22H post XXX challenge
C1544036|T201|COMP|40023-4|LNC|Glucose^23.5H post XXX challenge|Glucose^23.5H post XXX challenge
C1544037|T201|COMP|40024-2|LNC|Glucose^1D post XXX challenge|Glucose^1D post XXX challenge
C1544038|T201|COMP|40025-9|LNC|Glucose^3M post XXX challenge|Glucose^3M post XXX challenge
C1544039|T201|COMP|40026-7|LNC|Glucose^ 6M post XXX challenge|Glucose^ 6M post XXX challenge
C1544040|T201|COMP|40027-5|LNC|Glucose^9M post XXX challenge|Glucose^9M post XXX challenge
C1544041|T201|COMP|40028-3|LNC|Glucose^12M post XXX challenge|Glucose^12M post XXX challenge
C1544042|T201|COMP|40029-1|LNC|Glucose^14M post XXX challenge|Glucose^14M post XXX challenge
C1544043|T201|COMP|40030-9|LNC|Glucose^16M post XXX challenge|Glucose^16M post XXX challenge
C1544044|T201|COMP|40031-7|LNC|Glucose^19M post XXX challenge|Glucose^19M post XXX challenge
C1544045|T201|COMP|40032-5|LNC|Glucose^22M post XXX challenge|Glucose^22M post XXX challenge
C1544046|T201|COMP|40033-3|LNC|Glucose^25M post XXX challenge|Glucose^25M post XXX challenge
C1544047|T201|COMP|40034-1|LNC|Glucose^27M post XXX challenge|Glucose^27M post XXX challenge
C1544048|T201|COMP|40035-8|LNC|Glucose^4.5H post XXX challenge|Glucose^4.5H post XXX challenge
C1544049|T201|COMP|40036-6|LNC|Glucose^5.5H post XXX challenge|Glucose^5.5H post XXX challenge
C1544050|T201|COMP|40037-4|LNC|Glucose^25H post XXX challenge|Glucose^25H post XXX challenge
C1544051|T201|COMP|40038-2|LNC|Glucose^26H post XXX challenge|Glucose^26H post XXX challenge
C1544052|T201|COMP|40048-1|LNC|Albumin^30M post XXX challenge|Albumin^30M post XXX challenge
C1544053|T201|COMP|40049-9|LNC|Albumin^45M post XXX challenge|Albumin^45M post XXX challenge
C1544054|T201|COMP|40050-7|LNC|Albumin^1H post XXX challenge|Albumin^1H post XXX challenge
C1544055|T201|COMP|40051-5|LNC|Albumin^1.5H post XXX challenge|Albumin^1.5H post XXX challenge
C1544056|T201|COMP|40052-3|LNC|Albumin^2H post XXX challenge|Albumin^2H post XXX challenge
C1544057|T201|COMP|40053-1|LNC|Albumin^3H post XXX challenge|Albumin^3H post XXX challenge
C1544058|T201|COMP|40054-9|LNC|Albumin^4H post XXX challenge|Albumin^4H post XXX challenge
C1544059|T201|COMP|40055-6|LNC|Albumin^5H post XXX challenge|Albumin^5H post XXX challenge
C1544060|T201|COMP|40056-4|LNC|Albumin^6H post XXX challenge|Albumin^6H post XXX challenge
C1544061|T201|COMP|40057-2|LNC|Albumin^6.5H post XXX challenge|Albumin^6.5H post XXX challenge
C1544062|T201|COMP|40058-0|LNC|Albumin^8H post XXX challenge|Albumin^8H post XXX challenge
C1544063|T201|COMP|40059-8|LNC|Albumin^12H post XXX challenge|Albumin^12H post XXX challenge
C1544064|T201|COMP|40060-6|LNC|Albumin^1D post XXX challenge|Albumin^1D post XXX challenge
C1544065|T201|COMP|40061-4|LNC|Albumin^2D post XXX challenge|Albumin^2D post XXX challenge
C1544066|T201|COMP|40062-2|LNC|Albumin^3D post XXX challenge|Albumin^3D post XXX challenge
C1544067|T201|COMP|40063-0|LNC|Albumin^4D post XXX challenge|Albumin^4D post XXX challenge
C1544068|T201|COMP|40064-8|LNC|Calcium^pre XXX challenge|Calcium^pre XXX challenge
C1544069|T201|COMP|40065-5|LNC|Calcium^45M pre XXX challenge|Calcium^45M pre XXX challenge
C1544070|T201|COMP|40066-3|LNC|Calcium^15M pre XXX challenge|Calcium^15M pre XXX challenge
C1544071|T201|COMP|40067-1|LNC|Calcium^baseline|Calcium^baseline
C1544072|T201|COMP|40068-9|LNC|Calcium^45M post XXX challenge|Calcium^45M post XXX challenge
C1544073|T201|COMP|40069-7|LNC|Calcium^1.5H post XXX challenge|Calcium^1.5H post XXX challenge
C1544074|T201|COMP|40070-5|LNC|Calcium^2.5H post XXX challenge|Calcium^2.5H post XXX challenge
C1544075|T201|COMP|40071-3|LNC|Calcium^3H post XXX challenge|Calcium^3H post XXX challenge
C1544076|T201|COMP|40072-1|LNC|Calcium^4H post XXX challenge|Calcium^4H post XXX challenge
C1544077|T201|COMP|40073-9|LNC|Calcium^5H post XXX challenge|Calcium^5H post XXX challenge
C1544078|T201|COMP|40074-7|LNC|Calcium^6H post XXX challenge|Calcium^6H post XXX challenge
C1544079|T201|COMP|40075-4|LNC|Calcium^6.5H post XXX challenge|Calcium^6.5H post XXX challenge
C1544080|T201|COMP|40076-2|LNC|Calcium^7.5H post XXX challenge|Calcium^7.5H post XXX challenge
C1544081|T201|COMP|40077-0|LNC|Calcium^8H post XXX challenge|Calcium^8H post XXX challenge
C1544082|T201|COMP|40078-8|LNC|Calcium^12H post XXX challenge|Calcium^12H post XXX challenge
C1544083|T201|COMP|40079-6|LNC|Calcium^13H post XXX challenge|Calcium^13H post XXX challenge
C1544084|T201|COMP|40080-4|LNC|Calcium^14H post XXX challenge|Calcium^14H post XXX challenge
C1544085|T201|COMP|40081-2|LNC|Calcium^16H post XXX challenge|Calcium^16H post XXX challenge
C1544086|T201|COMP|40082-0|LNC|Calcium^20H post XXX challenge|Calcium^20H post XXX challenge
C1544087|T201|COMP|40083-8|LNC|Calcium^1D post XXX challenge|Calcium^1D post XXX challenge
C1544088|T201|COMP|40084-6|LNC|Calcium^36H post XXX challenge|Calcium^36H post XXX challenge
C1544089|T201|COMP|40085-3|LNC|Calcium^2D post XXX challenge|Calcium^2D post XXX challenge
C1544090|T201|COMP|40086-1|LNC|Calcium^3D post XXX challenge|Calcium^3D post XXX challenge
C1544092|T201|COMP|40088-7|LNC|Coagulation tissue factor induced^baseline|Coagulation tissue factor induced^baseline
C1544103|T201|COMP|40099-4|LNC|Coagulation surface induced^2H pre XXX challenge|Coagulation surface induced^2H pre XXX challenge
C1544104|T201|COMP|40100-0|LNC|Coagulation surface induced^baseline|Coagulation surface induced^baseline
C1544106|T201|COMP|40102-6|LNC|Coagulation surface induced^1H post XXX challenge|Coagulation surface induced^1H post XXX challenge
C1544108|T201|COMP|40104-2|LNC|Coagulation surface induced^2H post XXX challenge|Coagulation surface induced^2H post XXX challenge
C1544109|T201|COMP|40105-9|LNC|Coagulation surface induced^3H post XXX challenge|Coagulation surface induced^3H post XXX challenge
C1544110|T201|COMP|40106-7|LNC|Coagulation surface induced^4H post XXX challenge|Coagulation surface induced^4H post XXX challenge
C1544111|T201|COMP|40107-5|LNC|Coagulation surface induced^6H post XXX challenge|Coagulation surface induced^6H post XXX challenge
C1544112|T201|COMP|40108-3|LNC|Coagulation surface induced^8H post XXX challenge|Coagulation surface induced^8H post XXX challenge
C1544114|T201|COMP|40110-9|LNC|Coagulation surface induced^1D post XXX challenge|Coagulation surface induced^1D post XXX challenge
C1544115|T201|COMP|40120-8|LNC|Creatinine^8H post XXX challenge|Creatinine^8H post XXX challenge
C1544116|T201|COMP|40121-6|LNC|Creatinine^9H post XXX challenge|Creatinine^9H post XXX challenge
C1544117|T201|COMP|40122-4|LNC|Creatinine^10H post XXX challenge|Creatinine^10H post XXX challenge
C1544118|T201|COMP|40123-2|LNC|Creatinine^12H post XXX challenge|Creatinine^12H post XXX challenge
C1544119|T201|COMP|40124-0|LNC|Creatinine^16H post XXX challenge|Creatinine^16H post XXX challenge
C1544120|T201|COMP|40125-7|LNC|Creatinine^18H post XXX challenge|Creatinine^18H post XXX challenge
C1544121|T201|COMP|40126-5|LNC|Creatinine^2D post XXX challenge|Creatinine^2D post XXX challenge
C1544122|T201|COMP|40127-3|LNC|Creatinine^4D post XXX challenge|Creatinine^4D post XXX challenge
C1544123|T201|COMP|40128-1|LNC|Creatinine^7D post XXX challenge|Creatinine^7D post XXX challenge
C1544124|T201|COMP|40129-9|LNC|Creatinine^pre XXX challenge|Creatinine^pre XXX challenge
C1544125|T201|COMP|40130-7|LNC|Creatinine^1.5H pre XXX challenge|Creatinine^1.5H pre XXX challenge
C1544126|T201|COMP|40131-5|LNC|Creatinine^1H pre XXX challenge|Creatinine^1H pre XXX challenge
C1544127|T201|COMP|40132-3|LNC|Creatinine^30M pre XXX challenge|Creatinine^30M pre XXX challenge
C1544128|T201|COMP|40133-1|LNC|Creatinine^baseline|Creatinine^baseline
C1544129|T201|COMP|40134-9|LNC|Creatinine^30M post XXX challenge|Creatinine^30M post XXX challenge
C1544130|T201|COMP|40135-6|LNC|Creatinine^1H post XXX challenge|Creatinine^1H post XXX challenge
C1544131|T201|COMP|40136-4|LNC|Creatinine^1.5H post XXX challenge|Creatinine^1.5H post XXX challenge
C1544132|T201|COMP|40137-2|LNC|Creatinine^2H post XXX challenge|Creatinine^2H post XXX challenge
C1544133|T201|COMP|40138-0|LNC|Creatinine^2.5H post XXX challenge|Creatinine^2.5H post XXX challenge
C1544134|T201|COMP|40139-8|LNC|Creatinine^3H post XXX challenge|Creatinine^3H post XXX challenge
C1544135|T201|COMP|40140-6|LNC|Creatinine^3.5H post XXX challenge|Creatinine^3.5H post XXX challenge
C1544136|T201|COMP|40141-4|LNC|Creatinine^4H post XXX challenge|Creatinine^4H post XXX challenge
C1544137|T201|COMP|40142-2|LNC|Creatinine^4.5H post XXX challenge|Creatinine^4.5H post XXX challenge
C1544138|T201|COMP|40143-0|LNC|Creatinine^5H post XXX challenge|Creatinine^5H post XXX challenge
C1544139|T201|COMP|40144-8|LNC|Creatinine^5.5H post XXX challenge|Creatinine^5.5H post XXX challenge
C1544140|T201|COMP|40145-5|LNC|Creatinine^6H post XXX challenge|Creatinine^6H post XXX challenge
C1544141|T201|COMP|40146-3|LNC|Creatinine^8H post XXX challenge|Creatinine^8H post XXX challenge
C1544142|T201|COMP|40147-1|LNC|Creatinine^1D post XXX challenge|Creatinine^1D post XXX challenge
C1544143|T201|COMP|40148-9|LNC|Glucose^pre XXX challenge|Glucose^pre XXX challenge
C1544144|T201|COMP|40149-7|LNC|Glucose^30M pre XXX challenge|Glucose^30M pre XXX challenge
C1544145|T201|COMP|40150-5|LNC|Glucose^15M pre XXX challenge|Glucose^15M pre XXX challenge
C1544146|T201|COMP|40151-3|LNC|Glucose^10M pre XXX challenge|Glucose^10M pre XXX challenge
C1544147|T201|COMP|40152-1|LNC|Glucose^5M pre XXX challenge|Glucose^5M pre XXX challenge
C1544148|T201|COMP|40153-9|LNC|Glucose^5M post XXX challenge|Glucose^5M post XXX challenge
C1544149|T201|COMP|40154-7|LNC|Glucose^10M post XXX challenge|Glucose^10M post XXX challenge
C1544150|T201|COMP|40155-4|LNC|Glucose^15M post XXX challenge|Glucose^15M post XXX challenge
C1544151|T201|COMP|40156-2|LNC|Glucose^20M post XXX challenge|Glucose^20M post XXX challenge
C1544152|T201|COMP|40157-0|LNC|Glucose^40M post XXX challenge|Glucose^40M post XXX challenge
C1544153|T201|COMP|40158-8|LNC|Glucose^50M post XXX challenge|Glucose^50M post XXX challenge
C1544154|T201|COMP|40159-6|LNC|Glucose^70M post XXX challenge|Glucose^70M post XXX challenge
C1544155|T201|COMP|40160-4|LNC|Glucose^75M post XXX challenge|Glucose^75M post XXX challenge
C1544156|T201|COMP|40161-2|LNC|Glucose^2.5H post XXX challenge|Glucose^2.5H post XXX challenge
C1544157|T201|COMP|40162-0|LNC|Glucose^3H post XXX challenge|Glucose^3H post XXX challenge
C1544158|T201|COMP|40172-9|LNC|Glucose^9.5H post XXX challenge|Glucose^9.5H post XXX challenge
C1544159|T201|COMP|40173-7|LNC|Glucose^10H post XXX challenge|Glucose^10H post XXX challenge
C1544160|T201|COMP|40174-5|LNC|Glucose^10.75H post XXX challenge|Glucose^10.75H post XXX challenge
C1544161|T201|COMP|40175-2|LNC|Glucose^11.5H post XXX challenge|Glucose^11.5H post XXX challenge
C1544162|T201|COMP|40176-0|LNC|Glucose^12H post XXX challenge|Glucose^12H post XXX challenge
C1544163|T201|COMP|40177-8|LNC|Glucose^12.5H post XXX challenge|Glucose^12.5H post XXX challenge
C1544164|T201|COMP|40178-6|LNC|Glucose^13H post XXX challenge|Glucose^13H post XXX challenge
C1544165|T201|COMP|40179-4|LNC|Glucose^13.5H post XXX challenge|Glucose^13.5H post XXX challenge
C1544166|T201|COMP|40180-2|LNC|Glucose^14H post XXX challenge|Glucose^14H post XXX challenge
C1544167|T201|COMP|40181-0|LNC|Glucose^15.5H post XXX challenge|Glucose^15.5H post XXX challenge
C1544168|T201|COMP|40182-8|LNC|Glucose^16H post XXX challenge|Glucose^16H post XXX challenge
C1544169|T201|COMP|40183-6|LNC|Glucose^17.5H post XXX challenge|Glucose^17.5H post XXX challenge
C1544170|T201|COMP|40184-4|LNC|Glucose^18H post XXX challenge|Glucose^18H post XXX challenge
C1544171|T201|COMP|40185-1|LNC|Glucose^18.5H post XXX challenge|Glucose^18.5H post XXX challenge
C1544172|T201|COMP|40186-9|LNC|Glucose^19.5H post XXX challenge|Glucose^19.5H post XXX challenge
C1544173|T201|COMP|40187-7|LNC|Glucose^20H post XXX challenge|Glucose^20H post XXX challenge
C1544174|T201|COMP|40188-5|LNC|Glucose^20.5H post XXX challenge|Glucose^20.5H post XXX challenge
C1544175|T201|COMP|40189-3|LNC|Glucose^21.5H post XXX challenge|Glucose^21.5H post XXX challenge
C1544176|T201|COMP|40190-1|LNC|Glucose^22H post XXX challenge|Glucose^22H post XXX challenge
C1544177|T201|COMP|40191-9|LNC|Glucose^23.5H post XXX challenge|Glucose^23.5H post XXX challenge
C1544178|T201|COMP|40192-7|LNC|Glucose^1D post XXX challenge|Glucose^1D post XXX challenge
C1544179|T201|COMP|40193-5|LNC|Glucose^pre-meal|Glucose^pre-meal
C1544180|T201|COMP|40194-3|LNC|Glucose^20M pre XXX challenge|Glucose^20M pre XXX challenge
C1544181|T201|COMP|40195-0|LNC|Glucose^13M pre XXX challenge|Glucose^13M pre XXX challenge
C1544182|T201|COMP|40196-8|LNC|Glucose^8M pre XXX challenge|Glucose^8M pre XXX challenge
C1544183|T201|COMP|40197-6|LNC|Glucose^3M pre XXX challenge|Glucose^3M pre XXX challenge
C1544184|T201|COMP|40198-4|LNC|Glucose^2M post XXX challenge|Glucose^2M post XXX challenge
C1544185|T201|COMP|40199-2|LNC|Glucose^3M post XXX challenge|Glucose^3M post XXX challenge
C1544186|T201|COMP|40200-8|LNC|Glucose^4M post XXX challenge|Glucose^4M post XXX challenge
C1544187|T201|COMP|40201-6|LNC|Glucose^6M post XXX challenge|Glucose^6M post XXX challenge
C1544188|T201|COMP|40211-5|LNC|Glucose^3.5H post XXX challenge|Glucose^3.5H post XXX challenge
C1544189|T201|COMP|40212-3|LNC|Glucose^4.5H post XXX challenge|Glucose^4.5H post XXX challenge
C1544190|T201|COMP|40213-1|LNC|Glucose^5.5H post XXX challenge|Glucose^5.5H post XXX challenge
C1544191|T201|COMP|40214-9|LNC|Glucose^25H post XXX challenge|Glucose^25H post XXX challenge
C1544192|T201|COMP|40215-6|LNC|Glucose^26H post XXX challenge|Glucose^26H post XXX challenge
C1544193|T201|COMP|40216-4|LNC|Glucose^27H post XXX challenge|Glucose^27H post XXX challenge
C1544194|T201|COMP|40217-2|LNC|Glucose^28H post XXX challenge|Glucose^28H post XXX challenge
C1544195|T201|COMP|40218-0|LNC|Glucose^29H post XXX challenge|Glucose^29H post XXX challenge
C1544196|T201|COMP|40219-8|LNC|Glucose^30H post XXX challenge|Glucose^30H post XXX challenge
C1544197|T201|COMP|40220-6|LNC|Glucose^31H post XXX challenge|Glucose^31H post XXX challenge
C1544198|T201|COMP|40221-4|LNC|Glucose^36H post XXX challenge|Glucose^36H post XXX challenge
C1544199|T201|COMP|40222-2|LNC|Glucose^2D post XXX challenge|Glucose^2D post XXX challenge
C1544200|T201|COMP|40223-0|LNC|Calcium^pre XXX challenge|Calcium^pre XXX challenge
C1544201|T201|COMP|40224-8|LNC|Calcium^45M pre XXX challenge|Calcium^45M pre XXX challenge
C1544202|T201|COMP|40225-5|LNC|Calcium^15M pre XXX challenge|Calcium^15M pre XXX challenge
C1544203|T201|COMP|40226-3|LNC|Calcium^baseline|Calcium^baseline
C1544204|T201|COMP|40227-1|LNC|Calcium^30M post XXX challenge|Calcium^30M post XXX challenge
C1544205|T201|COMP|40228-9|LNC|Calcium^45M post XXX challenge|Calcium^45M post XXX challenge
C1544206|T201|COMP|40229-7|LNC|Calcium^1H post XXX challenge|Calcium^1H post XXX challenge
C1544207|T201|COMP|40230-5|LNC|Calcium^1.5H post XXX challenge|Calcium^1.5H post XXX challenge
C1544208|T201|COMP|40231-3|LNC|Calcium^2H post XXX challenge|Calcium^2H post XXX challenge
C1544209|T201|COMP|40232-1|LNC|Calcium^2.5H post XXX challenge|Calcium^2.5H post XXX challenge
C1544210|T201|COMP|40233-9|LNC|Calcium^3H post XXX challenge|Calcium^3H post XXX challenge
C1544211|T201|COMP|40234-7|LNC|Calcium^4H post XXX challenge|Calcium^4H post XXX challenge
C1544212|T201|COMP|40235-4|LNC|Calcium^5H post XXX challenge|Calcium^5H post XXX challenge
C1544213|T201|COMP|40236-2|LNC|Calcium^6.5H post XXX challenge|Calcium^6.5H post XXX challenge
C1544214|T201|COMP|40237-0|LNC|Calcium^7.5H post XXX challenge|Calcium^7.5H post XXX challenge
C1544215|T201|COMP|40238-8|LNC|Calcium^8H post XXX challenge|Calcium^8H post XXX challenge
C1544216|T201|COMP|40239-6|LNC|Calcium^12H post XXX challenge|Calcium^12H post XXX challenge
C1544217|T201|COMP|40240-4|LNC|Calcium^13H post XXX challenge|Calcium^13H post XXX challenge
C1544218|T201|COMP|40241-2|LNC|Calcium^14H post XXX challenge|Calcium^14H post XXX challenge
C1544219|T201|COMP|40242-0|LNC|Calcium^16H post XXX challenge|Calcium^16H post XXX challenge
C1544220|T201|COMP|40243-8|LNC|Calcium^20H post XXX challenge|Calcium^20H post XXX challenge
C1544221|T201|COMP|40244-6|LNC|Calcium^1D post XXX challenge|Calcium^1D post XXX challenge
C1544222|T201|COMP|40245-3|LNC|Calcium^36H post XXX challenge|Calcium^36H post XXX challenge
C1544223|T201|COMP|40246-1|LNC|Calcium^2D post XXX challenge|Calcium^2D post XXX challenge
C1544224|T201|COMP|40247-9|LNC|Calcium^3D post XXX challenge|Calcium^3D post XXX challenge
C1544225|T201|COMP|40248-7|LNC|Creatinine^baseline|Creatinine^baseline
C1544226|T201|COMP|40249-5|LNC|Creatinine^30M post XXX challenge|Creatinine^30M post XXX challenge
C1544227|T201|COMP|40250-3|LNC|Creatinine^1H post XXX challenge|Creatinine^1H post XXX challenge
C1544228|T201|COMP|40251-1|LNC|Creatinine^1.5H post XXX challenge|Creatinine^1.5H post XXX challenge
C1544229|T201|COMP|40252-9|LNC|Creatinine^2H post XXX challenge|Creatinine^2H post XXX challenge
C1544230|T201|COMP|40254-5|LNC|Creatinine^2.5H post XXX challenge|Creatinine^2.5H post XXX challenge
C1544231|T201|COMP|40255-2|LNC|Creatinine^3H post XXX challenge|Creatinine^3H post XXX challenge
C1544232|T201|COMP|40256-0|LNC|Creatinine^5H post XXX challenge|Creatinine^5H post XXX challenge
C1544233|T201|COMP|40257-8|LNC|Creatinine^6H post XXX challenge|Creatinine^6H post XXX challenge
C1544234|T201|COMP|40258-6|LNC|Creatinine^1D post XXX challenge|Creatinine^1D post XXX challenge
C1544235|T201|COMP|40259-4|LNC|Glucose^10.5H post XXX challenge|Glucose^10.5H post XXX challenge
C1544236|T201|COMP|40260-2|LNC|Glucose^10.75H post XXX challenge|Glucose^10.75H post XXX challenge
C1544237|T201|COMP|40261-0|LNC|Glucose^13M pre XXX challenge|Glucose^13M pre XXX challenge
C1544238|T201|COMP|40262-8|LNC|Glucose^3M pre XXX challenge|Glucose^3M pre XXX challenge
C1544239|T201|COMP|40263-6|LNC|Glucose^30M post XXX challenge|Glucose^30M post XXX challenge
C1544240|T201|COMP|40264-4|LNC|Creatinine^baseline|Creatinine^baseline
C1544241|T201|COMP|40265-1|LNC|Creatinine^30M post XXX challenge|Creatinine^30M post XXX challenge
C1544242|T201|COMP|40266-9|LNC|Creatinine^1H post XXX challenge|Creatinine^1H post XXX challenge
C1544243|T201|COMP|40267-7|LNC|Creatinine^1.5H post XXX challenge|Creatinine^1.5H post XXX challenge
C1544244|T201|COMP|40268-5|LNC|Creatinine^2H post XXX challenge|Creatinine^2H post XXX challenge
C1544245|T201|COMP|40269-3|LNC|Creatinine^2.5H post XXX challenge|Creatinine^2.5H post XXX challenge
C1544246|T201|COMP|40270-1|LNC|Creatinine^3H post XXX challenge|Creatinine^3H post XXX challenge
C1544247|T201|COMP|40271-9|LNC|Creatinine^5H post XXX challenge|Creatinine^5H post XXX challenge
C1544248|T201|COMP|40272-7|LNC|Creatinine^6H post XXX challenge|Creatinine^6H post XXX challenge
C1544249|T201|COMP|40273-5|LNC|Creatinine^1D post XXX challenge|Creatinine^1D post XXX challenge
C1544250|T201|COMP|40274-3|LNC|Cortisol^15M post XXX challenge|Cortisol^15M post XXX challenge
C1544251|T201|COMP|40275-0|LNC|Cortisol^45M post XXX challenge|Cortisol^45M post XXX challenge
C1544252|T201|COMP|40276-8|LNC|Glucose^30M post dose lactose PO|Glucose^30M post dose lactose PO
C1544253|T201|COMP|40277-6|LNC|Glucose^1H post dose lactose PO|Glucose^1H post dose lactose PO
C1544254|T201|COMP|40278-4|LNC|Glucose^1.5H post dose lactose PO|Glucose^1.5H post dose lactose PO
C1544255|T201|COMP|40279-2|LNC|Glucose^2H post dose lactose PO|Glucose^2H post dose lactose PO
C1544256|T201|COMP|40280-0|LNC|Glucose^3H post dose lactose PO|Glucose^3H post dose lactose PO
C1544257|T201|COMP|40281-8|LNC|Lactose^30M post dose lactose PO|Lactose^30M post dose lactose PO
C1544258|T201|COMP|40282-6|LNC|Lactose^1H post dose lactose PO|Lactose^1H post dose lactose PO
C1544259|T201|COMP|40283-4|LNC|Lactose^1.5H post dose lactose PO|Lactose^1.5H post dose lactose PO
C1544260|T201|COMP|40284-2|LNC|Lactose^2H post dose lactose PO|Lactose^2H post dose lactose PO
C1544261|T201|COMP|40285-9|LNC|Glucose^75M post dose glucose|Glucose^75M post dose glucose
C1544262|T201|COMP|40286-7|LNC|Glucose^105M post dose glucose|Glucose^105M post dose glucose
C1544263|T201|COMP|40287-5|LNC|Glucose^1H post meal|Glucose^1H post meal
C1544264|T201|COMP|40288-3|LNC|Insulin^30M post XXX challenge|Insulin^30M post XXX challenge
C1544265|T201|COMP|40289-1|LNC|Insulin^1H post XXX challenge|Insulin^1H post XXX challenge
C1544266|T201|COMP|40290-9|LNC|Insulin^1.5H post XXX challenge|Insulin^1.5H post XXX challenge
C1544267|T201|COMP|40291-7|LNC|Insulin^2H post XXX challenge|Insulin^2H post XXX challenge
C1544268|T201|COMP|40292-5|LNC|Insulin^2.5H post XXX challenge|Insulin^2.5H post XXX challenge
C1544269|T201|COMP|40293-3|LNC|Insulin^3H post XXX challenge|Insulin^3H post XXX challenge
C1544270|T201|COMP|40295-8|LNC|Triiodothyronine.free^2H post XXX challenge|Triiodothyronine.free^2H post XXX challenge
C1544271|T201|COMP|40296-6|LNC|Xylose^post CFst|Xylose^post CFst
C1544272|T201|COMP|40297-4|LNC|Somatotropin^3.5H post XXX challenge|Somatotropin^3.5H post XXX challenge
C1544273|T201|COMP|40298-2|LNC|Somatotropin^pre dose cloNIDine|Somatotropin^pre dose cloNIDine
C1544274|T201|COMP|40299-0|LNC|Somatotropin^1H post dose cloNIDine|Somatotropin^1H post dose cloNIDine
C1544275|T201|COMP|40300-6|LNC|Somatotropin^1.5H post dose cloNIDine|Somatotropin^1.5H post dose cloNIDine
C1544276|T201|COMP|40301-4|LNC|Somatotropin^2H post dose cloNIDine|Somatotropin^2H post dose cloNIDine
C1544277|T201|COMP|40302-2|LNC|Somatotropin^pre dose arginine|Somatotropin^pre dose arginine
C1544278|T201|COMP|40303-0|LNC|Somatotropin^1H post dose arginine|Somatotropin^1H post dose arginine
C1544279|T201|COMP|40304-8|LNC|Somatotropin^1.5H post dose arginine|Somatotropin^1.5H post dose arginine
C1544280|T201|COMP|40305-5|LNC|Somatotropin^2H post dose arginine|Somatotropin^2H post dose arginine
C1544281|T201|COMP|40306-3|LNC|Somatotropin^3H post dose arginine|Somatotropin^3H post dose arginine
C1544282|T201|COMP|40307-1|LNC|Somatotropin^3.5H post dose arginine|Somatotropin^3.5H post dose arginine
C1544283|T201|COMP|40308-9|LNC|Somatotropin^4H post dose arginine|Somatotropin^4H post dose arginine
C1544284|T201|COMP|40309-7|LNC|Somatotropin^pre or post dose glucose|Somatotropin^pre or post dose glucose
C1544285|T201|COMP|40310-5|LNC|Cortisol^pre dose triple bolus|Cortisol^pre dose triple bolus
C1544286|T201|COMP|40311-3|LNC|Cortisol^15M post dose triple bolus|Cortisol^15M post dose triple bolus
C1544287|T201|COMP|40312-1|LNC|Cortisol^30M post dose triple bolus|Cortisol^30M post dose triple bolus
C1544288|T201|COMP|40313-9|LNC|Cortisol^45M post dose triple bolus|Cortisol^45M post dose triple bolus
C1544289|T201|COMP|40314-7|LNC|Cortisol^1H post dose triple bolus|Cortisol^1H post dose triple bolus
C1544290|T201|COMP|40315-4|LNC|Cortisol^1.5H post dose triple bolus|Cortisol^1.5H post dose triple bolus
C1544291|T201|COMP|40316-2|LNC|Cortisol^2H post dose triple bolus|Cortisol^2H post dose triple bolus
C1544292|T201|COMP|40317-0|LNC|Cortisol^3H post dose triple bolus|Cortisol^3H post dose triple bolus
C1544293|T201|COMP|40318-8|LNC|Glucose^pre dose triple bolus|Glucose^pre dose triple bolus
C1544294|T201|COMP|40319-6|LNC|Glucose^15M post dose triple bolus|Glucose^15M post dose triple bolus
C1544295|T201|COMP|40320-4|LNC|Glucose^30M post dose triple bolus|Glucose^30M post dose triple bolus
C1544296|T201|COMP|40321-2|LNC|Glucose^45M post dose triple bolus|Glucose^45M post dose triple bolus
C1544297|T201|COMP|40322-0|LNC|Glucose^1H post dose triple bolus|Glucose^1H post dose triple bolus
C1544298|T201|COMP|40323-8|LNC|Glucose^2H post dose triple bolus|Glucose^2H post dose triple bolus
C1544299|T201|COMP|40324-6|LNC|Glucose^3H post dose triple bolus|Glucose^3H post dose triple bolus
C1544300|T201|COMP|40325-3|LNC|Testosterone^pre dose triple bolus|Testosterone^pre dose triple bolus
C1544301|T201|COMP|40326-1|LNC|Testosterone^3H post dose triple bolus|Testosterone^3H post dose triple bolus
C1544302|T201|COMP|40327-9|LNC|Triiodothyronine.free^pre dose triple bolus|Triiodothyronine.free^pre dose triple bolus
C1544303|T201|COMP|40328-7|LNC|Triiodothyronine.free^2H post dose triple bolus|Triiodothyronine.free^2H post dose triple bolus
C1544304|T201|COMP|40329-5|LNC|Prolactin^pre dose triple bolus|Prolactin^pre dose triple bolus
C1544305|T201|COMP|40330-3|LNC|Prolactin^15M post dose triple bolus|Prolactin^15M post dose triple bolus
C1544306|T201|COMP|40331-1|LNC|Prolactin^20M post dose triple bolus|Prolactin^20M post dose triple bolus
C1544307|T201|COMP|40332-9|LNC|Prolactin^30M post dose triple bolus|Prolactin^30M post dose triple bolus
C1544308|T201|COMP|40333-7|LNC|Prolactin^1H post dose triple bolus|Prolactin^1H post dose triple bolus
C1544309|T201|COMP|40334-5|LNC|Somatotropin^pre dose triple bolus|Somatotropin^pre dose triple bolus
C1544310|T201|COMP|40335-2|LNC|Somatotropin^15M post dose triple bolus|Somatotropin^15M post dose triple bolus
C1544311|T201|COMP|40336-0|LNC|Somatotropin^30M post dose triple bolus|Somatotropin^30M post dose triple bolus
C1544312|T201|COMP|40337-8|LNC|Somatotropin^45M post dose triple bolus|Somatotropin^45M post dose triple bolus
C1544313|T201|COMP|40338-6|LNC|Somatotropin^1H post dose triple bolus|Somatotropin^1H post dose triple bolus
C1544314|T201|COMP|40339-4|LNC|Somatotropin^2H post dose triple bolus|Somatotropin^2H post dose triple bolus
C1544315|T201|COMP|40340-2|LNC|Somatotropin^3H post dose triple bolus|Somatotropin^3H post dose triple bolus
C1544316|T201|COMP|40341-0|LNC|MT-ATP6 gene.m.8993T>G|MT-ATP6 gene.m.8993T>G
C1544317|T201|COMP|40342-8|LNC|MT-TL1 gene.m.3271T>C|MT-TL1 gene.m.3271T>C
C1544318|T201|COMP|40343-6|LNC|MT-TK gene.m.8296A>G|MT-TK gene.m.8296A>G
C1544319|T201|COMP|40344-4|LNC|Mttl1 gene.c.A3243G|Mttl1 gene.c.A3243G
C1544320|T201|COMP|40345-1|LNC|MT-TK gene.m.8356T>C|MT-TK gene.m.8356T>C
C1544321|T201|COMP|40346-9|LNC|MT-CO1 gene.m.7445A>G|MT-CO1 gene.m.7445A>G
C1544322|T201|COMP|40347-7|LNC|MT-TL1 gene.m.3256C>T|MT-TL1 gene.m.3256C>T
C1544323|T201|COMP|40348-5|LNC|MT-TL1 gene.m.3252T>C|MT-TL1 gene.m.3252T>C
C1544324|T201|COMP|40349-3|LNC|MT-TK gene.m.8363G>A|MT-TK gene.m.8363G>A
C1544325|T201|COMP|40350-1|LNC|MT-TL1 gene.m.3291T>C|MT-TL1 gene.m.3291T>C
C1544326|T201|COMP|40351-9|LNC|MT-ND4 gene.m.11778G>A|MT-ND4 gene.m.11778G>A
C1544327|T201|COMP|40352-7|LNC|MT-ND5 gene.m.13513G>A|MT-ND5 gene.m.13513G>A
C1544328|T201|COMP|40353-5|LNC|MT-ND6 gene.m.14484T>C|MT-ND6 gene.m.14484T>C
C1544329|T201|COMP|40354-3|LNC|MT-ND1 gene.m.3460G>A|MT-ND1 gene.m.3460G>A
C1544330|T201|COMP|40355-0|LNC|Cotinine|Cotinine
C1544331|T201|COMP|40356-8|LNC|Creatinine|Creatinine
C1544332|T201|COMP|40357-6|LNC|Creatinine|Creatinine
C1544333|T201|COMP|40358-4|LNC|Desipramine|Desipramine
C1544334|T201|COMP|40359-2|LNC|Dextromethorphan|Dextromethorphan
C1544335|T201|COMP|40360-0|LNC|Follitropin^15M post dose triple bolus|Follitropin^15M post dose triple bolus
C1544336|T201|COMP|40361-8|LNC|Follitropin^1H post dose triple bolus|Follitropin^1H post dose triple bolus
C1544337|T201|COMP|40362-6|LNC|Follitropin^20M post dose triple bolus|Follitropin^20M post dose triple bolus
C1544338|T201|COMP|40363-4|LNC|Follitropin^2H post dose triple bolus|Follitropin^2H post dose triple bolus
C1544339|T201|COMP|40364-2|LNC|Follitropin^30M post dose triple bolus|Follitropin^30M post dose triple bolus
C1544340|T201|COMP|40365-9|LNC|Follitropin^pre dose triple bolus|Follitropin^pre dose triple bolus
C1544341|T201|COMP|40366-7|LNC|Glucose|Glucose
C1544342|T201|COMP|40367-5|LNC|Heptacarboxylate|Heptacarboxylate
C1544343|T201|COMP|40368-3|LNC|Hexacarboxylate|Hexacarboxylate
C1544344|T201|COMP|40369-1|LNC|HYDROmorphone|HYDROmorphone
C1544345|T201|COMP|40370-9|LNC|Imipramine|Imipramine
C1544346|T201|COMP|40371-7|LNC|Isoniazid|Isoniazid
C1544347|T201|COMP|40372-5|LNC|Isopropanol|Isopropanol
C1544348|T201|COMP|40373-3|LNC|Lutropin^15M post dose triple bolus|Lutropin^15M post dose triple bolus
C1544349|T201|COMP|40374-1|LNC|Lutropin^1H post dose triple bolus|Lutropin^1H post dose triple bolus
C1544350|T201|COMP|40375-8|LNC|Lutropin^20M post dose triple bolus|Lutropin^20M post dose triple bolus
C1544351|T201|COMP|40376-6|LNC|Lutropin^2H post dose triple bolus|Lutropin^2H post dose triple bolus
C1544352|T201|COMP|40377-4|LNC|Lutropin^30M post dose triple bolus|Lutropin^30M post dose triple bolus
C1544353|T201|COMP|40378-2|LNC|Lutropin^pre dose triple bolus|Lutropin^pre dose triple bolus
C1544354|T201|COMP|40379-0|LNC|Maprotiline|Maprotiline
C1544355|T201|COMP|40380-8|LNC|Meprobamate|Meprobamate
C1544356|T201|COMP|40381-6|LNC|Methamphetamine|Methamphetamine
C1544357|T201|COMP|40382-4|LNC|Methaqualone|Methaqualone
C1544358|T201|COMP|40383-2|LNC|Methyprylon|Methyprylon
C1544359|T201|COMP|40384-0|LNC|Morphine|Morphine
C1544360|T201|COMP|40385-7|LNC|Nicotine|Nicotine
C1544361|T201|COMP|40386-5|LNC|Nicotine|Nicotine
C1544362|T201|COMP|40387-3|LNC|Nicotine|Nicotine
C1544363|T201|COMP|40388-1|LNC|Nitrogen|Nitrogen
C1544364|T201|COMP|40389-9|LNC|Nortriptyline|Nortriptyline
C1544365|T201|COMP|40390-7|LNC|OLANZapine|OLANZapine
C1544366|T201|COMP|40391-5|LNC|Para aminobenzoate.free|Para aminobenzoate.free
C1544367|T201|COMP|40392-3|LNC|Pentacarboxylate|Pentacarboxylate
C1544368|T201|COMP|40393-1|LNC|Pentazocine|Pentazocine
C1544369|T201|COMP|40394-9|LNC|Phencyclidine|Phencyclidine
C1544370|T201|COMP|40395-6|LNC|Phentermine|Phentermine
C1544371|T201|COMP|40396-4|LNC|Porphyrins|Porphyrins
C1544372|T201|COMP|40397-2|LNC|Thyrotropin^15M post dose triple bolus|Thyrotropin^15M post dose triple bolus
C1544373|T201|COMP|40398-0|LNC|Thyrotropin^1H post dose triple bolus|Thyrotropin^1H post dose triple bolus
C1544374|T201|COMP|40399-8|LNC|Thyrotropin^20M post dose triple bolus|Thyrotropin^20M post dose triple bolus
C1544375|T201|COMP|40400-4|LNC|Thyrotropin^30M post dose triple bolus|Thyrotropin^30M post dose triple bolus
C1544376|T201|COMP|40401-2|LNC|Thyrotropin^pre dose triple bolus|Thyrotropin^pre dose triple bolus
C1544377|T201|COMP|40402-0|LNC|traZODone|traZODone
C1544378|T201|COMP|40403-8|LNC|Trimipramine|Trimipramine
C1544379|T201|COMP|40404-6|LNC|Tripelennamine|Tripelennamine
C1544380|T201|COMP|40405-3|LNC|Urea|Urea
C1544381|T201|COMP|40406-1|LNC|Urea|Urea
C1544382|T201|COMP|40407-9|LNC|Uroporphyrin 1 isomer|Uroporphyrin 1 isomer
C1544383|T201|COMP|40408-7|LNC|Uroporphyrin 3 isomer|Uroporphyrin 3 isomer
C1544384|T201|COMP|40409-5|LNC|3-Methoxytyramine|3-Methoxytyramine
C1544385|T201|COMP|40410-3|LNC|Alkaline phosphatase|Alkaline phosphatase
C1544386|T201|COMP|40411-1|LNC|Amitriptyline|Amitriptyline
C1544387|T201|COMP|40412-9|LNC|Barbiturates|Barbiturates
C1544388|T201|COMP|40413-7|LNC|Barbiturates|Barbiturates
C1544389|T201|COMP|40414-5|LNC|Benzodiazepines|Benzodiazepines
C1544390|T201|COMP|40415-2|LNC|Benzodiazepines|Benzodiazepines
C1544391|T201|COMP|40416-0|LNC|Caffeine|Caffeine
C1544392|T201|COMP|40417-8|LNC|Chromium|Chromium
C1544393|T201|COMP|40418-6|LNC|Cotinine|Cotinine
C1544394|T201|COMP|40419-4|LNC|Amphetamine+Methamphetamine|Amphetamine+Methamphetamine
C1544395|T201|COMP|40420-2|LNC|Amphetamine+Methamphetamine|Amphetamine+Methamphetamine
C1544396|T201|COMP|40421-0|LNC|Amphetamine+Methamphetamine|Amphetamine+Methamphetamine
C1544397|T201|COMP|40422-8|LNC|Methotrimeprazine|Methotrimeprazine
C1544398|T201|COMP|40423-6|LNC|Methotrimeprazine|Methotrimeprazine
C1544399|T201|COMP|40424-4|LNC|Methotrimeprazine|Methotrimeprazine
C1544400|T201|COMP|40425-1|LNC|CYP2D6 gene targeted mutation analysis|CYP2D6 gene targeted mutation analysis
C1544401|T201|COMP|40426-9|LNC|FGD1 gene targeted mutation analysis|FGD1 gene targeted mutation analysis
C1544402|T201|COMP|40427-7|LNC|FGF23 gene targeted mutation analysis|FGF23 gene targeted mutation analysis
C1544403|T201|COMP|40428-5|LNC|NIPBL gene targeted mutation analysis|NIPBL gene targeted mutation analysis
C1544404|T201|COMP|40429-3|LNC|NOD2 gene targeted mutation analysis|NOD2 gene targeted mutation analysis
C1544405|T201|COMP|40430-1|LNC|TH gene targeted mutation analysis|TH gene targeted mutation analysis
C1544406|T201|COMP|40431-9|LNC|Osmotic fragility^fresh|Osmotic fragility^fresh
C1544407|T201|COMP|40432-7|LNC|Osmotic fragility^incubated|Osmotic fragility^incubated
C1544408|T201|COMP|40433-5|LNC|Sucrose hemolysis|Sucrose hemolysis
C1544409|T201|COMP|40434-3|LNC|APTX gene targeted mutation analysis|APTX gene targeted mutation analysis
C1544410|T201|COMP|40435-0|LNC|Fungus identified|Fungus identified
C1544411|T201|COMP|40436-8|LNC|Parainfluenza virus identified|Parainfluenza virus identified
C1544412|T201|COMP|40437-6|LNC|HIV 1 p24 Ab|HIV 1 p24 Ab
C1544413|T201|COMP|40438-4|LNC|HIV 1 gp41 Ab|HIV 1 gp41 Ab
C1544414|T201|COMP|40439-2|LNC|HIV 1 gp120+gp160 Ab|HIV 1 gp120+gp160 Ab
C1544415|T201|COMP|40440-0|LNC|XXX microorganism serotype|XXX microorganism serotype
C1544419|T201|COMP|40444-2|LNC|Cytomegalovirus gene mutations detected|Cytomegalovirus gene mutations detected
C1544426|T201|COMP|40451-7|LNC|Lead|Lead
C1544427|T201|COMP|40452-5|LNC|Sialate/Creatinine|Sialate/Creatinine
C1544428|T201|COMP|40453-3|LNC|Sialooligosaccharides|Sialooligosaccharides
C1544429|T201|COMP|40454-1|LNC|Coagulum lysis|Coagulum lysis
C1544430|T201|COMP|40455-8|LNC|Ceruloplasmin actual/Normal|Ceruloplasmin actual/Normal
C1544431|T201|COMP|40456-6|LNC|Beta 2 glycoprotein 1 Ab|Beta 2 glycoprotein 1 Ab
C1544432|T201|COMP|40457-4|LNC|Prothrombin Ab|Prothrombin Ab
C1544434|T201|COMP|40459-0|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1544435|T201|COMP|40460-8|LNC|Phenytoin.bound|Phenytoin.bound
C1544436|T201|COMP|40461-6|LNC|GJB1 gene allele 1|GJB1 gene allele 1
C1544437|T201|COMP|40462-4|LNC|GJB1 gene allele 2|GJB1 gene allele 2
C1544438|T201|COMP|40463-2|LNC|TNFRSF1A gene targeted mutation analysis|TNFRSF1A gene targeted mutation analysis
C1544439|T201|COMP|40464-0|LNC|Drugs identified|Drugs identified
C1544440|T201|COMP|40465-7|LNC|Glimepiride|Glimepiride
C1544441|T201|COMP|40466-5|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C1544442|T201|COMP|40467-3|LNC|U1 small nuclear ribonucleoprotein Ab.IgG|U1 small nuclear ribonucleoprotein Ab.IgG
C1544443|T201|COMP|40468-1|LNC|SLC26A4 gene targeted mutation analysis|SLC26A4 gene targeted mutation analysis
C1544444|T201|COMP|40469-9|LNC|Hydroflumethiazide|Hydroflumethiazide
C1544445|T201|COMP|40470-7|LNC|Lymphocytes|Lymphocytes
C1544446|T201|COMP|40471-5|LNC|FBN1 gene targeted mutation analysis|FBN1 gene targeted mutation analysis
C1544447|T201|COMP|40472-3|LNC|Tetradecadienoate/Creatinine|Tetradecadienoate/Creatinine
C1544448|T201|COMP|40473-1|LNC|Thermoactinomyces vulgaris 1 Ab|Thermoactinomyces vulgaris 1 Ab
C1544449|T201|COMP|40474-9|LNC|Volatiles|Volatiles
C1544450|T201|COMP|40475-6|LNC|WFS1 gene targeted mutation analysis|WFS1 gene targeted mutation analysis
C1544451|T201|COMP|40476-4|LNC|PARK2 gene targeted mutation analysis|PARK2 gene targeted mutation analysis
C1544452|T201|COMP|40477-2|LNC|L1CAM gene targeted mutation analysis|L1CAM gene targeted mutation analysis
C1544453|T201|COMP|40478-0|LNC|MAPT gene targeted mutation analysis|MAPT gene targeted mutation analysis
C1544454|T201|COMP|40479-8|LNC|Virus identified|Virus identified
C1544455|T201|COMP|40480-6|LNC|Virus identified|Virus identified
C1544456|T201|COMP|40481-4|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C1544457|T201|COMP|40482-2|LNC|Crystals.unidentified|Crystals.unidentified
C1544458|T201|COMP|40483-0|LNC|Phosphate crystals.amorphous|Phosphate crystals.amorphous
C1544459|T201|COMP|40484-8|LNC|Urate crystals.amorphous|Urate crystals.amorphous
C1544460|T201|COMP|40485-5|LNC|Urate crystals|Urate crystals
C1544461|T201|COMP|40486-3|LNC|Protein/Creatinine|Protein/Creatinine
C1544462|T201|COMP|40487-1|LNC|Urea/Creatinine|Urea/Creatinine
C1544463|T201|COMP|40488-9|LNC|Glucose/Creatinine|Glucose/Creatinine
C1544464|T201|COMP|40489-7|LNC|Histiocytes/100 cells|Histiocytes/100 cells
C1544465|T201|COMP|40490-5|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C1544466|T201|COMP|40492-1|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C1544467|T201|COMP|40493-9|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C1544468|T201|COMP|40494-7|LNC|Yersinia pseudotuberculosis Ab|Yersinia pseudotuberculosis Ab
C1544469|T201|COMP|40495-4|LNC|Yersinia pseudotuberculosis 3 Ab|Yersinia pseudotuberculosis 3 Ab
C1544470|T201|COMP|40496-2|LNC|Yersinia pseudotuberculosis 2 Ab|Yersinia pseudotuberculosis 2 Ab
C1544471|T201|COMP|40497-0|LNC|Yersinia pseudotuberculosis 1 Ab|Yersinia pseudotuberculosis 1 Ab
C1544472|T201|COMP|40498-8|LNC|Yersinia enterocolitica Ab|Yersinia enterocolitica Ab
C1544473|T201|COMP|40499-6|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C1544474|T201|COMP|40500-1|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C1544475|T201|COMP|40501-9|LNC|Candida sp Ab|Candida sp Ab
C1544476|T201|COMP|40502-7|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C1544477|T201|COMP|40503-5|LNC|Sindbis virus Ab|Sindbis virus Ab
C1544478|T201|COMP|40504-3|LNC|Powassan virus Ab|Powassan virus Ab
C1544479|T201|COMP|40505-0|LNC|Chikungunya virus Ab|Chikungunya virus Ab
C1544480|T201|COMP|40506-8|LNC|Jamestown canyon virus Ab|Jamestown canyon virus Ab
C1544481|T201|COMP|40507-6|LNC|Jamestown canyon virus Ab|Jamestown canyon virus Ab
C1544482|T201|COMP|40508-4|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1544483|T201|COMP|40509-2|LNC|Snowshoe hare virus Ab.IgM|Snowshoe hare virus Ab.IgM
C1544484|T201|COMP|40510-0|LNC|Snowshoe hare virus Ab|Snowshoe hare virus Ab
C1544485|T201|COMP|40511-8|LNC|Snowshoe hare virus Ab|Snowshoe hare virus Ab
C1544486|T201|COMP|40512-6|LNC|Semliki forest virus Ab|Semliki forest virus Ab
C1544487|T201|COMP|40513-4|LNC|Powassan virus Ab|Powassan virus Ab
C1544488|T201|COMP|40514-2|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C1544489|T201|COMP|40515-9|LNC|Dengue virus Ab|Dengue virus Ab
C1544490|T201|COMP|40516-7|LNC|Histiocytes/100 cells|Histiocytes/100 cells
C1544491|T201|COMP|40517-5|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C1544492|T201|COMP|40518-3|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C1544493|T201|COMP|40519-1|LNC|Histiocytes/100 cells|Histiocytes/100 cells
C1544494|T201|COMP|40520-9|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C1544495|T201|COMP|40521-7|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C1544496|T201|COMP|40522-5|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C1544497|T201|COMP|40523-3|LNC|Histiocytes/100 cells|Histiocytes/100 cells
C1544498|T201|COMP|40534-0|LNC|Erythrocytes|Erythrocytes
C1544499|T201|COMP|40535-7|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C1544500|T201|COMP|40536-5|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C1544501|T201|COMP|40537-3|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C1544502|T201|COMP|40538-1|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C1544503|T201|COMP|40539-9|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1544504|T201|COMP|40540-7|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1544505|T201|COMP|40541-5|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C1544506|T201|COMP|40542-3|LNC|Rubella virus Ab|Rubella virus Ab
C1544507|T201|COMP|40543-1|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C1544508|T201|COMP|40544-9|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C1544509|T201|COMP|40545-6|LNC|Hemoglobin C|Hemoglobin C
C1544510|T201|COMP|40546-4|LNC|Hemoglobin E|Hemoglobin E
C1544511|T201|COMP|40547-2|LNC|Hemoglobin H|Hemoglobin H
C1544512|T201|COMP|40548-0|LNC|Mononuclear cells.atypical|Mononuclear cells.atypical
C1544513|T201|COMP|40549-8|LNC|Hemoglobin F|Hemoglobin F
C1544514|T201|COMP|40550-6|LNC|Hemoglobin H|Hemoglobin H
C1544515|T201|COMP|40551-4|LNC|CD10 Ag|CD10 Ag
C1544516|T201|COMP|40552-2|LNC|CD117 Ag|CD117 Ag
C1544517|T201|COMP|40553-0|LNC|CD19 Ag|CD19 Ag
C1544518|T201|COMP|40554-8|LNC|CD45 Ag|CD45 Ag
C1544519|T201|COMP|40555-5|LNC|CD66e Ag|CD66e Ag
C1544520|T201|COMP|40556-3|LNC|Estrogen receptor Ag|Estrogen receptor Ag
C1544521|T201|COMP|40557-1|LNC|Progesterone receptor Ag|Progesterone receptor Ag
C1544522|T201|COMP|40558-9|LNC|Cytokeratin 20 Ag|Cytokeratin 20 Ag
C1544523|T201|COMP|40559-7|LNC|Cytokeratin 7 Ag|Cytokeratin 7 Ag
C1544524|T201|COMP|40560-5|LNC|Cytokeratin AE1+AE3 Ag|Cytokeratin AE1+AE3 Ag
C1544525|T201|COMP|40561-3|LNC|Cytokeratin Cam5.2 Ag|Cytokeratin Cam5.2 Ag
C1544526|T201|COMP|40562-1|LNC|Actin.muscle specific Ag|Actin.muscle specific Ag
C1544527|T201|COMP|40563-9|LNC|Actin.smooth muscle Ag|Actin.smooth muscle Ag
C1544528|T201|COMP|40564-7|LNC|Thyroid transcription factor 1 Ag|Thyroid transcription factor 1 Ag
C1544529|T201|COMP|40565-4|LNC|Promyelocytes|Promyelocytes
C1544530|T201|COMP|40567-0|LNC|Myelocytes|Myelocytes
C1544531|T201|COMP|40574-6|LNC|Platelets|Platelets
C1544532|T201|COMP|40575-3|LNC|Yersinia enterocolitica O:5,27 Ab|Yersinia enterocolitica O:5,27 Ab
C1544533|T201|COMP|40576-1|LNC|Yersinia enterocolitica O:8 Ab|Yersinia enterocolitica O:8 Ab
C1544534|T201|COMP|40577-9|LNC|Yersinia enterocolitica O:3 Ab|Yersinia enterocolitica O:3 Ab
C1544535|T201|COMP|40578-7|LNC|Cryoglobulin.IgM|Cryoglobulin.IgM
C1544536|T201|COMP|40579-5|LNC|Cryoglobulin.IgG|Cryoglobulin.IgG
C1544537|T201|COMP|40580-3|LNC|Cryoglobulin.IgA|Cryoglobulin.IgA
C1544538|T201|COMP|40581-1|LNC|Cryoglobulin.IgM|Cryoglobulin.IgM
C1544539|T201|COMP|40582-9|LNC|Cryoglobulin.IgG|Cryoglobulin.IgG
C1544540|T201|COMP|40583-7|LNC|Invasive trophoblast Ag|Invasive trophoblast Ag
C1544541|T201|COMP|40584-5|LNC|Arbovirus Ab.IgM|Arbovirus Ab.IgM
C1544542|T201|COMP|40585-2|LNC|Drugs identified|Drugs identified
C1544545|T201|COMP|40588-6|LNC|Inulin|Inulin
C1544552|T201|COMP|40595-1|LNC|Prothrombin Ab.IgG|Prothrombin Ab.IgG
C1544553|T201|COMP|40596-9|LNC|Prothrombin Ab.IgM|Prothrombin Ab.IgM
C1544554|T201|COMP|40597-7|LNC|7-Dehydrocholesterol|7-Dehydrocholesterol
C1544555|T201|COMP|40598-5|LNC|Acetone|Acetone
C1544556|T201|COMP|40599-3|LNC|Albumin|Albumin
C1544557|T201|COMP|40600-9|LNC|Alpha-1-Acid glycoprotein|Alpha-1-Acid glycoprotein
C1544558|T201|COMP|40601-7|LNC|Alpha-1-Acid glycoprotein|Alpha-1-Acid glycoprotein
C1544559|T201|COMP|40602-5|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C1544560|T201|COMP|40603-3|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C1544561|T201|COMP|40604-1|LNC|Alpha-2-Macroglobulin|Alpha-2-Macroglobulin
C1544562|T201|COMP|40605-8|LNC|Alpha-2-Macroglobulin|Alpha-2-Macroglobulin
C1544563|T201|COMP|40606-6|LNC|Appearance|Appearance
C1544564|T201|COMP|40607-4|LNC|Ascaris lumbricoides Ab.IgG|Ascaris lumbricoides Ab.IgG
C1544565|T201|COMP|40608-2|LNC|Ascaris lumbricoides Ab.IgM|Ascaris lumbricoides Ab.IgM
C1544566|T201|COMP|40609-0|LNC|Benzoylecgonine|Benzoylecgonine
C1544567|T201|COMP|40610-8|LNC|Beta-2 transferrin|Beta-2 transferrin
C1544568|T201|COMP|40612-4|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C1544569|T201|COMP|40613-2|LNC|Brucella sp Ab|Brucella sp Ab
C1544570|T201|COMP|40614-0|LNC|Brucella sp Ab|Brucella sp Ab
C1544571|T201|COMP|40615-7|LNC|Calcium oxalate crystals|Calcium oxalate crystals
C1544572|T201|COMP|40616-5|LNC|Campylobacter sp Ab.IgA|Campylobacter sp Ab.IgA
C1544573|T201|COMP|40617-3|LNC|Campylobacter sp Ab.IgG|Campylobacter sp Ab.IgG
C1544574|T201|COMP|40618-1|LNC|Cancer Ag 125|Cancer Ag 125
C1544577|T201|COMP|40621-5|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C1544578|T201|COMP|40622-3|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C1544579|T201|COMP|40623-1|LNC|Cells.CD3+CD4+/100 cells|Cells.CD3+CD4+/100 cells
C1544580|T201|COMP|40624-9|LNC|Cells.CD3+CD8+/100 cells|Cells.CD3+CD8+/100 cells
C1544581|T201|COMP|40625-6|LNC|Cocaine|Cocaine
C1544582|T201|COMP|40626-4|LNC|Codeine|Codeine
C1544583|T201|COMP|40627-2|LNC|Coproporphyrin|Coproporphyrin
C1544584|T201|COMP|40628-0|LNC|Cryoglobulin.IgA|Cryoglobulin.IgA
C1544585|T201|COMP|40629-8|LNC|Doxepin|Doxepin
C1544586|T201|COMP|40630-6|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C1544587|T201|COMP|40631-4|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C1544588|T201|COMP|40632-2|LNC|Gamma globulin/Beta globulin|Gamma globulin/Beta globulin
C1544589|T201|COMP|40633-0|LNC|Hemopexin|Hemopexin
C1544590|T201|COMP|40634-8|LNC|HYDROcodone|HYDROcodone
C1544591|T201|COMP|40635-5|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C1544592|T201|COMP|40636-3|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C1544593|T201|COMP|40637-1|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C1544594|T201|COMP|40638-9|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C1544595|T201|COMP|40639-7|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C1544596|T201|COMP|40640-5|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C1544597|T201|COMP|40641-3|LNC|Ketones|Ketones
C1544598|T201|COMP|40642-1|LNC|Leptospira autumnalis Ab|Leptospira autumnalis Ab
C1544599|T201|COMP|40643-9|LNC|Leptospira borgpetersenii serovar Ballum Ab|Leptospira borgpetersenii serovar Ballum Ab
C1544600|T201|COMP|40644-7|LNC|Leptospira borgpetersenii serovar Sejroe Ab|Leptospira borgpetersenii serovar Sejroe Ab
C1544601|T201|COMP|40645-4|LNC|Leptospira borgpetersenii serovar Tarrasovi Ab|Leptospira borgpetersenii serovar Tarrasovi Ab
C1544602|T201|COMP|40647-0|LNC|Lupus anticoagulant neutralization.platelet|Lupus anticoagulant neutralization.platelet
C1544603|T201|COMP|40648-8|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C1544604|T201|COMP|40649-6|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C1544605|T201|COMP|40650-4|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C1544606|T201|COMP|40651-2|LNC|Metamyelocytes|Metamyelocytes
C1544607|T201|COMP|40652-0|LNC|Methamphetamine|Methamphetamine
C1544608|T201|COMP|40653-8|LNC|Myelocytes/100 leukocytes|Myelocytes/100 leukocytes
C1544609|T201|COMP|40654-6|LNC|Neutrophils.hypogranulated|Neutrophils.hypogranulated
C1544610|T201|COMP|40655-3|LNC|Nuclear Ab|Nuclear Ab
C1544611|T201|COMP|40656-1|LNC|Parasite identified|Parasite identified
C1544612|T201|COMP|40657-9|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C1544613|T201|COMP|40658-7|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C1544614|T201|COMP|40659-5|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C1544615|T201|COMP|40660-3|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C1544616|T201|COMP|40661-1|LNC|Protein.monoclonal|Protein.monoclonal
C1544617|T201|COMP|40662-9|LNC|Protein^resting|Protein^resting
C1544618|T201|COMP|40663-7|LNC|Protein^upright|Protein^upright
C1544619|T201|COMP|40664-5|LNC|Pyrophosphate crystals|Pyrophosphate crystals
C1544620|T201|COMP|40665-2|LNC|Reticulocytes|Reticulocytes
C1544621|T201|COMP|40666-0|LNC|Rubella virus Ab|Rubella virus Ab
C1544622|T201|COMP|40667-8|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C1544623|T201|COMP|40668-6|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C1544624|T201|COMP|40669-4|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C1544625|T201|COMP|40670-2|LNC|Smudge cells/100 leukocytes|Smudge cells/100 leukocytes
C1544626|T201|COMP|40671-0|LNC|Specimen volume|Specimen volume
C1544627|T201|COMP|40672-8|LNC|Sucrose|Sucrose
C1544628|T201|COMP|40673-6|LNC|Thyrotropin binding inhibitory immunoglobulins|Thyrotropin binding inhibitory immunoglobulins
C1544629|T201|COMP|40674-4|LNC|Toxocara canis Ab.IgG|Toxocara canis Ab.IgG
C1544630|T201|COMP|40675-1|LNC|Toxocara canis Ab.IgM|Toxocara canis Ab.IgM
C1544631|T201|COMP|40676-9|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C1544632|T201|COMP|40677-7|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C1544633|T201|COMP|40678-5|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C1544634|T201|COMP|40679-3|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C1544635|T201|COMP|40680-1|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C1544636|T201|COMP|40681-9|LNC|Turbidity|Turbidity
C1544637|T201|COMP|40682-7|LNC|Urate crystals|Urate crystals
C1544638|T201|COMP|40683-5|LNC|Bentiromide|Bentiromide
C1544639|T201|COMP|40684-3|LNC|Acinetobacter sp.multidrug resistant identified|Acinetobacter sp.multidrug resistant identified
C1544640|T201|COMP|40685-0|LNC|Interpretation|Interpretation
C1544641|T201|COMP|40686-8|LNC|Platelet factor 3|Platelet factor 3
C1544642|T201|COMP|40687-6|LNC|Myeloid cells/100 cells|Myeloid cells/100 cells
C1544643|T201|COMP|40688-4|LNC|Megakaryocytes|Megakaryocytes
C1544644|T201|COMP|40689-2|LNC|Erythroid cells/100 cells|Erythroid cells/100 cells
C1544645|T201|COMP|40690-0|LNC|Tumor Ag 90|Tumor Ag 90
C1544646|T201|COMP|40691-8|LNC|Specimen volume^post washing|Specimen volume^post washing
C1544647|T201|COMP|40692-6|LNC|Specimen volume^pre washing|Specimen volume^pre washing
C1544648|T201|COMP|40693-4|LNC|RET gene targeted mutation analysis|RET gene targeted mutation analysis
C1544649|T201|COMP|40694-2|LNC|Sulfamethoxazole Ab.IgE|Sulfamethoxazole Ab.IgE
C1544650|T201|COMP|40695-9|LNC|Spermatozoa^post concentration|Spermatozoa^post concentration
C1544651|T201|COMP|40696-7|LNC|Spermatozoa.motile^post concentration|Spermatozoa.motile^post concentration
C1544652|T201|COMP|40697-5|LNC|Toxoplasma gondii Ab.IgM index|Toxoplasma gondii Ab.IgM index
C1544653|T201|COMP|40698-3|LNC|Mycoplasma sp identified|Mycoplasma sp identified
C1544654|T201|COMP|40699-1|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C1544655|T201|COMP|40700-7|LNC|Aromatic solvents|Aromatic solvents
C1544656|T201|COMP|40701-5|LNC|Arsenic|Arsenic
C1544657|T201|COMP|40702-3|LNC|Fibrin monomer|Fibrin monomer
C1544658|T201|COMP|40703-1|LNC|Lactoferrin|Lactoferrin
C1544659|T201|COMP|40704-9|LNC|Maternal cell contamination|Maternal cell contamination
C1544660|T201|COMP|40705-6|LNC|Brodifacoum|Brodifacoum
C1544661|T201|COMP|40706-4|LNC|Colchicine|Colchicine
C1544662|T201|COMP|40707-2|LNC|Amphotericin B^peak|Amphotericin B^peak
C1544663|T201|COMP|40708-0|LNC|Polio virus Ab.IgG^2nd specimen|Polio virus Ab.IgG^2nd specimen
C1544664|T201|COMP|40709-8|LNC|Polio virus Ab|Polio virus Ab
C1544665|T201|COMP|40710-6|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C1544666|T201|COMP|40711-4|LNC|Clostridium tetani Ab|Clostridium tetani Ab
C1544667|T201|COMP|40712-2|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C1544668|T201|COMP|40713-0|LNC|Giardia lamblia Ab.IgG|Giardia lamblia Ab.IgG
C1544669|T201|COMP|40714-8|LNC|Giardia lamblia Ab.IgM|Giardia lamblia Ab.IgM
C1544670|T201|COMP|40715-5|LNC|Granulocytes.immature|Granulocytes.immature
C1544671|T201|COMP|40716-3|LNC|Hairy cells|Hairy cells
C1544672|T201|COMP|40717-1|LNC|Haptoglobin|Haptoglobin
C1544673|T201|COMP|40718-9|LNC|Heinz bodies/100 erythrocytes|Heinz bodies/100 erythrocytes
C1544674|T201|COMP|40719-7|LNC|Hemoglobin|Hemoglobin
C1544675|T201|COMP|40720-5|LNC|Hemoglobin C|Hemoglobin C
C1544676|T201|COMP|40721-3|LNC|Hemoglobin F|Hemoglobin F
C1544677|T201|COMP|40722-1|LNC|Hemosiderin|Hemosiderin
C1544678|T201|COMP|40723-9|LNC|Heparin Ab|Heparin Ab
C1544679|T201|COMP|40724-7|LNC|Hepatitis A virus Ab.IgG|Hepatitis A virus Ab.IgG
C1544680|T201|COMP|40725-4|LNC|Hepatitis B virus core Ab.IgG|Hepatitis B virus core Ab.IgG
C1544681|T201|COMP|40726-2|LNC|Hepatitis C virus Ab.IgG|Hepatitis C virus Ab.IgG
C1544682|T201|COMP|40727-0|LNC|Hepatitis D virus Ab|Hepatitis D virus Ab
C1544683|T201|COMP|40728-8|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C1544684|T201|COMP|40729-6|LNC|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C1544685|T201|COMP|40730-4|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C1544686|T201|COMP|40731-2|LNC|Herpes virus 6 Ab.IgM|Herpes virus 6 Ab.IgM
C1544687|T201|COMP|40732-0|LNC|HIV 1 Ab.IgG|HIV 1 Ab.IgG
C1544688|T201|COMP|40733-8|LNC|HIV 1+2 Ab.IgG|HIV 1+2 Ab.IgG
C1544689|T201|COMP|40734-6|LNC|HLA Ab|HLA Ab
C1544690|T201|COMP|40735-3|LNC|HTLV I+II Ab.IgG|HTLV I+II Ab.IgG
C1544691|T201|COMP|40736-1|LNC|La Crosse virus Ab|La Crosse virus Ab
C1544692|T201|COMP|40737-9|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C1544693|T201|COMP|40738-7|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C1544694|T201|COMP|40739-5|LNC|Osmotic fragility^unincubated|Osmotic fragility^unincubated
C1544695|T201|COMP|40740-3|LNC|Osmotic fragility^incubated|Osmotic fragility^incubated
C1544696|T201|COMP|40741-1|LNC|Platelet clump|Platelet clump
C1544697|T201|COMP|40742-9|LNC|Rabies virus Ab.IgG|Rabies virus Ab.IgG
C1544698|T201|COMP|40743-7|LNC|Plasma cells|Plasma cells
C1544699|T201|COMP|40744-5|LNC|Factor inhibitor XXX|Factor inhibitor XXX
C1544700|T201|COMP|40745-2|LNC|Filaria identified|Filaria identified
C1544701|T201|COMP|40746-0|LNC|Fragments|Fragments
C1544702|T201|COMP|40747-8|LNC|Complement C2|Complement C2
C1544703|T201|COMP|40748-6|LNC|Dengue virus Ab|Dengue virus Ab
C1544704|T201|COMP|40749-4|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C1544705|T201|COMP|40750-2|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C1544706|T201|COMP|40751-0|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C1544707|T201|COMP|40752-8|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C1544708|T201|COMP|40753-6|LNC|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C1544709|T201|COMP|40754-4|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C1544710|T201|COMP|40755-1|LNC|Amiodarone^peak|Amiodarone^peak
C1544711|T201|COMP|40756-9|LNC|Amiodarone^trough|Amiodarone^trough
C1544712|T201|COMP|40757-7|LNC|Amphotericin B^trough|Amphotericin B^trough
C1544713|T201|COMP|40758-5|LNC|Coxsackievirus A Ab|Coxsackievirus A Ab
C1544714|T201|COMP|40759-3|LNC|Coxsackievirus A Ab.IgM^1st specimen|Coxsackievirus A Ab.IgM^1st specimen
C1544715|T201|COMP|40760-1|LNC|Coxsackievirus A Ab^2nd specimen|Coxsackievirus A Ab^2nd specimen
C1544716|T201|COMP|40761-9|LNC|Coxsackievirus A Ab^2nd specimen|Coxsackievirus A Ab^2nd specimen
C1544717|T201|COMP|40762-7|LNC|Coxsackievirus A Ab^1st specimen|Coxsackievirus A Ab^1st specimen
C1544718|T201|COMP|40763-5|LNC|Coxsackievirus B Ab.IgM^1st specimen|Coxsackievirus B Ab.IgM^1st specimen
C1544719|T201|COMP|40764-3|LNC|Coxsackievirus B Ab.IgG^2nd specimen|Coxsackievirus B Ab.IgG^2nd specimen
C1544720|T201|COMP|40765-0|LNC|Coxsackievirus B Ab|Coxsackievirus B Ab
C1544721|T201|COMP|40766-8|LNC|Coxsackievirus B Ab.IgM^1st specimen|Coxsackievirus B Ab.IgM^1st specimen
C1544722|T201|COMP|40767-6|LNC|Coxsackievirus B Ab.IgG^2nd specimen|Coxsackievirus B Ab.IgG^2nd specimen
C1544723|T201|COMP|40768-4|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1544724|T201|COMP|40769-2|LNC|Ethosuximide^peak|Ethosuximide^peak
C1544725|T201|COMP|40770-0|LNC|Ethosuximide^trough|Ethosuximide^trough
C1544726|T201|COMP|40771-8|LNC|Haemophilus influenzae Ag|Haemophilus influenzae Ag
C1544727|T201|COMP|40772-6|LNC|Heavy metals|Heavy metals
C1544728|T201|COMP|40773-4|LNC|Histoplasma capsulatum Ab.IgM^1st specimen|Histoplasma capsulatum Ab.IgM^1st specimen
C1544729|T201|COMP|40774-2|LNC|Histoplasma capsulatum Ab.IgG^2nd specimen|Histoplasma capsulatum Ab.IgG^2nd specimen
C1544730|T201|COMP|40775-9|LNC|Histoplasma capsulatum Ab.IgM^1st specimen|Histoplasma capsulatum Ab.IgM^1st specimen
C1544731|T201|COMP|40776-7|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1544732|T201|COMP|40777-5|LNC|Histoplasma sp Ab|Histoplasma sp Ab
C1544733|T201|COMP|40778-3|LNC|Histoplasma capsulatum Ab.IgG^2nd specimen|Histoplasma capsulatum Ab.IgG^2nd specimen
C1544734|T201|COMP|40779-1|LNC|Mexiletine^trough|Mexiletine^trough
C1544735|T201|COMP|40780-9|LNC|Mexiletine^peak|Mexiletine^peak
C1544736|T201|COMP|40781-7|LNC|Polio virus Ab.IgM^1st specimen|Polio virus Ab.IgM^1st specimen
C1544737|T201|COMP|40782-5|LNC|Polio virus Ab.IgM^1st specimen|Polio virus Ab.IgM^1st specimen
C1544738|T201|COMP|40783-3|LNC|Polio virus Ab.IgG^2nd specimen|Polio virus Ab.IgG^2nd specimen
C1544739|T201|COMP|40784-1|LNC|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C1544740|T201|COMP|40785-8|LNC|Toxoplasma gondii Ab.IgM^1st specimen|Toxoplasma gondii Ab.IgM^1st specimen
C1544741|T201|COMP|40786-6|LNC|Toxoplasma gondii Ab.IgG^2nd specimen|Toxoplasma gondii Ab.IgG^2nd specimen
C1544742|T201|COMP|40787-4|LNC|Calculus analysis|Calculus analysis
C1544743|T201|COMP|40788-2|LNC|Chamaecyparis obtusa Ab.IgE|Chamaecyparis obtusa Ab.IgE
C1544744|T201|COMP|40789-0|LNC|Humulus japonicus Ab.IgE|Humulus japonicus Ab.IgE
C1544745|T201|COMP|40790-8|LNC|Elaeis guineensis Ab.IgE|Elaeis guineensis Ab.IgE
C1544746|T201|COMP|40791-6|LNC|Coproporphyrin 3|Coproporphyrin 3
C1544747|T201|COMP|40792-4|LNC|Coproporphyrin 1|Coproporphyrin 1
C1544748|T201|COMP|40793-2|LNC|Alkaline phosphatase.placental|Alkaline phosphatase.placental
C1544749|T201|COMP|40794-0|LNC|Alkaline phosphatase.intestinal|Alkaline phosphatase.intestinal
C1544750|T201|COMP|40795-7|LNC|Alkaline phosphatase.liver 2|Alkaline phosphatase.liver 2
C1544751|T201|COMP|40796-5|LNC|Alkaline phosphatase.liver 1|Alkaline phosphatase.liver 1
C1544752|T201|COMP|40797-3|LNC|Alkaline phosphatase.bone|Alkaline phosphatase.bone
C1544753|T201|COMP|40798-1|LNC|Amphetamines|Amphetamines
C1544754|T201|COMP|40799-9|LNC|Amphetamines|Amphetamines
C1544755|T201|COMP|40800-5|LNC|Cannabinoids|Cannabinoids
C1544756|T201|COMP|40801-3|LNC|Cannabinoids|Cannabinoids
C1544757|T201|COMP|40802-1|LNC|Cocaine|Cocaine
C1544758|T201|COMP|40803-9|LNC|Methamphetamine|Methamphetamine
C1544759|T201|COMP|40804-7|LNC|Methamphetamine|Methamphetamine
C1544760|T201|COMP|40805-4|LNC|Opiates|Opiates
C1544761|T201|COMP|40806-2|LNC|Opiates|Opiates
C1544762|T201|COMP|40807-0|LNC|Phencyclidine|Phencyclidine
C1544763|T201|COMP|40808-8|LNC|Phencyclidine|Phencyclidine
C1544764|T201|COMP|40809-6|LNC|11-Deoxycortisol^1H post XXX challenge|11-Deoxycortisol^1H post XXX challenge
C1544765|T201|COMP|40810-4|LNC|11-Deoxycortisol^baseline|11-Deoxycortisol^baseline
C1544766|T201|COMP|40811-2|LNC|11-Deoxycorticosterone|11-Deoxycorticosterone
C1544767|T201|COMP|40812-0|LNC|11-Hydroxyandrosterone/Creatinine|11-Hydroxyandrosterone/Creatinine
C1544768|T201|COMP|40813-8|LNC|11-Hydroxyetiocholanolone/Creatinine|11-Hydroxyetiocholanolone/Creatinine
C1544769|T201|COMP|40814-6|LNC|11-Ketoandrosterone/Creatinine|11-Ketoandrosterone/Creatinine
C1544770|T201|COMP|40815-3|LNC|11-Ketoetiocholanolone/Creatinine|11-Ketoetiocholanolone/Creatinine
C1544771|T201|COMP|40816-1|LNC|11-Deoxycorticosterone^1H post XXX challenge|11-Deoxycorticosterone^1H post XXX challenge
C1544772|T201|COMP|40817-9|LNC|Tetrachlorodiphenylethane|Tetrachlorodiphenylethane
C1544773|T201|COMP|40818-7|LNC|11-Deoxycorticosterone|11-Deoxycorticosterone
C1544774|T201|COMP|40819-5|LNC|Disialylganglioside GD1a Ab.IgM|Disialylganglioside GD1a Ab.IgM
C1544775|T201|COMP|40820-3|LNC|Helicobacter pylori Ab.IgA|Helicobacter pylori Ab.IgA
C1544776|T201|COMP|40821-1|LNC|Helicobacter pylori Ab.IgM|Helicobacter pylori Ab.IgM
C1544777|T201|COMP|40822-9|LNC|HTLV I Ab|HTLV I Ab
C1544778|T201|COMP|40823-7|LNC|HTLV II Ab|HTLV II Ab
C1544779|T201|COMP|40824-5|LNC|von Willebrand factor cleaving protease inhibitor|von Willebrand factor cleaving protease inhibitor
C1544780|T201|COMP|40825-2|LNC|Candida sp Ab.IgG|Candida sp Ab.IgG
C1544781|T201|COMP|40826-0|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C1544782|T201|COMP|40827-8|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C1544783|T201|COMP|40828-6|LNC|Aspergillus fumigatus Ab|Aspergillus fumigatus Ab
C1544784|T201|COMP|40829-4|LNC|Ornithine|Ornithine
C1544785|T201|COMP|40830-2|LNC|Toxocara sp Ab|Toxocara sp Ab
C1544786|T201|COMP|40831-0|LNC|Adenovirus+Rotavirus Ag|Adenovirus+Rotavirus Ag
C1544787|T201|COMP|40832-8|LNC|Pistacia vera Ab.IgE/IgE.total|Pistacia vera Ab.IgE/IgE.total
C1544788|T201|COMP|40833-6|LNC|SOD1 gene allele 1|SOD1 gene allele 1
C1544789|T201|COMP|40834-4|LNC|Herpes virus 8 Ab.IgG|Herpes virus 8 Ab.IgG
C1544790|T201|COMP|40835-1|LNC|Fragaria vesca Ab.IgG|Fragaria vesca Ab.IgG
C1544791|T201|COMP|40836-9|LNC|Sulfonamide crystals|Sulfonamide crystals
C1544792|T201|COMP|40837-7|LNC|Alternaria sp Ab.IgG|Alternaria sp Ab.IgG
C1544793|T201|COMP|40838-5|LNC|Argininosuccinate|Argininosuccinate
C1544794|T201|COMP|40839-3|LNC|fentaNYL|fentaNYL
C1544795|T201|COMP|40840-1|LNC|Legionella pneumophila 1 Ab|Legionella pneumophila 1 Ab
C1544796|T201|COMP|40841-9|LNC|Lycopersicon lycopersicum Ab.IgE/IgE.total|Lycopersicon lycopersicum Ab.IgE/IgE.total
C1544797|T201|COMP|40842-7|LNC|Galactose 1 phosphate|Galactose 1 phosphate
C1544798|T201|COMP|40843-5|LNC|Chicken meat Ab.IgE/IgE.total|Chicken meat Ab.IgE/IgE.total
C1544800|T201|COMP|40845-0|LNC|Turkey meat Ab.IgE/IgE.total|Turkey meat Ab.IgE/IgE.total
C1544801|T201|COMP|40846-8|LNC|Homovanillate|Homovanillate
C1544802|T201|COMP|40847-6|LNC|Bromus inermis Ab.IgG4|Bromus inermis Ab.IgG4
C1544803|T201|COMP|40848-4|LNC|3-Methylcrotonylglycine|3-Methylcrotonylglycine
C1544804|T201|COMP|40849-2|LNC|Glucose^1st specimen post XXX challenge|Glucose^1st specimen post XXX challenge
C1544805|T201|COMP|40850-0|LNC|Glucose^2nd specimen post XXX challenge|Glucose^2nd specimen post XXX challenge
C1544806|T201|COMP|40851-8|LNC|Normetanephrine.free|Normetanephrine.free
C1544807|T201|COMP|40852-6|LNC|Leishmania sp Ab.IgG|Leishmania sp Ab.IgG
C1544808|T201|COMP|40853-4|LNC|Leishmania sp Ab.IgG|Leishmania sp Ab.IgG
C1544809|T201|COMP|40854-2|LNC|Chlamydia trachomatis L2 Ab.IgG|Chlamydia trachomatis L2 Ab.IgG
C1544810|T201|COMP|40855-9|LNC|Chlamydia trachomatis L2 Ab.IgA|Chlamydia trachomatis L2 Ab.IgA
C1544811|T201|COMP|40856-7|LNC|Chlamydia trachomatis L2 Ab.IgM|Chlamydia trachomatis L2 Ab.IgM
C1544812|T201|COMP|40857-5|LNC|Prealbumin|Prealbumin
C1544813|T201|COMP|40858-3|LNC|Glucose^baseline|Glucose^baseline
C1544814|T201|COMP|40859-1|LNC|SOD1 gene allele 2|SOD1 gene allele 2
C1544815|T201|COMP|40860-9|LNC|Cytokines|Cytokines
C1544816|T201|COMP|40861-7|LNC|Cells.CD103/100 cells|Cells.CD103/100 cells
C1544817|T201|COMP|40862-5|LNC|Methylparaben Ab.IgE|Methylparaben Ab.IgE
C1544818|T201|COMP|40863-3|LNC|Norovirus Genogroup I Ag|Norovirus Genogroup I Ag
C1544819|T201|COMP|40864-1|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C1544820|T201|COMP|40865-8|LNC|11-Oxo-Androsterone|11-Oxo-Androsterone
C1544821|T201|COMP|40866-6|LNC|11-Oxo-Androsterone/Creatinine|11-Oxo-Androsterone/Creatinine
C1544822|T201|COMP|40867-4|LNC|11-Oxo-Etiocholanolone|11-Oxo-Etiocholanolone
C1544823|T201|COMP|40868-2|LNC|11-Oxo-Etiocholanolone/Creatinine|11-Oxo-Etiocholanolone/Creatinine
C1544824|T201|COMP|40869-0|LNC|Carnitine esters/Carnitine.free (C0)|Carnitine esters/Carnitine.free (C0)
C1544825|T201|COMP|40870-8|LNC|Cystine.free|Cystine.free
C1544826|T201|COMP|40871-6|LNC|CNBP gene targeted mutation analysis|CNBP gene targeted mutation analysis
C1544827|T201|COMP|40872-4|LNC|CBS gene.c.833T>C|CBS gene.c.833T>C
C1544828|T201|COMP|40873-2|LNC|CBS gene.c.919G>A|CBS gene.c.919G>A
C1544829|T201|COMP|40874-0|LNC|Glucose^1st specimen|Glucose^1st specimen
C1544830|T201|COMP|40875-7|LNC|Glucose^3rd specimen|Glucose^3rd specimen
C1544831|T201|COMP|40876-5|LNC|AMPD1 gene.p.Gln12Ter+AMPD1 gene.p.Pro48Leu|AMPD1 gene.p.Gln12Ter+AMPD1 gene.p.Pro48Leu
C1544832|T201|COMP|40877-3|LNC|CPT2 gene.p.Pro50His+Ser113Leu|CPT2 gene.p.Pro50His+Ser113Leu
C1544833|T201|COMP|40878-1|LNC|CPT2 gene.p.Gln413FSer+Gly549Asp|CPT2 gene.p.Gln413FSer+Gly549Asp
C1544834|T201|COMP|40879-9|LNC|Chicken Ab.IgE|Chicken Ab.IgE
C1544835|T201|COMP|40880-7|LNC|Cells.CD3-CD56+/100 cells|Cells.CD3-CD56+/100 cells
C1544836|T201|COMP|40881-5|LNC|Cells.CD3-CD57+/100 cells|Cells.CD3-CD57+/100 cells
C1544837|T201|COMP|40882-3|LNC|Cells.CD3-CD57+/100 cells|Cells.CD3-CD57+/100 cells
C1544838|T201|COMP|40883-1|LNC|Cells.CD19+CD103+/100 cells|Cells.CD19+CD103+/100 cells
C1544839|T201|COMP|40884-9|LNC|Cells.CD19+CD103+/100 cells|Cells.CD19+CD103+/100 cells
C1544840|T201|COMP|40885-6|LNC|Cells.CD19+CD103+/100 cells|Cells.CD19+CD103+/100 cells
C1544841|T201|COMP|40886-4|LNC|Cells.CD19+CD103+/100 cells|Cells.CD19+CD103+/100 cells
C1544842|T201|COMP|40887-2|LNC|Cells.CD11c+CD19+/100 cells|Cells.CD11c+CD19+/100 cells
C1544843|T201|COMP|40888-0|LNC|Cells.CD11c+CD19+/100 cells|Cells.CD11c+CD19+/100 cells
C1544844|T201|COMP|40889-8|LNC|Cells.CD25+CD19+/100 cells|Cells.CD25+CD19+/100 cells
C1544845|T201|COMP|40890-6|LNC|Cells.CD25+CD19+/100 cells|Cells.CD25+CD19+/100 cells
C1544846|T201|COMP|40891-4|LNC|Cells.CD3-CD57+|Cells.CD3-CD57+
C1544847|T201|COMP|40892-2|LNC|Cells.CD3-CD16+/100 cells|Cells.CD3-CD16+/100 cells
C1544848|T201|COMP|40893-0|LNC|Cells.CD3-CD16+/100 cells|Cells.CD3-CD16+/100 cells
C1544849|T201|COMP|40894-8|LNC|Cells.CD3-CD16+/100 cells|Cells.CD3-CD16+/100 cells
C1544850|T201|COMP|40895-5|LNC|Cells.CD3+CD56+|Cells.CD3+CD56+
C1544851|T201|COMP|40896-3|LNC|Cells.CD3+CD56+|Cells.CD3+CD56+
C1544852|T201|COMP|40897-1|LNC|Cells.CD3+CD56+|Cells.CD3+CD56+
C1544853|T201|COMP|40898-9|LNC|Cells.CD3+CD4+|Cells.CD3+CD4+
C1544854|T201|COMP|40899-7|LNC|Cells.CD3+CD8+|Cells.CD3+CD8+
C1544855|T201|COMP|40900-3|LNC|Cells.CD3+CD4+/Cells.CD3+CD8+|Cells.CD3+CD4+/Cells.CD3+CD8+
C1544856|T201|COMP|40901-1|LNC|3-Hydroxybenzoylecgonine|3-Hydroxybenzoylecgonine
C1544857|T201|COMP|40902-9|LNC|Streptococcus pneumoniae 12 Ab.IgG^2nd specimen|Streptococcus pneumoniae 12 Ab.IgG^2nd specimen
C1544858|T201|COMP|40903-7|LNC|Streptococcus pneumoniae 12 Ab.IgG|Streptococcus pneumoniae 12 Ab.IgG
C1544859|T201|COMP|40904-5|LNC|Streptococcus pneumoniae 12 Ab.IgG^1st specimen|Streptococcus pneumoniae 12 Ab.IgG^1st specimen
C1544863|T201|COMP|40908-6|LNC|Streptococcus pneumoniae 4 Ab.IgG|Streptococcus pneumoniae 4 Ab.IgG
C1544867|T201|COMP|40920-1|LNC|Streptococcus pneumoniae 8 Ab.IgG|Streptococcus pneumoniae 8 Ab.IgG
C1544868|T201|COMP|40921-9|LNC|Streptococcus pneumoniae 8 Ab.IgG^1st specimen|Streptococcus pneumoniae 8 Ab.IgG^1st specimen
C1544869|T201|COMP|40922-7|LNC|Streptococcus pneumoniae 8 Ab.IgG^2nd specimen|Streptococcus pneumoniae 8 Ab.IgG^2nd specimen
C1544870|T201|COMP|40923-5|LNC|Streptococcus pneumoniae 9 Ab.IgG|Streptococcus pneumoniae 9 Ab.IgG
C1544871|T201|COMP|40924-3|LNC|Streptococcus pneumoniae 9 Ab.IgG^1st specimen|Streptococcus pneumoniae 9 Ab.IgG^1st specimen
C1544872|T201|COMP|40925-0|LNC|Streptococcus pneumoniae 9 Ab.IgG^2nd specimen|Streptococcus pneumoniae 9 Ab.IgG^2nd specimen
C1544874|T201|COMP|40927-6|LNC|3-Methylcrotonylglycine|3-Methylcrotonylglycine
C1544875|T201|COMP|40928-4|LNC|Cortisol^pre dose dexamethasone|Cortisol^pre dose dexamethasone
C1544876|T201|COMP|40929-2|LNC|Parathyrin.intact^10M post excision|Parathyrin.intact^10M post excision
C1544877|T201|COMP|40930-0|LNC|PYGM gene.p.Arg50Ter+Gly205Ser|PYGM gene.p.Arg50Ter+Gly205Ser
C1544878|T201|COMP|40931-8|LNC|Yersinia sp Ab|Yersinia sp Ab
C1544879|T201|COMP|40932-6|LNC|Yersinia enterocolitica O:3 Ab|Yersinia enterocolitica O:3 Ab
C1544880|T201|COMP|40933-4|LNC|Yersinia enterocolitica O:5 Ab|Yersinia enterocolitica O:5 Ab
C1544881|T201|COMP|40934-2|LNC|Yersinia enterocolitica O:8 Ab|Yersinia enterocolitica O:8 Ab
C1544882|T201|COMP|40935-9|LNC|Yersinia enterocolitica O:9 Ab|Yersinia enterocolitica O:9 Ab
C1544883|T201|COMP|40936-7|LNC|Yersinia pseudotuberculosis Ab|Yersinia pseudotuberculosis Ab
C1544884|T201|COMP|40937-5|LNC|Zinc|Zinc
C1544885|T201|COMP|40938-3|LNC|Yersinia sp Ab.IgG|Yersinia sp Ab.IgG
C1544886|T201|COMP|40939-1|LNC|Yersinia sp Ab.IgM|Yersinia sp Ab.IgM
C1544887|T201|COMP|40940-9|LNC|Yersinia sp Ab|Yersinia sp Ab
C1544888|T201|COMP|40941-7|LNC|Yersinia enterocolitica Ab|Yersinia enterocolitica Ab
C1544889|T201|COMP|40942-5|LNC|Yersinia sp Ab.IgM|Yersinia sp Ab.IgM
C1544890|T201|COMP|40943-3|LNC|Vespula spp Ab.IgE|Vespula spp Ab.IgE
C1544891|T201|COMP|40944-1|LNC|Yohimbine|Yohimbine
C1544892|T201|COMP|40945-8|LNC|Yersinia enterocolitica Ab.IgA|Yersinia enterocolitica Ab.IgA
C1544893|T201|COMP|40946-6|LNC|Yersinia enterocolitica Ab.IgG|Yersinia enterocolitica Ab.IgG
C1544894|T201|COMP|40947-4|LNC|Zinc|Zinc
C1544895|T201|COMP|40948-2|LNC|Yersinia enterocolitica O:3 Ab|Yersinia enterocolitica O:3 Ab
C1544896|T201|COMP|40949-0|LNC|Yersinia enterocolitica O:5 Ab|Yersinia enterocolitica O:5 Ab
C1544897|T201|COMP|40950-8|LNC|Yersinia enterocolitica O:8 Ab|Yersinia enterocolitica O:8 Ab
C1544898|T201|COMP|40951-6|LNC|Yersinia enterocolitica O:9 Ab|Yersinia enterocolitica O:9 Ab
C1544899|T201|COMP|40952-4|LNC|Vespula spp Ab.IgG4|Vespula spp Ab.IgG4
C1544900|T201|COMP|40953-2|LNC|Yersinia enterocolitica O:3 Ab|Yersinia enterocolitica O:3 Ab
C1544901|T201|COMP|40954-0|LNC|Yersinia enterocolitica O:8 Ab|Yersinia enterocolitica O:8 Ab
C1544902|T201|COMP|40955-7|LNC|Yersinia enterocolitica O:9 Ab|Yersinia enterocolitica O:9 Ab
C1544903|T201|COMP|40956-5|LNC|Yersinia sp Ab|Yersinia sp Ab
C1544904|T201|COMP|40957-3|LNC|Zinc|Zinc
C1544905|T201|COMP|40958-1|LNC|Cryptosporidium parvum identified|Cryptosporidium parvum identified
C1544906|T201|COMP|40959-9|LNC|MUTYH gene targeted mutation analysis|MUTYH gene targeted mutation analysis
C1544907|T201|COMP|40960-7|LNC|Parietal cell Ab.IgG|Parietal cell Ab.IgG
C1544908|T201|COMP|40961-5|LNC|SFTPB gene targeted mutation analysis|SFTPB gene targeted mutation analysis
C1544909|T201|COMP|40962-3|LNC|SFTPC gene targeted mutation analysis|SFTPC gene targeted mutation analysis
C1544910|T201|COMP|40963-1|LNC|Streptococcus pneumoniae 17 Ab.IgG|Streptococcus pneumoniae 17 Ab.IgG
C1544911|T201|COMP|40964-9|LNC|Streptococcus pneumoniae 2 Ab.IgG|Streptococcus pneumoniae 2 Ab.IgG
C1544912|T201|COMP|40965-6|LNC|Streptococcus pneumoniae 20 Ab.IgG|Streptococcus pneumoniae 20 Ab.IgG
C1544913|T201|COMP|40966-4|LNC|Streptococcus pneumoniae 22 Ab.IgG|Streptococcus pneumoniae 22 Ab.IgG
C1544914|T201|COMP|40967-2|LNC|Streptococcus pneumoniae 34 Ab.IgG|Streptococcus pneumoniae 34 Ab.IgG
C1544915|T201|COMP|40968-0|LNC|Streptococcus pneumoniae 43 Ab.IgG|Streptococcus pneumoniae 43 Ab.IgG
C1544917|T201|COMP|40970-6|LNC|VWF gene targeted mutation analysis|VWF gene targeted mutation analysis
C1544918|T201|COMP|40971-4|LNC|XXX microorganism DNA|XXX microorganism DNA
C1544919|T201|COMP|40972-2|LNC|XXX microorganism DNA|XXX microorganism DNA
C1544922|T201|COMP|40975-5|LNC|Adenovirus DNA|Adenovirus DNA
C1544923|T201|COMP|40976-3|LNC|Adenovirus DNA|Adenovirus DNA
C1544924|T201|COMP|40977-1|LNC|Adenovirus Ab.IgG|Adenovirus Ab.IgG
C1544925|T201|COMP|40978-9|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C1544926|T201|COMP|40979-7|LNC|Human metapneumovirus Ag|Human metapneumovirus Ag
C1544927|T201|COMP|40980-5|LNC|Human metapneumovirus Ab.IgG|Human metapneumovirus Ab.IgG
C1544928|T201|COMP|40981-3|LNC|Influenza virus A RNA|Influenza virus A RNA
C1544929|T201|COMP|40982-1|LNC|Influenza virus B RNA|Influenza virus B RNA
C1544930|T201|COMP|40983-9|LNC|Parainfluenza virus 1 Ab.IgG|Parainfluenza virus 1 Ab.IgG
C1544931|T201|COMP|40984-7|LNC|Parainfluenza virus 2 Ab.IgG|Parainfluenza virus 2 Ab.IgG
C1544932|T201|COMP|40985-4|LNC|Parainfluenza virus 3 Ab.IgG|Parainfluenza virus 3 Ab.IgG
C1544933|T201|COMP|40986-2|LNC|Parainfluenza virus 4 Ag|Parainfluenza virus 4 Ag
C1544934|T201|COMP|40987-0|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C1544935|T201|COMP|40988-8|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C1544936|T201|COMP|40989-6|LNC|Respiratory syncytial virus Ab.IgG|Respiratory syncytial virus Ab.IgG
C1544937|T201|COMP|40990-4|LNC|Rhinovirus RNA|Rhinovirus RNA
C1544938|T201|COMP|40991-2|LNC|Rhinovirus+Enterovirus RNA|Rhinovirus+Enterovirus RNA
C1544939|T201|COMP|40992-0|LNC|Rhinovirus+Enterovirus Ag|Rhinovirus+Enterovirus Ag
C1544940|T201|COMP|40993-8|LNC|Rhinovirus Ag|Rhinovirus Ag
C1544941|T201|COMP|40994-6|LNC|CPEO syndrome gene targeted mutation analysis|CPEO syndrome gene targeted mutation analysis
C1544942|T201|COMP|40995-3|LNC|Mitochondria DNA targeted mutation analysis|Mitochondria DNA targeted mutation analysis
C1544943|T201|COMP|40996-1|LNC|Alternaria alternata Ab.IgE/IgE.total|Alternaria alternata Ab.IgE/IgE.total
C1544944|T201|COMP|40997-9|LNC|Apis mellifera Ab.IgE/IgE.total|Apis mellifera Ab.IgE/IgE.total
C1544945|T201|COMP|40998-7|LNC|Calcium hydrogen phosphate dihydrate/Total|Calcium hydrogen phosphate dihydrate/Total
C1544946|T201|COMP|40999-5|LNC|Calcium hydrogen phosphate dihydrate|Calcium hydrogen phosphate dihydrate
C1544947|T201|COMP|41000-1|LNC|Human coronavirus RNA|Human coronavirus RNA
C1544948|T201|COMP|41001-9|LNC|Human coronavirus RNA|Human coronavirus RNA
C1544949|T201|COMP|41002-7|LNC|Human coronavirus 229E Ab.IgG|Human coronavirus 229E Ab.IgG
C1544950|T201|COMP|41003-5|LNC|Human coronavirus 229E RNA|Human coronavirus 229E RNA
C1544951|T201|COMP|41004-3|LNC|Human coronavirus 229E Ag|Human coronavirus 229E Ag
C1544952|T201|COMP|41005-0|LNC|Human coronavirus NL63 RNA|Human coronavirus NL63 RNA
C1544953|T201|COMP|41006-8|LNC|Human coronavirus NL63 Ab.IgG|Human coronavirus NL63 Ab.IgG
C1544954|T201|COMP|41007-6|LNC|Human coronavirus OC43 Ag|Human coronavirus OC43 Ag
C1544955|T201|COMP|41008-4|LNC|Human coronavirus OC43 Ab.IgG|Human coronavirus OC43 Ab.IgG
C1544956|T201|COMP|41009-2|LNC|Human coronavirus OC43 RNA|Human coronavirus OC43 RNA
C1544957|T201|COMP|41010-0|LNC|Parainfluenza virus 4 RNA|Parainfluenza virus 4 RNA
C1544958|T201|COMP|41011-8|LNC|Human metapneumovirus Ab.IgG|Human metapneumovirus Ab.IgG
C1544959|T201|COMP|41012-6|LNC|Respiratory syncytial virus Ab.IgG|Respiratory syncytial virus Ab.IgG
C1544960|T201|COMP|41013-4|LNC|Human coronavirus 229E Ab.IgG|Human coronavirus 229E Ab.IgG
C1544961|T201|COMP|41014-2|LNC|Human coronavirus NL63 Ab.IgG|Human coronavirus NL63 Ab.IgG
C1544962|T201|COMP|41015-9|LNC|Human coronavirus OC43 Ab.IgG|Human coronavirus OC43 Ab.IgG
C1544963|T201|COMP|41016-7|LNC|Bilirubin|Bilirubin
C1544964|T201|COMP|41017-5|LNC|Protoporphyrin|Protoporphyrin
C1544965|T201|COMP|41018-3|LNC|Testosterone.free+weakly bound|Testosterone.free+weakly bound
C1544966|T201|COMP|41019-1|LNC|Beta endorphin|Beta endorphin
C1544967|T201|COMP|41020-9|LNC|Flunitrazepam|Flunitrazepam
C1544968|T201|COMP|41021-7|LNC|Cocaine|Cocaine
C1544969|T201|COMP|41022-5|LNC|Citrate|Citrate
C1544970|T201|COMP|41023-3|LNC|Aldosterone|Aldosterone
C1544971|T201|COMP|41024-1|LNC|Glucose^2H post 50 g glucose PO|Glucose^2H post 50 g glucose PO
C1544972|T201|COMP|41025-8|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C1544973|T201|COMP|41026-6|LNC|Fungus identified|Fungus identified
C1544974|T201|COMP|41027-4|LNC|Tau protein/Amyloid beta 42 peptide|Tau protein/Amyloid beta 42 peptide
C1544975|T201|COMP|41028-2|LNC|Listeria monocytogenes O1 Ab|Listeria monocytogenes O1 Ab
C1544976|T201|COMP|41029-0|LNC|Listeria monocytogenes H1 Ab|Listeria monocytogenes H1 Ab
C1544977|T201|COMP|41030-8|LNC|Listeria monocytogenes O4b Ab|Listeria monocytogenes O4b Ab
C1544978|T201|COMP|41031-6|LNC|Lopinavir|Lopinavir
C1544979|T201|COMP|41032-4|LNC|Uroporphyrin|Uroporphyrin
C1544980|T201|COMP|41033-2|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C1544981|T201|COMP|41034-0|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C1544982|T201|COMP|41035-7|LNC|Norovirus RNA|Norovirus RNA
C1544983|T201|COMP|41036-5|LNC|Cocaine|Cocaine
C1544984|T201|COMP|41037-3|LNC|Cocaine|Cocaine
C1544985|T201|COMP|41038-1|LNC|Codeine|Codeine
C1544986|T201|COMP|41039-9|LNC|3-Methylcrotonylglycine|3-Methylcrotonylglycine
C1544987|T201|COMP|41040-7|LNC|Palmitoylcarnitine (C16)|Palmitoylcarnitine (C16)
C1544988|T201|COMP|41041-5|LNC|3-Hydroxypalmitoylcarnitine (C16-OH)|3-Hydroxypalmitoylcarnitine (C16-OH)
C1544989|T201|COMP|41042-3|LNC|WFS1 gene targeted mutation analysis|WFS1 gene targeted mutation analysis
C1544990|T201|COMP|41043-1|LNC|VHL gene targeted mutation analysis|VHL gene targeted mutation analysis
C1544991|T201|COMP|41044-9|LNC|UGT1A1 gene targeted mutation analysis|UGT1A1 gene targeted mutation analysis
C1544992|T201|COMP|41045-6|LNC|TYR gene targeted mutation analysis|TYR gene targeted mutation analysis
C1544993|T201|COMP|41046-4|LNC|TWIST1 gene targeted mutation analysis|TWIST1 gene targeted mutation analysis
C1544994|T201|COMP|41047-2|LNC|TSC gene targeted mutation analysis|TSC gene targeted mutation analysis
C1544995|T201|COMP|41049-8|LNC|TNFRSF1A gene targeted mutation analysis|TNFRSF1A gene targeted mutation analysis
C1544996|T201|COMP|41050-6|LNC|TH gene targeted mutation analysis|TH gene targeted mutation analysis
C1544997|T201|COMP|41051-4|LNC|SPINK1 gene targeted mutation analysis|SPINK1 gene targeted mutation analysis
C1544998|T201|COMP|41053-0|LNC|SMN1 gene targeted mutation analysis|SMN1 gene targeted mutation analysis
C1545000|T201|COMP|41114-0|LNC|CATCH22 syndrome gene targeted mutation analysis|CATCH22 syndrome gene targeted mutation analysis
C1545001|T201|COMP|41115-7|LNC|NOD2 gene targeted mutation analysis|NOD2 gene targeted mutation analysis
C1545002|T201|COMP|41116-5|LNC|ATP7A gene targeted mutation analysis|ATP7A gene targeted mutation analysis
C1545003|T201|COMP|41118-1|LNC|AR gene targeted mutation analysis|AR gene targeted mutation analysis
C1545004|T201|COMP|41119-9|LNC|APTX gene targeted mutation analysis|APTX gene targeted mutation analysis
C1545005|T201|COMP|41121-5|LNC|ACADS gene targeted mutation analysis|ACADS gene targeted mutation analysis
C1545006|T201|COMP|41122-3|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1545007|T201|COMP|41123-1|LNC|Toxoplasma gondii HS Ab|Toxoplasma gondii HS Ab
C1545008|T201|COMP|41055-5|LNC|SLC26A4 gene targeted mutation analysis|SLC26A4 gene targeted mutation analysis
C1545009|T201|COMP|41056-3|LNC|SLC22A18 gene targeted mutation analysis|SLC22A18 gene targeted mutation analysis
C1545010|T201|COMP|41057-1|LNC|SHOX gene targeted mutation analysis|SHOX gene targeted mutation analysis
C1545011|T201|COMP|41058-9|LNC|SH2D1A gene targeted mutation analysis|SH2D1A gene targeted mutation analysis
C1545012|T201|COMP|41059-7|LNC|SFTPC gene targeted mutation analysis|SFTPC gene targeted mutation analysis
C1545013|T201|COMP|41060-5|LNC|SFTPB gene targeted mutation analysis|SFTPB gene targeted mutation analysis
C1545014|T201|COMP|41062-1|LNC|SDHB gene targeted mutation analysis|SDHB gene targeted mutation analysis
C1545015|T201|COMP|41063-9|LNC|RPS6KA3 gene targeted mutation analysis|RPS6KA3 gene targeted mutation analysis
C1545016|T201|COMP|41064-7|LNC|PYGM gene targeted mutation analysis|PYGM gene targeted mutation analysis
C1545017|T201|COMP|41065-4|LNC|PTPN11 gene targeted mutation analysis|PTPN11 gene targeted mutation analysis
C1545018|T201|COMP|41066-2|LNC|PRX gene targeted mutation analysis|PRX gene targeted mutation analysis
C1545019|T201|COMP|41067-0|LNC|PRF1 gene targeted mutation analysis|PRF1 gene targeted mutation analysis
C1545020|T201|COMP|41069-6|LNC|PPT1 gene targeted mutation analysis|PPT1 gene targeted mutation analysis
C1545022|T201|COMP|41071-2|LNC|PARK2 gene targeted mutation analysis|PARK2 gene targeted mutation analysis
C1545023|T201|COMP|41072-0|LNC|PANK2 gene targeted mutation analysis|PANK2 gene targeted mutation analysis
C1545024|T201|COMP|41073-8|LNC|NR0B1 gene targeted mutation analysis|NR0B1 gene targeted mutation analysis
C1545025|T201|COMP|41074-6|LNC|NPHS1 gene targeted mutation analysis|NPHS1 gene targeted mutation analysis
C1545026|T201|COMP|41076-1|LNC|NPDC gene targeted mutation analysis|NPDC gene targeted mutation analysis
C1545027|T201|COMP|41077-9|LNC|NOTCH3 gene targeted mutation analysis|NOTCH3 gene targeted mutation analysis
C1545028|T201|COMP|41078-7|LNC|NIPBL gene targeted mutation analysis|NIPBL gene targeted mutation analysis
C1545029|T201|COMP|41079-5|LNC|NEFL gene targeted mutation analysis|NEFL gene targeted mutation analysis
C1545031|T201|COMP|41081-1|LNC|MUTYH gene targeted mutation analysis|MUTYH gene targeted mutation analysis
C1545032|T201|COMP|41083-7|LNC|MTM1 gene targeted mutation analysis|MTM1 gene targeted mutation analysis
C1545033|T201|COMP|41085-2|LNC|MPZ gene targeted mutation analysis|MPZ gene targeted mutation analysis
C1545034|T201|COMP|41086-0|LNC|MLH1 gene targeted mutation analysis|MLH1 gene targeted mutation analysis
C1545036|T201|COMP|41089-4|LNC|MEN1 gene targeted mutation analysis|MEN1 gene targeted mutation analysis
C1545037|T201|COMP|41090-2|LNC|MELAS gene targeted mutation analysis|MELAS gene targeted mutation analysis
C1545038|T201|COMP|41091-0|LNC|MEFV gene targeted mutation analysis|MEFV gene targeted mutation analysis
C1545039|T201|COMP|41092-8|LNC|MAPT gene targeted mutation analysis|MAPT gene targeted mutation analysis
C1545040|T201|COMP|41093-6|LNC|LHON syndrome gene targeted mutation analysis|LHON syndrome gene targeted mutation analysis
C1545041|T201|COMP|41095-1|LNC|L1CAM gene targeted mutation analysis|L1CAM gene targeted mutation analysis
C1545042|T201|COMP|41096-9|LNC|KEL gene targeted mutation analysis|KEL gene targeted mutation analysis
C1545043|T201|COMP|41097-7|LNC|HADHA gene.c.1528G>C|HADHA gene.c.1528G>C
C1545044|T201|COMP|41098-5|LNC|GPC3 gene targeted mutation analysis|GPC3 gene targeted mutation analysis
C1545045|T201|COMP|41100-9|LNC|GJB6 gene targeted mutation analysis|GJB6 gene targeted mutation analysis
C1545046|T201|COMP|41102-5|LNC|GJB1 gene targeted mutation analysis|GJB1 gene targeted mutation analysis
C1545047|T201|COMP|41103-3|LNC|Gene XXX targeted mutation analysis|Gene XXX targeted mutation analysis
C1545048|T201|COMP|41105-8|LNC|FSHD gene targeted mutation analysis|FSHD gene targeted mutation analysis
C1545049|T201|COMP|41106-6|LNC|FXN gene targeted mutation analysis|FXN gene targeted mutation analysis
C1545050|T201|COMP|41108-2|LNC|FGF23 gene targeted mutation analysis|FGF23 gene targeted mutation analysis
C1545051|T201|COMP|41109-0|LNC|FGD1 gene targeted mutation analysis|FGD1 gene targeted mutation analysis
C1545052|T201|COMP|41124-9|LNC|Toxoplasma gondii AC Ab|Toxoplasma gondii AC Ab
C1545053|T201|COMP|41125-6|LNC|Strongyloides sp Ab.IgG|Strongyloides sp Ab.IgG
C1545054|T201|COMP|41126-4|LNC|Salmonella typhi O D Ab|Salmonella typhi O D Ab
C1545055|T201|COMP|41127-2|LNC|Salmonella gallinarum Ab|Salmonella gallinarum Ab
C1545056|T201|COMP|41128-0|LNC|Rabies virus Ab.IgG|Rabies virus Ab.IgG
C1545057|T201|COMP|41129-8|LNC|Parvovirus B19 Ab.IgM^1st specimen|Parvovirus B19 Ab.IgM^1st specimen
C1545059|T201|COMP|41131-4|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C1545060|T201|COMP|41132-2|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C1545061|T201|COMP|41133-0|LNC|Jamestown canyon virus Ab|Jamestown canyon virus Ab
C1545062|T201|COMP|41134-8|LNC|Influenza virus A N9 Ab|Influenza virus A N9 Ab
C1545063|T201|COMP|41135-5|LNC|Influenza virus A N8 Ab|Influenza virus A N8 Ab
C1545064|T201|COMP|41136-3|LNC|Influenza virus A N7 Ab|Influenza virus A N7 Ab
C1545065|T201|COMP|41137-1|LNC|Influenza virus A N6 Ab|Influenza virus A N6 Ab
C1545066|T201|COMP|41138-9|LNC|Influenza virus A N5 Ab|Influenza virus A N5 Ab
C1545067|T201|COMP|41139-7|LNC|Influenza virus A N4 Ab|Influenza virus A N4 Ab
C1545068|T201|COMP|41140-5|LNC|Influenza virus A N3 Ab|Influenza virus A N3 Ab
C1545069|T201|COMP|41141-3|LNC|Influenza virus A N2 Ab|Influenza virus A N2 Ab
C1545070|T201|COMP|41142-1|LNC|Influenza virus A N1 Ab|Influenza virus A N1 Ab
C1545071|T201|COMP|41143-9|LNC|HIV 1 Ab|HIV 1 Ab
C1545072|T201|COMP|41144-7|LNC|HIV 1 Ab|HIV 1 Ab
C1545073|T201|COMP|41145-4|LNC|HIV 1 Ab|HIV 1 Ab
C1545074|T201|COMP|41146-2|LNC|Herpes virus 8 Ab.IgG|Herpes virus 8 Ab.IgG
C1545075|T201|COMP|41147-0|LNC|Herpes virus 6 Ab.IgM|Herpes virus 6 Ab.IgM
C1545076|T201|COMP|41148-8|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C1545077|T201|COMP|41149-6|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1545078|T201|COMP|41150-4|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1545079|T201|COMP|41151-2|LNC|Hepatitis B virus little e Ab.IgG|Hepatitis B virus little e Ab.IgG
C1545080|T201|COMP|41152-0|LNC|Haemophilus paragallinarum Ab|Haemophilus paragallinarum Ab
C1545081|T201|COMP|41153-8|LNC|Giardia lamblia Ab.IgM|Giardia lamblia Ab.IgM
C1545082|T201|COMP|41154-6|LNC|Giardia lamblia Ab.IgG|Giardia lamblia Ab.IgG
C1545083|T201|COMP|41155-3|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C1545084|T201|COMP|41156-1|LNC|Coccidioides sp Ab.IgG|Coccidioides sp Ab.IgG
C1545085|T201|COMP|41157-9|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C1545086|T201|COMP|41158-7|LNC|Canine herpesvirus Ab|Canine herpesvirus Ab
C1545087|T201|COMP|41159-5|LNC|Campylobacter sp Ab.IgG|Campylobacter sp Ab.IgG
C1545088|T201|COMP|41160-3|LNC|Ascaris lumbricoides Ab.IgM|Ascaris lumbricoides Ab.IgM
C1545089|T201|COMP|41161-1|LNC|Ascaris lumbricoides Ab.IgG|Ascaris lumbricoides Ab.IgG
C1545090|T201|COMP|41162-9|LNC|Adenovirus Ab.IgG|Adenovirus Ab.IgG
C1545091|T201|COMP|41163-7|LNC|Treponema pallidum DNA|Treponema pallidum DNA
C1545092|T201|COMP|41164-5|LNC|Uranium.depleted|Uranium.depleted
C1545093|T201|COMP|41165-2|LNC|Uranium 235/Uranium 238|Uranium 235/Uranium 238
C1545094|T201|COMP|41166-0|LNC|Uranium.depleted/Creatinine|Uranium.depleted/Creatinine
C1545095|T201|COMP|41167-8|LNC|Listeria monocytogenes H Ab|Listeria monocytogenes H Ab
C1545096|T201|COMP|41168-6|LNC|Arginine|Arginine
C1545097|T201|COMP|41169-4|LNC|Valine|Valine
C1545098|T201|COMP|41170-2|LNC|Phenylalanine+Tyrosine|Phenylalanine+Tyrosine
C1545099|T201|COMP|41171-0|LNC|Collagen crosslinked C-telopeptide|Collagen crosslinked C-telopeptide
C1545100|T201|COMP|41172-8|LNC|Yeast.budding|Yeast.budding
C1545101|T201|COMP|41173-6|LNC|Xylose^2H post dose xylose PO|Xylose^2H post dose xylose PO
C1545102|T201|COMP|41174-4|LNC|Waxy casts.broad|Waxy casts.broad
C1545103|T201|COMP|41175-1|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C1545107|T201|COMP|41183-5|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C1545108|T201|COMP|41184-3|LNC|Warfarin|Warfarin
C1545109|T201|COMP|41185-0|LNC|Xylose^5H post dose xylose PO|Xylose^5H post dose xylose PO
C1545110|T201|COMP|41186-8|LNC|Yeast|Yeast
C1545111|T201|COMP|41187-6|LNC|Waxy casts|Waxy casts
C1545112|T201|COMP|41188-4|LNC|Xylose^post CFst|Xylose^post CFst
C1545113|T201|COMP|41189-2|LNC|Xylose^post CFst|Xylose^post CFst
C1545114|T201|COMP|41190-0|LNC|Waxy casts|Waxy casts
C1545115|T201|COMP|41191-8|LNC|Xylose^2H post dose xylose PO|Xylose^2H post dose xylose PO
C1545116|T201|COMP|41192-6|LNC|Dolichovespula arenaria Ab.IgG4|Dolichovespula arenaria Ab.IgG4
C1545117|T201|COMP|41193-4|LNC|Dolichovespula maculata Ab.IgG4|Dolichovespula maculata Ab.IgG4
C1545118|T201|COMP|41194-2|LNC|West Nile virus Ab|West Nile virus Ab
C1545119|T201|COMP|41195-9|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1545120|T201|COMP|41196-7|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C1545121|T201|COMP|41198-3|LNC|Juglans spp Ab.IgE/IgE.total|Juglans spp Ab.IgE/IgE.total
C1545122|T201|COMP|41199-1|LNC|Voriconazole|Voriconazole
C1545123|T201|COMP|41200-7|LNC|Voriconazole|Voriconazole
C1545124|T201|COMP|41201-5|LNC|Voltage-gated calcium channel Ab.IgG|Voltage-gated calcium channel Ab.IgG
C1545125|T201|COMP|41202-3|LNC|Saccharomyces cerevisiae Ab.IgE/IgE.total|Saccharomyces cerevisiae Ab.IgE/IgE.total
C1545126|T201|COMP|41203-1|LNC|Vespula spp Ab.IgE/IgE.total|Vespula spp Ab.IgE/IgE.total
C1545127|T201|COMP|41204-9|LNC|Polistes spp Ab.IgE/IgE.total|Polistes spp Ab.IgE/IgE.total
C1545128|T201|COMP|41205-6|LNC|Citrullus lanatus Ab.IgG|Citrullus lanatus Ab.IgG
C1545129|T201|COMP|41206-4|LNC|West Nile virus Ab|West Nile virus Ab
C1545130|T201|COMP|41207-2|LNC|Triticum aestivum Ab.IgE/IgE.total|Triticum aestivum Ab.IgE/IgE.total
C1545131|T201|COMP|41208-0|LNC|Viscosity+Liquefaction|Viscosity+Liquefaction
C1545132|T201|COMP|41209-8|LNC|VWF gene.p.Arg854Gln|VWF gene.p.Arg854Gln
C1545133|T201|COMP|41210-6|LNC|VWF gene.p.Arg816Trp|VWF gene.p.Arg816Trp
C1545134|T201|COMP|41211-4|LNC|West Nile virus Ab.IgG+IgM|West Nile virus Ab.IgG+IgM
C1545135|T201|COMP|41212-2|LNC|West Nile virus RNA|West Nile virus RNA
C1545136|T201|COMP|41213-0|LNC|Xanthan gum Ab.IgE|Xanthan gum Ab.IgE
C1545137|T201|COMP|41214-8|LNC|Volatiles|Volatiles
C1545138|T201|COMP|41215-5|LNC|Yeast|Yeast
C1545139|T201|COMP|41216-3|LNC|Yellow fever virus Ab.IgM|Yellow fever virus Ab.IgM
C1545140|T201|COMP|41217-1|LNC|Yellow fever virus Ab.IgG|Yellow fever virus Ab.IgG
C1545141|T201|COMP|41218-9|LNC|Xipamid|Xipamid
C1545142|T201|COMP|41219-7|LNC|Polistes spp Ab.IgG|Polistes spp Ab.IgG
C1545143|T201|COMP|41220-5|LNC|Xanthurenate|Xanthurenate
C1545144|T201|COMP|41221-3|LNC|Xanthurenate+Kynurenate|Xanthurenate+Kynurenate
C1545145|T201|COMP|41222-1|LNC|Yeast|Yeast
C1545146|T201|COMP|41223-9|LNC|Waxy casts|Waxy casts
C1545147|T201|COMP|41224-7|LNC|West Nile virus Ab|West Nile virus Ab
C1545148|T201|COMP|41225-4|LNC|West Nile virus Ab|West Nile virus Ab
C1545149|T201|COMP|41226-2|LNC|Viscosity|Viscosity
C1545150|T201|COMP|41227-0|LNC|Xanthine|Xanthine
C1545151|T201|COMP|41228-8|LNC|Xanthine|Xanthine
C1545152|T201|COMP|41229-6|LNC|Vespula spp Ab.IgG|Vespula spp Ab.IgG
C1545153|T201|COMP|41230-4|LNC|Xanthine|Xanthine
C1545154|T201|COMP|41231-2|LNC|Xanthurenate+Kynurenate|Xanthurenate+Kynurenate
C1545155|T201|COMP|41232-0|LNC|West Nile virus Ab|West Nile virus Ab
C1545158|T201|COMP|41235-3|LNC|Polistes spp Ab.IgE|Polistes spp Ab.IgE
C1545159|T201|COMP|41236-1|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C1545160|T201|COMP|41237-9|LNC|Xylose^5H post dose xylose PO|Xylose^5H post dose xylose PO
C1545161|T201|COMP|41238-7|LNC|Viscosity|Viscosity
C1545162|T201|COMP|41239-5|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C1545163|T201|COMP|41240-3|LNC|Xanthurenate|Xanthurenate
C1545164|T201|COMP|41241-1|LNC|Viscosity|Viscosity
C1545165|T201|COMP|41242-9|LNC|Yeast|Yeast
C1545166|T201|COMP|41243-7|LNC|Yeast|Yeast
C1545167|T201|COMP|41244-5|LNC|Western equine encephalitis virus Ab.IgG|Western equine encephalitis virus Ab.IgG
C1545168|T201|COMP|41245-2|LNC|Viscosity|Viscosity
C1545169|T201|COMP|41246-0|LNC|Yellow fever virus Ab^2nd specimen|Yellow fever virus Ab^2nd specimen
C1545170|T201|COMP|41247-8|LNC|Yellow fever virus Ab^1st specimen|Yellow fever virus Ab^1st specimen
C1545171|T201|COMP|41248-6|LNC|Xanthurenate|Xanthurenate
C1545172|T201|COMP|41249-4|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C1545173|T201|COMP|41250-2|LNC|Xylose^baseline|Xylose^baseline
C1545174|T201|COMP|41251-0|LNC|Xylose^5H post 25 g xylose PO|Xylose^5H post 25 g xylose PO
C1545175|T201|COMP|41252-8|LNC|Xylose^5H post 25 g xylose PO|Xylose^5H post 25 g xylose PO
C1545176|T201|COMP|41253-6|LNC|Xylose^4H post 25 g xylose PO|Xylose^4H post 25 g xylose PO
C1545177|T201|COMP|41254-4|LNC|Xylose^4H post 25 g xylose PO|Xylose^4H post 25 g xylose PO
C1545178|T201|COMP|41255-1|LNC|Xylose^3H post 25 g xylose PO|Xylose^3H post 25 g xylose PO
C1545179|T201|COMP|41256-9|LNC|Xylose^3H post 25 g xylose PO|Xylose^3H post 25 g xylose PO
C1545180|T201|COMP|41257-7|LNC|Xylose^2H post 25 g xylose PO|Xylose^2H post 25 g xylose PO
C1545181|T201|COMP|41258-5|LNC|Xylose^1H post 25 g xylose PO|Xylose^1H post 25 g xylose PO
C1545182|T201|COMP|41259-3|LNC|Western equine encephalitis virus Ab.IgM|Western equine encephalitis virus Ab.IgM
C1545183|T201|COMP|41260-1|LNC|Western equine encephalitis virus Ab.IgG|Western equine encephalitis virus Ab.IgG
C1545184|T201|COMP|41261-9|LNC|Voltage-gated calcium channel Ab.IgG|Voltage-gated calcium channel Ab.IgG
C1545185|T201|COMP|41262-7|LNC|Viscosity|Viscosity
C1545186|T201|COMP|41263-5|LNC|Viscosity|Viscosity
C1545187|T201|COMP|41264-3|LNC|Viscosity|Viscosity
C1545188|T201|COMP|41265-0|LNC|Width|Width
C1545189|T201|COMP|41266-8|LNC|Volatiles|Volatiles
C1545190|T201|COMP|41267-6|LNC|Xylose^post dose xylose PO|Xylose^post dose xylose PO
C1545191|T201|COMP|41268-4|LNC|VWF gene.p.Thr791Met|VWF gene.p.Thr791Met
C1545192|T201|COMP|41269-2|LNC|Beta hydroxybutyrate+Gamma aminobutyrate|Beta hydroxybutyrate+Gamma aminobutyrate
C1545193|T201|COMP|41270-0|LNC|Drugs identified|Drugs identified
C1545194|T201|COMP|41271-8|LNC|Dermatophagoides sp Ab.IgE|Dermatophagoides sp Ab.IgE
C1545195|T201|COMP|41272-6|LNC|Dog dander+Dog epithelium Ab.IgE.RAST class|Dog dander+Dog epithelium Ab.IgE.RAST class
C1545196|T201|COMP|41273-4|LNC|Alpha-1-Fetoprotein interpretation|Alpha-1-Fetoprotein interpretation
C1545197|T201|COMP|41274-2|LNC|Alpha-1-Fetoprotein interpretation|Alpha-1-Fetoprotein interpretation
C1545198|T201|COMP|41275-9|LNC|Amino acids intense band position|Amino acids intense band position
C1545199|T201|COMP|41276-7|LNC|Anion gap|Anion gap
C1545200|T201|COMP|41277-5|LNC|Gross blood|Gross blood
C1545201|T201|COMP|41278-3|LNC|Gross blood|Gross blood
C1545203|T201|COMP|41280-9|LNC|Appearance|Appearance
C1545204|T201|COMP|41281-7|LNC|Burr cells|Burr cells
C1545205|T201|COMP|41282-5|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C1545206|T201|COMP|41283-3|LNC|HLA-DQ8|HLA-DQ8
C1545207|T201|COMP|41284-1|LNC|Epithelial cells.non-squamous|Epithelial cells.non-squamous
C1545208|T201|COMP|41285-8|LNC|Uranium.depleted/Creatinine|Uranium.depleted/Creatinine
C1545209|T201|COMP|41286-6|LNC|Uranium 235/Uranium 238|Uranium 235/Uranium 238
C1545210|T201|COMP|41287-4|LNC|Epithelial cells.parabasal|Epithelial cells.parabasal
C1545211|T201|COMP|41288-2|LNC|Egg whole Ab.IgE/IgE.total|Egg whole Ab.IgE/IgE.total
C1545212|T201|COMP|41289-0|LNC|11-Deoxycortisol^post dose metyraPONE|11-Deoxycortisol^post dose metyraPONE
C1546313|T201|COMP|40253-7|LNC|Creatinine^2.25H post XXX challenge|Creatinine^2.25H post XXX challenge
C1546339|T201|COMP|41084-5|LNC|MSH2 gene targeted mutation analysis|MSH2 gene targeted mutation analysis
C1546340|T201|COMP|41082-9|LNC|MT-TK gene targeted mutation analysis|MT-TK gene targeted mutation analysis
C1546342|T201|COMP|40568-8|LNC|Metamyelocytes|Metamyelocytes
C1546343|T201|COMP|41179-3|LNC|Mumps reaction wheal^1D post mumps ID|Mumps reaction wheal^1D post mumps ID
C1546344|T201|COMP|41178-5|LNC|Mumps reaction wheal^2D post dose mumps ID|Mumps reaction wheal^2D post dose mumps ID
C1621247|T201|COMP|42961-3|LNC|Salmonella pullorum Ab|Salmonella pullorum Ab
C1621808|T201|COMP|42506-6|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C1622349|T201|COMP|42773-2|LNC|Multiple drug resistant organism identified|Multiple drug resistant organism identified
C1623566|T201|COMP|41992-9|LNC|Arsenic.inorganic|Arsenic.inorganic
C1623567|T201|COMP|41993-7|LNC|Atazanavir|Atazanavir
C1623568|T201|COMP|41994-5|LNC|Cells.CD4+CD45RO+/100 cells|Cells.CD4+CD45RO+/100 cells
C1623569|T201|COMP|41996-0|LNC|Hepatitis C virus DNA|Hepatitis C virus DNA
C1623570|T201|COMP|41999-4|LNC|Lipoprotein.pre-beta|Lipoprotein.pre-beta
C1623571|T201|COMP|42000-0|LNC|Lopinavir+Ritonavir|Lopinavir+Ritonavir
C1623572|T201|COMP|42001-8|LNC|Nickel/Creatinine|Nickel/Creatinine
C1623573|T201|COMP|42003-4|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1623583|T201|COMP|43101-5|LNC|Phosphatidylserine Ab.IgA & IgG & IgM panel|Phosphatidylserine Ab.IgA & IgG & IgM panel
C1623584|T201|COMP|43105-6|LNC|Acetaldehyde & Paraldehyde panel|Acetaldehyde & Paraldehyde panel
C1623585|T201|COMP|43111-4|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C1623586|T201|COMP|43123-9|LNC|Imipramine & Desipramine panel|Imipramine & Desipramine panel
C1623587|T201|COMP|43127-0|LNC|Clomipramine & Norclomipramine panel|Clomipramine & Norclomipramine panel
C1623593|T201|COMP|43154-4|LNC|Spermatozoa^post concentration|Spermatozoa^post concentration
C1623595|T201|COMP|42672-6|LNC|Debris|Debris
C1623600|T201|COMP|42719-5|LNC|Bilirubin|Bilirubin
C1623601|T201|COMP|42724-5|LNC|OmpC Ab|OmpC Ab
C1623602|T201|COMP|42729-4|LNC|Cardiolipin Ab.IgA.B2GP1 dependent|Cardiolipin Ab.IgA.B2GP1 dependent
C1623603|T201|COMP|42732-8|LNC|Cardiolipin Ab.IgG.B2GP1 independent|Cardiolipin Ab.IgG.B2GP1 independent
C1623604|T201|COMP|42735-1|LNC|Cells.CD20+CD117+/100 cells|Cells.CD20+CD117+/100 cells
C1623605|T201|COMP|42739-3|LNC|Phosphatidylcholine Ab.IgA.B2GP1 dependent|Phosphatidylcholine Ab.IgA.B2GP1 dependent
C1623606|T201|COMP|42746-8|LNC|Phosphatidylethanolamine Ab.IgA.B2GP1 independent|Phosphatidylethanolamine Ab.IgA.B2GP1 independent
C1623607|T201|COMP|42747-6|LNC|Phosphatidylethanolamine Ab.IgG.B2GP1 dependent|Phosphatidylethanolamine Ab.IgG.B2GP1 dependent
C1623608|T201|COMP|42750-0|LNC|Phosphatidylethanolamine Ab.IgM.B2GP1 independent|Phosphatidylethanolamine Ab.IgM.B2GP1 independent
C1623609|T201|COMP|42753-4|LNC|Phosphatidylserine Ab.IgG.B2GP1 dependent|Phosphatidylserine Ab.IgG.B2GP1 dependent
C1623610|T201|COMP|42760-9|LNC|Inflammatory bowel disease Ab panel|Inflammatory bowel disease Ab panel
C1623611|T201|COMP|42770-8|LNC|Human papilloma virus high & Low risk DNA panel|Human papilloma virus high & Low risk DNA panel
C1623612|T201|COMP|42775-7|LNC|Multiple drug resistant organism identified|Multiple drug resistant organism identified
C1623613|T201|COMP|42929-0|LNC|Lactate dehydrogenase panel|Lactate dehydrogenase panel
C1623614|T201|COMP|42941-5|LNC|GALT gene allele 2|GALT gene allele 2
C1623615|T201|COMP|42944-9|LNC|Vesicular stomatitis New Jersey virus Ab|Vesicular stomatitis New Jersey virus Ab
C1623616|T201|COMP|42979-5|LNC|Polio virus 3 Ab|Polio virus 3 Ab
C1623617|T201|COMP|42982-9|LNC|Parainfluenza virus Ab|Parainfluenza virus Ab
C1623618|T201|COMP|43000-9|LNC|Leishmania braziliensis Ab|Leishmania braziliensis Ab
C1623619|T201|COMP|43002-5|LNC|Legionella pneumophila 1 Ab.IgM|Legionella pneumophila 1 Ab.IgM
C1623620|T201|COMP|43005-8|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C1623621|T201|COMP|43009-0|LNC|HIV 1+2 Ab.IgG|HIV 1+2 Ab.IgG
C1623622|T201|COMP|43022-3|LNC|Herpes virus 7 Ab.IgM|Herpes virus 7 Ab.IgM
C1623623|T201|COMP|43023-1|LNC|Herpes virus 7 Ab.IgG|Herpes virus 7 Ab.IgG
C1624104|T201|COMP|41995-2|LNC|Hemoglobin A1c|Hemoglobin A1c
C1624105|T201|COMP|41997-8|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C1624106|T201|COMP|42004-2|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C1624107|T201|COMP|42006-7|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C1624115|T201|COMP|43099-1|LNC|Vanillylmandelate & Creatinine panel|Vanillylmandelate & Creatinine panel
C1624116|T201|COMP|43102-3|LNC|Neuronal nuclear type 3 Ab|Neuronal nuclear type 3 Ab
C1624117|T201|COMP|43103-1|LNC|CV2 Ab.IgG|CV2 Ab.IgG
C1624118|T201|COMP|43110-6|LNC|Immunoglobulin light chains panel|Immunoglobulin light chains panel
C1624119|T201|COMP|43113-0|LNC|Hemoglobin panel|Hemoglobin panel
C1624120|T201|COMP|43114-8|LNC|Porphyrin fractions|Porphyrin fractions
C1624121|T201|COMP|43130-4|LNC|Bile acid fractions panel|Bile acid fractions panel
C1624122|T201|COMP|43132-0|LNC|California encephalitis virus Ab|California encephalitis virus Ab
C1624125|T201|COMP|42673-4|LNC|Calcium hydrogen phosphate dihydrate|Calcium hydrogen phosphate dihydrate
C1624126|T201|COMP|42676-7|LNC|Spermatozoa.normal.motile|Spermatozoa.normal.motile
C1624127|T201|COMP|42678-3|LNC|Urate|Urate
C1624136|T201|COMP|42712-0|LNC|AML+MDS gene 7q31 deletion|AML+MDS gene 7q31 deletion
C1624137|T201|COMP|42713-8|LNC|AML+MDS gene CEP 8 trisomy|AML+MDS gene CEP 8 trisomy
C1624139|T201|COMP|42720-3|LNC|Clindamycin.induced|Clindamycin.induced
C1624140|T201|COMP|42726-0|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C1624141|T201|COMP|42730-2|LNC|Cardiolipin Ab.IgA.B2GP1 independent|Cardiolipin Ab.IgA.B2GP1 independent
C1624142|T201|COMP|42738-5|LNC|Cells.CD7+CD8+/100 cells|Cells.CD7+CD8+/100 cells
C1624143|T201|COMP|42742-7|LNC|Phosphatidylcholine Ab.IgG.B2GP1 independent|Phosphatidylcholine Ab.IgG.B2GP1 independent
C1624144|T201|COMP|42744-3|LNC|Phosphatidylcholine Ab.IgM.B2GP1 independent|Phosphatidylcholine Ab.IgM.B2GP1 independent
C1624145|T201|COMP|42748-4|LNC|Phosphatidylethanolamine Ab.IgG.B2GP1 independent|Phosphatidylethanolamine Ab.IgG.B2GP1 independent
C1624146|T201|COMP|42759-1|LNC|Lymphocytes B|Lymphocytes B
C1624147|T201|COMP|42768-2|LNC|HIV 1 & 2 Ab|HIV 1 & 2 Ab
C1624148|T201|COMP|42772-4|LNC|Fibrinogen Ag|Fibrinogen Ag
C1624149|T201|COMP|42779-9|LNC|BRCA2 Ag|BRCA2 Ag
C1624151|T201|COMP|42783-1|LNC|ERBB2 gene targeted mutation analysis|ERBB2 gene targeted mutation analysis
C1624153|T201|COMP|42787-2|LNC|HER4 Ag|HER4 Ag
C1624154|T201|COMP|42791-4|LNC|Mitogen-Activated protein kinase 3 Ag|Mitogen-Activated protein kinase 3 Ag
C1624155|T201|COMP|42794-8|LNC|MYC gene targeted mutation analysis|MYC gene targeted mutation analysis
C1624156|T201|COMP|42921-7|LNC|JC virus DNA|JC virus DNA
C1624157|T201|COMP|42925-8|LNC|Myeloid cells/100 cells|Myeloid cells/100 cells
C1624158|T201|COMP|42930-8|LNC|Cells.CD11+CD18+|Cells.CD11+CD18+
C1624159|T201|COMP|42942-3|LNC|Yersinia sp Ab.IgM|Yersinia sp Ab.IgM
C1624160|T201|COMP|42943-1|LNC|Yersinia enterocolitica O:5,27 Ab|Yersinia enterocolitica O:5,27 Ab
C1624161|T201|COMP|42945-6|LNC|Vesicular stomatitis Indiana virus Ab|Vesicular stomatitis Indiana virus Ab
C1624162|T201|COMP|42946-4|LNC|Trypanosoma brucei rhodesiense Ab|Trypanosoma brucei rhodesiense Ab
C1624163|T201|COMP|42948-0|LNC|Toxoplasma sp Ab.IgM|Toxoplasma sp Ab.IgM
C1624164|T201|COMP|42949-8|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C1624165|T201|COMP|42960-5|LNC|Salmonella typhi H Ab|Salmonella typhi H Ab
C1624167|T201|COMP|42984-5|LNC|Parainfluenza virus 1 Ab^2nd specimen|Parainfluenza virus 1 Ab^2nd specimen
C1624168|T201|COMP|42987-8|LNC|Neisseria gonorrhoeae Ab|Neisseria gonorrhoeae Ab
C1624169|T201|COMP|43010-8|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C1624170|T201|COMP|43011-6|LNC|HIV 1 p24 Ab|HIV 1 p24 Ab
C1624171|T201|COMP|43012-4|LNC|HIV 1 gp41 Ab|HIV 1 gp41 Ab
C1624172|T201|COMP|43019-9|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C1624663|T201|COMP|42002-6|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C1624664|T201|COMP|42005-9|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C1624676|T201|COMP|43104-9|LNC|Paraneoplastic Ab panel|Paraneoplastic Ab panel
C1624677|T201|COMP|43115-5|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C1624678|T201|COMP|43117-1|LNC|Fluoxetine & Norfluoxetine panel|Fluoxetine & Norfluoxetine panel
C1624679|T201|COMP|43120-5|LNC|Echovirus Ab panel|Echovirus Ab panel
C1624680|T201|COMP|43121-3|LNC|Echovirus 6 Ab|Echovirus 6 Ab
C1624681|T201|COMP|43122-1|LNC|Doxepin & Nordoxepin panel|Doxepin & Nordoxepin panel
C1624682|T201|COMP|43124-7|LNC|Cystine panel|Cystine panel
C1624683|T201|COMP|43125-4|LNC|Nicotine & Metabolites panel|Nicotine & Metabolites panel
C1624684|T201|COMP|43126-2|LNC|Cortisol.free panel|Cortisol.free panel
C1624685|T201|COMP|43128-8|LNC|Chloride panel|Chloride panel
C1624686|T201|COMP|43129-6|LNC|Brucella abortus Ab.IgG & IgM panel|Brucella abortus Ab.IgG & IgM panel
C1624687|T201|COMP|43134-6|LNC|Calcidiol & Calciferol & Calcitriol panel|Calcidiol & Calciferol & Calcitriol panel
C1624693|T201|COMP|42671-8|LNC|Serotonin|Serotonin
C1624694|T201|COMP|42677-5|LNC|Succinylacetone|Succinylacetone
C1624695|T201|COMP|42679-1|LNC|Heparin|Heparin
C1624701|T201|COMP|42715-3|LNC|Del(5)(q12-35) gene deletion|Del(5)(q12-35) gene deletion
C1624702|T201|COMP|42716-1|LNC|Mycobacterium sp rRNA|Mycobacterium sp rRNA
C1624703|T201|COMP|42717-9|LNC|Mycobacterium tuberculosis complex genotype|Mycobacterium tuberculosis complex genotype
C1624705|T201|COMP|42721-1|LNC|Staphylococcus sp.oxacillin resistant isolate|Staphylococcus sp.oxacillin resistant isolate
C1624706|T201|COMP|42727-8|LNC|Fibrin D-dimer DDU|Fibrin D-dimer DDU
C1624707|T201|COMP|42734-4|LNC|Cardiolipin Ab.IgM.B2GP1 independent|Cardiolipin Ab.IgM.B2GP1 independent
C1624708|T201|COMP|42737-7|LNC|Cells.CD4+CD7+/100 cells|Cells.CD4+CD7+/100 cells
C1624709|T201|COMP|42741-9|LNC|Phosphatidylcholine Ab.IgG.B2GP1 dependent|Phosphatidylcholine Ab.IgG.B2GP1 dependent
C1624710|T201|COMP|42743-5|LNC|Phosphatidylcholine Ab.IgM.B2GP1 dependent|Phosphatidylcholine Ab.IgM.B2GP1 dependent
C1624711|T201|COMP|42754-2|LNC|Phosphatidylserine Ab.IgG.B2GP1 independent|Phosphatidylserine Ab.IgG.B2GP1 independent
C1624712|T201|COMP|42755-9|LNC|Phosphatidylserine Ab.IgM.B2GP1 dependent|Phosphatidylserine Ab.IgM.B2GP1 dependent
C1624713|T201|COMP|42756-7|LNC|Phosphatidylserine Ab.IgM.B2GP1 independent|Phosphatidylserine Ab.IgM.B2GP1 independent
C1624714|T201|COMP|42758-3|LNC|Reticulocytes|Reticulocytes
C1624715|T201|COMP|42766-6|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C1624716|T201|COMP|42769-0|LNC|HTLV I+II Ab|HTLV I+II Ab
C1624717|T201|COMP|42771-6|LNC|Streptococcus pneumoniae serotype Ab.IgG|Streptococcus pneumoniae serotype Ab.IgG
C1624718|T201|COMP|42774-0|LNC|Multiple drug resistant organism identified|Multiple drug resistant organism identified
C1624719|T201|COMP|42923-3|LNC|Kochia scoparia Ab.IgE/IgE.total|Kochia scoparia Ab.IgE/IgE.total
C1624720|T201|COMP|42926-6|LNC|Myeloid cells/100 cells|Myeloid cells/100 cells
C1624721|T201|COMP|42947-2|LNC|Trypanosoma brucei Ab|Trypanosoma brucei Ab
C1624722|T201|COMP|42980-3|LNC|Polio virus Ab|Polio virus Ab
C1624723|T201|COMP|42985-2|LNC|Neisseria meningitidis serogroup C Ab.IgG|Neisseria meningitidis serogroup C Ab.IgG
C1624724|T201|COMP|43006-6|LNC|Jamestown canyon virus Ab|Jamestown canyon virus Ab
C1624725|T201|COMP|43007-4|LNC|HTLV I+II Ab|HTLV I+II Ab
C1624726|T201|COMP|43008-2|LNC|HIV 1+2 Ab.IgM|HIV 1+2 Ab.IgM
C1624727|T201|COMP|43017-3|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C1624728|T201|COMP|43020-7|LNC|Heterophile Ab|Heterophile Ab
C1625198|T201|COMP|41998-6|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C1625207|T201|COMP|43106-4|LNC|Amitriptyline & Nortriptyline panel|Amitriptyline & Nortriptyline panel
C1625208|T201|COMP|43107-2|LNC|Mycoplasma sp & Ureaplasma sp panel|Mycoplasma sp & Ureaplasma sp panel
C1625209|T201|COMP|43108-0|LNC|Metanephrine & Normetanephrine panel|Metanephrine & Normetanephrine panel
C1625210|T201|COMP|43116-3|LNC|Porphyrin fractions panel|Porphyrin fractions panel
C1625211|T201|COMP|43118-9|LNC|Fat panel|Fat panel
C1625212|T201|COMP|43119-7|LNC|Extractable nuclear Ab panel|Extractable nuclear Ab panel
C1625215|T201|COMP|42674-2|LNC|Fat.neutral|Fat.neutral
C1625216|T201|COMP|42682-5|LNC|Succinyladenosine|Succinyladenosine
C1625221|T201|COMP|42733-6|LNC|Cardiolipin Ab.IgM.B2GP1 dependent|Cardiolipin Ab.IgM.B2GP1 dependent
C1625222|T201|COMP|42736-9|LNC|Cells.CD20+CD23+/100 cells|Cells.CD20+CD23+/100 cells
C1625223|T201|COMP|42745-0|LNC|Phosphatidylethanolamine Ab.IgA.B2GP1 dependent|Phosphatidylethanolamine Ab.IgA.B2GP1 dependent
C1625224|T201|COMP|42749-2|LNC|Phosphatidylethanolamine Ab.IgM.B2GP1 dependent|Phosphatidylethanolamine Ab.IgM.B2GP1 dependent
C1625225|T201|COMP|42752-6|LNC|Phosphatidylserine Ab.IgA.B2GP1 independent|Phosphatidylserine Ab.IgA.B2GP1 independent
C1625226|T201|COMP|42764-1|LNC|Crystals|Crystals
C1625227|T201|COMP|42767-4|LNC|Borrelia burgdorferi Ab.IgG & IgM|Borrelia burgdorferi Ab.IgG & IgM
C1625229|T201|COMP|42780-7|LNC|CCND1 gene targeted mutation analysis|CCND1 gene targeted mutation analysis
C1625231|T201|COMP|42786-4|LNC|HER3 Ag|HER3 Ag
C1625232|T201|COMP|42788-0|LNC|Insulin-like growth factor-I receptor Ag|Insulin-like growth factor-I receptor Ag
C1625233|T201|COMP|42789-8|LNC|Mitogen-Activated protein kinase 14 Ag|Mitogen-Activated protein kinase 14 Ag
C1625234|T201|COMP|42792-2|LNC|Mitogen-Activated protein kinase 8 Ag|Mitogen-Activated protein kinase 8 Ag
C1625235|T201|COMP|42793-0|LNC|Mitogen-Activated protein kinase 9 Ag|Mitogen-Activated protein kinase 9 Ag
C1625236|T201|COMP|42795-5|LNC|Retinoblastoma protein|Retinoblastoma protein
C1625238|T201|COMP|42924-1|LNC|Lactoferrin|Lactoferrin
C1625239|T201|COMP|42927-4|LNC|Myeloid cells/100 cells|Myeloid cells/100 cells
C1625240|T201|COMP|42928-2|LNC|Filaria Ag|Filaria Ag
C1625241|T201|COMP|42978-7|LNC|Polio virus 2 Ab|Polio virus 2 Ab
C1625242|T201|COMP|42983-7|LNC|Parainfluenza virus 4 Ab.IgG|Parainfluenza virus 4 Ab.IgG
C1625243|T201|COMP|42986-0|LNC|Neisseria meningitidis serogroup A Ab.IgG|Neisseria meningitidis serogroup A Ab.IgG
C1625244|T201|COMP|43001-7|LNC|Legionella sp Ab|Legionella sp Ab
C1625245|T201|COMP|43003-3|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C1625246|T201|COMP|43004-1|LNC|Jamestown canyon virus Ab.IgG|Jamestown canyon virus Ab.IgG
C1625247|T201|COMP|43014-0|LNC|Histoplasma sp Ab|Histoplasma sp Ab
C1625248|T201|COMP|43015-7|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C1625249|T201|COMP|43021-5|LNC|Herpes virus 8 Ab.IgG|Herpes virus 8 Ab.IgG
C1625665|T201|COMP|43160-1|LNC|Glutaraldehyde|Glutaraldehyde
C1625666|T201|COMP|43162-7|LNC|Monochloramine|Monochloramine
C1625667|T201|COMP|43169-2|LNC|Bromide|Bromide
C1625668|T201|COMP|42801-1|LNC|Histology grade|Histology grade
C1625751|T201|COMP|43159-3|LNC|Formaldehyde|Formaldehyde
C1625752|T201|COMP|43164-3|LNC|Silica|Silica
C1625753|T201|COMP|43165-0|LNC|Dissolved solids|Dissolved solids
C1625754|T201|COMP|42802-9|LNC|Age at menopause|Age at menopause
C1625755|T201|COMP|42805-2|LNC|Fungus identified|Fungus identified
C1625756|T201|COMP|42806-0|LNC|Bacteria identified|Bacteria identified
C1625757|T201|COMP|42815-1|LNC|Stachybotrys chartarum Ab.IgE|Stachybotrys chartarum Ab.IgE
C1625763|T201|COMP|42856-5|LNC|Benzoylecgonine|Benzoylecgonine
C1625764|T201|COMP|43030-6|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1625765|T201|COMP|43031-4|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C1625766|T201|COMP|43033-0|LNC|Herpes simplex virus 1+2 Ab|Herpes simplex virus 1+2 Ab
C1625767|T201|COMP|43034-8|LNC|Feline leukemia virus Ab|Feline leukemia virus Ab
C1625768|T201|COMP|43045-4|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C1625769|T201|COMP|43051-2|LNC|Colorado tick fever virus Ab.IgG|Colorado tick fever virus Ab.IgG
C1625770|T201|COMP|43053-8|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C1625771|T201|COMP|43055-3|LNC|Clostridioides difficile toxin Ab|Clostridioides difficile toxin Ab
C1625772|T201|COMP|43063-7|LNC|Chlamydia sp Ab.IgA|Chlamydia sp Ab.IgA
C1625793|T201|COMP|42539-7|LNC|Hydroxyperhexiline/Perhexiline|Hydroxyperhexiline/Perhexiline
C1625794|T201|COMP|41623-0|LNC|Bacillus anthracis DNA|Bacillus anthracis DNA
C1626179|T201|COMP|42180-0|LNC|C peptide^post CFst|C peptide^post CFst
C1626180|T201|COMP|42183-4|LNC|Gossypol.negative isomer|Gossypol.negative isomer
C1626181|T201|COMP|42186-7|LNC|Number of specimens received|Number of specimens received
C1626182|T201|COMP|42188-3|LNC|Cells.CD3+CD16+CD56+|Cells.CD3+CD16+CD56+
C1626183|T201|COMP|42189-1|LNC|Cells.CD3+CD16+CD56+/100 cells|Cells.CD3+CD16+CD56+/100 cells
C1626184|T201|COMP|42198-2|LNC|Curvularia specifera Ab.IgE|Curvularia specifera Ab.IgE
C1626185|T201|COMP|42200-6|LNC|DNA double strand Ab|DNA double strand Ab
C1626187|T201|COMP|42870-6|LNC|Cells.CD138/100 cells|Cells.CD138/100 cells
C1626188|T201|COMP|42882-1|LNC|Cells.CD3-CD57+/100 cells|Cells.CD3-CD57+/100 cells
C1626189|T201|COMP|42886-2|LNC|Cells.CD52/100 cells|Cells.CD52/100 cells
C1626190|T201|COMP|42889-6|LNC|Cells.CD79b/100 cells|Cells.CD79b/100 cells
C1626191|T201|COMP|42897-9|LNC|Coxiella burnetii phase 1 Ab.IgM|Coxiella burnetii phase 1 Ab.IgM
C1626192|T201|COMP|42899-5|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C1626193|T201|COMP|42904-3|LNC|Epicoccum purpurascens Ab.IgG|Epicoccum purpurascens Ab.IgG
C1626272|T201|COMP|43158-5|LNC|Chlorine.free|Chlorine.free
C1626273|T201|COMP|43161-9|LNC|Microorganism|Microorganism
C1626274|T201|COMP|43166-8|LNC|Carbon.organic|Carbon.organic
C1626275|T201|COMP|42797-1|LNC|Age at first pregnancy|Age at first pregnancy
C1626276|T201|COMP|42798-9|LNC|Age at menarche|Age at menarche
C1626279|T201|COMP|42803-7|LNC|Bacteria identified|Bacteria identified
C1626280|T201|COMP|42807-8|LNC|Parasite identified|Parasite identified
C1626281|T201|COMP|42808-6|LNC|Virus identified|Virus identified
C1626283|T201|COMP|42818-5|LNC|Cells.CD38+Lambda+/100 cells|Cells.CD38+Lambda+/100 cells
C1626287|T201|COMP|42855-7|LNC|11-Deoxycorticosterone|11-Deoxycorticosterone
C1626288|T201|COMP|42859-9|LNC|Candida albicans Ab|Candida albicans Ab
C1626289|T201|COMP|43027-2|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C1626290|T201|COMP|43029-8|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C1626291|T201|COMP|43037-1|LNC|Fasciola hepatica Ab|Fasciola hepatica Ab
C1626292|T201|COMP|43040-5|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C1626293|T201|COMP|43048-8|LNC|Coxsackievirus A9 Ab|Coxsackievirus A9 Ab
C1626294|T201|COMP|43049-6|LNC|Coxsackievirus A10 Ab|Coxsackievirus A10 Ab
C1626295|T201|COMP|43050-4|LNC|Coxiella burnetii phase 1 Ab|Coxiella burnetii phase 1 Ab
C1626296|T201|COMP|43056-1|LNC|Cladosporium sp Ab.IgG|Cladosporium sp Ab.IgG
C1626297|T201|COMP|43058-7|LNC|Chlamydia trachomatis D+K Ab.IgM|Chlamydia trachomatis D+K Ab.IgM
C1626298|T201|COMP|43066-0|LNC|Canine distemper virus Ab.IgG|Canine distemper virus Ab.IgG
C1626321|T201|COMP|41434-2|LNC|Cryptosporidium parvum DNA|Cryptosporidium parvum DNA
C1626323|T201|COMP|42533-0|LNC|Saccharomonospora viridis Ab|Saccharomonospora viridis Ab
C1626324|T201|COMP|41511-7|LNC|Trichomonas vaginalis Ag|Trichomonas vaginalis Ag
C1626771|T201|COMP|42178-4|LNC|Lipoprotein.X|Lipoprotein.X
C1626772|T201|COMP|42185-9|LNC|Number of specimens obtained|Number of specimens obtained
C1626773|T201|COMP|42190-9|LNC|Shigella sp DNA|Shigella sp DNA
C1626810|T201|COMP|42860-7|LNC|Cannabinoids|Cannabinoids
C1626811|T201|COMP|43024-9|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C1626812|T201|COMP|43025-6|LNC|Herpes virus 6 Ab.IgM|Herpes virus 6 Ab.IgM
C1626813|T201|COMP|43026-4|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C1626814|T201|COMP|43028-0|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C1626815|T201|COMP|43038-9|LNC|Enterovirus NOS Ab|Enterovirus NOS Ab
C1626816|T201|COMP|43039-7|LNC|Ehrlichia sp Ab|Ehrlichia sp Ab
C1626817|T201|COMP|43043-9|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C1626818|T201|COMP|43046-2|LNC|Coxsackievirus A16 Ab|Coxsackievirus A16 Ab
C1626819|T201|COMP|43059-5|LNC|Chlamydia trachomatis D+K Ab.IgG|Chlamydia trachomatis D+K Ab.IgG
C1626820|T201|COMP|43060-3|LNC|Chlamydia trachomatis D+K Ab.IgA|Chlamydia trachomatis D+K Ab.IgA
C1626821|T201|COMP|43061-1|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C1626822|T201|COMP|43062-9|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C1626823|T201|COMP|43065-2|LNC|Canine distemper virus Ab.IgM|Canine distemper virus Ab.IgM
C1626824|T201|COMP|43068-6|LNC|Campylobacter sp Ab.IgA|Campylobacter sp Ab.IgA
C1626825|T201|COMP|43069-4|LNC|Burkholderia pseudomallei Ab.IgM|Burkholderia pseudomallei Ab.IgM
C1626842|T201|COMP|42988-6|LNC|Mycoplasma synoviae Ab|Mycoplasma synoviae Ab
C1626844|T201|COMP|41445-8|LNC|Ova+Parasites identified|Ova+Parasites identified
C1626845|T201|COMP|41484-7|LNC|Coxsackievirus A Ab panel|Coxsackievirus A Ab panel
C1626846|T201|COMP|41507-5|LNC|Rabies virus Ab|Rabies virus Ab
C1627302|T201|COMP|42176-8|LNC|1,3 beta glucan|1,3 beta glucan
C1627303|T201|COMP|42187-5|LNC|Number of specimens tested|Number of specimens tested
C1627304|T201|COMP|42193-3|LNC|Cells.CD3/100 cells|Cells.CD3/100 cells
C1627305|T201|COMP|42196-6|LNC|Centromere Ab|Centromere Ab
C1627306|T201|COMP|42203-0|LNC|Ganglioside GM1 Ab|Ganglioside GM1 Ab
C1627308|T201|COMP|42219-6|LNC|Chromium|Chromium
C1627309|T201|COMP|42866-4|LNC|Cells.CD117/100 cells|Cells.CD117/100 cells
C1627310|T201|COMP|42867-2|LNC|Cells.CD117/100 cells|Cells.CD117/100 cells
C1627311|T201|COMP|42869-8|LNC|Cells.CD138/100 cells|Cells.CD138/100 cells
C1627312|T201|COMP|42874-8|LNC|Cells.CD18/100 cells|Cells.CD18/100 cells
C1627313|T201|COMP|42891-2|LNC|Choriogonadotropin|Choriogonadotropin
C1627314|T201|COMP|42902-7|LNC|Elastase.pancreatic|Elastase.pancreatic
C1627315|T201|COMP|42903-5|LNC|Enterovirus NOS Ab|Enterovirus NOS Ab
C1627316|T201|COMP|42905-0|LNC|Formate/Creatinine|Formate/Creatinine
C1627317|T201|COMP|42910-0|LNC|Hemoglobin.gastrointestinal^2nd specimen|Hemoglobin.gastrointestinal^2nd specimen
C1627318|T201|COMP|42911-8|LNC|Hemoglobin.gastrointestinal^3rd specimen|Hemoglobin.gastrointestinal^3rd specimen
C1627319|T201|COMP|42912-6|LNC|Hemoglobin.gastrointestinal^2nd specimen|Hemoglobin.gastrointestinal^2nd specimen
C1627320|T201|COMP|42919-1|LNC|Insulin^pre 100 g glucose PO|Insulin^pre 100 g glucose PO
C1627321|T201|COMP|42920-9|LNC|Isovalerylcarnitine (C5)|Isovalerylcarnitine (C5)
C1627322|T201|COMP|43072-8|LNC|Brucella canis Ab.IgG|Brucella canis Ab.IgG
C1627323|T201|COMP|43073-6|LNC|Bovine leukemia virus Ab|Bovine leukemia virus Ab
C1627324|T201|COMP|43092-6|LNC|Arbovirus NOS Ab|Arbovirus NOS Ab
C1627327|T201|COMP|42804-5|LNC|Fungus identified|Fungus identified
C1627328|T201|COMP|42809-4|LNC|Fungus identified|Fungus identified
C1627329|T201|COMP|42810-2|LNC|Hemoglobin|Hemoglobin
C1627373|T201|COMP|42817-7|LNC|Cells.CD38+Kappa+/100 cells|Cells.CD38+Kappa+/100 cells
C1627381|T201|COMP|42862-3|LNC|Carbofuran|Carbofuran
C1627382|T201|COMP|42863-1|LNC|Libocedrus decurrens Ab.IgE/IgE.total|Libocedrus decurrens Ab.IgE/IgE.total
C1627383|T201|COMP|43032-2|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C1627384|T201|COMP|43036-3|LNC|Feline herpesvirus Ab|Feline herpesvirus Ab
C1627385|T201|COMP|43042-1|LNC|Echovirus 4 Ab|Echovirus 4 Ab
C1627386|T201|COMP|43044-7|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C1627387|T201|COMP|43052-0|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1627388|T201|COMP|43054-6|LNC|Clostridium tetani toxin Ab|Clostridium tetani toxin Ab
C1627422|T201|COMP|42993-6|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C1627423|T201|COMP|41479-7|LNC|BK virus DNA|BK virus DNA
C1627424|T201|COMP|42481-2|LNC|Human papilloma virus 6+11+42+43+44 DNA|Human papilloma virus 6+11+42+43+44 DNA
C1627425|T201|COMP|41490-4|LNC|Echovirus 16 Ab|Echovirus 16 Ab
C1627426|T201|COMP|41618-0|LNC|HLA Ab|HLA Ab
C1627427|T201|COMP|41628-9|LNC|Burkholderia sp DNA|Burkholderia sp DNA
C1627910|T201|COMP|42908-4|LNC|Hematocrit|Hematocrit
C1627911|T201|COMP|42909-2|LNC|Hemoglobin.gastrointestinal^1st specimen|Hemoglobin.gastrointestinal^1st specimen
C1627912|T201|COMP|42913-4|LNC|Hemoglobin.gastrointestinal^1st specimen|Hemoglobin.gastrointestinal^1st specimen
C1627913|T201|COMP|42914-2|LNC|HER2|HER2
C1627914|T201|COMP|42918-3|LNC|Hydroflumethiazide|Hydroflumethiazide
C1627915|T201|COMP|43074-4|LNC|Borrelia burgdorferi C6 Ab|Borrelia burgdorferi C6 Ab
C1627916|T201|COMP|43077-7|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C1627917|T201|COMP|43078-5|LNC|Bluetongue virus 2 Ab|Bluetongue virus 2 Ab
C1627918|T201|COMP|43079-3|LNC|Bluetongue virus 17 Ab|Bluetongue virus 17 Ab
C1627919|T201|COMP|43082-7|LNC|Bluetongue virus 10 Ab|Bluetongue virus 10 Ab
C1627920|T201|COMP|43084-3|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C1627921|T201|COMP|43086-8|LNC|Babesia divergens Ab|Babesia divergens Ab
C1627922|T201|COMP|43087-6|LNC|Babesia canis Ab|Babesia canis Ab
C1627923|T201|COMP|43090-0|LNC|Aspergillus flavus Ab|Aspergillus flavus Ab
C1627924|T201|COMP|43097-5|LNC|COL3A1 gene targeted mutation analysis|COL3A1 gene targeted mutation analysis
C1627925|T201|COMP|43109-8|LNC|Leishmania sp Ab.IgG & IgM panel|Leishmania sp Ab.IgG & IgM panel
C1627926|T201|COMP|43112-2|LNC|Herpes simplex virus Ab panel|Herpes simplex virus Ab panel
C1628433|T201|COMP|42191-7|LNC|Hepatitis A & B & C 7a panel|Hepatitis A & B & C 7a panel
C1628434|T201|COMP|42192-5|LNC|Nidus|Nidus
C1628435|T201|COMP|42195-8|LNC|Cells.CD8/100 cells|Cells.CD8/100 cells
C1628436|T201|COMP|42205-5|LNC|Human antimouse Ab.IgG|Human antimouse Ab.IgG
C1628437|T201|COMP|42208-9|LNC|IgM.CSF/IgM.serum|IgM.CSF/IgM.serum
C1628439|T201|COMP|42213-9|LNC|Nuclear Ab pattern.rim|Nuclear Ab pattern.rim
C1628440|T201|COMP|42864-9|LNC|Cells.CD103/100 cells|Cells.CD103/100 cells
C1628441|T201|COMP|42865-6|LNC|Cells.CD117/100 cells|Cells.CD117/100 cells
C1628442|T201|COMP|42868-0|LNC|Cells.CD11c+CD19+/100 cells|Cells.CD11c+CD19+/100 cells
C1628443|T201|COMP|42871-4|LNC|Cells.CD138/100 cells|Cells.CD138/100 cells
C1628444|T201|COMP|42872-2|LNC|Cells.CD138/100 cells|Cells.CD138/100 cells
C1628445|T201|COMP|42877-1|LNC|Cells.CD3-CD16+|Cells.CD3-CD16+
C1628446|T201|COMP|42880-5|LNC|Cells.CD3-CD57+|Cells.CD3-CD57+
C1628447|T201|COMP|42881-3|LNC|Cells.CD3-CD57+|Cells.CD3-CD57+
C1628448|T201|COMP|42885-4|LNC|Cells.CD52/100 cells|Cells.CD52/100 cells
C1628449|T201|COMP|42888-8|LNC|Cells.CD79b/100 cells|Cells.CD79b/100 cells
C1628450|T201|COMP|42893-8|LNC|Cladosporium herbarum Ab.IgG|Cladosporium herbarum Ab.IgG
C1628451|T201|COMP|42898-7|LNC|Cyclic citrullinated peptide Ab.IgG|Cyclic citrullinated peptide Ab.IgG
C1628452|T201|COMP|42907-6|LNC|Helminthosporium sp Ab.IgG|Helminthosporium sp Ab.IgG
C1628453|T201|COMP|43071-0|LNC|Brucella canis Ab.IgM|Brucella canis Ab.IgM
C1628454|T201|COMP|43075-1|LNC|Borrelia burgdorferi C6 Ab|Borrelia burgdorferi C6 Ab
C1628455|T201|COMP|43076-9|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C1628456|T201|COMP|43081-9|LNC|Bluetongue virus 11 Ab|Bluetongue virus 11 Ab
C1628457|T201|COMP|43083-5|LNC|Blastomyces sp Ab|Blastomyces sp Ab
C1628458|T201|COMP|43085-0|LNC|Babesia duncani Ab|Babesia duncani Ab
C1628459|T201|COMP|43089-2|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C1628460|T201|COMP|43091-8|LNC|Ascaris sp Ab|Ascaris sp Ab
C1628461|T201|COMP|43093-4|LNC|Angiostrongylus costaricensis Ab|Angiostrongylus costaricensis Ab
C1628462|T201|COMP|43094-2|LNC|Angiostrongylus cantonensis Ab|Angiostrongylus cantonensis Ab
C1628463|T201|COMP|43095-9|LNC|Anaplasma marginale Ab|Anaplasma marginale Ab
C1628464|T201|COMP|43098-3|LNC|Yersinia sp Ab panel|Yersinia sp Ab panel
C1628562|T201|COMP|42325-1|LNC|RHD+RHC gene targeted mutation analysis|RHD+RHC gene targeted mutation analysis
C1628563|T201|COMP|42330-1|LNC|Bordetella pertussis Ab.IgG|Bordetella pertussis Ab.IgG
C1628564|T201|COMP|42353-3|LNC|Cefepime+Clavulanate|Cefepime+Clavulanate
C1629068|T201|COMP|42317-8|LNC|Foscarnet|Foscarnet
C1629069|T201|COMP|42342-6|LNC|Rickettsia (Proteus) Ab panel|Rickettsia (Proteus) Ab panel
C1629575|T201|COMP|42177-6|LNC|Fc epsilon RI Ab|Fc epsilon RI Ab
C1629576|T201|COMP|42179-2|LNC|PLP1 gene duplication|PLP1 gene duplication
C1629577|T201|COMP|42184-2|LNC|Gossypol.positive isomer|Gossypol.positive isomer
C1629578|T201|COMP|42197-4|LNC|Centromere Ab|Centromere Ab
C1629579|T201|COMP|42202-2|LNC|GALOP Ab.IgM|GALOP Ab.IgM
C1629580|T201|COMP|42207-1|LNC|IgG.CSF/IgG.serum|IgG.CSF/IgG.serum
C1629581|T201|COMP|42214-7|LNC|Nuclear Ab pattern.speckled|Nuclear Ab pattern.speckled
C1629582|T201|COMP|42216-2|LNC|Reference lab name|Reference lab name
C1629583|T201|COMP|42218-8|LNC|Sulfatide Ab.IgG & Ab.IgM panel|Sulfatide Ab.IgG & Ab.IgM panel
C1629584|T201|COMP|42873-0|LNC|Cells.CD18/100 cells|Cells.CD18/100 cells
C1629585|T201|COMP|42875-5|LNC|Cells.CD22/100 cells|Cells.CD22/100 cells
C1629586|T201|COMP|42876-3|LNC|Cells.CD25+CD19+/100 cells|Cells.CD25+CD19+/100 cells
C1629587|T201|COMP|42878-9|LNC|Cells.CD3-CD16+|Cells.CD3-CD16+
C1629588|T201|COMP|42879-7|LNC|Cells.CD3-CD16+|Cells.CD3-CD16+
C1629589|T201|COMP|42884-7|LNC|Cells.CD52/100 cells|Cells.CD52/100 cells
C1629590|T201|COMP|42887-0|LNC|Cells.CD79b/100 cells|Cells.CD79b/100 cells
C1629591|T201|COMP|42892-0|LNC|Citrulline|Citrulline
C1629592|T201|COMP|42896-1|LNC|Colorado tick fever virus Ab.IgM|Colorado tick fever virus Ab.IgM
C1629593|T201|COMP|42906-8|LNC|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C1629594|T201|COMP|42915-9|LNC|Herpes virus 6 Ab.IgM|Herpes virus 6 Ab.IgM
C1629595|T201|COMP|42916-7|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1629596|T201|COMP|43088-4|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C1629597|T201|COMP|43096-7|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C1629626|T201|COMP|42322-8|LNC|Hepatitis B virus S+pol gene|Hepatitis B virus S+pol gene
C1629627|T201|COMP|42339-2|LNC|HIV 1 p24 Ag|HIV 1 p24 Ag
C1630168|T201|COMP|42223-8|LNC|Manganese/Creatinine|Manganese/Creatinine
C1630170|T201|COMP|42245-1|LNC|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C1630171|T201|COMP|42246-9|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C1630172|T201|COMP|42248-5|LNC|Hemoglobin.other/Hemoglobin.total|Hemoglobin.other/Hemoglobin.total
C1630173|T201|COMP|42257-6|LNC|Shigella dysenteriae Ag|Shigella dysenteriae Ag
C1630189|T201|COMP|42790-6|LNC|MAP kinase 14|MAP kinase 14
C1630740|T201|COMP|17625-5|LNC|Streptococcus pneumoniae 23f Ab^2nd specimen|Streptococcus pneumoniae 23f Ab^2nd specimen
C1630741|T201|COMP|42225-3|LNC|Thallium|Thallium
C1630744|T201|COMP|42233-7|LNC|Acetylcholine receptor ganglionic neuronal Ab|Acetylcholine receptor ganglionic neuronal Ab
C1630745|T201|COMP|42249-3|LNC|levETIRAcetam|levETIRAcetam
C1630746|T201|COMP|42254-3|LNC|Nuclear Ab|Nuclear Ab
C1630747|T201|COMP|42255-0|LNC|Salmonella & Shigella sp identified|Salmonella & Shigella sp identified
C1630748|T201|COMP|42258-4|LNC|Shigella flexneri Ag|Shigella flexneri Ag
C1630752|T201|COMP|43133-8|LNC|Allopurinol & Oxipurinol panel|Allopurinol & Oxipurinol panel
C1630767|T201|COMP|42519-9|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C1630768|T201|COMP|42625-4|LNC|Coxsackievirus A6 Ab|Coxsackievirus A6 Ab
C1630770|T201|COMP|42484-6|LNC|Protein.monoclonal/Protein.total|Protein.monoclonal/Protein.total
C1630771|T201|COMP|42489-5|LNC|Aureobasidium pullulans Ab|Aureobasidium pullulans Ab
C1631248|T201|COMP|42221-2|LNC|Manganese|Manganese
C1631251|T201|COMP|42250-1|LNC|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C1631252|T201|COMP|42259-2|LNC|Shigella sonnei Ag|Shigella sonnei Ag
C1631262|T201|COMP|43135-3|LNC|17-Ketosteroids & 17-Ketogenic steroids panel|17-Ketosteroids & 17-Ketogenic steroids panel
C1631263|T201|COMP|43141-1|LNC|Synthetic glucocorticoid panel|Synthetic glucocorticoid panel
C1631264|T201|COMP|43163-5|LNC|Quaternary ammonium compound|Quaternary ammonium compound
C1631777|T201|COMP|42224-6|LNC|Thallium|Thallium
C1631778|T201|COMP|42234-5|LNC|Alpha subunit.free|Alpha subunit.free
C1631779|T201|COMP|42247-7|LNC|Hemoglobin pattern|Hemoglobin pattern
C1631780|T201|COMP|42252-7|LNC|Methaqualone+Metabolite|Methaqualone+Metabolite
C1631781|T201|COMP|42253-5|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C1631782|T201|COMP|42256-8|LNC|Shigella boydii Ag|Shigella boydii Ag
C1631788|T201|COMP|43131-2|LNC|Bacterial Ag panel|Bacterial Ag panel
C1631817|T201|COMP|42494-5|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C1631820|T201|COMP|42957-1|LNC|SARS coronavirus Ab.IgG|SARS coronavirus Ab.IgG
C1632232|T201|COMP|42315-2|LNC|APOE gene alleles e2 & e3 & e4|APOE gene alleles e2 & e3 & e4
C1632233|T201|COMP|42501-7|LNC|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C1632234|T201|COMP|42503-3|LNC|Hantavirus Ab|Hantavirus Ab
C1632235|T201|COMP|42963-9|LNC|Salmonella paratyphi C H Ab|Salmonella paratyphi C H Ab
C1632236|T201|COMP|42318-6|LNC|GALT gene targeted mutation analysis|GALT gene targeted mutation analysis
C1632237|T201|COMP|42319-4|LNC|Glucose-6-Phosphate dehydrogenase phenotype|Glucose-6-Phosphate dehydrogenase phenotype
C1632260|T201|COMP|42644-5|LNC|Ciprofloxacin 2.0 ug/mL|Ciprofloxacin 2.0 ug/mL
C1632261|T201|COMP|42675-9|LNC|HLA Ag|HLA Ag
C1632263|T201|COMP|42731-0|LNC|Cardiolipin Ab.IgG.B2GP1 dependent|Cardiolipin Ab.IgG.B2GP1 dependent
C1632264|T201|COMP|41722-0|LNC|Telithromycin|Telithromycin
C1632266|T201|COMP|42894-6|LNC|Clindamycin Ab.IgE|Clindamycin Ab.IgE
C1632267|T201|COMP|43013-2|LNC|HIV 1 gp120+gp160 Ab|HIV 1 gp120+gp160 Ab
C1632336|T201|COMP|42354-1|LNC|Tigecycline|Tigecycline
C1632341|T201|COMP|42316-0|LNC|RHD gene targeted mutation analysis|RHD gene targeted mutation analysis
C1632342|T201|COMP|42500-9|LNC|Fosamprenavir|Fosamprenavir
C1632343|T201|COMP|42504-1|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C1632344|T201|COMP|42505-8|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C1632345|T201|COMP|42965-4|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C1632346|T201|COMP|42968-8|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C1632347|T201|COMP|42975-3|LNC|Powassan virus Ab|Powassan virus Ab
C1632348|T201|COMP|42321-0|LNC|HTT gene targeted mutation analysis|HTT gene targeted mutation analysis
C1632349|T201|COMP|42324-4|LNC|I group phenotype|I group phenotype
C1632362|T201|COMP|42956-3|LNC|SARS coronavirus Ab.IgM|SARS coronavirus Ab.IgM
C1632363|T201|COMP|42765-8|LNC|Tube number|Tube number
C1632364|T201|COMP|41493-8|LNC|Febrile agglutinin Ab panel|Febrile agglutinin Ab panel
C1632366|T201|COMP|42995-1|LNC|Leptospira borgpetersenii serovar Tarrasovi Ab|Leptospira borgpetersenii serovar Tarrasovi Ab
C1632367|T201|COMP|42524-9|LNC|Mucus|Mucus
C1632368|T201|COMP|41862-4|LNC|Viscosity^20M post collection|Viscosity^20M post collection
C1632370|T201|COMP|42935-7|LNC|Pyrazinamide 100.0 ug/mL|Pyrazinamide 100.0 ug/mL
C1632371|T201|COMP|43047-0|LNC|Coxsackievirus A7 Ab|Coxsackievirus A7 Ab
C1632374|T201|COMP|42601-5|LNC|Immune complex.IgG|Immune complex.IgG
C1632378|T201|COMP|41654-5|LNC|Hematocrit|Hematocrit
C1632379|T201|COMP|42900-1|LNC|Daucus carota Ab.IgE/IgE.total|Daucus carota Ab.IgE/IgE.total
C1632381|T201|COMP|42931-6|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1632384|T201|COMP|42206-3|LNC|IgA.CSF/IgA.serum|IgA.CSF/IgA.serum
C1632385|T201|COMP|42212-1|LNC|Nuclear Ab pattern.nucleolar|Nuclear Ab pattern.nucleolar
C1632386|T201|COMP|42217-0|LNC|Striated muscle Ab.IgG|Striated muscle Ab.IgG
C1632387|T201|COMP|42222-0|LNC|Manganese|Manganese
C1632389|T201|COMP|43041-3|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C1632390|T201|COMP|42502-5|LNC|Glycolate|Glycolate
C1632391|T201|COMP|42966-2|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C1632392|T201|COMP|42352-5|LNC|cefTAZidime+Clavulanate|cefTAZidime+Clavulanate
C1632783|T201|COMP|42952-2|LNC|Snowshoe hare virus Ab|Snowshoe hare virus Ab
C1632784|T201|COMP|42958-9|LNC|Salmonella typhimurium Ab|Salmonella typhimurium Ab
C1632787|T201|COMP|42329-3|LNC|Bordetella pertussis Ab.IgM|Bordetella pertussis Ab.IgM
C1632788|T201|COMP|42331-9|LNC|Nuclear Ab.IgG|Nuclear Ab.IgG
C1632791|T201|COMP|42337-6|LNC|Herpes simplex virus 1 glycoprotein G Ab.IgG|Herpes simplex virus 1 glycoprotein G Ab.IgG
C1632792|T201|COMP|42340-0|LNC|HTLV I p42 Ab|HTLV I p42 Ab
C1632793|T201|COMP|42341-8|LNC|Neisseria meningitidis serogroups A+w135 Ag|Neisseria meningitidis serogroups A+w135 Ag
C1632795|T201|COMP|42365-7|LNC|Streptococcus pneumoniae 4 serotypes Ab.IgG panel|Streptococcus pneumoniae 4 serotypes Ab.IgG panel
C1632796|T201|COMP|42370-7|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C1632797|T201|COMP|42374-9|LNC|Neisseria meningitidis serogroup Y Ag|Neisseria meningitidis serogroup Y Ag
C1632957|T201|COMP|42499-4|LNC|Fibrin D-dimer|Fibrin D-dimer
C1632958|T201|COMP|42508-2|LNC|Herpes virus 8 Ab.IgG|Herpes virus 8 Ab.IgG
C1632959|T201|COMP|42509-0|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C1632960|T201|COMP|42510-8|LNC|IgD|IgD
C1632961|T201|COMP|42971-2|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1632962|T201|COMP|42972-0|LNC|Powassan virus Ab.IgM|Powassan virus Ab.IgM
C1632963|T201|COMP|42974-6|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1632977|T201|COMP|41841-8|LNC|Coxiella burnetii phase 1 & 2 Ab.IgM panel|Coxiella burnetii phase 1 & 2 Ab.IgM panel
C1632978|T201|COMP|41856-6|LNC|Variola virus DNA|Variola virus DNA
C1632979|T201|COMP|41687-5|LNC|Clavulanate|Clavulanate
C1632990|T201|COMP|42372-3|LNC|Neisseria meningitidis serogroup D Ag|Neisseria meningitidis serogroup D Ag
C1633391|T201|COMP|42953-0|LNC|Snowshoe hare virus Ab.IgM|Snowshoe hare virus Ab.IgM
C1633392|T201|COMP|42955-5|LNC|Semliki forest virus Ab|Semliki forest virus Ab
C1633393|T201|COMP|41494-6|LNC|Gatifloxacin|Gatifloxacin
C1633394|T201|COMP|41498-7|LNC|HIV 1 RNA|HIV 1 RNA
C1633395|T201|COMP|41502-6|LNC|Moxifloxacin|Moxifloxacin
C1633396|T201|COMP|41503-4|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C1633397|T201|COMP|41504-2|LNC|Norfloxacin|Norfloxacin
C1633405|T201|COMP|42343-4|LNC|Toxoplasma gondii identified|Toxoplasma gondii identified
C1633445|T201|COMP|42355-8|LNC|Tigecycline|Tigecycline
C1633449|T201|COMP|42964-7|LNC|Salmonella paratyphi B O Ab|Salmonella paratyphi B O Ab
C1633450|T201|COMP|42967-0|LNC|Rubella virus Ab|Rubella virus Ab
C1633451|T201|COMP|42969-6|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C1633452|T201|COMP|42320-2|LNC|Glutathione reductase phenotype|Glutathione reductase phenotype
C1633453|T201|COMP|42323-6|LNC|HLA-DR Ag|HLA-DR Ag
C1633468|T201|COMP|41394-8|LNC|Collection date|Collection date
C1633476|T201|COMP|42857-3|LNC|Calcium|Calcium
C1633479|T201|COMP|42201-4|LNC|DNA single strand Ab.IgG|DNA single strand Ab.IgG
C1633480|T201|COMP|43080-1|LNC|Bluetongue virus 13 Ab|Bluetongue virus 13 Ab
C1634494|T201|COMP|42951-4|LNC|Taylorella equigenitalis Ab|Taylorella equigenitalis Ab
C1634495|T201|COMP|42954-8|LNC|Sindbis virus Ab|Sindbis virus Ab
C1634496|T201|COMP|41496-1|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C1634497|T201|COMP|41497-9|LNC|HIV 1 RNA|HIV 1 RNA
C1634498|T201|COMP|41499-5|LNC|Legionella pneumophila 1 Ag|Legionella pneumophila 1 Ag
C1634499|T201|COMP|41501-8|LNC|Measles virus Ab|Measles virus Ab
C1634505|T201|COMP|42368-1|LNC|Neisseria meningitidis serogroup w135 Ag|Neisseria meningitidis serogroup w135 Ag
C1634995|T201|COMP|42236-0|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C1634996|T201|COMP|42238-6|LNC|Borrelia burgdorferi 23kD Ab|Borrelia burgdorferi 23kD Ab
C1634997|T201|COMP|42243-6|LNC|Hemoglobin|Hemoglobin
C1635003|T201|COMP|41290-8|LNC|HIV 1+2 Ab.IgM|HIV 1+2 Ab.IgM
C1635066|T201|COMP|42350-9|LNC|Cefepime+Clavulanate|Cefepime+Clavulanate
C1635610|T201|COMP|42240-2|LNC|CHD7 gene targeted mutation analysis|CHD7 gene targeted mutation analysis
C1635612|T201|COMP|42933-2|LNC|Cells.CD79a/100 cells|Cells.CD79a/100 cells
C1635613|T201|COMP|42934-0|LNC|Cells.CD83/100 cells|Cells.CD83/100 cells
C1635614|T201|COMP|42938-1|LNC|CFTR gene allele 1|CFTR gene allele 1
C1635615|T201|COMP|42940-7|LNC|GALT gene allele 1|GALT gene allele 1
C1635644|T201|COMP|42356-6|LNC|Tigecycline|Tigecycline
C1635645|T201|COMP|42358-2|LNC|HLA-B*57:01|HLA-B*57:01
C1635646|T201|COMP|42950-6|LNC|Toxocara canis Ab|Toxocara canis Ab
C1635647|T201|COMP|41495-3|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C1635648|T201|COMP|41500-0|LNC|Linezolid|Linezolid
C1635649|T201|COMP|41505-9|LNC|Parainfluenza virus Ag panel|Parainfluenza virus Ag panel
C1635653|T201|COMP|42326-9|LNC|Drugs identified|Drugs identified
C1635654|T201|COMP|42328-5|LNC|Bordetella pertussis Ab.IgA|Bordetella pertussis Ab.IgA
C1635655|T201|COMP|42336-8|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C1635656|T201|COMP|42338-4|LNC|Herpes simplex virus 2 glycoprotein G Ab.IgG|Herpes simplex virus 2 glycoprotein G Ab.IgG
C1635658|T201|COMP|42351-7|LNC|Cefepime+Clavulanate|Cefepime+Clavulanate
C1635659|T201|COMP|42369-9|LNC|Neisseria meningitidis serogroup A Ag|Neisseria meningitidis serogroup A Ag
C1635660|T201|COMP|42373-1|LNC|Neisseria meningitidis serogroup X Ag|Neisseria meningitidis serogroup X Ag
C1635661|T201|COMP|42376-4|LNC|Neisseria meningitidis serogroup Z' Ag|Neisseria meningitidis serogroup Z' Ag
C1636058|T201|COMP|42242-8|LNC|Ethanol|Ethanol
C1636064|T201|COMP|42936-5|LNC|Intercellular substance Ab.IgA|Intercellular substance Ab.IgA
C1637219|T201|COMP|22553-2|LNC|Streptococcus pneumoniae 7f Ab^1st specimen|Streptococcus pneumoniae 7f Ab^1st specimen
C1637228|T201|COMP|41397-1|LNC|Beta lactoglobulin Ab.IgE|Beta lactoglobulin Ab.IgE
C1637232|T201|COMP|42482-0|LNC|Protein.monoclonal|Protein.monoclonal
C1637233|T201|COMP|42486-1|LNC|Aspergillus fumigatus 1 Ab|Aspergillus fumigatus 1 Ab
C1637234|T201|COMP|42492-9|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C1637235|T201|COMP|42498-6|LNC|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C1637236|T201|COMP|42513-2|LNC|IgE|IgE
C1637237|T201|COMP|42518-1|LNC|Leptospira sp Ab|Leptospira sp Ab
C1637238|T201|COMP|42521-5|LNC|Saccharopolyspora rectivirgula Ab|Saccharopolyspora rectivirgula Ab
C1637239|T201|COMP|42525-6|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C1637240|T201|COMP|42528-0|LNC|Phenothiazines|Phenothiazines
C1637241|T201|COMP|42534-8|LNC|Thermoactinomyces vulgaris Ab|Thermoactinomyces vulgaris Ab
C1637274|T201|COMP|41294-0|LNC|Cells.S phase|Cells.S phase
C1637791|T201|COMP|41396-3|LNC|Tenofovir|Tenofovir
C1637792|T201|COMP|41398-9|LNC|Alloisoleucine|Alloisoleucine
C1637793|T201|COMP|41399-7|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1638282|T201|COMP|42488-7|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C1638283|T201|COMP|42493-7|LNC|Catecholamines.free fractionated|Catecholamines.free fractionated
C1638284|T201|COMP|42520-7|LNC|Methylmalonate|Methylmalonate
C1638285|T201|COMP|42523-1|LNC|Molindone|Molindone
C1638286|T201|COMP|42526-4|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C1638287|T201|COMP|42538-9|LNC|Hydroxyperhexiline|Hydroxyperhexiline
C1638453|T201|COMP|42237-8|LNC|Borrelia burgdorferi 18kD Ab.IgG|Borrelia burgdorferi 18kD Ab.IgG
C1638454|T201|COMP|42244-4|LNC|Hemoglobin A/Hemoglobin.total|Hemoglobin A/Hemoglobin.total
C1638460|T201|COMP|42939-9|LNC|CFTR gene allele 2|CFTR gene allele 2
C1638461|T201|COMP|41293-2|LNC|Clot|Clot
C1638885|T201|COMP|41395-5|LNC|Collection date|Collection date
C1638887|T201|COMP|42490-3|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C1638888|T201|COMP|42491-1|LNC|Cannabinoids|Cannabinoids
C1638889|T201|COMP|42511-6|LNC|IgD|IgD
C1638890|T201|COMP|42512-4|LNC|IgE|IgE
C1638891|T201|COMP|42515-7|LNC|Jamestown canyon virus RNA|Jamestown canyon virus RNA
C1638892|T201|COMP|42536-3|LNC|Tropheryma whippelii DNA|Tropheryma whippelii DNA
C1638893|T201|COMP|42537-1|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C1639387|T201|COMP|42990-2|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C1639388|T201|COMP|42992-8|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C1639389|T201|COMP|42997-7|LNC|Leptospira autumnalis Ab|Leptospira autumnalis Ab
C1639390|T201|COMP|41400-3|LNC|Yersinia sp Ab.IgA|Yersinia sp Ab.IgA
C1639391|T201|COMP|41411-0|LNC|Angiostrongylus cantonensis Ab|Angiostrongylus cantonensis Ab
C1639392|T201|COMP|41413-6|LNC|Babesia divergens Ab|Babesia divergens Ab
C1639393|T201|COMP|41422-7|LNC|Schistosoma haematobium Ab|Schistosoma haematobium Ab
C1639394|T201|COMP|41425-0|LNC|Toxocara canis Ab|Toxocara canis Ab
C1639395|T201|COMP|41426-8|LNC|Trichinella spiralis Ab|Trichinella spiralis Ab
C1639401|T201|COMP|42575-1|LNC|Amoxicillin Ab.IgE/IgE.total|Amoxicillin Ab.IgE/IgE.total
C1639402|T201|COMP|42585-0|LNC|Bendiocarb|Bendiocarb
C1639403|T201|COMP|42596-7|LNC|Corticotropin^30M post XXX challenge|Corticotropin^30M post XXX challenge
C1639404|T201|COMP|42600-7|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C1639405|T201|COMP|42603-1|LNC|Coxsackievirus A6 Ab|Coxsackievirus A6 Ab
C1639534|T201|COMP|42483-8|LNC|Protein.monoclonal/Protein.total|Protein.monoclonal/Protein.total
C1639535|T201|COMP|42485-3|LNC|Anion gap|Anion gap
C1639536|T201|COMP|42487-9|LNC|Aspergillus fumigatus 6 Ab|Aspergillus fumigatus 6 Ab
C1639537|T201|COMP|42495-2|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C1639538|T201|COMP|42514-0|LNC|Inhibin Ag|Inhibin Ag
C1639539|T201|COMP|42516-5|LNC|Legionella sp Ab|Legionella sp Ab
C1639540|T201|COMP|42517-3|LNC|Leishmania sp Ab|Leishmania sp Ab
C1639541|T201|COMP|42522-3|LNC|Mitochondria Ab|Mitochondria Ab
C1639542|T201|COMP|42529-8|LNC|Pigeon serum Ab|Pigeon serum Ab
C1639543|T201|COMP|42530-6|LNC|Smooth muscle Ab|Smooth muscle Ab
C1639544|T201|COMP|42531-4|LNC|Spermatozoa.motile|Spermatozoa.motile
C1639910|T201|COMP|41401-1|LNC|Yersinia sp Ab.IgG|Yersinia sp Ab.IgG
C1639911|T201|COMP|41402-9|LNC|Emtricitabine|Emtricitabine
C1639912|T201|COMP|41403-7|LNC|Atazanavir|Atazanavir
C1639913|T201|COMP|41404-5|LNC|17-Hydroxycorticosteroids/Creatinine|17-Hydroxycorticosteroids/Creatinine
C1639914|T201|COMP|41405-2|LNC|Parainfluenza virus 2 Ab.IgG|Parainfluenza virus 2 Ab.IgG
C1639915|T201|COMP|41408-6|LNC|Ofloxacin 1.0 ug/mL|Ofloxacin 1.0 ug/mL
C1639916|T201|COMP|41409-4|LNC|Ofloxacin 2.0 ug/mL|Ofloxacin 2.0 ug/mL
C1639917|T201|COMP|41414-4|LNC|Babesia microti Ab|Babesia microti Ab
C1639918|T201|COMP|41417-7|LNC|Filaria Ab|Filaria Ab
C1639919|T201|COMP|41419-3|LNC|Leishmania braziliensis Ab|Leishmania braziliensis Ab
C1639920|T201|COMP|41420-1|LNC|Leishmania tropica Ab|Leishmania tropica Ab
C1639921|T201|COMP|41421-9|LNC|Paragonimus sp Ab|Paragonimus sp Ab
C1639922|T201|COMP|41423-5|LNC|Schistosoma japonicum Ab|Schistosoma japonicum Ab
C1639923|T201|COMP|41427-6|LNC|Trypanosoma brucei gambiense Ab|Trypanosoma brucei gambiense Ab
C1639932|T201|COMP|42572-8|LNC|11-Deoxycortisol|11-Deoxycortisol
C1639933|T201|COMP|42573-6|LNC|18-Hydroxycorticosterone|18-Hydroxycorticosterone
C1639934|T201|COMP|42574-4|LNC|1-Naphthol|1-Naphthol
C1639935|T201|COMP|42576-9|LNC|Amphetamine|Amphetamine
C1639936|T201|COMP|42578-5|LNC|Artifact|Artifact
C1639937|T201|COMP|42581-9|LNC|Babesia sp Ab.IgG|Babesia sp Ab.IgG
C1639938|T201|COMP|42593-4|LNC|Calcium|Calcium
C1640452|T201|COMP|42989-4|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C1640453|T201|COMP|42991-0|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C1640454|T201|COMP|42996-9|LNC|Leptospira borgpetersenii serovar Ballum Ab|Leptospira borgpetersenii serovar Ballum Ab
C1640455|T201|COMP|42998-5|LNC|Leishmania tropica Ab|Leishmania tropica Ab
C1640456|T201|COMP|41406-0|LNC|Meropenem|Meropenem
C1640457|T201|COMP|41412-8|LNC|Angiostrongylus costaricensis Ab|Angiostrongylus costaricensis Ab
C1640458|T201|COMP|41416-9|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C1640459|T201|COMP|41429-2|LNC|Acanthamoeba sp DNA|Acanthamoeba sp DNA
C1640464|T201|COMP|42570-2|LNC|Sodium|Sodium
C1640465|T201|COMP|42579-3|LNC|Aspergillus fumigatus Ab.IgM|Aspergillus fumigatus Ab.IgM
C1640466|T201|COMP|42580-1|LNC|Babesia sp Ab.IgM|Babesia sp Ab.IgM
C1640467|T201|COMP|42595-9|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1640468|T201|COMP|42597-5|LNC|Corticotropin^1.5H post XXX challenge|Corticotropin^1.5H post XXX challenge
C1640469|T201|COMP|42598-3|LNC|Corticotropin^baseline|Corticotropin^baseline
C1640470|T201|COMP|42604-9|LNC|Glucose^3H post dose lactose PO|Glucose^3H post dose lactose PO
C1640471|T201|COMP|42606-4|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C1640472|T201|COMP|42357-4|LNC|Tigecycline|Tigecycline
C1640473|T201|COMP|42239-4|LNC|Borrelia burgdorferi 39kD Ab.IgG|Borrelia burgdorferi 39kD Ab.IgG
C1641049|T201|COMP|42994-4|LNC|Leptospira sp Ab|Leptospira sp Ab
C1641050|T201|COMP|42999-3|LNC|Leishmania sp Ab|Leishmania sp Ab
C1641051|T201|COMP|41418-5|LNC|Gnathostoma sp Ab|Gnathostoma sp Ab
C1641052|T201|COMP|41428-4|LNC|Trypanosoma brucei rhodesiense Ab|Trypanosoma brucei rhodesiense Ab
C1641056|T201|COMP|42577-7|LNC|Ampicillin Ab.IgE/IgE.total|Ampicillin Ab.IgE/IgE.total
C1641057|T201|COMP|42582-7|LNC|Barbiturates|Barbiturates
C1641058|T201|COMP|42586-8|LNC|Benzodiazepines|Benzodiazepines
C1641059|T201|COMP|42587-6|LNC|BK virus DNA|BK virus DNA
C1641060|T201|COMP|42588-4|LNC|Bordetella parapertussis DNA|Bordetella parapertussis DNA
C1641061|T201|COMP|42590-0|LNC|Borrelia sp Ab|Borrelia sp Ab
C1641062|T201|COMP|42591-8|LNC|Botrytis cinerea Ab.IgG|Botrytis cinerea Ab.IgG
C1641063|T201|COMP|42602-3|LNC|Tropheryma whippelii DNA|Tropheryma whippelii DNA
C1641480|T201|COMP|41432-6|LNC|Balamuthia mandrillaris DNA|Balamuthia mandrillaris DNA
C1641481|T201|COMP|41442-5|LNC|Entamoeba dispar DNA|Entamoeba dispar DNA
C1641482|T201|COMP|41443-3|LNC|Enterocytozoon bieneusi DNA|Enterocytozoon bieneusi DNA
C1641483|T201|COMP|41446-6|LNC|Parasite identified|Parasite identified
C1641484|T201|COMP|41448-2|LNC|Plasmodium malariae DNA|Plasmodium malariae DNA
C1641485|T201|COMP|41461-5|LNC|Virus identified|Virus identified
C1641486|T201|COMP|41463-1|LNC|Wuchereria bancrofti+Brugia malayi Ag|Wuchereria bancrofti+Brugia malayi Ag
C1641487|T201|COMP|41467-2|LNC|Benzodiazepines/Creatinine|Benzodiazepines/Creatinine
C1641488|T201|COMP|41469-8|LNC|Ribavirin|Ribavirin
C1641489|T201|COMP|41475-5|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C1641490|T201|COMP|41476-3|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C1641491|T201|COMP|41478-9|LNC|Bartonella henselae Ab.IgG & IgM panel|Bartonella henselae Ab.IgG & IgM panel
C1641492|T201|COMP|42610-6|LNC|Salicylurate|Salicylurate
C1641493|T201|COMP|42611-4|LNC|Glucose^1H post dose lactose PO|Glucose^1H post dose lactose PO
C1641494|T201|COMP|42614-8|LNC|Colorado tick fever virus Ab|Colorado tick fever virus Ab
C1641495|T201|COMP|42623-9|LNC|Coxsackievirus A3 Ab|Coxsackievirus A3 Ab
C1641496|T201|COMP|42629-6|LNC|Glucose^4H post dose lactose PO|Glucose^4H post dose lactose PO
C1641497|T201|COMP|42643-7|LNC|Capreomycin 10.0 ug/mL|Capreomycin 10.0 ug/mL
C1641498|T201|COMP|42646-0|LNC|Ethambutol 5.0 ug/mL|Ethambutol 5.0 ug/mL
C1641499|T201|COMP|42656-9|LNC|Rifabutin 2.0 ug/mL|Rifabutin 2.0 ug/mL
C1641500|T201|COMP|42666-8|LNC|Fat.neutral|Fat.neutral
C1641501|T201|COMP|41424-3|LNC|Schistosoma mansoni Ab|Schistosoma mansoni Ab
C1641502|T201|COMP|41440-9|LNC|Encephalitozoon hellem DNA|Encephalitozoon hellem DNA
C1641503|T201|COMP|41453-2|LNC|Human coronavirus Ag|Human coronavirus Ag
C1641504|T201|COMP|41509-1|LNC|Toxoplasma sp Ab.IgG|Toxoplasma sp Ab.IgG
C1641505|T201|COMP|41512-5|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C1641506|T201|COMP|41598-4|LNC|Bacteria|Bacteria
C1641507|T201|COMP|41607-3|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C1641508|T201|COMP|41611-5|LNC|Tube number|Tube number
C1641509|T201|COMP|41613-1|LNC|Tube number|Tube number
C1641510|T201|COMP|41619-8|LNC|Hemoglobin.unstable|Hemoglobin.unstable
C1641511|T201|COMP|41625-5|LNC|Brucella sp DNA|Brucella sp DNA
C1641512|T201|COMP|41630-5|LNC|Clostridium botulinum toxin A|Clostridium botulinum toxin A
C1641513|T201|COMP|41633-9|LNC|Clostridium botulinum toxin B botB gene|Clostridium botulinum toxin B botB gene
C1641514|T201|COMP|41646-1|LNC|Calcium.ionized|Calcium.ionized
C1641515|T201|COMP|41647-9|LNC|Carbon dioxide|Carbon dioxide
C1641516|T201|COMP|41648-7|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C1641517|T201|COMP|41650-3|LNC|Chloride|Chloride
C1641518|T201|COMP|41652-9|LNC|Glucose|Glucose
C1641519|T201|COMP|41724-6|LNC|Thiamphenicol|Thiamphenicol
C1641520|T201|COMP|41733-7|LNC|Clavulanate|Clavulanate
C1641521|T201|COMP|41736-0|LNC|Oritavancin|Oritavancin
C1641522|T201|COMP|41737-8|LNC|Ramoplanin|Ramoplanin
C1641523|T201|COMP|41744-4|LNC|Beclomethasone dipropionate|Beclomethasone dipropionate
C1641524|T201|COMP|41747-7|LNC|Budesonide|Budesonide
C1641525|T201|COMP|41754-3|LNC|Fludrocortisone|Fludrocortisone
C1641526|T201|COMP|41762-6|LNC|Megestrol acetate|Megestrol acetate
C1641527|T201|COMP|41764-2|LNC|SBDS gene targeted mutation analysis|SBDS gene targeted mutation analysis
C1641528|T201|COMP|41766-7|LNC|Triamcinolone|Triamcinolone
C1642048|T201|COMP|41435-9|LNC|Cyclospora carcopitheci DNA|Cyclospora carcopitheci DNA
C1642049|T201|COMP|41438-3|LNC|Cyclospora papionis DNA|Cyclospora papionis DNA
C1642050|T201|COMP|41447-4|LNC|Plasmodium falciparum DNA|Plasmodium falciparum DNA
C1642051|T201|COMP|41452-4|LNC|Adenovirus serotype|Adenovirus serotype
C1642052|T201|COMP|41458-1|LNC|SARS coronavirus RNA|SARS coronavirus RNA
C1642053|T201|COMP|41473-0|LNC|carBAMazepine 10,11-Epoxide|carBAMazepine 10,11-Epoxide
C1642054|T201|COMP|41491-2|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C1642055|T201|COMP|42613-0|LNC|Glucose^2H post dose lactose PO|Glucose^2H post dose lactose PO
C1642056|T201|COMP|42616-3|LNC|Magnesium|Magnesium
C1642057|T201|COMP|42618-9|LNC|Naloxone|Naloxone
C1642059|T201|COMP|42621-3|LNC|Mycoplasma hominis DNA|Mycoplasma hominis DNA
C1642060|T201|COMP|42624-7|LNC|Gastrin^2M post XXX challenge|Gastrin^2M post XXX challenge
C1642061|T201|COMP|42634-6|LNC|1p & 19q chromosome deletion|1p & 19q chromosome deletion
C1642062|T201|COMP|42639-5|LNC|Immune complex.IgG|Immune complex.IgG
C1642063|T201|COMP|42652-8|LNC|Kanamycin 5.0 ug/mL|Kanamycin 5.0 ug/mL
C1642064|T201|COMP|42653-6|LNC|Ofloxacin 2.0 ug/mL|Ofloxacin 2.0 ug/mL
C1642065|T201|COMP|42660-1|LNC|Alpha 2 laminin|Alpha 2 laminin
C1642066|T201|COMP|42663-5|LNC|HLA-Cw locus|HLA-Cw locus
C1642067|T201|COMP|42667-6|LNC|Fatty acids|Fatty acids
C1642069|T201|COMP|41510-9|LNC|Toxoplasma sp Ab.IgM|Toxoplasma sp Ab.IgM
C1642070|T201|COMP|41514-1|LNC|HIV 1 RNA|HIV 1 RNA
C1642071|T201|COMP|41600-8|LNC|Bacteria|Bacteria
C1642072|T201|COMP|41605-7|LNC|Lactose^pre CFst|Lactose^pre CFst
C1642073|T201|COMP|41606-5|LNC|Lactose^3H post dose lactose PO|Lactose^3H post dose lactose PO
C1642074|T201|COMP|41610-7|LNC|Tube number|Tube number
C1642075|T201|COMP|41624-8|LNC|Brucella sp Ag|Brucella sp Ag
C1642076|T201|COMP|41638-8|LNC|Marburg virus RNA|Marburg virus RNA
C1642077|T201|COMP|41643-8|LNC|West Nile virus Ag|West Nile virus Ag
C1642078|T201|COMP|41655-2|LNC|Hematocrit|Hematocrit
C1642079|T201|COMP|41725-3|LNC|Thiamphenicol|Thiamphenicol
C1642080|T201|COMP|41729-5|LNC|cefoTEtan+Clavulanate|cefoTEtan+Clavulanate
C1642081|T201|COMP|41732-9|LNC|cefTRIAXone+Clavulanate|cefTRIAXone+Clavulanate
C1642082|T201|COMP|41735-2|LNC|Everninomicin|Everninomicin
C1642083|T201|COMP|41739-4|LNC|Sulbactam|Sulbactam
C1642540|T201|COMP|41431-8|LNC|Angiostrongylus costaricensis DNA|Angiostrongylus costaricensis DNA
C1642541|T201|COMP|41436-7|LNC|Cyclospora cayetanensis DNA|Cyclospora cayetanensis DNA
C1642542|T201|COMP|41437-5|LNC|Cyclospora colobi DNA|Cyclospora colobi DNA
C1642543|T201|COMP|41444-1|LNC|Naegleria fowleri DNA|Naegleria fowleri DNA
C1642544|T201|COMP|41449-0|LNC|Plasmodium ovale DNA|Plasmodium ovale DNA
C1642545|T201|COMP|41450-8|LNC|Plasmodium vivax DNA|Plasmodium vivax DNA
C1642546|T201|COMP|41454-0|LNC|Human coronavirus identified|Human coronavirus identified
C1642547|T201|COMP|41462-3|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C1642548|T201|COMP|41470-6|LNC|Atazanavir|Atazanavir
C1642549|T201|COMP|41477-1|LNC|Bacterial sialidase|Bacterial sialidase
C1642550|T201|COMP|41485-4|LNC|Coxsackievirus B Ab panel|Coxsackievirus B Ab panel
C1642551|T201|COMP|41486-2|LNC|Coxsackievirus B Ab panel|Coxsackievirus B Ab panel
C1642552|T201|COMP|41487-0|LNC|Cryptosporidium parvum Ag|Cryptosporidium parvum Ag
C1642553|T201|COMP|41489-6|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C1642554|T201|COMP|42609-8|LNC|Glucose^6H post dose lactose PO|Glucose^6H post dose lactose PO
C1642555|T201|COMP|42628-8|LNC|Cells.CD9+CD41+/100 cells|Cells.CD9+CD41+/100 cells
C1642556|T201|COMP|42631-2|LNC|Glucose^5H post dose lactose PO|Glucose^5H post dose lactose PO
C1642558|T201|COMP|42635-3|LNC|Chromosome 12p tetrasomy|Chromosome 12p tetrasomy
C1642559|T201|COMP|42637-9|LNC|Natriuretic peptide.B|Natriuretic peptide.B
C1642560|T201|COMP|42648-6|LNC|Ethionamide 5.0 ug/mL|Ethionamide 5.0 ug/mL
C1642561|T201|COMP|42651-0|LNC|Isoniazid 5.0 ug/mL|Isoniazid 5.0 ug/mL
C1642562|T201|COMP|42659-3|LNC|Streptomycin 2.0 ug/mL|Streptomycin 2.0 ug/mL
C1642563|T201|COMP|42662-7|LNC|Benzodiazepines|Benzodiazepines
C1642565|T201|COMP|41410-2|LNC|Ofloxacin 4.0 ug/mL|Ofloxacin 4.0 ug/mL
C1642566|T201|COMP|41464-9|LNC|Amphetamines/Creatinine|Amphetamines/Creatinine
C1642567|T201|COMP|41465-6|LNC|Opiates/Creatinine|Opiates/Creatinine
C1642568|T201|COMP|41482-1|LNC|Chlamydia sp Ab.IgG & IgM panel|Chlamydia sp Ab.IgG & IgM panel
C1642569|T201|COMP|41513-3|LNC|HIV 1 RNA|HIV 1 RNA
C1642570|T201|COMP|41599-2|LNC|Bacteria|Bacteria
C1642571|T201|COMP|41602-4|LNC|Bacteria|Bacteria
C1642572|T201|COMP|41603-2|LNC|Bacteria|Bacteria
C1642573|T201|COMP|41608-1|LNC|Prolactin^30M post XXX challenge|Prolactin^30M post XXX challenge
C1642574|T201|COMP|41612-3|LNC|Tube number|Tube number
C1642575|T201|COMP|41615-6|LNC|Xanthurenate|Xanthurenate
C1642576|T201|COMP|41634-7|LNC|Clostridium botulinum toxin E|Clostridium botulinum toxin E
C1642577|T201|COMP|41636-2|LNC|Ebola virus RNA|Ebola virus RNA
C1642578|T201|COMP|41640-4|LNC|Ricin toxin Ab.IgG|Ricin toxin Ab.IgG
C1642579|T201|COMP|41641-2|LNC|Ricin toxin|Ricin toxin
C1642580|T201|COMP|41642-0|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1642581|T201|COMP|41644-6|LNC|Calcium.ionized|Calcium.ionized
C1642582|T201|COMP|41728-7|LNC|Biapenem|Biapenem
C1642583|T201|COMP|41730-3|LNC|cefOXitin+Clavulanate|cefOXitin+Clavulanate
C1642584|T201|COMP|41734-5|LNC|Dalbavancin|Dalbavancin
C1642585|T201|COMP|41740-2|LNC|Tazobactam|Tazobactam
C1642586|T201|COMP|41750-1|LNC|COCH gene targeted mutation analysis|COCH gene targeted mutation analysis
C1642587|T201|COMP|41752-7|LNC|Ehrlichia chaffeensis Ab|Ehrlichia chaffeensis Ab
C1642588|T201|COMP|41758-4|LNC|GNAS1 gene targeted mutation analysis|GNAS1 gene targeted mutation analysis
C1642589|T201|COMP|41763-4|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C1642590|T201|COMP|41767-5|LNC|Triamcinolone acetonide|Triamcinolone acetonide
C1643172|T201|COMP|41433-4|LNC|Cryptosporidium hominis DNA|Cryptosporidium hominis DNA
C1643173|T201|COMP|41441-7|LNC|Encephalitozoon intestinalis DNA|Encephalitozoon intestinalis DNA
C1643174|T201|COMP|41451-6|LNC|Plasmodium stage|Plasmodium stage
C1643175|T201|COMP|41455-7|LNC|Human metapneumovirus genotype|Human metapneumovirus genotype
C1643176|T201|COMP|41456-5|LNC|Respiratory syncytial virus genotype|Respiratory syncytial virus genotype
C1643177|T201|COMP|41457-3|LNC|Rhinovirus serotype|Rhinovirus serotype
C1643178|T201|COMP|41459-9|LNC|SARS coronavirus|SARS coronavirus
C1643179|T201|COMP|41460-7|LNC|SARS coronavirus Ab.IgG|SARS coronavirus Ab.IgG
C1643180|T201|COMP|41466-4|LNC|Methadone/Creatinine|Methadone/Creatinine
C1643181|T201|COMP|41468-0|LNC|Barbiturates/Creatinine|Barbiturates/Creatinine
C1643182|T201|COMP|41471-4|LNC|Phenethicillin|Phenethicillin
C1643183|T201|COMP|41472-2|LNC|carBAMazepine|carBAMazepine
C1643184|T201|COMP|41480-5|LNC|BK virus DNA|BK virus DNA
C1643185|T201|COMP|41481-3|LNC|Blastomyces sp Ab|Blastomyces sp Ab
C1643186|T201|COMP|41483-9|LNC|Clostridium tetani toxoid Ab|Clostridium tetani toxoid Ab
C1643187|T201|COMP|41488-8|LNC|Cryptosporidium sp|Cryptosporidium sp
C1643188|T201|COMP|41492-0|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C1643189|T201|COMP|42608-0|LNC|Cells.CD10+CD20+/100 cells|Cells.CD10+CD20+/100 cells
C1643190|T201|COMP|42612-2|LNC|Salicylurate|Salicylurate
C1643191|T201|COMP|42617-1|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1643192|T201|COMP|42622-1|LNC|Cells.CD13+CD56+/100 cells|Cells.CD13+CD56+/100 cells
C1643193|T201|COMP|42626-2|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1643194|T201|COMP|42630-4|LNC|Cannabinoids|Cannabinoids
C1643196|T201|COMP|42638-7|LNC|Coagulation tissue factor induced|Coagulation tissue factor induced
C1643197|T201|COMP|42641-1|LNC|Babesia sp DNA|Babesia sp DNA
C1643198|T201|COMP|42647-8|LNC|Ethionamide 10.0 ug/mL|Ethionamide 10.0 ug/mL
C1643199|T201|COMP|42649-4|LNC|Isoniazid 0.2 ug/mL|Isoniazid 0.2 ug/mL
C1643200|T201|COMP|42654-4|LNC|Para aminosalicylate 2.0 ug/mL|Para aminosalicylate 2.0 ug/mL
C1643201|T201|COMP|42657-7|LNC|rifAMPin 1.0 ug/mL|rifAMPin 1.0 ug/mL
C1643202|T201|COMP|42658-5|LNC|Streptomycin 10.0 ug/mL|Streptomycin 10.0 ug/mL
C1643203|T201|COMP|42661-9|LNC|Bacteria identified|Bacteria identified
C1643204|T201|COMP|42664-3|LNC|HLA-Cw|HLA-Cw
C1643205|T201|COMP|42665-0|LNC|Dantron|Dantron
C1643206|T201|COMP|41292-4|LNC|Soluble mesothelin related proteins|Soluble mesothelin related proteins
C1643208|T201|COMP|41439-1|LNC|Encephalitozoon cuniculi DNA|Encephalitozoon cuniculi DNA
C1643225|T201|COMP|41506-7|LNC|Polio virus Ab panel|Polio virus Ab panel
C1643226|T201|COMP|41508-3|LNC|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C1643227|T201|COMP|41515-8|LNC|HIV 1 RNA|HIV 1 RNA
C1643228|T201|COMP|41616-4|LNC|Platelet Ab|Platelet Ab
C1643229|T201|COMP|41620-6|LNC|Xylose^5H post 5 g xylose PO|Xylose^5H post 5 g xylose PO
C1643230|T201|COMP|41629-7|LNC|Burkholderia sp DNA|Burkholderia sp DNA
C1643231|T201|COMP|41632-1|LNC|Clostridium botulinum toxin B|Clostridium botulinum toxin B
C1643232|T201|COMP|41637-0|LNC|Ebola virus Ag|Ebola virus Ag
C1643233|T201|COMP|41651-1|LNC|Glucose|Glucose
C1643234|T201|COMP|41727-9|LNC|Aztreonam+Clavulanate|Aztreonam+Clavulanate
C1643235|T201|COMP|41731-1|LNC|Cefpodoxime+Clavulanate|Cefpodoxime+Clavulanate
C1643236|T201|COMP|41738-6|LNC|Rosamicin|Rosamicin
C1643238|T201|COMP|41746-9|LNC|Blastomyces dermatitidis Ag|Blastomyces dermatitidis Ag
C1643239|T201|COMP|41751-9|LNC|COL3A1 gene targeted mutation analysis|COL3A1 gene targeted mutation analysis
C1643240|T201|COMP|41755-0|LNC|Flunisolide|Flunisolide
C1643241|T201|COMP|41756-8|LNC|Fluorometholone|Fluorometholone
C1643580|T201|COMP|41617-2|LNC|Neutrophil Ab|Neutrophil Ab
C1643581|T201|COMP|41622-2|LNC|Bacillus anthracis DNA|Bacillus anthracis DNA
C1643582|T201|COMP|41631-3|LNC|Clostridium botulinum toxin A botA gene|Clostridium botulinum toxin A botA gene
C1643583|T201|COMP|41649-5|LNC|Chloride|Chloride
C1643584|T201|COMP|41663-6|LNC|Aztreonam+Clavulanate|Aztreonam+Clavulanate
C1643585|T201|COMP|41666-9|LNC|Biapenem|Biapenem
C1643586|T201|COMP|41667-7|LNC|Biapenem|Biapenem
C1643587|T201|COMP|41674-3|LNC|cefoTEtan+Clavulanate|cefoTEtan+Clavulanate
C1643588|T201|COMP|41690-9|LNC|Dalbavancin|Dalbavancin
C1643589|T201|COMP|41698-2|LNC|Josamycine|Josamycine
C1643590|T201|COMP|41707-1|LNC|Oritavancin|Oritavancin
C1643591|T201|COMP|41712-1|LNC|Ramoplanin|Ramoplanin
C1643592|T201|COMP|41713-9|LNC|Rosamicin|Rosamicin
C1643593|T201|COMP|41714-7|LNC|Rosamicin|Rosamicin
C1643594|T201|COMP|41716-2|LNC|Sulbactam|Sulbactam
C1643595|T201|COMP|41719-6|LNC|Tazobactam|Tazobactam
C1643601|T201|COMP|41839-2|LNC|Burkholderia pseudomallei Ab.IgG & IgM panel|Burkholderia pseudomallei Ab.IgG & IgM panel
C1643602|T201|COMP|41840-0|LNC|Coxiella burnetii phase 1 & 2 Ab.IgG panel|Coxiella burnetii phase 1 & 2 Ab.IgG panel
C1643603|T201|COMP|41849-1|LNC|Curry Ab.IgG|Curry Ab.IgG
C1643604|T201|COMP|41851-7|LNC|Thymus vulgaris Ab.IgG|Thymus vulgaris Ab.IgG
C1643605|T201|COMP|41853-3|LNC|Orthopoxvirus DNA|Orthopoxvirus DNA
C1643606|T201|COMP|41865-7|LNC|Yeast.hyphae|Yeast.hyphae
C1643607|T201|COMP|41871-5|LNC|Voltage-gated potassium channel Ab|Voltage-gated potassium channel Ab
C1643610|T201|COMP|41877-2|LNC|Bordetella pertussis Ab.IgA & IgG & IgM panel|Bordetella pertussis Ab.IgA & IgG & IgM panel
C1644135|T201|COMP|41614-9|LNC|Tube number|Tube number
C1644136|T201|COMP|41627-1|LNC|Burkholderia sp Ag|Burkholderia sp Ag
C1644137|T201|COMP|41662-8|LNC|Aztreonam+Clavulanate|Aztreonam+Clavulanate
C1644138|T201|COMP|41665-1|LNC|Biapenem|Biapenem
C1644139|T201|COMP|41670-1|LNC|ceFAZolin|ceFAZolin
C1644140|T201|COMP|41678-4|LNC|Cefpodoxime+Clavulanate|Cefpodoxime+Clavulanate
C1644141|T201|COMP|41684-2|LNC|Cephaloridine|Cephaloridine
C1644142|T201|COMP|41686-7|LNC|Clavulanate|Clavulanate
C1644143|T201|COMP|41696-6|LNC|Everninomicin|Everninomicin
C1644144|T201|COMP|41704-8|LNC|Nafcillin|Nafcillin
C1644145|T201|COMP|41710-5|LNC|Ramoplanin|Ramoplanin
C1644146|T201|COMP|41720-4|LNC|Tazobactam|Tazobactam
C1644157|T201|COMP|41848-3|LNC|Capsicum annuum Ab.IgG|Capsicum annuum Ab.IgG
C1644158|T201|COMP|41852-5|LNC|Microorganism or agent identified|Microorganism or agent identified
C1644159|T201|COMP|41855-8|LNC|Staphylococcus aureus enterotoxin B|Staphylococcus aureus enterotoxin B
C1644160|T201|COMP|41859-0|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C1644161|T201|COMP|41860-8|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C1644162|T201|COMP|41868-1|LNC|Waxy casts|Waxy casts
C1644163|T201|COMP|41870-7|LNC|Tryptase.mature|Tryptase.mature
C1644164|T201|COMP|41873-1|LNC|Alnus rugosa Ab.IgG|Alnus rugosa Ab.IgG
C1644165|T201|COMP|42182-6|LNC|Gossypol.bound|Gossypol.bound
C1644166|T201|COMP|42220-4|LNC|Chromium/Creatinine|Chromium/Creatinine
C1644167|T201|COMP|42235-2|LNC|Benzodiazepine metabolites|Benzodiazepine metabolites
C1644626|T201|COMP|41516-6|LNC|HIV 1 RNA|HIV 1 RNA
C1644627|T201|COMP|41604-0|LNC|Glucose^post CFst|Glucose^post CFst
C1644628|T201|COMP|41621-4|LNC|Arenavirus RNA|Arenavirus RNA
C1644629|T201|COMP|41626-3|LNC|Brucella sp DNA|Brucella sp DNA
C1644630|T201|COMP|42669-2|LNC|Fatty acids|Fatty acids
C1644632|T201|COMP|42722-9|LNC|OmpC Ab|OmpC Ab
C1644633|T201|COMP|42723-7|LNC|OmpC Ab|OmpC Ab
C1644634|T201|COMP|41668-5|LNC|Carbenicillin|Carbenicillin
C1644635|T201|COMP|41671-9|LNC|Cefotaxime+Clavulanate|Cefotaxime+Clavulanate
C1644636|T201|COMP|41679-2|LNC|Cefpodoxime+Clavulanate|Cefpodoxime+Clavulanate
C1644637|T201|COMP|41681-8|LNC|cefTRIAXone+Clavulanate|cefTRIAXone+Clavulanate
C1644638|T201|COMP|41689-1|LNC|Dalbavancin|Dalbavancin
C1644639|T201|COMP|41691-7|LNC|DAPTOmycin|DAPTOmycin
C1644640|T201|COMP|41693-3|LNC|Ethionamide|Ethionamide
C1644641|T201|COMP|41702-2|LNC|Mezlocillin|Mezlocillin
C1644642|T201|COMP|41711-3|LNC|Ramoplanin|Ramoplanin
C1644643|T201|COMP|41721-2|LNC|Tazobactam|Tazobactam
C1644649|T201|COMP|41842-6|LNC|Herpes virus 7 Ab.IgG & IgM panel|Herpes virus 7 Ab.IgG & IgM panel
C1644651|T201|COMP|41864-0|LNC|Yeast.hyphae|Yeast.hyphae
C1644652|T201|COMP|41866-5|LNC|von Willebrand factor Ag actual/Normal|von Willebrand factor Ag actual/Normal
C1644653|T201|COMP|41867-3|LNC|von Willebrand factor Ag|von Willebrand factor Ag
C1644654|T201|COMP|41869-9|LNC|Testosterone.bioavailable+Free/Testosterone.total|Testosterone.bioavailable+Free/Testosterone.total
C1644655|T201|COMP|41878-0|LNC|Dengue virus Ab.IgG & IgM panel|Dengue virus Ab.IgG & IgM panel
C1644656|T201|COMP|41898-8|LNC|Vendor device model code|Vendor device model code
C1644660|T201|COMP|42194-1|LNC|Cells.CD4/100 cells|Cells.CD4/100 cells
C1644661|T201|COMP|42199-0|LNC|Soluble liver Ab|Soluble liver Ab
C1645294|T201|COMP|41601-6|LNC|Bacteria|Bacteria
C1645295|T201|COMP|41609-9|LNC|Prolactin^1H post XXX challenge|Prolactin^1H post XXX challenge
C1645296|T201|COMP|41635-4|LNC|Clostridium botulinum toxin F|Clostridium botulinum toxin F
C1645297|T201|COMP|41656-0|LNC|Potassium|Potassium
C1645298|T201|COMP|41658-6|LNC|ABT492|ABT492
C1645299|T201|COMP|41659-4|LNC|ABT492|ABT492
C1645300|T201|COMP|41660-2|LNC|ABT492|ABT492
C1645301|T201|COMP|41661-0|LNC|Azlocillin|Azlocillin
C1645302|T201|COMP|41664-4|LNC|Aztreonam+Clavulanate|Aztreonam+Clavulanate
C1645303|T201|COMP|41669-3|LNC|Cefamandole|Cefamandole
C1645304|T201|COMP|41673-5|LNC|cefoTEtan+Clavulanate|cefoTEtan+Clavulanate
C1645305|T201|COMP|41682-6|LNC|cefTRIAXone+Clavulanate|cefTRIAXone+Clavulanate
C1645306|T201|COMP|41685-9|LNC|Clavulanate|Clavulanate
C1645307|T201|COMP|41695-8|LNC|Everninomicin|Everninomicin
C1645308|T201|COMP|41701-4|LNC|Lomefloxacin|Lomefloxacin
C1645309|T201|COMP|41703-0|LNC|Moxalactam|Moxalactam
C1645310|T201|COMP|41706-3|LNC|Novobiocin|Novobiocin
C1645311|T201|COMP|41709-7|LNC|Oritavancin|Oritavancin
C1645312|T201|COMP|41715-4|LNC|Rosamicin|Rosamicin
C1645320|T201|COMP|41854-1|LNC|Ricinus communis DNA|Ricinus communis DNA
C1645321|T201|COMP|41858-2|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C1645322|T201|COMP|41861-6|LNC|Yeast.hyphae|Yeast.hyphae
C1645323|T201|COMP|41872-3|LNC|PDCD10 gene targeted mutation analysis|PDCD10 gene targeted mutation analysis
C1645324|T201|COMP|41874-9|LNC|Betula populifolia Ab.IgE|Betula populifolia Ab.IgE
C1645326|T201|COMP|42215-4|LNC|Erythrocytes.nucleated/100 cells|Erythrocytes.nucleated/100 cells
C1645327|T201|COMP|42226-1|LNC|Thallium/Creatinine|Thallium/Creatinine
C1645723|T201|COMP|41653-7|LNC|Glucose|Glucose
C1645724|T201|COMP|41676-8|LNC|cefOXitin+Clavulanate|cefOXitin+Clavulanate
C1645725|T201|COMP|41677-6|LNC|cefOXitin+Clavulanate|cefOXitin+Clavulanate
C1645726|T201|COMP|41680-0|LNC|Cefpodoxime+Clavulanate|Cefpodoxime+Clavulanate
C1645727|T201|COMP|41697-4|LNC|Gemifloxacin|Gemifloxacin
C1645728|T201|COMP|41700-6|LNC|Lincomycin|Lincomycin
C1645729|T201|COMP|41708-9|LNC|Oritavancin|Oritavancin
C1645730|T201|COMP|42327-7|LNC|Leukocytes|Leukocytes
C1645731|T201|COMP|42332-7|LNC|Alpha-1-Fetoprotein.L3/Alpha-1-Fetoprotein.total|Alpha-1-Fetoprotein.L3/Alpha-1-Fetoprotein.total
C1645733|T201|COMP|42496-0|LNC|Echinococcus sp Ab|Echinococcus sp Ab
C1645734|T201|COMP|42527-2|LNC|Parietal cell Ab|Parietal cell Ab
C1645735|T201|COMP|42584-3|LNC|Beet Ab.IgG|Beet Ab.IgG
C1645736|T201|COMP|42607-2|LNC|Prolactin.monomeric|Prolactin.monomeric
C1645737|T201|COMP|42977-9|LNC|Porcine influenza virus A Ab|Porcine influenza virus A Ab
C1645738|T201|COMP|41748-5|LNC|CAPN3 gene targeted mutation analysis|CAPN3 gene targeted mutation analysis
C1645739|T201|COMP|41761-8|LNC|lamoTRIgine|lamoTRIgine
C1645740|T201|COMP|41765-9|LNC|SCN1A gene targeted mutation analysis|SCN1A gene targeted mutation analysis
C1646205|T201|COMP|41675-0|LNC|cefOXitin+Clavulanate|cefOXitin+Clavulanate
C1646206|T201|COMP|42751-8|LNC|Phosphatidylserine Ab.IgA.B2GP1 dependent|Phosphatidylserine Ab.IgA.B2GP1 dependent
C1646207|T201|COMP|42777-3|LNC|AKT1 gene targeted mutation analysis|AKT1 gene targeted mutation analysis
C1646208|T201|COMP|42778-1|LNC|BRCA1 Ag|BRCA1 Ag
C1646314|T201|COMP|42973-8|LNC|Powassan virus Ab.IgG|Powassan virus Ab.IgG
C1646315|T201|COMP|42364-0|LNC|Streptococcus pneumoniae 6 serotypes Ab.IgG panel|Streptococcus pneumoniae 6 serotypes Ab.IgG panel
C1646318|T201|COMP|42583-5|LNC|Bean string Ab.IgE.RAST class|Bean string Ab.IgE.RAST class
C1646319|T201|COMP|42594-2|LNC|Fraxinus americana Ab.IgE/IgE.total|Fraxinus americana Ab.IgE/IgE.total
C1646320|T201|COMP|42605-6|LNC|Dialysis bag number|Dialysis bag number
C1646321|T201|COMP|42619-7|LNC|Cells.CD28/100 cells|Cells.CD28/100 cells
C1646322|T201|COMP|42640-3|LNC|Urease^1D post incubation|Urease^1D post incubation
C1646323|T201|COMP|42645-2|LNC|Ethambutol 10.0 ug/mL|Ethambutol 10.0 ug/mL
C1646324|T201|COMP|42668-4|LNC|Fatty acids|Fatty acids
C1646325|T201|COMP|42917-5|LNC|HIV 1 RNA|HIV 1 RNA
C1646327|T201|COMP|41749-3|LNC|CHIC2 gene targeted mutation analysis|CHIC2 gene targeted mutation analysis
C1646328|T201|COMP|41757-6|LNC|Fluticasone propionate|Fluticasone propionate
C1646768|T201|COMP|41657-8|LNC|Sodium|Sodium
C1646769|T201|COMP|41692-5|LNC|Enoxacin|Enoxacin
C1646770|T201|COMP|41705-5|LNC|Neomycin|Neomycin
C1646771|T201|COMP|42740-1|LNC|Phosphatidylcholine Ab.IgA.B2GP1 independent|Phosphatidylcholine Ab.IgA.B2GP1 independent
C1646772|T201|COMP|42757-5|LNC|Troponin I.cardiac|Troponin I.cardiac
C1646774|T201|COMP|42497-8|LNC|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C1646775|T201|COMP|42589-2|LNC|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C1646776|T201|COMP|42901-9|LNC|Dihydrocodeine|Dihydrocodeine
C1646777|T201|COMP|42959-7|LNC|Salmonella typhi O Ab|Salmonella typhi O Ab
C1646778|T201|COMP|41393-0|LNC|Collection date|Collection date
C1646779|T201|COMP|41741-0|LNC|Bacteria identified|Bacteria identified
C1646780|T201|COMP|41753-5|LNC|FKRP gene targeted mutation analysis|FKRP gene targeted mutation analysis
C1646781|T201|COMP|41760-0|LNC|Interleukin 12|Interleukin 12
C1647447|T201|COMP|41688-3|LNC|Dalbavancin|Dalbavancin
C1647448|T201|COMP|41699-0|LNC|Josamycine|Josamycine
C1647449|T201|COMP|42785-6|LNC|FGFR1 gene targeted mutation analysis|FGFR1 gene targeted mutation analysis
C1647450|T201|COMP|42375-6|LNC|Neisseria meningitidis serogroup Z Ag|Neisseria meningitidis serogroup Z Ag
C1647451|T201|COMP|42532-2|LNC|Thermoactinomyces candidus Ab|Thermoactinomyces candidus Ab
C1647452|T201|COMP|42535-5|LNC|Tipranavir|Tipranavir
C1647453|T201|COMP|42615-5|LNC|Glucose^30M post dose lactose PO|Glucose^30M post dose lactose PO
C1647454|T201|COMP|42627-0|LNC|HIV 1 Ab|HIV 1 Ab
C1647455|T201|COMP|42655-1|LNC|Rifabutin 0.5 ug/mL|Rifabutin 0.5 ug/mL
C1647456|T201|COMP|42981-1|LNC|Polio virus 1 Ab|Polio virus 1 Ab
C1647457|T201|COMP|41768-3|LNC|VWF gene targeted mutation analysis|VWF gene targeted mutation analysis
C1647458|T201|COMP|41769-1|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C1647880|T201|COMP|41718-8|LNC|Sulbactam|Sulbactam
C1647881|T201|COMP|41745-1|LNC|Betamethasone|Betamethasone
C1647883|T201|COMP|42895-3|LNC|Colorado tick fever virus Ab.IgG|Colorado tick fever virus Ab.IgG
C1647884|T201|COMP|43016-5|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C1647885|T201|COMP|43067-8|LNC|Candida sp Ab|Candida sp Ab
C1647886|T201|COMP|43070-2|LNC|Burkholderia pseudomallei Ab.IgG|Burkholderia pseudomallei Ab.IgG
C1647893|T201|COMP|22561-5|LNC|Streptococcus pneumoniae 9n Ab^2nd specimen|Streptococcus pneumoniae 9n Ab^2nd specimen
C1648316|T201|COMP|42507-4|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C1648358|T201|COMP|41430-0|LNC|Angiostrongylus cantonensis DNA|Angiostrongylus cantonensis DNA
C1648838|T201|COMP|41474-8|LNC|Diethylcarbamazepine|Diethylcarbamazepine
C1648839|T201|COMP|41857-4|LNC|Vibrio parahaemolyticus DNA|Vibrio parahaemolyticus DNA
C1648935|T201|COMP|41717-0|LNC|Sulbactam|Sulbactam
C1648936|T201|COMP|41723-8|LNC|Thiamphenicol|Thiamphenicol
C1648939|T201|COMP|42861-5|LNC|Carbaryl|Carbaryl
C1648940|T201|COMP|42883-9|LNC|Cells.CD52/100 cells|Cells.CD52/100 cells
C1648941|T201|COMP|42890-4|LNC|Cells.myeloperoxidase/100 cells|Cells.myeloperoxidase/100 cells
C1648953|T201|COMP|41847-5|LNC|Armoracia rusticana Ab.IgG|Armoracia rusticana Ab.IgG
C1648954|T201|COMP|41850-9|LNC|Lidocaine Ab.IgE|Lidocaine Ab.IgE
C1649472|T201|COMP|43064-5|LNC|Chikungunya virus Ab|Chikungunya virus Ab
C1649478|T201|COMP|41407-8|LNC|Cortisol^pre dose corticotropin|Cortisol^pre dose corticotropin
C1649479|T201|COMP|41415-1|LNC|Babesia duncani Ab|Babesia duncani Ab
C1650343|T201|COMP|43018-1|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C1650493|T201|COMP|42204-8|LNC|Hairy cells/100 leukocytes|Hairy cells/100 leukocytes
C1650896|T201|COMP|42371-5|LNC|Neisseria meningitidis serogroup C Ag|Neisseria meningitidis serogroup C Ag
C1651089|T201|COMP|42962-1|LNC|Salmonella paratyphi C O Ab|Salmonella paratyphi C O Ab
C1651090|T201|COMP|42970-4|LNC|Pseudallescheria boydii Ab.IgG|Pseudallescheria boydii Ab.IgG
C1651491|T201|COMP|41645-3|LNC|Calcium.ionized|Calcium.ionized
C1651657|T201|COMP|42922-5|LNC|Ketamine|Ketamine
C1651672|T201|COMP|41863-2|LNC|Yeast.pseudohyphae|Yeast.pseudohyphae
C1651680|T201|COMP|42181-8|LNC|Myocardium Ab|Myocardium Ab
C1652145|T201|COMP|42251-9|LNC|Methadone+Metabolite|Methadone+Metabolite
C1652657|T201|COMP|41639-6|LNC|Ricin toxin Ab.IgM|Ricin toxin Ab.IgM
C1652658|T201|COMP|42816-9|LNC|Stachybotrys chartarum Ab.IgG|Stachybotrys chartarum Ab.IgG
C1652660|T201|COMP|42642-9|LNC|Amikacin 2.0 ug/mL|Amikacin 2.0 ug/mL
C1652983|T201|COMP|43035-5|LNC|Feline immunodeficiency virus Ab|Feline immunodeficiency virus Ab
C1652984|T201|COMP|43057-9|LNC|Chlamydophila psittaci Ab.IgM|Chlamydophila psittaci Ab.IgM
C1652985|T201|COMP|41683-4|LNC|cefTRIAXone+Clavulanate|cefTRIAXone+Clavulanate
C1652986|T201|COMP|41694-1|LNC|Everninomicin|Everninomicin
C1652988|T201|COMP|41672-7|LNC|cefoTEtan+Clavulanate|cefoTEtan+Clavulanate
C1652992|T201|COMP|42636-1|LNC|Urease^3H post incubation|Urease^3H post incubation
C1653514|T201|COMP|17636-2|LNC|Streptococcus pneumoniae 6b Ab^1st specimen|Streptococcus pneumoniae 6b Ab^1st specimen
C1653515|T201|COMP|41743-6|LNC|BBS1 gene targeted mutation analysis|BBS1 gene targeted mutation analysis
C1653519|T201|COMP|42241-0|LNC|Cocaine+Benzoylecgonine|Cocaine+Benzoylecgonine
C1654323|T201|COMP|41990-3|LNC|Parainfluenza virus 4 Ab.IgG|Parainfluenza virus 4 Ab.IgG
C1654324|T201|COMP|41991-1|LNC|SARS coronavirus Ab.IgM|SARS coronavirus Ab.IgM
C1654325|T201|COMP|42599-1|LNC|Corticotropin^1H post XXX challenge|Corticotropin^1H post XXX challenge
C1654326|T201|COMP|42650-2|LNC|Isoniazid 1.0 ug/mL|Isoniazid 1.0 ug/mL
C1654330|T201|COMP|42932-4|LNC|Cells.CD40/100 cells|Cells.CD40/100 cells
C1654331|T201|COMP|41726-1|LNC|ABT492|ABT492
C1655382|T201|COMP|42725-2|LNC|Bromide|Bromide
C1657622|T201|COMP|42592-6|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C1704252|T201|COMP|6028-3|LNC|Parrot australian droppings Ab.IgE|Parrot australian droppings Ab.IgE
C1704283|T201|COMP|13095-5|LNC|Monosialoganglioside GM1 Ab.IgA|Monosialoganglioside GM1 Ab.IgA
C1704284|T201|COMP|13124-3|LNC|Sulfate-3-Glucuronyl paragloboside Ab|Sulfate-3-Glucuronyl paragloboside Ab
C1704286|T201|COMP|13109-4|LNC|Disialylganglioside GD1b Ab|Disialylganglioside GD1b Ab
C1704287|T201|COMP|13113-6|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C1704288|T201|COMP|13108-6|LNC|Tetrasialylganglioside GQ1b Ab|Tetrasialylganglioside GQ1b Ab
C1704357|T201|COMP|13122-7|LNC|Sulfatide Ab.IgM|Sulfatide Ab.IgM
C1704395|T201|COMP|45349-8|LNC|Condition of tick|Condition of tick
C1705870|T201|COMP|43191-6|LNC|FANCC gene targeted mutation analysis|FANCC gene targeted mutation analysis
C1705906|T201|COMP|45191-4|LNC|CAPN3 gene targeted mutation analysis|CAPN3 gene targeted mutation analysis
C1706065|T201|COMP|43268-2|LNC|Cells.CD3-CD57+/100 cells|Cells.CD3-CD57+/100 cells
C1706300|T201|COMP|44290-5|LNC|Adenovirus Ab|Adenovirus Ab
C1706356|T201|COMP|44421-6|LNC|PKD1 gene+PKD2 gene targeted mutation analysis|PKD1 gene+PKD2 gene targeted mutation analysis
C1706361|T201|COMP|46207-7|LNC|PKD1 gene+PKD2 gene targeted mutation analysis|PKD1 gene+PKD2 gene targeted mutation analysis
C1706521|T201|COMP|45078-3|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1706522|T201|COMP|45082-5|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1706523|T201|COMP|45077-5|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1706524|T201|COMP|45080-9|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1706525|T201|COMP|45083-3|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1706557|T201|COMP|45079-1|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1706558|T201|COMP|45081-7|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1706580|T201|COMP|43812-7|LNC|Influenza virus A Ab|Influenza virus A Ab
C1706581|T201|COMP|44091-7|LNC|Influenza virus A hemagglutinin H5 RNA|Influenza virus A hemagglutinin H5 RNA
C1706594|T201|COMP|44937-1|LNC|Thyrotropin^pre dose TRH IV|Thyrotropin^pre dose TRH IV
C1714476|T201|COMP|43270-8|LNC|Ceftobiprole|Ceftobiprole
C1714477|T201|COMP|43271-6|LNC|Ceftobiprole|Ceftobiprole
C1714478|T201|COMP|43272-4|LNC|Ceftobiprole|Ceftobiprole
C1714479|T201|COMP|43273-2|LNC|Cells.CD19+CD27+IgD+/100 cells|Cells.CD19+CD27+IgD+/100 cells
C1714480|T201|COMP|43274-0|LNC|Cells.CD1c+CD22+/100 cells|Cells.CD1c+CD22+/100 cells
C1714481|T201|COMP|43275-7|LNC|Cells.CD3/Cells.CD4|Cells.CD3/Cells.CD4
C1714482|T201|COMP|43276-5|LNC|Dermatophagoides sp Ab.IgE.RAST class|Dermatophagoides sp Ab.IgE.RAST class
C1714483|T201|COMP|43277-3|LNC|GDAP1 gene targeted mutation analysis|GDAP1 gene targeted mutation analysis
C1714484|T201|COMP|43278-1|LNC|Glucose^2H post meal|Glucose^2H post meal
C1714485|T201|COMP|43279-9|LNC|Hepatitis B virus YMDD mutation|Hepatitis B virus YMDD mutation
C1714486|T201|COMP|43280-7|LNC|Hepatitis D virus Ag|Hepatitis D virus Ag
C1714487|T201|COMP|43575-0|LNC|Complement C3|Complement C3
C1714488|T201|COMP|43576-8|LNC|Acylcarnitine/Carnitine.free (C0)|Acylcarnitine/Carnitine.free (C0)
C1714489|T201|COMP|43577-6|LNC|Histamine/Creatinine|Histamine/Creatinine
C1714490|T201|COMP|43578-4|LNC|Complement C3|Complement C3
C1714491|T201|COMP|43579-2|LNC|Complement C3|Complement C3
C1714492|T201|COMP|43580-0|LNC|Complement C4|Complement C4
C1714493|T201|COMP|43581-8|LNC|Complement C4|Complement C4
C1714494|T201|COMP|43582-6|LNC|Complement C4|Complement C4
C1714502|T201|COMP|43752-5|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C1714503|T201|COMP|43753-3|LNC|Spermatozoa IgM binding location|Spermatozoa IgM binding location
C1714504|T201|COMP|43754-1|LNC|Sulfate|Sulfate
C1714505|T201|COMP|43755-8|LNC|Casts|Casts
C1714509|T201|COMP|43921-6|LNC|Bartonella sp Ab.IgM|Bartonella sp Ab.IgM
C1714510|T201|COMP|43922-4|LNC|Beta endorphin|Beta endorphin
C1714511|T201|COMP|43923-2|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C1714512|T201|COMP|43924-0|LNC|azaTHIOprine|azaTHIOprine
C1714513|T201|COMP|43925-7|LNC|Bordetella parapertussis|Bordetella parapertussis
C1714514|T201|COMP|43926-5|LNC|Babesia sp Ab|Babesia sp Ab
C1714515|T201|COMP|43927-3|LNC|Arginine|Arginine
C1714516|T201|COMP|43928-1|LNC|Coxiella burnetii phase 2 Ab.IgM|Coxiella burnetii phase 2 Ab.IgM
C1714517|T201|COMP|43929-9|LNC|Anthraquinone|Anthraquinone
C1714518|T201|COMP|43175-9|LNC|Chlamydia trachomatis L2 Ab.IgM|Chlamydia trachomatis L2 Ab.IgM
C1714519|T201|COMP|43177-5|LNC|Phenmetrazine|Phenmetrazine
C1714520|T201|COMP|43178-3|LNC|Phentermine|Phentermine
C1714521|T201|COMP|43179-1|LNC|Asialoganglioside GM1 Ab.IgM|Asialoganglioside GM1 Ab.IgM
C1714522|T201|COMP|43180-9|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C1714523|T201|COMP|43181-7|LNC|Arsenic.organic|Arsenic.organic
C1714524|T201|COMP|43182-5|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C1714525|T201|COMP|43183-3|LNC|Cyanide|Cyanide
C1714531|T201|COMP|43739-2|LNC|Blood group Ag|Blood group Ag
C1714532|T201|COMP|43740-0|LNC|Glucose/Insulin|Glucose/Insulin
C1714533|T201|COMP|43741-8|LNC|Temperature|Temperature
C1714534|T201|COMP|43742-6|LNC|Time next dose|Time next dose
C1714535|T201|COMP|43743-4|LNC|Lymphocytes.variant|Lymphocytes.variant
C1714536|T201|COMP|43744-2|LNC|COX10 gene targeted mutation analysis|COX10 gene targeted mutation analysis
C1714537|T201|COMP|43822-6|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C1714538|T201|COMP|43823-4|LNC|Aspergillus glaucus Ab|Aspergillus glaucus Ab
C1714539|T201|COMP|43824-2|LNC|Bilirubin|Bilirubin
C1714540|T201|COMP|43825-9|LNC|Arsenic|Arsenic
C1714541|T201|COMP|43827-5|LNC|Barbiturates|Barbiturates
C1714542|T201|COMP|43828-3|LNC|Benzodiazepines|Benzodiazepines
C1714543|T201|COMP|43829-1|LNC|Caffeine|Caffeine
C1714544|T201|COMP|43830-9|LNC|Nicotine|Nicotine
C1714549|T201|COMP|44977-7|LNC|Chlamydophila psittaci Ab.IgM|Chlamydophila psittaci Ab.IgM
C1714550|T201|COMP|44978-5|LNC|Chlamydophila psittaci Ab.IgA|Chlamydophila psittaci Ab.IgA
C1714551|T201|COMP|44979-3|LNC|Chlamydophila pneumoniae Ab^2nd specimen|Chlamydophila pneumoniae Ab^2nd specimen
C1714552|T201|COMP|44980-1|LNC|Chlamydophila pneumoniae Ab^1st specimen|Chlamydophila pneumoniae Ab^1st specimen
C1714553|T201|COMP|44981-9|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C1714554|T201|COMP|43170-0|LNC|Human papilloma virus 31+33 DNA|Human papilloma virus 31+33 DNA
C1714555|T201|COMP|43171-8|LNC|Interleukin 2 receptor|Interleukin 2 receptor
C1714556|T201|COMP|43172-6|LNC|Triiodothyronine Ab|Triiodothyronine Ab
C1714557|T201|COMP|43173-4|LNC|Chlamydia trachomatis L2 Ab.IgG|Chlamydia trachomatis L2 Ab.IgG
C1714558|T201|COMP|43184-1|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C1714559|T201|COMP|43185-8|LNC|HIV 1 & 2 Ab band pattern|HIV 1 & 2 Ab band pattern
C1714560|T201|COMP|43186-6|LNC|Acylcarnitine/Carnitine.free (C0)|Acylcarnitine/Carnitine.free (C0)
C1714561|T201|COMP|43187-4|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C1714562|T201|COMP|43188-2|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C1714563|T201|COMP|43189-0|LNC|Saccharomyces cerevisiae Ab.IgA|Saccharomyces cerevisiae Ab.IgA
C1714564|T201|COMP|43192-4|LNC|Legionella pneumophila 2+3+4+5+6+8 Ab|Legionella pneumophila 2+3+4+5+6+8 Ab
C1714565|T201|COMP|43193-2|LNC|Legionella non pneumophila sp Ab|Legionella non pneumophila sp Ab
C1714566|T201|COMP|43194-0|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C1714567|T201|COMP|43195-7|LNC|Nicotine|Nicotine
C1714568|T201|COMP|43196-5|LNC|Cotinine|Cotinine
C1714569|T201|COMP|43197-3|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C1714570|T201|COMP|43198-1|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C1714571|T201|COMP|43199-9|LNC|Norfentanyl|Norfentanyl
C1714572|T201|COMP|43200-5|LNC|Norfentanyl|Norfentanyl
C1714573|T201|COMP|43201-3|LNC|BK virus DNA|BK virus DNA
C1714574|T201|COMP|43202-1|LNC|Liver kidney microsomal 1 Ab.IgG|Liver kidney microsomal 1 Ab.IgG
C1714575|T201|COMP|43203-9|LNC|Parainfluenza virus 1 Ab|Parainfluenza virus 1 Ab
C1714576|T201|COMP|43205-4|LNC|Parainfluenza virus 3 Ab|Parainfluenza virus 3 Ab
C1714577|T201|COMP|43206-2|LNC|Tetrachloroethylene|Tetrachloroethylene
C1714578|T201|COMP|43207-0|LNC|Invasive trophoblast Ag|Invasive trophoblast Ag
C1714579|T201|COMP|43208-8|LNC|Invasive trophoblast Ag|Invasive trophoblast Ag
C1714582|T201|COMP|43211-2|LNC|Human papilloma virus 6+11+42+43+44 DNA|Human papilloma virus 6+11+42+43+44 DNA
C1714583|T201|COMP|43212-0|LNC|Albumin|Albumin
C1714584|T201|COMP|43213-8|LNC|Polychlorinated biphenyl|Polychlorinated biphenyl
C1714585|T201|COMP|43214-6|LNC|Bacteria identified|Bacteria identified
C1714586|T201|COMP|43215-3|LNC|Cortisol^baseline|Cortisol^baseline
C1714588|T201|COMP|43218-7|LNC|Nicotine+Cotinine|Nicotine+Cotinine
C1714589|T201|COMP|43219-5|LNC|traMADol|traMADol
C1714590|T201|COMP|43220-3|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C1714591|T201|COMP|43222-9|LNC|Potassium/Creatinine|Potassium/Creatinine
C1714592|T201|COMP|43223-7|LNC|Sodium/Creatinine|Sodium/Creatinine
C1714593|T201|COMP|43224-5|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1714594|T201|COMP|43225-2|LNC|Toxocara sp Ab|Toxocara sp Ab
C1714595|T201|COMP|43226-0|LNC|2-Hydroxyisocaproate|2-Hydroxyisocaproate
C1714596|T201|COMP|43227-8|LNC|Ova & parasites identified|Ova & parasites identified
C1714597|T201|COMP|43228-6|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1714598|T201|COMP|43229-4|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1714599|T201|COMP|43230-2|LNC|Benzoylecgonine|Benzoylecgonine
C1714600|T201|COMP|43231-0|LNC|Histone Ab|Histone Ab
C1714601|T201|COMP|43233-6|LNC|OTC gene targeted mutation analysis|OTC gene targeted mutation analysis
C1714602|T201|COMP|43234-4|LNC|Liver kidney microsomal 1 Ab.IgG|Liver kidney microsomal 1 Ab.IgG
C1714603|T201|COMP|43235-1|LNC|Acrylylcarnitine (C3:1)|Acrylylcarnitine (C3:1)
C1714604|T201|COMP|43236-9|LNC|Streptococcus pneumoniae Ab.IgG|Streptococcus pneumoniae Ab.IgG
C1714605|T201|COMP|43237-7|LNC|Thrombopoietin|Thrombopoietin
C1714606|T201|COMP|43238-5|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1714607|T201|COMP|43240-1|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C1714608|T201|COMP|43241-9|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C1714609|T201|COMP|43242-7|LNC|ACADM gene targeted mutation analysis|ACADM gene targeted mutation analysis
C1714610|T201|COMP|43243-5|LNC|Isobutyrylcarnitine (C4)|Isobutyrylcarnitine (C4)
C1714611|T201|COMP|43244-3|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1714612|T201|COMP|43245-0|LNC|Erythrocytes|Erythrocytes
C1714613|T201|COMP|43246-8|LNC|PHOX2B gene targeted mutation analysis|PHOX2B gene targeted mutation analysis
C1714614|T201|COMP|43247-6|LNC|Catecholamines/Creatinine|Catecholamines/Creatinine
C1714615|T201|COMP|43248-4|LNC|EPINEPHrine/Creatinine|EPINEPHrine/Creatinine
C1714616|T201|COMP|43249-2|LNC|X ray dye crystals|X ray dye crystals
C1714617|T201|COMP|43250-0|LNC|Xanthine derivatives|Xanthine derivatives
C1714632|T201|COMP|43265-8|LNC|Benztropine|Benztropine
C1714633|T201|COMP|43267-4|LNC|Uranium.depleted cutoff|Uranium.depleted cutoff
C1714634|T201|COMP|43281-5|LNC|Hepatitis D virus Ag|Hepatitis D virus Ag
C1714635|T201|COMP|43282-3|LNC|Heterophile Ab|Heterophile Ab
C1714636|T201|COMP|43283-1|LNC|Myeloid cells/100 cells|Myeloid cells/100 cells
C1714637|T201|COMP|43284-9|LNC|Spermatozoa IgA binding location|Spermatozoa IgA binding location
C1714638|T201|COMP|43285-6|LNC|Spermatozoa Ab.IgM/100 spermatozoa|Spermatozoa Ab.IgM/100 spermatozoa
C1714639|T201|COMP|43286-4|LNC|Spermatozoa Ab.IgG/100 spermatozoa|Spermatozoa Ab.IgG/100 spermatozoa
C1714640|T201|COMP|43287-2|LNC|Spermatozoa IgG binding location|Spermatozoa IgG binding location
C1714641|T201|COMP|43288-0|LNC|Spermatozoa Ab.IgA/100 spermatozoa|Spermatozoa Ab.IgA/100 spermatozoa
C1714642|T201|COMP|43289-8|LNC|Methylcrotonylcarnitine (C5:1)|Methylcrotonylcarnitine (C5:1)
C1714643|T201|COMP|43290-6|LNC|HLA-DRB1|HLA-DRB1
C1714644|T201|COMP|43291-4|LNC|HLA-DQB1|HLA-DQB1
C1714646|T201|COMP|43293-0|LNC|HTLV I+II p28 Ab|HTLV I+II p28 Ab
C1714647|T201|COMP|43294-8|LNC|HTLV I+II p26 Ab|HTLV I+II p26 Ab
C1714648|T201|COMP|43295-5|LNC|HTLV I+II p53 Ab|HTLV I+II p53 Ab
C1714649|T201|COMP|43297-1|LNC|HTLV I+II p32 Ab|HTLV I+II p32 Ab
C1714650|T201|COMP|43298-9|LNC|HTLV I+II rgp21 Ab|HTLV I+II rgp21 Ab
C1714651|T201|COMP|43299-7|LNC|HTLV I+II p19 Ab|HTLV I+II p19 Ab
C1714652|T201|COMP|43300-3|LNC|HTLV I+II p24 Ab|HTLV I+II p24 Ab
C1714653|T201|COMP|43301-1|LNC|HTLV I+II p36 Ab|HTLV I+II p36 Ab
C1714654|T201|COMP|43302-9|LNC|Platelet glycoprotein Ab|Platelet glycoprotein Ab
C1714655|T201|COMP|43303-7|LNC|Immune complex.C3d|Immune complex.C3d
C1714656|T201|COMP|43304-5|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1714657|T201|COMP|43305-2|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1714658|T201|COMP|43306-0|LNC|Chromosome 21 trisomy|Chromosome 21 trisomy
C1714659|T201|COMP|43307-8|LNC|Bacteria identified|Bacteria identified
C1714660|T201|COMP|43308-6|LNC|Lupus anticoagulant neutralization.buffer|Lupus anticoagulant neutralization.buffer
C1714661|T201|COMP|43309-4|LNC|Desmoglein 1 & Desmoglein 3 Ab panel|Desmoglein 1 & Desmoglein 3 Ab panel
C1714662|T201|COMP|43310-2|LNC|FBN2 gene targeted mutation analysis|FBN2 gene targeted mutation analysis
C1714663|T201|COMP|43311-0|LNC|Desmoglein 1 Ab|Desmoglein 1 Ab
C1714664|T201|COMP|43312-8|LNC|Desmoglein 3 Ab|Desmoglein 3 Ab
C1714665|T201|COMP|43313-6|LNC|Avian adenovirus 127 Ab|Avian adenovirus 127 Ab
C1714666|T201|COMP|43314-4|LNC|Avian paramyxovirus 6 Ab|Avian paramyxovirus 6 Ab
C1714667|T201|COMP|43315-1|LNC|Avian paramyxovirus 7 Ab|Avian paramyxovirus 7 Ab
C1714668|T201|COMP|43316-9|LNC|Avian paramyxovirus 8 Ab|Avian paramyxovirus 8 Ab
C1714669|T201|COMP|43317-7|LNC|Avian paramyxovirus 9 Ab|Avian paramyxovirus 9 Ab
C1714670|T201|COMP|43318-5|LNC|Avian metapneumovirus A Ab|Avian metapneumovirus A Ab
C1714671|T201|COMP|43321-9|LNC|Avian metapneumovirus B Ab|Avian metapneumovirus B Ab
C1714672|T201|COMP|43322-7|LNC|Avian metapneumovirus C Ab|Avian metapneumovirus C Ab
C1714673|T201|COMP|43323-5|LNC|Avian metapneumovirus C Ab|Avian metapneumovirus C Ab
C1714674|T201|COMP|43324-3|LNC|Avian reovirus Ab|Avian reovirus Ab
C1714675|T201|COMP|43325-0|LNC|Chicken anemia virus Ab|Chicken anemia virus Ab
C1714676|T201|COMP|43326-8|LNC|Classical swine fever virus Ab|Classical swine fever virus Ab
C1714677|T201|COMP|43327-6|LNC|Classical swine fever virus Ag|Classical swine fever virus Ag
C1714678|T201|COMP|43328-4|LNC|Duck enteritis virus Ab|Duck enteritis virus Ab
C1714679|T201|COMP|43329-2|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C1714680|T201|COMP|43330-0|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C1714681|T201|COMP|43331-8|LNC|Ehrlichia risticii Ab|Ehrlichia risticii Ab
C1714682|T201|COMP|43332-6|LNC|Equine herpesvirus 1 Ab|Equine herpesvirus 1 Ab
C1714683|T201|COMP|43334-2|LNC|Equine herpesvirus 3 Ab|Equine herpesvirus 3 Ab
C1714684|T201|COMP|43335-9|LNC|Fowl adenovirus 1 Ab|Fowl adenovirus 1 Ab
C1714685|T201|COMP|43336-7|LNC|Goose parvovirus Ab|Goose parvovirus Ab
C1714686|T201|COMP|43337-5|LNC|Goose parvovirus RNA|Goose parvovirus RNA
C1714687|T201|COMP|43339-1|LNC|Porcine adenovirus Ab|Porcine adenovirus Ab
C1714688|T201|COMP|43340-9|LNC|Psittacid herpesvirus 1 Ab|Psittacid herpesvirus 1 Ab
C1714689|T201|COMP|43341-7|LNC|Venezuelan equine encephalitis virus Ab|Venezuelan equine encephalitis virus Ab
C1714690|T201|COMP|43342-5|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1714691|T201|COMP|43343-3|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C1714692|T201|COMP|43344-1|LNC|Avian adenovirus 127 Ab|Avian adenovirus 127 Ab
C1714693|T201|COMP|43345-8|LNC|Avian paramyxovirus 6 Ab|Avian paramyxovirus 6 Ab
C1714694|T201|COMP|43346-6|LNC|Avian paramyxovirus 7 Ab|Avian paramyxovirus 7 Ab
C1714695|T201|COMP|43347-4|LNC|Avian paramyxovirus 8 Ab|Avian paramyxovirus 8 Ab
C1714696|T201|COMP|43348-2|LNC|Avian paramyxovirus 9 Ab|Avian paramyxovirus 9 Ab
C1714697|T201|COMP|43349-0|LNC|Avian metapneumovirus A Ab|Avian metapneumovirus A Ab
C1714698|T201|COMP|43350-8|LNC|Avian metapneumovirus A Ab|Avian metapneumovirus A Ab
C1714699|T201|COMP|43351-6|LNC|Avian metapneumovirus B Ab|Avian metapneumovirus B Ab
C1714700|T201|COMP|43352-4|LNC|Avian metapneumovirus B Ab|Avian metapneumovirus B Ab
C1714701|T201|COMP|43354-0|LNC|Avian metapneumovirus C Ab|Avian metapneumovirus C Ab
C1714702|T201|COMP|43355-7|LNC|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgG|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgG
C1714703|T201|COMP|43356-5|LNC|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgA|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgA
C1714704|T201|COMP|43357-3|LNC|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgM|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgM
C1714705|T201|COMP|43358-1|LNC|UNC13D gene targeted mutation analysis|UNC13D gene targeted mutation analysis
C1714706|T201|COMP|43359-9|LNC|11-Ketoetiocholanolone|11-Ketoetiocholanolone
C1714707|T201|COMP|43360-7|LNC|Bordetella sp Ag|Bordetella sp Ag
C1714708|T201|COMP|43361-5|LNC|Cardiolipin Ab.IgA|Cardiolipin Ab.IgA
C1714709|T201|COMP|43362-3|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C1714710|T201|COMP|43363-1|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C1714711|T201|COMP|43364-9|LNC|Enterovirus identified|Enterovirus identified
C1714712|T201|COMP|43365-6|LNC|Nocardia sp identified|Nocardia sp identified
C1714713|T201|COMP|43366-4|LNC|Parainfluenza virus Ag|Parainfluenza virus Ag
C1714714|T201|COMP|43367-2|LNC|Trichomonas sp|Trichomonas sp
C1714715|T201|COMP|43368-0|LNC|Microsatellite instability|Microsatellite instability
C1714716|T201|COMP|43369-8|LNC|PlA1 Ab|PlA1 Ab
C1714717|T201|COMP|43370-6|LNC|CFTR gene.p.IVS8 polyT|CFTR gene.p.IVS8 polyT
C1714718|T201|COMP|43371-4|LNC|Salmonella & Shigella sp identified|Salmonella & Shigella sp identified
C1714720|T201|COMP|43374-8|LNC|Parietaria officinalis Ab.IgE.RAST class|Parietaria officinalis Ab.IgE.RAST class
C1714721|T201|COMP|43375-5|LNC|Phoenix dactylifera Ab.IgE.RAST class|Phoenix dactylifera Ab.IgE.RAST class
C1714722|T201|COMP|43376-3|LNC|Spermatozoa.progressive^post washing|Spermatozoa.progressive^post washing
C1714723|T201|COMP|43377-1|LNC|Spermatozoa.progressive^pre washing|Spermatozoa.progressive^pre washing
C1714724|T201|COMP|43378-9|LNC|Spermatozoa.motile^post washing|Spermatozoa.motile^post washing
C1714725|T201|COMP|43379-7|LNC|HLA-DRB3|HLA-DRB3
C1714726|T201|COMP|43380-5|LNC|Coccidioides immitis Ab.IgG|Coccidioides immitis Ab.IgG
C1714727|T201|COMP|43381-3|LNC|Bordetella pertussis Ab|Bordetella pertussis Ab
C1714729|T201|COMP|43383-9|LNC|Neisseria sp identified|Neisseria sp identified
C1714730|T201|COMP|43384-7|LNC|Neisseria sp identified|Neisseria sp identified
C1714731|T201|COMP|43385-4|LNC|Neisseria sp identified|Neisseria sp identified
C1714732|T201|COMP|43386-2|LNC|Neisseria sp identified|Neisseria sp identified
C1714733|T201|COMP|43387-0|LNC|Neisseria sp identified|Neisseria sp identified
C1714734|T201|COMP|43390-4|LNC|Streptococcus sp identified|Streptococcus sp identified
C1714735|T201|COMP|43391-2|LNC|Bacterial vaginosis score|Bacterial vaginosis score
C1714736|T201|COMP|43392-0|LNC|LDL 1|LDL 1
C1714737|T201|COMP|43393-8|LNC|LDL 4|LDL 4
C1714738|T201|COMP|43394-6|LNC|Cholesterol.in LDL.acetylated|Cholesterol.in LDL.acetylated
C1714739|T201|COMP|43395-3|LNC|Cholesterol.in VLDL.acetylated|Cholesterol.in VLDL.acetylated
C1714740|T201|COMP|43396-1|LNC|Cholesterol.non HDL|Cholesterol.non HDL
C1714741|T201|COMP|43398-7|LNC|Gardnerella vaginalis+Prevotella sp morphotypes|Gardnerella vaginalis+Prevotella sp morphotypes
C1714742|T201|COMP|43399-5|LNC|JAK2 gene.p.Val617Phe|JAK2 gene.p.Val617Phe
C1714743|T201|COMP|43400-1|LNC|Lactobacillus sp morphotypes|Lactobacillus sp morphotypes
C1714744|T201|COMP|43401-9|LNC|Cryofibrinogen|Cryofibrinogen
C1714745|T201|COMP|43403-5|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C1714746|T201|COMP|43404-3|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1714747|T201|COMP|43405-0|LNC|Chlamydia trachomatis & Neisseria gonorrhoeae DNA|Chlamydia trachomatis & Neisseria gonorrhoeae DNA
C1714748|T201|COMP|43406-8|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae DNA|Chlamydia trachomatis+Neisseria gonorrhoeae DNA
C1714749|T201|COMP|43407-6|LNC|Bacteria identified|Bacteria identified
C1714750|T201|COMP|43408-4|LNC|Bacteria identified|Bacteria identified
C1714751|T201|COMP|43409-2|LNC|Bacteria identified|Bacteria identified
C1714752|T201|COMP|43411-8|LNC|Bacteria identified|Bacteria identified
C1714753|T201|COMP|43412-6|LNC|Blood product units issued|Blood product units issued
C1714754|T201|COMP|43413-4|LNC|Blood product units requested|Blood product units requested
C1714755|T201|COMP|43414-2|LNC|Blood product units available|Blood product units available
C1714756|T201|COMP|43415-9|LNC|Unidentified cells/100 cells|Unidentified cells/100 cells
C1714757|T201|COMP|43416-7|LNC|Hematocrit|Hematocrit
C1714759|T201|COMP|43419-1|LNC|Tuberculosis reaction wheal^3D post 1 TU ID|Tuberculosis reaction wheal^3D post 1 TU ID
C1714760|T201|COMP|43420-9|LNC|Uranium dose assessment|Uranium dose assessment
C1714761|T201|COMP|43421-7|LNC|Thiopurine methyltransferase|Thiopurine methyltransferase
C1714762|T201|COMP|43422-5|LNC|Rabbit dander Ab.IgE|Rabbit dander Ab.IgE
C1714763|T201|COMP|43423-3|LNC|Sodium urate|Sodium urate
C1714764|T201|COMP|43424-1|LNC|Bartonella sp Ab.IgM|Bartonella sp Ab.IgM
C1714765|T201|COMP|43425-8|LNC|Bartonella sp Ab.IgG|Bartonella sp Ab.IgG
C1714766|T201|COMP|43426-6|LNC|Bacteria identified|Bacteria identified
C1714768|T201|COMP|43428-2|LNC|Bilirubin.microscopic observation|Bilirubin.microscopic observation
C1714769|T201|COMP|43429-0|LNC|Haemophilus influenzae B Ag|Haemophilus influenzae B Ag
C1714770|T201|COMP|43430-8|LNC|Neisseria meningitidis serogroup B Ag|Neisseria meningitidis serogroup B Ag
C1714771|T201|COMP|43431-6|LNC|Escherichia coli K1 Ag|Escherichia coli K1 Ag
C1714772|T201|COMP|43432-4|LNC|Escherichia coli K1 Ag|Escherichia coli K1 Ag
C1714773|T201|COMP|43433-2|LNC|Acylcarnitine panel|Acylcarnitine panel
C1714774|T201|COMP|43434-0|LNC|Bacterial Ag panel|Bacterial Ag panel
C1714780|T201|COMP|43441-5|LNC|Bacteria identified|Bacteria identified
C1714781|T201|COMP|43442-3|LNC|Bacteria identified|Bacteria identified
C1714782|T201|COMP|43443-1|LNC|Bacterial Ag panel|Bacterial Ag panel
C1714828|T201|COMP|43686-5|LNC|Salivary gland Ab.IgA|Salivary gland Ab.IgA
C1714829|T201|COMP|43687-3|LNC|Powassan virus polyvalent E Ab|Powassan virus polyvalent E Ab
C1714830|T201|COMP|43689-9|LNC|HLA-DQ2 & HLA-DQ8|HLA-DQ2 & HLA-DQ8
C1714831|T201|COMP|43690-7|LNC|Triamterene/Total|Triamterene/Total
C1714832|T201|COMP|44318-4|LNC|Insulin porcine Ab|Insulin porcine Ab
C1714833|T201|COMP|44319-2|LNC|Insulin.bound|Insulin.bound
C1714834|T201|COMP|44320-0|LNC|Interferon.alpha|Interferon.alpha
C1714835|T201|COMP|44321-8|LNC|Interleukin 5|Interleukin 5
C1714836|T201|COMP|44322-6|LNC|Interleukin 6|Interleukin 6
C1714837|T201|COMP|44323-4|LNC|Iodine|Iodine
C1714838|T201|COMP|44324-2|LNC|Iodine.inorganic|Iodine.inorganic
C1714839|T201|COMP|44325-9|LNC|Iron|Iron
C1714840|T201|COMP|44326-7|LNC|Iron|Iron
C1714841|T201|COMP|44327-5|LNC|Iron|Iron
C1714842|T201|COMP|44328-3|LNC|Isocitrate|Isocitrate
C1714843|T201|COMP|44329-1|LNC|Isoleucine/Creatinine|Isoleucine/Creatinine
C1714844|T201|COMP|44723-5|LNC|Histiocytes|Histiocytes
C1714845|T201|COMP|44724-3|LNC|HLA-A29|HLA-A29
C1714846|T201|COMP|44725-0|LNC|HLA-B1|HLA-B1
C1714847|T201|COMP|44727-6|LNC|HLA-DP2|HLA-DP2
C1714848|T201|COMP|44728-4|LNC|HLA-DQA1|HLA-DQA1
C1714849|T201|COMP|44729-2|LNC|Progesterone/11-Deoxycorticosterone|Progesterone/11-Deoxycorticosterone
C1714850|T201|COMP|44730-0|LNC|Progesterone/Estradiol|Progesterone/Estradiol
C1714853|T201|COMP|44733-4|LNC|Triglyceride/Cholesterol.in HDL|Triglyceride/Cholesterol.in HDL
C1714854|T201|COMP|44734-2|LNC|Urea nitrogen/Creatinine|Urea nitrogen/Creatinine
C1714855|T201|COMP|44735-9|LNC|Urea nitrogen/Creatinine|Urea nitrogen/Creatinine
C1714856|T201|COMP|44736-7|LNC|Asialoganglioside GM1 Ab|Asialoganglioside GM1 Ab
C1714857|T201|COMP|44737-5|LNC|Asialoganglioside GM1 Ab|Asialoganglioside GM1 Ab
C1714858|T201|COMP|44738-3|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C1714859|T201|COMP|44739-1|LNC|Beta tubulin Ab.IgM|Beta tubulin Ab.IgM
C1714860|T201|COMP|44741-7|LNC|Disialylganglioside GD1b Ab|Disialylganglioside GD1b Ab
C1714861|T201|COMP|44742-5|LNC|Disialylganglioside GD1b Ab.IgG|Disialylganglioside GD1b Ab.IgG
C1714862|T201|COMP|44744-1|LNC|La Crosse virus Ab|La Crosse virus Ab
C1714863|T201|COMP|44745-8|LNC|La Crosse virus Ab|La Crosse virus Ab
C1714864|T201|COMP|44746-6|LNC|La Crosse virus Ab|La Crosse virus Ab
C1714865|T201|COMP|44747-4|LNC|La Crosse virus Ab|La Crosse virus Ab
C1714866|T201|COMP|44949-6|LNC|Borrelia burgdorferi 34kD Ab.IgG|Borrelia burgdorferi 34kD Ab.IgG
C1714888|T201|COMP|44982-7|LNC|Chlamydophila pneumoniae Ab.IgA|Chlamydophila pneumoniae Ab.IgA
C1714889|T201|COMP|44983-5|LNC|Chlamydia trachomatis L2 Ab.IgM|Chlamydia trachomatis L2 Ab.IgM
C1714890|T201|COMP|44984-3|LNC|Chlamydia trachomatis L2 Ab.IgG|Chlamydia trachomatis L2 Ab.IgG
C1714891|T201|COMP|44985-0|LNC|Chlamydia trachomatis L2 Ab.IgA|Chlamydia trachomatis L2 Ab.IgA
C1714892|T201|COMP|44986-8|LNC|Chlamydia trachomatis G+F+K Ab.IgM|Chlamydia trachomatis G+F+K Ab.IgM
C1714893|T201|COMP|44987-6|LNC|Chlamydia trachomatis G+F+K Ab.IgA|Chlamydia trachomatis G+F+K Ab.IgA
C1714894|T201|COMP|44988-4|LNC|Chlamydia trachomatis D+K Ab.IgM|Chlamydia trachomatis D+K Ab.IgM
C1714895|T201|COMP|44990-0|LNC|Chlamydia trachomatis D+K Ab.IgA|Chlamydia trachomatis D+K Ab.IgA
C1714896|T201|COMP|44991-8|LNC|Chlamydia trachomatis C Ab.IgM|Chlamydia trachomatis C Ab.IgM
C1714897|T201|COMP|44992-6|LNC|Chlamydia trachomatis C Ab.IgG|Chlamydia trachomatis C Ab.IgG
C1714898|T201|COMP|44993-4|LNC|Chlamydia trachomatis C Ab.IgA|Chlamydia trachomatis C Ab.IgA
C1714960|T201|COMP|43573-5|LNC|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C1714962|T201|COMP|43584-2|LNC|Bizarre cells|Bizarre cells
C1714963|T201|COMP|43585-9|LNC|TYMP gene targeted mutation analysis|TYMP gene targeted mutation analysis
C1714964|T201|COMP|43586-7|LNC|Yersinia pseudotuberculosis Ab|Yersinia pseudotuberculosis Ab
C1714965|T201|COMP|43587-5|LNC|Vitis vinifera Ab.IgE/IgE.total|Vitis vinifera Ab.IgE/IgE.total
C1714966|T201|COMP|43588-3|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C1714967|T201|COMP|43589-1|LNC|Shigella sp Ab|Shigella sp Ab
C1714968|T201|COMP|43590-9|LNC|Rabies virus Ab|Rabies virus Ab
C1714969|T201|COMP|43592-5|LNC|Prunus domestica Ab.IgE/IgE.total|Prunus domestica Ab.IgE/IgE.total
C1714970|T201|COMP|43593-3|LNC|Plasmodium malariae Ab.IgG|Plasmodium malariae Ab.IgG
C1714971|T201|COMP|43594-1|LNC|Nidus|Nidus
C1714972|T201|COMP|43595-8|LNC|Methadone|Methadone
C1714973|T201|COMP|43596-6|LNC|Malus sylvestris Ab.IgE/IgE.total|Malus sylvestris Ab.IgE/IgE.total
C1714974|T201|COMP|43597-4|LNC|Inner Ear 68kD Ab|Inner Ear 68kD Ab
C1714975|T201|COMP|43598-2|LNC|Indicans|Indicans
C1714976|T201|COMP|43599-0|LNC|HIV 1 Ab|HIV 1 Ab
C1714977|T201|COMP|43600-6|LNC|Ganglioside GD1b Ab.IgM|Ganglioside GD1b Ab.IgM
C1714978|T201|COMP|43601-4|LNC|Ganglioside GD1b Ab.IgG|Ganglioside GD1b Ab.IgG
C1714979|T201|COMP|43602-2|LNC|Echinococcus granulosus Ab|Echinococcus granulosus Ab
C1714980|T201|COMP|43603-0|LNC|Androstenedione^1st specimen post XXX challenge|Androstenedione^1st specimen post XXX challenge
C1714981|T201|COMP|43604-8|LNC|Aldosterone^1st specimen post XXX challenge|Aldosterone^1st specimen post XXX challenge
C1714982|T201|COMP|43605-5|LNC|Albumin|Albumin
C1714983|T201|COMP|43606-3|LNC|Albumin|Albumin
C1714984|T201|COMP|43608-9|LNC|Adrenal cortex Ab|Adrenal cortex Ab
C1714985|T201|COMP|43609-7|LNC|Adipate|Adipate
C1714986|T201|COMP|43610-5|LNC|Adenovirus Ag|Adenovirus Ag
C1714987|T201|COMP|43611-3|LNC|Adenovirus Ag|Adenovirus Ag
C1714988|T201|COMP|43612-1|LNC|Adenovirus Ag|Adenovirus Ag
C1714989|T201|COMP|43614-7|LNC|Adenovirus Ag|Adenovirus Ag
C1714990|T201|COMP|43615-4|LNC|Adenovirus Ag|Adenovirus Ag
C1714991|T201|COMP|43616-2|LNC|Adenovirus Ab|Adenovirus Ab
C1714992|T201|COMP|43617-0|LNC|Adenovirus Ab|Adenovirus Ab
C1714993|T201|COMP|43618-8|LNC|Adenovirus Ab|Adenovirus Ab
C1714994|T201|COMP|43619-6|LNC|Actinomyces sp Ab|Actinomyces sp Ab
C1714995|T201|COMP|43620-4|LNC|Actinomyces israelii Ab|Actinomyces israelii Ab
C1714996|T201|COMP|43621-2|LNC|Actinomyces bovis Ab|Actinomyces bovis Ab
C1714997|T201|COMP|43622-0|LNC|Aconitate|Aconitate
C1714998|T201|COMP|43623-8|LNC|Acetylcholine receptor blocking Ab|Acetylcholine receptor blocking Ab
C1714999|T201|COMP|43624-6|LNC|Acetylcholine receptor binding Ab|Acetylcholine receptor binding Ab
C1715000|T201|COMP|43625-3|LNC|Acetylcholine receptor Ab|Acetylcholine receptor Ab
C1715001|T201|COMP|43626-1|LNC|acetoHEXAMIDE|acetoHEXAMIDE
C1715002|T201|COMP|43627-9|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C1715003|T201|COMP|43628-7|LNC|Acetaminophen crystals|Acetaminophen crystals
C1715004|T201|COMP|43630-3|LNC|6-Thioguanine|6-Thioguanine
C1715005|T201|COMP|43631-1|LNC|6-Methylmercaptopurine metabolite|6-Methylmercaptopurine metabolite
C1715006|T201|COMP|43632-9|LNC|6-Methylmercaptopurine|6-Methylmercaptopurine
C1715007|T201|COMP|43633-7|LNC|5-Oxoproline|5-Oxoproline
C1715008|T201|COMP|43634-5|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C1715009|T201|COMP|43635-2|LNC|2-Hydroxyglutarate|2-Hydroxyglutarate
C1715010|T201|COMP|43636-0|LNC|Plasminogen activator tissue type|Plasminogen activator tissue type
C1715011|T201|COMP|43637-8|LNC|Parrot droppings Ab.IgG|Parrot droppings Ab.IgG
C1715012|T201|COMP|43638-6|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C1715013|T201|COMP|43639-4|LNC|Mercaptopurine|Mercaptopurine
C1715014|T201|COMP|43640-2|LNC|Aldosterone-18-glucuronide|Aldosterone-18-glucuronide
C1715038|T201|COMP|43674-1|LNC|Fatty acid panel.comprehensive C8-C26|Fatty acid panel.comprehensive C8-C26
C1715039|T201|COMP|43675-8|LNC|Fatty acid panel.mitochondrial C8-C18|Fatty acid panel.mitochondrial C8-C18
C1715040|T201|COMP|43676-6|LNC|Fatty acid panel.essential C12-C22|Fatty acid panel.essential C12-C22
C1715041|T201|COMP|43677-4|LNC|Fatty acid panel.very long chain C22-C26|Fatty acid panel.very long chain C22-C26
C1715042|T201|COMP|43691-5|LNC|Cladosporium sp Ab.IgE|Cladosporium sp Ab.IgE
C1715043|T201|COMP|43692-3|LNC|Fusarium sp Ab.IgE.RAST class|Fusarium sp Ab.IgE.RAST class
C1715044|T201|COMP|43693-1|LNC|Varicella zoster virus identified|Varicella zoster virus identified
C1715045|T201|COMP|43694-9|LNC|Inner Ear 68kD Ab|Inner Ear 68kD Ab
C1715046|T201|COMP|43695-6|LNC|Herpes virus identified|Herpes virus identified
C1715047|T201|COMP|43697-2|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1715048|T201|COMP|43698-0|LNC|Enterovirus identified|Enterovirus identified
C1715049|T201|COMP|43699-8|LNC|Enterovirus identified|Enterovirus identified
C1715050|T201|COMP|43700-4|LNC|Cytomegalovirus|Cytomegalovirus
C1715051|T201|COMP|43701-2|LNC|Cytomegalovirus|Cytomegalovirus
C1715052|T201|COMP|43702-0|LNC|Cytomegalovirus|Cytomegalovirus
C1715053|T201|COMP|43703-8|LNC|Cytomegalovirus|Cytomegalovirus
C1715054|T201|COMP|43704-6|LNC|Cytomegalovirus|Cytomegalovirus
C1715055|T201|COMP|43705-3|LNC|Cytomegalovirus|Cytomegalovirus
C1715056|T201|COMP|43706-1|LNC|Cytomegalovirus|Cytomegalovirus
C1715057|T201|COMP|43707-9|LNC|Cytomegalovirus|Cytomegalovirus
C1715058|T201|COMP|43708-7|LNC|Alkaline phosphatase.liver+bone|Alkaline phosphatase.liver+bone
C1715059|T201|COMP|43709-5|LNC|Alkaline phosphatase.intestinal+renal|Alkaline phosphatase.intestinal+renal
C1715060|T201|COMP|43710-3|LNC|Alkaline phosphatase.heat stable|Alkaline phosphatase.heat stable
C1715061|T201|COMP|43711-1|LNC|Albumin|Albumin
C1715062|T201|COMP|43712-9|LNC|Albumin|Albumin
C1715063|T201|COMP|43714-5|LNC|Adenovirus Ab|Adenovirus Ab
C1715064|T201|COMP|43715-2|LNC|Acylcarnitine|Acylcarnitine
C1715065|T201|COMP|43716-0|LNC|Acylcarnitine|Acylcarnitine
C1715066|T201|COMP|43717-8|LNC|Acylcarnitine|Acylcarnitine
C1715067|T201|COMP|43718-6|LNC|Acid phosphatase.prostatic|Acid phosphatase.prostatic
C1715068|T201|COMP|43720-2|LNC|Acetaminophen+Codeine|Acetaminophen+Codeine
C1715069|T201|COMP|43721-0|LNC|Acetaldehyde+Paraldehyde|Acetaldehyde+Paraldehyde
C1715070|T201|COMP|43722-8|LNC|5-Ethyl-5-Phenylhydantoin|5-Ethyl-5-Phenylhydantoin
C1715071|T201|COMP|43723-6|LNC|5,10-Methylenetetrahydrofolate reductase|5,10-Methylenetetrahydrofolate reductase
C1715072|T201|COMP|43724-4|LNC|2,5-Dichlorophenol|2,5-Dichlorophenol
C1715073|T201|COMP|43725-1|LNC|2,4-Dichlorophenol|2,4-Dichlorophenol
C1715074|T201|COMP|43726-9|LNC|17-Ketogenic steroids|17-Ketogenic steroids
C1715075|T201|COMP|43727-7|LNC|Lipoprotein.beta.subparticle.small|Lipoprotein.beta.subparticle.small
C1715076|T201|COMP|43728-5|LNC|Lipoprotein.pre-beta.subparticle.large|Lipoprotein.pre-beta.subparticle.large
C1715077|T201|COMP|43729-3|LNC|Lipoprotein.alpha.subparticle.large|Lipoprotein.alpha.subparticle.large
C1715078|T201|COMP|43730-1|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1715079|T201|COMP|43731-9|LNC|Alkaline phosphatase.fetal+lung+lymphocyte|Alkaline phosphatase.fetal+lung+lymphocyte
C1715080|T201|COMP|43732-7|LNC|4-Hydroxybenzoate|4-Hydroxybenzoate
C1715081|T201|COMP|43733-5|LNC|4-Hydroxybenzoate|4-Hydroxybenzoate
C1715082|T201|COMP|43734-3|LNC|Coagulation surface induced|Coagulation surface induced
C1715083|T201|COMP|43745-9|LNC|DYS gene mutations tested for|DYS gene mutations tested for
C1715084|T201|COMP|43746-7|LNC|KCNQ1 gene targeted mutation analysis|KCNQ1 gene targeted mutation analysis
C1715085|T201|COMP|43747-5|LNC|OCA2 gene targeted mutation analysis|OCA2 gene targeted mutation analysis
C1715086|T201|COMP|43748-3|LNC|SCO1 gene targeted mutation analysis|SCO1 gene targeted mutation analysis
C1715087|T201|COMP|43749-1|LNC|SCO2 gene targeted mutation analysis|SCO2 gene targeted mutation analysis
C1715088|T201|COMP|43751-7|LNC|Moxifloxacin|Moxifloxacin
C1715124|T201|COMP|43800-2|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C1715125|T201|COMP|43801-0|LNC|Choriogonadotropin.intact|Choriogonadotropin.intact
C1715126|T201|COMP|43802-8|LNC|Estriol|Estriol
C1715127|T201|COMP|43803-6|LNC|Estriol^^adjusted|Estriol^^adjusted
C1715128|T201|COMP|43804-4|LNC|Amino acid pattern|Amino acid pattern
C1715129|T201|COMP|43805-1|LNC|Urease^1H post incubation|Urease^1H post incubation
C1715130|T201|COMP|43806-9|LNC|Urease^20M post incubation|Urease^20M post incubation
C1715131|T201|COMP|43807-7|LNC|Urease^4H post incubation|Urease^4H post incubation
C1715132|T201|COMP|43808-5|LNC|Urease^30M post incubation|Urease^30M post incubation
C1715133|T201|COMP|43809-3|LNC|Arsenic|Arsenic
C1715134|T201|COMP|43810-1|LNC|Rubella virus Ab|Rubella virus Ab
C1715135|T201|COMP|43811-9|LNC|Propoxyphene|Propoxyphene
C1715136|T201|COMP|43813-5|LNC|Reagin Ab|Reagin Ab
C1715137|T201|COMP|43814-3|LNC|Basement membrane Ab.IgG|Basement membrane Ab.IgG
C1715138|T201|COMP|43817-6|LNC|Androstenedione|Androstenedione
C1715139|T201|COMP|43818-4|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C1715140|T201|COMP|43819-2|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C1715141|T201|COMP|43820-0|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C1715142|T201|COMP|43821-8|LNC|Amylase|Amylase
C1715143|T201|COMP|43831-7|LNC|Phenytoin|Phenytoin
C1715144|T201|COMP|43832-5|LNC|quiNIDine|quiNIDine
C1715145|T201|COMP|43833-3|LNC|quiNINE|quiNINE
C1715146|T201|COMP|43834-1|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C1715147|T201|COMP|43835-8|LNC|Apolipoprotein E|Apolipoprotein E
C1715148|T201|COMP|43836-6|LNC|Beta globulin|Beta globulin
C1715149|T201|COMP|43838-2|LNC|Influenza virus A Ab.IgM|Influenza virus A Ab.IgM
C1715150|T201|COMP|43840-8|LNC|Influenza virus B Ab.IgM|Influenza virus B Ab.IgM
C1715151|T201|COMP|43841-6|LNC|Betula populifolia Ab.IgE.RAST class|Betula populifolia Ab.IgE.RAST class
C1715152|T201|COMP|43842-4|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C1715153|T201|COMP|43843-2|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C1715154|T201|COMP|43844-0|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C1715155|T201|COMP|43845-7|LNC|Chlamydophila pneumoniae Ab|Chlamydophila pneumoniae Ab
C1715156|T201|COMP|43846-5|LNC|Chlamydophila sp Ab|Chlamydophila sp Ab
C1715157|T201|COMP|43847-3|LNC|Chlamydophila sp Ab|Chlamydophila sp Ab
C1715158|T201|COMP|43848-1|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C1715159|T201|COMP|43849-9|LNC|Coccidioides sp Ab.IgG|Coccidioides sp Ab.IgG
C1715160|T201|COMP|43850-7|LNC|Coccidioides sp Ab.IgM|Coccidioides sp Ab.IgM
C1715161|T201|COMP|43851-5|LNC|Influenza virus A Ab.IgA|Influenza virus A Ab.IgA
C1715162|T201|COMP|43852-3|LNC|Influenza virus B Ab.IgA|Influenza virus B Ab.IgA
C1715163|T201|COMP|43853-1|LNC|Legionella pneumophila 1+3+4+5+6+8 Ab.IgM|Legionella pneumophila 1+3+4+5+6+8 Ab.IgM
C1715164|T201|COMP|43854-9|LNC|Mycobacterium sp rRNA|Mycobacterium sp rRNA
C1715165|T201|COMP|43857-2|LNC|Benztropine|Benztropine
C1715166|T201|COMP|43858-0|LNC|Beta-2 transferrin|Beta-2 transferrin
C1715167|T201|COMP|43859-8|LNC|Bolasterone|Bolasterone
C1715168|T201|COMP|43860-6|LNC|Amphetamine+Methamphetamine|Amphetamine+Methamphetamine
C1715169|T201|COMP|43861-4|LNC|Asialoganglioside GM1 Ab|Asialoganglioside GM1 Ab
C1715170|T201|COMP|43862-2|LNC|Aspergillus sp Ab.IgE.RAST class|Aspergillus sp Ab.IgE.RAST class
C1715171|T201|COMP|43863-0|LNC|Benzthiazide|Benzthiazide
C1715172|T201|COMP|43864-8|LNC|Blastomyces dermatitidis Ab.IgG|Blastomyces dermatitidis Ab.IgG
C1715173|T201|COMP|43865-5|LNC|Blastomyces dermatitidis Ab.IgG|Blastomyces dermatitidis Ab.IgG
C1715174|T201|COMP|43866-3|LNC|Bartonella sp Ab|Bartonella sp Ab
C1715175|T201|COMP|43867-1|LNC|Beta-2 transferrin|Beta-2 transferrin
C1715176|T201|COMP|43868-9|LNC|Chlamydophila psittaci Ab.IgG|Chlamydophila psittaci Ab.IgG
C1715177|T201|COMP|43869-7|LNC|Antithrombin Ag|Antithrombin Ag
C1715178|T201|COMP|43870-5|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C1715179|T201|COMP|43871-3|LNC|Aspergillus sp Ab.IgA|Aspergillus sp Ab.IgA
C1715180|T201|COMP|43872-1|LNC|Aspergillus sp Ab.IgG|Aspergillus sp Ab.IgG
C1715181|T201|COMP|43875-4|LNC|Basement membrane Ab.IgM|Basement membrane Ab.IgM
C1715182|T201|COMP|43877-0|LNC|Bile acid|Bile acid
C1715183|T201|COMP|43878-8|LNC|Bismuth|Bismuth
C1715184|T201|COMP|43879-6|LNC|Bordetella parapertussis|Bordetella parapertussis
C1715188|T201|COMP|43883-8|LNC|Ampicillin|Ampicillin
C1715189|T201|COMP|43884-6|LNC|Ampicillin|Ampicillin
C1715190|T201|COMP|43885-3|LNC|Beryllium|Beryllium
C1715191|T201|COMP|43886-1|LNC|Bismuth|Bismuth
C1715192|T201|COMP|43887-9|LNC|Bilirubin|Bilirubin
C1715193|T201|COMP|43888-7|LNC|Bile acid|Bile acid
C1715194|T201|COMP|43889-5|LNC|Bile acid|Bile acid
C1715195|T201|COMP|43890-3|LNC|Bordetella pertussis|Bordetella pertussis
C1715196|T201|COMP|43891-1|LNC|Bordetella pertussis Ag|Bordetella pertussis Ag
C1715197|T201|COMP|43893-7|LNC|Babesia microti Ab.IgG|Babesia microti Ab.IgG
C1715198|T201|COMP|43895-2|LNC|Influenza virus B Ag|Influenza virus B Ag
C1715199|T201|COMP|43896-0|LNC|Bordetella pertussis|Bordetella pertussis
C1715200|T201|COMP|43897-8|LNC|Baclofen|Baclofen
C1715201|T201|COMP|43898-6|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C1715202|T201|COMP|43899-4|LNC|Beta lipotropin|Beta lipotropin
C1715203|T201|COMP|43900-0|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C1715204|T201|COMP|43901-8|LNC|Barium|Barium
C1715205|T201|COMP|43902-6|LNC|Azinphos-methyl|Azinphos-methyl
C1715206|T201|COMP|43904-2|LNC|Azinphos-methyl|Azinphos-methyl
C1715207|T201|COMP|43905-9|LNC|Arbovirus Ab.IgG|Arbovirus Ab.IgG
C1715208|T201|COMP|43906-7|LNC|Anserine|Anserine
C1715209|T201|COMP|43907-5|LNC|Argininosuccinate|Argininosuccinate
C1715210|T201|COMP|43908-3|LNC|Avian encephalomyelitis virus Ab|Avian encephalomyelitis virus Ab
C1715211|T201|COMP|43910-9|LNC|Ascaris sp Ab.IgM|Ascaris sp Ab.IgM
C1715212|T201|COMP|43911-7|LNC|Aspergillus versicolor Ab|Aspergillus versicolor Ab
C1715213|T201|COMP|43912-5|LNC|Bisacodyl|Bisacodyl
C1715214|T201|COMP|43913-3|LNC|Bordetella pertussis DNA|Bordetella pertussis DNA
C1715215|T201|COMP|43914-1|LNC|Beta 2 glycoprotein 1 Ab.IgG|Beta 2 glycoprotein 1 Ab.IgG
C1715216|T201|COMP|43915-8|LNC|Beta 2 glycoprotein 1 Ab.IgA|Beta 2 glycoprotein 1 Ab.IgA
C1715217|T201|COMP|43916-6|LNC|Beta 2 glycoprotein 1 Ab.IgM|Beta 2 glycoprotein 1 Ab.IgM
C1715218|T201|COMP|43917-4|LNC|Benzene|Benzene
C1715219|T201|COMP|43918-2|LNC|Babesia microti Ab|Babesia microti Ab
C1715220|T201|COMP|43919-0|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C1715221|T201|COMP|43920-8|LNC|Bartonella sp Ab.IgG|Bartonella sp Ab.IgG
C1715222|T201|COMP|43930-7|LNC|Yersinia enterocolitica Ab|Yersinia enterocolitica Ab
C1715223|T201|COMP|43931-5|LNC|California encephalitis virus Ab|California encephalitis virus Ab
C1715224|T201|COMP|43933-1|LNC|Cathine|Cathine
C1715225|T201|COMP|43934-9|LNC|Amphetamines|Amphetamines
C1715226|T201|COMP|43935-6|LNC|Cells.CD55/100 cells|Cells.CD55/100 cells
C1715227|T201|COMP|43936-4|LNC|Cells.CD55/100 cells|Cells.CD55/100 cells
C1715228|T201|COMP|43937-2|LNC|Cells.CD59/100 cells|Cells.CD59/100 cells
C1715229|T201|COMP|43939-8|LNC|Alkaline phosphatase.liver|Alkaline phosphatase.liver
C1715230|T201|COMP|43940-6|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C1715231|T201|COMP|43941-4|LNC|Agrostis stolonifera Ab.IgE/IgE.total|Agrostis stolonifera Ab.IgE/IgE.total
C1715232|T201|COMP|43942-2|LNC|Insulin.free|Insulin.free
C1715233|T201|COMP|43943-0|LNC|Cat epithelium Ab.IgE|Cat epithelium Ab.IgE
C1715234|T201|COMP|43944-8|LNC|Cells.CD4+CD45+/100 cells|Cells.CD4+CD45+/100 cells
C1715235|T201|COMP|43945-5|LNC|Cells.CD4+CD45RO+/100 cells|Cells.CD4+CD45RO+/100 cells
C1715236|T201|COMP|43946-3|LNC|Cells.CD4+CD45RO+/100 cells|Cells.CD4+CD45RO+/100 cells
C1715237|T201|COMP|43947-1|LNC|Cells.CD4+CD45+/100 cells|Cells.CD4+CD45+/100 cells
C1715238|T201|COMP|43948-9|LNC|Cells.CD4+CD45RO+/100 cells|Cells.CD4+CD45RO+/100 cells
C1715239|T201|COMP|43949-7|LNC|Cells.CD2|Cells.CD2
C1715240|T201|COMP|43950-5|LNC|Cells.CD2|Cells.CD2
C1715241|T201|COMP|43951-3|LNC|Cells.CD2|Cells.CD2
C1715242|T201|COMP|43952-1|LNC|Cells.CD4+CD45RO+|Cells.CD4+CD45RO+
C1715243|T201|COMP|43953-9|LNC|Cells.CD4+CD45RO+|Cells.CD4+CD45RO+
C1715244|T201|COMP|43956-2|LNC|Cells.CD4+CD45RO+|Cells.CD4+CD45RO+
C1715245|T201|COMP|43957-0|LNC|Cells.CD3+HLA-DR+|Cells.CD3+HLA-DR+
C1715246|T201|COMP|43958-8|LNC|Cells.CD3+HLA-DR+|Cells.CD3+HLA-DR+
C1715247|T201|COMP|43959-6|LNC|Cells.CD3+HLA-DR+|Cells.CD3+HLA-DR+
C1715248|T201|COMP|43960-4|LNC|Cells.CD3+HLA-DR+|Cells.CD3+HLA-DR+
C1715249|T201|COMP|43961-2|LNC|Cells.CD3+HLA-DR+|Cells.CD3+HLA-DR+
C1715250|T201|COMP|43962-0|LNC|Cells.CD4+CD45RA+/100 cells|Cells.CD4+CD45RA+/100 cells
C1715251|T201|COMP|43963-8|LNC|Cells.CD4+CD45RA+/100 cells|Cells.CD4+CD45RA+/100 cells
C1715252|T201|COMP|43964-6|LNC|Cells.CD4+CD45RA+/100 cells|Cells.CD4+CD45RA+/100 cells
C1715253|T201|COMP|43965-3|LNC|Cells.CD4+CD45RA+/100 cells|Cells.CD4+CD45RA+/100 cells
C1715254|T201|COMP|43967-9|LNC|Cells.CD3+CD25+/100 cells|Cells.CD3+CD25+/100 cells
C1715255|T201|COMP|43968-7|LNC|Cells.CD3+HLA-DR+/100 cells|Cells.CD3+HLA-DR+/100 cells
C1715256|T201|COMP|43969-5|LNC|Cells.CD3+CD25+|Cells.CD3+CD25+
C1715257|T201|COMP|43970-3|LNC|Cells.CD3+CD4+/100 cells|Cells.CD3+CD4+/100 cells
C1715258|T201|COMP|43971-1|LNC|Cells.CD3+CD8+/100 cells|Cells.CD3+CD8+/100 cells
C1715259|T201|COMP|43973-7|LNC|Zinc|Zinc
C1715260|T201|COMP|43974-5|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1715261|T201|COMP|43975-2|LNC|Aprobarbital|Aprobarbital
C1715262|T201|COMP|43976-0|LNC|Measles virus Ab|Measles virus Ab
C1715263|T201|COMP|43977-8|LNC|Anabolic steroids|Anabolic steroids
C1715264|T201|COMP|43978-6|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C1715265|T201|COMP|43979-4|LNC|Aspergillus sp identified|Aspergillus sp identified
C1715266|T201|COMP|43980-2|LNC|Rabies virus Ab|Rabies virus Ab
C1715267|T201|COMP|43981-0|LNC|Choriogonadotropin.intact^^adjusted|Choriogonadotropin.intact^^adjusted
C1715268|T201|COMP|43982-8|LNC|Choriogonadotropin.intact|Choriogonadotropin.intact
C1715269|T201|COMP|43983-6|LNC|Amphetamines|Amphetamines
C1715270|T201|COMP|43984-4|LNC|Benzoylecgonine|Benzoylecgonine
C1715271|T201|COMP|43985-1|LNC|Benzoylecgonine|Benzoylecgonine
C1715272|T201|COMP|43986-9|LNC|Clofazimine 2.0 ug/mL|Clofazimine 2.0 ug/mL
C1715273|T201|COMP|43987-7|LNC|Clarithromycin 12.0 ug/mL|Clarithromycin 12.0 ug/mL
C1715274|T201|COMP|43988-5|LNC|Clofazimine 0.5 ug/mL|Clofazimine 0.5 ug/mL
C1715275|T201|COMP|43989-3|LNC|Clofazimine 1.0 ug/mL|Clofazimine 1.0 ug/mL
C1715276|T201|COMP|43991-9|LNC|Clarithromycin 6.0 ug/mL|Clarithromycin 6.0 ug/mL
C1715277|T201|COMP|43992-7|LNC|Anaplasma phagocytophilum Ab|Anaplasma phagocytophilum Ab
C1715279|T201|COMP|43994-3|LNC|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C1715280|T201|COMP|43995-0|LNC|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C1715281|T201|COMP|43996-8|LNC|Alpha-1-Fetoprotein^^adjusted for diabetes+weight|Alpha-1-Fetoprotein^^adjusted for diabetes+weight
C1715282|T201|COMP|43997-6|LNC|Alpha-1-Fetoprotein^^adjusted for weight|Alpha-1-Fetoprotein^^adjusted for weight
C1715283|T201|COMP|43998-4|LNC|Alpha-1-Fetoprotein^^adjusted for diabetes|Alpha-1-Fetoprotein^^adjusted for diabetes
C1715284|T201|COMP|43999-2|LNC|Choriogonadotropin|Choriogonadotropin
C1715285|T201|COMP|44000-8|LNC|Choriogonadotropin|Choriogonadotropin
C1715286|T201|COMP|44001-6|LNC|Choriogonadotropin|Choriogonadotropin
C1715287|T201|COMP|44002-4|LNC|Choriogonadotropin^^adjusted|Choriogonadotropin^^adjusted
C1715288|T201|COMP|44003-2|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C1715289|T201|COMP|44004-0|LNC|Estriol.unconjugated|Estriol.unconjugated
C1715290|T201|COMP|44005-7|LNC|Chlamydia trachomatis D & K Ab.IgA & IgG & IgM|Chlamydia trachomatis D & K Ab.IgA & IgG & IgM
C1715291|T201|COMP|44006-5|LNC|Coxiella burnetii phase 1 & 2 Ab.IgG & IgM|Coxiella burnetii phase 1 & 2 Ab.IgG & IgM
C1715292|T201|COMP|44008-1|LNC|Herpes simplex virus 1 & 2 Ab.IgM|Herpes simplex virus 1 & 2 Ab.IgM
C1715293|T201|COMP|44009-9|LNC|Herpes simplex virus 1 & 2 Ab.IgG|Herpes simplex virus 1 & 2 Ab.IgG
C1715294|T201|COMP|44010-7|LNC|Influenza virus A & B Ab|Influenza virus A & B Ab
C1715295|T201|COMP|44011-5|LNC|Measles virus Ab.IgG & IgM|Measles virus Ab.IgG & IgM
C1715296|T201|COMP|44012-3|LNC|Measles virus Ab.IgG & IgM|Measles virus Ab.IgG & IgM
C1715297|T201|COMP|44013-1|LNC|Metanephrine & Normetanephrine|Metanephrine & Normetanephrine
C1715298|T201|COMP|44014-9|LNC|Porphyrins|Porphyrins
C1715299|T201|COMP|44015-6|LNC|Helicobacter pylori|Helicobacter pylori
C1715300|T201|COMP|44016-4|LNC|Bile|Bile
C1715301|T201|COMP|44018-0|LNC|Basophils|Basophils
C1715302|T201|COMP|44019-8|LNC|Bordetella parapertussis Ab|Bordetella parapertussis Ab
C1715303|T201|COMP|44020-6|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C1715304|T201|COMP|44021-4|LNC|Coxiella burnetii Ab|Coxiella burnetii Ab
C1715305|T201|COMP|44022-2|LNC|Bacteria|Bacteria
C1715306|T201|COMP|44023-0|LNC|Bacteria|Bacteria
C1715307|T201|COMP|44024-8|LNC|Boldenone|Boldenone
C1715308|T201|COMP|44026-3|LNC|Aspergillus flavus H Ab|Aspergillus flavus H Ab
C1715309|T201|COMP|44028-9|LNC|Aspergillus fumigatus H Ab|Aspergillus fumigatus H Ab
C1715310|T201|COMP|44029-7|LNC|Aspergillus nidulans B Ab|Aspergillus nidulans B Ab
C1715311|T201|COMP|44031-3|LNC|Aspergillus niger B Ab|Aspergillus niger B Ab
C1715312|T201|COMP|44032-1|LNC|Aspergillus niger H Ab|Aspergillus niger H Ab
C1715313|T201|COMP|44033-9|LNC|Bilirubin|Bilirubin
C1715314|T201|COMP|44034-7|LNC|Bile canalicular Ab|Bile canalicular Ab
C1715315|T201|COMP|44035-4|LNC|Analgesics.non-narcotic|Analgesics.non-narcotic
C1715316|T201|COMP|44036-2|LNC|Analgesics.non-narcotic|Analgesics.non-narcotic
C1715317|T201|COMP|44037-0|LNC|Glucosylceramidase|Glucosylceramidase
C1715318|T201|COMP|44038-8|LNC|Bacteria|Bacteria
C1715319|T201|COMP|44039-6|LNC|Bacteria|Bacteria
C1715320|T201|COMP|44040-4|LNC|Basophils|Basophils
C1715321|T201|COMP|44042-0|LNC|Basophils|Basophils
C1715322|T201|COMP|44043-8|LNC|Basophils|Basophils
C1715323|T201|COMP|44044-6|LNC|Basophils|Basophils
C1715324|T201|COMP|44045-3|LNC|Aspergillus fumigatus O Ab|Aspergillus fumigatus O Ab
C1715325|T201|COMP|44046-1|LNC|Bordetella pertussis Higashi-Hama Ab|Bordetella pertussis Higashi-Hama Ab
C1715326|T201|COMP|44047-9|LNC|Bordetella pertussis Yamaguchi Ab|Bordetella pertussis Yamaguchi Ab
C1715327|T201|COMP|44048-7|LNC|Basophils|Basophils
C1715328|T201|COMP|44049-5|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C1715329|T201|COMP|44051-1|LNC|Adenylate kinase|Adenylate kinase
C1715330|T201|COMP|44052-9|LNC|Phosphofructokinase|Phosphofructokinase
C1715331|T201|COMP|44053-7|LNC|Phosphoglycerate kinase|Phosphoglycerate kinase
C1715332|T201|COMP|44054-5|LNC|Triosephosphate isomerase|Triosephosphate isomerase
C1715333|T201|COMP|44055-2|LNC|Pyrimidine-5'-Nucleotidase|Pyrimidine-5'-Nucleotidase
C1715334|T201|COMP|44056-0|LNC|Cells.CD4+CD45RA+CD45RB+CD45RC+|Cells.CD4+CD45RA+CD45RB+CD45RC+
C1715335|T201|COMP|44057-8|LNC|Cells.CD4+CD45RA+CD45RB+CD45RC+|Cells.CD4+CD45RA+CD45RB+CD45RC+
C1715336|T201|COMP|44058-6|LNC|Cells.CD4+CD45RA+CD45RB+CD45RC+|Cells.CD4+CD45RA+CD45RB+CD45RC+
C1715337|T201|COMP|44059-4|LNC|Cells.CD4+CD45RA+CD45RB+CD45RC+|Cells.CD4+CD45RA+CD45RB+CD45RC+
C1715338|T201|COMP|44060-2|LNC|Cells.CD4+CD45RA+CD45RB+CD45RC+|Cells.CD4+CD45RA+CD45RB+CD45RC+
C1715339|T201|COMP|44061-0|LNC|Cells.CD20+FMC7+/100 cells|Cells.CD20+FMC7+/100 cells
C1715340|T201|COMP|44062-8|LNC|Cells.CD20+FMC7+/100 cells|Cells.CD20+FMC7+/100 cells
C1715341|T201|COMP|44063-6|LNC|Cells.CD20+FMC7+/100 cells|Cells.CD20+FMC7+/100 cells
C1715342|T201|COMP|44064-4|LNC|Cells.CD20+FMC7+/100 cells|Cells.CD20+FMC7+/100 cells
C1715343|T201|COMP|44065-1|LNC|Cells.CD20+FMC7+|Cells.CD20+FMC7+
C1715344|T201|COMP|44066-9|LNC|Cells.CD20+FMC7+|Cells.CD20+FMC7+
C1715345|T201|COMP|44068-5|LNC|Cells.CD20+FMC7+|Cells.CD20+FMC7+
C1715346|T201|COMP|44069-3|LNC|Cells.CD20+FMC7+|Cells.CD20+FMC7+
C1715347|T201|COMP|44070-1|LNC|Cells.CD20+CD52+/100 cells|Cells.CD20+CD52+/100 cells
C1715348|T201|COMP|44071-9|LNC|Cells.CD20+CD52+/100 cells|Cells.CD20+CD52+/100 cells
C1715349|T201|COMP|44072-7|LNC|Cells.CD20+CD52+/100 cells|Cells.CD20+CD52+/100 cells
C1715350|T201|COMP|44073-5|LNC|Cells.CD20+CD52+/100 cells|Cells.CD20+CD52+/100 cells
C1715351|T201|COMP|44075-0|LNC|Bilirubin casts|Bilirubin casts
C1715352|T201|COMP|44076-8|LNC|Alpha tocopherol & Beta+gamma tocopherol|Alpha tocopherol & Beta+gamma tocopherol
C1715353|T201|COMP|44077-6|LNC|Brucella canis Ab.IgG & IgM|Brucella canis Ab.IgG & IgM
C1715354|T201|COMP|44078-4|LNC|Catecholamines|Catecholamines
C1715355|T201|COMP|44080-0|LNC|Chlamydophila pneumoniae Ab.IgG & IgM|Chlamydophila pneumoniae Ab.IgG & IgM
C1715356|T201|COMP|44081-8|LNC|Chlamydophila psittaci Ab.IgA & IgG & IgM|Chlamydophila psittaci Ab.IgA & IgG & IgM
C1715357|T201|COMP|44082-6|LNC|Cryoglobulin IgA & IgG & IgM|Cryoglobulin IgA & IgG & IgM
C1715358|T201|COMP|44083-4|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C1715359|T201|COMP|44084-2|LNC|Fatty acids pattern|Fatty acids pattern
C1715360|T201|COMP|44085-9|LNC|Xylose absorption|Xylose absorption
C1715361|T201|COMP|44086-7|LNC|ABO & Rh group|ABO & Rh group
C1715362|T201|COMP|44087-5|LNC|Escherichia coli O157 Ag|Escherichia coli O157 Ag
C1715363|T201|COMP|44088-3|LNC|Escherichia coli O157:H7 DNA|Escherichia coli O157:H7 DNA
C1715364|T201|COMP|44089-1|LNC|Escherichia coli O157:H7|Escherichia coli O157:H7
C1715365|T201|COMP|44090-9|LNC|Escherichia coli O157:H7|Escherichia coli O157:H7
C1715366|T201|COMP|44092-5|LNC|Leukocytes|Leukocytes
C1715367|T201|COMP|44093-3|LNC|Neisseria meningitidis|Neisseria meningitidis
C1715368|T201|COMP|44094-1|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C1715369|T201|COMP|44095-8|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C1715370|T201|COMP|44096-6|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C1715371|T201|COMP|44097-4|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C1715499|T201|COMP|44241-8|LNC|Clue cells|Clue cells
C1715500|T201|COMP|44242-6|LNC|Erythrocytes|Erythrocytes
C1715501|T201|COMP|44243-4|LNC|Bacteria|Bacteria
C1715502|T201|COMP|44244-2|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C1715503|T201|COMP|44245-9|LNC|Fungi.filamentous|Fungi.filamentous
C1715504|T201|COMP|44246-7|LNC|Yeast|Yeast
C1715505|T201|COMP|44247-5|LNC|Spermatozoa.motile|Spermatozoa.motile
C1715506|T201|COMP|44248-3|LNC|Spermatozoa.immotile|Spermatozoa.immotile
C1715520|T201|COMP|44263-2|LNC|Influenza virus A RNA|Influenza virus A RNA
C1715521|T201|COMP|44264-0|LNC|Influenza virus A H5 RNA|Influenza virus A H5 RNA
C1715522|T201|COMP|44266-5|LNC|Influenza virus A H7 RNA|Influenza virus A H7 RNA
C1715523|T201|COMP|44267-3|LNC|Avian paramyxovirus 1 RNA|Avian paramyxovirus 1 RNA
C1715524|T201|COMP|44268-1|LNC|Avian paramyxovirus 1.exotic RNA|Avian paramyxovirus 1.exotic RNA
C1715525|T201|COMP|44269-9|LNC|Bacillus anthracis cell wall Ag|Bacillus anthracis cell wall Ag
C1715526|T201|COMP|44270-7|LNC|Bacillus anthracis spore Ag|Bacillus anthracis spore Ag
C1715527|T201|COMP|44271-5|LNC|Brucella sp Ag|Brucella sp Ag
C1715528|T201|COMP|44272-3|LNC|Cache valley virus Ab|Cache valley virus Ab
C1715529|T201|COMP|44273-1|LNC|Classical swine fever virus RNA|Classical swine fever virus RNA
C1715530|T201|COMP|44274-9|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C1715531|T201|COMP|44275-6|LNC|Coxiella burnetii|Coxiella burnetii
C1715532|T201|COMP|44276-4|LNC|Equine adenovirus Ag|Equine adenovirus Ag
C1715534|T201|COMP|44278-0|LNC|16-Alpha hydroxydehydroepiandrosterone/Creatinine|16-Alpha hydroxydehydroepiandrosterone/Creatinine
C1715536|T201|COMP|44280-6|LNC|17 alpha-Hydroxypregnanolone/Creatinine|17 alpha-Hydroxypregnanolone/Creatinine
C1715537|T201|COMP|44281-4|LNC|17-Ketosteroids/Creatinine|17-Ketosteroids/Creatinine
C1715538|T201|COMP|44282-2|LNC|2-Hydroxyisocaproate/Creatinine|2-Hydroxyisocaproate/Creatinine
C1715539|T201|COMP|44283-0|LNC|2-Hydroxyphenylacetate/Creatinine|2-Hydroxyphenylacetate/Creatinine
C1715540|T201|COMP|44284-8|LNC|2-Methylcitrate/Creatinine|2-Methylcitrate/Creatinine
C1715541|T201|COMP|44286-3|LNC|3-Methylhistidine/Creatinine|3-Methylhistidine/Creatinine
C1715542|T201|COMP|44287-1|LNC|5-Hydroxyhexanoate/Creatinine|5-Hydroxyhexanoate/Creatinine
C1715543|T201|COMP|44288-9|LNC|5-Hydroxyindoleacetate/Creatinine|5-Hydroxyindoleacetate/Creatinine
C1715544|T201|COMP|44289-7|LNC|Adenovirus Ab|Adenovirus Ab
C1715545|T201|COMP|44291-3|LNC|Alanine/Creatinine|Alanine/Creatinine
C1715546|T201|COMP|44292-1|LNC|Albumin/Creatinine|Albumin/Creatinine
C1715547|T201|COMP|44293-9|LNC|Albumin/Globulin|Albumin/Globulin
C1715548|T201|COMP|44294-7|LNC|Albumin/Globulin|Albumin/Globulin
C1715549|T201|COMP|44295-4|LNC|Aldosterone/Creatinine|Aldosterone/Creatinine
C1715550|T201|COMP|44296-2|LNC|Alpha aminobutyrate/Creatinine|Alpha aminobutyrate/Creatinine
C1715551|T201|COMP|44297-0|LNC|Androsterone/Creatinine|Androsterone/Creatinine
C1715552|T201|COMP|44298-8|LNC|Apis mellifera Ab.IgG.RAST class|Apis mellifera Ab.IgG.RAST class
C1715553|T201|COMP|44299-6|LNC|Arginine/Creatinine|Arginine/Creatinine
C1715554|T201|COMP|44300-2|LNC|Arsenic.inorganic/Creatinine|Arsenic.inorganic/Creatinine
C1715555|T201|COMP|44301-0|LNC|Asparagine/Creatinine|Asparagine/Creatinine
C1715556|T201|COMP|44302-8|LNC|Aspartate/Creatinine|Aspartate/Creatinine
C1715557|T201|COMP|44303-6|LNC|Beta-2-Microglobulin/Creatinine|Beta-2-Microglobulin/Creatinine
C1715558|T201|COMP|44304-4|LNC|Carnosine/Creatinine|Carnosine/Creatinine
C1715559|T201|COMP|44306-9|LNC|Citrate/Creatinine|Citrate/Creatinine
C1715560|T201|COMP|44308-5|LNC|Collagen crosslinked N-telopeptide/Creatinine|Collagen crosslinked N-telopeptide/Creatinine
C1715561|T201|COMP|44309-3|LNC|Cortisol.free/Creatinine|Cortisol.free/Creatinine
C1715562|T201|COMP|44310-1|LNC|Cortisol/Creatinine|Cortisol/Creatinine
C1715563|T201|COMP|44311-9|LNC|Cotinine/Creatinine|Cotinine/Creatinine
C1715564|T201|COMP|44312-7|LNC|Cystine/Creatinine|Cystine/Creatinine
C1715565|T201|COMP|44313-5|LNC|Delta aminolevulinate/Creatinine|Delta aminolevulinate/Creatinine
C1715566|T201|COMP|44314-3|LNC|D-lactate/Creatinine|D-lactate/Creatinine
C1715567|T201|COMP|44315-0|LNC|Dolichovespula maculata Ab.IgG.RAST class|Dolichovespula maculata Ab.IgG.RAST class
C1715568|T201|COMP|44316-8|LNC|DOPamine/Creatinine|DOPamine/Creatinine
C1715569|T201|COMP|44330-9|LNC|Isospora belli|Isospora belli
C1715570|T201|COMP|44331-7|LNC|Isovalerylglycine/Creatinine|Isovalerylglycine/Creatinine
C1715571|T201|COMP|44332-5|LNC|Jo-1 extractable nuclear Ab.IgG|Jo-1 extractable nuclear Ab.IgG
C1715572|T201|COMP|44333-3|LNC|Lactate/Creatinine|Lactate/Creatinine
C1715573|T201|COMP|44334-1|LNC|Leucine/Creatinine|Leucine/Creatinine
C1715574|T201|COMP|44335-8|LNC|Lysine/Creatinine|Lysine/Creatinine
C1715575|T201|COMP|44336-6|LNC|Magnesium/Creatinine|Magnesium/Creatinine
C1715576|T201|COMP|44338-2|LNC|Methionine/Creatinine|Methionine/Creatinine
C1715577|T201|COMP|44340-8|LNC|N-methylhistamine/Creatinine|N-methylhistamine/Creatinine
C1715578|T201|COMP|44341-6|LNC|Norepinephrine/Creatinine|Norepinephrine/Creatinine
C1715579|T201|COMP|44342-4|LNC|Normetanephrine/Creatinine|Normetanephrine/Creatinine
C1715580|T201|COMP|44343-2|LNC|Organic acids/Creatinine|Organic acids/Creatinine
C1715581|T201|COMP|44344-0|LNC|Ornithine/Creatinine|Ornithine/Creatinine
C1715582|T201|COMP|44345-7|LNC|Orotate/Creatinine|Orotate/Creatinine
C1715583|T201|COMP|44346-5|LNC|Phenol/Creatinine|Phenol/Creatinine
C1715584|T201|COMP|44347-3|LNC|Phenol/Creatinine|Phenol/Creatinine
C1715585|T201|COMP|44348-1|LNC|Phenylalanine/Creatinine|Phenylalanine/Creatinine
C1715586|T201|COMP|44349-9|LNC|Phenylalanine/Creatinine|Phenylalanine/Creatinine
C1715587|T201|COMP|44350-7|LNC|Phenylpropionylglycine/Creatinine|Phenylpropionylglycine/Creatinine
C1715588|T201|COMP|44351-5|LNC|Phosphoethanolamine/Creatinine|Phosphoethanolamine/Creatinine
C1715589|T201|COMP|44352-3|LNC|Phosphoethanolamine/Creatinine|Phosphoethanolamine/Creatinine
C1715590|T201|COMP|44354-9|LNC|Ethylmalonate/Creatinine|Ethylmalonate/Creatinine
C1715591|T201|COMP|44355-6|LNC|Etiocholanolone/Creatinine|Etiocholanolone/Creatinine
C1715592|T201|COMP|44357-2|LNC|Galactomannan Ag|Galactomannan Ag
C1715593|T201|COMP|44358-0|LNC|Gamma hydroxybutyrate/Creatinine|Gamma hydroxybutyrate/Creatinine
C1715594|T201|COMP|44359-8|LNC|Glutamate/Creatinine|Glutamate/Creatinine
C1715595|T201|COMP|44360-6|LNC|Glutamate+Glutamine/Creatinine|Glutamate+Glutamine/Creatinine
C1715596|T201|COMP|44361-4|LNC|Glutamate+Glutamine/Creatinine|Glutamate+Glutamine/Creatinine
C1715597|T201|COMP|44362-2|LNC|Glutamine/Creatinine|Glutamine/Creatinine
C1715598|T201|COMP|44363-0|LNC|Glutarate/Creatinine|Glutarate/Creatinine
C1715599|T201|COMP|44365-5|LNC|Glycine/Creatinine|Glycine/Creatinine
C1715600|T201|COMP|44366-3|LNC|Glycosaminoglycans/Creatinine|Glycosaminoglycans/Creatinine
C1715601|T201|COMP|44367-1|LNC|Glycosaminoglycans/Creatinine|Glycosaminoglycans/Creatinine
C1715602|T201|COMP|44368-9|LNC|Hexanoylglycine/Creatinine|Hexanoylglycine/Creatinine
C1715603|T201|COMP|44369-7|LNC|Hexokinase|Hexokinase
C1715604|T201|COMP|44370-5|LNC|Hippurate/Creatinine|Hippurate/Creatinine
C1715605|T201|COMP|44371-3|LNC|Histamine/Creatinine|Histamine/Creatinine
C1715606|T201|COMP|44372-1|LNC|Histidine/Creatinine|Histidine/Creatinine
C1715607|T201|COMP|44373-9|LNC|Homocysteine|Homocysteine
C1715608|T201|COMP|44374-7|LNC|Homocysteine|Homocysteine
C1715609|T201|COMP|44375-4|LNC|Homocysteine|Homocysteine
C1715610|T201|COMP|44376-2|LNC|Homocysteine|Homocysteine
C1715611|T201|COMP|44378-8|LNC|Homocystine/Creatinine|Homocystine/Creatinine
C1715612|T201|COMP|44379-6|LNC|Horse hair+Horse dander Ab.IgE.RAST class|Horse hair+Horse dander Ab.IgE.RAST class
C1715613|T201|COMP|44380-4|LNC|House dust Hollister Stier Ab.IgG.RAST class|House dust Hollister Stier Ab.IgG.RAST class
C1715614|T201|COMP|44381-2|LNC|Humulus japonicus Ab.IgE.RAST class|Humulus japonicus Ab.IgE.RAST class
C1715615|T201|COMP|44383-8|LNC|Hyaluronate|Hyaluronate
C1715616|T201|COMP|44384-6|LNC|hydroCHLOROthiazide|hydroCHLOROthiazide
C1715617|T201|COMP|44385-3|LNC|Hydroflumethiazide|Hydroflumethiazide
C1715618|T201|COMP|44386-1|LNC|Hydroxyproline/Creatinine|Hydroxyproline/Creatinine
C1715619|T201|COMP|44387-9|LNC|Hypnotics|Hypnotics
C1715620|T201|COMP|44388-7|LNC|IgA|IgA
C1715621|T201|COMP|44389-5|LNC|IgA|IgA
C1715622|T201|COMP|44390-3|LNC|Imipramine|Imipramine
C1715623|T201|COMP|44391-1|LNC|Immune complex|Immune complex
C1715624|T201|COMP|44393-7|LNC|Immune complex|Immune complex
C1715625|T201|COMP|44394-5|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C1715626|T201|COMP|44395-2|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C1715627|T201|COMP|44396-0|LNC|Insulin|Insulin
C1715628|T201|COMP|44397-8|LNC|Insulin bovine Ab|Insulin bovine Ab
C1715629|T201|COMP|44398-6|LNC|Proline/Creatinine|Proline/Creatinine
C1715630|T201|COMP|44399-4|LNC|Propionylglycine/Creatinine|Propionylglycine/Creatinine
C1715631|T201|COMP|44400-0|LNC|Pyruvate/Creatinine|Pyruvate/Creatinine
C1715632|T201|COMP|44402-6|LNC|Selenium/Creatinine|Selenium/Creatinine
C1715633|T201|COMP|44403-4|LNC|Serine/Creatinine|Serine/Creatinine
C1715634|T201|COMP|44404-2|LNC|Silicon/Creatinine|Silicon/Creatinine
C1715635|T201|COMP|44405-9|LNC|Sodium/Creatinine|Sodium/Creatinine
C1715636|T201|COMP|44406-7|LNC|Sodium/Potassium|Sodium/Potassium
C1715637|T201|COMP|44407-5|LNC|Somatotropin/Creatinine|Somatotropin/Creatinine
C1715638|T201|COMP|44409-1|LNC|Succinate/Creatinine|Succinate/Creatinine
C1715639|T201|COMP|44410-9|LNC|Superoxide dismutase|Superoxide dismutase
C1715640|T201|COMP|44411-7|LNC|Taurine/Creatinine|Taurine/Creatinine
C1715641|T201|COMP|44413-3|LNC|Threonine/Creatinine|Threonine/Creatinine
C1715642|T201|COMP|44414-1|LNC|Tryptophan/Creatinine|Tryptophan/Creatinine
C1715643|T201|COMP|44415-8|LNC|Tyrosine/Creatinine|Tyrosine/Creatinine
C1715644|T201|COMP|44416-6|LNC|Urea nitrogen/Creatinine|Urea nitrogen/Creatinine
C1715645|T201|COMP|44417-4|LNC|Valine/Creatinine|Valine/Creatinine
C1715646|T201|COMP|44418-2|LNC|Vanillylmandelate/Creatine|Vanillylmandelate/Creatine
C1715647|T201|COMP|44420-8|LNC|CACNA1A gene targeted mutation analysis|CACNA1A gene targeted mutation analysis
C1715648|T201|COMP|44422-4|LNC|Interleukin 2 receptor alpha chain.soluble|Interleukin 2 receptor alpha chain.soluble
C1715649|T201|COMP|44423-2|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C1715650|T201|COMP|44424-0|LNC|Methylenedioxymethamphetamine/Creatinine|Methylenedioxymethamphetamine/Creatinine
C1715652|T201|COMP|44426-5|LNC|3-Hydroxyphenylacetate/Creatinine|3-Hydroxyphenylacetate/Creatinine
C1715653|T201|COMP|44427-3|LNC|3-Hydroxyphenylacetate/Creatinine|3-Hydroxyphenylacetate/Creatinine
C1715655|T201|COMP|44429-9|LNC|Albumin/Globulin|Albumin/Globulin
C1715656|T201|COMP|44430-7|LNC|Alpha cortolone/Creatinine|Alpha cortolone/Creatinine
C1715657|T201|COMP|44431-5|LNC|Annexin V Ab.IgG|Annexin V Ab.IgG
C1715658|T201|COMP|44432-3|LNC|Annexin V Ab.IgM|Annexin V Ab.IgM
C1715659|T201|COMP|44433-1|LNC|Antibiotic XXX^peak|Antibiotic XXX^peak
C1715660|T201|COMP|44434-9|LNC|Antibiotic XXX^trough|Antibiotic XXX^trough
C1715661|T201|COMP|44435-6|LNC|Ascaris lumbricoides adult Ab.IgG|Ascaris lumbricoides adult Ab.IgG
C1715662|T201|COMP|44436-4|LNC|Ascaris lumbricoides larva Ab.IgG|Ascaris lumbricoides larva Ab.IgG
C1715663|T201|COMP|44438-0|LNC|Aspergillus fumigatus 1 Ab|Aspergillus fumigatus 1 Ab
C1715664|T201|COMP|44439-8|LNC|Aspergillus fumigatus 3 Ab|Aspergillus fumigatus 3 Ab
C1715665|T201|COMP|44440-6|LNC|Aspergillus fumigatus 6 Ab|Aspergillus fumigatus 6 Ab
C1715666|T201|COMP|44441-4|LNC|Aspergillus niger Ab|Aspergillus niger Ab
C1715667|T201|COMP|44442-2|LNC|Bartonella henselae Ab|Bartonella henselae Ab
C1715668|T201|COMP|44443-0|LNC|Bartonella sp Ab.IgG|Bartonella sp Ab.IgG
C1715669|T201|COMP|44444-8|LNC|Bartonella sp Ab.IgM|Bartonella sp Ab.IgM
C1715670|T201|COMP|44445-5|LNC|Basement membrane Ab.IgA|Basement membrane Ab.IgA
C1715671|T201|COMP|44446-3|LNC|Basement membrane Ab.IgG|Basement membrane Ab.IgG
C1715672|T201|COMP|44447-1|LNC|Beta 2 glycoprotein 1 Ab.IgA|Beta 2 glycoprotein 1 Ab.IgA
C1715673|T201|COMP|44449-7|LNC|Beta 2 glycoprotein 1 Ab.IgM|Beta 2 glycoprotein 1 Ab.IgM
C1715674|T201|COMP|44450-5|LNC|Beta cortolone/Creatinine|Beta cortolone/Creatinine
C1715675|T201|COMP|44451-3|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C1715676|T201|COMP|44452-1|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C1715677|T201|COMP|44453-9|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C1715678|T201|COMP|44454-7|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C1715679|T201|COMP|44456-2|LNC|Borrelia burgdorferi Ab^1st specimen|Borrelia burgdorferi Ab^1st specimen
C1715680|T201|COMP|44457-0|LNC|Borrelia sp Ab|Borrelia sp Ab
C1715681|T201|COMP|44458-8|LNC|Brucella abortus Ab.IgG+IgM|Brucella abortus Ab.IgG+IgM
C1715683|T201|COMP|44460-4|LNC|Cladosporium herbarum Ab|Cladosporium herbarum Ab
C1715684|T201|COMP|44461-2|LNC|Dermatophagoides farinae Ab|Dermatophagoides farinae Ab
C1715685|T201|COMP|44462-0|LNC|Insulin.free+Bound|Insulin.free+Bound
C1715686|T201|COMP|44464-6|LNC|Herpes simplex virus 1|Herpes simplex virus 1
C1715687|T201|COMP|44465-3|LNC|Herpes simplex virus 1|Herpes simplex virus 1
C1715688|T201|COMP|44466-1|LNC|Herpes simplex virus 1|Herpes simplex virus 1
C1715689|T201|COMP|44467-9|LNC|Herpes simplex virus 1|Herpes simplex virus 1
C1715690|T201|COMP|44468-7|LNC|Herpes simplex virus 1|Herpes simplex virus 1
C1715691|T201|COMP|44470-3|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1715692|T201|COMP|44471-1|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1715693|T201|COMP|44472-9|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1715694|T201|COMP|44473-7|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1715695|T201|COMP|44474-5|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1715696|T201|COMP|44475-2|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1715697|T201|COMP|44476-0|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1715698|T201|COMP|44477-8|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C1715699|T201|COMP|44478-6|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C1715700|T201|COMP|44479-4|LNC|Herpes simplex virus 1+2 Ab|Herpes simplex virus 1+2 Ab
C1715701|T201|COMP|44480-2|LNC|Herpes simplex virus 1+2 Ab|Herpes simplex virus 1+2 Ab
C1715702|T201|COMP|44481-0|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C1715703|T201|COMP|44482-8|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C1715704|T201|COMP|44483-6|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1715705|T201|COMP|44484-4|LNC|Herpes simplex virus 2|Herpes simplex virus 2
C1715706|T201|COMP|44485-1|LNC|Herpes simplex virus 2|Herpes simplex virus 2
C1715707|T201|COMP|44486-9|LNC|Herpes simplex virus 2|Herpes simplex virus 2
C1715708|T201|COMP|44488-5|LNC|Herpes simplex virus 2|Herpes simplex virus 2
C1715709|T201|COMP|44489-3|LNC|Herpes simplex virus 2|Herpes simplex virus 2
C1715710|T201|COMP|44490-1|LNC|Herpes simplex virus 2|Herpes simplex virus 2
C1715711|T201|COMP|44491-9|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C1715712|T201|COMP|44492-7|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C1715713|T201|COMP|44493-5|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C1715714|T201|COMP|44494-3|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C1715715|T201|COMP|44495-0|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1715716|T201|COMP|44496-8|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1715717|T201|COMP|44497-6|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1715718|T201|COMP|44498-4|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1715719|T201|COMP|44499-2|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1715720|T201|COMP|44500-7|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1715721|T201|COMP|44501-5|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1715722|T201|COMP|44502-3|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C1715723|T201|COMP|44503-1|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C1715724|T201|COMP|44504-9|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C1715725|T201|COMP|44505-6|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C1715726|T201|COMP|44506-4|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C1715727|T201|COMP|44507-2|LNC|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C1715728|T201|COMP|44508-0|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1715729|T201|COMP|44509-8|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1715730|T201|COMP|44510-6|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1715731|T201|COMP|44511-4|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1715732|T201|COMP|44512-2|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1715733|T201|COMP|44513-0|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1715734|T201|COMP|44514-8|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1715735|T201|COMP|44515-5|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1715736|T201|COMP|44517-1|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C1715737|T201|COMP|44518-9|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C1715738|T201|COMP|44519-7|LNC|Herpes virus 6 Ab|Herpes virus 6 Ab
C1715739|T201|COMP|44520-5|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C1715740|T201|COMP|44522-1|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C1715741|T201|COMP|44523-9|LNC|Histoplasma capsulatum Ab.IgG|Histoplasma capsulatum Ab.IgG
C1715742|T201|COMP|44524-7|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1715743|T201|COMP|44525-4|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1715744|T201|COMP|44526-2|LNC|Histoplasma capsulatum H Ab|Histoplasma capsulatum H Ab
C1715745|T201|COMP|44527-0|LNC|Histoplasma capsulatum H Ab|Histoplasma capsulatum H Ab
C1715746|T201|COMP|44528-8|LNC|Histoplasma capsulatum M Ab|Histoplasma capsulatum M Ab
C1715747|T201|COMP|44529-6|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C1715748|T201|COMP|44530-4|LNC|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C1715749|T201|COMP|44531-2|LNC|HIV 1 Ag|HIV 1 Ag
C1715750|T201|COMP|44532-0|LNC|HIV 1 gp120 Ab|HIV 1 gp120 Ab
C1715751|T201|COMP|44533-8|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C1715752|T201|COMP|44535-3|LNC|HTLV I Ab|HTLV I Ab
C1715753|T201|COMP|44536-1|LNC|HTLV I DNA|HTLV I DNA
C1715754|T201|COMP|44538-7|LNC|HTLV I+II Ab|HTLV I+II Ab
C1715755|T201|COMP|44539-5|LNC|HTLV II Ab|HTLV II Ab
C1715756|T201|COMP|44540-3|LNC|HTLV II Ab.IgG|HTLV II Ab.IgG
C1715757|T201|COMP|44541-1|LNC|HTLV II DNA|HTLV II DNA
C1715758|T201|COMP|44542-9|LNC|HTLV II DNA|HTLV II DNA
C1715759|T201|COMP|44543-7|LNC|Human papilloma virus 31+33 Ag|Human papilloma virus 31+33 Ag
C1715760|T201|COMP|44544-5|LNC|Human papilloma virus 35 Ag|Human papilloma virus 35 Ag
C1715761|T201|COMP|44545-2|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C1715762|T201|COMP|44546-0|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C1715763|T201|COMP|44547-8|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C1715764|T201|COMP|44548-6|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C1715765|T201|COMP|44549-4|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C1715766|T201|COMP|44550-2|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C1715767|T201|COMP|44551-0|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C1715768|T201|COMP|44552-8|LNC|hydroCHLOROthiazide|hydroCHLOROthiazide
C1715769|T201|COMP|44553-6|LNC|Hydroxyitraconazole|Hydroxyitraconazole
C1715770|T201|COMP|44555-1|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C1715771|T201|COMP|44556-9|LNC|Influenza virus A Ab|Influenza virus A Ab
C1715772|T201|COMP|44557-7|LNC|Influenza virus A Ab|Influenza virus A Ab
C1715773|T201|COMP|44558-5|LNC|Influenza virus A Ag|Influenza virus A Ag
C1715774|T201|COMP|44559-3|LNC|Influenza virus A Ag|Influenza virus A Ag
C1715775|T201|COMP|44560-1|LNC|Influenza virus A Ag|Influenza virus A Ag
C1715776|T201|COMP|44561-9|LNC|Influenza virus A Ag|Influenza virus A Ag
C1715777|T201|COMP|44562-7|LNC|Influenza virus A Ag|Influenza virus A Ag
C1715778|T201|COMP|44563-5|LNC|Influenza virus A Ag|Influenza virus A Ag
C1715779|T201|COMP|44564-3|LNC|Influenza virus A Ag|Influenza virus A Ag
C1715780|T201|COMP|44565-0|LNC|Influenza virus A+B Ab|Influenza virus A+B Ab
C1715781|T201|COMP|44566-8|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C1715782|T201|COMP|44567-6|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C1715783|T201|COMP|44568-4|LNC|Influenza virus B Ab|Influenza virus B Ab
C1715784|T201|COMP|44569-2|LNC|Influenza virus B Ab|Influenza virus B Ab
C1715785|T201|COMP|44669-0|LNC|Margin involvement|Margin involvement
C1715786|T201|COMP|44671-6|LNC|Margin involvement|Margin involvement
C1715787|T201|COMP|44673-2|LNC|DCIS.uninvolved margin distance.closest|DCIS.uninvolved margin distance.closest
C1715788|T201|COMP|44674-0|LNC|Invasive carcinoma.uninvolved margin.closest|Invasive carcinoma.uninvolved margin.closest
C1715789|T201|COMP|44675-7|LNC|DCIS.uninvolved margin.closest|DCIS.uninvolved margin.closest
C1715790|T201|COMP|44676-5|LNC|Margin(s) involved by invasive carcinoma|Margin(s) involved by invasive carcinoma
C1715791|T201|COMP|44677-3|LNC|Margin(s) involved by DCIS|Margin(s) involved by DCIS
C1715796|T201|COMP|44768-0|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C1715797|T201|COMP|44769-8|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C1715798|T201|COMP|44770-6|LNC|Neuronal nuclear Ab.IgG|Neuronal nuclear Ab.IgG
C1715799|T201|COMP|44771-4|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C1715800|T201|COMP|45181-5|LNC|19q chromosome deletion|19q chromosome deletion
C1715801|T201|COMP|45182-3|LNC|HIV phenotype|HIV phenotype
C1715802|T201|COMP|45183-1|LNC|Neisseria meningitidis|Neisseria meningitidis
C1715803|T201|COMP|45184-9|LNC|11-Deoxycortisol/Cortisol|11-Deoxycortisol/Cortisol
C1715804|T201|COMP|45185-6|LNC|2-Oxo-3-Hydroxy-Lysergate diethylamide|2-Oxo-3-Hydroxy-Lysergate diethylamide
C1715805|T201|COMP|45186-4|LNC|Actinidia chinensis Ab.IgE/IgE.total|Actinidia chinensis Ab.IgE/IgE.total
C1715806|T201|COMP|45187-2|LNC|Antibiotic XXX|Antibiotic XXX
C1715807|T201|COMP|45188-0|LNC|Basement membrane zone BP180 Ab|Basement membrane zone BP180 Ab
C1715808|T201|COMP|45358-9|LNC|Length of calorie fast|Length of calorie fast
C1715809|T201|COMP|45359-7|LNC|Length of time post dose|Length of time post dose
C1715831|T201|COMP|46110-3|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C1715832|T201|COMP|46111-1|LNC|Mycoplasma sp DNA|Mycoplasma sp DNA
C1715833|T201|COMP|46112-9|LNC|Borrelia burgdorferi 18kD Ab.IgG|Borrelia burgdorferi 18kD Ab.IgG
C1715834|T201|COMP|46113-7|LNC|Borrelia burgdorferi 23kD Ab.IgM|Borrelia burgdorferi 23kD Ab.IgM
C1715835|T201|COMP|46114-5|LNC|Borrelia burgdorferi 23kD Ab.IgG|Borrelia burgdorferi 23kD Ab.IgG
C1715836|T201|COMP|46115-2|LNC|Borrelia burgdorferi 28kD Ab.IgG|Borrelia burgdorferi 28kD Ab.IgG
C1715837|T201|COMP|46116-0|LNC|Borrelia burgdorferi 30kD Ab.IgG|Borrelia burgdorferi 30kD Ab.IgG
C1715838|T201|COMP|46117-8|LNC|Borrelia burgdorferi 39kD Ab.IgM|Borrelia burgdorferi 39kD Ab.IgM
C1715839|T201|COMP|46118-6|LNC|Borrelia burgdorferi 39kD Ab.IgG|Borrelia burgdorferi 39kD Ab.IgG
C1715840|T201|COMP|44570-0|LNC|Influenza virus B Ab|Influenza virus B Ab
C1715841|T201|COMP|44571-8|LNC|Influenza virus B Ag|Influenza virus B Ag
C1715842|T201|COMP|44572-6|LNC|Influenza virus B Ag|Influenza virus B Ag
C1715843|T201|COMP|44573-4|LNC|Influenza virus B Ag|Influenza virus B Ag
C1715844|T201|COMP|44574-2|LNC|Influenza virus B Ag|Influenza virus B Ag
C1715845|T201|COMP|44575-9|LNC|Influenza virus B Ag|Influenza virus B Ag
C1715846|T201|COMP|44576-7|LNC|Influenza virus B Ag|Influenza virus B Ag
C1715847|T201|COMP|44577-5|LNC|Influenza virus B Ag|Influenza virus B Ag
C1715848|T201|COMP|44578-3|LNC|Influenza virus C Ab|Influenza virus C Ab
C1715849|T201|COMP|44579-1|LNC|Influenza virus C Ab|Influenza virus C Ab
C1715850|T201|COMP|44580-9|LNC|HTLV I+II p21 env Ab|HTLV I+II p21 env Ab
C1715851|T201|COMP|44581-7|LNC|HTLV I+II p38 tax Ab|HTLV I+II p38 tax Ab
C1715852|T201|COMP|44582-5|LNC|IgA|IgA
C1715853|T201|COMP|44583-3|LNC|IgA Ab|IgA Ab
C1715854|T201|COMP|44584-1|LNC|IgA Ab|IgA Ab
C1715855|T201|COMP|44585-8|LNC|IgA Ab.IgG|IgA Ab.IgG
C1715856|T201|COMP|44586-6|LNC|IgA Ab.IgM|IgA Ab.IgM
C1715857|T201|COMP|44587-4|LNC|IgA.monoclonal|IgA.monoclonal
C1715858|T201|COMP|44588-2|LNC|IgA.monoclonal|IgA.monoclonal
C1715859|T201|COMP|44589-0|LNC|IgA.monoclonal|IgA.monoclonal
C1715860|T201|COMP|44590-8|LNC|IgA.secretory|IgA.secretory
C1715861|T201|COMP|44591-6|LNC|IgD|IgD
C1715862|T201|COMP|44592-4|LNC|IgD|IgD
C1715863|T201|COMP|44594-0|LNC|IgE|IgE
C1715864|T201|COMP|44596-5|LNC|IgG Ag|IgG Ag
C1715865|T201|COMP|44597-3|LNC|IgG.monoclonal|IgG.monoclonal
C1715866|T201|COMP|44598-1|LNC|IgG.monoclonal|IgG.monoclonal
C1715867|T201|COMP|44599-9|LNC|IgG.monoclonal|IgG.monoclonal
C1715868|T201|COMP|44600-5|LNC|IgM|IgM
C1715869|T201|COMP|44601-3|LNC|IgM.monoclonal|IgM.monoclonal
C1715870|T201|COMP|44602-1|LNC|IgM.monoclonal|IgM.monoclonal
C1715871|T201|COMP|44603-9|LNC|IgM.monoclonal|IgM.monoclonal
C1715872|T201|COMP|44604-7|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C1715873|T201|COMP|44605-4|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C1715874|T201|COMP|44606-2|LNC|ALOX3+ALOX12B gene targeted mutation analysis|ALOX3+ALOX12B gene targeted mutation analysis
C1715875|T201|COMP|44607-0|LNC|HIV 1|HIV 1
C1715876|T201|COMP|44608-8|LNC|KCNQ1 gene mutations tested for|KCNQ1 gene mutations tested for
C1715884|T201|COMP|44617-9|LNC|PWS gene targeted mutation analysis|PWS gene targeted mutation analysis
C1715885|T201|COMP|44618-7|LNC|Total linear mm of carcinoma|Total linear mm of carcinoma
C1715886|T201|COMP|44619-5|LNC|Length of tissue core(s)|Length of tissue core(s)
C1715887|T201|COMP|44620-3|LNC|Other quantitation|Other quantitation
C1715888|T201|COMP|44621-1|LNC|Regional lymph nodes examined|Regional lymph nodes examined
C1715889|T201|COMP|44622-9|LNC|Regional lymph nodes containing metastases|Regional lymph nodes containing metastases
C1715890|T201|COMP|44623-7|LNC|Matted nodes|Matted nodes
C1715891|T201|COMP|44624-5|LNC|Additional pathological findings|Additional pathological findings
C1715892|T201|COMP|44626-0|LNC|Seminal vesicle invasion|Seminal vesicle invasion
C1715893|T201|COMP|44627-8|LNC|Extraprostatic extension|Extraprostatic extension
C1715894|T201|COMP|44628-6|LNC|Reason specimen size cannot be determined|Reason specimen size cannot be determined
C1715895|T201|COMP|44629-4|LNC|Specimen size.max dimension|Specimen size.max dimension
C1715896|T201|COMP|44630-2|LNC|Specimen size.additional dimension 1|Specimen size.additional dimension 1
C1715897|T201|COMP|44631-0|LNC|Specimen size.additional dimension 2|Specimen size.additional dimension 2
C1715898|T201|COMP|44632-8|LNC|Satellite nodule presence|Satellite nodule presence
C1715899|T201|COMP|44633-6|LNC|Tumor pigmentation|Tumor pigmentation
C1715901|T201|COMP|44635-1|LNC|Invasive component size.max.dimension|Invasive component size.max.dimension
C1715902|T201|COMP|44636-9|LNC|Invasive component size.additional dimension 1|Invasive component size.additional dimension 1
C1715903|T201|COMP|44637-7|LNC|Invasive component size.additional dimension 2|Invasive component size.additional dimension 2
C1715904|T201|COMP|44638-5|LNC|Histologic type|Histologic type
C1715905|T201|COMP|44639-3|LNC|Histologic type|Histologic type
C1715906|T201|COMP|44641-9|LNC|Gleason pattern.primary|Gleason pattern.primary
C1715907|T201|COMP|44642-7|LNC|Gleason pattern.secondary|Gleason pattern.secondary
C1715908|T201|COMP|44643-5|LNC|Gleason pattern.tertiary|Gleason pattern.tertiary
C1715909|T201|COMP|44644-3|LNC|Tubule formation|Tubule formation
C1715910|T201|COMP|44645-0|LNC|Nuclear pleomorphism|Nuclear pleomorphism
C1715911|T201|COMP|44646-8|LNC|Nottingham mitotic count.25x obj|Nottingham mitotic count.25x obj
C1715912|T201|COMP|44647-6|LNC|Nottingham mitotic count.40x obj|Nottingham mitotic count.40x obj
C1715913|T201|COMP|44648-4|LNC|Histologic grade|Histologic grade
C1715914|T201|COMP|44649-2|LNC|Grading system|Grading system
C1715915|T201|COMP|44650-0|LNC|Mitotic count per 10 HPF|Mitotic count per 10 HPF
C1715916|T201|COMP|44651-8|LNC|Tissue cores.positive.carcinoma|Tissue cores.positive.carcinoma
C1715917|T201|COMP|44652-6|LNC|Total number of cores|Total number of cores
C1715918|T201|COMP|44653-4|LNC|Tumor quantitation.incidental|Tumor quantitation.incidental
C1715919|T201|COMP|44654-2|LNC|Prostatic tissue involved by tumor|Prostatic tissue involved by tumor
C1715920|T201|COMP|44655-9|LNC|Tissue chips.positive.carcinoma|Tissue chips.positive.carcinoma
C1715921|T201|COMP|44656-7|LNC|Number of tissue chips|Number of tissue chips
C1715922|T201|COMP|44657-5|LNC|Dominant nodule.max.dimension|Dominant nodule.max.dimension
C1715923|T201|COMP|44658-3|LNC|Dominant nodule.additional dimension 1|Dominant nodule.additional dimension 1
C1715924|T201|COMP|44660-9|LNC|Tumor involved by ulceration|Tumor involved by ulceration
C1715925|T201|COMP|44661-7|LNC|Depth of invasion by tumor|Depth of invasion by tumor
C1715927|T201|COMP|44663-3|LNC|T classification|T classification
C1715928|T201|COMP|44664-1|LNC|T classification|T classification
C1715929|T201|COMP|44665-8|LNC|T classification|T classification
C1715930|T201|COMP|44666-6|LNC|M stage of distant metastasis|M stage of distant metastasis
C1715931|T201|COMP|44667-4|LNC|Site of distant metastasis|Site of distant metastasis
C1715932|T201|COMP|44668-2|LNC|M stage of distant metastasis|M stage of distant metastasis
C1715933|T201|COMP|44679-9|LNC|Margin(s) involved by invasive melanoma|Margin(s) involved by invasive melanoma
C1715934|T201|COMP|44680-7|LNC|Margin(s) involved by melanoma in situ|Margin(s) involved by melanoma in situ
C1715935|T201|COMP|44681-5|LNC|Invasive melanoma.uninvolved margin.closest|Invasive melanoma.uninvolved margin.closest
C1715946|T201|COMP|44692-2|LNC|Microcalcifications|Microcalcifications
C1715947|T201|COMP|44693-0|LNC|Tumor infiltrating lymphocytes|Tumor infiltrating lymphocytes
C1715948|T201|COMP|44694-8|LNC|Tumor regression|Tumor regression
C1715949|T201|COMP|44695-5|LNC|Mitotic index|Mitotic index
C1715950|T201|COMP|44696-3|LNC|Inflammation type|Inflammation type
C1715951|T201|COMP|44697-1|LNC|Lesion size.max.dimension|Lesion size.max.dimension
C1715952|T201|COMP|44698-9|LNC|Lesion size.additional dimension 1|Lesion size.additional dimension 1
C1715953|T201|COMP|44699-7|LNC|Extent of margin involvement|Extent of margin involvement
C1715954|T201|COMP|44700-3|LNC|ACTA1 gene targeted mutation analysis|ACTA1 gene targeted mutation analysis
C1715955|T201|COMP|44701-1|LNC|BHD gene targeted mutation analysis|BHD gene targeted mutation analysis
C1715956|T201|COMP|44703-7|LNC|MC4R gene targeted mutation analysis|MC4R gene targeted mutation analysis
C1715957|T201|COMP|44704-5|LNC|NEB gene targeted mutation analysis|NEB gene targeted mutation analysis
C1715958|T201|COMP|44705-2|LNC|ALS4 gene targeted mutation analysis|ALS4 gene targeted mutation analysis
C1715959|T201|COMP|44706-0|LNC|Actin.smooth muscle Ab.IgG|Actin.smooth muscle Ab.IgG
C1715960|T201|COMP|44707-8|LNC|Albumin/Creatinine|Albumin/Creatinine
C1715961|T201|COMP|44708-6|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C1715962|T201|COMP|44709-4|LNC|Asialoganglioside GM1 Ab.IgM|Asialoganglioside GM1 Ab.IgM
C1715963|T201|COMP|44710-2|LNC|Carnitine/Acylcarnitine|Carnitine/Acylcarnitine
C1715964|T201|COMP|44711-0|LNC|Cholesterol.in LDL/Apolipoprotein B|Cholesterol.in LDL/Apolipoprotein B
C1715965|T201|COMP|44712-8|LNC|Collagen crosslinked N-telopeptide/Creatinine|Collagen crosslinked N-telopeptide/Creatinine
C1715966|T201|COMP|44713-6|LNC|Collagen crosslinked N-telopeptide/Creatinine|Collagen crosslinked N-telopeptide/Creatinine
C1715967|T201|COMP|44714-4|LNC|Complement C3/Protein|Complement C3/Protein
C1715968|T201|COMP|44715-1|LNC|Complement C4/Protein|Complement C4/Protein
C1715969|T201|COMP|44716-9|LNC|Creatinine/Calcium|Creatinine/Calcium
C1715970|T201|COMP|44717-7|LNC|Lipoprotein.beta/Lipoprotein.alpha|Lipoprotein.beta/Lipoprotein.alpha
C1715971|T201|COMP|44719-3|LNC|Methylmalonate/Homocysteine|Methylmalonate/Homocysteine
C1715972|T201|COMP|44720-1|LNC|Methylmalonate/Homocystine|Methylmalonate/Homocystine
C1715973|T201|COMP|44721-9|LNC|Histiocytes|Histiocytes
C1715974|T201|COMP|44722-7|LNC|Histiocytes|Histiocytes
C1715975|T201|COMP|44748-2|LNC|La Crosse virus Ab|La Crosse virus Ab
C1715976|T201|COMP|44749-0|LNC|Ganglioside GM1 Ab.IgA|Ganglioside GM1 Ab.IgA
C1715977|T201|COMP|44750-8|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C1715978|T201|COMP|44751-6|LNC|Nuclear Ab|Nuclear Ab
C1715979|T201|COMP|44752-4|LNC|Nuclear Ab|Nuclear Ab
C1715980|T201|COMP|44753-2|LNC|Sulfatide Ab.IgM|Sulfatide Ab.IgM
C1715981|T201|COMP|44754-0|LNC|Hepatitis D virus Ag|Hepatitis D virus Ag
C1715982|T201|COMP|44755-7|LNC|Hepatitis D virus Ag|Hepatitis D virus Ag
C1715984|T201|COMP|44757-3|LNC|Blood product units given|Blood product units given
C1716000|T201|COMP|44783-9|LNC|Sodium|Sodium
C1716001|T201|COMP|44784-7|LNC|Creatinine|Creatinine
C1716002|T201|COMP|44785-4|LNC|Alanine aminotransferase|Alanine aminotransferase
C1716003|T201|COMP|44786-2|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C1716005|T201|COMP|44789-6|LNC|Amylase & Creatinine clearance panel|Amylase & Creatinine clearance panel
C1716006|T201|COMP|44790-4|LNC|Iodide|Iodide
C1716007|T201|COMP|44791-2|LNC|Menorrhagia coagulation panel|Menorrhagia coagulation panel
C1716008|T201|COMP|44792-0|LNC|Immunoglobulin light chains panel|Immunoglobulin light chains panel
C1716009|T201|COMP|44793-8|LNC|Immunoglobulin light chains panel|Immunoglobulin light chains panel
C1716010|T201|COMP|44794-6|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C1716011|T201|COMP|44795-3|LNC|Influenza virus A H5 Asian RNA|Influenza virus A H5 Asian RNA
C1716012|T201|COMP|44796-1|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C1716013|T201|COMP|44797-9|LNC|Brucella sp|Brucella sp
C1716014|T201|COMP|44798-7|LNC|Burkholderia sp identified|Burkholderia sp identified
C1716015|T201|COMP|44799-5|LNC|Coxiella burnetii|Coxiella burnetii
C1716016|T201|COMP|44801-9|LNC|Aldolase|Aldolase
C1716017|T201|COMP|44802-7|LNC|Enolase.neuron specific|Enolase.neuron specific
C1716018|T201|COMP|44804-3|LNC|Taenia solium Ab.IgG|Taenia solium Ab.IgG
C1716019|T201|COMP|44805-0|LNC|BK virus DNA|BK virus DNA
C1716020|T201|COMP|44806-8|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae DNA|Chlamydia trachomatis+Neisseria gonorrhoeae DNA
C1716021|T201|COMP|44807-6|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae DNA|Chlamydia trachomatis+Neisseria gonorrhoeae DNA
C1716022|T201|COMP|44808-4|LNC|Histoplasma capsulatum H Ab band pattern|Histoplasma capsulatum H Ab band pattern
C1716023|T201|COMP|44809-2|LNC|Histoplasma capsulatum M Ab band pattern|Histoplasma capsulatum M Ab band pattern
C1716024|T201|COMP|44810-0|LNC|HTLV I gp21e Ab|HTLV I gp21e Ab
C1716025|T201|COMP|44811-8|LNC|Coccidioides sp Ab.IgA|Coccidioides sp Ab.IgA
C1716026|T201|COMP|44812-6|LNC|Yeast.hyphae|Yeast.hyphae
C1716027|T201|COMP|44813-4|LNC|Hepatitis C virus c22p Ab|Hepatitis C virus c22p Ab
C1716028|T201|COMP|44814-2|LNC|Coxiella burnetii phase 2 Ab.IgM|Coxiella burnetii phase 2 Ab.IgM
C1716029|T201|COMP|44815-9|LNC|Brucella abortus Ab.IgM|Brucella abortus Ab.IgM
C1716030|T201|COMP|44816-7|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C1716031|T201|COMP|44817-5|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C1716032|T201|COMP|44818-3|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C1716033|T201|COMP|44819-1|LNC|Leishmania donovani Ab.IgM|Leishmania donovani Ab.IgM
C1716034|T201|COMP|44820-9|LNC|Leishmania braziliensis Ab.IgM|Leishmania braziliensis Ab.IgM
C1716035|T201|COMP|44821-7|LNC|Leishmania braziliensis Ab.IgG|Leishmania braziliensis Ab.IgG
C1716036|T201|COMP|44823-3|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C1716037|T201|COMP|44824-1|LNC|Leishmania donovani Ab.IgG|Leishmania donovani Ab.IgG
C1716038|T201|COMP|44825-8|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C1716039|T201|COMP|44826-6|LNC|Hepatitis D virus Ab.IgM|Hepatitis D virus Ab.IgM
C1716040|T201|COMP|44827-4|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C1716041|T201|COMP|44828-2|LNC|Teriflunomide|Teriflunomide
C1716042|T201|COMP|44829-0|LNC|Acremonium sp Ab.IgG.RAST class|Acremonium sp Ab.IgG.RAST class
C1716043|T201|COMP|44830-8|LNC|Phosphorylase|Phosphorylase
C1716044|T201|COMP|44831-6|LNC|Hepatitis C virus c100p+5-1-1 Ab|Hepatitis C virus c100p+5-1-1 Ab
C1716045|T201|COMP|44832-4|LNC|Glycogen synthase I/Glycogen synthase.total|Glycogen synthase I/Glycogen synthase.total
C1716047|T201|COMP|44834-0|LNC|Acid phosphatase.tartrate resistant|Acid phosphatase.tartrate resistant
C1716048|T201|COMP|44835-7|LNC|Acid phosphatase.tartrate resistant|Acid phosphatase.tartrate resistant
C1716049|T201|COMP|44836-5|LNC|5-Hydroxymethyl-2-Furoate|5-Hydroxymethyl-2-Furoate
C1716050|T201|COMP|44837-3|LNC|Epinephrine+Norepinephrine|Epinephrine+Norepinephrine
C1716051|T201|COMP|44838-1|LNC|Catecholamines|Catecholamines
C1716052|T201|COMP|44840-7|LNC|Fungus identified^^^5|Fungus identified^^^5
C1716053|T201|COMP|44841-5|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1716054|T201|COMP|44842-3|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1716055|T201|COMP|44843-1|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1716056|T201|COMP|44844-9|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1716057|T201|COMP|44845-6|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1716058|T201|COMP|44846-4|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C1716059|T201|COMP|44847-2|LNC|Bacteria identified^^^7|Bacteria identified^^^7
C1716060|T201|COMP|44848-0|LNC|Bacteria identified^^^7|Bacteria identified^^^7
C1716061|T201|COMP|44849-8|LNC|Bacteria identified^^^8|Bacteria identified^^^8
C1716062|T201|COMP|44850-6|LNC|Bacteria identified^^^8|Bacteria identified^^^8
C1716063|T201|COMP|44851-4|LNC|Mycobacterium sp identified^^^2|Mycobacterium sp identified^^^2
C1716064|T201|COMP|44852-2|LNC|Mycobacterium sp identified^^^3|Mycobacterium sp identified^^^3
C1716065|T201|COMP|44853-0|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1716066|T201|COMP|44854-8|LNC|Mycobacterium sp identified^^^4|Mycobacterium sp identified^^^4
C1716067|T201|COMP|44855-5|LNC|Mycobacterium sp identified^^^5|Mycobacterium sp identified^^^5
C1716068|T201|COMP|44856-3|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1716069|T201|COMP|44858-9|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C1716070|T201|COMP|44859-7|LNC|Bacteria identified^^^7|Bacteria identified^^^7
C1716071|T201|COMP|44860-5|LNC|Methoxyacetate/Creatinine|Methoxyacetate/Creatinine
C1716075|T201|COMP|44865-4|LNC|Ammonium urate|Ammonium urate
C1716076|T201|COMP|44867-0|LNC|Iron.microscopic observation|Iron.microscopic observation
C1716077|T201|COMP|44868-8|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1716078|T201|COMP|44869-6|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C1716079|T201|COMP|44870-4|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1716080|T201|COMP|44871-2|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C1716081|T201|COMP|44872-0|LNC|HIV 1 p24 Ag|HIV 1 p24 Ag
C1716082|T201|COMP|44873-8|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C1716083|T201|COMP|44874-6|LNC|HTLV I+II RNA|HTLV I+II RNA
C1716084|T201|COMP|44875-3|LNC|IgM Ag|IgM Ag
C1716085|T201|COMP|44876-1|LNC|Influenza virus A Ab|Influenza virus A Ab
C1716086|T201|COMP|44878-7|LNC|Staphylococcus aureus enterotoxin A sea gene|Staphylococcus aureus enterotoxin A sea gene
C1716087|T201|COMP|44879-5|LNC|Staphylococcus aureus enterotoxin E see gene|Staphylococcus aureus enterotoxin E see gene
C1716088|T201|COMP|44880-3|LNC|Staphylococcus aureus enterotoxin B seb gene|Staphylococcus aureus enterotoxin B seb gene
C1716090|T201|COMP|44882-9|LNC|Malignant cells|Malignant cells
C1716091|T201|COMP|44883-7|LNC|Malignant cells|Malignant cells
C1716092|T201|COMP|44884-5|LNC|Malignant cells|Malignant cells
C1716093|T201|COMP|44885-2|LNC|Malignant cells|Malignant cells
C1716094|T201|COMP|44886-0|LNC|Malignant cells|Malignant cells
C1716095|T201|COMP|44887-8|LNC|Malignant cells|Malignant cells
C1716096|T201|COMP|44888-6|LNC|Malignant cells|Malignant cells
C1716097|T201|COMP|44889-4|LNC|Malignant cells|Malignant cells
C1716098|T201|COMP|44890-2|LNC|Malignant cells|Malignant cells
C1716099|T201|COMP|44891-0|LNC|Malignant cells|Malignant cells
C1716100|T201|COMP|44893-6|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716101|T201|COMP|44894-4|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716102|T201|COMP|44895-1|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716103|T201|COMP|44896-9|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716104|T201|COMP|44897-7|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716105|T201|COMP|44898-5|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716106|T201|COMP|44899-3|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716107|T201|COMP|44900-9|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716108|T201|COMP|44901-7|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716109|T201|COMP|44902-5|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716110|T201|COMP|44903-3|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716111|T201|COMP|44904-1|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716112|T201|COMP|44905-8|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1716113|T201|COMP|44906-6|LNC|Homovanillate panel|Homovanillate panel
C1716114|T201|COMP|44907-4|LNC|5-Hydroxyindoleacetate panel|5-Hydroxyindoleacetate panel
C1716115|T201|COMP|44908-2|LNC|Homovanillate & Creatinine|Homovanillate & Creatinine
C1716116|T201|COMP|44909-0|LNC|5-Hydroxyindoleacetate & Creatinine|5-Hydroxyindoleacetate & Creatinine
C1716117|T201|COMP|44910-8|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C1716118|T201|COMP|44911-6|LNC|Beta 2 globulin+Gamma globulin|Beta 2 globulin+Gamma globulin
C1716119|T201|COMP|44912-4|LNC|Beta 2 globulin+Gamma globulin/Protein.total|Beta 2 globulin+Gamma globulin/Protein.total
C1716120|T201|COMP|44913-2|LNC|Beta globulin+Gamma globulin|Beta globulin+Gamma globulin
C1716121|T201|COMP|44915-7|LNC|Cholesterol.in LDL/Cholesterol.in HDL|Cholesterol.in LDL/Cholesterol.in HDL
C1716122|T201|COMP|44916-5|LNC|Cortisol^pre XXX challenge|Cortisol^pre XXX challenge
C1716123|T201|COMP|44917-3|LNC|Cortisol^post dose dexamethasone|Cortisol^post dose dexamethasone
C1716124|T201|COMP|44918-1|LNC|DOPamine/Creatinine|DOPamine/Creatinine
C1716125|T201|COMP|44919-9|LNC|Glucose^1.5H post meal|Glucose^1.5H post meal
C1716126|T201|COMP|44920-7|LNC|Hemoglobin C/Hemoglobin.total|Hemoglobin C/Hemoglobin.total
C1716127|T201|COMP|44921-5|LNC|Hemoglobin D/Hemoglobin.total|Hemoglobin D/Hemoglobin.total
C1716128|T201|COMP|44922-3|LNC|Hemoglobin E/Hemoglobin.total|Hemoglobin E/Hemoglobin.total
C1716129|T201|COMP|44923-1|LNC|Hemoglobin S/Hemoglobin.total|Hemoglobin S/Hemoglobin.total
C1716130|T201|COMP|44924-9|LNC|Normetanephrine/Creatinine|Normetanephrine/Creatinine
C1716131|T201|COMP|44926-4|LNC|Prolactin^1.5H post dose TRH IV|Prolactin^1.5H post dose TRH IV
C1716132|T201|COMP|44927-2|LNC|Prolactin^30M post dose TRH IV|Prolactin^30M post dose TRH IV
C1716133|T201|COMP|44928-0|LNC|Prolactin^15M pre dose TRH IV|Prolactin^15M pre dose TRH IV
C1716134|T201|COMP|44930-6|LNC|Prolactin^2H post dose TRH IV|Prolactin^2H post dose TRH IV
C1716135|T201|COMP|44931-4|LNC|Prolactin^pre dose TRH IV|Prolactin^pre dose TRH IV
C1716136|T201|COMP|44932-2|LNC|Protein.monoclonal band 2/Protein.total|Protein.monoclonal band 2/Protein.total
C1716137|T201|COMP|44933-0|LNC|Specific gravity|Specific gravity
C1716138|T201|COMP|44934-8|LNC|Thymidine kinase|Thymidine kinase
C1716139|T201|COMP|44935-5|LNC|Thyrotropin^15M post dose TRH IV|Thyrotropin^15M post dose TRH IV
C1716140|T201|COMP|44936-3|LNC|Thyrotropin^15M pre dose TRH IV|Thyrotropin^15M pre dose TRH IV
C1716141|T201|COMP|44938-9|LNC|Hepatitis D virus Ab.IgM|Hepatitis D virus Ab.IgM
C1716148|T201|COMP|44945-4|LNC|Australian cervix cytology code|Australian cervix cytology code
C1716149|T201|COMP|44946-2|LNC|Borrelia burgdorferi 31kD Ab.IgG|Borrelia burgdorferi 31kD Ab.IgG
C1716150|T201|COMP|44994-2|LNC|Chlamydia trachomatis B Ab.IgM|Chlamydia trachomatis B Ab.IgM
C1716151|T201|COMP|44995-9|LNC|Chlamydia trachomatis B Ab.IgG|Chlamydia trachomatis B Ab.IgG
C1716152|T201|COMP|44996-7|LNC|Chlamydia trachomatis B Ab.IgA|Chlamydia trachomatis B Ab.IgA
C1716153|T201|COMP|44997-5|LNC|Chlamydia trachomatis Ab^2nd specimen|Chlamydia trachomatis Ab^2nd specimen
C1716154|T201|COMP|44998-3|LNC|Chlamydia trachomatis Ab^1st specimen|Chlamydia trachomatis Ab^1st specimen
C1716155|T201|COMP|44999-1|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C1716156|T201|COMP|45000-7|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C1716157|T201|COMP|45001-5|LNC|Chlamydia trachomatis Ab.IgM|Chlamydia trachomatis Ab.IgM
C1716158|T201|COMP|45002-3|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C1716159|T201|COMP|45003-1|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C1716160|T201|COMP|45004-9|LNC|Chlamydia trachomatis Ab.IgA|Chlamydia trachomatis Ab.IgA
C1716161|T201|COMP|45005-6|LNC|Chlamydia trachomatis Ab.IgA|Chlamydia trachomatis Ab.IgA
C1716162|T201|COMP|45007-2|LNC|Chlamydia trachomatis Ab|Chlamydia trachomatis Ab
C1716163|T201|COMP|45008-0|LNC|Chlamydia trachomatis Ab|Chlamydia trachomatis Ab
C1716164|T201|COMP|45009-8|LNC|Chlamydia trachomatis Ab|Chlamydia trachomatis Ab
C1716165|T201|COMP|45010-6|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C1716166|T201|COMP|45011-4|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C1716169|T201|COMP|45015-5|LNC|Adenosine monophosphate.cyclic^baseline|Adenosine monophosphate.cyclic^baseline
C1716174|T201|COMP|45021-3|LNC|Metanephrine & Normetanephrine|Metanephrine & Normetanephrine
C1716175|T201|COMP|45022-1|LNC|Methadone+Metabolite|Methadone+Metabolite
C1716176|T201|COMP|45023-9|LNC|HLA typing for celiac disease panel|HLA typing for celiac disease panel
C1716177|T201|COMP|45024-7|LNC|HLA typing for narcolepsy panel|HLA typing for narcolepsy panel
C1716178|T201|COMP|45025-4|LNC|HLA-A SBT|HLA-A SBT
C1716179|T201|COMP|45026-2|LNC|HLA-A2 SBT|HLA-A2 SBT
C1716180|T201|COMP|45027-0|LNC|HLA-A2 panel|HLA-A2 panel
C1716181|T201|COMP|45028-8|LNC|HLA-B SBT|HLA-B SBT
C1716182|T201|COMP|45029-6|LNC|HLA-DQB1 SBT|HLA-DQB1 SBT
C1716183|T201|COMP|45030-4|LNC|HLA-DRB1 SBT|HLA-DRB1 SBT
C1716184|T201|COMP|45031-2|LNC|HLA-C SBT|HLA-C SBT
C1716185|T201|COMP|45032-0|LNC|Tyrosine|Tyrosine
C1716187|T201|COMP|45034-6|LNC|Bacteria producing catalase|Bacteria producing catalase
C1716188|T201|COMP|45035-3|LNC|Bacterial virulence|Bacterial virulence
C1716189|T201|COMP|45036-1|LNC|Bacteria producing oxidase|Bacteria producing oxidase
C1716190|T201|COMP|45037-9|LNC|Bacteria producing urease|Bacteria producing urease
C1716191|T201|COMP|45038-7|LNC|Bacteria producing arginine decarboxylase|Bacteria producing arginine decarboxylase
C1716192|T201|COMP|45039-5|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C1716193|T201|COMP|45040-3|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C1716195|T201|COMP|45044-5|LNC|Bacteria producing indole|Bacteria producing indole
C1716196|T201|COMP|45045-2|LNC|Yersinia pestis Ab|Yersinia pestis Ab
C1716197|T201|COMP|45046-0|LNC|Bacteria producing X & V factors|Bacteria producing X & V factors
C1716198|T201|COMP|45047-8|LNC|Cortisol^12 AM specimen|Cortisol^12 AM specimen
C1716199|T201|COMP|45048-6|LNC|Cortisol^12 PM specimen|Cortisol^12 PM specimen
C1716200|T201|COMP|45049-4|LNC|Cortisol^4 PM specimen|Cortisol^4 PM specimen
C1716201|T201|COMP|45050-2|LNC|Cortisol^8 AM specimen|Cortisol^8 AM specimen
C1716202|T201|COMP|45051-0|LNC|Cortisol^8 PM specimen|Cortisol^8 PM specimen
C1716203|T201|COMP|45052-8|LNC|Glucose^12 AM specimen|Glucose^12 AM specimen
C1716204|T201|COMP|45053-6|LNC|Glucose^8 AM specimen|Glucose^8 AM specimen
C1716205|T201|COMP|45054-4|LNC|Glucose^12 PM specimen|Glucose^12 PM specimen
C1716206|T201|COMP|45055-1|LNC|Glucose^4 PM specimen|Glucose^4 PM specimen
C1716214|T201|COMP|46195-4|LNC|Legionella pneumophila 2+3+4+5+6+8 Ab|Legionella pneumophila 2+3+4+5+6+8 Ab
C1716215|T201|COMP|46196-2|LNC|Leptospira interrogans Ab.IgG|Leptospira interrogans Ab.IgG
C1716216|T201|COMP|46197-0|LNC|Measles virus Ab|Measles virus Ab
C1716217|T201|COMP|46198-8|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C1716218|T201|COMP|46199-6|LNC|Parainfluenza virus 1 Ab|Parainfluenza virus 1 Ab
C1716219|T201|COMP|46200-2|LNC|Parainfluenza virus 3 Ab|Parainfluenza virus 3 Ab
C1716220|T201|COMP|46201-0|LNC|Porcine adenovirus Ab|Porcine adenovirus Ab
C1716221|T201|COMP|46202-8|LNC|Psittacid herpesvirus 1 Ab|Psittacid herpesvirus 1 Ab
C1716222|T201|COMP|46203-6|LNC|Reagin Ab|Reagin Ab
C1716223|T201|COMP|45056-9|LNC|Glucose^8 PM specimen|Glucose^8 PM specimen
C1716224|T201|COMP|45057-7|LNC|Cardiolipin Ab.IgA & IgG & IgM panel|Cardiolipin Ab.IgA & IgG & IgM panel
C1716225|T201|COMP|45058-5|LNC|cycloSPORINE.monoclonal & polyclonal panel|cycloSPORINE.monoclonal & polyclonal panel
C1716226|T201|COMP|45061-9|LNC|Spermatozoa Ab.IgA & IgG & IgM panel|Spermatozoa Ab.IgA & IgG & IgM panel
C1716227|T201|COMP|45062-7|LNC|C reactive protein|C reactive protein
C1716228|T201|COMP|45063-5|LNC|Varicella zoster virus Ab.IgG & IgM panel|Varicella zoster virus Ab.IgG & IgM panel
C1716232|T201|COMP|45068-4|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae DNA|Chlamydia trachomatis+Neisseria gonorrhoeae DNA
C1716233|T201|COMP|45069-2|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1716234|T201|COMP|45070-0|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1716235|T201|COMP|45071-8|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1716236|T201|COMP|45072-6|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1716237|T201|COMP|45073-4|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1716238|T201|COMP|45074-2|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1716239|T201|COMP|45075-9|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1716240|T201|COMP|45076-7|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1716241|T201|COMP|45084-1|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1716242|T201|COMP|45085-8|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1716243|T201|COMP|45086-6|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1716244|T201|COMP|45089-0|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1716245|T201|COMP|45090-8|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1716246|T201|COMP|45091-6|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1716247|T201|COMP|45092-4|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1716248|T201|COMP|45093-2|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C1716249|T201|COMP|45094-0|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C1716250|T201|COMP|45095-7|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C1716251|T201|COMP|45096-5|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C1716252|T201|COMP|45097-3|LNC|Chlamydia sp identified|Chlamydia sp identified
C1716253|T201|COMP|45098-1|LNC|Chlamydia sp identified|Chlamydia sp identified
C1716254|T201|COMP|45099-9|LNC|Chlamydia sp identified|Chlamydia sp identified
C1716255|T201|COMP|45100-5|LNC|Chlamydia sp identified|Chlamydia sp identified
C1716256|T201|COMP|45101-3|LNC|Chlamydia sp identified|Chlamydia sp identified
C1716257|T201|COMP|45102-1|LNC|Chlamydia sp identified|Chlamydia sp identified
C1716258|T201|COMP|45103-9|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716259|T201|COMP|45104-7|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716260|T201|COMP|45105-4|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716261|T201|COMP|45106-2|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716262|T201|COMP|45107-0|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716263|T201|COMP|45108-8|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716264|T201|COMP|45109-6|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716265|T201|COMP|45111-2|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716266|T201|COMP|45112-0|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716267|T201|COMP|45113-8|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716268|T201|COMP|45114-6|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716269|T201|COMP|45116-1|LNC|Mycobacterium gordonae rRNA|Mycobacterium gordonae rRNA
C1716270|T201|COMP|45117-9|LNC|Mycobacterium kansasii rRNA|Mycobacterium kansasii rRNA
C1716271|T201|COMP|45118-7|LNC|Vesicular stomatitis Indiana virus Ag|Vesicular stomatitis Indiana virus Ag
C1716272|T201|COMP|45119-5|LNC|Vesicular stomatitis Indiana virus 1 Ab|Vesicular stomatitis Indiana virus 1 Ab
C1716273|T201|COMP|45120-3|LNC|Vesicular stomatitis Indiana virus Ag|Vesicular stomatitis Indiana virus Ag
C1716274|T201|COMP|45122-9|LNC|Cocal virus Ag|Cocal virus Ag
C1716275|T201|COMP|45123-7|LNC|Cocal virus Ab|Cocal virus Ab
C1716276|T201|COMP|45124-5|LNC|Vesicular stomatitis Alagoas virus Ab|Vesicular stomatitis Alagoas virus Ab
C1716277|T201|COMP|45125-2|LNC|Vesicular stomatitis Alagoas virus Ag|Vesicular stomatitis Alagoas virus Ag
C1716278|T201|COMP|45126-0|LNC|Vesicular stomatitis Alagoas virus Ag|Vesicular stomatitis Alagoas virus Ag
C1716279|T201|COMP|45127-8|LNC|Vesicular stomatitis New Jersey virus Ag|Vesicular stomatitis New Jersey virus Ag
C1716280|T201|COMP|45128-6|LNC|Vesicular stomatitis New Jersey virus Ag|Vesicular stomatitis New Jersey virus Ag
C1716282|T201|COMP|45130-2|LNC|Chlamydia trachomatis Ab|Chlamydia trachomatis Ab
C1716283|T201|COMP|45131-0|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716284|T201|COMP|45132-8|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1716285|T201|COMP|45134-4|LNC|Campylobacter jejuni Ab.IgM|Campylobacter jejuni Ab.IgM
C1716286|T201|COMP|45135-1|LNC|Chlamydia trachomatis Ab.IgG|Chlamydia trachomatis Ab.IgG
C1716287|T201|COMP|45136-9|LNC|Endomysium Ab.IgG|Endomysium Ab.IgG
C1716288|T201|COMP|45137-7|LNC|IgA.secretory|IgA.secretory
C1716289|T201|COMP|45138-5|LNC|Listeria monocytogenes O4b Ab.IgG|Listeria monocytogenes O4b Ab.IgG
C1716290|T201|COMP|45139-3|LNC|Listeria monocytogenes O4b Ab.IgM|Listeria monocytogenes O4b Ab.IgM
C1716291|T201|COMP|45140-1|LNC|Phenols|Phenols
C1716292|T201|COMP|45141-9|LNC|Platelet associated Ab|Platelet associated Ab
C1716293|T201|COMP|45143-5|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C1716294|T201|COMP|45144-3|LNC|clomiPRAMINE|clomiPRAMINE
C1716295|T201|COMP|45145-0|LNC|Methdilazine|Methdilazine
C1716296|T201|COMP|45146-8|LNC|Triflupromazine|Triflupromazine
C1716297|T201|COMP|45147-6|LNC|Propiomazine|Propiomazine
C1716298|T201|COMP|45148-4|LNC|OmpC Ab.IgA|OmpC Ab.IgA
C1716299|T201|COMP|45150-0|LNC|Neutrophil Ab|Neutrophil Ab
C1716300|T201|COMP|45151-8|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C1716301|T201|COMP|45152-6|LNC|OJ Ab|OJ Ab
C1716302|T201|COMP|45153-4|LNC|HLA Ab|HLA Ab
C1716303|T201|COMP|45154-2|LNC|Phenylalanine hydroxylase Ab|Phenylalanine hydroxylase Ab
C1716304|T201|COMP|45155-9|LNC|Platelet factor 4 heparin complex induced Ab|Platelet factor 4 heparin complex induced Ab
C1716305|T201|COMP|45156-7|LNC|Rheumatoid factor|Rheumatoid factor
C1716306|T201|COMP|45157-5|LNC|U2 small nuclear ribonucleoprotein Ab.IgG|U2 small nuclear ribonucleoprotein Ab.IgG
C1716307|T201|COMP|45158-3|LNC|Immune complex|Immune complex
C1716308|T201|COMP|45159-1|LNC|Hepatitis B virus & Hepatitis D virus Ab|Hepatitis B virus & Hepatitis D virus Ab
C1716309|T201|COMP|45160-9|LNC|Acremonium sp Ab|Acremonium sp Ab
C1716310|T201|COMP|45161-7|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1716311|T201|COMP|45162-5|LNC|Escherichia coli O157 Ag|Escherichia coli O157 Ag
C1716312|T201|COMP|45163-3|LNC|Alternaria alternata Ab|Alternaria alternata Ab
C1716313|T201|COMP|45164-1|LNC|Asialoganglioside GM2 Ab|Asialoganglioside GM2 Ab
C1716314|T201|COMP|45165-8|LNC|Borrelia burgdorferi Ab.IgA|Borrelia burgdorferi Ab.IgA
C1716315|T201|COMP|45168-2|LNC|Malonate|Malonate
C1716316|T201|COMP|45169-0|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C1716317|T201|COMP|45170-8|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C1716318|T201|COMP|45171-6|LNC|Pancreatic islet cell Ab|Pancreatic islet cell Ab
C1716319|T201|COMP|45172-4|LNC|Purkinje cells Ab|Purkinje cells Ab
C1716320|T201|COMP|45173-2|LNC|Thyrotropin.alpha subunit|Thyrotropin.alpha subunit
C1716321|T201|COMP|45174-0|LNC|Herpes gestationis Ab panel|Herpes gestationis Ab panel
C1716324|T201|COMP|45177-3|LNC|Herpes gestationis Ab.IgG.non-complement fixing|Herpes gestationis Ab.IgG.non-complement fixing
C1716325|T201|COMP|45178-1|LNC|Basement membrane zone Ab.IgG|Basement membrane zone Ab.IgG
C1716326|T201|COMP|45179-9|LNC|Herpes gestationis Ab.IgG.complement fixing|Herpes gestationis Ab.IgG.complement fixing
C1716327|T201|COMP|45180-7|LNC|1p chromosome deletion|1p chromosome deletion
C1716328|T201|COMP|45189-8|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C1716329|T201|COMP|45192-2|LNC|Carnitine esters/Carnitine.free (C0)|Carnitine esters/Carnitine.free (C0)
C1716330|T201|COMP|45193-0|LNC|Cells.CD20+CD52+/100 cells|Cells.CD20+CD52+/100 cells
C1716331|T201|COMP|45194-8|LNC|Choriogonadotropin.intact+Beta subunit|Choriogonadotropin.intact+Beta subunit
C1716332|T201|COMP|45195-5|LNC|Cow epithelium+Cow dander Ab.IgE|Cow epithelium+Cow dander Ab.IgE
C1716333|T201|COMP|45196-3|LNC|Cytokines|Cytokines
C1716334|T201|COMP|45197-1|LNC|Decanoylcarnitine (C10)|Decanoylcarnitine (C10)
C1716335|T201|COMP|45198-9|LNC|Decenoylcarnitine (C10:1)|Decenoylcarnitine (C10:1)
C1716336|T201|COMP|45199-7|LNC|Dodecanoylcarnitine (C12)|Dodecanoylcarnitine (C12)
C1716337|T201|COMP|45200-3|LNC|Dodecenoylcarnitine (C12:1)|Dodecenoylcarnitine (C12:1)
C1716338|T201|COMP|45201-1|LNC|Egg whole Ab.IgG|Egg whole Ab.IgG
C1716339|T201|COMP|45202-9|LNC|Ganglioside GD1a Ab|Ganglioside GD1a Ab
C1716340|T201|COMP|45203-7|LNC|Ganglioside GQ1b Ab|Ganglioside GQ1b Ab
C1716341|T201|COMP|45204-5|LNC|Glucose^3rd specimen post XXX challenge|Glucose^3rd specimen post XXX challenge
C1716342|T201|COMP|45205-2|LNC|Glucose^4th specimen post XXX challenge|Glucose^4th specimen post XXX challenge
C1716343|T201|COMP|45206-0|LNC|Glucose^5th specimen post XXX challenge|Glucose^5th specimen post XXX challenge
C1716344|T201|COMP|45207-8|LNC|Glutarylcarnitine (C5-DC)|Glutarylcarnitine (C5-DC)
C1716345|T201|COMP|45208-6|LNC|Hemoglobin A|Hemoglobin A
C1716346|T201|COMP|45209-4|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C1716347|T201|COMP|45210-2|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C1716348|T201|COMP|45211-0|LNC|Hexanoylcarnitine (C6)|Hexanoylcarnitine (C6)
C1716349|T201|COMP|45212-8|LNC|HIV 2 p31+p34 Ab|HIV 2 p31+p34 Ab
C1716350|T201|COMP|45213-6|LNC|Isobutyrylcarnitine (C4)|Isobutyrylcarnitine (C4)
C1716351|T201|COMP|45214-4|LNC|Isoleucine+Leucine|Isoleucine+Leucine
C1716352|T201|COMP|45216-9|LNC|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)
C1716353|T201|COMP|45217-7|LNC|Linoleoylcarnitine (C18:2)|Linoleoylcarnitine (C18:2)
C1716354|T201|COMP|45218-5|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C1716355|T201|COMP|45219-3|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C1716356|T201|COMP|45220-1|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C1716357|T201|COMP|45221-9|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C1716358|T201|COMP|45222-7|LNC|Methylmalonylcarnitine (C4-DC)|Methylmalonylcarnitine (C4-DC)
C1716359|T201|COMP|45223-5|LNC|Moxifloxacin|Moxifloxacin
C1716360|T201|COMP|45224-3|LNC|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C1716361|T201|COMP|45225-0|LNC|Pancreatic islet cell complement fixing Ab|Pancreatic islet cell complement fixing Ab
C1716362|T201|COMP|45226-8|LNC|Ribosomal P Ab.IgG|Ribosomal P Ab.IgG
C1716363|T201|COMP|45227-6|LNC|Rubus fruticosus Ab.IgE/IgE.total|Rubus fruticosus Ab.IgE/IgE.total
C1716364|T201|COMP|45228-4|LNC|Streptolysin O Ab|Streptolysin O Ab
C1716365|T201|COMP|45229-2|LNC|Toxocara cati Ab|Toxocara cati Ab
C1716398|T201|COMP|45265-6|LNC|Immunodeficiency markers|Immunodeficiency markers
C1716399|T201|COMP|45266-4|LNC|Chronic leukemia markers|Chronic leukemia markers
C1716400|T201|COMP|45268-0|LNC|Immunodeficiency panel|Immunodeficiency panel
C1716401|T201|COMP|45269-8|LNC|Chronic leukemia panel|Chronic leukemia panel
C1716402|T201|COMP|45270-6|LNC|Acute leukemia panel|Acute leukemia panel
C1716403|T201|COMP|45271-4|LNC|Bordetella bronchiseptica DNA|Bordetella bronchiseptica DNA
C1716404|T201|COMP|45272-2|LNC|Sympathomimetics|Sympathomimetics
C1716406|T201|COMP|45274-8|LNC|Low molecular weight heparin induced platelet Ab|Low molecular weight heparin induced platelet Ab
C1716407|T201|COMP|45275-5|LNC|Bacteria identified|Bacteria identified
C1716408|T201|COMP|45276-3|LNC|Bacteria identified|Bacteria identified
C1716409|T201|COMP|45277-1|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C1716410|T201|COMP|45278-9|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C1716411|T201|COMP|45279-7|LNC|Influenza virus A+B Ab|Influenza virus A+B Ab
C1716412|T201|COMP|45280-5|LNC|Echovirus 9 Ab|Echovirus 9 Ab
C1716413|T201|COMP|45281-3|LNC|Echovirus 7 Ab|Echovirus 7 Ab
C1716414|T201|COMP|45282-1|LNC|Echovirus 30 Ab|Echovirus 30 Ab
C1716415|T201|COMP|45284-7|LNC|DPYD gene targeted mutation analysis|DPYD gene targeted mutation analysis
C1716416|T201|COMP|45285-4|LNC|Date and time|Date and time
C1716417|T201|COMP|45286-2|LNC|Cytomegalovirus Ab.IgA|Cytomegalovirus Ab.IgA
C1716418|T201|COMP|45287-0|LNC|Coxsackievirus B6 Ab|Coxsackievirus B6 Ab
C1716419|T201|COMP|45288-8|LNC|Coxsackievirus B5 Ab|Coxsackievirus B5 Ab
C1716420|T201|COMP|45289-6|LNC|Coxsackievirus B4 Ab|Coxsackievirus B4 Ab
C1716421|T201|COMP|45290-4|LNC|Coxsackievirus B3 Ab|Coxsackievirus B3 Ab
C1716422|T201|COMP|45291-2|LNC|Coxsackievirus B2 Ab|Coxsackievirus B2 Ab
C1716423|T201|COMP|45292-0|LNC|Coxsackievirus B1 Ab|Coxsackievirus B1 Ab
C1716424|T201|COMP|45294-6|LNC|Bordetella bronchiseptica DNA|Bordetella bronchiseptica DNA
C1716425|T201|COMP|45296-1|LNC|Cortisol^pre dose dexamethasone|Cortisol^pre dose dexamethasone
C1716426|T201|COMP|45297-9|LNC|Glucose|Glucose
C1716427|T201|COMP|45298-7|LNC|Glucose^2.5H post 50 g lactose PO|Glucose^2.5H post 50 g lactose PO
C1716428|T201|COMP|45299-5|LNC|Glucose^45M post dose lactose PO|Glucose^45M post dose lactose PO
C1716429|T201|COMP|45300-1|LNC|Glycerol|Glycerol
C1716430|T201|COMP|45301-9|LNC|Nortriptyline|Nortriptyline
C1716431|T201|COMP|45302-7|LNC|Urea|Urea
C1716432|T201|COMP|45303-5|LNC|Urea^2H specimen|Urea^2H specimen
C1716433|T201|COMP|45304-3|LNC|Urea^4H specimen|Urea^4H specimen
C1716434|T201|COMP|45305-0|LNC|Coproporphyrin 1|Coproporphyrin 1
C1716435|T201|COMP|45307-6|LNC|Deuteroporphyrin|Deuteroporphyrin
C1716436|T201|COMP|45308-4|LNC|Heptacarboxylate|Heptacarboxylate
C1716437|T201|COMP|45309-2|LNC|Hexacarboxylate|Hexacarboxylate
C1716438|T201|COMP|45310-0|LNC|Mesoporphyrin|Mesoporphyrin
C1716439|T201|COMP|45311-8|LNC|Pentacarboxylate|Pentacarboxylate
C1716440|T201|COMP|45312-6|LNC|Uroporphyrin 3 isomer|Uroporphyrin 3 isomer
C1716441|T201|COMP|45313-4|LNC|Coproporphyrin 1/Creatinine|Coproporphyrin 1/Creatinine
C1716442|T201|COMP|45314-2|LNC|Coproporphyrin 3/Coproporphyrin 1|Coproporphyrin 3/Coproporphyrin 1
C1716443|T201|COMP|45316-7|LNC|Hexacarboxylate/Creatinine|Hexacarboxylate/Creatinine
C1716444|T201|COMP|45317-5|LNC|Pentacarboxylate/Creatinine|Pentacarboxylate/Creatinine
C1716445|T201|COMP|45318-3|LNC|Uroporphyrin 3 isomer/Creatinine|Uroporphyrin 3 isomer/Creatinine
C1716446|T201|COMP|45320-9|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C1716447|T201|COMP|45321-7|LNC|FMR1 gene allele 1.CGG repeats|FMR1 gene allele 1.CGG repeats
C1716448|T201|COMP|45322-5|LNC|FMR1 gene allele 2.CGG repeats|FMR1 gene allele 2.CGG repeats
C1716450|T201|COMP|45324-1|LNC|Ethyl glucuronide|Ethyl glucuronide
C1716451|T201|COMP|45325-8|LNC|Campylobacter jejuni Ab.IgG|Campylobacter jejuni Ab.IgG
C1716452|T201|COMP|45326-6|LNC|Cytomegalovirus Ab.IgG avidity|Cytomegalovirus Ab.IgG avidity
C1716453|T201|COMP|45327-4|LNC|FMR1 gene targeted mutation analysis|FMR1 gene targeted mutation analysis
C1716454|T201|COMP|45328-2|LNC|Glutathione peroxidase|Glutathione peroxidase
C1716455|T201|COMP|45329-0|LNC|Glutathione reductase|Glutathione reductase
C1716456|T201|COMP|45330-8|LNC|Leptospira interrogans Ab.IgG|Leptospira interrogans Ab.IgG
C1716457|T201|COMP|45331-6|LNC|NF1 gene targeted mutation analysis|NF1 gene targeted mutation analysis
C1716458|T201|COMP|45332-4|LNC|NF2 gene targeted mutation analysis|NF2 gene targeted mutation analysis
C1716459|T201|COMP|45334-0|LNC|Tryptase|Tryptase
C1716460|T201|COMP|45335-7|LNC|Bacteria identification test|Bacteria identification test
C1716461|T201|COMP|45336-5|LNC|Bacteria producing hemolysis|Bacteria producing hemolysis
C1716462|T201|COMP|45337-3|LNC|Bacterial biochemical profile|Bacterial biochemical profile
C1716463|T201|COMP|45338-1|LNC|Proinsulin/Insulin|Proinsulin/Insulin
C1716464|T201|COMP|45339-9|LNC|Tick identified^^^4|Tick identified^^^4
C1716465|T201|COMP|45340-7|LNC|Tick identified^^^3|Tick identified^^^3
C1716466|T201|COMP|45341-5|LNC|Tick identified^^^2|Tick identified^^^2
C1716467|T201|COMP|45342-3|LNC|Tick identified|Tick identified
C1716468|T201|COMP|45343-1|LNC|Sex&Stage|Sex&Stage
C1716469|T201|COMP|45344-9|LNC|Mouth intact|Mouth intact
C1716470|T201|COMP|45345-6|LNC|Engorgement|Engorgement
C1716471|T201|COMP|45346-4|LNC|Date tick removed|Date tick removed
C1716472|T201|COMP|45347-2|LNC|Date tick attached|Date tick attached
C1716473|T201|COMP|45348-0|LNC|Date tick acquired|Date tick acquired
C1716474|T201|COMP|45350-6|LNC|Tick identification panel|Tick identification panel
C1716475|T201|COMP|45351-4|LNC|Date of skin test|Date of skin test
C1716476|T201|COMP|45352-2|LNC|Date skin test interpreted|Date skin test interpreted
C1716477|T201|COMP|45353-0|LNC|Date of analysis|Date of analysis
C1716479|T201|COMP|45356-3|LNC|Time Rh immune globulin given|Time Rh immune globulin given
C1716480|T201|COMP|45357-1|LNC|Erythrocytes.filamented|Erythrocytes.filamented
C1716483|T201|COMP|45370-4|LNC|Platelet crossmatch|Platelet crossmatch
C1716486|T201|COMP|45373-8|LNC|Medication route|Medication route
C1716487|T201|COMP|45374-6|LNC|Specimen expiration date|Specimen expiration date
C1716488|T201|COMP|45375-3|LNC|Time of analysis|Time of analysis
C1716489|T201|COMP|45377-9|LNC|Time of transfusion reaction|Time of transfusion reaction
C1716490|T201|COMP|45378-7|LNC|Glutathione peroxidase|Glutathione peroxidase
C1716491|T201|COMP|45379-5|LNC|Eosinophils|Eosinophils
C1716492|T201|COMP|45380-3|LNC|Basophilic stippling.fine|Basophilic stippling.fine
C1716493|T201|COMP|45381-1|LNC|Basophilic stippling.coarse|Basophilic stippling.coarse
C1716494|T201|COMP|45382-9|LNC|Epidermis Ab|Epidermis Ab
C1716495|T201|COMP|45383-7|LNC|Leukocytes|Leukocytes
C1716510|T201|COMP|46080-8|LNC|Erythrocytes.CD55/100 erythrocytes|Erythrocytes.CD55/100 erythrocytes
C1716511|T201|COMP|46081-6|LNC|Theophylline|Theophylline
C1716512|T201|COMP|46082-4|LNC|Influenza virus A Ag|Influenza virus A Ag
C1716513|T201|COMP|46083-2|LNC|Influenza virus B Ag|Influenza virus B Ag
C1716514|T201|COMP|46084-0|LNC|Immunoglobulin light chains|Immunoglobulin light chains
C1716515|T201|COMP|46086-5|LNC|Creatinine^2H specimen|Creatinine^2H specimen
C1716516|T201|COMP|46087-3|LNC|Erythrocytes^2nd tube|Erythrocytes^2nd tube
C1716517|T201|COMP|46088-1|LNC|Leukocytes^2nd tube|Leukocytes^2nd tube
C1716518|T201|COMP|45384-5|LNC|Leucine crystals|Leucine crystals
C1716519|T201|COMP|45385-2|LNC|Hippurate crystals|Hippurate crystals
C1716520|T201|COMP|45386-0|LNC|Epithelial casts|Epithelial casts
C1716521|T201|COMP|45387-8|LNC|Cystine crystals|Cystine crystals
C1716522|T201|COMP|45388-6|LNC|Calcium phosphate crystals|Calcium phosphate crystals
C1716523|T201|COMP|45389-4|LNC|Calcium carbonate crystals|Calcium carbonate crystals
C1716524|T201|COMP|45390-2|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C1716525|T201|COMP|45391-0|LNC|Epithelial cells.renal|Epithelial cells.renal
C1717124|T201|COMP|46089-9|LNC|Leukocytes^3rd tube|Leukocytes^3rd tube
C1717125|T201|COMP|46091-5|LNC|Erythrocytes^3rd tube|Erythrocytes^3rd tube
C1717126|T201|COMP|46092-3|LNC|Erythrocytes^4th tube|Erythrocytes^4th tube
C1717127|T201|COMP|46093-1|LNC|Calcium.ionized|Calcium.ionized
C1717128|T201|COMP|46094-9|LNC|Plasmodium sp Ag|Plasmodium sp Ag
C1717129|T201|COMP|46095-6|LNC|Anabolic steroids|Anabolic steroids
C1717130|T201|COMP|46096-4|LNC|Arsenic|Arsenic
C1717131|T201|COMP|46097-2|LNC|Time corticotropin given|Time corticotropin given
C1717133|T201|COMP|46099-8|LNC|Calcium^^corrected for albumin|Calcium^^corrected for albumin
C1717134|T201|COMP|46100-4|LNC|Pregnenolone^1H post 250 ug corticotropin|Pregnenolone^1H post 250 ug corticotropin
C1717141|T201|COMP|46108-7|LNC|18q chromosome deletion|18q chromosome deletion
C1717142|T201|COMP|46109-5|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C1717143|T201|COMP|46120-2|LNC|Borrelia burgdorferi 41kD Ab.IgG|Borrelia burgdorferi 41kD Ab.IgG
C1717144|T201|COMP|46121-0|LNC|Borrelia burgdorferi 45kD Ab.IgG|Borrelia burgdorferi 45kD Ab.IgG
C1717145|T201|COMP|46122-8|LNC|Borrelia burgdorferi 58kD Ab.IgG|Borrelia burgdorferi 58kD Ab.IgG
C1717146|T201|COMP|46123-6|LNC|Borrelia burgdorferi 66kD Ab.IgG|Borrelia burgdorferi 66kD Ab.IgG
C1717147|T201|COMP|46124-4|LNC|Borrelia burgdorferi 93kD Ab.IgG|Borrelia burgdorferi 93kD Ab.IgG
C1717148|T201|COMP|46126-9|LNC|Endomysium Ab.IgA|Endomysium Ab.IgA
C1717149|T201|COMP|46128-5|LNC|Tissue transglutaminase Ab.IgA|Tissue transglutaminase Ab.IgA
C1717150|T201|COMP|46129-3|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C1717151|T201|COMP|46130-1|LNC|Prealbumin|Prealbumin
C1717152|T201|COMP|46131-9|LNC|Clostridioides difficile toxin B|Clostridioides difficile toxin B
C1717153|T201|COMP|46132-7|LNC|Glycosaminoglycans/Creatinine|Glycosaminoglycans/Creatinine
C1717154|T201|COMP|46133-5|LNC|Epithelial cells|Epithelial cells
C1717155|T201|COMP|46134-3|LNC|Granular casts|Granular casts
C1717156|T201|COMP|46135-0|LNC|Hyaline casts|Hyaline casts
C1717157|T201|COMP|46136-8|LNC|Transitional cells|Transitional cells
C1717158|T201|COMP|46137-6|LNC|Triple phosphate crystals|Triple phosphate crystals
C1717159|T201|COMP|46138-4|LNC|Urate crystals|Urate crystals
C1717174|T201|COMP|46154-1|LNC|Trichomonas vaginalis rRNA|Trichomonas vaginalis rRNA
C1717175|T201|COMP|46156-6|LNC|Ascaris lumbricoides larva Ab.IgG|Ascaris lumbricoides larva Ab.IgG
C1717176|T201|COMP|46157-4|LNC|Aspergillus glaucus Ab|Aspergillus glaucus Ab
C1717177|T201|COMP|46158-2|LNC|Bartonella sp Ab.IgG|Bartonella sp Ab.IgG
C1717178|T201|COMP|46159-0|LNC|Bartonella sp Ab.IgM|Bartonella sp Ab.IgM
C1717179|T201|COMP|46161-6|LNC|Borrelia burgdorferi 18kD Ab.IgG|Borrelia burgdorferi 18kD Ab.IgG
C1717180|T201|COMP|46162-4|LNC|Borrelia burgdorferi 23kD Ab.IgG|Borrelia burgdorferi 23kD Ab.IgG
C1717181|T201|COMP|46163-2|LNC|Borrelia burgdorferi 23kD Ab.IgM|Borrelia burgdorferi 23kD Ab.IgM
C1717182|T201|COMP|46164-0|LNC|Borrelia burgdorferi 28kD Ab.IgG|Borrelia burgdorferi 28kD Ab.IgG
C1717183|T201|COMP|46165-7|LNC|Borrelia burgdorferi 30kD Ab.IgG|Borrelia burgdorferi 30kD Ab.IgG
C1717184|T201|COMP|46166-5|LNC|Borrelia burgdorferi 39kD Ab.IgG|Borrelia burgdorferi 39kD Ab.IgG
C1717185|T201|COMP|46167-3|LNC|Borrelia burgdorferi 39kD Ab.IgM|Borrelia burgdorferi 39kD Ab.IgM
C1717186|T201|COMP|46168-1|LNC|Borrelia burgdorferi 41kD Ab.IgG|Borrelia burgdorferi 41kD Ab.IgG
C1717187|T201|COMP|46169-9|LNC|Borrelia burgdorferi 41kD Ab.IgM|Borrelia burgdorferi 41kD Ab.IgM
C1717188|T201|COMP|46170-7|LNC|Borrelia burgdorferi 45kD Ab.IgG|Borrelia burgdorferi 45kD Ab.IgG
C1717189|T201|COMP|46171-5|LNC|Borrelia burgdorferi 58kD Ab.IgG|Borrelia burgdorferi 58kD Ab.IgG
C1717190|T201|COMP|46172-3|LNC|Borrelia burgdorferi 66kD Ab.IgG|Borrelia burgdorferi 66kD Ab.IgG
C1717191|T201|COMP|46173-1|LNC|Borrelia burgdorferi 93kD Ab.IgG|Borrelia burgdorferi 93kD Ab.IgG
C1717192|T201|COMP|46174-9|LNC|Borrelia burgdorferi Ab.IgA|Borrelia burgdorferi Ab.IgA
C1717193|T201|COMP|46175-6|LNC|Cache valley virus Ab|Cache valley virus Ab
C1717194|T201|COMP|46176-4|LNC|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgA|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgA
C1717195|T201|COMP|46179-8|LNC|Chlamydophila sp Ab|Chlamydophila sp Ab
C1717196|T201|COMP|46180-6|LNC|Classical swine fever virus Ab|Classical swine fever virus Ab
C1717197|T201|COMP|46181-4|LNC|Coccidioides sp Ab.IgA|Coccidioides sp Ab.IgA
C1717198|T201|COMP|46182-2|LNC|Coccidioides sp Ab.IgG|Coccidioides sp Ab.IgG
C1717199|T201|COMP|46183-0|LNC|Coccidioides sp Ab.IgM|Coccidioides sp Ab.IgM
C1717200|T201|COMP|46184-8|LNC|Echinococcus granulosus Ab|Echinococcus granulosus Ab
C1717201|T201|COMP|46185-5|LNC|Ehrlichia risticii Ab|Ehrlichia risticii Ab
C1717202|T201|COMP|46186-3|LNC|Equine herpesvirus 1 Ab|Equine herpesvirus 1 Ab
C1717203|T201|COMP|46187-1|LNC|Equine herpesvirus 2 Ab|Equine herpesvirus 2 Ab
C1717204|T201|COMP|46188-9|LNC|Equine herpesvirus 3 Ab|Equine herpesvirus 3 Ab
C1717205|T201|COMP|46189-7|LNC|Goose parvovirus Ab|Goose parvovirus Ab
C1717206|T201|COMP|46190-5|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C1717207|T201|COMP|46192-1|LNC|HTLV II Ab.IgG|HTLV II Ab.IgG
C1717208|T201|COMP|46193-9|LNC|Infectious bronchitis virus JMK Ab|Infectious bronchitis virus JMK Ab
C1717209|T201|COMP|46194-7|LNC|Legionella non pneumophila sp Ab|Legionella non pneumophila sp Ab
C1717210|T201|COMP|46204-4|LNC|Salmonella typhi O D Ab|Salmonella typhi O D Ab
C1717211|T201|COMP|46205-1|LNC|Streptococcus pneumoniae Ab.IgG|Streptococcus pneumoniae Ab.IgG
C1717212|T201|COMP|46206-9|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1717220|T201|COMP|43269-0|LNC|Ceftobiprole|Ceftobiprole
C1717223|T201|COMP|43176-7|LNC|Lithium|Lithium
C1717225|T201|COMP|43737-6|LNC|Tipranavir|Tipranavir
C1717226|T201|COMP|43826-7|LNC|Androstanolone|Androstanolone
C1717227|T201|COMP|43174-2|LNC|Chlamydia trachomatis L2 Ab.IgA|Chlamydia trachomatis L2 Ab.IgA
C1717229|T201|COMP|43204-7|LNC|Parainfluenza virus 2 Ab|Parainfluenza virus 2 Ab
C1717230|T201|COMP|43217-9|LNC|Cortisol^15M post dose corticotropin IM|Cortisol^15M post dose corticotropin IM
C1717231|T201|COMP|43221-1|LNC|Chloride/Creatinine|Chloride/Creatinine
C1717232|T201|COMP|43232-8|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C1717233|T201|COMP|43239-3|LNC|Norsildenafil|Norsildenafil
C1717234|T201|COMP|43266-6|LNC|Leishmania chagasi K39 Ab|Leishmania chagasi K39 Ab
C1717235|T201|COMP|43296-3|LNC|HTLV I+II gp46 Ab|HTLV I+II gp46 Ab
C1717236|T201|COMP|43319-3|LNC|Avian metapneumovirus A Ab|Avian metapneumovirus A Ab
C1717237|T201|COMP|43320-1|LNC|Avian metapneumovirus B Ab|Avian metapneumovirus B Ab
C1717238|T201|COMP|43333-4|LNC|Equine herpesvirus 2 Ab|Equine herpesvirus 2 Ab
C1717239|T201|COMP|43338-3|LNC|Infectious bronchitis virus JMK Ab|Infectious bronchitis virus JMK Ab
C1717240|T201|COMP|43353-2|LNC|Avian metapneumovirus C Ab|Avian metapneumovirus C Ab
C1717241|T201|COMP|43372-2|LNC|Figure associated with report or note|Figure associated with report or note
C1717242|T201|COMP|43389-6|LNC|Streptococcus sp identified|Streptococcus sp identified
C1717243|T201|COMP|43402-7|LNC|Erythrocyte sedimentation rate|Erythrocyte sedimentation rate
C1717244|T201|COMP|43410-0|LNC|Bacteria identified|Bacteria identified
C1717245|T201|COMP|43418-3|LNC|Stem cell product given|Stem cell product given
C1717250|T201|COMP|43688-1|LNC|16-Alpha hydroxypregnenolone/Creatinine|16-Alpha hydroxypregnenolone/Creatinine
C1717251|T201|COMP|44317-6|LNC|Insulin human Ab|Insulin human Ab
C1717252|T201|COMP|44740-9|LNC|Ganglioside GD1a Ab|Ganglioside GD1a Ab
C1717253|T201|COMP|44743-3|LNC|Disialylganglioside GD1b Ab.IgM|Disialylganglioside GD1b Ab.IgM
C1717256|T201|COMP|44989-2|LNC|Chlamydia trachomatis D+K Ab.IgG|Chlamydia trachomatis D+K Ab.IgG
C1717263|T201|COMP|43591-7|LNC|Prunus persica Ab.IgE/IgE.total|Prunus persica Ab.IgE/IgE.total
C1717264|T201|COMP|43607-1|LNC|Albumin|Albumin
C1717265|T201|COMP|43613-9|LNC|Adenovirus Ag|Adenovirus Ag
C1717266|T201|COMP|43629-5|LNC|8-Hydroxyamoxapine|8-Hydroxyamoxapine
C1717270|T201|COMP|43696-4|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C1717271|T201|COMP|43713-7|LNC|Albumin|Albumin
C1717272|T201|COMP|43719-4|LNC|Acetaminophen+oxyCODONE|Acetaminophen+oxyCODONE
C1717273|T201|COMP|43736-8|LNC|Fosamprenavir|Fosamprenavir
C1717274|T201|COMP|43750-9|LNC|SURF1 gene targeted mutation analysis|SURF1 gene targeted mutation analysis
C1717277|T201|COMP|43798-8|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C1717278|T201|COMP|43799-6|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C1717279|T201|COMP|43815-0|LNC|Arsenic|Arsenic
C1717280|T201|COMP|43816-8|LNC|Amylase|Amylase
C1717281|T201|COMP|43837-4|LNC|Influenza virus A Ab.IgG|Influenza virus A Ab.IgG
C1717282|T201|COMP|43839-0|LNC|Influenza virus B Ab.IgG|Influenza virus B Ab.IgG
C1717283|T201|COMP|43855-6|LNC|Urease^2H post incubation|Urease^2H post incubation
C1717284|T201|COMP|43856-4|LNC|Cells.CD3+CD25+/100 cells|Cells.CD3+CD25+/100 cells
C1717285|T201|COMP|43873-9|LNC|Aspergillus sp Ab.IgM|Aspergillus sp Ab.IgM
C1717286|T201|COMP|43874-7|LNC|Influenza virus A Ag|Influenza virus A Ag
C1717287|T201|COMP|43876-2|LNC|Antimony|Antimony
C1717288|T201|COMP|43892-9|LNC|Borate|Borate
C1717289|T201|COMP|43894-5|LNC|Bismuth|Bismuth
C1717290|T201|COMP|43903-4|LNC|Azinphos-methyl|Azinphos-methyl
C1717291|T201|COMP|43909-1|LNC|Bordetella pertussis Ag|Bordetella pertussis Ag
C1717292|T201|COMP|43932-3|LNC|Rheumatoid factor|Rheumatoid factor
C1717293|T201|COMP|43938-0|LNC|Cells.CD59/100 cells|Cells.CD59/100 cells
C1717294|T201|COMP|43954-7|LNC|Cells.CD4+CD45RO+|Cells.CD4+CD45RO+
C1717295|T201|COMP|43955-4|LNC|Cells.CD4+CD45RO+|Cells.CD4+CD45RO+
C1717296|T201|COMP|43966-1|LNC|Cells.CD4+CD45RA+/100 cells|Cells.CD4+CD45RA+/100 cells
C1717297|T201|COMP|43972-9|LNC|Cells.CD19|Cells.CD19
C1717298|T201|COMP|43990-1|LNC|Clarithromycin 3.0 ug/mL|Clarithromycin 3.0 ug/mL
C1717299|T201|COMP|44007-3|LNC|Erythrocytes.CD55 & CD59|Erythrocytes.CD55 & CD59
C1717300|T201|COMP|44017-2|LNC|Blasts|Blasts
C1717301|T201|COMP|44025-5|LNC|Aspergillus flavus B Ab|Aspergillus flavus B Ab
C1717302|T201|COMP|44027-1|LNC|Aspergillus fumigatus B Ab|Aspergillus fumigatus B Ab
C1717303|T201|COMP|44030-5|LNC|Aspergillus nidulans H Ab|Aspergillus nidulans H Ab
C1717304|T201|COMP|44041-2|LNC|Basophils|Basophils
C1717305|T201|COMP|44050-3|LNC|Glucose phosphate isomerase|Glucose phosphate isomerase
C1717306|T201|COMP|44067-7|LNC|Cells.CD20+FMC7+|Cells.CD20+FMC7+
C1717307|T201|COMP|44074-3|LNC|Arbovirus Ab|Arbovirus Ab
C1717308|T201|COMP|44079-2|LNC|Chlamydia trachomatis Ab.IgA & IgG & IgM|Chlamydia trachomatis Ab.IgA & IgG & IgM
C1717310|T201|COMP|44099-0|LNC|Galactomannan Ag|Galactomannan Ag
C1717325|T201|COMP|44265-7|LNC|Influenza virus A H6 RNA|Influenza virus A H6 RNA
C1717326|T201|COMP|44285-5|LNC|3-Methylcrotonylglycine/Creatinine|3-Methylcrotonylglycine/Creatinine
C1717327|T201|COMP|44305-1|LNC|Chloral hydrate/Creatinine|Chloral hydrate/Creatinine
C1717328|T201|COMP|44307-7|LNC|Citrulline/Creatinine|Citrulline/Creatinine
C1717329|T201|COMP|44337-4|LNC|Metanephrine.free/Creatinine|Metanephrine.free/Creatinine
C1717330|T201|COMP|44353-1|LNC|Porphyrins/Creatinine|Porphyrins/Creatinine
C1717331|T201|COMP|44356-4|LNC|Follitropin/Creatinine|Follitropin/Creatinine
C1717332|T201|COMP|44364-8|LNC|Glutarate/Creatinine|Glutarate/Creatinine
C1717333|T201|COMP|44377-0|LNC|Homocysteine/Creatinine|Homocysteine/Creatinine
C1717334|T201|COMP|44382-0|LNC|Hyaline casts.broad|Hyaline casts.broad
C1717335|T201|COMP|44392-9|LNC|Immune complex|Immune complex
C1717336|T201|COMP|44401-8|LNC|Sarcosine/Creatinine|Sarcosine/Creatinine
C1717337|T201|COMP|44408-3|LNC|Suberate/Creatinine|Suberate/Creatinine
C1717338|T201|COMP|44412-5|LNC|Tetrahydrodeoxycortisol/Creatinine|Tetrahydrodeoxycortisol/Creatinine
C1717339|T201|COMP|44437-2|LNC|Ascaris sp Ab.IgG|Ascaris sp Ab.IgG
C1717340|T201|COMP|44448-9|LNC|Beta 2 glycoprotein 1 Ab.IgG|Beta 2 glycoprotein 1 Ab.IgG
C1717341|T201|COMP|44455-4|LNC|Borrelia burgdorferi Ab^1st specimen|Borrelia burgdorferi Ab^1st specimen
C1717342|T201|COMP|44463-8|LNC|Herpes simplex virus 1|Herpes simplex virus 1
C1717343|T201|COMP|44469-5|LNC|Herpes simplex virus 1 Ab|Herpes simplex virus 1 Ab
C1717344|T201|COMP|44487-7|LNC|Herpes simplex virus 2|Herpes simplex virus 2
C1717345|T201|COMP|44516-3|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1717346|T201|COMP|44521-3|LNC|Herpes virus 6 Ab.IgG|Herpes virus 6 Ab.IgG
C1717347|T201|COMP|44534-6|LNC|HLA Ab|HLA Ab
C1717348|T201|COMP|44537-9|LNC|HTLV I DNA|HTLV I DNA
C1717349|T201|COMP|44554-4|LNC|Hymenopterase Ab.IgE.RAST class|Hymenopterase Ab.IgE.RAST class
C1717350|T201|COMP|44670-8|LNC|Margin involvement|Margin involvement
C1717354|T201|COMP|46119-4|LNC|Borrelia burgdorferi 41kD Ab.IgM|Borrelia burgdorferi 41kD Ab.IgM
C1717355|T201|COMP|44593-2|LNC|IgE|IgE
C1717356|T201|COMP|44595-7|LNC|IgG|IgG
C1717358|T201|COMP|44625-2|LNC|Periprostatic fat invasion|Periprostatic fat invasion
C1717359|T201|COMP|44640-1|LNC|Histologic type|Histologic type
C1717360|T201|COMP|44659-1|LNC|Dominant nodule.additional dimension 2|Dominant nodule.additional dimension 2
C1717361|T201|COMP|44678-1|LNC|Margin(s) involved by invasive carcinoma|Margin(s) involved by invasive carcinoma
C1717362|T201|COMP|44702-9|LNC|Complement C1q Ab|Complement C1q Ab
C1717363|T201|COMP|44718-5|LNC|Lipoprotein.pre-beta/Triglyceride|Lipoprotein.pre-beta/Triglyceride
C1717367|T201|COMP|44800-1|LNC|Burkholderia sp|Burkholderia sp
C1717368|T201|COMP|44803-5|LNC|GNE gene targeted mutation analysis|GNE gene targeted mutation analysis
C1717369|T201|COMP|44822-5|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C1717370|T201|COMP|44839-9|LNC|Choriogonadotropin|Choriogonadotropin
C1717371|T201|COMP|44857-1|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1717372|T201|COMP|44861-3|LNC|4-Hydroxymandelate/Creatinine|4-Hydroxymandelate/Creatinine
C1717373|T201|COMP|44877-9|LNC|Insulin dependent diabetes mellitus|Insulin dependent diabetes mellitus
C1717374|T201|COMP|44892-8|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C1717375|T201|COMP|44914-0|LNC|Beta globulin+Gamma globulin/Protein.total|Beta globulin+Gamma globulin/Protein.total
C1717376|T201|COMP|44925-6|LNC|Prolactin^1H post dose TRH IV|Prolactin^1H post dose TRH IV
C1717377|T201|COMP|44929-8|LNC|Prolactin^15M post dose TRH IV|Prolactin^15M post dose TRH IV
C1717378|T201|COMP|44947-0|LNC|Borrelia burgdorferi 31kD Ab.IgM|Borrelia burgdorferi 31kD Ab.IgM
C1717379|T201|COMP|44948-8|LNC|Borrelia burgdorferi 34kD Ab.IgM|Borrelia burgdorferi 34kD Ab.IgM
C1717380|T201|COMP|45006-4|LNC|Chlamydia trachomatis Ab.IgA|Chlamydia trachomatis Ab.IgA
C1717381|T201|COMP|45012-2|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C1717383|T201|COMP|45041-1|LNC|Francisella tularensis Ag|Francisella tularensis Ag
C1717384|T201|COMP|45042-9|LNC|XXX microorganism Ag|XXX microorganism Ag
C1717386|T201|COMP|45059-3|LNC|Ehrlichia chaffeensis Ab.IgG & IgM panel|Ehrlichia chaffeensis Ab.IgG & IgM panel
C1717387|T201|COMP|45060-1|LNC|Protein & Glucose panel|Protein & Glucose panel
C1717388|T201|COMP|45067-6|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1717389|T201|COMP|45087-4|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1717390|T201|COMP|45088-2|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1717391|T201|COMP|45110-4|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1717392|T201|COMP|45115-3|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1717393|T201|COMP|45121-1|LNC|Cocal virus Ag|Cocal virus Ag
C1717394|T201|COMP|45133-6|LNC|Chlamydia sp Ag|Chlamydia sp Ag
C1717395|T201|COMP|45142-7|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C1717396|T201|COMP|45149-2|LNC|Ej Ab|Ej Ab
C1717397|T201|COMP|45166-6|LNC|Corynebacterium diphtheriae Ab.IgG|Corynebacterium diphtheriae Ab.IgG
C1717398|T201|COMP|45167-4|LNC|IgE|IgE
C1717399|T201|COMP|45190-6|LNC|CASR gene targeted mutation analysis|CASR gene targeted mutation analysis
C1717400|T201|COMP|45215-1|LNC|Isoniazid 2.0 ug/mL|Isoniazid 2.0 ug/mL
C1717404|T201|COMP|45267-2|LNC|Acute leukemia markers|Acute leukemia markers
C1717405|T201|COMP|45283-9|LNC|Echovirus 11 Ab|Echovirus 11 Ab
C1717407|T201|COMP|45295-3|LNC|Acetylcholinesterase/Cholinesterase|Acetylcholinesterase/Cholinesterase
C1717408|T201|COMP|45306-8|LNC|Coproporphyrin 3|Coproporphyrin 3
C1717409|T201|COMP|45315-9|LNC|Coproporphyrin 3/Creatinine|Coproporphyrin 3/Creatinine
C1717410|T201|COMP|45319-1|LNC|Uroporphyrin/Creatinine|Uroporphyrin/Creatinine
C1717411|T201|COMP|45355-5|LNC|Date Rh immune globulin given|Date Rh immune globulin given
C1717414|T201|COMP|45376-1|LNC|Date of transfusion reaction|Date of transfusion reaction
C1717416|T201|COMP|46085-7|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C1717466|T201|COMP|46090-7|LNC|Leukocytes^4th tube|Leukocytes^4th tube
C1717468|T201|COMP|46125-1|LNC|Cardiolipin Ab|Cardiolipin Ab
C1717469|T201|COMP|46127-7|LNC|Haptoglobin|Haptoglobin
C1717471|T201|COMP|46155-8|LNC|Ascaris lumbricoides adult Ab.IgG|Ascaris lumbricoides adult Ab.IgG
C1717472|T201|COMP|46160-8|LNC|Blastomyces dermatitidis Ab.IgG|Blastomyces dermatitidis Ab.IgG
C1717473|T201|COMP|46177-2|LNC|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgG|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgG
C1717474|T201|COMP|46178-0|LNC|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgM|Chlamydia trachomatis D+E+F+G+H+I+J+K Ab.IgM
C1717475|T201|COMP|46191-3|LNC|Histoplasma capsulatum Ab.IgG|Histoplasma capsulatum Ab.IgG
C1718546|T201|COMP|43583-4|LNC|Lipoprotein (little a)|Lipoprotein (little a)
C1718547|T201|COMP|44726-8|LNC|HLA-B51|HLA-B51
C1718548|T201|COMP|45333-2|LNC|Superoxide dismutase|Superoxide dismutase
C1719212|T201|COMP|44419-0|LNC|CIAS1 gene targeted mutation analysis|CIAS1 gene targeted mutation analysis
C1744597|T201|COMP|40491-3|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C1744598|T201|COMP|1197-3|LNC|Little NOS Ab|Little NOS Ab
C1744599|T201|COMP|1198-1|LNC|Little NOS Ab|Little NOS Ab
C1744600|T201|COMP|2758-1|LNC|Phenol|Phenol
C1744633|T201|COMP|24122-4|LNC|Leukocytes|Leukocytes
C1744636|T201|COMP|25441-7|LNC|Homocystine|Homocystine
C1744683|T201|COMP|14832-0|LNC|Metanephrines|Metanephrines
C1744689|T201|COMP|32655-3|LNC|Metanephrines/Creatinine|Metanephrines/Creatinine
C1764750|T201|COMP|21616-8|LNC|APC gene mutation analysis|APC gene mutation analysis
C1764752|T201|COMP|16574-6|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C1764753|T201|COMP|21745-5|LNC|BCL2 gene rearrangements|BCL2 gene rearrangements
C1764754|T201|COMP|13520-2|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C1764755|T201|COMP|40571-2|LNC|Basophils|Basophils
C1764756|T201|COMP|19280-7|LNC|Benzodiazepines tested for|Benzodiazepines tested for
C1764757|T201|COMP|11132-8|LNC|Bilirubin|Bilirubin
C1764758|T201|COMP|6336-2|LNC|Candida albicans Ab|Candida albicans Ab
C1764759|T201|COMP|24473-1|LNC|Cells.CD23/100 cells|Cells.CD23/100 cells
C1764760|T201|COMP|33776-6|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C1764761|T201|COMP|10440-6|LNC|CD30 Ag|CD30 Ag
C1764762|T201|COMP|9560-4|LNC|Lymphocytes.CD5|Lymphocytes.CD5
C1764763|T201|COMP|9562-0|LNC|Lymphocytes.CD5+CD19+|Lymphocytes.CD5+CD19+
C1764764|T201|COMP|24466-5|LNC|Cells.CD56/100 cells|Cells.CD56/100 cells
C1764765|T201|COMP|21177-1|LNC|CFTR gene mutation analysis|CFTR gene mutation analysis
C1764766|T201|COMP|22242-2|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C1764767|T201|COMP|5123-5|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C1764768|T201|COMP|13541-8|LNC|Carbon dioxide|Carbon dioxide
C1764769|T201|COMP|6335-4|LNC|Campylobacter sp identified|Campylobacter sp identified
C1764770|T201|COMP|9841-8|LNC|Casts|Casts
C1764771|T201|COMP|6645-7|LNC|Cefepime|Cefepime
C1764772|T201|COMP|6649-9|LNC|Cefpirome|Cefpirome
C1764773|T201|COMP|6342-0|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C1764774|T201|COMP|12531-0|LNC|Cholesterol|Cholesterol
C1764775|T201|COMP|14440-2|LNC|Cholesterol|Cholesterol
C1764776|T201|COMP|19361-5|LNC|Cocaine|Cocaine
C1764777|T201|COMP|14659-7|LNC|Collection duration|Collection duration
C1764778|T201|COMP|19085-0|LNC|Collection duration|Collection duration
C1764779|T201|COMP|12571-6|LNC|Creatinine|Creatinine
C1764780|T201|COMP|1309-4|LNC|D NOS Ab|D NOS Ab
C1764781|T201|COMP|975-3|LNC|D Ab|D Ab
C1764784|T201|COMP|22262-0|LNC|Eastern equine encephalitis virus Ab|Eastern equine encephalitis virus Ab
C1764785|T201|COMP|13353-8|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C1764786|T201|COMP|40569-6|LNC|Eosinophils|Eosinophils
C1764787|T201|COMP|2244-2|LNC|Estradiol|Estradiol
C1764788|T201|COMP|22311-5|LNC|Helicobacter pylori Ab|Helicobacter pylori Ab
C1764789|T201|COMP|10682-3|LNC|HIV 1 RNA|HIV 1 RNA
C1764790|T201|COMP|4673-0|LNC|HLA-B27|HLA-B27
C1764791|T201|COMP|4675-5|LNC|HLA-B35|HLA-B35
C1764792|T201|COMP|4676-3|LNC|HLA-B35|HLA-B35
C1764793|T201|COMP|6415-5|LNC|Haemophilus influenzae C Ag|Haemophilus influenzae C Ag
C1764794|T201|COMP|20834-8|LNC|Herbicide|Herbicide
C1764795|T201|COMP|27940-6|LNC|Insulin^1.5H post 75 g glucose PO|Insulin^1.5H post 75 g glucose PO
C1764796|T201|COMP|22374-3|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C1764797|T201|COMP|22376-8|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C1764798|T201|COMP|20494-1|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C1764799|T201|COMP|6491-5|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1764800|T201|COMP|23317-1|LNC|Nairobi sheep disease virus Ab|Nairobi sheep disease virus Ab
C1764801|T201|COMP|752-6|LNC|Neutrophils|Neutrophils
C1764802|T201|COMP|13352-0|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C1764803|T201|COMP|40566-2|LNC|Neutrophils|Neutrophils
C1764804|T201|COMP|23348-6|LNC|Pasteurella multocida serotype|Pasteurella multocida serotype
C1764805|T201|COMP|13543-4|LNC|Phosphate|Phosphate
C1764806|T201|COMP|5907-1|LNC|Platelets|Platelets
C1764807|T201|COMP|6530-0|LNC|Rabies virus Ag|Rabies virus Ag
C1764807|T201|COMP|6531-8|LNC|Rabies virus Ag|Rabies virus Ag
C1764808|T201|COMP|6534-2|LNC|Rabies virus Ag|Rabies virus Ag
C1764808|T201|COMP|6535-9|LNC|Rabies virus Ag|Rabies virus Ag
C1764809|T201|COMP|6537-5|LNC|Rabies virus identified|Rabies virus identified
C1764809|T201|COMP|6538-3|LNC|Rabies virus identified|Rabies virus identified
C1764810|T201|COMP|6540-9|LNC|Rabies virus identified|Rabies virus identified
C1764810|T201|COMP|6541-7|LNC|Rabies virus identified|Rabies virus identified
C1764811|T201|COMP|20954-4|LNC|Salmonella sp identified|Salmonella sp identified
C1764812|T201|COMP|19770-7|LNC|Specimen source|Specimen source
C1764813|T201|COMP|10595-7|LNC|Spermatozoa|Spermatozoa
C1764814|T201|COMP|12279-6|LNC|Spermatozoa Ab|Spermatozoa Ab
C1764815|T201|COMP|13628-3|LNC|Spermatozoa.motile/100 spermatozoa|Spermatozoa.motile/100 spermatozoa
C1764816|T201|COMP|23457-5|LNC|Taylorella equigenitalis Ag|Taylorella equigenitalis Ag
C1764818|T201|COMP|12980-9|LNC|Urate|Urate
C1764819|T201|COMP|22612-6|LNC|Western equine encephalitis virus Ab|Western equine encephalitis virus Ab
C1764820|T201|COMP|6520-1|LNC|Pneumocystis carinii Ag|Pneumocystis carinii Ag
C1764821|T201|COMP|21811-5|LNC|t(15,17) (PML,RARA) gene translocation|t(15,17) (PML,RARA) gene translocation
C1764826|T201|COMP|23902-0|LNC|Monocyte+Macrophage/100 leukocytes|Monocyte+Macrophage/100 leukocytes
C1765327|T201|COMP|21019-5|LNC|Metanephrine|Metanephrine
C1765328|T201|COMP|2608-8|LNC|Metanephrines|Metanephrines
C1765329|T201|COMP|19297-1|LNC|Opiates tested for|Opiates tested for
C1765333|T201|COMP|14638-1|LNC|Calculus analysis|Calculus analysis
C1765334|T201|COMP|3427-2|LNC|Cannabinoids|Cannabinoids
C1830044|T201|COMP|47198-7|LNC|Vasopressin^1st specimen post XXX challenge|Vasopressin^1st specimen post XXX challenge
C1830045|T201|COMP|47199-5|LNC|Methionine|Methionine
C1830046|T201|COMP|47200-1|LNC|Methionine+Homocysteine|Methionine+Homocysteine
C1830047|T201|COMP|47201-9|LNC|Bentiromide|Bentiromide
C1830048|T201|COMP|47202-7|LNC|Sincalide|Sincalide
C1830049|T201|COMP|47203-5|LNC|Pyridoxine|Pyridoxine
C1830050|T201|COMP|47204-3|LNC|glipiZIDE|glipiZIDE
C1830051|T201|COMP|47205-0|LNC|metyraPONE|metyraPONE
C1830052|T201|COMP|47206-8|LNC|Corticotropin|Corticotropin
C1830053|T201|COMP|47207-6|LNC|Secretin|Secretin
C1830054|T201|COMP|47208-4|LNC|Arginine|Arginine
C1830055|T201|COMP|47209-2|LNC|Glucagon|Glucagon
C1830056|T201|COMP|47210-0|LNC|Triglyceride^post CFst|Triglyceride^post CFst
C1830057|T201|COMP|47211-8|LNC|Chlamydia trachomatis L2 DNA|Chlamydia trachomatis L2 DNA
C1830058|T201|COMP|47212-6|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1830059|T201|COMP|47213-4|LNC|Cholesterol.in LDL real size pattern|Cholesterol.in LDL real size pattern
C1830060|T201|COMP|47214-2|LNC|Homeostasis model assessment|Homeostasis model assessment
C1830061|T201|COMP|47215-9|LNC|Lipoprotein.beta.subparticle.intermediate|Lipoprotein.beta.subparticle.intermediate
C1830062|T201|COMP|47216-7|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1830063|T201|COMP|47217-5|LNC|Immune complex.C3d|Immune complex.C3d
C1830064|T201|COMP|47218-3|LNC|Cholesterol.in VLDL 3+4|Cholesterol.in VLDL 3+4
C1830065|T201|COMP|47219-1|LNC|Cholesterol.in VLDL 5+6|Cholesterol.in VLDL 5+6
C1830066|T201|COMP|47220-9|LNC|Cholesterol.in HDL 4+5|Cholesterol.in HDL 4+5
C1830067|T201|COMP|47221-7|LNC|Cholesterol.in HDL 1+2|Cholesterol.in HDL 1+2
C1830068|T201|COMP|47365-2|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C1830077|T201|COMP|47383-5|LNC|Nuclear Ab|Nuclear Ab
C1830078|T201|COMP|47384-3|LNC|Cephalosporine mold Ab.IgE.RAST class|Cephalosporine mold Ab.IgE.RAST class
C1830080|T201|COMP|47385-0|LNC|Netilmicin|Netilmicin
C1830095|T201|COMP|46265-5|LNC|Cryofibrinogen|Cryofibrinogen
C1830096|T201|COMP|46266-3|LNC|Myeloperoxidase Ab|Myeloperoxidase Ab
C1830097|T201|COMP|46267-1|LNC|Proteinase 3 Ab|Proteinase 3 Ab
C1830098|T201|COMP|46268-9|LNC|ABO & Rh group^post transfusion reaction|ABO & Rh group^post transfusion reaction
C1830099|T201|COMP|46269-7|LNC|25-Hydroxycalciferol|25-Hydroxycalciferol
C1830100|T201|COMP|46270-5|LNC|ABO group^post transfusion reaction|ABO group^post transfusion reaction
C1830102|T201|COMP|46272-1|LNC|Appearance^post transfusion reaction|Appearance^post transfusion reaction
C1830103|T201|COMP|46425-5|LNC|Lipemic index|Lipemic index
C1830104|T201|COMP|46426-3|LNC|Icteric index|Icteric index
C1830105|T201|COMP|46427-1|LNC|Beta fructofuranosidase|Beta fructofuranosidase
C1830106|T201|COMP|46428-9|LNC|Xylose^15M post 25 g xylose PO|Xylose^15M post 25 g xylose PO
C1830107|T201|COMP|46429-7|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C1830108|T201|COMP|46430-5|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C1830109|T201|COMP|46431-3|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C1830110|T201|COMP|47168-0|LNC|Norepinephrine^4th specimen post XXX challenge|Norepinephrine^4th specimen post XXX challenge
C1830111|T201|COMP|47169-8|LNC|Norepinephrine^5th specimen post XXX challenge|Norepinephrine^5th specimen post XXX challenge
C1830112|T201|COMP|47170-6|LNC|Norepinephrine^5th specimen post XXX challenge|Norepinephrine^5th specimen post XXX challenge
C1830113|T201|COMP|47171-4|LNC|Norepinephrine^6th specimen post XXX challenge|Norepinephrine^6th specimen post XXX challenge
C1830114|T201|COMP|47172-2|LNC|Norepinephrine^6th specimen post XXX challenge|Norepinephrine^6th specimen post XXX challenge
C1830115|T201|COMP|47173-0|LNC|Catecholamines^7th specimen post XXX challenge|Catecholamines^7th specimen post XXX challenge
C1830116|T201|COMP|47174-8|LNC|Norepinephrine^7th specimen post XXX challenge|Norepinephrine^7th specimen post XXX challenge
C1830119|T201|COMP|46218-4|LNC|5-Fluorocytosine|5-Fluorocytosine
C1830120|T201|COMP|46219-2|LNC|Creatinine^4H specimen|Creatinine^4H specimen
C1830121|T201|COMP|46220-0|LNC|Creatinine^overnight|Creatinine^overnight
C1830122|T201|COMP|46221-8|LNC|Glucose^2H specimen|Glucose^2H specimen
C1830123|T201|COMP|46222-6|LNC|Glucose^4H specimen|Glucose^4H specimen
C1830124|T201|COMP|46223-4|LNC|Glucose^overnight|Glucose^overnight
C1830126|T201|COMP|46225-9|LNC|ABCA3 gene targeted mutation analysis|ABCA3 gene targeted mutation analysis
C1830128|T201|COMP|46226-7|LNC|SGCA gene targeted mutation analysis|SGCA gene targeted mutation analysis
C1830130|T201|COMP|46227-5|LNC|DULoxetine|DULoxetine
C1830131|T201|COMP|46228-3|LNC|Clenbuterol|Clenbuterol
C1830132|T201|COMP|46229-1|LNC|Furazabol|Furazabol
C1830133|T201|COMP|46230-9|LNC|Methanolone|Methanolone
C1830134|T201|COMP|46231-7|LNC|Cells.ZAP70/100 cells|Cells.ZAP70/100 cells
C1830136|T201|COMP|46232-5|LNC|Cells.ZAP70/100 cells|Cells.ZAP70/100 cells
C1830137|T201|COMP|46233-3|LNC|Cells.ZAP70/100 cells|Cells.ZAP70/100 cells
C1830138|T201|COMP|46234-1|LNC|Cells.ZAP70/100 cells|Cells.ZAP70/100 cells
C1830139|T201|COMP|46235-8|LNC|Cells.ZAP70/100 cells|Cells.ZAP70/100 cells
C1830140|T201|COMP|46236-6|LNC|HLA-B*51|HLA-B*51
C1830141|T201|COMP|46237-4|LNC|Lymphocytes.kappa/100 lymphocytes|Lymphocytes.kappa/100 lymphocytes
C1830142|T201|COMP|46238-2|LNC|Lymphocytes.kappa/100 lymphocytes|Lymphocytes.kappa/100 lymphocytes
C1830149|T201|COMP|46243-2|LNC|Urea^overnight|Urea^overnight
C1830154|T201|COMP|46248-1|LNC|Borrelia burgdorferi Ab.IgG & IgM|Borrelia burgdorferi Ab.IgG & IgM
C1830160|T201|COMP|46252-3|LNC|Acylcarnitine pattern|Acylcarnitine pattern
C1830162|T201|COMP|46254-9|LNC|Bordetella pertussis.pertussis toxin Ab.IgG|Bordetella pertussis.pertussis toxin Ab.IgG
C1830163|T201|COMP|46255-6|LNC|Methyl ethyl ketone|Methyl ethyl ketone
C1830164|T201|COMP|46256-4|LNC|oxyCODONE.free|oxyCODONE.free
C1830165|T201|COMP|46257-2|LNC|Dihydrocodeine+Hydrocodol|Dihydrocodeine+Hydrocodol
C1830166|T201|COMP|46258-0|LNC|oxyMORphone.free|oxyMORphone.free
C1830167|T201|COMP|46259-8|LNC|Morphine.free|Morphine.free
C1830168|T201|COMP|46260-6|LNC|HYDROmorphone.free|HYDROmorphone.free
C1830169|T201|COMP|46261-4|LNC|HYDROcodone.free|HYDROcodone.free
C1830170|T201|COMP|46262-2|LNC|Codeine.free|Codeine.free
C1830171|T201|COMP|46263-0|LNC|6-Monoacetylmorphine.free|6-Monoacetylmorphine.free
C1830174|T201|COMP|46273-9|LNC|Appearance^post transfusion reaction|Appearance^post transfusion reaction
C1830176|T201|COMP|46275-4|LNC|Major crossmatch^post transfusion reaction|Major crossmatch^post transfusion reaction
C1830177|T201|COMP|46276-2|LNC|Rh^post transfusion reaction|Rh^post transfusion reaction
C1830178|T201|COMP|46277-0|LNC|Rh immune globulin given by|Rh immune globulin given by
C1830286|T201|COMP|46397-6|LNC|Cortisol^15M post 1 ug/kg CRH IV|Cortisol^15M post 1 ug/kg CRH IV
C1830287|T201|COMP|46398-4|LNC|Cortisol^1.5H post 1 ug/kg CRH IV|Cortisol^1.5H post 1 ug/kg CRH IV
C1830288|T201|COMP|46399-2|LNC|Cortisol^2H post 1 ug/kg CRH IV|Cortisol^2H post 1 ug/kg CRH IV
C1830289|T201|COMP|46400-8|LNC|Corticotropin^15M post 1 ug/kg CRH IV|Corticotropin^15M post 1 ug/kg CRH IV
C1830290|T201|COMP|46401-6|LNC|Corticotropin^1.5H post 1 ug/kg CRH IV|Corticotropin^1.5H post 1 ug/kg CRH IV
C1830291|T201|COMP|46402-4|LNC|Corticotropin^2H post 1 ug/kg CRH IV|Corticotropin^2H post 1 ug/kg CRH IV
C1830292|T201|COMP|46403-2|LNC|Cortisol^2H post dose insulin IV|Cortisol^2H post dose insulin IV
C1830293|T201|COMP|46404-0|LNC|Somatotropin^2H post dose insulin IV|Somatotropin^2H post dose insulin IV
C1830294|T201|COMP|46405-7|LNC|Somatotropin^30M pre 1 g/kg glucose PO|Somatotropin^30M pre 1 g/kg glucose PO
C1830295|T201|COMP|46406-5|LNC|Somatotropin^30M post 1 g/kg glucose PO|Somatotropin^30M post 1 g/kg glucose PO
C1830296|T201|COMP|46407-3|LNC|Somatotropin^1.5H post 1 g/kg glucose PO|Somatotropin^1.5H post 1 g/kg glucose PO
C1830297|T201|COMP|46408-1|LNC|Somatotropin^15M pre dose arginine|Somatotropin^15M pre dose arginine
C1830298|T201|COMP|46409-9|LNC|Somatotropin^15M post dose arginine|Somatotropin^15M post dose arginine
C1830299|T201|COMP|46410-7|LNC|Somatotropin^30M post dose arginine|Somatotropin^30M post dose arginine
C1830300|T201|COMP|46411-5|LNC|Somatotropin^45M post dose arginine|Somatotropin^45M post dose arginine
C1830301|T201|COMP|46412-3|LNC|Somatotropin^105M post dose arginine|Somatotropin^105M post dose arginine
C1830302|T201|COMP|46413-1|LNC|Calcitonin^7M post 0.5 ug/kg pentagastrin IV|Calcitonin^7M post 0.5 ug/kg pentagastrin IV
C1830306|T201|COMP|46417-2|LNC|Coagulation tissue factor induced|Coagulation tissue factor induced
C1830307|T201|COMP|46418-0|LNC|Coagulation tissue factor induced.INR|Coagulation tissue factor induced.INR
C1830308|T201|COMP|46419-8|LNC|Erythrocytes|Erythrocytes
C1830309|T201|COMP|46420-6|LNC|Leukocyte clumps|Leukocyte clumps
C1830310|T201|COMP|46421-4|LNC|Mucus|Mucus
C1830311|T201|COMP|46422-2|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C1830312|T201|COMP|46423-0|LNC|Hemoglobin distribution width|Hemoglobin distribution width
C1830313|T201|COMP|46424-8|LNC|Hemolysis index|Hemolysis index
C1830314|T201|COMP|46432-1|LNC|Hydrogen/Expired gas^post 50 g lactose PO|Hydrogen/Expired gas^post 50 g lactose PO
C1830315|T201|COMP|46433-9|LNC|Hydrogen/Expired gas^post 10 g lactulose PO|Hydrogen/Expired gas^post 10 g lactulose PO
C1830318|T201|COMP|46436-2|LNC|Histamine|Histamine
C1830352|T201|COMP|46454-5|LNC|Shigella sp|Shigella sp
C1830353|T201|COMP|46455-2|LNC|Shigella sp DNA|Shigella sp DNA
C1830493|T201|COMP|29626-9|LNC|3-Hydroxysebacate|3-Hydroxysebacate
C1830772|T201|COMP|46698-7|LNC|Cyanide|Cyanide
C1830773|T201|COMP|46699-5|LNC|Fibroblast growth factor 23|Fibroblast growth factor 23
C1830774|T201|COMP|46700-1|LNC|7-Dehydrocholesterol|7-Dehydrocholesterol
C1830775|T201|COMP|46701-9|LNC|Adenosine triphosphate|Adenosine triphosphate
C1830776|T201|COMP|46702-7|LNC|Leukocytes|Leukocytes
C1830777|T201|COMP|46703-5|LNC|Dihydrocodeine.free+Hydrocodol.free|Dihydrocodeine.free+Hydrocodol.free
C1830778|T201|COMP|46704-3|LNC|Dihydrocodeine.free+Hydrocodol.free|Dihydrocodeine.free+Hydrocodol.free
C1830779|T201|COMP|46705-0|LNC|Clostridium botulinum toxin gene|Clostridium botulinum toxin gene
C1830780|T201|COMP|46706-8|LNC|Clostridium perfringens toxin gene|Clostridium perfringens toxin gene
C1830784|T201|COMP|46710-0|LNC|(Beef+Chicken meat+Pork+Turkey meat) Ab.IgE|(Beef+Chicken meat+Pork+Turkey meat) Ab.IgE
C1830789|T201|COMP|46715-9|LNC|B cell crossmatch|B cell crossmatch
C1830790|T201|COMP|46716-7|LNC|Ceruloplasmin|Ceruloplasmin
C1830792|T201|COMP|46718-3|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C1830793|T201|COMP|46719-1|LNC|Streptomycin 4.0 ug/mL|Streptomycin 4.0 ug/mL
C1830795|T201|COMP|46720-9|LNC|T cell crossmatch|T cell crossmatch
C1830796|T201|COMP|46721-7|LNC|Ustilago nuda Ab.IgE|Ustilago nuda Ab.IgE
C1830798|T201|COMP|46722-5|LNC|Cells.ZAP70|Cells.ZAP70
C1830799|T201|COMP|46723-3|LNC|Alpha-1-Microglobulin|Alpha-1-Microglobulin
C1830800|T201|COMP|46724-1|LNC|CYP2C9 gene targeted mutation analysis|CYP2C9 gene targeted mutation analysis
C1830802|T201|COMP|46725-8|LNC|Tropheryma whippelii DNA|Tropheryma whippelii DNA
C1830803|T201|COMP|46726-6|LNC|HTR2A gene+HTR2C gene targeted mutation analysis|HTR2A gene+HTR2C gene targeted mutation analysis
C1830805|T201|COMP|46727-4|LNC|Prolactin.monomeric|Prolactin.monomeric
C1830806|T201|COMP|46728-2|LNC|Weight|Weight
C1830807|T201|COMP|46729-0|LNC|Weight container+Specimen|Weight container+Specimen
C1830808|T201|COMP|46730-8|LNC|Bacterial vaginosis whiff test|Bacterial vaginosis whiff test
C1830809|T201|COMP|46731-6|LNC|RHC gene targeted mutation analysis|RHC gene targeted mutation analysis
C1830810|T201|COMP|46732-4|LNC|Francisella tularensis subtype|Francisella tularensis subtype
C1830811|T201|COMP|46733-2|LNC|Amino acidemias|Amino acidemias
C1830812|T201|COMP|46734-0|LNC|Citrullinemias &or arginosuccinic aciduria|Citrullinemias &or arginosuccinic aciduria
C1830813|T201|COMP|46735-7|LNC|Endocrine disorders|Endocrine disorders
C1830814|T201|COMP|46736-5|LNC|Fatty acid oxidation defects|Fatty acid oxidation defects
C1830815|T201|COMP|46737-3|LNC|Galactosemias|Galactosemias
C1830816|T201|COMP|46738-1|LNC|Genetic disorders|Genetic disorders
C1830817|T201|COMP|46739-9|LNC|Glutaric acidemia type 1|Glutaric acidemia type 1
C1830818|T201|COMP|46740-7|LNC|Hemoglobin disorders|Hemoglobin disorders
C1830819|T201|COMP|46741-5|LNC|Homocystinuria &or other hypermethioninemias|Homocystinuria &or other hypermethioninemias
C1830820|T201|COMP|46742-3|LNC|Isovaleric acidemia &or 2-Methylbutyric acidemia|Isovaleric acidemia &or 2-Methylbutyric acidemia
C1830821|T201|COMP|46743-1|LNC|Maple syrup urine disease|Maple syrup urine disease
C1830822|T201|COMP|46744-9|LNC|Organic acidemias|Organic acidemias
C1830823|T201|COMP|46745-6|LNC|Other amino acidopathies|Other amino acidopathies
C1830825|T201|COMP|46747-2|LNC|Propionic &or methylmalonic acidemias|Propionic &or methylmalonic acidemias
C1830826|T201|COMP|46748-0|LNC|Tyrosinemias|Tyrosinemias
C1830829|T201|COMP|46751-4|LNC|Other organic acidemias|Other organic acidemias
C1830833|T201|COMP|46755-5|LNC|Carnitine uptake defect &or CPT1 deficiency|Carnitine uptake defect &or CPT1 deficiency
C1830834|T201|COMP|46756-3|LNC|Other fatty acid oxidation disorders|Other fatty acid oxidation disorders
C1830835|T201|COMP|46757-1|LNC|Congenital hypothyroidism|Congenital hypothyroidism
C1830836|T201|COMP|46758-9|LNC|Congenital adrenal hyperplasia|Congenital adrenal hyperplasia
C1830837|T201|COMP|46759-7|LNC|Hb SS, Hb SC, Hb SB thal|Hb SS, Hb SC, Hb SB thal
C1830838|T201|COMP|46760-5|LNC|Other hemoglobinopathies|Other hemoglobinopathies
C1830839|T201|COMP|46761-3|LNC|Biotinidase deficiency|Biotinidase deficiency
C1830840|T201|COMP|46762-1|LNC|Congenital hypothyroidism|Congenital hypothyroidism
C1830841|T201|COMP|46763-9|LNC|Secondary congenital hypothyroidism|Secondary congenital hypothyroidism
C1830842|T201|COMP|46764-7|LNC|Thyroid binding globulin deficiency|Thyroid binding globulin deficiency
C1830843|T201|COMP|46765-4|LNC|Sickle cell anemia|Sickle cell anemia
C1830844|T201|COMP|46766-2|LNC|Hemoglobin SC disease|Hemoglobin SC disease
C1830845|T201|COMP|46767-0|LNC|Hemoglobin S beta thalassemia|Hemoglobin S beta thalassemia
C1830846|T201|COMP|46768-8|LNC|Sickle cell carrier (trait)|Sickle cell carrier (trait)
C1830847|T201|COMP|46769-6|LNC|Cystic fibrosis|Cystic fibrosis
C1830848|T201|COMP|46770-4|LNC|Hearing loss|Hearing loss
C1830849|T201|COMP|46771-2|LNC|Classical galactosemia|Classical galactosemia
C1830850|T201|COMP|46772-0|LNC|Galactokinase deficiency|Galactokinase deficiency
C1830851|T201|COMP|46773-8|LNC|Galactose epimerase deficiency|Galactose epimerase deficiency
C1830852|T201|COMP|46774-6|LNC|Carnitine uptake deficiency|Carnitine uptake deficiency
C1830853|T201|COMP|46775-3|LNC|Carnitine palmitoyltransferase 1 deficiency|Carnitine palmitoyltransferase 1 deficiency
C1830854|T201|COMP|46776-1|LNC|CPT2 &or CACT|CPT2 &or CACT
C1830856|T201|COMP|46778-7|LNC|MCAD|MCAD
C1830859|T201|COMP|46781-1|LNC|Malonic acidemia|Malonic acidemia
C1830860|T201|COMP|46782-9|LNC|Argininemia|Argininemia
C1831023|T201|COMP|46945-2|LNC|Beclomethasone dipropionate|Beclomethasone dipropionate
C1831024|T201|COMP|46946-0|LNC|Betamethasone|Betamethasone
C1831025|T201|COMP|46947-8|LNC|Budesonide|Budesonide
C1831026|T201|COMP|46948-6|LNC|Dexamethasone|Dexamethasone
C1831027|T201|COMP|46949-4|LNC|Fludrocortisone|Fludrocortisone
C1831028|T201|COMP|46950-2|LNC|Flunisolide|Flunisolide
C1831029|T201|COMP|46951-0|LNC|Fluorometholone|Fluorometholone
C1831030|T201|COMP|46952-8|LNC|Fluticasone propionate|Fluticasone propionate
C1831031|T201|COMP|46953-6|LNC|Megestrol acetate|Megestrol acetate
C1831032|T201|COMP|46954-4|LNC|Methylprednisolone|Methylprednisolone
C1831033|T201|COMP|46955-1|LNC|prednisoLONE|prednisoLONE
C1831034|T201|COMP|46956-9|LNC|predniSONE|predniSONE
C1831035|T201|COMP|46957-7|LNC|Triamcinolone|Triamcinolone
C1831036|T201|COMP|46958-5|LNC|Triamcinolone acetonide|Triamcinolone acetonide
C1831037|T201|COMP|46959-3|LNC|Synthetic glucocorticoid panel|Synthetic glucocorticoid panel
C1831038|T201|COMP|46960-1|LNC|TCR alpha beta Ag|TCR alpha beta Ag
C1831039|T201|COMP|46961-9|LNC|TCR gamma delta Ag|TCR gamma delta Ag
C1831040|T201|COMP|46962-7|LNC|Vasoactive intestinal peptide Ag|Vasoactive intestinal peptide Ag
C1831042|T201|COMP|46963-5|LNC|Tube number|Tube number
C1831043|T201|COMP|46964-3|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C1831044|T201|COMP|46965-0|LNC|MCOLN1 gene targeted mutation analysis|MCOLN1 gene targeted mutation analysis
C1831045|T201|COMP|46966-8|LNC|Cells.CD69|Cells.CD69
C1831046|T201|COMP|46967-6|LNC|Cells.CD40|Cells.CD40
C1831047|T201|COMP|46968-4|LNC|Cells.CD122|Cells.CD122
C1831048|T201|COMP|46969-2|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C1831049|T201|COMP|46970-0|LNC|BK virus DNA|BK virus DNA
C1831050|T201|COMP|46971-8|LNC|HYDROmorphone.free|HYDROmorphone.free
C1831051|T201|COMP|46973-4|LNC|oxyCODONE.free|oxyCODONE.free
C1831052|T201|COMP|46974-2|LNC|oxyMORphone.free|oxyMORphone.free
C1831053|T201|COMP|46975-9|LNC|oxyMORphone.free|oxyMORphone.free
C1831054|T201|COMP|46976-7|LNC|Benzodiazepines|Benzodiazepines
C1831055|T201|COMP|46977-5|LNC|Benzodiazepines|Benzodiazepines
C1831056|T201|COMP|46978-3|LNC|Salicylates|Salicylates
C1831057|T201|COMP|46979-1|LNC|Flurazepam|Flurazepam
C1831058|T201|COMP|46980-9|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C1831059|T201|COMP|46981-7|LNC|Silicon|Silicon
C1831061|T201|COMP|47310-8|LNC|Haemophilus influenzae B Ab.IgG^1st specimen|Haemophilus influenzae B Ab.IgG^1st specimen
C1831062|T201|COMP|47311-6|LNC|Haemophilus influenzae B Ab.IgG^2nd specimen|Haemophilus influenzae B Ab.IgG^2nd specimen
C1831063|T201|COMP|47312-4|LNC|Influenza virus A Ab.IgM|Influenza virus A Ab.IgM
C1831064|T201|COMP|47313-2|LNC|Influenza virus A Ab.IgG|Influenza virus A Ab.IgG
C1831065|T201|COMP|47314-0|LNC|Influenza virus B Ab.IgG|Influenza virus B Ab.IgG
C1831066|T201|COMP|47315-7|LNC|Influenza virus B Ab.IgM|Influenza virus B Ab.IgM
C1831067|T201|COMP|47369-4|LNC|Calcitonin|Calcitonin
C1831076|T201|COMP|46982-5|LNC|Liver kidney microsomal Ab.IgG|Liver kidney microsomal Ab.IgG
C1831078|T201|COMP|46983-3|LNC|Ethanol|Ethanol
C1831079|T201|COMP|46984-1|LNC|LDL 2|LDL 2
C1831080|T201|COMP|46985-8|LNC|LDL 3|LDL 3
C1831081|T201|COMP|46986-6|LNC|Cholesterol.in VLDL 3|Cholesterol.in VLDL 3
C1831082|T201|COMP|46987-4|LNC|Helicobacter pylori Ab.IgM|Helicobacter pylori Ab.IgM
C1831083|T201|COMP|46988-2|LNC|GBA gene mutations tested for|GBA gene mutations tested for
C1831085|T201|COMP|46989-0|LNC|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C1831086|T201|COMP|46990-8|LNC|ASPA gene targeted mutation analysis|ASPA gene targeted mutation analysis
C1831087|T201|COMP|46991-6|LNC|BLM gene targeted mutation analysis|BLM gene targeted mutation analysis
C1831088|T201|COMP|46992-4|LNC|DYS gene targeted mutation analysis|DYS gene targeted mutation analysis
C1831089|T201|COMP|46993-2|LNC|HLA Ab panel|HLA Ab panel
C1831090|T201|COMP|46994-0|LNC|HLA-A+B+C Ab|HLA-A+B+C Ab
C1831092|T201|COMP|46995-7|LNC|HLA-DP+DQ+DR Ab|HLA-DP+DQ+DR Ab
C1831093|T201|COMP|46996-5|LNC|HLA Ab positive cells|HLA Ab positive cells
C1831095|T201|COMP|46997-3|LNC|HLA Ab cells tested|HLA Ab cells tested
C1831098|T201|COMP|46999-9|LNC|Bacterial vaginosis & vaginitis rRNA panel|Bacterial vaginosis & vaginitis rRNA panel
C1831099|T201|COMP|47000-5|LNC|Candida sp rRNA|Candida sp rRNA
C1831101|T201|COMP|47001-3|LNC|Brucella sp Ag|Brucella sp Ag
C1831102|T201|COMP|47002-1|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1831103|T201|COMP|47003-9|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1831104|T201|COMP|47004-7|LNC|6-Monoacetylmorphine.free|6-Monoacetylmorphine.free
C1831105|T201|COMP|47005-4|LNC|Spermatozoa Ab.IgM/100 spermatozoa|Spermatozoa Ab.IgM/100 spermatozoa
C1831106|T201|COMP|47006-2|LNC|Spermatozoa Ab.IgG/100 spermatozoa|Spermatozoa Ab.IgG/100 spermatozoa
C1831107|T201|COMP|47007-0|LNC|Spermatozoa Ab.IgA/100 spermatozoa|Spermatozoa Ab.IgA/100 spermatozoa
C1831108|T201|COMP|47008-8|LNC|Platelet associated Ab.IgG|Platelet associated Ab.IgG
C1831109|T201|COMP|47009-6|LNC|BCL6 Ag|BCL6 Ag
C1831110|T201|COMP|47010-4|LNC|Ber-EP4 Ag|Ber-EP4 Ag
C1831111|T201|COMP|47011-2|LNC|Calretinin Ag|Calretinin Ag
C1831112|T201|COMP|47012-0|LNC|Cancer Ag 72-4|Cancer Ag 72-4
C1831113|T201|COMP|47013-8|LNC|CD1a Ag|CD1a Ag
C1831114|T201|COMP|47014-6|LNC|CD21 Ag|CD21 Ag
C1831115|T201|COMP|47015-3|LNC|CD31 Ag|CD31 Ag
C1831116|T201|COMP|47016-1|LNC|CD4 Ag|CD4 Ag
C1831117|T201|COMP|47017-9|LNC|CD68 Ag|CD68 Ag
C1831118|T201|COMP|47018-7|LNC|CD79a Ag|CD79a Ag
C1831119|T201|COMP|47019-5|LNC|CD8 Ag|CD8 Ag
C1831120|T201|COMP|47020-3|LNC|CD99 Ag|CD99 Ag
C1831121|T201|COMP|47021-1|LNC|CDX2 Ag|CDX2 Ag
C1831122|T201|COMP|47022-9|LNC|Cells.CD11c+CD19+/100 cells|Cells.CD11c+CD19+/100 cells
C1831123|T201|COMP|47023-7|LNC|Cells.CD19+CD23+/100 cells|Cells.CD19+CD23+/100 cells
C1831124|T201|COMP|47024-5|LNC|Choriogonadotropin.beta subunit Ag|Choriogonadotropin.beta subunit Ag
C1831125|T201|COMP|47025-2|LNC|Cytokeratin 5+6 Ag|Cytokeratin 5+6 Ag
C1831126|T201|COMP|47026-0|LNC|Cytokeratin HMW Ag|Cytokeratin HMW Ag
C1831127|T201|COMP|47027-8|LNC|DBA44 Ag|DBA44 Ag
C1831128|T201|COMP|47028-6|LNC|Follitropin Ag|Follitropin Ag
C1831129|T201|COMP|47029-4|LNC|HIV 2 Ab|HIV 2 Ab
C1831130|T201|COMP|47030-2|LNC|Phosphatidate Ab.IgA|Phosphatidate Ab.IgA
C1831131|T201|COMP|47031-0|LNC|Melan-A Ag|Melan-A Ag
C1831132|T201|COMP|47032-8|LNC|MyoD1 Ag|MyoD1 Ag
C1831133|T201|COMP|47033-6|LNC|Myogenin Ag|Myogenin Ag
C1831134|T201|COMP|47034-4|LNC|Neurofilament Ag|Neurofilament Ag
C1831135|T201|COMP|47035-1|LNC|NKI-C3 Ag|NKI-C3 Ag
C1831136|T201|COMP|47036-9|LNC|Streptococcus pneumoniae 34 Ab.IgG^1st specimen|Streptococcus pneumoniae 34 Ab.IgG^1st specimen
C1831138|T201|COMP|47038-5|LNC|Villin Ag|Villin Ag
C1831151|T201|COMP|47050-0|LNC|Herpes virus 8 Ab.IgG|Herpes virus 8 Ab.IgG
C1831152|T201|COMP|47051-8|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C1831153|T201|COMP|47052-6|LNC|Chlamydophila pneumoniae Ab|Chlamydophila pneumoniae Ab
C1831154|T201|COMP|47053-4|LNC|Enolase.neuron specific|Enolase.neuron specific
C1831155|T201|COMP|47054-2|LNC|Legionella pneumophila 10 Ab.IgM|Legionella pneumophila 10 Ab.IgM
C1831156|T201|COMP|47055-9|LNC|Legionella pneumophila 11 Ab.IgG|Legionella pneumophila 11 Ab.IgG
C1831157|T201|COMP|47056-7|LNC|Legionella pneumophila 11 Ab.IgM|Legionella pneumophila 11 Ab.IgM
C1831158|T201|COMP|47057-5|LNC|Legionella pneumophila 12 Ab.IgG|Legionella pneumophila 12 Ab.IgG
C1831159|T201|COMP|47058-3|LNC|Legionella pneumophila 12 Ab.IgM|Legionella pneumophila 12 Ab.IgM
C1831160|T201|COMP|47059-1|LNC|Legionella pneumophila 13 Ab.IgG|Legionella pneumophila 13 Ab.IgG
C1831161|T201|COMP|47060-9|LNC|Legionella pneumophila 13 Ab.IgM|Legionella pneumophila 13 Ab.IgM
C1831162|T201|COMP|47061-7|LNC|Legionella pneumophila 14 Ab.IgG|Legionella pneumophila 14 Ab.IgG
C1831163|T201|COMP|47062-5|LNC|Legionella pneumophila 14 Ab.IgM|Legionella pneumophila 14 Ab.IgM
C1831164|T201|COMP|47063-3|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C1831165|T201|COMP|47064-1|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C1831166|T201|COMP|47065-8|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C1831167|T201|COMP|47066-6|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C1831168|T201|COMP|47067-4|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C1831169|T201|COMP|47068-2|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C1831170|T201|COMP|47069-0|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C1831171|T201|COMP|47070-8|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C1831172|T201|COMP|47071-6|LNC|Babesia microti Ab.IgG|Babesia microti Ab.IgG
C1831173|T201|COMP|47072-4|LNC|Epstein Barr virus early Ab.IgA|Epstein Barr virus early Ab.IgA
C1831175|T201|COMP|47073-2|LNC|Babesia microti Ab.IgM|Babesia microti Ab.IgM
C1831176|T201|COMP|47074-0|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C1831177|T201|COMP|47075-7|LNC|Coxiella burnetii phase 1 Ab.IgM|Coxiella burnetii phase 1 Ab.IgM
C1831178|T201|COMP|47076-5|LNC|Legionella pneumophila 7 Ab.IgG|Legionella pneumophila 7 Ab.IgG
C1831180|T201|COMP|47077-3|LNC|Legionella pneumophila 7 Ab.IgM|Legionella pneumophila 7 Ab.IgM
C1831182|T201|COMP|47078-1|LNC|Legionella pneumophila 8 Ab.IgG|Legionella pneumophila 8 Ab.IgG
C1831184|T201|COMP|47079-9|LNC|Legionella pneumophila 8 Ab.IgM|Legionella pneumophila 8 Ab.IgM
C1831186|T201|COMP|47080-7|LNC|Legionella pneumophila 9 Ab.IgG|Legionella pneumophila 9 Ab.IgG
C1831188|T201|COMP|47081-5|LNC|Legionella pneumophila 9 Ab.IgM|Legionella pneumophila 9 Ab.IgM
C1831190|T201|COMP|47082-3|LNC|Legionella pneumophila 10 Ab.IgG|Legionella pneumophila 10 Ab.IgG
C1831191|T201|COMP|47083-1|LNC|IgG|IgG
C1831192|T201|COMP|47084-9|LNC|Platelet glycoprotein Ia-IIa Ab|Platelet glycoprotein Ia-IIa Ab
C1831193|T201|COMP|47085-6|LNC|Plasmodium sp DNA|Plasmodium sp DNA
C1831194|T201|COMP|47086-4|LNC|11-Hydroxyandrostenedione|11-Hydroxyandrostenedione
C1831195|T201|COMP|47087-2|LNC|Angiotensinogen|Angiotensinogen
C1831196|T201|COMP|47088-0|LNC|Delta aminolevulinate|Delta aminolevulinate
C1831197|T201|COMP|47089-8|LNC|Indicans|Indicans
C1831198|T201|COMP|47090-6|LNC|Indicans/Creatinine|Indicans/Creatinine
C1831200|T201|COMP|47091-4|LNC|Methylmalonate|Methylmalonate
C1831201|T201|COMP|47092-2|LNC|Natriuretic peptide.B|Natriuretic peptide.B
C1831202|T201|COMP|47093-0|LNC|Parathyrin.biointact|Parathyrin.biointact
C1831203|T201|COMP|47094-8|LNC|Calciferol|Calciferol
C1831204|T201|COMP|47095-5|LNC|Acetaminophen|Acetaminophen
C1831205|T201|COMP|47096-3|LNC|Aluminum|Aluminum
C1831206|T201|COMP|47097-1|LNC|carBAMazepine 10,11-Epoxide.free|carBAMazepine 10,11-Epoxide.free
C1831207|T201|COMP|47098-9|LNC|Chromium|Chromium
C1831208|T201|COMP|47099-7|LNC|Chromium|Chromium
C1831209|T201|COMP|47100-3|LNC|Copper|Copper
C1831210|T201|COMP|47101-1|LNC|Copper|Copper
C1831211|T201|COMP|47102-9|LNC|Copper|Copper
C1831212|T201|COMP|47103-7|LNC|Copper|Copper
C1831213|T201|COMP|47104-5|LNC|Doxepin|Doxepin
C1831214|T201|COMP|47105-2|LNC|ePHEDrine|ePHEDrine
C1831215|T201|COMP|47106-0|LNC|ePHEDrine|ePHEDrine
C1831216|T201|COMP|47107-8|LNC|Ethanol|Ethanol
C1831217|T201|COMP|47108-6|LNC|Furosemide|Furosemide
C1831218|T201|COMP|47109-4|LNC|Gentamicin|Gentamicin
C1831219|T201|COMP|47110-2|LNC|Glutethimide|Glutethimide
C1831220|T201|COMP|47111-0|LNC|Glutethimide|Glutethimide
C1831221|T201|COMP|47112-8|LNC|Gold|Gold
C1831222|T201|COMP|47113-6|LNC|Gold/Creatinine|Gold/Creatinine
C1831223|T201|COMP|47114-4|LNC|LORazepam|LORazepam
C1831224|T201|COMP|47115-1|LNC|LORazepam|LORazepam
C1831225|T201|COMP|47116-9|LNC|Manganese|Manganese
C1831226|T201|COMP|47117-7|LNC|Maprotiline|Maprotiline
C1831227|T201|COMP|47118-5|LNC|Maprotiline|Maprotiline
C1831228|T201|COMP|47119-3|LNC|Meprobamate|Meprobamate
C1831229|T201|COMP|47120-1|LNC|Meprobamate|Meprobamate
C1831230|T201|COMP|47121-9|LNC|Mercury|Mercury
C1831231|T201|COMP|47122-7|LNC|Methyprylon|Methyprylon
C1831232|T201|COMP|47123-5|LNC|Nickel|Nickel
C1831233|T201|COMP|47124-3|LNC|PHENobarbital|PHENobarbital
C1831234|T201|COMP|47125-0|LNC|Primidone|Primidone
C1831235|T201|COMP|47126-8|LNC|Protriptyline|Protriptyline
C1831236|T201|COMP|47127-6|LNC|Protriptyline|Protriptyline
C1831237|T201|COMP|47128-4|LNC|Salicylates|Salicylates
C1831238|T201|COMP|47129-2|LNC|Silver|Silver
C1831239|T201|COMP|47130-0|LNC|Thallium|Thallium
C1831240|T201|COMP|47131-8|LNC|Thioridazine|Thioridazine
C1831241|T201|COMP|47132-6|LNC|Thioridazine|Thioridazine
C1831242|T201|COMP|47133-4|LNC|Trimipramine|Trimipramine
C1831243|T201|COMP|47134-2|LNC|Trimipramine|Trimipramine
C1831244|T201|COMP|47135-9|LNC|Ascorbate^post dose|Ascorbate^post dose
C1831245|T201|COMP|47136-7|LNC|Epinephrine^1H post 300 ug cloNIDine PO|Epinephrine^1H post 300 ug cloNIDine PO
C1831246|T201|COMP|47137-5|LNC|Epinephrine^2H post 300 ug cloNIDine PO|Epinephrine^2H post 300 ug cloNIDine PO
C1831247|T201|COMP|47138-3|LNC|EPINEPHrine^2H post XXX challenge|EPINEPHrine^2H post XXX challenge
C1831248|T201|COMP|47139-1|LNC|EPINEPHrine^2nd specimen post XXX challenge|EPINEPHrine^2nd specimen post XXX challenge
C1831249|T201|COMP|47140-9|LNC|EPINEPHrine^2nd specimen post XXX challenge|EPINEPHrine^2nd specimen post XXX challenge
C1831250|T201|COMP|47141-7|LNC|Epinephrine^3H post 300 ug cloNIDine PO|Epinephrine^3H post 300 ug cloNIDine PO
C1831251|T201|COMP|47142-5|LNC|EPINEPHrine^3rd specimen post XXX challenge|EPINEPHrine^3rd specimen post XXX challenge
C1831252|T201|COMP|47143-3|LNC|EPINEPHrine^3rd specimen post XXX challenge|EPINEPHrine^3rd specimen post XXX challenge
C1831253|T201|COMP|47144-1|LNC|EPINEPHrine^4H post XXX challenge|EPINEPHrine^4H post XXX challenge
C1831254|T201|COMP|47145-8|LNC|EPINEPHrine^4th specimen post XXX challenge|EPINEPHrine^4th specimen post XXX challenge
C1831255|T201|COMP|47146-6|LNC|EPINEPHrine^4th specimen post XXX challenge|EPINEPHrine^4th specimen post XXX challenge
C1831256|T201|COMP|47147-4|LNC|EPINEPHrine^5th specimen post XXX challenge|EPINEPHrine^5th specimen post XXX challenge
C1831257|T201|COMP|47148-2|LNC|EPINEPHrine^5th specimen post XXX challenge|EPINEPHrine^5th specimen post XXX challenge
C1831258|T201|COMP|47149-0|LNC|EPINEPHrine^6th specimen post XXX challenge|EPINEPHrine^6th specimen post XXX challenge
C1831259|T201|COMP|47150-8|LNC|EPINEPHrine^6th specimen post XXX challenge|EPINEPHrine^6th specimen post XXX challenge
C1831260|T201|COMP|47151-6|LNC|EPINEPHrine^7th specimen post XXX challenge|EPINEPHrine^7th specimen post XXX challenge
C1831261|T201|COMP|47152-4|LNC|EPINEPHrine^7th specimen post XXX challenge|EPINEPHrine^7th specimen post XXX challenge
C1831262|T201|COMP|47153-2|LNC|Epinephrine^pre 300 ug cloNIDine PO|Epinephrine^pre 300 ug cloNIDine PO
C1831263|T201|COMP|47154-0|LNC|Lead^post EDTA therapy|Lead^post EDTA therapy
C1831264|T201|COMP|47155-7|LNC|Norepinephrine^10M post standing|Norepinephrine^10M post standing
C1831265|T201|COMP|47156-5|LNC|Norepinephrine^1H post 300 ug clonidine PO|Norepinephrine^1H post 300 ug clonidine PO
C1831266|T201|COMP|47157-3|LNC|Norepinephrine^1H post XXX challenge|Norepinephrine^1H post XXX challenge
C1831267|T201|COMP|47158-1|LNC|Norepinephrine^2H post 300 ug clonidine PO|Norepinephrine^2H post 300 ug clonidine PO
C1831268|T201|COMP|47159-9|LNC|Norepinephrine^2H post XXX challenge|Norepinephrine^2H post XXX challenge
C1831269|T201|COMP|47160-7|LNC|Norepinephrine^2nd specimen post XXX challenge|Norepinephrine^2nd specimen post XXX challenge
C1831270|T201|COMP|47161-5|LNC|Norepinephrine^2nd specimen post XXX challenge|Norepinephrine^2nd specimen post XXX challenge
C1831271|T201|COMP|47162-3|LNC|Norepinephrine^3H post 300 ug clonidine PO|Norepinephrine^3H post 300 ug clonidine PO
C1831272|T201|COMP|47163-1|LNC|Norepinephrine^3H post XXX challenge|Norepinephrine^3H post XXX challenge
C1831273|T201|COMP|47164-9|LNC|Norepinephrine^3rd specimen post XXX challenge|Norepinephrine^3rd specimen post XXX challenge
C1831274|T201|COMP|47165-6|LNC|Norepinephrine^3rd specimen post XXX challenge|Norepinephrine^3rd specimen post XXX challenge
C1831275|T201|COMP|47166-4|LNC|Norepinephrine^4H post XXX challenge|Norepinephrine^4H post XXX challenge
C1831276|T201|COMP|47167-2|LNC|Norepinephrine^4th specimen post XXX challenge|Norepinephrine^4th specimen post XXX challenge
C1831277|T201|COMP|47175-5|LNC|Norepinephrine^pre 300 ug clonidine PO|Norepinephrine^pre 300 ug clonidine PO
C1831278|T201|COMP|47176-3|LNC|Parathyrin.intact^10M post excision|Parathyrin.intact^10M post excision
C1831279|T201|COMP|47177-1|LNC|Parathyrin.intact^5M post excision|Parathyrin.intact^5M post excision
C1831280|T201|COMP|47178-9|LNC|Parathyrin.intact^baseline|Parathyrin.intact^baseline
C1831281|T201|COMP|47179-7|LNC|Parathyrin^10M post excision|Parathyrin^10M post excision
C1831282|T201|COMP|47180-5|LNC|Parathyrin^baseline|Parathyrin^baseline
C1831283|T201|COMP|47181-3|LNC|Progesterone^1.5H post XXX challenge|Progesterone^1.5H post XXX challenge
C1831284|T201|COMP|47182-1|LNC|Progesterone^10th specimen post XXX challenge|Progesterone^10th specimen post XXX challenge
C1831285|T201|COMP|47183-9|LNC|Progesterone^15M post XXX challenge|Progesterone^15M post XXX challenge
C1831286|T201|COMP|47184-7|LNC|Progesterone^1H post XXX challenge|Progesterone^1H post XXX challenge
C1831287|T201|COMP|47185-4|LNC|Progesterone^2H post XXX challenge|Progesterone^2H post XXX challenge
C1831288|T201|COMP|47186-2|LNC|Progesterone^30M post XXX challenge|Progesterone^30M post XXX challenge
C1831289|T201|COMP|47187-0|LNC|Progesterone^45M post XXX challenge|Progesterone^45M post XXX challenge
C1831290|T201|COMP|47188-8|LNC|Progesterone^5th specimen post XXX challenge|Progesterone^5th specimen post XXX challenge
C1831291|T201|COMP|47189-6|LNC|Progesterone^baseline|Progesterone^baseline
C1831292|T201|COMP|47190-4|LNC|Proinsulin^baseline|Proinsulin^baseline
C1831293|T201|COMP|47191-2|LNC|Triiodothyronine^2nd specimen post XXX challenge|Triiodothyronine^2nd specimen post XXX challenge
C1831294|T201|COMP|47192-0|LNC|Triiodothyronine^3rd specimen post XXX challenge|Triiodothyronine^3rd specimen post XXX challenge
C1831295|T201|COMP|47193-8|LNC|Triiodothyronine^4th specimen post XXX challenge|Triiodothyronine^4th specimen post XXX challenge
C1831296|T201|COMP|47194-6|LNC|Triiodothyronine^5th specimen post XXX challenge|Triiodothyronine^5th specimen post XXX challenge
C1831297|T201|COMP|47195-3|LNC|Triiodothyronine^6th specimen post XXX challenge|Triiodothyronine^6th specimen post XXX challenge
C1831298|T201|COMP|47196-1|LNC|Triiodothyronine^7th specimen post XXX challenge|Triiodothyronine^7th specimen post XXX challenge
C1831299|T201|COMP|47197-9|LNC|Triiodothyronine^8th specimen post XXX challenge|Triiodothyronine^8th specimen post XXX challenge
C1831301|T201|COMP|47223-3|LNC|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C1831303|T201|COMP|47225-8|LNC|Bilirubin|Bilirubin
C1831304|T201|COMP|47226-6|LNC|Fetal lung maturity|Fetal lung maturity
C1831305|T201|COMP|47227-4|LNC|Blood.dried|Blood.dried
C1831306|T201|COMP|47228-2|LNC|Cholesterol.non HDL/Cholesterol.total|Cholesterol.non HDL/Cholesterol.total
C1831308|T201|COMP|47229-0|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C1831309|T201|COMP|47230-8|LNC|Herpes simplex virus glycoprotein G Ab.IgG|Herpes simplex virus glycoprotein G Ab.IgG
C1831310|T201|COMP|47231-6|LNC|IgM Ab|IgM Ab
C1831311|T201|COMP|47232-4|LNC|Influenza virus A Ab^1st specimen|Influenza virus A Ab^1st specimen
C1831312|T201|COMP|47233-2|LNC|Influenza virus A Ab^2nd specimen|Influenza virus A Ab^2nd specimen
C1831313|T201|COMP|47234-0|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C1831314|T201|COMP|47235-7|LNC|Reagin Ab|Reagin Ab
C1831315|T201|COMP|47236-5|LNC|Treponema pallidum Ab.IgG+IgM|Treponema pallidum Ab.IgG+IgM
C1831316|T201|COMP|47237-3|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C1831317|T201|COMP|47238-1|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C1831319|T201|COMP|47251-4|LNC|BK virus DNA|BK virus DNA
C1831320|T201|COMP|47252-2|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1831321|T201|COMP|47253-0|LNC|Coproporphyrin 1|Coproporphyrin 1
C1831322|T201|COMP|47254-8|LNC|Coproporphyrin 3|Coproporphyrin 3
C1831323|T201|COMP|47255-5|LNC|Procollagen type I.N-terminal propeptide|Procollagen type I.N-terminal propeptide
C1831324|T201|COMP|47256-3|LNC|Creatinine^2nd specimen post XXX challenge|Creatinine^2nd specimen post XXX challenge
C1831325|T201|COMP|47257-1|LNC|Creatinine^1st specimen post XXX challenge|Creatinine^1st specimen post XXX challenge
C1831326|T201|COMP|47258-9|LNC|Creatinine^3rd specimen post XXX challenge|Creatinine^3rd specimen post XXX challenge
C1831327|T201|COMP|47259-7|LNC|Creatinine^4th specimen post XXX challenge|Creatinine^4th specimen post XXX challenge
C1831328|T201|COMP|47260-5|LNC|Plasmodium sp DNA|Plasmodium sp DNA
C1831329|T201|COMP|47261-3|LNC|Creatinine^6th specimen post XXX challenge|Creatinine^6th specimen post XXX challenge
C1831341|T201|COMP|47273-8|LNC|Creatinine^5th specimen post XXX challenge|Creatinine^5th specimen post XXX challenge
C1831342|T201|COMP|47274-6|LNC|S100 calcium binding protein B|S100 calcium binding protein B
C1831343|T201|COMP|47275-3|LNC|S100 calcium binding protein B|S100 calcium binding protein B
C1831344|T201|COMP|47276-1|LNC|Complement Sc5b-9 Ab|Complement Sc5b-9 Ab
C1831345|T201|COMP|47277-9|LNC|Erythrocyte distribution width|Erythrocyte distribution width
C1831346|T201|COMP|47278-7|LNC|Erythrocyte mean corpuscular hemoglobin|Erythrocyte mean corpuscular hemoglobin
C1831348|T201|COMP|47280-3|LNC|Erythrocytes|Erythrocytes
C1831349|T201|COMP|47281-1|LNC|Leukocytes|Leukocytes
C1831350|T201|COMP|47282-9|LNC|Erythrocyte mean corpuscular volume|Erythrocyte mean corpuscular volume
C1831351|T201|COMP|47283-7|LNC|Platelet mean volume|Platelet mean volume
C1831352|T201|COMP|47284-5|LNC|Platelets|Platelets
C1831353|T201|COMP|47285-2|LNC|Heparin cofactor II Ag|Heparin cofactor II Ag
C1831354|T201|COMP|47286-0|LNC|Differential panel|Differential panel
C1831355|T201|COMP|47287-8|LNC|Hemogram WO platelets panel|Hemogram WO platelets panel
C1831356|T201|COMP|47288-6|LNC|CBC WO Differential panel|CBC WO Differential panel
C1831357|T201|COMP|47289-4|LNC|IgG & IgG subclass panel|IgG & IgG subclass panel
C1831358|T201|COMP|47290-2|LNC|IgG subclass panel|IgG subclass panel
C1831359|T201|COMP|47291-0|LNC|Fungus identified^^^6|Fungus identified^^^6
C1831360|T201|COMP|47292-8|LNC|Fungus identified^^^7|Fungus identified^^^7
C1831361|T201|COMP|47293-6|LNC|Bacteria identified^^^7|Bacteria identified^^^7
C1831362|T201|COMP|47294-4|LNC|Bacteria identified^^^7|Bacteria identified^^^7
C1831363|T201|COMP|47295-1|LNC|Bacteria identified^^^8|Bacteria identified^^^8
C1831365|T201|COMP|47297-7|LNC|Corynebacterium diphtheriae toxin Ab^1st specimen|Corynebacterium diphtheriae toxin Ab^1st specimen
C1831367|T201|COMP|47300-9|LNC|Phosphatidate Ab.IgM|Phosphatidate Ab.IgM
C1831368|T201|COMP|47301-7|LNC|Ribosomal P Ab|Ribosomal P Ab
C1831370|T201|COMP|47303-3|LNC|Anaplastic lymphoma kinase Ag|Anaplastic lymphoma kinase Ag
C1831371|T201|COMP|47304-1|LNC|Borrelia burgdorferi Ab.IgG index|Borrelia burgdorferi Ab.IgG index
C1831373|T201|COMP|47305-8|LNC|BRST 2 Ag|BRST 2 Ag
C1831374|T201|COMP|47306-6|LNC|Cartilage oligomeric matrix protein|Cartilage oligomeric matrix protein
C1831375|T201|COMP|47307-4|LNC|Cytomegalovirus Ab.IgG Index|Cytomegalovirus Ab.IgG Index
C1831377|T201|COMP|47308-2|LNC|Echinococcus granulosus Ab.IgG|Echinococcus granulosus Ab.IgG
C1831378|T201|COMP|47316-5|LNC|Inner Ear 68kD Ab|Inner Ear 68kD Ab
C1831379|T201|COMP|47317-3|LNC|Interleukin 12|Interleukin 12
C1831380|T201|COMP|47318-1|LNC|Liver kidney microsomal 1 Ab.IgG|Liver kidney microsomal 1 Ab.IgG
C1831381|T201|COMP|47319-9|LNC|Myelin basic protein Ab|Myelin basic protein Ab
C1831382|T201|COMP|47320-7|LNC|Saccharomyces cerevisiae Ab.IgA|Saccharomyces cerevisiae Ab.IgA
C1831383|T201|COMP|47321-5|LNC|Saccharomyces cerevisiae Ab.IgG|Saccharomyces cerevisiae Ab.IgG
C1831384|T201|COMP|47322-3|LNC|SCL-70 extractable nuclear Ab.IgG|SCL-70 extractable nuclear Ab.IgG
C1831385|T201|COMP|47323-1|LNC|Streptococcus pneumoniae 17 Ab.IgG|Streptococcus pneumoniae 17 Ab.IgG
C1831386|T201|COMP|47324-9|LNC|Streptococcus pneumoniae 17 Ab.IgG^1st specimen|Streptococcus pneumoniae 17 Ab.IgG^1st specimen
C1831387|T201|COMP|47325-6|LNC|Streptococcus pneumoniae 17 Ab.IgG^2nd specimen|Streptococcus pneumoniae 17 Ab.IgG^2nd specimen
C1831389|T201|COMP|47327-2|LNC|Streptococcus pneumoniae 2 Ab.IgG|Streptococcus pneumoniae 2 Ab.IgG
C1831390|T201|COMP|47328-0|LNC|Streptococcus pneumoniae 2 Ab.IgG^1st specimen|Streptococcus pneumoniae 2 Ab.IgG^1st specimen
C1831391|T201|COMP|47329-8|LNC|Streptococcus pneumoniae 2 Ab.IgG^2nd specimen|Streptococcus pneumoniae 2 Ab.IgG^2nd specimen
C1831393|T201|COMP|47331-4|LNC|Streptococcus pneumoniae 20 Ab.IgG|Streptococcus pneumoniae 20 Ab.IgG
C1831394|T201|COMP|47332-2|LNC|Streptococcus pneumoniae 20 Ab.IgG^1st specimen|Streptococcus pneumoniae 20 Ab.IgG^1st specimen
C1831395|T201|COMP|47333-0|LNC|Streptococcus pneumoniae 20 Ab.IgG^2nd specimen|Streptococcus pneumoniae 20 Ab.IgG^2nd specimen
C1831397|T201|COMP|47335-5|LNC|Streptococcus pneumoniae 22 Ab.IgG|Streptococcus pneumoniae 22 Ab.IgG
C1831398|T201|COMP|47336-3|LNC|Streptococcus pneumoniae 22 Ab.IgG^1st specimen|Streptococcus pneumoniae 22 Ab.IgG^1st specimen
C1831399|T201|COMP|47337-1|LNC|Streptococcus pneumoniae 22 Ab.IgG^2nd specimen|Streptococcus pneumoniae 22 Ab.IgG^2nd specimen
C1831401|T201|COMP|47339-7|LNC|Streptococcus pneumoniae 34 Ab.IgG|Streptococcus pneumoniae 34 Ab.IgG
C1831402|T201|COMP|47340-5|LNC|Streptococcus pneumoniae 34 Ab.IgG^2nd specimen|Streptococcus pneumoniae 34 Ab.IgG^2nd specimen
C1831404|T201|COMP|47342-1|LNC|Streptococcus pneumoniae 43 Ab.IgG|Streptococcus pneumoniae 43 Ab.IgG
C1831405|T201|COMP|47343-9|LNC|Streptococcus pneumoniae 43 Ab.IgG^1st specimen|Streptococcus pneumoniae 43 Ab.IgG^1st specimen
C1831406|T201|COMP|47344-7|LNC|Streptococcus pneumoniae 43 Ab.IgG^2nd specimen|Streptococcus pneumoniae 43 Ab.IgG^2nd specimen
C1831415|T201|COMP|47353-8|LNC|Streptococcus pneumoniae 5 Ab.IgG^1st specimen|Streptococcus pneumoniae 5 Ab.IgG^1st specimen
C1831416|T201|COMP|47354-6|LNC|Streptococcus pneumoniae 5 Ab.IgG^2nd specimen|Streptococcus pneumoniae 5 Ab.IgG^2nd specimen
C1831420|T201|COMP|47358-7|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C1831421|T201|COMP|47359-5|LNC|HIV 1 RNA|HIV 1 RNA
C1831422|T201|COMP|47360-3|LNC|Reagin Ab|Reagin Ab
C1831423|T201|COMP|47361-1|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C1831424|T201|COMP|47362-9|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C1831425|T201|COMP|47363-7|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C1831426|T201|COMP|47364-5|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C1831427|T201|COMP|47386-8|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C1831428|T201|COMP|47387-6|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C1831429|T201|COMP|47388-4|LNC|Salmonella typhi H D Ab|Salmonella typhi H D Ab
C1831430|T201|COMP|47389-2|LNC|Toxoplasma gondii Ab.IgG avidity|Toxoplasma gondii Ab.IgG avidity
C1831431|T201|COMP|47390-0|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C1831432|T201|COMP|47391-8|LNC|Sulfonylurea|Sulfonylurea
C1831433|T201|COMP|47392-6|LNC|chlorproPAMIDE|chlorproPAMIDE
C1831434|T201|COMP|47393-4|LNC|Gliadin peptide Ab.IgA|Gliadin peptide Ab.IgA
C1831435|T201|COMP|47394-2|LNC|Gliadin peptide Ab.IgG|Gliadin peptide Ab.IgG
C1831436|T201|COMP|47395-9|LNC|Kanamycin|Kanamycin
C1831437|T201|COMP|47396-7|LNC|Babesia microti DNA|Babesia microti DNA
C1831438|T201|COMP|47397-5|LNC|BCS1L gene targeted mutation analysis|BCS1L gene targeted mutation analysis
C1831440|T201|COMP|47398-3|LNC|Beta mannosidase actual/Normal|Beta mannosidase actual/Normal
C1831442|T201|COMP|47399-1|LNC|Cells.ZAP70+CD19+/100 cells|Cells.ZAP70+CD19+/100 cells
C1831444|T201|COMP|47400-7|LNC|Cocaine+Benzoylecgonine|Cocaine+Benzoylecgonine
C1831445|T201|COMP|47401-5|LNC|CV2 Ab.IgG|CV2 Ab.IgG
C1831446|T201|COMP|47402-3|LNC|CV2 Ab|CV2 Ab
C1831447|T201|COMP|47403-1|LNC|CYP2D6 gene targeted mutation analysis|CYP2D6 gene targeted mutation analysis
C1831448|T201|COMP|47404-9|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C1831449|T201|COMP|47405-6|LNC|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C1831450|T201|COMP|47406-4|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C1831451|T201|COMP|47407-2|LNC|Fibers|Fibers
C1831452|T201|COMP|47408-0|LNC|Fosphenytoin|Fosphenytoin
C1831453|T201|COMP|47409-8|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1831454|T201|COMP|47410-6|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1831455|T201|COMP|47411-4|LNC|Methadone|Methadone
C1831456|T201|COMP|47412-2|LNC|Mumps virus Ab|Mumps virus Ab
C1831457|T201|COMP|47413-0|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C1831458|T201|COMP|47414-8|LNC|Pregabalin|Pregabalin
C1831459|T201|COMP|47415-5|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C1831460|T201|COMP|47416-3|LNC|RB1 gene targeted mutation analysis|RB1 gene targeted mutation analysis
C1831461|T201|COMP|47417-1|LNC|Red dye Ab.IgE.RAST class|Red dye Ab.IgE.RAST class
C1831463|T201|COMP|47418-9|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C1831464|T201|COMP|47419-7|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C1831467|T201|COMP|47421-3|LNC|Aspergillus flavus B Ab|Aspergillus flavus B Ab
C1831468|T201|COMP|47422-1|LNC|Aspergillus flavus H Ab|Aspergillus flavus H Ab
C1831469|T201|COMP|47423-9|LNC|Aspergillus fumigatus B Ab|Aspergillus fumigatus B Ab
C1831470|T201|COMP|47424-7|LNC|Aspergillus fumigatus H Ab|Aspergillus fumigatus H Ab
C1831471|T201|COMP|47425-4|LNC|Aspergillus nidulans B Ab|Aspergillus nidulans B Ab
C1831472|T201|COMP|47426-2|LNC|Aspergillus nidulans H Ab|Aspergillus nidulans H Ab
C1831473|T201|COMP|47427-0|LNC|Aspergillus niger B Ab|Aspergillus niger B Ab
C1831474|T201|COMP|47428-8|LNC|Aspergillus niger H Ab|Aspergillus niger H Ab
C1831475|T201|COMP|47429-6|LNC|Corynebacterium diphtheriae toxin Ab^1st specimen|Corynebacterium diphtheriae toxin Ab^1st specimen
C1831476|T201|COMP|47430-4|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C1831477|T201|COMP|47431-2|LNC|Echinococcus granulosus Ab.IgG|Echinococcus granulosus Ab.IgG
C1831478|T201|COMP|47432-0|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C1831479|T201|COMP|47433-8|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C1831480|T201|COMP|47434-6|LNC|Epstein Barr virus early diffuse Ab|Epstein Barr virus early diffuse Ab
C1831481|T201|COMP|47435-3|LNC|Epstein Barr virus early Ab.IgA|Epstein Barr virus early Ab.IgA
C1831482|T201|COMP|47436-1|LNC|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C1831483|T201|COMP|47437-9|LNC|Epstein Barr virus early restricted Ab|Epstein Barr virus early restricted Ab
C1831484|T201|COMP|47438-7|LNC|Fowl adenovirus 1 Ab|Fowl adenovirus 1 Ab
C1831485|T201|COMP|47439-5|LNC|Haemophilus influenzae B Ab.IgG^1st specimen|Haemophilus influenzae B Ab.IgG^1st specimen
C1831486|T201|COMP|47440-3|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C1831487|T201|COMP|47441-1|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C1831488|T201|COMP|47442-9|LNC|Herpes virus 8 Ab.IgG|Herpes virus 8 Ab.IgG
C1831489|T201|COMP|47443-7|LNC|Influenza virus A Ab|Influenza virus A Ab
C1831490|T201|COMP|47444-5|LNC|Influenza virus A H1 Ab|Influenza virus A H1 Ab
C1831491|T201|COMP|47445-2|LNC|Influenza virus A H10 Ab|Influenza virus A H10 Ab
C1831492|T201|COMP|47446-0|LNC|Influenza virus A H11 Ab|Influenza virus A H11 Ab
C1831493|T201|COMP|47447-8|LNC|Influenza virus A H12 Ab|Influenza virus A H12 Ab
C1831494|T201|COMP|47448-6|LNC|Influenza virus A H13 Ab|Influenza virus A H13 Ab
C1831495|T201|COMP|47449-4|LNC|Influenza virus A H14 Ab|Influenza virus A H14 Ab
C1831496|T201|COMP|47450-2|LNC|Influenza virus A H15 Ab|Influenza virus A H15 Ab
C1831497|T201|COMP|47451-0|LNC|Influenza virus A H2 Ab|Influenza virus A H2 Ab
C1831498|T201|COMP|47452-8|LNC|Influenza virus A H3 Ab|Influenza virus A H3 Ab
C1831499|T201|COMP|47453-6|LNC|Influenza virus A H4 Ab|Influenza virus A H4 Ab
C1831500|T201|COMP|47454-4|LNC|Influenza virus A H5 Ab|Influenza virus A H5 Ab
C1831501|T201|COMP|47455-1|LNC|Influenza virus A H6 Ab|Influenza virus A H6 Ab
C1831502|T201|COMP|47456-9|LNC|Influenza virus A H7 Ab|Influenza virus A H7 Ab
C1831503|T201|COMP|47457-7|LNC|Influenza virus A H8 Ab|Influenza virus A H8 Ab
C1831504|T201|COMP|47458-5|LNC|Influenza virus A H9 Ab|Influenza virus A H9 Ab
C1831505|T201|COMP|47459-3|LNC|Legionella pneumophila 10 Ab.IgG|Legionella pneumophila 10 Ab.IgG
C1831506|T201|COMP|47460-1|LNC|Legionella pneumophila 10 Ab.IgM|Legionella pneumophila 10 Ab.IgM
C1831507|T201|COMP|47461-9|LNC|Legionella pneumophila 11 Ab.IgG|Legionella pneumophila 11 Ab.IgG
C1831508|T201|COMP|47462-7|LNC|Legionella pneumophila 11 Ab.IgM|Legionella pneumophila 11 Ab.IgM
C1831509|T201|COMP|47463-5|LNC|Legionella pneumophila 12 Ab.IgG|Legionella pneumophila 12 Ab.IgG
C1831510|T201|COMP|47464-3|LNC|Legionella pneumophila 12 Ab.IgM|Legionella pneumophila 12 Ab.IgM
C1831511|T201|COMP|47465-0|LNC|Legionella pneumophila 13 Ab.IgG|Legionella pneumophila 13 Ab.IgG
C1831512|T201|COMP|47466-8|LNC|Legionella pneumophila 13 Ab.IgM|Legionella pneumophila 13 Ab.IgM
C1831513|T201|COMP|47467-6|LNC|Legionella pneumophila 14 Ab.IgG|Legionella pneumophila 14 Ab.IgG
C1831514|T201|COMP|47468-4|LNC|Legionella pneumophila 14 Ab.IgM|Legionella pneumophila 14 Ab.IgM
C1831515|T201|COMP|47469-2|LNC|Legionella pneumophila 7 Ab.IgG|Legionella pneumophila 7 Ab.IgG
C1831516|T201|COMP|47470-0|LNC|Legionella pneumophila 7 Ab.IgM|Legionella pneumophila 7 Ab.IgM
C1831517|T201|COMP|47471-8|LNC|Legionella pneumophila 8 Ab.IgG|Legionella pneumophila 8 Ab.IgG
C1831518|T201|COMP|47472-6|LNC|Legionella pneumophila 8 Ab.IgM|Legionella pneumophila 8 Ab.IgM
C1831519|T201|COMP|47473-4|LNC|Legionella pneumophila 9 Ab.IgG|Legionella pneumophila 9 Ab.IgG
C1831520|T201|COMP|47474-2|LNC|Legionella pneumophila 9 Ab.IgM|Legionella pneumophila 9 Ab.IgM
C1831521|T201|COMP|47475-9|LNC|Powassan virus polyvalent E Ab|Powassan virus polyvalent E Ab
C1831522|T201|COMP|47476-7|LNC|Reagin Ab|Reagin Ab
C1831523|T201|COMP|47477-5|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C1831524|T201|COMP|47478-3|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C1831525|T201|COMP|47479-1|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C1831526|T201|COMP|47480-9|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C1831527|T201|COMP|47481-7|LNC|Streptococcus pneumoniae 1 Ab.IgG^1st specimen|Streptococcus pneumoniae 1 Ab.IgG^1st specimen
C1831528|T201|COMP|47482-5|LNC|Streptococcus pneumoniae 1 Ab.IgG^2nd specimen|Streptococcus pneumoniae 1 Ab.IgG^2nd specimen
C1831529|T201|COMP|47483-3|LNC|Streptococcus pneumoniae 14 Ab.IgG^1st specimen|Streptococcus pneumoniae 14 Ab.IgG^1st specimen
C1831530|T201|COMP|47484-1|LNC|Streptococcus pneumoniae 14 Ab.IgG^2nd specimen|Streptococcus pneumoniae 14 Ab.IgG^2nd specimen
C1831531|T201|COMP|47485-8|LNC|Streptococcus pneumoniae 17 Ab.IgG^1st specimen|Streptococcus pneumoniae 17 Ab.IgG^1st specimen
C1831532|T201|COMP|47486-6|LNC|Streptococcus pneumoniae 17 Ab.IgG^2nd specimen|Streptococcus pneumoniae 17 Ab.IgG^2nd specimen
C1831533|T201|COMP|47487-4|LNC|Streptococcus pneumoniae 2 Ab.IgG^1st specimen|Streptococcus pneumoniae 2 Ab.IgG^1st specimen
C1831534|T201|COMP|47488-2|LNC|Streptococcus pneumoniae 2 Ab.IgG^2nd specimen|Streptococcus pneumoniae 2 Ab.IgG^2nd specimen
C1831535|T201|COMP|47489-0|LNC|Streptococcus pneumoniae 20 Ab.IgG^1st specimen|Streptococcus pneumoniae 20 Ab.IgG^1st specimen
C1831536|T201|COMP|47490-8|LNC|Streptococcus pneumoniae 20 Ab.IgG^2nd specimen|Streptococcus pneumoniae 20 Ab.IgG^2nd specimen
C1831537|T201|COMP|47491-6|LNC|Streptococcus pneumoniae 22 Ab.IgG^1st specimen|Streptococcus pneumoniae 22 Ab.IgG^1st specimen
C1831538|T201|COMP|47492-4|LNC|Streptococcus pneumoniae 22 Ab.IgG^2nd specimen|Streptococcus pneumoniae 22 Ab.IgG^2nd specimen
C1831539|T201|COMP|47493-2|LNC|Streptococcus pneumoniae 3 Ab.IgG^1st specimen|Streptococcus pneumoniae 3 Ab.IgG^1st specimen
C1831540|T201|COMP|47494-0|LNC|Streptococcus pneumoniae 3 Ab.IgG^2nd specimen|Streptococcus pneumoniae 3 Ab.IgG^2nd specimen
C1831541|T201|COMP|47495-7|LNC|Streptococcus pneumoniae 34 Ab.IgG^1st specimen|Streptococcus pneumoniae 34 Ab.IgG^1st specimen
C1831542|T201|COMP|47496-5|LNC|Streptococcus pneumoniae 34 Ab.IgG^2nd specimen|Streptococcus pneumoniae 34 Ab.IgG^2nd specimen
C1831543|T201|COMP|47497-3|LNC|Streptococcus pneumoniae 43 Ab.IgG^1st specimen|Streptococcus pneumoniae 43 Ab.IgG^1st specimen
C1831544|T201|COMP|47498-1|LNC|Streptococcus pneumoniae 43 Ab.IgG^2nd specimen|Streptococcus pneumoniae 43 Ab.IgG^2nd specimen
C1831545|T201|COMP|47499-9|LNC|Streptococcus pneumoniae 5 Ab.IgG^1st specimen|Streptococcus pneumoniae 5 Ab.IgG^1st specimen
C1831546|T201|COMP|47500-4|LNC|Streptococcus pneumoniae 5 Ab.IgG^2nd specimen|Streptococcus pneumoniae 5 Ab.IgG^2nd specimen
C1831551|T201|COMP|47505-3|LNC|Streptococcus pneumoniae 6 Ab.IgG|Streptococcus pneumoniae 6 Ab.IgG
C1831557|T201|COMP|47511-1|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1831558|T201|COMP|47512-9|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C1831559|T201|COMP|47513-7|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C1831560|T201|COMP|47514-5|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C1831561|T201|COMP|47515-2|LNC|Vesicular stomatitis Indiana virus 1 Ab|Vesicular stomatitis Indiana virus 1 Ab
C1831562|T201|COMP|47516-0|LNC|Cocal virus Ab|Cocal virus Ab
C1831563|T201|COMP|47517-8|LNC|Vesicular stomatitis Alagoas virus Ab|Vesicular stomatitis Alagoas virus Ab
C1831564|T201|COMP|47518-6|LNC|Yersinia pestis Ab|Yersinia pestis Ab
C1831567|T201|COMP|47520-2|LNC|Cytology report|Cytology report
C1831568|T201|COMP|47521-0|LNC|Cytology report|Cytology report
C1831569|T201|COMP|47522-8|LNC|Cytology report|Cytology report
C1831570|T201|COMP|47523-6|LNC|Cytology report|Cytology report
C1831571|T201|COMP|47524-4|LNC|Cytology report|Cytology report
C1831572|T201|COMP|47525-1|LNC|Cytology report|Cytology report
C1831573|T201|COMP|47526-9|LNC|Cytology report|Cytology report
C1831574|T201|COMP|47527-7|LNC|Cytology report|Cytology report
C1831575|T201|COMP|47528-5|LNC|Cytology report|Cytology report
C1831576|T201|COMP|47529-3|LNC|Cytology report|Cytology report
C1831577|T201|COMP|47530-1|LNC|Cytology report|Cytology report
C1831578|T201|COMP|47531-9|LNC|Wet mount panel|Wet mount panel
C1831586|T201|COMP|46972-6|LNC|6-Monoacetylmorphine.free|6-Monoacetylmorphine.free
C1831587|T201|COMP|47299-3|LNC|DNA double strand Ab|DNA double strand Ab
C1879319|T201|COMP|1187-4|LNC|little i NOS Ag|little i NOS Ag
C1952627|T201|COMP|47667-1|LNC|Insulin^6M post dose glucagon|Insulin^6M post dose glucagon
C1952628|T201|COMP|47668-9|LNC|Insulin^pre dose glucose|Insulin^pre dose glucose
C1952629|T201|COMP|47669-7|LNC|Insulin^pre dose glucagon|Insulin^pre dose glucagon
C1952630|T201|COMP|47670-5|LNC|Insulin^pre-meal|Insulin^pre-meal
C1952631|T201|COMP|47671-3|LNC|Isoleucine|Isoleucine
C1952632|T201|COMP|47672-1|LNC|Isoleucine/Amino acids.total|Isoleucine/Amino acids.total
C1952634|T201|COMP|47673-9|LNC|Isoleucine/Amino acids.total|Isoleucine/Amino acids.total
C1952644|T201|COMP|47666-3|LNC|Insulin^5M pre dose glucose|Insulin^5M pre dose glucose
C1952645|T201|COMP|47838-8|LNC|Carnitine acyltransferase II|Carnitine acyltransferase II
C1952646|T201|COMP|47839-6|LNC|Carnitine acyltransferase II|Carnitine acyltransferase II
C1952647|T201|COMP|47840-4|LNC|Carnitine acyltransferase II|Carnitine acyltransferase II
C1952648|T201|COMP|47841-2|LNC|Citrate synthase|Citrate synthase
C1952649|T201|COMP|47842-0|LNC|Collection duration|Collection duration
C1952650|T201|COMP|47843-8|LNC|Corticotropin^post dose dexamethasone|Corticotropin^post dose dexamethasone
C1952651|T201|COMP|47844-6|LNC|Cortisol^post 1 mg dexamethasone PO overnight|Cortisol^post 1 mg dexamethasone PO overnight
C1952658|T201|COMP|47563-2|LNC|Arginine/Amino acids.total|Arginine/Amino acids.total
C1952660|T201|COMP|47564-0|LNC|Arginine/Amino acids.total|Arginine/Amino acids.total
C1952661|T201|COMP|47565-7|LNC|Arginine/Amino acids.total|Arginine/Amino acids.total
C1952662|T201|COMP|47566-5|LNC|Arginine/Amino acids.total|Arginine/Amino acids.total
C1952663|T201|COMP|47567-3|LNC|Arginine/Amino acids.total|Arginine/Amino acids.total
C1952664|T201|COMP|47568-1|LNC|Arginine/Amino acids.total|Arginine/Amino acids.total
C1952665|T201|COMP|47569-9|LNC|Argininosuccinate lyase|Argininosuccinate lyase
C1952666|T201|COMP|47570-7|LNC|Argininosuccinate lyase|Argininosuccinate lyase
C1952667|T201|COMP|47571-5|LNC|Argininosuccinate synthase|Argininosuccinate synthase
C1952668|T201|COMP|47572-3|LNC|Asparagine|Asparagine
C1952669|T201|COMP|47573-1|LNC|Aspartate|Aspartate
C1952670|T201|COMP|47574-9|LNC|Aspartate/Amino acids.total|Aspartate/Amino acids.total
C1952672|T201|COMP|47575-6|LNC|Aspartate/Amino acids.total|Aspartate/Amino acids.total
C1952673|T201|COMP|48126-7|LNC|Somatotropin^15M pre dose ornithine|Somatotropin^15M pre dose ornithine
C1952674|T201|COMP|48127-5|LNC|Somatotropin^15M pre dose TRH|Somatotropin^15M pre dose TRH
C1952675|T201|COMP|48128-3|LNC|Somatotropin^1H post dose arginine+insulin|Somatotropin^1H post dose arginine+insulin
C1952676|T201|COMP|48129-1|LNC|Somatotropin^30M pre dose betaxolol+glucagon|Somatotropin^30M pre dose betaxolol+glucagon
C1952677|T201|COMP|48130-9|LNC|Somatotropin^30M pre dose propranolol+glucagon|Somatotropin^30M pre dose propranolol+glucagon
C1952678|T201|COMP|48131-7|LNC|Somatotropin^30M pre dose TRH|Somatotropin^30M pre dose TRH
C1952679|T201|COMP|48132-5|LNC|Xylitol/Creatinine|Xylitol/Creatinine
C1952681|T201|COMP|48133-3|LNC|3-Oxovalerate|3-Oxovalerate
C1952683|T201|COMP|48134-1|LNC|Alanine aminotransferase.macromolecular|Alanine aminotransferase.macromolecular
C1952685|T201|COMP|48135-8|LNC|Acadesine|Acadesine
C1952686|T201|COMP|48136-6|LNC|Aspartate aminotransferase.macromolecular|Aspartate aminotransferase.macromolecular
C1952688|T201|COMP|48137-4|LNC|4,5-Dihydroxyhexanoate/Creatinine|4,5-Dihydroxyhexanoate/Creatinine
C1952690|T201|COMP|48364-4|LNC|Morphine-3-Glucuronide|Morphine-3-Glucuronide
C1952691|T201|COMP|48365-1|LNC|Methadone.R|Methadone.R
C1952692|T201|COMP|48366-9|LNC|Pentadecanoate|Pentadecanoate
C1952694|T201|COMP|48367-7|LNC|cis-Vaccenate|cis-Vaccenate
C1952696|T201|COMP|48368-5|LNC|trans-Octadecanoate|trans-Octadecanoate
C1952698|T201|COMP|48369-3|LNC|trans-Vaccenate|trans-Vaccenate
C1952700|T201|COMP|48370-1|LNC|Dihomogammalinolenate|Dihomogammalinolenate
C1952702|T201|COMP|48379-2|LNC|Zopiclone|Zopiclone
C1952703|T201|COMP|48380-0|LNC|3-Methoxytyramine|3-Methoxytyramine
C1952704|T201|COMP|48381-8|LNC|3-Methoxytyramine/Creatinine|3-Methoxytyramine/Creatinine
C1952706|T201|COMP|48382-6|LNC|Fatty acids.omega 6/Fatty acids.omega 3|Fatty acids.omega 6/Fatty acids.omega 3
C1952708|T201|COMP|48383-4|LNC|Collagen.bovine type 1 Ab|Collagen.bovine type 1 Ab
C1952710|T201|COMP|48384-2|LNC|Collagen.bovine type 2 Ab|Collagen.bovine type 2 Ab
C1952714|T201|COMP|48493-1|LNC|Beta-trace protein|Beta-trace protein
C1952715|T201|COMP|48984-9|LNC|Glucose^10M post dose glucose|Glucose^10M post dose glucose
C1952716|T201|COMP|48985-6|LNC|Glucose^20M post dose glucose|Glucose^20M post dose glucose
C1952717|T201|COMP|48986-4|LNC|Glucose^8 AM specimen|Glucose^8 AM specimen
C1952718|T201|COMP|48987-2|LNC|Pyridinoline.free/Creatinine|Pyridinoline.free/Creatinine
C1952720|T201|COMP|48988-0|LNC|Glucose^12 PM specimen|Glucose^12 PM specimen
C1952721|T201|COMP|48989-8|LNC|Glucose^6 PM specimen|Glucose^6 PM specimen
C1952722|T201|COMP|48990-6|LNC|Glucose^8 PM specimen|Glucose^8 PM specimen
C1952723|T201|COMP|49208-2|LNC|Bartonella elizabethae Ab.IgG|Bartonella elizabethae Ab.IgG
C1952725|T201|COMP|49209-0|LNC|Bartonella bacilliformis Ab.IgM|Bartonella bacilliformis Ab.IgM
C1952727|T201|COMP|49210-8|LNC|Bartonella bacilliformis Ab.IgG|Bartonella bacilliformis Ab.IgG
C1952729|T201|COMP|49211-6|LNC|Bartonella bacilliformis Ab.IgM|Bartonella bacilliformis Ab.IgM
C1952730|T201|COMP|49212-4|LNC|Bartonella bacilliformis Ab.IgG|Bartonella bacilliformis Ab.IgG
C1952731|T201|COMP|49213-2|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1952732|T201|COMP|49214-0|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1952733|T201|COMP|49215-7|LNC|PKHD1 gene targeted mutation analysis|PKHD1 gene targeted mutation analysis
C1952735|T201|COMP|47532-7|LNC|Mumps virus RNA|Mumps virus RNA
C1952737|T201|COMP|47534-3|LNC|2-Hydroxyphenylacetate/Creatinine|2-Hydroxyphenylacetate/Creatinine
C1952738|T201|COMP|47535-0|LNC|2-Methyl,3-Hydroxybutyrate/Creatinine|2-Methyl,3-Hydroxybutyrate/Creatinine
C1952740|T201|COMP|47536-8|LNC|3-Hydroxypropionate|3-Hydroxypropionate
C1952741|T201|COMP|47537-6|LNC|3-Hydroxysebacate/Creatinine|3-Hydroxysebacate/Creatinine
C1952743|T201|COMP|47538-4|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C1952744|T201|COMP|47539-2|LNC|3-Methylhistidine|3-Methylhistidine
C1952745|T201|COMP|47540-0|LNC|3-Methylhistidine|3-Methylhistidine
C1952746|T201|COMP|47541-8|LNC|4-Hydroxybenzoate/Creatinine|4-Hydroxybenzoate/Creatinine
C1952748|T201|COMP|47542-6|LNC|Gamma hydroxybutyrate/Creatinine|Gamma hydroxybutyrate/Creatinine
C1952749|T201|COMP|47543-4|LNC|4-Hydroxymandelate/Creatinine|4-Hydroxymandelate/Creatinine
C1952750|T201|COMP|47544-2|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C1952751|T201|COMP|47545-9|LNC|5-Hydroxyindoleacetate/Creatinine|5-Hydroxyindoleacetate/Creatinine
C1952752|T201|COMP|47546-7|LNC|5-Hydroxytryptophan|5-Hydroxytryptophan
C1952753|T201|COMP|47547-5|LNC|5-Methyltetrahydrofolate|5-Methyltetrahydrofolate
C1952754|T201|COMP|47548-3|LNC|Adenosine deaminase|Adenosine deaminase
C1952755|T201|COMP|47549-1|LNC|Adenosine deaminase|Adenosine deaminase
C1952756|T201|COMP|47550-9|LNC|Adenosine deaminase|Adenosine deaminase
C1952757|T201|COMP|47551-7|LNC|Alanine|Alanine
C1952758|T201|COMP|48119-2|LNC|Pentadecanoate/Creatinine|Pentadecanoate/Creatinine
C1952760|T201|COMP|48120-0|LNC|Prolactin^15M pre dose TRH IV|Prolactin^15M pre dose TRH IV
C1952761|T201|COMP|48121-8|LNC|Quinolinate/Creatinine|Quinolinate/Creatinine
C1952763|T201|COMP|48122-6|LNC|Somatotropin^15M post dose TRH|Somatotropin^15M post dose TRH
C1952764|T201|COMP|48123-4|LNC|Somatotropin^15M pre dose arginine+insulin|Somatotropin^15M pre dose arginine+insulin
C1952765|T201|COMP|48124-2|LNC|Somatotropin^15M pre dose glucagon|Somatotropin^15M pre dose glucagon
C1952766|T201|COMP|48125-9|LNC|Somatotropin^15M pre dose insulin IV|Somatotropin^15M pre dose insulin IV
C1952767|T201|COMP|48199-4|LNC|Ampicillin leukotriene release|Ampicillin leukotriene release
C1952769|T201|COMP|48200-0|LNC|Penicillin V leukotriene release|Penicillin V leukotriene release
C1952771|T201|COMP|48201-8|LNC|Penicillin G leukotriene release|Penicillin G leukotriene release
C1952775|T201|COMP|48203-4|LNC|Apium graveolens leukotriene release|Apium graveolens leukotriene release
C1952777|T201|COMP|48204-2|LNC|Casein leukotriene release|Casein leukotriene release
C1952779|T201|COMP|48205-9|LNC|Beta lactoglobulin leukotriene release|Beta lactoglobulin leukotriene release
C1952781|T201|COMP|49110-0|LNC|Mycoplasma sp identified|Mycoplasma sp identified
C1952782|T201|COMP|49111-8|LNC|Spermatozoa|Spermatozoa
C1952783|T201|COMP|49112-6|LNC|Borna disease virus Ab|Borna disease virus Ab
C1952785|T201|COMP|49113-4|LNC|ZAP70 Ag|ZAP70 Ag
C1952787|T201|COMP|49114-2|LNC|Flavivirus rRNA|Flavivirus rRNA
C1952789|T201|COMP|49115-9|LNC|Thiamine.free|Thiamine.free
C1952791|T201|COMP|49116-7|LNC|Trichosporon sp DNA|Trichosporon sp DNA
C1952793|T201|COMP|49117-5|LNC|Norovirus Ag|Norovirus Ag
C1952794|T201|COMP|47552-5|LNC|Alanine/Amino acids.total|Alanine/Amino acids.total
C1952796|T201|COMP|47553-3|LNC|Alanine/Amino acids.total|Alanine/Amino acids.total
C1952797|T201|COMP|47554-1|LNC|Alanine/Amino acids.total|Alanine/Amino acids.total
C1952798|T201|COMP|47555-8|LNC|Alanine/Amino acids.total|Alanine/Amino acids.total
C1952799|T201|COMP|47556-6|LNC|Alanine/Amino acids.total|Alanine/Amino acids.total
C1952800|T201|COMP|47557-4|LNC|Alanine/Amino acids.total|Alanine/Amino acids.total
C1952801|T201|COMP|47558-2|LNC|Albumin/Protein.total|Albumin/Protein.total
C1952802|T201|COMP|47559-0|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C1952803|T201|COMP|47560-8|LNC|Androstenedione^pre 250 ug corticotropin IM|Androstenedione^pre 250 ug corticotropin IM
C1952804|T201|COMP|47561-6|LNC|Anion gap|Anion gap
C1952805|T201|COMP|47562-4|LNC|Arginine|Arginine
C1952806|T201|COMP|47576-4|LNC|Aspartate/Amino acids.total|Aspartate/Amino acids.total
C1952807|T201|COMP|47577-2|LNC|Aspartate/Amino acids.total|Aspartate/Amino acids.total
C1952808|T201|COMP|47578-0|LNC|Aspartate/Amino acids.total|Aspartate/Amino acids.total
C1952809|T201|COMP|47579-8|LNC|Bicarbonate|Bicarbonate
C1952810|T201|COMP|47580-6|LNC|Bicarbonate|Bicarbonate
C1952811|T201|COMP|47581-4|LNC|Biopterin|Biopterin
C1952812|T201|COMP|47582-2|LNC|Biopterin/Creatinine|Biopterin/Creatinine
C1952814|T201|COMP|47583-0|LNC|C peptide^1.5H post dose glucose|C peptide^1.5H post dose glucose
C1952815|T201|COMP|47584-8|LNC|C peptide^10M post dose glucose|C peptide^10M post dose glucose
C1952816|T201|COMP|47585-5|LNC|C peptide^15M post dose glucose|C peptide^15M post dose glucose
C1952817|T201|COMP|47586-3|LNC|C peptide^1H post dose glucose|C peptide^1H post dose glucose
C1952818|T201|COMP|47587-1|LNC|C peptide^1M post dose glucose|C peptide^1M post dose glucose
C1952819|T201|COMP|47588-9|LNC|C peptide^2H post dose glucose|C peptide^2H post dose glucose
C1952820|T201|COMP|47589-7|LNC|C peptide^30M post dose glucose|C peptide^30M post dose glucose
C1952821|T201|COMP|47590-5|LNC|C peptide^3H post dose glucose|C peptide^3H post dose glucose
C1952822|T201|COMP|47591-3|LNC|C peptide^3M post dose glucose|C peptide^3M post dose glucose
C1952823|T201|COMP|47592-1|LNC|C peptide^5M post dose glucose|C peptide^5M post dose glucose
C1952824|T201|COMP|47593-9|LNC|C peptide^5M pre dose glucose|C peptide^5M pre dose glucose
C1952825|T201|COMP|47594-7|LNC|C peptide^pre dose glucagon|C peptide^pre dose glucagon
C1952826|T201|COMP|47595-4|LNC|C peptide^pre dose glucose|C peptide^pre dose glucose
C1952827|T201|COMP|47596-2|LNC|Calcium.ionized|Calcium.ionized
C1952828|T201|COMP|47597-0|LNC|Calcium^^corrected for total protein|Calcium^^corrected for total protein
C1952829|T201|COMP|47598-8|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C1952831|T201|COMP|47600-2|LNC|Ceruloplasmin|Ceruloplasmin
C1952832|T201|COMP|47601-0|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C1952833|T201|COMP|47602-8|LNC|Citrate synthase|Citrate synthase
C1952834|T201|COMP|47603-6|LNC|Citrate synthase|Citrate synthase
C1952835|T201|COMP|47604-4|LNC|Cortisol^1.5H post 1 ug/kg CRH IV|Cortisol^1.5H post 1 ug/kg CRH IV
C1952836|T201|COMP|47605-1|LNC|Cortisol^15M post 1 ug/kg CRH IV|Cortisol^15M post 1 ug/kg CRH IV
C1952837|T201|COMP|47606-9|LNC|Cortisol^1H post 1 ug/kg CRH IV|Cortisol^1H post 1 ug/kg CRH IV
C1952838|T201|COMP|47607-7|LNC|Cortisol^30M post 1 ug/kg CRH IV|Cortisol^30M post 1 ug/kg CRH IV
C1952839|T201|COMP|47608-5|LNC|Cortisol^pre dose corticotropin|Cortisol^pre dose corticotropin
C1952840|T201|COMP|47609-3|LNC|Cortisol^pre 1 ug/kg CRH IV|Cortisol^pre 1 ug/kg CRH IV
C1952841|T201|COMP|47610-1|LNC|Creatinine|Creatinine
C1952842|T201|COMP|47611-9|LNC|Crystals|Crystals
C1952843|T201|COMP|47612-7|LNC|Cystatin C|Cystatin C
C1952844|T201|COMP|47613-5|LNC|Decanoate/Creatinine|Decanoate/Creatinine
C1952846|T201|COMP|47614-3|LNC|Decenoate/Creatinine|Decenoate/Creatinine
C1952848|T201|COMP|47615-0|LNC|Dermatan sulfate|Dermatan sulfate
C1952849|T201|COMP|47616-8|LNC|Estradiol^1H post dose corticotropin|Estradiol^1H post dose corticotropin
C1952850|T201|COMP|47617-6|LNC|Estradiol^pre dose corticotropin|Estradiol^pre dose corticotropin
C1952853|T201|COMP|47620-0|LNC|Glucose|Glucose
C1952854|T201|COMP|47621-8|LNC|Glucose.IV|Glucose.IV
C1952856|T201|COMP|47622-6|LNC|Glucose^pre dose glucose|Glucose^pre dose glucose
C1952857|T201|COMP|47623-4|LNC|Glutamate|Glutamate
C1952858|T201|COMP|47624-2|LNC|Glutamate/Amino acids.total|Glutamate/Amino acids.total
C1952860|T201|COMP|47625-9|LNC|Glutamate/Amino acids.total|Glutamate/Amino acids.total
C1952861|T201|COMP|47626-7|LNC|Glutamate/Amino acids.total|Glutamate/Amino acids.total
C1952862|T201|COMP|47627-5|LNC|Glutamate/Amino acids.total|Glutamate/Amino acids.total
C1952863|T201|COMP|47628-3|LNC|Glutamate/Amino acids.total|Glutamate/Amino acids.total
C1952864|T201|COMP|47629-1|LNC|Glutamate/Amino acids.total|Glutamate/Amino acids.total
C1952865|T201|COMP|47630-9|LNC|Glutamine|Glutamine
C1952866|T201|COMP|47631-7|LNC|Glutathione.oxidized|Glutathione.oxidized
C1952867|T201|COMP|47632-5|LNC|Glycerol/Creatinine|Glycerol/Creatinine
C1952869|T201|COMP|47633-3|LNC|Glycine|Glycine
C1952870|T201|COMP|47634-1|LNC|Glycine/Amino acids.total|Glycine/Amino acids.total
C1952872|T201|COMP|47635-8|LNC|Glycine/Amino acids.total|Glycine/Amino acids.total
C1952873|T201|COMP|47636-6|LNC|Glycine/Amino acids.total|Glycine/Amino acids.total
C1952874|T201|COMP|47637-4|LNC|Glycine/Amino acids.total|Glycine/Amino acids.total
C1952875|T201|COMP|47638-2|LNC|Glycine/Amino acids.total|Glycine/Amino acids.total
C1952876|T201|COMP|47639-0|LNC|Glycine/Amino acids.total|Glycine/Amino acids.total
C1952877|T201|COMP|47640-8|LNC|Hematocrit|Hematocrit
C1952878|T201|COMP|47641-6|LNC|Palmitate/Creatinine|Palmitate/Creatinine
C1952880|T201|COMP|47642-4|LNC|Hexadecenoate/Creatinine|Hexadecenoate/Creatinine
C1952882|T201|COMP|47643-2|LNC|Histidine|Histidine
C1952883|T201|COMP|47644-0|LNC|Histidine/Amino acids.total|Histidine/Amino acids.total
C1952885|T201|COMP|47645-7|LNC|Histidine/Amino acids.total|Histidine/Amino acids.total
C1952886|T201|COMP|47646-5|LNC|Histidine/Amino acids.total|Histidine/Amino acids.total
C1952887|T201|COMP|47647-3|LNC|Histidine/Amino acids.total|Histidine/Amino acids.total
C1952888|T201|COMP|47648-1|LNC|Histidine/Amino acids.total|Histidine/Amino acids.total
C1952889|T201|COMP|47649-9|LNC|Histidine/Amino acids.total|Histidine/Amino acids.total
C1952890|T201|COMP|47650-7|LNC|Homogentisate/Creatinine|Homogentisate/Creatinine
C1952892|T201|COMP|47651-5|LNC|Hydroxyproline|Hydroxyproline
C1952893|T201|COMP|47652-3|LNC|Hypoxanthine phosphoribosyltransferase|Hypoxanthine phosphoribosyltransferase
C1952894|T201|COMP|47653-1|LNC|Insulin^10M post dose glucagon|Insulin^10M post dose glucagon
C1952895|T201|COMP|47654-9|LNC|Insulin^10M post dose glucose|Insulin^10M post dose glucose
C1952896|T201|COMP|47655-6|LNC|Insulin^15M post dose glucagon|Insulin^15M post dose glucagon
C1952897|T201|COMP|47656-4|LNC|Insulin^1M post dose glucose|Insulin^1M post dose glucose
C1952898|T201|COMP|47657-2|LNC|Insulin^1H post dose glucose|Insulin^1H post dose glucose
C1952899|T201|COMP|47658-0|LNC|Insulin^1.5H post dose glucose|Insulin^1.5H post dose glucose
C1952900|T201|COMP|47659-8|LNC|Insulin^2H post dose glucose|Insulin^2H post dose glucose
C1952901|T201|COMP|47660-6|LNC|Insulin^2.5H post dose glucose|Insulin^2.5H post dose glucose
C1952902|T201|COMP|47661-4|LNC|Insulin^20M post dose glucose|Insulin^20M post dose glucose
C1952903|T201|COMP|47662-2|LNC|Insulin^3H post dose glucose|Insulin^3H post dose glucose
C1952904|T201|COMP|47663-0|LNC|Insulin^30M post dose glucose|Insulin^30M post dose glucose
C1952905|T201|COMP|47664-8|LNC|Insulin^3M post dose glucose|Insulin^3M post dose glucose
C1952906|T201|COMP|47665-5|LNC|Insulin^5M post dose glucose|Insulin^5M post dose glucose
C1952907|T201|COMP|47674-7|LNC|Isoleucine/Amino acids.total|Isoleucine/Amino acids.total
C1952908|T201|COMP|47675-4|LNC|Isoleucine/Amino acids.total|Isoleucine/Amino acids.total
C1952909|T201|COMP|47676-2|LNC|Isoleucine/Amino acids.total|Isoleucine/Amino acids.total
C1952910|T201|COMP|47677-0|LNC|Isoleucine/Amino acids.total|Isoleucine/Amino acids.total
C1952911|T201|COMP|47678-8|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C1952912|T201|COMP|47679-6|LNC|Leucine|Leucine
C1952913|T201|COMP|47680-4|LNC|Leucine/Amino acids.total|Leucine/Amino acids.total
C1952915|T201|COMP|47681-2|LNC|Leucine/Amino acids.total|Leucine/Amino acids.total
C1952916|T201|COMP|47682-0|LNC|Leucine/Amino acids.total|Leucine/Amino acids.total
C1952917|T201|COMP|47683-8|LNC|Leucine/Amino acids.total|Leucine/Amino acids.total
C1952918|T201|COMP|47684-6|LNC|Leucine/Amino acids.total|Leucine/Amino acids.total
C1952919|T201|COMP|47685-3|LNC|Leucine/Amino acids.total|Leucine/Amino acids.total
C1952920|T201|COMP|47686-1|LNC|Linoleate/Creatinine|Linoleate/Creatinine
C1952924|T201|COMP|47689-5|LNC|Lysine|Lysine
C1952925|T201|COMP|47690-3|LNC|Lysine/Amino acids.total|Lysine/Amino acids.total
C1952927|T201|COMP|47691-1|LNC|Lysine/Amino acids.total|Lysine/Amino acids.total
C1952928|T201|COMP|47692-9|LNC|Lysine/Amino acids.total|Lysine/Amino acids.total
C1952929|T201|COMP|47693-7|LNC|Lysine/Amino acids.total|Lysine/Amino acids.total
C1952930|T201|COMP|47694-5|LNC|Lysine/Amino acids.total|Lysine/Amino acids.total
C1952931|T201|COMP|47695-2|LNC|Lysine/Amino acids.total|Lysine/Amino acids.total
C1952932|T201|COMP|47696-0|LNC|Malonate/Creatinine|Malonate/Creatinine
C1952934|T201|COMP|47697-8|LNC|Mandelate/Creatinine|Mandelate/Creatinine
C1952935|T201|COMP|47698-6|LNC|Mannitol/Creatinine|Mannitol/Creatinine
C1952937|T201|COMP|47699-4|LNC|Metanephrine/Creatinine|Metanephrine/Creatinine
C1952938|T201|COMP|47700-0|LNC|Methionine|Methionine
C1952939|T201|COMP|47701-8|LNC|Methionine/Amino acids.total|Methionine/Amino acids.total
C1952941|T201|COMP|47702-6|LNC|Methionine/Amino acids.total|Methionine/Amino acids.total
C1952942|T201|COMP|47703-4|LNC|Methionine/Amino acids.total|Methionine/Amino acids.total
C1952943|T201|COMP|47704-2|LNC|Methionine/Amino acids.total|Methionine/Amino acids.total
C1952944|T201|COMP|47705-9|LNC|Methionine/Amino acids.total|Methionine/Amino acids.total
C1952945|T201|COMP|47706-7|LNC|Methionine/Amino acids.total|Methionine/Amino acids.total
C1952946|T201|COMP|47707-5|LNC|Methylmalonate/Urea|Methylmalonate/Urea
C1952948|T201|COMP|47708-3|LNC|Methylmalonate/Urea|Methylmalonate/Urea
C1952949|T201|COMP|47709-1|LNC|Methylmalonate/Urea|Methylmalonate/Urea
C1952950|T201|COMP|47710-9|LNC|N-acetylaspartate/Creatinine|N-acetylaspartate/Creatinine
C1952951|T201|COMP|47711-7|LNC|Neopterin/Creatinine|Neopterin/Creatinine
C1952952|T201|COMP|47712-5|LNC|Nitrogen|Nitrogen
C1952953|T201|COMP|47713-3|LNC|Oleate/Creatinine|Oleate/Creatinine
C1952955|T201|COMP|47714-1|LNC|Ornithine|Ornithine
C1952956|T201|COMP|47715-8|LNC|Oxalate|Oxalate
C1952957|T201|COMP|47716-6|LNC|Oxygen^^adjusted to patient's actual temperature|Oxygen^^adjusted to patient's actual temperature
C1952958|T201|COMP|47717-4|LNC|Parathyrin^2H post dose calcium|Parathyrin^2H post dose calcium
C1952959|T201|COMP|47718-2|LNC|Parathyrin^4H post dose calcium|Parathyrin^4H post dose calcium
C1952960|T201|COMP|47719-0|LNC|Parathyrin^pre dose calcium|Parathyrin^pre dose calcium
C1952961|T201|COMP|47720-8|LNC|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1952962|T201|COMP|47721-6|LNC|Phenylalanine/Amino acids.total|Phenylalanine/Amino acids.total
C1952964|T201|COMP|47722-4|LNC|Phenylalanine/Amino acids.total|Phenylalanine/Amino acids.total
C1952965|T201|COMP|47723-2|LNC|Phenylalanine/Amino acids.total|Phenylalanine/Amino acids.total
C1952966|T201|COMP|47724-0|LNC|Phenylalanine/Amino acids.total|Phenylalanine/Amino acids.total
C1952967|T201|COMP|47725-7|LNC|Phenylalanine/Amino acids.total|Phenylalanine/Amino acids.total
C1952968|T201|COMP|47726-5|LNC|Phytanate/Creatinine|Phytanate/Creatinine
C1952970|T201|COMP|47727-3|LNC|Pipecolate/Creatinine|Pipecolate/Creatinine
C1952971|T201|COMP|47728-1|LNC|Procollagen type III/Creatinine|Procollagen type III/Creatinine
C1952973|T201|COMP|47729-9|LNC|Prolactin^1.5H post dose TRH IV|Prolactin^1.5H post dose TRH IV
C1952974|T201|COMP|47730-7|LNC|Prolactin^15M post dose TRH IV|Prolactin^15M post dose TRH IV
C1952975|T201|COMP|47731-5|LNC|Prolactin^2H post dose TRH IV|Prolactin^2H post dose TRH IV
C1952976|T201|COMP|47732-3|LNC|Proline|Proline
C1952977|T201|COMP|47733-1|LNC|Proline/Amino acids.total|Proline/Amino acids.total
C1952979|T201|COMP|47734-9|LNC|Proline/Amino acids.total|Proline/Amino acids.total
C1952980|T201|COMP|47735-6|LNC|Proline/Amino acids.total|Proline/Amino acids.total
C1952981|T201|COMP|47736-4|LNC|Proline/Amino acids.total|Proline/Amino acids.total
C1952982|T201|COMP|47737-2|LNC|Proline/Amino acids.total|Proline/Amino acids.total
C1952983|T201|COMP|47738-0|LNC|Prostate specific Ag|Prostate specific Ag
C1952984|T201|COMP|47739-8|LNC|Protein|Protein
C1952985|T201|COMP|47740-6|LNC|Purine nucleoside phosphorylase|Purine nucleoside phosphorylase
C1952986|T201|COMP|47741-4|LNC|Purine nucleoside phosphorylase|Purine nucleoside phosphorylase
C1952987|T201|COMP|47742-2|LNC|Serine|Serine
C1952988|T201|COMP|47743-0|LNC|Serine/Amino acids.total|Serine/Amino acids.total
C1952990|T201|COMP|47744-8|LNC|Serine/Amino acids.total|Serine/Amino acids.total
C1952991|T201|COMP|47745-5|LNC|Serine/Amino acids.total|Serine/Amino acids.total
C1952992|T201|COMP|47746-3|LNC|Serine/Amino acids.total|Serine/Amino acids.total
C1952993|T201|COMP|47747-1|LNC|Serine/Amino acids.total|Serine/Amino acids.total
C1952994|T201|COMP|47748-9|LNC|Serine/Amino acids.total|Serine/Amino acids.total
C1952995|T201|COMP|47749-7|LNC|Somatotropin^1.5H post dose glucagon|Somatotropin^1.5H post dose glucagon
C1952996|T201|COMP|47750-5|LNC|Somatotropin^1.5H post dose glucose PO|Somatotropin^1.5H post dose glucose PO
C1952997|T201|COMP|47751-3|LNC|Somatotropin^1.5H post dose TRH|Somatotropin^1.5H post dose TRH
C1952998|T201|COMP|47752-1|LNC|Somatotropin^1.5H post dose arginine|Somatotropin^1.5H post dose arginine
C1952999|T201|COMP|47753-9|LNC|Somatotropin^1.5H post dose insulin IV|Somatotropin^1.5H post dose insulin IV
C1953000|T201|COMP|47754-7|LNC|Somatotropin^10M post dose TRH|Somatotropin^10M post dose TRH
C1953001|T201|COMP|47755-4|LNC|Somatotropin^10th specimen post XXX challenge|Somatotropin^10th specimen post XXX challenge
C1953002|T201|COMP|47756-2|LNC|Somatotropin^15M pre dose arginine|Somatotropin^15M pre dose arginine
C1953003|T201|COMP|47757-0|LNC|Somatotropin^15M post dose arginine|Somatotropin^15M post dose arginine
C1953004|T201|COMP|47758-8|LNC|Somatotropin^15M post dose glucagon|Somatotropin^15M post dose glucagon
C1953005|T201|COMP|47759-6|LNC|Somatotropin^15M post dose insulin IV|Somatotropin^15M post dose insulin IV
C1953006|T201|COMP|47760-4|LNC|Somatotropin^1H post dose arginine|Somatotropin^1H post dose arginine
C1953007|T201|COMP|47761-2|LNC|Somatotropin^1H post dose glucose PO|Somatotropin^1H post dose glucose PO
C1953008|T201|COMP|47762-0|LNC|Somatotropin^1H post dose insulin IV|Somatotropin^1H post dose insulin IV
C1953009|T201|COMP|47763-8|LNC|Somatotropin^1st specimen post XXX challenge|Somatotropin^1st specimen post XXX challenge
C1953010|T201|COMP|48289-3|LNC|Sodium benzoate leukotriene release|Sodium benzoate leukotriene release
C1953012|T201|COMP|48290-1|LNC|Sodium nitrite leukotriene release|Sodium nitrite leukotriene release
C1953014|T201|COMP|48291-9|LNC|Potassium metabisulfite leukotriene release|Potassium metabisulfite leukotriene release
C1953016|T201|COMP|48292-7|LNC|Sodium salicylate leukotriene release|Sodium salicylate leukotriene release
C1953018|T201|COMP|48293-5|LNC|Tartrazine leukotriene release|Tartrazine leukotriene release
C1953020|T201|COMP|48294-3|LNC|Food colorant mix I leukotriene release|Food colorant mix I leukotriene release
C1953022|T201|COMP|48295-0|LNC|Food colorant mix II leukotriene release|Food colorant mix II leukotriene release
C1953024|T201|COMP|48296-8|LNC|Quinoline yellow leukotriene release|Quinoline yellow leukotriene release
C1953026|T201|COMP|48297-6|LNC|Chromotrope 2B leukotriene release|Chromotrope 2B leukotriene release
C1953028|T201|COMP|48371-9|LNC|Docosapentaenoate|Docosapentaenoate
C1953030|T201|COMP|48372-7|LNC|Spermatozoa.isolated head/100 spermatozoa|Spermatozoa.isolated head/100 spermatozoa
C1953032|T201|COMP|48373-5|LNC|Spermatozoa.angled midpiece/100 spermatozoa|Spermatozoa.angled midpiece/100 spermatozoa
C1953034|T201|COMP|48374-3|LNC|Spermatozoa.isolated tail/100 spermatozoa|Spermatozoa.isolated tail/100 spermatozoa
C1953036|T201|COMP|48375-0|LNC|Spermatozoa.short tail/100 spermatozoa|Spermatozoa.short tail/100 spermatozoa
C1953038|T201|COMP|48376-8|LNC|Collagen type 1 Ab|Collagen type 1 Ab
C1953039|T201|COMP|48377-6|LNC|Mullerian inhibiting substance|Mullerian inhibiting substance
C1953043|T201|COMP|48750-4|LNC|3-Hydroxy fatty acids pattern|3-Hydroxy fatty acids pattern
C1953045|T201|COMP|48751-2|LNC|3-Hydroxypalmitate.free|3-Hydroxypalmitate.free
C1953047|T201|COMP|48752-0|LNC|3-Hydroxymyristate.free|3-Hydroxymyristate.free
C1953049|T201|COMP|48753-8|LNC|3-Hydroxydodecanoate.free|3-Hydroxydodecanoate.free
C1953051|T201|COMP|48754-6|LNC|3-Hydroxydodecanoate|3-Hydroxydodecanoate
C1953052|T201|COMP|48755-3|LNC|3-Hydroxydecanoate.free|3-Hydroxydecanoate.free
C1953068|T201|COMP|47764-6|LNC|Somatotropin^2H post dose arginine|Somatotropin^2H post dose arginine
C1953069|T201|COMP|47765-3|LNC|Somatotropin^2H post dose glucose PO|Somatotropin^2H post dose glucose PO
C1953070|T201|COMP|47766-1|LNC|Somatotropin^2H post dose insulin IV|Somatotropin^2H post dose insulin IV
C1953071|T201|COMP|47767-9|LNC|Somatotropin^2nd specimen post XXX challenge|Somatotropin^2nd specimen post XXX challenge
C1953072|T201|COMP|47768-7|LNC|Somatotropin^30M post dose arginine|Somatotropin^30M post dose arginine
C1953073|T201|COMP|47769-5|LNC|Somatotropin^30M post dose glucose PO|Somatotropin^30M post dose glucose PO
C1953074|T201|COMP|47770-3|LNC|Somatotropin^30M post dose insulin IV|Somatotropin^30M post dose insulin IV
C1953075|T201|COMP|47771-1|LNC|Somatotropin^3H post dose glucose PO|Somatotropin^3H post dose glucose PO
C1953076|T201|COMP|47772-9|LNC|Somatotropin^45M post dose arginine|Somatotropin^45M post dose arginine
C1953077|T201|COMP|47773-7|LNC|Somatotropin^45M post dose insulin IV|Somatotropin^45M post dose insulin IV
C1953078|T201|COMP|47774-5|LNC|Somatotropin^pre dose arginine|Somatotropin^pre dose arginine
C1953079|T201|COMP|47775-2|LNC|Somatotropin^pre dose glucagon|Somatotropin^pre dose glucagon
C1953080|T201|COMP|47776-0|LNC|Somatotropin^pre dose glucose PO|Somatotropin^pre dose glucose PO
C1953081|T201|COMP|47777-8|LNC|Somatotropin^pre dose insulin IV|Somatotropin^pre dose insulin IV
C1953082|T201|COMP|47778-6|LNC|Somatotropin^pre dose TRH|Somatotropin^pre dose TRH
C1953083|T201|COMP|47779-4|LNC|Octadecanoate/Creatinine|Octadecanoate/Creatinine
C1953085|T201|COMP|47780-2|LNC|Sulfate|Sulfate
C1953086|T201|COMP|47781-0|LNC|Sulfocysteine|Sulfocysteine
C1953087|T201|COMP|47782-8|LNC|Taurine|Taurine
C1953088|T201|COMP|47783-6|LNC|Myristate/Creatinine|Myristate/Creatinine
C1953090|T201|COMP|47784-4|LNC|Threonine|Threonine
C1953091|T201|COMP|47785-1|LNC|Threonine/Amino acids.total|Threonine/Amino acids.total
C1953093|T201|COMP|47786-9|LNC|Threonine/Amino acids.total|Threonine/Amino acids.total
C1953094|T201|COMP|47787-7|LNC|Threonine/Amino acids.total|Threonine/Amino acids.total
C1953095|T201|COMP|47788-5|LNC|Threonine/Amino acids.total|Threonine/Amino acids.total
C1953096|T201|COMP|47789-3|LNC|Threonine/Amino acids.total|Threonine/Amino acids.total
C1953097|T201|COMP|47790-1|LNC|Threonine/Amino acids.total|Threonine/Amino acids.total
C1953098|T201|COMP|47791-9|LNC|Tocopherols|Tocopherols
C1953099|T201|COMP|47792-7|LNC|Tyrosine/Amino acids.total|Tyrosine/Amino acids.total
C1953101|T201|COMP|47793-5|LNC|Tyrosine/Amino acids.total|Tyrosine/Amino acids.total
C1953102|T201|COMP|47794-3|LNC|Tyrosine/Amino acids.total|Tyrosine/Amino acids.total
C1953103|T201|COMP|47795-0|LNC|Tyrosine/Amino acids.total|Tyrosine/Amino acids.total
C1953104|T201|COMP|47796-8|LNC|Tyrosine/Amino acids.total|Tyrosine/Amino acids.total
C1953105|T201|COMP|47797-6|LNC|Tyrosine/Amino acids.total|Tyrosine/Amino acids.total
C1953106|T201|COMP|47798-4|LNC|Urea|Urea
C1953107|T201|COMP|47799-2|LNC|Valine|Valine
C1953108|T201|COMP|47800-8|LNC|Valine/Amino acids.total|Valine/Amino acids.total
C1953110|T201|COMP|47801-6|LNC|Valine/Amino acids.total|Valine/Amino acids.total
C1953111|T201|COMP|47802-4|LNC|Valine/Amino acids.total|Valine/Amino acids.total
C1953112|T201|COMP|47803-2|LNC|Valine/Amino acids.total|Valine/Amino acids.total
C1953113|T201|COMP|47804-0|LNC|Valine/Amino acids.total|Valine/Amino acids.total
C1953114|T201|COMP|47805-7|LNC|Valine/Amino acids.total|Valine/Amino acids.total
C1953115|T201|COMP|47806-5|LNC|Xylose|Xylose
C1953116|T201|COMP|47807-3|LNC|2-Deoxytetronate/Creatinine|2-Deoxytetronate/Creatinine
C1953118|T201|COMP|47808-1|LNC|2-Ethylhydracrylate/Creatinine|2-Ethylhydracrylate/Creatinine
C1953120|T201|COMP|47809-9|LNC|2-Hydroxysebacate/Creatinine|2-Hydroxysebacate/Creatinine
C1953122|T201|COMP|47810-7|LNC|2-Methyl-3-Hydroxyvalerate|2-Methyl-3-Hydroxyvalerate
C1953123|T201|COMP|47811-5|LNC|2-Methyl-3-Oxobutyrate/Creatinine|2-Methyl-3-Oxobutyrate/Creatinine
C1953125|T201|COMP|47812-3|LNC|2-Methylglutaconate/Creatinine|2-Methylglutaconate/Creatinine
C1953127|T201|COMP|47813-1|LNC|2-Methylglutarate/Creatinine|2-Methylglutarate/Creatinine
C1953129|T201|COMP|47814-9|LNC|3,4-Dihydroxyphenyllactate/Creatinine|3,4-Dihydroxyphenyllactate/Creatinine
C1953131|T201|COMP|47815-6|LNC|3,4-Hydroxymandelate/Creatinine|3,4-Hydroxymandelate/Creatinine
C1953133|T201|COMP|47816-4|LNC|3-Deoxytetronate/Creatinine|3-Deoxytetronate/Creatinine
C1953135|T201|COMP|47817-2|LNC|3-Hydroxy,4-Methoxybenzoate/Creatinine|3-Hydroxy,4-Methoxybenzoate/Creatinine
C1953137|T201|COMP|47818-0|LNC|3-Hydroxyhexanoate/Creatinine|3-Hydroxyhexanoate/Creatinine
C1953139|T201|COMP|47819-8|LNC|3-Hydroxysuberate/Creatinine|3-Hydroxysuberate/Creatinine
C1953141|T201|COMP|47820-6|LNC|3-Hydroxyvalerate|3-Hydroxyvalerate
C1953142|T201|COMP|47821-4|LNC|3-Indolelactate/Creatinine|3-Indolelactate/Creatinine
C1953144|T201|COMP|47822-2|LNC|3-Methyladipate/Creatinine|3-Methyladipate/Creatinine
C1953146|T201|COMP|47823-0|LNC|4-Hydroxy-3-Methoxyphenyllactate/Creatinine|4-Hydroxy-3-Methoxyphenyllactate/Creatinine
C1953148|T201|COMP|47824-8|LNC|5-Hydroxycaproate/Creatinine|5-Hydroxycaproate/Creatinine
C1953150|T201|COMP|47825-5|LNC|7-Hydroxyoctanoate/Creatinine|7-Hydroxyoctanoate/Creatinine
C1953152|T201|COMP|47826-3|LNC|Adenosine deaminase|Adenosine deaminase
C1953153|T201|COMP|47827-1|LNC|Adenosyl homocysteine hydrolase|Adenosyl homocysteine hydrolase
C1953154|T201|COMP|47828-9|LNC|Adiponectin|Adiponectin
C1953155|T201|COMP|47829-7|LNC|Arabitol/Creatinine|Arabitol/Creatinine
C1953157|T201|COMP|47830-5|LNC|Argininosuccinate synthase|Argininosuccinate synthase
C1953158|T201|COMP|47831-3|LNC|Argininosuccinate synthase|Argininosuccinate synthase
C1953159|T201|COMP|47832-1|LNC|C peptide^4M post 1 mg glucagon|C peptide^4M post 1 mg glucagon
C1953160|T201|COMP|47833-9|LNC|C peptide^6M post dose glucagon|C peptide^6M post dose glucagon
C1953161|T201|COMP|47834-7|LNC|C peptide^8M post dose glucagon|C peptide^8M post dose glucagon
C1953162|T201|COMP|47835-4|LNC|Carnitine acyltransferase I|Carnitine acyltransferase I
C1953163|T201|COMP|47836-2|LNC|Carnitine acyltransferase I|Carnitine acyltransferase I
C1953164|T201|COMP|47837-0|LNC|Carnitine acyltransferase II|Carnitine acyltransferase II
C1953165|T201|COMP|47845-3|LNC|Cortisol^post 1 mg dexamethasone PO overnight|Cortisol^post 1 mg dexamethasone PO overnight
C1953170|T201|COMP|47850-3|LNC|Cortisol^post dose corticotropin|Cortisol^post dose corticotropin
C1953171|T201|COMP|47851-1|LNC|Cortisol^post dose dexamethasone|Cortisol^post dose dexamethasone
C1953172|T201|COMP|47852-9|LNC|Dehydroepiandrosterone^pre 250 ug corticotropin|Dehydroepiandrosterone^pre 250 ug corticotropin
C1953173|T201|COMP|47853-7|LNC|Diphosphoglycerate phosphatase|Diphosphoglycerate phosphatase
C1953174|T201|COMP|47854-5|LNC|Fibroblast growth factor 23.intact|Fibroblast growth factor 23.intact
C1953175|T201|COMP|47855-2|LNC|Fibroblast growth factor 23.C-terminal|Fibroblast growth factor 23.C-terminal
C1953177|T201|COMP|47857-8|LNC|Galactitol/Creatinine|Galactitol/Creatinine
C1953179|T201|COMP|47858-6|LNC|Gentisate/Creatinine|Gentisate/Creatinine
C1953181|T201|COMP|47859-4|LNC|Glucose^5M post dose glucose|Glucose^5M post dose glucose
C1953182|T201|COMP|47860-2|LNC|Glutamate dehydrogenase|Glutamate dehydrogenase
C1953183|T201|COMP|47861-0|LNC|Hypoxanthine phosphoribosyltransferase|Hypoxanthine phosphoribosyltransferase
C1953184|T201|COMP|47862-8|LNC|Insulin^post meal|Insulin^post meal
C1953185|T201|COMP|47863-6|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C1953187|T201|COMP|47865-1|LNC|Malondialdehyde|Malondialdehyde
C1953188|T201|COMP|47866-9|LNC|Phosphoribosylpyrophosphate synthetase|Phosphoribosylpyrophosphate synthetase
C1953189|T201|COMP|47867-7|LNC|Phosphoribosylpyrophosphate synthetase|Phosphoribosylpyrophosphate synthetase
C1953190|T201|COMP|47868-5|LNC|Prolactin^1.5H post dose metoclopramide|Prolactin^1.5H post dose metoclopramide
C1953191|T201|COMP|47869-3|LNC|Prolactin^1H post dose metoclopramide|Prolactin^1H post dose metoclopramide
C1953192|T201|COMP|47870-1|LNC|Prolactin^2.5H post dose TRH IV|Prolactin^2.5H post dose TRH IV
C1953193|T201|COMP|47871-9|LNC|Prolactin^30M post dose metoclopramide|Prolactin^30M post dose metoclopramide
C1953194|T201|COMP|47872-7|LNC|Prolactin^pre dose metoclopramide|Prolactin^pre dose metoclopramide
C1953195|T201|COMP|47873-5|LNC|Propionyl CO-A carboxylase|Propionyl CO-A carboxylase
C1953196|T201|COMP|47874-3|LNC|Propionyl CO-A carboxylase|Propionyl CO-A carboxylase
C1953197|T201|COMP|47875-0|LNC|Propionyl CO-A carboxylase|Propionyl CO-A carboxylase
C1953198|T201|COMP|47876-8|LNC|Propionyl CO-A carboxylase|Propionyl CO-A carboxylase
C1953199|T201|COMP|47877-6|LNC|Propionyl CO-A carboxylase|Propionyl CO-A carboxylase
C1953200|T201|COMP|47878-4|LNC|Propionylglycine|Propionylglycine
C1953201|T201|COMP|47879-2|LNC|Pyruvate carboxylase|Pyruvate carboxylase
C1953202|T201|COMP|47880-0|LNC|Pyruvate carboxylase|Pyruvate carboxylase
C1953203|T201|COMP|47881-8|LNC|Pyruvate carboxylase|Pyruvate carboxylase
C1953204|T201|COMP|47882-6|LNC|Pyruvate carboxylase|Pyruvate carboxylase
C1953205|T201|COMP|47883-4|LNC|Renin^upright|Renin^upright
C1953206|T201|COMP|47884-2|LNC|Ribitol/Creatinine|Ribitol/Creatinine
C1953208|T201|COMP|47885-9|LNC|Somatotropin^1.5H post dose arginine+insulin|Somatotropin^1.5H post dose arginine+insulin
C1953209|T201|COMP|47886-7|LNC|Somatotropin^1.5H post dose betaxolol+glucagon|Somatotropin^1.5H post dose betaxolol+glucagon
C1953210|T201|COMP|47887-5|LNC|Somatotropin^1.5H post dose ornithine|Somatotropin^1.5H post dose ornithine
C1953211|T201|COMP|47888-3|LNC|Somatotropin^1.75H post dose arginine+insulin|Somatotropin^1.75H post dose arginine+insulin
C1953212|T201|COMP|47889-1|LNC|Somatotropin^1.75H post dose ornithine|Somatotropin^1.75H post dose ornithine
C1953213|T201|COMP|47890-9|LNC|Somatotropin^15M post dose arginine+insulin|Somatotropin^15M post dose arginine+insulin
C1953215|T201|COMP|47892-5|LNC|Somatotropin^15M post dose ornithine|Somatotropin^15M post dose ornithine
C1953216|T201|COMP|47893-3|LNC|Somatotropin^1H post dose glucagon|Somatotropin^1H post dose glucagon
C1953218|T201|COMP|47895-8|LNC|Somatotropin^1H post dose ornithine|Somatotropin^1H post dose ornithine
C1953219|T201|COMP|47896-6|LNC|Somatotropin^1H post dose propranolol+glucagon|Somatotropin^1H post dose propranolol+glucagon
C1953220|T201|COMP|47897-4|LNC|Somatotropin^1H post dose TRH|Somatotropin^1H post dose TRH
C1953221|T201|COMP|47898-2|LNC|Somatotropin^2.25H post dose arginine+insulin|Somatotropin^2.25H post dose arginine+insulin
C1953222|T201|COMP|47899-0|LNC|Somatotropin^2.5H post dose propranolol+glucagon|Somatotropin^2.5H post dose propranolol+glucagon
C1953223|T201|COMP|47900-6|LNC|Somatotropin^20M post dose TRH|Somatotropin^20M post dose TRH
C1953224|T201|COMP|47901-4|LNC|Somatotropin^2H post dose arginine+insulin|Somatotropin^2H post dose arginine+insulin
C1953225|T201|COMP|47902-2|LNC|Somatotropin^2H post dose betaxolol+glucagon|Somatotropin^2H post dose betaxolol+glucagon
C1953226|T201|COMP|47903-0|LNC|Somatotropin^2H post dose glucagon|Somatotropin^2H post dose glucagon
C1953228|T201|COMP|47905-5|LNC|Somatotropin^2H post dose ornithine|Somatotropin^2H post dose ornithine
C1953229|T201|COMP|47906-3|LNC|Somatotropin^2H post dose propranolol+glucagon|Somatotropin^2H post dose propranolol+glucagon
C1953230|T201|COMP|47907-1|LNC|Somatotropin^2H post dose TRH|Somatotropin^2H post dose TRH
C1953231|T201|COMP|47908-9|LNC|Somatotropin^2H pre dose propranolol+glucagon|Somatotropin^2H pre dose propranolol+glucagon
C1953232|T201|COMP|47909-7|LNC|Somatotropin^30M post dose arginine+insulin|Somatotropin^30M post dose arginine+insulin
C1953233|T201|COMP|47910-5|LNC|Somatotropin^30M post dose betaxolol+glucagon|Somatotropin^30M post dose betaxolol+glucagon
C1953234|T201|COMP|47911-3|LNC|Somatotropin^30M post dose glucagon|Somatotropin^30M post dose glucagon
C1953236|T201|COMP|47913-9|LNC|Somatotropin^30M post dose ornithine|Somatotropin^30M post dose ornithine
C1953237|T201|COMP|47914-7|LNC|Somatotropin^30M post dose TRH|Somatotropin^30M post dose TRH
C1953238|T201|COMP|47915-4|LNC|Somatotropin^3H post dose betaxolol+glucagon|Somatotropin^3H post dose betaxolol+glucagon
C1953239|T201|COMP|47916-2|LNC|Somatotropin^3H post dose glucagon|Somatotropin^3H post dose glucagon
C1953240|T201|COMP|47917-0|LNC|Somatotropin^3H post dose propranolol+glucagon|Somatotropin^3H post dose propranolol+glucagon
C1953241|T201|COMP|47918-8|LNC|Somatotropin^3rd specimen post XXX challenge|Somatotropin^3rd specimen post XXX challenge
C1953242|T201|COMP|47919-6|LNC|Somatotropin^45M post dose arginine+insulin|Somatotropin^45M post dose arginine+insulin
C1953243|T201|COMP|47920-4|LNC|Somatotropin^45M post dose glucagon|Somatotropin^45M post dose glucagon
C1953245|T201|COMP|47922-0|LNC|Somatotropin^45M post dose ornithine|Somatotropin^45M post dose ornithine
C1953246|T201|COMP|47923-8|LNC|Somatotropin^4th specimen post XXX challenge|Somatotropin^4th specimen post XXX challenge
C1953247|T201|COMP|47924-6|LNC|Somatotropin^5M post dose arginine|Somatotropin^5M post dose arginine
C1953248|T201|COMP|47925-3|LNC|Somatotropin^5M post dose arginine+insulin|Somatotropin^5M post dose arginine+insulin
C1953249|T201|COMP|47926-1|LNC|Somatotropin^5M post dose ornithine|Somatotropin^5M post dose ornithine
C1953250|T201|COMP|47927-9|LNC|Somatotropin^5th specimen post XXX challenge|Somatotropin^5th specimen post XXX challenge
C1953251|T201|COMP|47928-7|LNC|Somatotropin^1H post dose betaxolol+glucagon|Somatotropin^1H post dose betaxolol+glucagon
C1953252|T201|COMP|47929-5|LNC|Somatotropin^6th specimen post XXX challenge|Somatotropin^6th specimen post XXX challenge
C1953253|T201|COMP|47930-3|LNC|Somatotropin^7th specimen post XXX challenge|Somatotropin^7th specimen post XXX challenge
C1953254|T201|COMP|47931-1|LNC|Somatotropin^8th specimen post XXX challenge|Somatotropin^8th specimen post XXX challenge
C1953255|T201|COMP|47932-9|LNC|Somatotropin^9th specimen post XXX challenge|Somatotropin^9th specimen post XXX challenge
C1953256|T201|COMP|47933-7|LNC|Somatotropin^pre dose arginine+insulin|Somatotropin^pre dose arginine+insulin
C1953257|T201|COMP|47934-5|LNC|Somatotropin^pre dose betaxolol+glucagon|Somatotropin^pre dose betaxolol+glucagon
C1953259|T201|COMP|47936-0|LNC|Somatotropin^pre dose ornithine|Somatotropin^pre dose ornithine
C1953260|T201|COMP|47937-8|LNC|Somatotropin^pre dose propranolol+glucagon|Somatotropin^pre dose propranolol+glucagon
C1953261|T201|COMP|47938-6|LNC|Specimen source|Specimen source
C1953262|T201|COMP|47939-4|LNC|Sulfocysteine|Sulfocysteine
C1953263|T201|COMP|47940-2|LNC|Testosterone^12H post 5000 U HCG IM|Testosterone^12H post 5000 U HCG IM
C1953264|T201|COMP|47941-0|LNC|Testosterone^1H post dose corticotropin|Testosterone^1H post dose corticotropin
C1953265|T201|COMP|47942-8|LNC|Testosterone^1D post 5000 U HCG IM|Testosterone^1D post 5000 U HCG IM
C1953266|T201|COMP|47943-6|LNC|Testosterone^2D post 5000 U HCG IM|Testosterone^2D post 5000 U HCG IM
C1953267|T201|COMP|47944-4|LNC|Testosterone^4H post 5000 U HCG IM|Testosterone^4H post 5000 U HCG IM
C1953268|T201|COMP|47945-1|LNC|Testosterone^3D post 5000 U HCG IM|Testosterone^3D post 5000 U HCG IM
C1953269|T201|COMP|47946-9|LNC|Testosterone^pre dose corticotropin|Testosterone^pre dose corticotropin
C1953277|T201|COMP|47954-3|LNC|Tiglylglycine|Tiglylglycine
C1953278|T201|COMP|47955-0|LNC|EYA1 gene targeted mutation analysis|EYA1 gene targeted mutation analysis
C1953280|T201|COMP|47956-8|LNC|CNR1 gene targeted mutation analysis|CNR1 gene targeted mutation analysis
C1953282|T201|COMP|47957-6|LNC|Deoxyuridine|Deoxyuridine
C1953283|T201|COMP|47958-4|LNC|FLT3 gene targeted mutation analysis|FLT3 gene targeted mutation analysis
C1953285|T201|COMP|47959-2|LNC|GFAP gene targeted mutation analysis|GFAP gene targeted mutation analysis
C1953287|T201|COMP|47960-0|LNC|GLRA1 gene targeted mutation analysis|GLRA1 gene targeted mutation analysis
C1953289|T201|COMP|47961-8|LNC|ACVRL1 gene targeted mutation analysis|ACVRL1 gene targeted mutation analysis
C1953291|T201|COMP|47962-6|LNC|JAG1 gene targeted mutation analysis|JAG1 gene targeted mutation analysis
C1953293|T201|COMP|47963-4|LNC|JAK3 gene targeted mutation analysis|JAK3 gene targeted mutation analysis
C1953295|T201|COMP|47964-2|LNC|MVK gene targeted mutation analysis|MVK gene targeted mutation analysis
C1953297|T201|COMP|47965-9|LNC|Mycoplasma penetrans DNA|Mycoplasma penetrans DNA
C1953298|T201|COMP|47966-7|LNC|NCF2 gene targeted mutation analysis|NCF2 gene targeted mutation analysis
C1953300|T201|COMP|47967-5|LNC|NSD1 gene targeted mutation analysis|NSD1 gene targeted mutation analysis
C1953302|T201|COMP|47968-3|LNC|PINK1 gene targeted mutation analysis|PINK1 gene targeted mutation analysis
C1953304|T201|COMP|47969-1|LNC|PTEN gene targeted mutation analysis|PTEN gene targeted mutation analysis
C1953306|T201|COMP|47970-9|LNC|SGCB gene targeted mutation analysis|SGCB gene targeted mutation analysis
C1953308|T201|COMP|47971-7|LNC|SGSH gene targeted mutation analysis|SGSH gene targeted mutation analysis
C1953310|T201|COMP|47972-5|LNC|TGFBR1 gene targeted mutation analysis|TGFBR1 gene targeted mutation analysis
C1953312|T201|COMP|47973-3|LNC|TGFBR2 gene targeted mutation analysis|TGFBR2 gene targeted mutation analysis
C1953314|T201|COMP|47974-1|LNC|THRB gene targeted mutation analysis|THRB gene targeted mutation analysis
C1953316|T201|COMP|47975-8|LNC|tiZANidine|tiZANidine
C1953317|T201|COMP|47976-6|LNC|Selenium|Selenium
C1953318|T201|COMP|47977-4|LNC|Smooth muscle Ab.IgG|Smooth muscle Ab.IgG
C1953319|T201|COMP|47978-2|LNC|17-Ketosteroids|17-Ketosteroids
C1953320|T201|COMP|47979-0|LNC|Tranylcypromine|Tranylcypromine
C1953321|T201|COMP|47980-8|LNC|Mirtazapine|Mirtazapine
C1953322|T201|COMP|47981-6|LNC|Phenylalanine/Creatinine|Phenylalanine/Creatinine
C1953323|T201|COMP|47982-4|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1953329|T201|COMP|47988-1|LNC|Progesterone^6th specimen post XXX challenge|Progesterone^6th specimen post XXX challenge
C1953330|T201|COMP|47989-9|LNC|Progesterone^7th specimen post XXX challenge|Progesterone^7th specimen post XXX challenge
C1953331|T201|COMP|47990-7|LNC|Progesterone^8th specimen post XXX challenge|Progesterone^8th specimen post XXX challenge
C1953332|T201|COMP|47991-5|LNC|Progesterone^9th specimen post XXX challenge|Progesterone^9th specimen post XXX challenge
C1953333|T201|COMP|47994-9|LNC|Bilirubin|Bilirubin
C1953334|T201|COMP|47995-6|LNC|Glucose|Glucose
C1953335|T201|COMP|47996-4|LNC|Adenosine deaminase binding protein|Adenosine deaminase binding protein
C1953336|T201|COMP|47997-2|LNC|Genetic variant clinical significance|Genetic variant clinical significance
C1953338|T201|COMP|47998-0|LNC|DNA sequence variation display name|DNA sequence variation display name
C1953340|T201|COMP|47999-8|LNC|DNA region name|DNA region name
C1953342|T201|COMP|48000-4|LNC|Chromosome|Chromosome
C1953344|T201|COMP|48001-2|LNC|Chromosome region|Chromosome region
C1953346|T201|COMP|48002-0|LNC|Genomic source class|Genomic source class
C1953348|T201|COMP|48003-8|LNC|DNA sequence variation identifier|DNA sequence variation identifier
C1953350|T201|COMP|48004-6|LNC|DNA change|DNA change
C1953352|T201|COMP|48005-3|LNC|Amino acid change|Amino acid change
C1953354|T201|COMP|48006-1|LNC|Amino acid change type|Amino acid change type
C1953356|T201|COMP|48007-9|LNC|Genetic variant allelic state|Genetic variant allelic state
C1953358|T201|COMP|48008-7|LNC|Allele name|Allele name
C1953360|T201|COMP|48009-5|LNC|Genechip manufacturer ID|Genechip manufacturer ID
C1953362|T201|COMP|48010-3|LNC|Genechip ID|Genechip ID
C1953364|T201|COMP|48011-1|LNC|Genechip version|Genechip version
C1953366|T201|COMP|48012-9|LNC|Reference sequence|Reference sequence
C1953368|T201|COMP|48013-7|LNC|Genomic reference sequence identifier|Genomic reference sequence identifier
C1953370|T201|COMP|48014-5|LNC|Sequence variation panel|Sequence variation panel
C1953372|T201|COMP|48015-2|LNC|Individual allele panel|Individual allele panel
C1953374|T201|COMP|48016-0|LNC|Genechip kit panel|Genechip kit panel
C1953376|T201|COMP|48017-8|LNC|Sequencing methodology panel|Sequencing methodology panel
C1953378|T201|COMP|48018-6|LNC|Gene identifier|Gene identifier
C1953379|T201|COMP|48019-4|LNC|DNA change type|DNA change type
C1953381|T201|COMP|48020-2|LNC|Forward primer|Forward primer
C1953383|T201|COMP|48021-0|LNC|Reverse primer|Reverse primer
C1953387|T201|COMP|48023-6|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C1953389|T201|COMP|48024-4|LNC|AS gene targeted mutation analysis|AS gene targeted mutation analysis
C1953391|T201|COMP|48025-1|LNC|Gene mutations tested for|Gene mutations tested for
C1953392|T201|COMP|48026-9|LNC|ITGA2B gene targeted mutation analysis|ITGA2B gene targeted mutation analysis
C1953394|T201|COMP|48027-7|LNC|MT-ND4 gene.c.G15257A|MT-ND4 gene.c.G15257A
C1953396|T201|COMP|48028-5|LNC|SERPINE1 gene targeted mutation analysis|SERPINE1 gene targeted mutation analysis
C1953398|T201|COMP|48029-3|LNC|PKLR gene targeted mutation analysis|PKLR gene targeted mutation analysis
C1953400|T201|COMP|48030-1|LNC|RHE gene targeted mutation analysis|RHE gene targeted mutation analysis
C1953402|T201|COMP|48031-9|LNC|SCA10 gene.CAG repeats|SCA10 gene.CAG repeats
C1953404|T201|COMP|48032-7|LNC|THRB gene.p.Ala317Thr|THRB gene.p.Ala317Thr
C1953406|T201|COMP|48033-5|LNC|TTR gene targeted mutation analysis|TTR gene targeted mutation analysis
C1953408|T201|COMP|48034-3|LNC|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C1953409|T201|COMP|48035-0|LNC|Hemoglobin|Hemoglobin
C1953410|T201|COMP|48036-8|LNC|Glucose|Glucose
C1953412|T201|COMP|48038-4|LNC|Pathologist interpretation|Pathologist interpretation
C1953413|T201|COMP|48039-2|LNC|Fibronectin.fetal|Fibronectin.fetal
C1953414|T201|COMP|48040-0|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C1953415|T201|COMP|48041-8|LNC|Anthraquinone cutoff|Anthraquinone cutoff
C1953417|T201|COMP|48042-6|LNC|Bisacodyl cutoff|Bisacodyl cutoff
C1953419|T201|COMP|48043-4|LNC|Oxyphenisatin cutoff|Oxyphenisatin cutoff
C1953421|T201|COMP|48044-2|LNC|Phenolphthalein cutoff|Phenolphthalein cutoff
C1953423|T201|COMP|48045-9|LNC|Magnesium cutoff|Magnesium cutoff
C1953425|T201|COMP|48046-7|LNC|Phosphate cutoff|Phosphate cutoff
C1953427|T201|COMP|48047-5|LNC|Hemoglobin.gastrointestinal|Hemoglobin.gastrointestinal
C1953428|T201|COMP|48048-3|LNC|Neutrophils|Neutrophils
C1953429|T201|COMP|48049-1|LNC|Eosinophils|Eosinophils
C1953430|T201|COMP|48050-9|LNC|Neutrophils|Neutrophils
C1953431|T201|COMP|48051-7|LNC|Erythrocytes|Erythrocytes
C1953432|T201|COMP|48052-5|LNC|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C1953433|T201|COMP|48053-3|LNC|Turbidity|Turbidity
C1953434|T201|COMP|48054-1|LNC|Coagulation kaolin induced|Coagulation kaolin induced
C1953435|T201|COMP|48055-8|LNC|Pneumocystis jiroveci|Pneumocystis jiroveci
C1953436|T201|COMP|48056-6|LNC|Human bocavirus Ag|Human bocavirus Ag
C1953438|T201|COMP|48057-4|LNC|Human bocavirus Ab.IgG|Human bocavirus Ab.IgG
C1953440|T201|COMP|48058-2|LNC|Fibrin D-dimer DDU|Fibrin D-dimer DDU
C1953441|T201|COMP|48059-0|LNC|Giardia lamblia+Cryptosporidium sp Ag|Giardia lamblia+Cryptosporidium sp Ag
C1953443|T201|COMP|48060-8|LNC|Giardia lamblia+Cryptosporidium sp Ag|Giardia lamblia+Cryptosporidium sp Ag
C1953444|T201|COMP|48061-6|LNC|Giardia lamblia+Cryptosporidium sp Ag|Giardia lamblia+Cryptosporidium sp Ag
C1953445|T201|COMP|48062-4|LNC|Giardia lamblia+Cryptosporidium parvum Ag|Giardia lamblia+Cryptosporidium parvum Ag
C1953447|T201|COMP|48063-2|LNC|Giardia lamblia+Cryptosporidium parvum Ag|Giardia lamblia+Cryptosporidium parvum Ag
C1953448|T201|COMP|48064-0|LNC|Giardia lamblia+Cryptosporidium parvum Ag|Giardia lamblia+Cryptosporidium parvum Ag
C1953449|T201|COMP|48065-7|LNC|Fibrin D-dimer FEU|Fibrin D-dimer FEU
C1953451|T201|COMP|48066-5|LNC|Fibrin D-dimer DDU|Fibrin D-dimer DDU
C1953452|T201|COMP|48067-3|LNC|Fibrin D-dimer FEU|Fibrin D-dimer FEU
C1953453|T201|COMP|48068-1|LNC|Heinz bodies|Heinz bodies
C1953454|T201|COMP|48069-9|LNC|Spherocytes.micro|Spherocytes.micro
C1953456|T201|COMP|48070-7|LNC|Hepatitis B virus surface Ab.IgG|Hepatitis B virus surface Ab.IgG
C1953458|T201|COMP|48071-5|LNC|Complement total hemolytic CH50|Complement total hemolytic CH50
C1953459|T201|COMP|48072-3|LNC|Synthetic glucocorticoid drug|Synthetic glucocorticoid drug
C1953461|T201|COMP|48073-1|LNC|Thyroxine binding globulin panel|Thyroxine binding globulin panel
C1953463|T201|COMP|48074-9|LNC|Somatotropin^2.5H post dose arginine+insulin|Somatotropin^2.5H post dose arginine+insulin
C1953464|T201|COMP|48075-6|LNC|Somatotropin^2.5H post dose betaxolol+glucagon|Somatotropin^2.5H post dose betaxolol+glucagon
C1953465|T201|COMP|48076-4|LNC|Somatotropin^2.5H post dose glucagon|Somatotropin^2.5H post dose glucagon
C1953467|T201|COMP|48078-0|LNC|3,6-Epoxydecanedioate/Creatinine|3,6-Epoxydecanedioate/Creatinine
C1953469|T201|COMP|48079-8|LNC|3,6-Epoxydodecanedioate/Creatinine|3,6-Epoxydodecanedioate/Creatinine
C1953471|T201|COMP|48080-6|LNC|3,6-Epoxyoctanedioate/Creatinine|3,6-Epoxyoctanedioate/Creatinine
C1953473|T201|COMP|48081-4|LNC|3,6-Epoxytetradecanedioate/Creatinine|3,6-Epoxytetradecanedioate/Creatinine
C1953475|T201|COMP|48082-2|LNC|3-Hydroxyadipate 3,6-lactone/Creatinine|3-Hydroxyadipate 3,6-lactone/Creatinine
C1953477|T201|COMP|48083-0|LNC|3-Hydroxydodecanedienedioate/Creatinine|3-Hydroxydodecanedienedioate/Creatinine
C1953479|T201|COMP|48084-8|LNC|3-Hydroxydodecanedioate/Creatinine|3-Hydroxydodecanedioate/Creatinine
C1953480|T201|COMP|48085-5|LNC|3-Hydroxydodecenedioate/Creatinine|3-Hydroxydodecenedioate/Creatinine
C1953482|T201|COMP|48086-3|LNC|3-Hydroxytetradecadienedioate/Creatinine|3-Hydroxytetradecadienedioate/Creatinine
C1953484|T201|COMP|48087-1|LNC|3-Hydroxytetradecanedioate/Creatinine|3-Hydroxytetradecanedioate/Creatinine
C1953486|T201|COMP|48088-9|LNC|3-Hydroxytetradecenedioate/Creatinine|3-Hydroxytetradecenedioate/Creatinine
C1953488|T201|COMP|48089-7|LNC|Cholesterol/Apolipoprotein B|Cholesterol/Apolipoprotein B
C1953492|T201|COMP|48091-3|LNC|Corticotropin^12 AM specimen|Corticotropin^12 AM specimen
C1953493|T201|COMP|48092-1|LNC|Corticotropin^12 PM specimen|Corticotropin^12 PM specimen
C1953494|T201|COMP|48093-9|LNC|Corticotropin^15M pre 1 ug/kg CRH IV|Corticotropin^15M pre 1 ug/kg CRH IV
C1953495|T201|COMP|48094-7|LNC|Corticotropin^4 AM specimen|Corticotropin^4 AM specimen
C1953496|T201|COMP|48095-4|LNC|Corticotropin^4 PM specimen|Corticotropin^4 PM specimen
C1953497|T201|COMP|48096-2|LNC|Corticotropin^8 AM specimen|Corticotropin^8 AM specimen
C1953498|T201|COMP|48097-0|LNC|Corticotropin^8 PM specimen|Corticotropin^8 PM specimen
C1953499|T201|COMP|48098-8|LNC|Cortisol^12 AM specimen|Cortisol^12 AM specimen
C1953500|T201|COMP|48099-6|LNC|Cortisol^12 PM specimen|Cortisol^12 PM specimen
C1953501|T201|COMP|48100-2|LNC|Cortisol^15M pre 1 ug/kg CRH IV|Cortisol^15M pre 1 ug/kg CRH IV
C1953502|T201|COMP|48101-0|LNC|Cortisol^15M pre 1 ug/kg CRH IV|Cortisol^15M pre 1 ug/kg CRH IV
C1953503|T201|COMP|48102-8|LNC|Cortisol^4 AM specimen|Cortisol^4 AM specimen
C1953504|T201|COMP|48103-6|LNC|Cortisol^4 AM specimen|Cortisol^4 AM specimen
C1953505|T201|COMP|48104-4|LNC|Cortisol^8 AM specimen|Cortisol^8 AM specimen
C1953506|T201|COMP|48105-1|LNC|Cortisol^8 PM specimen|Cortisol^8 PM specimen
C1953507|T201|COMP|48106-9|LNC|4,5-Dihydroxyhexanolactone/Creatinine|4,5-Dihydroxyhexanolactone/Creatinine
C1953509|T201|COMP|48107-7|LNC|Erythritol/Creatinine|Erythritol/Creatinine
C1953512|T201|COMP|48109-3|LNC|Glucose^15M pre dose glucose|Glucose^15M pre dose glucose
C1953513|T201|COMP|48110-1|LNC|Glutathione.oxidized/glutathione.reduced|Glutathione.oxidized/glutathione.reduced
C1953515|T201|COMP|48111-9|LNC|Glutathione.reduced|Glutathione.reduced
C1953516|T201|COMP|48112-7|LNC|Glutathione.reduced|Glutathione.reduced
C1953517|T201|COMP|48113-5|LNC|Heptadecenoate/Creatinine|Heptadecenoate/Creatinine
C1953519|T201|COMP|48114-3|LNC|Hexadecanedioate/Creatinine|Hexadecanedioate/Creatinine
C1953521|T201|COMP|48115-0|LNC|Homocysteine.free/Creatinine|Homocysteine.free/Creatinine
C1953523|T201|COMP|48116-8|LNC|Insulin^10M pre dose glucose|Insulin^10M pre dose glucose
C1953524|T201|COMP|48117-6|LNC|Isovalerylglycine/Urea|Isovalerylglycine/Urea
C1953527|T201|COMP|48138-2|LNC|Enolase.neuron specific|Enolase.neuron specific
C1953528|T201|COMP|48139-0|LNC|Erythro-4,5-Dihydroxyhexanoate/Creatinine|Erythro-4,5-Dihydroxyhexanoate/Creatinine
C1953530|T201|COMP|48140-8|LNC|Erythro-4-Deoxytetronate/Creatinine|Erythro-4-Deoxytetronate/Creatinine
C1953532|T201|COMP|48141-6|LNC|Ferritin|Ferritin
C1953533|T201|COMP|48142-4|LNC|Indole-3-Acetate/Creatinine|Indole-3-Acetate/Creatinine
C1953535|T201|COMP|48143-2|LNC|LDL.oxidized Ab|LDL.oxidized Ab
C1953537|T201|COMP|48144-0|LNC|Mannose|Mannose
C1953538|T201|COMP|48145-7|LNC|Mevalonolactone/Creatinine|Mevalonolactone/Creatinine
C1953540|T201|COMP|48146-5|LNC|Myeloperoxidase|Myeloperoxidase
C1953541|T201|COMP|48147-3|LNC|Oligosaccharides/Creatinine|Oligosaccharides/Creatinine
C1953543|T201|COMP|48148-1|LNC|Osmolality|Osmolality
C1953544|T201|COMP|48149-9|LNC|Osmolality.urine/Osmolality.ser|Osmolality.urine/Osmolality.ser
C1953546|T201|COMP|48150-7|LNC|Perseitol/Creatinine|Perseitol/Creatinine
C1953548|T201|COMP|48151-5|LNC|Sedoheptitol/Creatinine|Sedoheptitol/Creatinine
C1953550|T201|COMP|48152-3|LNC|Sorbitol/Creatinine|Sorbitol/Creatinine
C1953552|T201|COMP|48153-1|LNC|Threitol/Creatinine|Threitol/Creatinine
C1953554|T201|COMP|48154-9|LNC|Threo-4,5-Dihydrohexanoate/Creatinine|Threo-4,5-Dihydrohexanoate/Creatinine
C1953556|T201|COMP|48155-6|LNC|Threo-4,5-Dihydrohexanolactone/Creatinine|Threo-4,5-Dihydrohexanolactone/Creatinine
C1953558|T201|COMP|48156-4|LNC|Threo-4-Deoxytetronate/Creatinine|Threo-4-Deoxytetronate/Creatinine
C1953560|T201|COMP|48157-2|LNC|Thymine/Creatinine|Thymine/Creatinine
C1953562|T201|COMP|48158-0|LNC|Vanillate/Creatinine|Vanillate/Creatinine
C1953564|T201|COMP|48159-8|LNC|Hepatitis C virus Ab Signal/Cutoff|Hepatitis C virus Ab Signal/Cutoff
C1953566|T201|COMP|48160-6|LNC|HTLV I rgp21 Ab|HTLV I rgp21 Ab
C1953567|T201|COMP|48161-4|LNC|PROS1 gene targeted mutation analysis|PROS1 gene targeted mutation analysis
C1953569|T201|COMP|48162-2|LNC|Thymidine|Thymidine
C1953570|T201|COMP|48163-0|LNC|Cytokeratin 19|Cytokeratin 19
C1953571|T201|COMP|48164-8|LNC|Enolase.neuron specific|Enolase.neuron specific
C1953572|T201|COMP|48165-5|LNC|Squamous cell carcinoma Ag|Squamous cell carcinoma Ag
C1953573|T201|COMP|48166-3|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C1953574|T201|COMP|48167-1|LNC|Prostate specific Ag/Creatinine|Prostate specific Ag/Creatinine
C1953576|T201|COMP|48168-9|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C1953577|T201|COMP|48169-7|LNC|Amikacin 1.5 ug/mL|Amikacin 1.5 ug/mL
C1953579|T201|COMP|48170-5|LNC|Capreomycin 3.0 ug/mL|Capreomycin 3.0 ug/mL
C1953581|T201|COMP|48171-3|LNC|Isoniazid 0.1 ug/mL|Isoniazid 0.1 ug/mL
C1953582|T201|COMP|48172-1|LNC|Isoniazid 0.4 ug/mL|Isoniazid 0.4 ug/mL
C1953583|T201|COMP|48173-9|LNC|levoFLOXacin 1.5 ug/mL|levoFLOXacin 1.5 ug/mL
C1953585|T201|COMP|48174-7|LNC|Mycobacterium tuberculosis complex rRNA|Mycobacterium tuberculosis complex rRNA
C1953589|T201|COMP|48177-0|LNC|Streptomycin 1.0 ug/mL|Streptomycin 1.0 ug/mL
C1953591|T201|COMP|48178-8|LNC|Reference change value 0.99|Reference change value 0.99
C1953593|T201|COMP|48179-6|LNC|Reference change value 0.99|Reference change value 0.99
C1953594|T201|COMP|48180-4|LNC|Reference change value 0.95|Reference change value 0.95
C1953596|T201|COMP|48181-2|LNC|Reference change value 0.95|Reference change value 0.95
C1953597|T201|COMP|48182-0|LNC|Vespa crabro leukotriene release|Vespa crabro leukotriene release
C1953599|T201|COMP|48183-8|LNC|Polistes spp leukotriene release|Polistes spp leukotriene release
C1953601|T201|COMP|48184-6|LNC|Vespula spp leukotriene release|Vespula spp leukotriene release
C1953603|T201|COMP|48185-3|LNC|Apis mellifera leukotriene release|Apis mellifera leukotriene release
C1953605|T201|COMP|48186-1|LNC|Amylase leukotriene release|Amylase leukotriene release
C1953607|T201|COMP|48187-9|LNC|Chloramin T leukotriene release|Chloramin T leukotriene release
C1953609|T201|COMP|48188-7|LNC|Latex leukotriene release|Latex leukotriene release
C1953611|T201|COMP|48189-5|LNC|Formaldehyde leukotriene release|Formaldehyde leukotriene release
C1953613|T201|COMP|48190-3|LNC|Phthalic anhydride leukotriene release|Phthalic anhydride leukotriene release
C1953615|T201|COMP|48191-1|LNC|Monosodium glutamate leukotriene release|Monosodium glutamate leukotriene release
C1953617|T201|COMP|48192-9|LNC|Sunset yellow FCF leukotriene release|Sunset yellow FCF leukotriene release
C1953619|T201|COMP|48193-7|LNC|Succinylcholine leukotriene release|Succinylcholine leukotriene release
C1953621|T201|COMP|48194-5|LNC|Lidocaine leukotriene release|Lidocaine leukotriene release
C1953623|T201|COMP|48195-2|LNC|Trimethoprim leukotriene release|Trimethoprim leukotriene release
C1953625|T201|COMP|48196-0|LNC|Cephalosporin C leukotriene release|Cephalosporin C leukotriene release
C1953627|T201|COMP|48197-8|LNC|Cefuroxime leukotriene release|Cefuroxime leukotriene release
C1953629|T201|COMP|48198-6|LNC|Amoxicillin leukotriene release|Amoxicillin leukotriene release
C1953631|T201|COMP|48206-7|LNC|Lactalbumin alpha leukotriene release|Lactalbumin alpha leukotriene release
C1953633|T201|COMP|48207-5|LNC|Egg yolk leukotriene release|Egg yolk leukotriene release
C1953635|T201|COMP|48208-3|LNC|Saccharomyces cerevisiae leukotriene release|Saccharomyces cerevisiae leukotriene release
C1953637|T201|COMP|48209-1|LNC|Citrus sinensis leukotriene release|Citrus sinensis leukotriene release
C1953639|T201|COMP|48210-9|LNC|Daucus carota leukotriene release|Daucus carota leukotriene release
C1953641|T201|COMP|48211-7|LNC|Beef leukotriene release|Beef leukotriene release
C1953643|T201|COMP|48212-5|LNC|Pork leukotriene release|Pork leukotriene release
C1953645|T201|COMP|48213-3|LNC|Lycopersicon lycopersicum leukotriene release|Lycopersicon lycopersicum leukotriene release
C1953647|T201|COMP|48214-1|LNC|Pandalus borealis leukotriene release|Pandalus borealis leukotriene release
C1953649|T201|COMP|48215-8|LNC|Cancer pagurus leukotriene release|Cancer pagurus leukotriene release
C1953651|T201|COMP|48216-6|LNC|Corylus avellana leukotriene release|Corylus avellana leukotriene release
C1953653|T201|COMP|48217-4|LNC|Glycine max leukotriene release|Glycine max leukotriene release
C1953655|T201|COMP|48218-2|LNC|Arachis hypogaea leukotriene release|Arachis hypogaea leukotriene release
C1953657|T201|COMP|48219-0|LNC|Sesamum indicum leukotriene release|Sesamum indicum leukotriene release
C1953659|T201|COMP|48220-8|LNC|Avena sativa leukotriene release|Avena sativa leukotriene release
C1953661|T201|COMP|48221-6|LNC|Hordeum vulgare leukotriene release|Hordeum vulgare leukotriene release
C1953663|T201|COMP|48222-4|LNC|Secale cereale leukotriene release|Secale cereale leukotriene release
C1953665|T201|COMP|48223-2|LNC|Triticum aestivum leukotriene release|Triticum aestivum leukotriene release
C1953667|T201|COMP|48224-0|LNC|Gadus morhua leukotriene release|Gadus morhua leukotriene release
C1953669|T201|COMP|48225-7|LNC|Cow milk leukotriene release|Cow milk leukotriene release
C1953671|T201|COMP|48226-5|LNC|Egg white leukotriene release|Egg white leukotriene release
C1953673|T201|COMP|48227-3|LNC|Human serum albumin leukotriene release|Human serum albumin leukotriene release
C1953675|T201|COMP|48228-1|LNC|Bovine serum albumin leukotriene release|Bovine serum albumin leukotriene release
C1953677|T201|COMP|48229-9|LNC|Dog epithelium leukotriene release|Dog epithelium leukotriene release
C1953679|T201|COMP|48230-7|LNC|Cat dander leukotriene release|Cat dander leukotriene release
C1953681|T201|COMP|48231-5|LNC|Glycyphagus domesticus leukotriene release|Glycyphagus domesticus leukotriene release
C1953683|T201|COMP|48232-3|LNC|Tyrophagus putrescentiae leukotriene release|Tyrophagus putrescentiae leukotriene release
C1953685|T201|COMP|48233-1|LNC|Lepidoglyphus destructor leukotriene release|Lepidoglyphus destructor leukotriene release
C1953687|T201|COMP|48234-9|LNC|Acarus siro leukotriene release|Acarus siro leukotriene release
C1953689|T201|COMP|48235-6|LNC|Dermatophagoides farinae leukotriene release|Dermatophagoides farinae leukotriene release
C1953693|T201|COMP|48237-2|LNC|Ctenocephalides sp leukotriene release|Ctenocephalides sp leukotriene release
C1953695|T201|COMP|48238-0|LNC|Blatella germanica leukotriene release|Blatella germanica leukotriene release
C1953697|T201|COMP|48239-8|LNC|Alternaria alternata leukotriene release|Alternaria alternata leukotriene release
C1953699|T201|COMP|48240-6|LNC|Candida albicans leukotriene release|Candida albicans leukotriene release
C1953701|T201|COMP|48241-4|LNC|Aspergillus fumigatus leukotriene release|Aspergillus fumigatus leukotriene release
C1953703|T201|COMP|48242-2|LNC|Cladosporium herbarum leukotriene release|Cladosporium herbarum leukotriene release
C1953705|T201|COMP|48243-0|LNC|Penicillium notatum leukotriene release|Penicillium notatum leukotriene release
C1953707|T201|COMP|48244-8|LNC|Juniperus virginiana leukotriene release|Juniperus virginiana leukotriene release
C1953709|T201|COMP|48245-5|LNC|Cryptomeria japonica leukotriene release|Cryptomeria japonica leukotriene release
C1953711|T201|COMP|48246-3|LNC|Olea europaea pollen leukotriene release|Olea europaea pollen leukotriene release
C1953713|T201|COMP|48247-1|LNC|Quercus alba leukotriene release|Quercus alba leukotriene release
C1953715|T201|COMP|48248-9|LNC|Corylus avellana pollen leukotriene release|Corylus avellana pollen leukotriene release
C1953717|T201|COMP|48249-7|LNC|Betula verrucosa leukotriene release|Betula verrucosa leukotriene release
C1953719|T201|COMP|48250-5|LNC|Parietaria judaica leukotriene release|Parietaria judaica leukotriene release
C1953721|T201|COMP|48251-3|LNC|Parietaria officinalis leukotriene release|Parietaria officinalis leukotriene release
C1953723|T201|COMP|48252-1|LNC|Salsola kali leukotriene release|Salsola kali leukotriene release
C1953725|T201|COMP|48253-9|LNC|Plantago lanceolata leukotriene release|Plantago lanceolata leukotriene release
C1953727|T201|COMP|48254-7|LNC|Artemisia vulgaris leukotriene release|Artemisia vulgaris leukotriene release
C1953729|T201|COMP|48255-4|LNC|Ambrosia trifida leukotriene release|Ambrosia trifida leukotriene release
C1953731|T201|COMP|48256-2|LNC|Ambrosia elatior leukotriene release|Ambrosia elatior leukotriene release
C1953733|T201|COMP|48257-0|LNC|Holcus lanatus leukotriene release|Holcus lanatus leukotriene release
C1953735|T201|COMP|48258-8|LNC|Secale cereale pollen leukotriene release|Secale cereale pollen leukotriene release
C1953737|T201|COMP|48259-6|LNC|Poa pratensis leukotriene release|Poa pratensis leukotriene release
C1953739|T201|COMP|48260-4|LNC|Phleum pratense leukotriene release|Phleum pratense leukotriene release
C1953741|T201|COMP|48261-2|LNC|Lolium perenne leukotriene release|Lolium perenne leukotriene release
C1953743|T201|COMP|48262-0|LNC|Festuca elatior leukotriene release|Festuca elatior leukotriene release
C1953745|T201|COMP|48263-8|LNC|Dactylis glomerata leukotriene release|Dactylis glomerata leukotriene release
C1953747|T201|COMP|48264-6|LNC|Cynodon dactylon leukotriene release|Cynodon dactylon leukotriene release
C1953753|T201|COMP|48267-9|LNC|Benzylpenicilloyl-polylysine leukotriene release|Benzylpenicilloyl-polylysine leukotriene release
C1953755|T201|COMP|48268-7|LNC|Minor determinant mixture leukotriene release|Minor determinant mixture leukotriene release
C1953757|T201|COMP|48269-5|LNC|Cefamandole leukotriene release|Cefamandole leukotriene release
C1953759|T201|COMP|48270-3|LNC|ceFAZolin leukotriene release|ceFAZolin leukotriene release
C1953761|T201|COMP|48271-1|LNC|Tetracycline leukotriene release|Tetracycline leukotriene release
C1953763|T201|COMP|48272-9|LNC|Ciprofloxacin leukotriene release|Ciprofloxacin leukotriene release
C1953765|T201|COMP|48273-7|LNC|Lysine acetylsalicylate leukotriene release|Lysine acetylsalicylate leukotriene release
C1953767|T201|COMP|48274-5|LNC|Diclofenac leukotriene release|Diclofenac leukotriene release
C1953769|T201|COMP|48275-2|LNC|Ibuprofen leukotriene release|Ibuprofen leukotriene release
C1953771|T201|COMP|48276-0|LNC|Indomethacin leukotriene release|Indomethacin leukotriene release
C1953773|T201|COMP|48277-8|LNC|Acetaminophen leukotriene release|Acetaminophen leukotriene release
C1953775|T201|COMP|48278-6|LNC|Mefenamate leukotriene release|Mefenamate leukotriene release
C1953777|T201|COMP|48279-4|LNC|Propyphenazone leukotriene release|Propyphenazone leukotriene release
C1953779|T201|COMP|48280-2|LNC|Dipyrone leukotriene release|Dipyrone leukotriene release
C1953781|T201|COMP|48281-0|LNC|Sulfamethoxazole leukotriene release|Sulfamethoxazole leukotriene release
C1953783|T201|COMP|48282-8|LNC|Atracurium leukotriene release|Atracurium leukotriene release
C1953785|T201|COMP|48283-6|LNC|Mivacurium leukotriene release|Mivacurium leukotriene release
C1953787|T201|COMP|48284-4|LNC|Pancuronium leukotriene release|Pancuronium leukotriene release
C1953789|T201|COMP|48285-1|LNC|Propofol leukotriene release|Propofol leukotriene release
C1953791|T201|COMP|48286-9|LNC|Rocuronium leukotriene release|Rocuronium leukotriene release
C1953793|T201|COMP|48287-7|LNC|Suxamethonium leukotriene release|Suxamethonium leukotriene release
C1953795|T201|COMP|48288-5|LNC|Vecuronium leukotriene release|Vecuronium leukotriene release
C1953797|T201|COMP|48298-4|LNC|Pigweed leukotriene release|Pigweed leukotriene release
C1953799|T201|COMP|48299-2|LNC|New coccine leukotriene release|New coccine leukotriene release
C1953801|T201|COMP|48300-8|LNC|Erythrosine leukotriene release|Erythrosine leukotriene release
C1953803|T201|COMP|48301-6|LNC|Patent blue V leukotriene release|Patent blue V leukotriene release
C1953805|T201|COMP|48302-4|LNC|Indigo carmine leukotriene release|Indigo carmine leukotriene release
C1953807|T201|COMP|48303-2|LNC|Brilliant black BN leukotriene release|Brilliant black BN leukotriene release
C1953809|T201|COMP|48304-0|LNC|Glutamate leukotriene release|Glutamate leukotriene release
C1953811|T201|COMP|48305-7|LNC|Coproporphyrin 1/Creatinine|Coproporphyrin 1/Creatinine
C1953812|T201|COMP|48306-5|LNC|Coproporphyrin 3/Creatinine|Coproporphyrin 3/Creatinine
C1953813|T201|COMP|48307-3|LNC|Didanosine|Didanosine
C1953814|T201|COMP|48308-1|LNC|DNA double strand Ab|DNA double strand Ab
C1953815|T201|COMP|48309-9|LNC|BK virus DNA|BK virus DNA
C1953816|T201|COMP|48310-7|LNC|Influenza virus A|Influenza virus A
C1953817|T201|COMP|48311-5|LNC|Lysosomal enzymes screen|Lysosomal enzymes screen
C1953818|T201|COMP|48312-3|LNC|Yersinia enterocolitica O:5 Ab|Yersinia enterocolitica O:5 Ab
C1953819|T201|COMP|48313-1|LNC|Yersinia enterocolitica O:9 Ab|Yersinia enterocolitica O:9 Ab
C1953820|T201|COMP|48314-9|LNC|Leishmania mexicana Ab.IgG|Leishmania mexicana Ab.IgG
C1953821|T201|COMP|48315-6|LNC|Leishmania mexicana Ab.IgM|Leishmania mexicana Ab.IgM
C1953822|T201|COMP|48316-4|LNC|Leishmania tropica Ab.IgG|Leishmania tropica Ab.IgG
C1953823|T201|COMP|48317-2|LNC|Leishmania tropica Ab.IgM|Leishmania tropica Ab.IgM
C1953824|T201|COMP|48318-0|LNC|Cat hair+Cat epithelium Ab.IgE.RAST class|Cat hair+Cat epithelium Ab.IgE.RAST class
C1953826|T201|COMP|48319-8|LNC|glipiZIDE|glipiZIDE
C1953827|T201|COMP|48320-6|LNC|glyBURIDE|glyBURIDE
C1953828|T201|COMP|48321-4|LNC|TOLBUTamide|TOLBUTamide
C1953829|T201|COMP|48322-2|LNC|acetoHEXAMIDE|acetoHEXAMIDE
C1953830|T201|COMP|48323-0|LNC|TOLAZamide|TOLAZamide
C1953831|T201|COMP|48324-8|LNC|chlorproPAMIDE|chlorproPAMIDE
C1953832|T201|COMP|48325-5|LNC|Glimepiride|Glimepiride
C1953833|T201|COMP|48326-3|LNC|glipiZIDE|glipiZIDE
C1953834|T201|COMP|48327-1|LNC|glyBURIDE|glyBURIDE
C1953835|T201|COMP|48328-9|LNC|Repaglinide|Repaglinide
C1953836|T201|COMP|48329-7|LNC|chlorproPAMIDE|chlorproPAMIDE
C1953837|T201|COMP|48330-5|LNC|MCOLN1 gene mutations tested for|MCOLN1 gene mutations tested for
C1953839|T201|COMP|48331-3|LNC|BLM gene mutations tested for|BLM gene mutations tested for
C1953845|T201|COMP|48335-4|LNC|Aspergillus sp Ag|Aspergillus sp Ag
C1953847|T201|COMP|48336-2|LNC|Candida sp Ag|Candida sp Ag
C1953848|T201|COMP|48337-0|LNC|Cryptococcus neoformans Ag|Cryptococcus neoformans Ag
C1953849|T201|COMP|48338-8|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1953850|T201|COMP|48339-6|LNC|Sporothrix schenckii Ag|Sporothrix schenckii Ag
C1953851|T201|COMP|48340-4|LNC|17-Hydroxyprogesterone^30M post XXX challenge|17-Hydroxyprogesterone^30M post XXX challenge
C1953852|T201|COMP|48341-2|LNC|17-Hydroxyprogesterone^1H post XXX challenge|17-Hydroxyprogesterone^1H post XXX challenge
C1953853|T201|COMP|48342-0|LNC|Ethanol+Methanol+Isopropyl alcohol+Acetone|Ethanol+Methanol+Isopropyl alcohol+Acetone
C1953855|T201|COMP|48343-8|LNC|Hemoglobin.other/Hemoglobin.total|Hemoglobin.other/Hemoglobin.total
C1953856|T201|COMP|48344-6|LNC|Activated clotting time|Activated clotting time
C1953857|T201|COMP|48345-3|LNC|HIV 1+O+2 Ab|HIV 1+O+2 Ab
C1953859|T201|COMP|48346-1|LNC|HIV 1+O+2 Ab|HIV 1+O+2 Ab
C1953860|T201|COMP|48347-9|LNC|levETIRAcetam|levETIRAcetam
C1953861|T201|COMP|48348-7|LNC|10-Hydroxycarbazepine|10-Hydroxycarbazepine
C1953862|T201|COMP|48349-5|LNC|Pregabalin|Pregabalin
C1953863|T201|COMP|48350-3|LNC|Venlafaxine+Norvenlafaxine|Venlafaxine+Norvenlafaxine
C1953865|T201|COMP|48351-1|LNC|Methotrimeprazine|Methotrimeprazine
C1953866|T201|COMP|48352-9|LNC|Reboxetine|Reboxetine
C1953867|T201|COMP|48353-7|LNC|Chlorprothixene|Chlorprothixene
C1953868|T201|COMP|48354-5|LNC|ARIPiprazole|ARIPiprazole
C1953869|T201|COMP|48355-2|LNC|traMADol|traMADol
C1953870|T201|COMP|48356-0|LNC|Prazepam|Prazepam
C1953871|T201|COMP|48357-8|LNC|Testosterone|Testosterone
C1953872|T201|COMP|48358-6|LNC|Herpes virus 8 Ab.IgM|Herpes virus 8 Ab.IgM
C1953874|T201|COMP|48359-4|LNC|Echinococcus granulosus Ab|Echinococcus granulosus Ab
C1953875|T201|COMP|48360-2|LNC|Borrelia afzelii Ab.IgG|Borrelia afzelii Ab.IgG
C1953877|T201|COMP|48361-0|LNC|Borrelia valaisiana Ab.IgG|Borrelia valaisiana Ab.IgG
C1953879|T201|COMP|48362-8|LNC|Norvenlafaxine|Norvenlafaxine
C1953880|T201|COMP|48363-6|LNC|Morphine-6-Glucuronide|Morphine-6-Glucuronide
C1953881|T201|COMP|48385-9|LNC|Collagen.injectable Ab|Collagen.injectable Ab
C1953883|T201|COMP|48386-7|LNC|Platelets.large/Platelets|Platelets.large/Platelets
C1953885|T201|COMP|48387-5|LNC|Thyroglobulin recovery|Thyroglobulin recovery
C1953886|T201|COMP|48388-3|LNC|Heparin Ab.IgE|Heparin Ab.IgE
C1953888|T201|COMP|48389-1|LNC|Macroprolactin/Prolactin|Macroprolactin/Prolactin
C1953890|T201|COMP|48390-9|LNC|B cell crossmatch|B cell crossmatch
C1953891|T201|COMP|48391-7|LNC|Carbon dioxide|Carbon dioxide
C1953892|T201|COMP|48392-5|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C1953893|T201|COMP|48393-3|LNC|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C1953894|T201|COMP|48394-1|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1953895|T201|COMP|48395-8|LNC|Coproporphyrin/Creatinine|Coproporphyrin/Creatinine
C1953896|T201|COMP|48396-6|LNC|Ganglioside GD1b Ab|Ganglioside GD1b Ab
C1953898|T201|COMP|48398-2|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1953899|T201|COMP|48399-0|LNC|Herpes simplex virus 1 glycoprotein G Ab.IgG|Herpes simplex virus 1 glycoprotein G Ab.IgG
C1953900|T201|COMP|48400-6|LNC|Herpes simplex virus 1+2 Ag|Herpes simplex virus 1+2 Ag
C1953901|T201|COMP|48401-4|LNC|Herpes simplex virus 2 glycoprotein G Ab.IgG|Herpes simplex virus 2 glycoprotein G Ab.IgG
C1953902|T201|COMP|48402-2|LNC|Latex Ab.IgE/IgE.total|Latex Ab.IgE/IgE.total
C1953903|T201|COMP|48403-0|LNC|Methadone+Metabolite|Methadone+Metabolite
C1953904|T201|COMP|48404-8|LNC|Myeloperoxidase Ab.IgG|Myeloperoxidase Ab.IgG
C1953906|T201|COMP|48405-5|LNC|Neuronal nuclear Ab.IgG|Neuronal nuclear Ab.IgG
C1953907|T201|COMP|48406-3|LNC|Parietal cell Ab.IgG|Parietal cell Ab.IgG
C1953908|T201|COMP|48407-1|LNC|Pregnancy associated plasma protein A|Pregnancy associated plasma protein A
C1953909|T201|COMP|48408-9|LNC|Proteinase 3 Ab.IgG|Proteinase 3 Ab.IgG
C1953911|T201|COMP|48409-7|LNC|T cell crossmatch|T cell crossmatch
C1953912|T201|COMP|48410-5|LNC|Yersinia sp Ab.IgM|Yersinia sp Ab.IgM
C1953913|T201|COMP|48411-3|LNC|Fungus identified|Fungus identified
C1953914|T201|COMP|48412-1|LNC|Zygomycete sp Ag|Zygomycete sp Ag
C1953915|T201|COMP|48413-9|LNC|Alpha-1-Microglobulin|Alpha-1-Microglobulin
C1953916|T201|COMP|48414-7|LNC|Alpha-1-Microglobulin|Alpha-1-Microglobulin
C1953917|T201|COMP|48415-4|LNC|Alpha-1-Microglobulin/Creatinine|Alpha-1-Microglobulin/Creatinine
C1953919|T201|COMP|48416-2|LNC|Alpha-1-Acid glycoprotein|Alpha-1-Acid glycoprotein
C1953920|T201|COMP|48417-0|LNC|Staphylolysin Ab|Staphylolysin Ab
C1953921|T201|COMP|48418-8|LNC|Staphylolysin Ab|Staphylolysin Ab
C1953922|T201|COMP|48419-6|LNC|Immune complex.IgG|Immune complex.IgG
C1953923|T201|COMP|48420-4|LNC|Complement C3c|Complement C3c
C1953924|T201|COMP|48421-2|LNC|C reactive protein|C reactive protein
C1953925|T201|COMP|48422-0|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C1953926|T201|COMP|48423-8|LNC|Protein pattern|Protein pattern
C1953927|T201|COMP|48424-6|LNC|Protein pattern|Protein pattern
C1953928|T201|COMP|48425-3|LNC|Troponin T.cardiac|Troponin T.cardiac
C1953929|T201|COMP|48426-1|LNC|Troponin T.cardiac|Troponin T.cardiac
C1953932|T201|COMP|48428-7|LNC|Rumenate|Rumenate
C1953934|T201|COMP|48429-5|LNC|Lavandula angustifolia Ab.IgE|Lavandula angustifolia Ab.IgE
C1953936|T201|COMP|48430-3|LNC|Carnitine|Carnitine
C1953937|T201|COMP|48431-1|LNC|Zinc|Zinc
C1953938|T201|COMP|48432-9|LNC|Fructose|Fructose
C1953994|T201|COMP|48494-9|LNC|Complement C1 esterase inhibitor actual/Normal|Complement C1 esterase inhibitor actual/Normal
C1953998|T201|COMP|48496-4|LNC|Complement total hemolytic CH50 actual/Normal|Complement total hemolytic CH50 actual/Normal
C1954000|T201|COMP|48497-2|LNC|Pro-hepcidin|Pro-hepcidin
C1954002|T201|COMP|48498-0|LNC|Amyloid A|Amyloid A
C1954003|T201|COMP|48499-8|LNC|Beta-trace protein|Beta-trace protein
C1954004|T201|COMP|48500-3|LNC|Borrelia burgdorferi 18kD Ab.IgG|Borrelia burgdorferi 18kD Ab.IgG
C1954005|T201|COMP|48501-1|LNC|HLA Ab|HLA Ab
C1954006|T201|COMP|48502-9|LNC|Platelet glycoprotein Ia-IIa Ab.IgG|Platelet glycoprotein Ia-IIa Ab.IgG
C1954008|T201|COMP|48503-7|LNC|Platelet glycoprotein Ib-Ix Ab.IgG|Platelet glycoprotein Ib-Ix Ab.IgG
C1954010|T201|COMP|48504-5|LNC|Platelet glycoprotein IIb-IIIa Ab.IgG|Platelet glycoprotein IIb-IIIa Ab.IgG
C1954012|T201|COMP|48505-2|LNC|Platelet glycoprotein IIb-IIIa Ab|Platelet glycoprotein IIb-IIIa Ab
C1954014|T201|COMP|48506-0|LNC|Platelet glycoprotein Ib-Ix Ab|Platelet glycoprotein Ib-Ix Ab
C1954016|T201|COMP|48507-8|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C1954017|T201|COMP|48508-6|LNC|Measles virus RNA|Measles virus RNA
C1954018|T201|COMP|48509-4|LNC|Influenza virus A & B RNA|Influenza virus A & B RNA
C1954020|T201|COMP|48510-2|LNC|HIV 1 RNA|HIV 1 RNA
C1954021|T201|COMP|48511-0|LNC|HIV 1 RNA|HIV 1 RNA
C1954112|T201|COMP|48551-6|LNC|HIV 1 RNA|HIV 1 RNA
C1954113|T201|COMP|48552-4|LNC|HIV 1 RNA|HIV 1 RNA
C1954114|T201|COMP|48553-2|LNC|Muscle sarcolemma Ab|Muscle sarcolemma Ab
C1954115|T201|COMP|48554-0|LNC|Myocardium Ab|Myocardium Ab
C1954116|T201|COMP|48555-7|LNC|Fetal blood|Fetal blood
C1954117|T201|COMP|48556-5|LNC|Erythrocytes.fetal/1000 erythrocytes|Erythrocytes.fetal/1000 erythrocytes
C1954119|T201|COMP|48557-3|LNC|Origin|Origin
C1954120|T201|COMP|48558-1|LNC|HIV genotype|HIV genotype
C1954122|T201|COMP|48559-9|LNC|HIV genotype|HIV genotype
C1954123|T201|COMP|48560-7|LNC|Human papilloma virus genotype|Human papilloma virus genotype
C1954125|T201|COMP|48561-5|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1954126|T201|COMP|48562-3|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1954127|T201|COMP|48563-1|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C1954128|T201|COMP|48564-9|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C1954129|T201|COMP|48565-6|LNC|Bacteria identified^^^6|Bacteria identified^^^6
C1954130|T201|COMP|48566-4|LNC|Bacteria identified^^^7|Bacteria identified^^^7
C1954131|T201|COMP|48567-2|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1954132|T201|COMP|48568-0|LNC|Bacteria identified^^^7|Bacteria identified^^^7
C1954133|T201|COMP|48569-8|LNC|Bacteria identified^^^8|Bacteria identified^^^8
C1954134|T201|COMP|48570-6|LNC|Follitropin^on cycle day 10|Follitropin^on cycle day 10
C1954135|T201|COMP|48571-4|LNC|Follitropin^on cycle day 11|Follitropin^on cycle day 11
C1954136|T201|COMP|48572-2|LNC|Follitropin^on cycle day 21|Follitropin^on cycle day 21
C1954137|T201|COMP|48573-0|LNC|Follitropin^on cycle day 3|Follitropin^on cycle day 3
C1954138|T201|COMP|48574-8|LNC|Hepatitis C virus genotype|Hepatitis C virus genotype
C1954139|T201|COMP|48575-5|LNC|Hepatitis C virus genotype|Hepatitis C virus genotype
C1954140|T201|COMP|48576-3|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1954143|T201|COMP|48578-9|LNC|HFE gene.c.187G>C|HFE gene.c.187G>C
C1954147|T201|COMP|48580-5|LNC|KCNQ1OT1 gene targeted mutation analysis|KCNQ1OT1 gene targeted mutation analysis
C1954149|T201|COMP|48581-3|LNC|Lutropin^on cycle day 11|Lutropin^on cycle day 11
C1954150|T201|COMP|48582-1|LNC|Lutropin^on cycle day 3|Lutropin^on cycle day 3
C1954151|T201|COMP|48583-9|LNC|Lutropin^on cycle day 21|Lutropin^on cycle day 21
C1954155|T201|COMP|48586-2|LNC|Collagen crosslinked C-telopeptide|Collagen crosslinked C-telopeptide
C1954156|T201|COMP|48587-0|LNC|Collagen crosslinked C-telopeptide/Creatinine|Collagen crosslinked C-telopeptide/Creatinine
C1954158|T201|COMP|48588-8|LNC|Coccidioides sp rRNA|Coccidioides sp rRNA
C1954160|T201|COMP|48589-6|LNC|Coccidioides sp rRNA|Coccidioides sp rRNA
C1954161|T201|COMP|48590-4|LNC|Coagulation surface induced^after addition of APC|Coagulation surface induced^after addition of APC
C1954162|T201|COMP|48591-2|LNC|Activated protein C resistance|Activated protein C resistance
C1954163|T201|COMP|48592-0|LNC|Fibrin+Fibrinogen fragments|Fibrin+Fibrinogen fragments
C1954164|T201|COMP|48593-8|LNC|von Willebrand panel|von Willebrand panel
C1954166|T201|COMP|48594-6|LNC|Platelet glycoprotein IIb-IIIa Ab|Platelet glycoprotein IIb-IIIa Ab
C1954167|T201|COMP|48595-3|LNC|von Willebrand evaluation|von Willebrand evaluation
C1954169|T201|COMP|48596-1|LNC|Activated protein C resistance panel|Activated protein C resistance panel
C1954171|T201|COMP|48597-9|LNC|cycloSPORINE^trough|cycloSPORINE^trough
C1954172|T201|COMP|48598-7|LNC|BBS2 gene targeted mutation analysis|BBS2 gene targeted mutation analysis
C1954174|T201|COMP|48599-5|LNC|CLCN1 gene targeted mutation analysis|CLCN1 gene targeted mutation analysis
C1954176|T201|COMP|48600-1|LNC|VPS13B gene targeted mutation analysis|VPS13B gene targeted mutation analysis
C1954178|T201|COMP|48601-9|LNC|OPA1 gene targeted mutation analysis|OPA1 gene targeted mutation analysis
C1954180|T201|COMP|48602-7|LNC|TGM1 gene targeted mutation analysis|TGM1 gene targeted mutation analysis
C1954182|T201|COMP|48604-3|LNC|Yellow dye Ab.IgE.RAST class|Yellow dye Ab.IgE.RAST class
C1954184|T201|COMP|48605-0|LNC|Glucose^1H post dose fructose PO|Glucose^1H post dose fructose PO
C1954185|T201|COMP|48606-8|LNC|Glucose^pre dose fructose PO|Glucose^pre dose fructose PO
C1954186|T201|COMP|48607-6|LNC|Glucose^30M post dose fructose PO|Glucose^30M post dose fructose PO
C1954187|T201|COMP|48608-4|LNC|2-Hydroxyvalerate/Creatinine|2-Hydroxyvalerate/Creatinine
C1954189|T201|COMP|48609-2|LNC|Adenovirus DNA|Adenovirus DNA
C1954190|T201|COMP|48610-0|LNC|7-Dehydrocholesterol|7-Dehydrocholesterol
C1954191|T201|COMP|48611-8|LNC|Antibiotic tested|Antibiotic tested
C1954192|T201|COMP|48612-6|LNC|Hydrogen/Expired gas^45M post dose lactose PO|Hydrogen/Expired gas^45M post dose lactose PO
C1954193|T201|COMP|48613-4|LNC|Hydrogen/Expired gas^15M post dose lactose PO|Hydrogen/Expired gas^15M post dose lactose PO
C1954194|T201|COMP|48614-2|LNC|Cryoglobulin|Cryoglobulin
C1954195|T201|COMP|48615-9|LNC|Insulin.free & Insulin.total panel|Insulin.free & Insulin.total panel
C1954197|T201|COMP|48616-7|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C1954198|T201|COMP|48617-5|LNC|Phosphate^post dialysis|Phosphate^post dialysis
C1954199|T201|COMP|48618-3|LNC|Cholesterol.in VLDL|Cholesterol.in VLDL
C1954200|T201|COMP|48619-1|LNC|Apolipoprotein E1|Apolipoprotein E1
C1954202|T201|COMP|48620-9|LNC|Cholesterol|Cholesterol
C1954203|T201|COMP|48621-7|LNC|Hexacarboxylporphyrin/Creatinine|Hexacarboxylporphyrin/Creatinine
C1954204|T201|COMP|48622-5|LNC|Urea nitrogen^24H post peritoneal dialysis|Urea nitrogen^24H post peritoneal dialysis
C1954205|T201|COMP|48623-3|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C1954206|T201|COMP|48624-1|LNC|Bilirubin|Bilirubin
C1954207|T201|COMP|48625-8|LNC|Choriogonadotropin.intact|Choriogonadotropin.intact
C1954208|T201|COMP|48626-6|LNC|Creatinine^24H post peritoneal dialysis|Creatinine^24H post peritoneal dialysis
C1954209|T201|COMP|48627-4|LNC|Protein.monoclonal|Protein.monoclonal
C1954210|T201|COMP|48628-2|LNC|Insulin-like growth factor binding protein 3|Insulin-like growth factor binding protein 3
C1954211|T201|COMP|48629-0|LNC|Urea nitrogen^post dialysis|Urea nitrogen^post dialysis
C1954212|T201|COMP|48630-8|LNC|Creatinine^pre dialysis|Creatinine^pre dialysis
C1954213|T201|COMP|48631-6|LNC|Bicarbonate^post dialysis|Bicarbonate^post dialysis
C1954214|T201|COMP|48632-4|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C1954215|T201|COMP|48633-2|LNC|Trypsinogen I.free|Trypsinogen I.free
C1954216|T201|COMP|48634-0|LNC|Coproporphyrin/Creatinine|Coproporphyrin/Creatinine
C1954217|T201|COMP|48635-7|LNC|Cholesterol.in LDL pattern A|Cholesterol.in LDL pattern A
C1954219|T201|COMP|48636-5|LNC|Cholesterol.in LDL pattern BII|Cholesterol.in LDL pattern BII
C1954221|T201|COMP|48637-3|LNC|Cholesterol.in LDL pattern BI|Cholesterol.in LDL pattern BI
C1954223|T201|COMP|48638-1|LNC|Cryoglobulin type|Cryoglobulin type
C1954224|T201|COMP|48639-9|LNC|Urea nitrogen^post dialysis|Urea nitrogen^post dialysis
C1954225|T201|COMP|48640-7|LNC|Second trimester triple maternal screen|Second trimester triple maternal screen
C1954227|T201|COMP|48641-5|LNC|Phosphate^pre dialysis|Phosphate^pre dialysis
C1954234|T201|COMP|48645-6|LNC|Pseudomonas sp DNA|Pseudomonas sp DNA
C1954236|T201|COMP|48646-4|LNC|Yersinia sp DNA|Yersinia sp DNA
C1954238|T201|COMP|48647-2|LNC|Ej Ab|Ej Ab
C1954239|T201|COMP|48648-0|LNC|MART-1|MART-1
C1954240|T201|COMP|48649-8|LNC|OJ Ab|OJ Ab
C1954241|T201|COMP|48650-6|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1954242|T201|COMP|48651-4|LNC|Borrelia burgdorferi Ab.IgM index|Borrelia burgdorferi Ab.IgM index
C1954244|T201|COMP|48652-2|LNC|Clostridium tetani toxoid Ab.IgG^2nd specimen|Clostridium tetani toxoid Ab.IgG^2nd specimen
C1954246|T201|COMP|48653-0|LNC|Clostridium tetani toxoid Ab.IgG^1st specimen|Clostridium tetani toxoid Ab.IgG^1st specimen
C1954247|T201|COMP|48654-8|LNC|Corynebacterium diphtheriae toxin Ab.IgG|Corynebacterium diphtheriae toxin Ab.IgG
C1954249|T201|COMP|48655-5|LNC|Corynebacterium diphtheriae toxin Ab^2nd specimen|Corynebacterium diphtheriae toxin Ab^2nd specimen
C1954250|T201|COMP|48656-3|LNC|Ganglioside GD1a Ab|Ganglioside GD1a Ab
C1954251|T201|COMP|48657-1|LNC|Ganglioside GM2 Ab|Ganglioside GM2 Ab
C1954253|T201|COMP|48658-9|LNC|Ganglioside GQ1b Ab|Ganglioside GQ1b Ab
C1954254|T201|COMP|48659-7|LNC|Hepatitis B virus precore codon 28|Hepatitis B virus precore codon 28
C1954256|T201|COMP|48660-5|LNC|Ganglioside GM1 Ab|Ganglioside GM1 Ab
C1954260|T201|COMP|48663-9|LNC|YKL-40|YKL-40
C1954262|T201|COMP|48664-7|LNC|Fibrinogen|Fibrinogen
C1954263|T201|COMP|48665-4|LNC|IgA.intrathecally synthesized|IgA.intrathecally synthesized
C1954265|T201|COMP|48666-2|LNC|IgG.intrathecally synthesized|IgG.intrathecally synthesized
C1954267|T201|COMP|48667-0|LNC|IgM.intrathecally synthesized|IgM.intrathecally synthesized
C1954269|T201|COMP|48668-8|LNC|Protein fractions.oligoclonal bands.IT|Protein fractions.oligoclonal bands.IT
C1954271|T201|COMP|48669-6|LNC|Albumin & Immunoglobulin Quotient|Albumin & Immunoglobulin Quotient
C1954273|T201|COMP|48670-4|LNC|IgVH gene targeted mutation analysis|IgVH gene targeted mutation analysis
C1954275|T201|COMP|48671-2|LNC|Prostate cancer risk|Prostate cancer risk
C1954277|T201|COMP|48672-0|LNC|Clinical cytogeneticist|Clinical cytogeneticist
C1954278|T201|COMP|48673-8|LNC|EBV-LMP Ag|EBV-LMP Ag
C1954280|T201|COMP|48674-6|LNC|Genetic diseases|Genetic diseases
C1954281|T201|COMP|48675-3|LNC|HER2|HER2
C1954282|T201|COMP|48676-1|LNC|HER2|HER2
C1954283|T201|COMP|48677-9|LNC|Cancer Ag 125|Cancer Ag 125
C1954284|T201|COMP|48678-7|LNC|P57 Ag|P57 Ag
C1954286|T201|COMP|48679-5|LNC|Pancytokeratin Ag|Pancytokeratin Ag
C1954288|T201|COMP|48680-3|LNC|PAX5 Ag|PAX5 Ag
C1954290|T201|COMP|48681-1|LNC|Plasma cell Ag|Plasma cell Ag
C1954292|T201|COMP|48682-9|LNC|Smooth muscle myosin heavy chain Ag|Smooth muscle myosin heavy chain Ag
C1954294|T201|COMP|48683-7|LNC|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C1954296|T201|COMP|48684-5|LNC|X & Y chromosome^post bone marrow transplant|X & Y chromosome^post bone marrow transplant
C1954298|T201|COMP|48685-2|LNC|Para aminosalicylate 10.0 ug/mL|Para aminosalicylate 10.0 ug/mL
C1954300|T201|COMP|48686-0|LNC|Salmonella paratyphi C Ab|Salmonella paratyphi C Ab
C1954316|T201|COMP|48700-9|LNC|Thyrotropin releasing hormone|Thyrotropin releasing hormone
C1954317|T201|COMP|48701-7|LNC|Lutenizing releasing hormone|Lutenizing releasing hormone
C1954319|T201|COMP|48702-5|LNC|Spermatozoa.immature/100 spermatozoa|Spermatozoa.immature/100 spermatozoa
C1954321|T201|COMP|48703-3|LNC|Hematocrit|Hematocrit
C1954322|T201|COMP|48704-1|LNC|Unidentified cells|Unidentified cells
C1954323|T201|COMP|48705-8|LNC|Leukocytes+Platelets|Leukocytes+Platelets
C1954325|T201|COMP|48706-6|LNC|Reticulocyte mean volume|Reticulocyte mean volume
C1954327|T201|COMP|48707-4|LNC|Hemoglobin C crystals|Hemoglobin C crystals
C1954328|T201|COMP|48708-2|LNC|Erythrocytes.fresh/100 erythrocytes|Erythrocytes.fresh/100 erythrocytes
C1954330|T201|COMP|48709-0|LNC|Burr cells/100 erythrocytes|Burr cells/100 erythrocytes
C1954332|T201|COMP|48710-8|LNC|Eosinophils|Eosinophils
C1954333|T201|COMP|48711-6|LNC|Hemoglobin.free^post transfusion reaction|Hemoglobin.free^post transfusion reaction
C1954335|T201|COMP|48713-2|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C1954336|T201|COMP|48714-0|LNC|Leishmania tropica Ab.IgM|Leishmania tropica Ab.IgM
C1954337|T201|COMP|48715-7|LNC|Leishmania tropica Ab.IgG|Leishmania tropica Ab.IgG
C1954338|T201|COMP|48716-5|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C1954339|T201|COMP|48717-3|LNC|Leishmania mexicana Ab.IgM|Leishmania mexicana Ab.IgM
C1954340|T201|COMP|48718-1|LNC|Leishmania mexicana Ab.IgG|Leishmania mexicana Ab.IgG
C1954341|T201|COMP|48719-9|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C1954342|T201|COMP|48720-7|LNC|Coxiella burnetii phase 1 Ab.IgG|Coxiella burnetii phase 1 Ab.IgG
C1954343|T201|COMP|48721-5|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C1954345|T201|COMP|48723-1|LNC|Epstein Barr virus Ab|Epstein Barr virus Ab
C1954346|T201|COMP|48724-9|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C1954347|T201|COMP|48725-6|LNC|Hemoglobin^pre therapeutic phlebotomy|Hemoglobin^pre therapeutic phlebotomy
C1954348|T201|COMP|48726-4|LNC|JAK2 gene targeted mutation analysis|JAK2 gene targeted mutation analysis
C1954350|T201|COMP|48727-2|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C1954351|T201|COMP|48728-0|LNC|NCF1+NCF2+CYBB gene targeted mutation analysis|NCF1+NCF2+CYBB gene targeted mutation analysis
C1954353|T201|COMP|48729-8|LNC|CYBA gene targeted mutation analysis|CYBA gene targeted mutation analysis
C1954355|T201|COMP|48730-6|LNC|X linked heterotaxy|X linked heterotaxy
C1954357|T201|COMP|48731-4|LNC|Complement C4|Complement C4
C1954358|T201|COMP|48732-2|LNC|NCF1 gene targeted mutation analysis|NCF1 gene targeted mutation analysis
C1954360|T201|COMP|48733-0|LNC|NCF2 gene targeted mutation analysis|NCF2 gene targeted mutation analysis
C1954361|T201|COMP|48734-8|LNC|CYBB gene targeted mutation analysis|CYBB gene targeted mutation analysis
C1954370|T201|COMP|48741-3|LNC|Bordetella pertussis|Bordetella pertussis
C1954377|T201|COMP|48756-1|LNC|3-Hydroxyoctanoate.free|3-Hydroxyoctanoate.free
C1954379|T201|COMP|48757-9|LNC|3-Hydroxyoctanoate|3-Hydroxyoctanoate
C1954380|T201|COMP|48758-7|LNC|3-Hydroxyhexanoate.free|3-Hydroxyhexanoate.free
C1954382|T201|COMP|48759-5|LNC|3-Hydroxyhexanoate|3-Hydroxyhexanoate
C1954383|T201|COMP|48760-3|LNC|3-Hydroxy fatty acid panel|3-Hydroxy fatty acid panel
C1954385|T201|COMP|48761-1|LNC|3-Hydroxypalmitate|3-Hydroxypalmitate
C1954387|T201|COMP|48762-9|LNC|3-Hydroxymyristate|3-Hydroxymyristate
C1954389|T201|COMP|48763-7|LNC|3-Hydroxydecanoate|3-Hydroxydecanoate
C1954403|T201|COMP|48771-0|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C1954404|T201|COMP|48772-8|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C1954406|T201|COMP|48774-4|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C1954407|T201|COMP|48775-1|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C1954409|T201|COMP|48777-7|LNC|Immunoglobulin light chains.kappa.free/Albumin|Immunoglobulin light chains.kappa.free/Albumin
C1954411|T201|COMP|48778-5|LNC|Erythrocytes.nucleated/100 cells|Erythrocytes.nucleated/100 cells
C1954416|T201|COMP|48781-9|LNC|CYP21A2 gene targeted mutation analysis|CYP21A2 gene targeted mutation analysis
C1954417|T201|COMP|48782-7|LNC|Dipyrone Ab.IgE.RAST class|Dipyrone Ab.IgE.RAST class
C1954419|T201|COMP|48783-5|LNC|Dipyrone Ab.IgE|Dipyrone Ab.IgE
C1954421|T201|COMP|48784-3|LNC|Herpes simplex virus 2 Ab|Herpes simplex virus 2 Ab
C1954422|T201|COMP|48785-0|LNC|Prostaglandin D2|Prostaglandin D2
C1954423|T201|COMP|48786-8|LNC|Renin^30M pre XXX challenge|Renin^30M pre XXX challenge
C1954424|T201|COMP|48787-6|LNC|Glucose^24H post peritoneal dialysis|Glucose^24H post peritoneal dialysis
C1954425|T201|COMP|48788-4|LNC|Creatinine peritoneal dialysis clearance|Creatinine peritoneal dialysis clearance
C1954427|T201|COMP|48790-0|LNC|Creatinine|Creatinine
C1954430|T201|COMP|48792-6|LNC|Necroinflammatory activity score|Necroinflammatory activity score
C1954432|T201|COMP|48793-4|LNC|Necroinflammatory activity grade|Necroinflammatory activity grade
C1954434|T201|COMP|48794-2|LNC|Fibrosis stage|Fibrosis stage
C1954436|T201|COMP|48795-9|LNC|Liver fibrosis score|Liver fibrosis score
C1954438|T201|COMP|48796-7|LNC|Hepatitis C virus FibroSURE panel|Hepatitis C virus FibroSURE panel
C1954440|T201|COMP|48797-5|LNC|Organic acids panel|Organic acids panel
C1954441|T201|COMP|48798-3|LNC|First trimester maternal screen panel|First trimester maternal screen panel
C1954443|T201|COMP|48799-1|LNC|Second trimester penta maternal screen panel|Second trimester penta maternal screen panel
C1954445|T201|COMP|48800-7|LNC|Second trimester quad maternal screen panel|Second trimester quad maternal screen panel
C1954447|T201|COMP|48802-3|LNC|Alpha-1-fetoprotein panel|Alpha-1-fetoprotein panel
C1954449|T201|COMP|48803-1|LNC|Neural tube defect risk|Neural tube defect risk
C1954451|T201|COMP|48804-9|LNC|Taenia solium Ag|Taenia solium Ag
C1954452|T201|COMP|48805-6|LNC|Platelet aggregation panel|Platelet aggregation panel
C1954458|T201|COMP|48808-0|LNC|Leukogram panel|Leukogram panel
C1954460|T201|COMP|48809-8|LNC|Erythrogram panel|Erythrogram panel
C1954462|T201|COMP|48810-6|LNC|Glucose^5H post 50 g glucose PO|Glucose^5H post 50 g glucose PO
C1954463|T201|COMP|48811-4|LNC|Protein fractions 3 panel|Protein fractions 3 panel
C1954465|T201|COMP|48812-2|LNC|Spermatozoa morphology panel|Spermatozoa morphology panel
C1954467|T201|COMP|48813-0|LNC|Bacterial methicillin resistance mecA gene|Bacterial methicillin resistance mecA gene
C1954469|T201|COMP|48814-8|LNC|Bacterial vancomycin resistance vanA gene|Bacterial vancomycin resistance vanA gene
C1954471|T201|COMP|48815-5|LNC|Herpes simplex virus+Varicella zoster virus DNA|Herpes simplex virus+Varicella zoster virus DNA
C1954474|T201|COMP|48817-1|LNC|Donath Landsteiner Ab|Donath Landsteiner Ab
C1954475|T201|COMP|48818-9|LNC|Karyotype|Karyotype
C1954476|T201|COMP|48819-7|LNC|Karyotype|Karyotype
C1954477|T201|COMP|48820-5|LNC|Karyotype|Karyotype
C1954478|T201|COMP|48821-3|LNC|t(12;21)(p13;q22.3)(ETV6,RUNX1) fusion transcript|t(12;21)(p13;q22.3)(ETV6,RUNX1) fusion transcript
C1954479|T201|COMP|48822-1|LNC|Tubular basement membrane Ab.IgG|Tubular basement membrane Ab.IgG
C1954481|T201|COMP|48823-9|LNC|Tubular basement membrane Ab.IgG|Tubular basement membrane Ab.IgG
C1954490|T201|COMP|48835-3|LNC|Respiratory allergen panel, US - Arid southwest|Respiratory allergen panel, US - Arid southwest
C1954502|T201|COMP|48841-1|LNC|Respiratory allergen panel, US - Alaska a|Respiratory allergen panel, US - Alaska a
C1954504|T201|COMP|48842-9|LNC|Bartonella bacilliformis Ab.IgG|Bartonella bacilliformis Ab.IgG
C1954505|T201|COMP|48843-7|LNC|Bartonella bacilliformis Ab.IgM|Bartonella bacilliformis Ab.IgM
C1954506|T201|COMP|48844-5|LNC|Bartonella elizabethae Ab.IgG|Bartonella elizabethae Ab.IgG
C1954507|T201|COMP|48845-2|LNC|Bartonella elizabethae Ab.IgM|Bartonella elizabethae Ab.IgM
C1954509|T201|COMP|48846-0|LNC|Bartonella vinsonii berkhoffii Ab.IgM|Bartonella vinsonii berkhoffii Ab.IgM
C1954511|T201|COMP|48847-8|LNC|Bartonella vinsonii berkhoffii Ab.IgG|Bartonella vinsonii berkhoffii Ab.IgG
C1954513|T201|COMP|48848-6|LNC|Coxiella burnetii phase 1 Ab.IgA|Coxiella burnetii phase 1 Ab.IgA
C1954514|T201|COMP|48849-4|LNC|Coxiella burnetii phase 2 Ab.IgA|Coxiella burnetii phase 2 Ab.IgA
C1954515|T201|COMP|48850-2|LNC|Ehrlichia chaffeensis Ab.IgM|Ehrlichia chaffeensis Ab.IgM
C1954516|T201|COMP|48851-0|LNC|Orientia tsutsugamushi Gilliam Ab.IgM|Orientia tsutsugamushi Gilliam Ab.IgM
C1954518|T201|COMP|48852-8|LNC|Orientia tsutsugamushi Gilliam Ab.IgG|Orientia tsutsugamushi Gilliam Ab.IgG
C1954520|T201|COMP|48853-6|LNC|Orientia tsutsugamushi Karp Ab.IgG|Orientia tsutsugamushi Karp Ab.IgG
C1954522|T201|COMP|48854-4|LNC|Orientia tsutsugamushi Karp Ab.IgM|Orientia tsutsugamushi Karp Ab.IgM
C1954524|T201|COMP|48855-1|LNC|Orientia tsutsugamushi Kato Ab.IgG|Orientia tsutsugamushi Kato Ab.IgG
C1954526|T201|COMP|48856-9|LNC|Orientia tsutsugamushi Kato Ab.IgM|Orientia tsutsugamushi Kato Ab.IgM
C1954528|T201|COMP|48857-7|LNC|Rickettsia africae Ab.IgM|Rickettsia africae Ab.IgM
C1954530|T201|COMP|48858-5|LNC|Rickettsia africae Ab.IgG|Rickettsia africae Ab.IgG
C1954532|T201|COMP|48859-3|LNC|Rickettsia akari Ab.IgG|Rickettsia akari Ab.IgG
C1954534|T201|COMP|48860-1|LNC|Rickettsia akari Ab.IgM|Rickettsia akari Ab.IgM
C1954536|T201|COMP|48861-9|LNC|Rickettsia parkeri Ab.IgM|Rickettsia parkeri Ab.IgM
C1954538|T201|COMP|48862-7|LNC|Rickettsia parkeri Ab.IgG|Rickettsia parkeri Ab.IgG
C1954540|T201|COMP|48863-5|LNC|Rickettsia sp DNA|Rickettsia sp DNA
C1954542|T201|COMP|48864-3|LNC|Bartonella sp DNA|Bartonella sp DNA
C1954543|T201|COMP|48865-0|LNC|Ehrlichia ewingii DNA|Ehrlichia ewingii DNA
C1954545|T201|COMP|48866-8|LNC|Ehrlichia sp DNA|Ehrlichia sp DNA
C1954547|T201|COMP|48867-6|LNC|Orientia tsutsugamushi DNA|Orientia tsutsugamushi DNA
C1954549|T201|COMP|48868-4|LNC|Rickettsia rickettsii DNA|Rickettsia rickettsii DNA
C1954551|T201|COMP|48869-2|LNC|Rickettsia sp DNA|Rickettsia sp DNA
C1954552|T201|COMP|48870-0|LNC|Rickettsia spotted fever group DNA|Rickettsia spotted fever group DNA
C1954554|T201|COMP|48871-8|LNC|Rickettsia typhus group DNA|Rickettsia typhus group DNA
C1954556|T201|COMP|48872-6|LNC|Anaplasma phagocytophilum|Anaplasma phagocytophilum
C1954557|T201|COMP|48873-4|LNC|Ehrlichia sp identified|Ehrlichia sp identified
C1954559|T201|COMP|48874-2|LNC|Neorickettsia sp|Neorickettsia sp
C1954561|T201|COMP|48875-9|LNC|Orientia tsutsugamushi|Orientia tsutsugamushi
C1954562|T201|COMP|48876-7|LNC|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C1954563|T201|COMP|48877-5|LNC|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C1954564|T201|COMP|48878-3|LNC|Bartonella bacilliformis Ab.IgG|Bartonella bacilliformis Ab.IgG
C1954565|T201|COMP|48879-1|LNC|Bartonella bacilliformis Ab.IgM|Bartonella bacilliformis Ab.IgM
C1954566|T201|COMP|48880-9|LNC|Bartonella elizabethae Ab.IgG|Bartonella elizabethae Ab.IgG
C1954567|T201|COMP|48881-7|LNC|Bartonella elizabethae Ab.IgM|Bartonella elizabethae Ab.IgM
C1954568|T201|COMP|48882-5|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C1954569|T201|COMP|48883-3|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C1954570|T201|COMP|48884-1|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C1954571|T201|COMP|48885-8|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C1954572|T201|COMP|48886-6|LNC|Bartonella vinsonii berkhoffii Ab.IgM|Bartonella vinsonii berkhoffii Ab.IgM
C1954573|T201|COMP|48887-4|LNC|Bartonella vinsonii berkhoffii Ab.IgG|Bartonella vinsonii berkhoffii Ab.IgG
C1954574|T201|COMP|48888-2|LNC|Coxiella burnetii phase 1 Ab.IgG|Coxiella burnetii phase 1 Ab.IgG
C1954575|T201|COMP|48889-0|LNC|Coxiella burnetii phase 1 Ab.IgA|Coxiella burnetii phase 1 Ab.IgA
C1954576|T201|COMP|48890-8|LNC|Coxiella burnetii phase 1 Ab.IgM|Coxiella burnetii phase 1 Ab.IgM
C1954577|T201|COMP|48891-6|LNC|Coxiella burnetii phase 2 Ab.IgA|Coxiella burnetii phase 2 Ab.IgA
C1954578|T201|COMP|48892-4|LNC|Coxiella burnetii phase 2 Ab.IgM|Coxiella burnetii phase 2 Ab.IgM
C1954579|T201|COMP|48893-2|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C1954580|T201|COMP|48894-0|LNC|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C1954581|T201|COMP|48895-7|LNC|Ehrlichia chaffeensis Ab.IgM|Ehrlichia chaffeensis Ab.IgM
C1954582|T201|COMP|48896-5|LNC|Orientia tsutsugamushi Gilliam Ab.IgM|Orientia tsutsugamushi Gilliam Ab.IgM
C1954583|T201|COMP|48897-3|LNC|Orientia tsutsugamushi Gilliam Ab.IgG|Orientia tsutsugamushi Gilliam Ab.IgG
C1954584|T201|COMP|48898-1|LNC|Orientia tsutsugamushi Karp Ab.IgG|Orientia tsutsugamushi Karp Ab.IgG
C1954585|T201|COMP|48899-9|LNC|Orientia tsutsugamushi Karp Ab.IgM|Orientia tsutsugamushi Karp Ab.IgM
C1954586|T201|COMP|48900-5|LNC|Orientia tsutsugamushi Kato Ab.IgG|Orientia tsutsugamushi Kato Ab.IgG
C1954587|T201|COMP|48901-3|LNC|Orientia tsutsugamushi Kato Ab.IgM|Orientia tsutsugamushi Kato Ab.IgM
C1954588|T201|COMP|48902-1|LNC|Rickettsia africae Ab.IgM|Rickettsia africae Ab.IgM
C1954589|T201|COMP|48903-9|LNC|Rickettsia africae Ab.IgG|Rickettsia africae Ab.IgG
C1954590|T201|COMP|48904-7|LNC|Rickettsia akari Ab.IgG|Rickettsia akari Ab.IgG
C1954591|T201|COMP|48905-4|LNC|Rickettsia akari Ab.IgM|Rickettsia akari Ab.IgM
C1954592|T201|COMP|48906-2|LNC|Rickettsia conorii Ab.IgM|Rickettsia conorii Ab.IgM
C1954593|T201|COMP|48907-0|LNC|Rickettsia conorii Ab.IgG|Rickettsia conorii Ab.IgG
C1954594|T201|COMP|48908-8|LNC|Rickettsia parkeri Ab.IgM|Rickettsia parkeri Ab.IgM
C1954595|T201|COMP|48909-6|LNC|Rickettsia parkeri Ab.IgG|Rickettsia parkeri Ab.IgG
C1954596|T201|COMP|48910-4|LNC|Rickettsia prowazekii Ab.IgM|Rickettsia prowazekii Ab.IgM
C1954597|T201|COMP|48911-2|LNC|Rickettsia prowazekii Ab.IgG|Rickettsia prowazekii Ab.IgG
C1954598|T201|COMP|48912-0|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C1954599|T201|COMP|48913-8|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C1954600|T201|COMP|48914-6|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C1954601|T201|COMP|48915-3|LNC|Rickettsia typhi Ab.IgM|Rickettsia typhi Ab.IgM
C1954608|T201|COMP|48919-5|LNC|Respiratory allergen panel, US - Central Florida|Respiratory allergen panel, US - Central Florida
C1954610|T201|COMP|48920-3|LNC|Respiratory allergen panel, US - Southern Florida|Respiratory allergen panel, US - Southern Florida
C1954612|T201|COMP|48921-1|LNC|Respiratory allergen panel, US - Southeast coast|Respiratory allergen panel, US - Southeast coast
C1954634|T201|COMP|48932-8|LNC|Respiratory allergen panel, US - Alaska b|Respiratory allergen panel, US - Alaska b
C1954636|T201|COMP|48933-6|LNC|Respiratory allergen panel, US - Hawaii|Respiratory allergen panel, US - Hawaii
C1954638|T201|COMP|48934-4|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C1954639|T201|COMP|48935-1|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C1954640|T201|COMP|48936-9|LNC|Acylcarnitine pattern|Acylcarnitine pattern
C1954641|T201|COMP|48937-7|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C1954642|T201|COMP|48938-5|LNC|ALPRAZolam|ALPRAZolam
C1954643|T201|COMP|48939-3|LNC|Amphetamines|Amphetamines
C1954644|T201|COMP|48940-1|LNC|Benzodiazepines|Benzodiazepines
C1954645|T201|COMP|48941-9|LNC|Benzodiazepines|Benzodiazepines
C1954646|T201|COMP|48942-7|LNC|Cannabinoids|Cannabinoids
C1954647|T201|COMP|48943-5|LNC|Cannabinoids|Cannabinoids
C1954648|T201|COMP|48944-3|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C1954649|T201|COMP|48945-0|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C1954650|T201|COMP|48946-8|LNC|Cocaethylene|Cocaethylene
C1954651|T201|COMP|48947-6|LNC|Cocaine|Cocaine
C1954652|T201|COMP|48948-4|LNC|diazePAM|diazePAM
C1954653|T201|COMP|48949-2|LNC|Estazolam|Estazolam
C1954654|T201|COMP|48950-0|LNC|Flurazepam|Flurazepam
C1954656|T201|COMP|48952-6|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1954657|T201|COMP|48953-4|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C1954658|T201|COMP|48954-2|LNC|Hydroxytriazolam|Hydroxytriazolam
C1954659|T201|COMP|48955-9|LNC|LORazepam|LORazepam
C1954660|T201|COMP|48956-7|LNC|Methadone|Methadone
C1954661|T201|COMP|48957-5|LNC|Methadone|Methadone
C1954662|T201|COMP|48958-3|LNC|Midazolam|Midazolam
C1954663|T201|COMP|48959-1|LNC|Nordiazepam|Nordiazepam
C1954664|T201|COMP|48960-9|LNC|Norpropoxyphene|Norpropoxyphene
C1954665|T201|COMP|48961-7|LNC|Opiates|Opiates
C1954666|T201|COMP|48962-5|LNC|Oxazepam|Oxazepam
C1954667|T201|COMP|48963-3|LNC|Propoxyphene|Propoxyphene
C1954668|T201|COMP|48964-1|LNC|Propoxyphene|Propoxyphene
C1954669|T201|COMP|48965-8|LNC|Temazepam|Temazepam
C1954670|T201|COMP|48966-6|LNC|Triazolam|Triazolam
C1954671|T201|COMP|48967-4|LNC|Brucella abortus Ab|Brucella abortus Ab
C1954672|T201|COMP|48968-2|LNC|PKHD1 gene targeted mutation analysis|PKHD1 gene targeted mutation analysis
C1954673|T201|COMP|48969-0|LNC|DCX gene targeted mutation analysis|DCX gene targeted mutation analysis
C1954675|T201|COMP|48970-8|LNC|ELN gene targeted mutation analysis|ELN gene targeted mutation analysis
C1954676|T201|COMP|48971-6|LNC|EYA1 gene targeted mutation analysis|EYA1 gene targeted mutation analysis
C1954678|T201|COMP|48972-4|LNC|FGFR2 gene+FGFR3 gene targeted mutation analysis|FGFR2 gene+FGFR3 gene targeted mutation analysis
C1954680|T201|COMP|48973-2|LNC|Leukocytes^2nd specimen|Leukocytes^2nd specimen
C1954681|T201|COMP|48974-0|LNC|MDCR gene targeted mutation analysis|MDCR gene targeted mutation analysis
C1954683|T201|COMP|48975-7|LNC|GPR143 gene targeted mutation analysis|GPR143 gene targeted mutation analysis
C1954685|T201|COMP|48976-5|LNC|POLG gene targeted mutation analysis|POLG gene targeted mutation analysis
C1954687|T201|COMP|48977-3|LNC|SGCG gene targeted mutation analysis|SGCG gene targeted mutation analysis
C1954689|T201|COMP|48978-1|LNC|CDKL5 gene targeted mutation analysis|CDKL5 gene targeted mutation analysis
C1954691|T201|COMP|48979-9|LNC|TSC1 gene targeted mutation analysis|TSC1 gene targeted mutation analysis
C1954693|T201|COMP|48980-7|LNC|TSC2 gene targeted mutation analysis|TSC2 gene targeted mutation analysis
C1954695|T201|COMP|48981-5|LNC|Anaplasma sp|Anaplasma sp
C1954696|T201|COMP|48982-3|LNC|Ehrlichia sp|Ehrlichia sp
C1954697|T201|COMP|48983-1|LNC|Glucose^20M pre XXX challenge|Glucose^20M pre XXX challenge
C1954698|T201|COMP|48991-4|LNC|Glucose^10 PM specimen|Glucose^10 PM specimen
C1954699|T201|COMP|48992-2|LNC|Glucose^12 AM specimen|Glucose^12 AM specimen
C1954700|T201|COMP|48993-0|LNC|Glucose^3 AM specimen|Glucose^3 AM specimen
C1954701|T201|COMP|48994-8|LNC|Glucose^6 AM specimen|Glucose^6 AM specimen
C1954702|T201|COMP|48995-5|LNC|N-acetyl-beta-glucosaminidase/Creatinine|N-acetyl-beta-glucosaminidase/Creatinine
C1954704|T201|COMP|48996-3|LNC|Amylase.pancreatic|Amylase.pancreatic
C1954705|T201|COMP|48997-1|LNC|Immune complex.IgG|Immune complex.IgG
C1954706|T201|COMP|48998-9|LNC|6-Phosphogluconate dehydrogenase|6-Phosphogluconate dehydrogenase
C1954707|T201|COMP|48999-7|LNC|Urea|Urea
C1954708|T201|COMP|49000-3|LNC|Hemoglobin.free|Hemoglobin.free
C1954709|T201|COMP|49001-1|LNC|Osmolality|Osmolality
C1954710|T201|COMP|49002-9|LNC|Albumin|Albumin
C1954711|T201|COMP|49003-7|LNC|Urate|Urate
C1954712|T201|COMP|49004-5|LNC|Creatinine|Creatinine
C1954713|T201|COMP|49005-2|LNC|Calcium|Calcium
C1954714|T201|COMP|49006-0|LNC|Phosphate|Phosphate
C1954715|T201|COMP|49007-8|LNC|Magnesium|Magnesium
C1954716|T201|COMP|49008-6|LNC|Coagulum retraction|Coagulum retraction
C1954717|T201|COMP|49009-4|LNC|Norepinephrine^7th specimen post XXX challenge|Norepinephrine^7th specimen post XXX challenge
C1954719|T201|COMP|49011-0|LNC|Platelet aggregation.arachidonate induced|Platelet aggregation.arachidonate induced
C1954720|T201|COMP|49012-8|LNC|Influenza virus A & B identified|Influenza virus A & B identified
C1954722|T201|COMP|49013-6|LNC|Pancreastatin|Pancreastatin
C1954723|T201|COMP|49014-4|LNC|PAH gene targeted mutation analysis|PAH gene targeted mutation analysis
C1954725|T201|COMP|49015-1|LNC|SCA15 gene.CAG repeats|SCA15 gene.CAG repeats
C1954727|T201|COMP|49016-9|LNC|Streptococcus sp exoenzyme Ab|Streptococcus sp exoenzyme Ab
C1954733|T201|COMP|49019-3|LNC|Respiratory allergen panel, US - Puerto Rico|Respiratory allergen panel, US - Puerto Rico
C1954741|T201|COMP|49023-5|LNC|Albumin|Albumin
C1954742|T201|COMP|49024-3|LNC|Differential cell count method|Differential cell count method
C1954744|T201|COMP|49025-0|LNC|Cells.CD25+CD127Low/Cells.CD4|Cells.CD25+CD127Low/Cells.CD4
C1954746|T201|COMP|49026-8|LNC|LDL 6|LDL 6
C1954748|T201|COMP|49027-6|LNC|LDL 7|LDL 7
C1954750|T201|COMP|49028-4|LNC|Microdeletion syndromes|Microdeletion syndromes
C1954752|T201|COMP|49029-2|LNC|Cortisol.free/Cortisone.free|Cortisol.free/Cortisone.free
C1954756|T201|COMP|49031-8|LNC|Erythrocytes.CD59/100 erythrocytes|Erythrocytes.CD59/100 erythrocytes
C1954758|T201|COMP|49032-6|LNC|Second trimester penta maternal screen|Second trimester penta maternal screen
C1954762|T201|COMP|49034-2|LNC|Microorganism identified|Microorganism identified
C1954765|T201|COMP|49036-7|LNC|Parathyrin.intact^post excision|Parathyrin.intact^post excision
C1954766|T201|COMP|49037-5|LNC|Respiratory syncytial virus Ab.IgG & IgM panel|Respiratory syncytial virus Ab.IgG & IgM panel
C1954768|T201|COMP|49038-3|LNC|Riboflavin|Riboflavin
C1954769|T201|COMP|49039-1|LNC|Subtelomere analysis|Subtelomere analysis
C1954771|T201|COMP|49040-9|LNC|Subtelomere analysis|Subtelomere analysis
C1954772|T201|COMP|49041-7|LNC|Testosterone|Testosterone
C1954773|T201|COMP|49042-5|LNC|Testosterone.free|Testosterone.free
C1954774|T201|COMP|49043-3|LNC|Testosterone.free/Testosterone.total|Testosterone.free/Testosterone.total
C1954775|T201|COMP|49044-1|LNC|Diazepam & Nordiazepam panel|Diazepam & Nordiazepam panel
C1954777|T201|COMP|49045-8|LNC|PT & aPTT & Fibrinogen panel|PT & aPTT & Fibrinogen panel
C1954779|T201|COMP|49046-6|LNC|Drugs of abuse panel|Drugs of abuse panel
C1954781|T201|COMP|49047-4|LNC|Globulin|Globulin
C1954782|T201|COMP|49048-2|LNC|Protein feed time|Protein feed time
C1954784|T201|COMP|49049-0|LNC|Collection time|Collection time
C1954793|T201|COMP|49054-0|LNC|25-Hydroxycalciferol|25-Hydroxycalciferol
C1954794|T201|COMP|49055-7|LNC|Ribonucleoprotein extractable nuclear 52kD Ab|Ribonucleoprotein extractable nuclear 52kD Ab
C1954796|T201|COMP|49056-5|LNC|Shigella sp serotype|Shigella sp serotype
C1954798|T201|COMP|49057-3|LNC|Blood group antibody score|Blood group antibody score
C1954800|T201|COMP|49058-1|LNC|Coagulation surface induced|Coagulation surface induced
C1954802|T201|COMP|49059-9|LNC|Trisomy 21+Trisomy 18 risk|Trisomy 21+Trisomy 18 risk
C1954804|T201|COMP|49060-7|LNC|Fondaparinux|Fondaparinux
C1954805|T201|COMP|49061-5|LNC|Hepatic iron index|Hepatic iron index
C1954807|T201|COMP|49062-3|LNC|Lipid risk factors|Lipid risk factors
C1954809|T201|COMP|49063-1|LNC|Microdeletion syndromes|Microdeletion syndromes
C1954810|T201|COMP|49064-9|LNC|Gamma 2 globulin|Gamma 2 globulin
C1954812|T201|COMP|49065-6|LNC|Eastern equine encephalitis virus Ab.IgG & IgM|Eastern equine encephalitis virus Ab.IgG & IgM
C1954813|T201|COMP|49066-4|LNC|Western equine encephalitis virus Ab.IgG & IgM|Western equine encephalitis virus Ab.IgG & IgM
C1954815|T201|COMP|49067-2|LNC|La Crosse virus Ab.IgG & IgM|La Crosse virus Ab.IgG & IgM
C1954817|T201|COMP|49068-0|LNC|Saint Louis encephalitis virus Ab.IgG & IgM|Saint Louis encephalitis virus Ab.IgG & IgM
C1954819|T201|COMP|49069-8|LNC|Epstein Barr virus Ab|Epstein Barr virus Ab
C1954820|T201|COMP|49070-6|LNC|Specimen drawn|Specimen drawn
C1954821|T201|COMP|49071-4|LNC|Urea nitrogen^post dialysis/pre dialysis|Urea nitrogen^post dialysis/pre dialysis
C1954822|T201|COMP|49072-2|LNC|Cocaethylene|Cocaethylene
C1954823|T201|COMP|49073-0|LNC|Influenza virus A Ab.IgG|Influenza virus A Ab.IgG
C1954824|T201|COMP|49074-8|LNC|Influenza virus A Ab.IgA|Influenza virus A Ab.IgA
C1954825|T201|COMP|49075-5|LNC|Influenza virus A Ab.IgM|Influenza virus A Ab.IgM
C1954826|T201|COMP|49076-3|LNC|Influenza virus B Ab.IgA|Influenza virus B Ab.IgA
C1954827|T201|COMP|49077-1|LNC|Influenza virus B Ab.IgG|Influenza virus B Ab.IgG
C1954828|T201|COMP|49078-9|LNC|Influenza virus B Ab.IgM|Influenza virus B Ab.IgM
C1954829|T201|COMP|49079-7|LNC|Periplaneta americana Ab.IgE.RAST class|Periplaneta americana Ab.IgE.RAST class
C1954831|T201|COMP|49080-5|LNC|Kanamycin 1.0 ug/mL|Kanamycin 1.0 ug/mL
C1954833|T201|COMP|49081-3|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C1954834|T201|COMP|49082-1|LNC|Western equine encephalitis virus Ab.IgG & IgM|Western equine encephalitis virus Ab.IgG & IgM
C1954843|T201|COMP|49087-0|LNC|Maternal screen clinical predictors panel|Maternal screen clinical predictors panel
C1954849|T201|COMP|49090-4|LNC|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C1954851|T201|COMP|49091-2|LNC|Neural tube defect risk|Neural tube defect risk
C1954853|T201|COMP|49092-0|LNC|Second trimester quad maternal screen|Second trimester quad maternal screen
C1954855|T201|COMP|49093-8|LNC|Arbovirus Ab.IgG & IgM panel|Arbovirus Ab.IgG & IgM panel
C1954857|T201|COMP|49094-6|LNC|Arbovirus Ab.IgG & IgM panel|Arbovirus Ab.IgG & IgM panel
C1954858|T201|COMP|49095-3|LNC|Saint Louis encephalitis virus Ab.IgG & IgM|Saint Louis encephalitis virus Ab.IgG & IgM
C1954859|T201|COMP|49096-1|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1954860|T201|COMP|49097-9|LNC|Creatine|Creatine
C1954861|T201|COMP|49098-7|LNC|Cryptococcus neoformans rRNA|Cryptococcus neoformans rRNA
C1954862|T201|COMP|49099-5|LNC|Gadus morhua Ab.IgG|Gadus morhua Ab.IgG
C1954863|T201|COMP|49100-1|LNC|H2a-H2b DNA Ab.IgG|H2a-H2b DNA Ab.IgG
C1954864|T201|COMP|49101-9|LNC|Helicobacter pylori DNA|Helicobacter pylori DNA
C1954866|T201|COMP|49102-7|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1954867|T201|COMP|49103-5|LNC|Leukocyte casts|Leukocyte casts
C1954868|T201|COMP|49104-3|LNC|Mycoplasma pneumoniae DNA|Mycoplasma pneumoniae DNA
C1954869|T201|COMP|49105-0|LNC|Phenolphthalein|Phenolphthalein
C1954870|T201|COMP|49106-8|LNC|Phenols|Phenols
C1954871|T201|COMP|49107-6|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C1954872|T201|COMP|49108-4|LNC|Titanium|Titanium
C1954873|T201|COMP|49109-2|LNC|Toxoplasma gondii Ab|Toxoplasma gondii Ab
C1954875|T201|COMP|49119-1|LNC|Monosaccharides.sulfated|Monosaccharides.sulfated
C1954877|T201|COMP|49120-9|LNC|Immunodeficiency follow-up panel|Immunodeficiency follow-up panel
C1954879|T201|COMP|49121-7|LNC|Erythrocyte inclusion bodies|Erythrocyte inclusion bodies
C1954881|T201|COMP|49122-5|LNC|Anaplasma sp identified|Anaplasma sp identified
C1954882|T201|COMP|49123-3|LNC|Bartonella sp identified|Bartonella sp identified
C1954883|T201|COMP|49124-1|LNC|Coxiella burnetii identified|Coxiella burnetii identified
C1954885|T201|COMP|49125-8|LNC|Ehrlichia sp identified|Ehrlichia sp identified
C1954886|T201|COMP|49126-6|LNC|Orientia tsutsugamushi identified|Orientia tsutsugamushi identified
C1954888|T201|COMP|49127-4|LNC|Rickettsia sp identified|Rickettsia sp identified
C1954889|T201|COMP|49128-2|LNC|Rickettsia typhus group identified|Rickettsia typhus group identified
C1954891|T201|COMP|49129-0|LNC|Creatine kinase.MiMi/Creatine kinase.total|Creatine kinase.MiMi/Creatine kinase.total
C1954893|T201|COMP|49130-8|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C1954894|T201|COMP|49131-6|LNC|Chylomicrons/Lipoprotein.total|Chylomicrons/Lipoprotein.total
C1954896|T201|COMP|49132-4|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C1954897|T201|COMP|49133-2|LNC|Cholesterol.in VLDL|Cholesterol.in VLDL
C1954898|T201|COMP|49134-0|LNC|Glucose^2H post dose glucose|Glucose^2H post dose glucose
C1954899|T201|COMP|49135-7|LNC|Fractional excretion of sodium|Fractional excretion of sodium
C1954900|T201|COMP|49136-5|LNC|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C1954901|T201|COMP|49137-3|LNC|Hemoglobin|Hemoglobin
C1954902|T201|COMP|49138-1|LNC|California encephalitis virus Ab.IgG|California encephalitis virus Ab.IgG
C1954903|T201|COMP|49139-9|LNC|California encephalitis virus Ab.IgM|California encephalitis virus Ab.IgM
C1954904|T201|COMP|49140-7|LNC|California encephalitis virus Ab.IgG|California encephalitis virus Ab.IgG
C1954905|T201|COMP|49141-5|LNC|California encephalitis virus Ab.IgM|California encephalitis virus Ab.IgM
C1954906|T201|COMP|49142-3|LNC|La Crosse virus Ab.IgG & IgM|La Crosse virus Ab.IgG & IgM
C1954909|T201|COMP|49144-9|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C1954910|T201|COMP|49145-6|LNC|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C1954911|T201|COMP|49146-4|LNC|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C1954912|T201|COMP|49147-2|LNC|Rickettsia prowazekii Ab.IgM|Rickettsia prowazekii Ab.IgM
C1954913|T201|COMP|49148-0|LNC|Rickettsia prowazekii Ab.IgG|Rickettsia prowazekii Ab.IgG
C1954914|T201|COMP|49149-8|LNC|Rickettsia parkeri Ab.IgG|Rickettsia parkeri Ab.IgG
C1954915|T201|COMP|49150-6|LNC|Rickettsia parkeri Ab.IgM|Rickettsia parkeri Ab.IgM
C1954916|T201|COMP|49151-4|LNC|Rickettsia parkeri Ab.IgG|Rickettsia parkeri Ab.IgG
C1954917|T201|COMP|49152-2|LNC|Rickettsia parkeri Ab.IgM|Rickettsia parkeri Ab.IgM
C1954918|T201|COMP|49153-0|LNC|Rickettsia conorii Ab.IgM|Rickettsia conorii Ab.IgM
C1954919|T201|COMP|49154-8|LNC|Rickettsia conorii Ab.IgG|Rickettsia conorii Ab.IgG
C1954920|T201|COMP|49155-5|LNC|Rickettsia akari Ab.IgM|Rickettsia akari Ab.IgM
C1954921|T201|COMP|49156-3|LNC|Rickettsia akari Ab.IgM|Rickettsia akari Ab.IgM
C1954922|T201|COMP|49157-1|LNC|Rickettsia akari Ab.IgG|Rickettsia akari Ab.IgG
C1954923|T201|COMP|49158-9|LNC|Rickettsia akari Ab.IgG|Rickettsia akari Ab.IgG
C1954924|T201|COMP|49159-7|LNC|Rickettsia africae Ab.IgG|Rickettsia africae Ab.IgG
C1954925|T201|COMP|49160-5|LNC|Rickettsia africae Ab.IgM|Rickettsia africae Ab.IgM
C1954926|T201|COMP|49161-3|LNC|Rickettsia africae Ab.IgG|Rickettsia africae Ab.IgG
C1954927|T201|COMP|49162-1|LNC|Rickettsia africae Ab.IgM|Rickettsia africae Ab.IgM
C1954928|T201|COMP|49163-9|LNC|Orientia tsutsugamushi Kato Ab.IgM|Orientia tsutsugamushi Kato Ab.IgM
C1954929|T201|COMP|49164-7|LNC|Orientia tsutsugamushi Kato Ab.IgM|Orientia tsutsugamushi Kato Ab.IgM
C1954930|T201|COMP|49165-4|LNC|Orientia tsutsugamushi Kato Ab.IgG|Orientia tsutsugamushi Kato Ab.IgG
C1954931|T201|COMP|49166-2|LNC|Orientia tsutsugamushi Kato Ab.IgG|Orientia tsutsugamushi Kato Ab.IgG
C1954932|T201|COMP|49167-0|LNC|Orientia tsutsugamushi Karp Ab.IgM|Orientia tsutsugamushi Karp Ab.IgM
C1954933|T201|COMP|49168-8|LNC|Orientia tsutsugamushi Karp Ab.IgM|Orientia tsutsugamushi Karp Ab.IgM
C1954934|T201|COMP|49169-6|LNC|Orientia tsutsugamushi Karp Ab.IgG|Orientia tsutsugamushi Karp Ab.IgG
C1954935|T201|COMP|49170-4|LNC|Orientia tsutsugamushi Karp Ab.IgG|Orientia tsutsugamushi Karp Ab.IgG
C1954936|T201|COMP|49171-2|LNC|Orientia tsutsugamushi Gilliam Ab.IgM|Orientia tsutsugamushi Gilliam Ab.IgM
C1954937|T201|COMP|49172-0|LNC|Orientia tsutsugamushi Gilliam Ab.IgM|Orientia tsutsugamushi Gilliam Ab.IgM
C1954938|T201|COMP|49173-8|LNC|Orientia tsutsugamushi Gilliam Ab.IgG|Orientia tsutsugamushi Gilliam Ab.IgG
C1954939|T201|COMP|49174-6|LNC|Orientia tsutsugamushi Gilliam Ab.IgG|Orientia tsutsugamushi Gilliam Ab.IgG
C1954940|T201|COMP|49175-3|LNC|Human bocavirus Ab.IgG|Human bocavirus Ab.IgG
C1954941|T201|COMP|49176-1|LNC|Herpes virus 8 Ab.IgM|Herpes virus 8 Ab.IgM
C1954942|T201|COMP|49177-9|LNC|Hepatitis B virus surface Ab.IgG|Hepatitis B virus surface Ab.IgG
C1954943|T201|COMP|49178-7|LNC|Epstein Barr virus Ab|Epstein Barr virus Ab
C1954944|T201|COMP|49179-5|LNC|Ehrlichia chaffeensis Ab.IgM|Ehrlichia chaffeensis Ab.IgM
C1954945|T201|COMP|49180-3|LNC|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C1954946|T201|COMP|49181-1|LNC|Echinococcus granulosus Ab|Echinococcus granulosus Ab
C1954947|T201|COMP|49182-9|LNC|Coxiella burnetii phase 2 Ab.IgM|Coxiella burnetii phase 2 Ab.IgM
C1954948|T201|COMP|49183-7|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C1954949|T201|COMP|49184-5|LNC|Coxiella burnetii phase 2 Ab.IgA|Coxiella burnetii phase 2 Ab.IgA
C1954950|T201|COMP|49185-2|LNC|Coxiella burnetii phase 1 Ab.IgM|Coxiella burnetii phase 1 Ab.IgM
C1954951|T201|COMP|49186-0|LNC|Coxiella burnetii phase 1 Ab.IgG|Coxiella burnetii phase 1 Ab.IgG
C1954952|T201|COMP|49187-8|LNC|Coxiella burnetii phase 1 Ab.IgA|Coxiella burnetii phase 1 Ab.IgA
C1954953|T201|COMP|49188-6|LNC|Corynebacterium diphtheriae toxin Ab^2nd specimen|Corynebacterium diphtheriae toxin Ab^2nd specimen
C1954954|T201|COMP|49189-4|LNC|Corynebacterium diphtheriae toxin Ab.IgG|Corynebacterium diphtheriae toxin Ab.IgG
C1954955|T201|COMP|49190-2|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1954956|T201|COMP|49191-0|LNC|Clostridium tetani toxoid Ab.IgG^1st specimen|Clostridium tetani toxoid Ab.IgG^1st specimen
C1954957|T201|COMP|49192-8|LNC|Clostridium tetani toxoid Ab.IgG^2nd specimen|Clostridium tetani toxoid Ab.IgG^2nd specimen
C1954958|T201|COMP|49193-6|LNC|California encephalitis virus Ab.IgM|California encephalitis virus Ab.IgM
C1954959|T201|COMP|49194-4|LNC|California encephalitis virus Ab.IgG|California encephalitis virus Ab.IgG
C1954960|T201|COMP|49195-1|LNC|California encephalitis virus Ab.IgG|California encephalitis virus Ab.IgG
C1954961|T201|COMP|49196-9|LNC|Brucella abortus Ab|Brucella abortus Ab
C1954962|T201|COMP|49197-7|LNC|Bartonella vinsonii berkhoffii Ab.IgG|Bartonella vinsonii berkhoffii Ab.IgG
C1954963|T201|COMP|49198-5|LNC|Bartonella vinsonii berkhoffii Ab.IgM|Bartonella vinsonii berkhoffii Ab.IgM
C1954964|T201|COMP|49199-3|LNC|Bartonella vinsonii berkhoffii Ab.IgG|Bartonella vinsonii berkhoffii Ab.IgG
C1954965|T201|COMP|49200-9|LNC|Bartonella vinsonii berkhoffii Ab.IgM|Bartonella vinsonii berkhoffii Ab.IgM
C1954966|T201|COMP|49201-7|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C1954967|T201|COMP|49202-5|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C1954968|T201|COMP|49203-3|LNC|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C1954969|T201|COMP|49204-1|LNC|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C1954970|T201|COMP|49205-8|LNC|Bartonella elizabethae Ab.IgM|Bartonella elizabethae Ab.IgM
C1954971|T201|COMP|49206-6|LNC|Bartonella elizabethae Ab.IgG|Bartonella elizabethae Ab.IgG
C1954972|T201|COMP|49207-4|LNC|Bartonella elizabethae Ab.IgM|Bartonella elizabethae Ab.IgM
C1954973|T201|COMP|49216-5|LNC|Hexokinase|Hexokinase
C1954974|T201|COMP|49217-3|LNC|2,3-Diphosphoglycerate|2,3-Diphosphoglycerate
C1954975|T201|COMP|49218-1|LNC|Phosphatidylinositol/Surfactant.total|Phosphatidylinositol/Surfactant.total
C1954977|T201|COMP|49219-9|LNC|Galactose|Galactose
C1954978|T201|COMP|49220-7|LNC|Prolactin|Prolactin
C1954979|T201|COMP|49221-5|LNC|Catalase|Catalase
C1954980|T201|COMP|49222-3|LNC|Food allergen panel|Food allergen panel
C1954982|T201|COMP|49223-1|LNC|Colony count|Colony count
C1954983|T201|COMP|49224-9|LNC|Leukocytes|Leukocytes
C1954984|T201|COMP|49225-6|LNC|Heptacarboxylate/Creatinine|Heptacarboxylate/Creatinine
C1954985|T201|COMP|49226-4|LNC|lamiVUDine|lamiVUDine
C1954986|T201|COMP|49227-2|LNC|Stavudine|Stavudine
C1954987|T201|COMP|49228-0|LNC|Porphobilinogen deaminase|Porphobilinogen deaminase
C1954988|T201|COMP|49229-8|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C1954989|T201|COMP|49230-6|LNC|Acetylcholinesterase|Acetylcholinesterase
C1954990|T201|COMP|49231-4|LNC|Cholinesterase|Cholinesterase
C1954991|T201|COMP|49232-2|LNC|Giardia lamblia+Cryptosporidium sp Ag|Giardia lamblia+Cryptosporidium sp Ag
C1954992|T201|COMP|49233-0|LNC|Giardia lamblia+Cryptosporidium parvum Ag|Giardia lamblia+Cryptosporidium parvum Ag
C1954993|T201|COMP|49234-8|LNC|Patient symptoms^1.5H post dose lactose PO|Patient symptoms^1.5H post dose lactose PO
C1954994|T201|COMP|49235-5|LNC|Patient symptoms^1H post dose lactose PO|Patient symptoms^1H post dose lactose PO
C1954995|T201|COMP|49236-3|LNC|Patient symptoms^2.5H post dose lactose PO|Patient symptoms^2.5H post dose lactose PO
C1954996|T201|COMP|49237-1|LNC|Patient symptoms^2H post dose lactose PO|Patient symptoms^2H post dose lactose PO
C1954997|T201|COMP|49238-9|LNC|Patient symptoms^30M post dose lactose PO|Patient symptoms^30M post dose lactose PO
C1954998|T201|COMP|49239-7|LNC|Patient symptoms^3H post dose lactose PO|Patient symptoms^3H post dose lactose PO
C1954999|T201|COMP|49240-5|LNC|Patient symptoms^pre dose lactose PO|Patient symptoms^pre dose lactose PO
C1955000|T201|COMP|49241-3|LNC|Xylose absorption|Xylose absorption
C1955001|T201|COMP|49242-1|LNC|Acylcarnitine pattern|Acylcarnitine pattern
C1955002|T201|COMP|49243-9|LNC|Alkaline phosphatase isoenzymes|Alkaline phosphatase isoenzymes
C1955003|T201|COMP|49244-7|LNC|Alpha 1 antitrypsin phenotyping|Alpha 1 antitrypsin phenotyping
C1955004|T201|COMP|49245-4|LNC|Alpha tocopherol & Beta+gamma tocopherol|Alpha tocopherol & Beta+gamma tocopherol
C1955005|T201|COMP|49246-2|LNC|Alpha-1-Fetoprotein interpretation|Alpha-1-Fetoprotein interpretation
C1955006|T201|COMP|49247-0|LNC|Amino acid pattern|Amino acid pattern
C1955007|T201|COMP|49248-8|LNC|Amino acid pattern|Amino acid pattern
C1955008|T201|COMP|49249-6|LNC|Amino acids|Amino acids
C1955009|T201|COMP|49250-4|LNC|Amino acids|Amino acids
C1955010|T201|COMP|49251-2|LNC|Amylase isoenzymes|Amylase isoenzymes
C1955011|T201|COMP|49252-0|LNC|Calculus analysis|Calculus analysis
C1955012|T201|COMP|49253-8|LNC|Beta-N-acetylhexosaminidase A & B|Beta-N-acetylhexosaminidase A & B
C1955013|T201|COMP|49254-6|LNC|Bile acid pattern|Bile acid pattern
C1955014|T201|COMP|49255-3|LNC|Calculus analysis|Calculus analysis
C1955015|T201|COMP|49256-1|LNC|Catecholamines|Catecholamines
C1955016|T201|COMP|49257-9|LNC|Catecholamines|Catecholamines
C1955017|T201|COMP|49258-7|LNC|Creatine kinase isoenzymes|Creatine kinase isoenzymes
C1955018|T201|COMP|49259-5|LNC|Creatine kinase isoenzymes|Creatine kinase isoenzymes
C1955019|T201|COMP|49260-3|LNC|Cryoglobulin IgA & IgG & IgM|Cryoglobulin IgA & IgG & IgM
C1955020|T201|COMP|49261-1|LNC|Cryoproteins|Cryoproteins
C1955021|T201|COMP|49262-9|LNC|Fatty acids pattern|Fatty acids pattern
C1955022|T201|COMP|49263-7|LNC|Fatty acids.very long chain pattern|Fatty acids.very long chain pattern
C1955023|T201|COMP|49264-5|LNC|Folate+Cyanocobalamin|Folate+Cyanocobalamin
C1955024|T201|COMP|49265-2|LNC|Gammopathy|Gammopathy
C1955025|T201|COMP|49266-0|LNC|Glucose-6-Phosphate dehydrogenase phenotype|Glucose-6-Phosphate dehydrogenase phenotype
C1955026|T201|COMP|49267-8|LNC|Glutathione reductase phenotype|Glutathione reductase phenotype
C1955027|T201|COMP|49268-6|LNC|Glycosaminoglycans pattern|Glycosaminoglycans pattern
C1955028|T201|COMP|49269-4|LNC|Homovanillate & Creatinine|Homovanillate & Creatinine
C1955029|T201|COMP|49270-2|LNC|Immunoglobulin light chains|Immunoglobulin light chains
C1955030|T201|COMP|49271-0|LNC|Interpretation|Interpretation
C1955031|T201|COMP|49272-8|LNC|Interpretation|Interpretation
C1955032|T201|COMP|49273-6|LNC|Interpretation|Interpretation
C1955033|T201|COMP|49274-4|LNC|Interpretation|Interpretation
C1955034|T201|COMP|49275-1|LNC|Interpretation|Interpretation
C1955035|T201|COMP|49276-9|LNC|Interpretation|Interpretation
C1955036|T201|COMP|49277-7|LNC|Interpretation|Interpretation
C1955037|T201|COMP|49278-5|LNC|Interpretation|Interpretation
C1955038|T201|COMP|49279-3|LNC|Lactate dehydrogenase isoenzymes|Lactate dehydrogenase isoenzymes
C1955039|T201|COMP|49280-1|LNC|Lipoprotein pattern|Lipoprotein pattern
C1955040|T201|COMP|49281-9|LNC|Lipoprotein pattern|Lipoprotein pattern
C1955041|T201|COMP|49282-7|LNC|Metanephrine & Normetanephrine|Metanephrine & Normetanephrine
C1955042|T201|COMP|49283-5|LNC|Metanephrine & Normetanephrine|Metanephrine & Normetanephrine
C1955043|T201|COMP|49284-3|LNC|Oligosaccharides pattern|Oligosaccharides pattern
C1955044|T201|COMP|49285-0|LNC|Organic acids pattern|Organic acids pattern
C1955045|T201|COMP|49286-8|LNC|Organic acids pattern|Organic acids pattern
C1955046|T201|COMP|49287-6|LNC|Organic acids pattern|Organic acids pattern
C1955047|T201|COMP|49288-4|LNC|Parathyrin|Parathyrin
C1955048|T201|COMP|49289-2|LNC|Porphyrins|Porphyrins
C1955049|T201|COMP|49290-0|LNC|Porphyrins|Porphyrins
C1955050|T201|COMP|49291-8|LNC|Porphyrins|Porphyrins
C1955051|T201|COMP|49292-6|LNC|Porphyrin fractions|Porphyrin fractions
C1955052|T201|COMP|49293-4|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C1955053|T201|COMP|49294-2|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C1955054|T201|COMP|49295-9|LNC|Protein pattern|Protein pattern
C1955055|T201|COMP|49296-7|LNC|Protein pattern|Protein pattern
C1955056|T201|COMP|49297-5|LNC|Protein pattern|Protein pattern
C1955057|T201|COMP|49298-3|LNC|Protein pattern|Protein pattern
C1955058|T201|COMP|49299-1|LNC|Protein pattern|Protein pattern
C1955059|T201|COMP|49300-7|LNC|Protein pattern|Protein pattern
C1955060|T201|COMP|49301-5|LNC|Protein pattern|Protein pattern
C1955061|T201|COMP|49302-3|LNC|Protein pattern|Protein pattern
C1955062|T201|COMP|49303-1|LNC|Amino acid pattern|Amino acid pattern
C1955063|T201|COMP|49304-9|LNC|Uranium dose assessment|Uranium dose assessment
C1955066|T201|COMP|49307-2|LNC|Myocardium Ab pattern|Myocardium Ab pattern
C1955067|T201|COMP|49308-0|LNC|Neutrophil cytoplasmic Ab pattern|Neutrophil cytoplasmic Ab pattern
C1955068|T201|COMP|49309-8|LNC|Nuclear Ab pattern|Nuclear Ab pattern
C1955069|T201|COMP|49310-6|LNC|Nuclear Ab pattern|Nuclear Ab pattern
C1955070|T201|COMP|49311-4|LNC|Nuclear Ab pattern|Nuclear Ab pattern
C1955071|T201|COMP|49312-2|LNC|Acute leukemia markers|Acute leukemia markers
C1955072|T201|COMP|49313-0|LNC|Chronic leukemia markers|Chronic leukemia markers
C1955073|T201|COMP|49314-8|LNC|Immunodeficiency markers|Immunodeficiency markers
C1955074|T201|COMP|49315-5|LNC|Hemolytic disease of newborn screen|Hemolytic disease of newborn screen
C1955075|T201|COMP|49316-3|LNC|Hemoglobin pattern|Hemoglobin pattern
C1955076|T201|COMP|49317-1|LNC|Hemoglobin pattern|Hemoglobin pattern
C1955077|T201|COMP|49318-9|LNC|Alpha-1-Fetoprotein interpretation|Alpha-1-Fetoprotein interpretation
C1955078|T201|COMP|49319-7|LNC|Beta glucosidase activator|Beta glucosidase activator
C1955079|T201|COMP|49320-5|LNC|Beta-N-acetylhexosaminidase.A activator|Beta-N-acetylhexosaminidase.A activator
C1955080|T201|COMP|49321-3|LNC|Cerebroside sulfatase activator|Cerebroside sulfatase activator
C1955081|T201|COMP|49322-1|LNC|Hemoglobin pattern|Hemoglobin pattern
C1955082|T201|COMP|49323-9|LNC|Hemoglobin pattern|Hemoglobin pattern
C1955484|T201|COMP|4257-2|LNC|5-Fluorocytosine|5-Fluorocytosine
C1955485|T201|COMP|17831-9|LNC|5-Fluorocytosine|5-Fluorocytosine
C1955486|T201|COMP|17832-7|LNC|5-Fluorocytosine|5-Fluorocytosine
C1955487|T201|COMP|18925-8|LNC|5-Fluorocytosine|5-Fluorocytosine
C1959619|T201|COMP|10408-3|LNC|little i Ag|little i Ag
C1959623|T201|COMP|10407-5|LNC|little i Ag|little i Ag
C1963619|T201|COMP|40646-2|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C1976776|T201|COMP|49554-9|LNC|Beta F1 Ag|Beta F1 Ag
C1976778|T201|COMP|49555-6|LNC|HLA-A+B+C Ag|HLA-A+B+C Ag
C1976779|T201|COMP|49556-4|LNC|p16INK4a Ag|p16INK4a Ag
C1976781|T201|COMP|49557-2|LNC|PDGFR-beta Ag|PDGFR-beta Ag
C1976783|T201|COMP|49558-0|LNC|TAU 3 Ag|TAU 3 Ag
C1976785|T201|COMP|49559-8|LNC|TAU 4 Ag|TAU 4 Ag
C1976792|T201|COMP|49426-0|LNC|Papova virus SV40 DNA|Papova virus SV40 DNA
C1976794|T201|COMP|49427-8|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1976795|T201|COMP|49428-6|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1976796|T201|COMP|49429-4|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1976797|T201|COMP|49430-2|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1976798|T201|COMP|49431-0|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1976799|T201|COMP|49432-8|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1976800|T201|COMP|49433-6|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1976801|T201|COMP|49726-3|LNC|Endomysium Ab.IgG|Endomysium Ab.IgG
C1976802|T201|COMP|49727-1|LNC|Homocysteine|Homocysteine
C1976803|T201|COMP|49728-9|LNC|Neurokinin A|Neurokinin A
C1976804|T201|COMP|49729-7|LNC|Penicillin G Ab.IgG|Penicillin G Ab.IgG
C1976806|T201|COMP|49730-5|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C1976807|T201|COMP|49731-3|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1976808|T201|COMP|49732-1|LNC|Interleukin 6|Interleukin 6
C1976809|T201|COMP|49733-9|LNC|Interleukin 10|Interleukin 10
C1976810|T201|COMP|49734-7|LNC|11-Dehydro thromboxane beta 2/Creatinine|11-Dehydro thromboxane beta 2/Creatinine
C1976812|T201|COMP|49735-4|LNC|FBN1 gene targeted mutation analysis|FBN1 gene targeted mutation analysis
C1976813|T201|COMP|49736-2|LNC|Clarity|Clarity
C1976814|T201|COMP|49737-0|LNC|Sirolimus|Sirolimus
C1976815|T201|COMP|49738-8|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C1976816|T201|COMP|49739-6|LNC|Apis mellifera Ab.IgG|Apis mellifera Ab.IgG
C1976817|T201|COMP|49740-4|LNC|Dolichovespula arenaria Ab.IgG|Dolichovespula arenaria Ab.IgG
C1976818|T201|COMP|49741-2|LNC|Plasmodium malariae Ab.IgG|Plasmodium malariae Ab.IgG
C1976819|T201|COMP|50518-0|LNC|Prolactin^2nd specimen|Prolactin^2nd specimen
C1976820|T201|COMP|50519-8|LNC|Prolactin^3rd specimen|Prolactin^3rd specimen
C1976821|T201|COMP|50520-6|LNC|Prolactin^4th specimen|Prolactin^4th specimen
C1976822|T201|COMP|50521-4|LNC|Prolactin^5th specimen|Prolactin^5th specimen
C1976823|T201|COMP|50522-2|LNC|Prolactin^6th specimen|Prolactin^6th specimen
C1976824|T201|COMP|50523-0|LNC|Prolactin^7th specimen|Prolactin^7th specimen
C1976825|T201|COMP|50524-8|LNC|Prolactin^8th specimen|Prolactin^8th specimen
C1976826|T201|COMP|50525-5|LNC|Parathyrin.intact^1st specimen|Parathyrin.intact^1st specimen
C1976827|T201|COMP|50526-3|LNC|Parathyrin.intact^2nd specimen|Parathyrin.intact^2nd specimen
C1976828|T201|COMP|50527-1|LNC|Parathyrin.intact^3rd specimen|Parathyrin.intact^3rd specimen
C1976829|T201|COMP|50528-9|LNC|Parathyrin.intact^4th specimen|Parathyrin.intact^4th specimen
C1976830|T201|COMP|50529-7|LNC|Parathyrin.intact^5th specimen|Parathyrin.intact^5th specimen
C1976831|T201|COMP|50530-5|LNC|Parathyrin.intact^6th specimen|Parathyrin.intact^6th specimen
C1976844|T201|COMP|49324-7|LNC|11-Deoxycortisol^2H post dose metyraPONE|11-Deoxycortisol^2H post dose metyraPONE
C1976845|T201|COMP|49325-4|LNC|17-Hydroxypregnenolone^1H post XXX challenge|17-Hydroxypregnenolone^1H post XXX challenge
C1976846|T201|COMP|49326-2|LNC|Aldosterone^2H post XXX challenge|Aldosterone^2H post XXX challenge
C1976847|T201|COMP|49626-5|LNC|Muscle sarcolemma Ab|Muscle sarcolemma Ab
C1976848|T201|COMP|49627-3|LNC|Muscle sarcolemma Ab|Muscle sarcolemma Ab
C1976849|T201|COMP|49628-1|LNC|Remnant lipoprotein|Remnant lipoprotein
C1976851|T201|COMP|49629-9|LNC|Citrulline|Citrulline
C1976852|T201|COMP|49630-7|LNC|Darunavir+Ritonavir|Darunavir+Ritonavir
C1976854|T201|COMP|49631-5|LNC|ATN1 gene allele 1.CAG repeats|ATN1 gene allele 1.CAG repeats
C1976856|T201|COMP|49632-3|LNC|ATN1 gene allele 2.CAG repeats|ATN1 gene allele 2.CAG repeats
C1976858|T201|COMP|49633-1|LNC|Ethanolamine|Ethanolamine
C1976859|T201|COMP|49634-9|LNC|FXN gene allele 1.GAA repeats|FXN gene allele 1.GAA repeats
C1976861|T201|COMP|49635-6|LNC|FXN gene allele 2.GAA repeats|FXN gene allele 2.GAA repeats
C1976863|T201|COMP|49636-4|LNC|Ganglioside GM1 Ab|Ganglioside GM1 Ab
C1976864|T201|COMP|49637-2|LNC|HTT gene allele 1.CAG repeats|HTT gene allele 1.CAG repeats
C1976866|T201|COMP|49638-0|LNC|HTT gene allele 2.CAG repeats|HTT gene allele 2.CAG repeats
C1976868|T201|COMP|49939-2|LNC|Dodecenedioate/Creatinine|Dodecenedioate/Creatinine
C1976870|T201|COMP|49940-0|LNC|Glutamate dehydrogenase|Glutamate dehydrogenase
C1976871|T201|COMP|49941-8|LNC|Sepiapterin|Sepiapterin
C1976872|T201|COMP|49942-6|LNC|Somatotropin^1 AM specimen|Somatotropin^1 AM specimen
C1976873|T201|COMP|49943-4|LNC|Somatotropin^1.30 AM specimen|Somatotropin^1.30 AM specimen
C1976874|T201|COMP|49944-2|LNC|Somatotropin^10 PM specimen|Somatotropin^10 PM specimen
C1976875|T201|COMP|49945-9|LNC|Somatotropin^10.30 PM specimen|Somatotropin^10.30 PM specimen
C1976876|T201|COMP|49946-7|LNC|Somatotropin^11 PM specimen|Somatotropin^11 PM specimen
C1976877|T201|COMP|49947-5|LNC|Somatotropin^11.30 PM specimen|Somatotropin^11.30 PM specimen
C1976878|T201|COMP|49948-3|LNC|Somatotropin^12 PM specimen|Somatotropin^12 PM specimen
C1976879|T201|COMP|49949-1|LNC|Somatotropin^12.30 PM specimen|Somatotropin^12.30 PM specimen
C1976880|T201|COMP|49950-9|LNC|Somatotropin^2 AM specimen|Somatotropin^2 AM specimen
C1976881|T201|COMP|49951-7|LNC|Somatotropin^2.30 AM specimen|Somatotropin^2.30 AM specimen
C1976882|T201|COMP|49952-5|LNC|Somatotropin^3 AM specimen|Somatotropin^3 AM specimen
C1976883|T201|COMP|49953-3|LNC|Somatotropin^3.30 AM specimen|Somatotropin^3.30 AM specimen
C1976884|T201|COMP|50174-2|LNC|Alloisoleucine|Alloisoleucine
C1976885|T201|COMP|50175-9|LNC|Alloisoleucine|Alloisoleucine
C1976886|T201|COMP|50176-7|LNC|Alpha-2-Macroglobulin/Protein.total|Alpha-2-Macroglobulin/Protein.total
C1976888|T201|COMP|50177-5|LNC|Hemicystine|Hemicystine
C1976891|T201|COMP|50186-6|LNC|Wine vinegar Ab.IgE|Wine vinegar Ab.IgE
C1976897|T201|COMP|50189-0|LNC|Neonatal bilirubin panel|Neonatal bilirubin panel
C1976899|T201|COMP|50190-8|LNC|Iron & Iron binding capacity panel|Iron & Iron binding capacity panel
C1976901|T201|COMP|50191-6|LNC|Occult blood panel|Occult blood panel
C1976903|T201|COMP|50192-4|LNC|Cholesterol.in VLDL 1+2+3|Cholesterol.in VLDL 1+2+3
C1976905|T201|COMP|50193-2|LNC|Cholesterol.in LDL.narrow density|Cholesterol.in LDL.narrow density
C1976907|T201|COMP|50194-0|LNC|Cholesterol.in IDL+Cholesterol.in VLDL 3|Cholesterol.in IDL+Cholesterol.in VLDL 3
C1976909|T201|COMP|49452-6|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1976910|T201|COMP|49453-4|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1976911|T201|COMP|49454-2|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1976912|T201|COMP|49455-9|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1976913|T201|COMP|49456-7|LNC|Alpha synuclein Ag|Alpha synuclein Ag
C1976914|T201|COMP|49457-5|LNC|Androgen receptor Ag|Androgen receptor Ag
C1976915|T201|COMP|49458-3|LNC|Annexin 1 Ag|Annexin 1 Ag
C1976916|T201|COMP|49459-1|LNC|Alzheimer precursor protein Ag|Alzheimer precursor protein Ag
C1976918|T201|COMP|49460-9|LNC|Beta catenin Ag|Beta catenin Ag
C1976920|T201|COMP|49461-7|LNC|C4d Ag|C4d Ag
C1976921|T201|COMP|49462-5|LNC|Calponin Ag|Calponin Ag
C1976922|T201|COMP|49463-3|LNC|CD1 Ag|CD1 Ag
C1976923|T201|COMP|49464-1|LNC|CD13 Ag|CD13 Ag
C1976924|T201|COMP|49465-8|LNC|CD14 Ag|CD14 Ag
C1976925|T201|COMP|49466-6|LNC|CD2 Ag|CD2 Ag
C1976926|T201|COMP|49467-4|LNC|CD22 Ag|CD22 Ag
C1976927|T201|COMP|49468-2|LNC|CD27 Ag|CD27 Ag
C1976928|T201|COMP|49469-0|LNC|CD33 Ag|CD33 Ag
C1976929|T201|COMP|49470-8|LNC|CD35 Ag|CD35 Ag
C1976930|T201|COMP|49471-6|LNC|IgG subclass 4 Ag|IgG subclass 4 Ag
C1976932|T201|COMP|49472-4|LNC|Mammaglobin Ag|Mammaglobin Ag
C1976933|T201|COMP|49473-2|LNC|CD123 Ag|CD123 Ag
C1976934|T201|COMP|49474-0|LNC|CD163 Ag|CD163 Ag
C1976935|T201|COMP|49475-7|LNC|CD41-Bf Ag|CD41-Bf Ag
C1976936|T201|COMP|49476-5|LNC|Cyclooxygenase 2 Ag|Cyclooxygenase 2 Ag
C1976937|T201|COMP|49477-3|LNC|CXCL13 Ag|CXCL13 Ag
C1976939|T201|COMP|49478-1|LNC|CXCR5 Ag|CXCR5 Ag
C1976941|T201|COMP|49479-9|LNC|FOXP3 Ag|FOXP3 Ag
C1976945|T201|COMP|49480-7|LNC|Herpes virus 8 latent nuclear Ag|Herpes virus 8 latent nuclear Ag
C1976946|T201|COMP|49481-5|LNC|TCL-1A Ag|TCL-1A Ag
C1976948|T201|COMP|49482-3|LNC|Vascular endothelial growth factor Ag|Vascular endothelial growth factor Ag
C1976950|T201|COMP|49483-1|LNC|HIV 1|HIV 1
C1976951|T201|COMP|49688-5|LNC|Glucose tolerance^post 75 g glucose PO|Glucose tolerance^post 75 g glucose PO
C1976952|T201|COMP|49689-3|LNC|Glucose tolerance^post 100 g glucose PO|Glucose tolerance^post 100 g glucose PO
C1976953|T201|COMP|49690-1|LNC|Mirtazapine|Mirtazapine
C1976954|T201|COMP|49691-9|LNC|Nortrimipramine|Nortrimipramine
C1976955|T201|COMP|49692-7|LNC|Striated muscle Ab.IgG|Striated muscle Ab.IgG
C1976956|T201|COMP|49693-5|LNC|Hepatitis E virus Ab.IgG|Hepatitis E virus Ab.IgG
C1976959|T201|COMP|49696-8|LNC|Oxygen^^adjusted to patient's actual temperature|Oxygen^^adjusted to patient's actual temperature
C1976960|T201|COMP|49697-6|LNC|Oxygen^^adjusted to patient's actual temperature|Oxygen^^adjusted to patient's actual temperature
C1976961|T201|COMP|49698-4|LNC|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1976962|T201|COMP|49699-2|LNC|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1976963|T201|COMP|49700-8|LNC|Metanephrine.free|Metanephrine.free
C1976964|T201|COMP|49836-0|LNC|Platelet function|Platelet function
C1976967|T201|COMP|49838-6|LNC|Neural tube defect risk|Neural tube defect risk
C1976968|T201|COMP|49839-4|LNC|Eosinophils|Eosinophils
C1976969|T201|COMP|49840-2|LNC|Cells.CD19+IgG+/100 cells|Cells.CD19+IgG+/100 cells
C1976971|T201|COMP|49841-0|LNC|Cells.CD19+IgM+/100 cells|Cells.CD19+IgM+/100 cells
C1976973|T201|COMP|49842-8|LNC|Cells.CD19+IgA+/100 cells|Cells.CD19+IgA+/100 cells
C1976978|T201|COMP|49846-9|LNC|Hepatitis C virus core Ag|Hepatitis C virus core Ag
C1976979|T201|COMP|49847-7|LNC|Enterovirus RNA|Enterovirus RNA
C1976980|T201|COMP|49848-5|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C1976981|T201|COMP|49849-3|LNC|Hydroxylysine.free/Creatinine|Hydroxylysine.free/Creatinine
C1976983|T201|COMP|49850-1|LNC|Insulin-like growth factor-I^baseline|Insulin-like growth factor-I^baseline
C1976984|T201|COMP|50025-6|LNC|Volatiles panel|Volatiles panel
C1976985|T201|COMP|50036-3|LNC|Dengue virus Ab|Dengue virus Ab
C1976986|T201|COMP|50037-1|LNC|Powassan virus Ab|Powassan virus Ab
C1976987|T201|COMP|50038-9|LNC|Snowshoe hare virus Ab|Snowshoe hare virus Ab
C1976988|T201|COMP|50039-7|LNC|5-Methyltetrahydrofolate/Folate|5-Methyltetrahydrofolate/Folate
C1976990|T201|COMP|50040-5|LNC|Advanced oxidation protein products|Advanced oxidation protein products
C1976992|T201|COMP|50041-3|LNC|Bilirubin+Urobilinogen|Bilirubin+Urobilinogen
C1976994|T201|COMP|50042-1|LNC|Basal metabolic rate index|Basal metabolic rate index
C1976996|T201|COMP|50043-9|LNC|Protein carbonyl/protein|Protein carbonyl/protein
C1976999|T201|COMP|50045-4|LNC|Hemicystine|Hemicystine
C1977000|T201|COMP|50046-2|LNC|Hemicystine|Hemicystine
C1977001|T201|COMP|50047-0|LNC|Hemicystine|Hemicystine
C1977002|T201|COMP|50048-8|LNC|Hemicystine|Hemicystine
C1977003|T201|COMP|50049-6|LNC|Hemicystine/Amino acids.total|Hemicystine/Amino acids.total
C1977005|T201|COMP|49767-7|LNC|Filaria Ab.IgG2|Filaria Ab.IgG2
C1977007|T201|COMP|49768-5|LNC|Filaria Ab.IgG3|Filaria Ab.IgG3
C1977009|T201|COMP|49769-3|LNC|Filaria Ab.IgG4|Filaria Ab.IgG4
C1977010|T201|COMP|49770-1|LNC|Filaria Ab.IgG1|Filaria Ab.IgG1
C1977012|T201|COMP|49771-9|LNC|Onchocerca sp Ab.IgG|Onchocerca sp Ab.IgG
C1977014|T201|COMP|49772-7|LNC|Fructose|Fructose
C1977015|T201|COMP|49773-5|LNC|Galactitol|Galactitol
C1977016|T201|COMP|49774-3|LNC|Glomerular basement membrane Ab|Glomerular basement membrane Ab
C1977017|T201|COMP|49853-5|LNC|Transforming growth factor beta 1|Transforming growth factor beta 1
C1977020|T201|COMP|49855-0|LNC|Tetracycline Ab.IgE|Tetracycline Ab.IgE
C1977022|T201|COMP|49856-8|LNC|methylTESTOSTERone|methylTESTOSTERone
C1977023|T201|COMP|49857-6|LNC|SMN1 gene+SMN2 gene targeted mutation analysis|SMN1 gene+SMN2 gene targeted mutation analysis
C1977025|T201|COMP|49858-4|LNC|Peptide YY|Peptide YY
C1977026|T201|COMP|49859-2|LNC|Amphotericin B|Amphotericin B
C1977029|T201|COMP|50027-2|LNC|Narcissus sp Ab.IgE|Narcissus sp Ab.IgE
C1977031|T201|COMP|50028-0|LNC|Escherichia coli Ab.IgE|Escherichia coli Ab.IgE
C1977033|T201|COMP|50029-8|LNC|Mahogany wood dust Ab.IgE|Mahogany wood dust Ab.IgE
C1977035|T201|COMP|50030-6|LNC|Oak wood dust Ab.IgE|Oak wood dust Ab.IgE
C1977037|T201|COMP|50031-4|LNC|Sulfamethoxazole Ab.IgE|Sulfamethoxazole Ab.IgE
C1977038|T201|COMP|50032-2|LNC|Callistephus chinesi Ab.IgE|Callistephus chinesi Ab.IgE
C1977040|T201|COMP|50033-0|LNC|Cephalosporin Ab.IgE|Cephalosporin Ab.IgE
C1977042|T201|COMP|50034-8|LNC|Arbovirus Ab|Arbovirus Ab
C1977043|T201|COMP|50035-5|LNC|Colorado tick fever virus Ab|Colorado tick fever virus Ab
C1977044|T201|COMP|50179-1|LNC|Calcitonin Calcium & Pentagastrin challenge panel|Calcitonin Calcium & Pentagastrin challenge panel
C1977051|T201|COMP|50185-8|LNC|Magnolia grandiflora Ab.IgE|Magnolia grandiflora Ab.IgE
C1977053|T201|COMP|50694-9|LNC|Rubella virus Ab|Rubella virus Ab
C1977054|T201|COMP|50695-6|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1977055|T201|COMP|50696-4|LNC|Influenza virus A Ab|Influenza virus A Ab
C1977056|T201|COMP|50697-2|LNC|Influenza virus A Ag|Influenza virus A Ag
C1977057|T201|COMP|50698-0|LNC|Influenza virus A.adamantane resistance|Influenza virus A.adamantane resistance
C1977059|T201|COMP|50699-8|LNC|Influenza virus A.adamantane resistance|Influenza virus A.adamantane resistance
C1977060|T201|COMP|50700-4|LNC|Influenza virus A.adamantane resistant RNA|Influenza virus A.adamantane resistant RNA
C1977062|T201|COMP|50701-2|LNC|Influenza virus A H1 Ag|Influenza virus A H1 Ag
C1977064|T201|COMP|50702-0|LNC|Influenza virus A matrix protein RNA|Influenza virus A matrix protein RNA
C1977066|T201|COMP|49577-0|LNC|Lecithin/Surfactant.total|Lecithin/Surfactant.total
C1977068|T201|COMP|49578-8|LNC|Aminocaproate cutoff|Aminocaproate cutoff
C1977070|T201|COMP|49579-6|LNC|Aminocaproate|Aminocaproate
C1977071|T201|COMP|49580-4|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C1977072|T201|COMP|49581-2|LNC|Reference lab test identifier and name|Reference lab test identifier and name
C1977074|T201|COMP|49582-0|LNC|Trisomy 18 risk cutoff|Trisomy 18 risk cutoff
C1977076|T201|COMP|49583-8|LNC|Trisomy 21 risk cutoff|Trisomy 21 risk cutoff
C1977078|T201|COMP|49584-6|LNC|Neural tube defect risk cutoff|Neural tube defect risk cutoff
C1977080|T201|COMP|49639-8|LNC|Protein C/Coagulation factor X|Protein C/Coagulation factor X
C1977082|T201|COMP|49640-6|LNC|Protein S Ag/Coagulation factor X Ag|Protein S Ag/Coagulation factor X Ag
C1977084|T201|COMP|49641-4|LNC|SCA1 gene allele 1.CAG repeats|SCA1 gene allele 1.CAG repeats
C1977085|T201|COMP|49642-2|LNC|SCA1 gene allele 2.CAG repeats|SCA1 gene allele 2.CAG repeats
C1977086|T201|COMP|49643-0|LNC|SCA10 gene allele 1.ATTCT repeats|SCA10 gene allele 1.ATTCT repeats
C1977088|T201|COMP|49644-8|LNC|SCA10 gene allele 2.ATTCT repeats|SCA10 gene allele 2.ATTCT repeats
C1977090|T201|COMP|49645-5|LNC|SCA2 gene allele 1.CAG repeats|SCA2 gene allele 1.CAG repeats
C1977091|T201|COMP|49709-9|LNC|predniSONE|predniSONE
C1977092|T201|COMP|49710-7|LNC|SOD1 gene targeted mutation analysis|SOD1 gene targeted mutation analysis
C1977094|T201|COMP|49711-5|LNC|Listeria sp Ab|Listeria sp Ab
C1977095|T201|COMP|49712-3|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C1977096|T201|COMP|49713-1|LNC|Parainfluenza virus Ab|Parainfluenza virus Ab
C1977097|T201|COMP|49714-9|LNC|Interleukin 8|Interleukin 8
C1977098|T201|COMP|49715-6|LNC|Musca domestica Ab.IgE|Musca domestica Ab.IgE
C1977100|T201|COMP|49716-4|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C1977101|T201|COMP|49717-2|LNC|Interleukin 1 beta|Interleukin 1 beta
C1977102|T201|COMP|49790-9|LNC|Sodium|Sodium
C1977103|T201|COMP|49791-7|LNC|Sodium|Sodium
C1977104|T201|COMP|49792-5|LNC|Somatostatin|Somatostatin
C1977111|T201|COMP|49327-0|LNC|Androstenedione^1H post XXX challenge|Androstenedione^1H post XXX challenge
C1977112|T201|COMP|49328-8|LNC|Clavulanate Ab.IgE|Clavulanate Ab.IgE
C1977114|T201|COMP|49329-6|LNC|Interferon.alpha Ab|Interferon.alpha Ab
C1977116|T201|COMP|49330-4|LNC|Renin^3H post XXX challenge|Renin^3H post XXX challenge
C1977117|T201|COMP|49331-2|LNC|Renin^2H post XXX challenge|Renin^2H post XXX challenge
C1977118|T201|COMP|49332-0|LNC|Vasopressin^30M post XXX challenge|Vasopressin^30M post XXX challenge
C1977119|T201|COMP|49333-8|LNC|Galactitol|Galactitol
C1977120|T201|COMP|49334-6|LNC|Adenovirus DNA|Adenovirus DNA
C1977121|T201|COMP|49335-3|LNC|Adenovirus DNA|Adenovirus DNA
C1977122|T201|COMP|49336-1|LNC|Adenovirus DNA|Adenovirus DNA
C1977123|T201|COMP|49337-9|LNC|Adenovirus DNA|Adenovirus DNA
C1977124|T201|COMP|49338-7|LNC|Adenovirus DNA|Adenovirus DNA
C1977125|T201|COMP|49339-5|LNC|Adenovirus DNA|Adenovirus DNA
C1977126|T201|COMP|49340-3|LNC|Adenovirus DNA|Adenovirus DNA
C1977127|T201|COMP|49341-1|LNC|Adenovirus DNA|Adenovirus DNA
C1977128|T201|COMP|49342-9|LNC|BK virus DNA|BK virus DNA
C1977129|T201|COMP|49343-7|LNC|BK virus DNA|BK virus DNA
C1977130|T201|COMP|49344-5|LNC|BK virus DNA|BK virus DNA
C1977131|T201|COMP|49345-2|LNC|BK virus DNA|BK virus DNA
C1977132|T201|COMP|49346-0|LNC|BK virus DNA|BK virus DNA
C1977133|T201|COMP|49347-8|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1977134|T201|COMP|49348-6|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1977135|T201|COMP|49349-4|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1977136|T201|COMP|49350-2|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1977137|T201|COMP|49351-0|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C1977138|T201|COMP|49352-8|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1977139|T201|COMP|49353-6|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1977140|T201|COMP|49354-4|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1977141|T201|COMP|49355-1|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1977142|T201|COMP|49356-9|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C1977143|T201|COMP|49357-7|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977144|T201|COMP|49358-5|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977145|T201|COMP|49359-3|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977146|T201|COMP|49360-1|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977147|T201|COMP|49361-9|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977148|T201|COMP|49362-7|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977149|T201|COMP|49363-5|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977150|T201|COMP|49364-3|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977151|T201|COMP|49365-0|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977152|T201|COMP|49366-8|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977153|T201|COMP|49367-6|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977154|T201|COMP|49368-4|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977155|T201|COMP|49369-2|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977156|T201|COMP|49370-0|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977157|T201|COMP|49371-8|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977158|T201|COMP|49372-6|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977159|T201|COMP|49373-4|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977160|T201|COMP|49374-2|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977161|T201|COMP|49375-9|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977162|T201|COMP|49376-7|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977163|T201|COMP|49377-5|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977164|T201|COMP|49378-3|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977165|T201|COMP|49379-1|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977166|T201|COMP|49380-9|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977167|T201|COMP|49381-7|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1977168|T201|COMP|49382-5|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1977169|T201|COMP|49383-3|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1977170|T201|COMP|49384-1|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1977171|T201|COMP|49385-8|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1977172|T201|COMP|49386-6|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C1977173|T201|COMP|49387-4|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1977174|T201|COMP|49388-2|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1977175|T201|COMP|49389-0|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1977176|T201|COMP|49390-8|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1977177|T201|COMP|49391-6|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1977178|T201|COMP|49392-4|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1977179|T201|COMP|49393-2|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C1977180|T201|COMP|49394-0|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C1977181|T201|COMP|49395-7|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C1977182|T201|COMP|49396-5|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C1977183|T201|COMP|49397-3|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C1977184|T201|COMP|49398-1|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C1977185|T201|COMP|49399-9|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C1977186|T201|COMP|49400-5|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C1977187|T201|COMP|49401-3|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C1977188|T201|COMP|49402-1|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1977189|T201|COMP|49403-9|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1977190|T201|COMP|49404-7|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1977191|T201|COMP|49405-4|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1977192|T201|COMP|49406-2|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1977193|T201|COMP|49407-0|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1977194|T201|COMP|49408-8|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1977195|T201|COMP|49409-6|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C1977196|T201|COMP|49410-4|LNC|JC virus DNA|JC virus DNA
C1977197|T201|COMP|49411-2|LNC|JC virus DNA|JC virus DNA
C1977198|T201|COMP|49412-0|LNC|JC virus DNA|JC virus DNA
C1977199|T201|COMP|49413-8|LNC|JC virus DNA|JC virus DNA
C1977200|T201|COMP|49414-6|LNC|JC virus DNA|JC virus DNA
C1977201|T201|COMP|49415-3|LNC|JC virus DNA|JC virus DNA
C1977202|T201|COMP|49416-1|LNC|JC virus DNA|JC virus DNA
C1977203|T201|COMP|49417-9|LNC|JC virus DNA|JC virus DNA
C1977204|T201|COMP|49418-7|LNC|Papova virus SV40 DNA|Papova virus SV40 DNA
C1977205|T201|COMP|49419-5|LNC|Papova virus SV40 DNA|Papova virus SV40 DNA
C1977206|T201|COMP|49420-3|LNC|Papova virus SV40 DNA|Papova virus SV40 DNA
C1977207|T201|COMP|49421-1|LNC|Papova virus SV40 DNA|Papova virus SV40 DNA
C1977208|T201|COMP|49422-9|LNC|Papova virus SV40 DNA|Papova virus SV40 DNA
C1977209|T201|COMP|49423-7|LNC|Papova virus SV40 DNA|Papova virus SV40 DNA
C1977210|T201|COMP|49424-5|LNC|Papova virus SV40 DNA|Papova virus SV40 DNA
C1977211|T201|COMP|49425-2|LNC|Papova virus SV40 DNA|Papova virus SV40 DNA
C1977212|T201|COMP|49434-4|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1977213|T201|COMP|49435-1|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1977214|T201|COMP|49436-9|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C1977215|T201|COMP|49437-7|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C1977216|T201|COMP|49438-5|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C1977217|T201|COMP|49439-3|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C1977218|T201|COMP|49440-1|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C1977219|T201|COMP|49441-9|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C1977220|T201|COMP|49442-7|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C1977221|T201|COMP|49443-5|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1977222|T201|COMP|49444-3|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1977223|T201|COMP|49445-0|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1977224|T201|COMP|49446-8|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1977225|T201|COMP|49447-6|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1977226|T201|COMP|49448-4|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1977227|T201|COMP|49449-2|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C1977228|T201|COMP|49450-0|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1977229|T201|COMP|49451-8|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C1977230|T201|COMP|49484-9|LNC|Phenylalanine|Phenylalanine
C1977232|T201|COMP|49486-4|LNC|Alphapinene|Alphapinene
C1977233|T201|COMP|49487-2|LNC|Nateglinide|Nateglinide
C1977234|T201|COMP|49488-0|LNC|Collection time|Collection time
C1977237|T201|COMP|49490-6|LNC|BCR-ABL1 b2a2 fusion protein|BCR-ABL1 b2a2 fusion protein
C1977238|T201|COMP|49491-4|LNC|BCR-ABL1 b3a2 fusion protein|BCR-ABL1 b3a2 fusion protein
C1977239|T201|COMP|49492-2|LNC|Leukemia markers|Leukemia markers
C1977240|T201|COMP|49493-0|LNC|Leukemia markers|Leukemia markers
C1977241|T201|COMP|49494-8|LNC|Leukemia markers|Leukemia markers
C1977244|T201|COMP|49496-3|LNC|BCR-ABL1 e1a1 fusion protein|BCR-ABL1 e1a1 fusion protein
C1977245|T201|COMP|49497-1|LNC|Platelets|Platelets
C1977246|T201|COMP|49498-9|LNC|Leukocytes|Leukocytes
C1977247|T201|COMP|49499-7|LNC|Blood.dried/Total|Blood.dried/Total
C1977248|T201|COMP|49500-2|LNC|Calcium oxalate dihydrate/Total|Calcium oxalate dihydrate/Total
C1977249|T201|COMP|49501-0|LNC|Calcium oxalate monohydrate/Total|Calcium oxalate monohydrate/Total
C1977250|T201|COMP|49502-8|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C1977251|T201|COMP|49503-6|LNC|Neutrophil cytoplasmic Ab.perinuclear.atypical|Neutrophil cytoplasmic Ab.perinuclear.atypical
C1977253|T201|COMP|49504-4|LNC|CMT demyelinating gene targeted mutation analysis|CMT demyelinating gene targeted mutation analysis
C1977255|T201|COMP|49505-1|LNC|Erythrocyte clumps|Erythrocyte clumps
C1977256|T201|COMP|49506-9|LNC|MYOC gene targeted mutation analysis|MYOC gene targeted mutation analysis
C1977265|T201|COMP|49514-3|LNC|Acetaldehyde|Acetaldehyde
C1977266|T201|COMP|49515-0|LNC|Bisacodyl|Bisacodyl
C1977267|T201|COMP|49516-8|LNC|Topiramate^peak|Topiramate^peak
C1977268|T201|COMP|49517-6|LNC|Topiramate^trough|Topiramate^trough
C1977269|T201|COMP|49518-4|LNC|Influenza virus Ab|Influenza virus Ab
C1977270|T201|COMP|49519-2|LNC|Influenza virus A H16 Ab|Influenza virus A H16 Ab
C1977272|T201|COMP|49520-0|LNC|Influenza virus A H1 RNA|Influenza virus A H1 RNA
C1977274|T201|COMP|49521-8|LNC|Influenza virus A H1 RNA|Influenza virus A H1 RNA
C1977275|T201|COMP|49522-6|LNC|Influenza virus A H3 Ag|Influenza virus A H3 Ag
C1977277|T201|COMP|49523-4|LNC|Influenza virus A H3 RNA|Influenza virus A H3 RNA
C1977279|T201|COMP|49524-2|LNC|Influenza virus A H3 RNA|Influenza virus A H3 RNA
C1977280|T201|COMP|49525-9|LNC|Influenza virus A H5 Ab|Influenza virus A H5 Ab
C1977281|T201|COMP|49526-7|LNC|Influenza virus A H5 RNA|Influenza virus A H5 RNA
C1977282|T201|COMP|49527-5|LNC|Influenza virus A H7 RNA|Influenza virus A H7 RNA
C1977283|T201|COMP|49528-3|LNC|Influenza virus A H9 RNA|Influenza virus A H9 RNA
C1977285|T201|COMP|49529-1|LNC|Influenza virus A Ag|Influenza virus A Ag
C1977286|T201|COMP|49530-9|LNC|Influenza virus A neuraminidase cDNA|Influenza virus A neuraminidase cDNA
C1977287|T201|COMP|49531-7|LNC|Influenza virus A RNA|Influenza virus A RNA
C1977288|T201|COMP|49532-5|LNC|Influenza virus A hemagglutinin type RNA|Influenza virus A hemagglutinin type RNA
C1977289|T201|COMP|49533-3|LNC|Influenza virus B Ab|Influenza virus B Ab
C1977290|T201|COMP|49534-1|LNC|Influenza virus B Ag|Influenza virus B Ag
C1977291|T201|COMP|49535-8|LNC|Influenza virus B RNA|Influenza virus B RNA
C1977292|T201|COMP|49536-6|LNC|Influenza virus B RNA|Influenza virus B RNA
C1977294|T201|COMP|49537-4|LNC|Influenza virus A & B RNA|Influenza virus A & B RNA
C1977295|T201|COMP|49538-2|LNC|Influenza virus identified|Influenza virus identified
C1977296|T201|COMP|49539-0|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C1977297|T201|COMP|49540-8|LNC|Acid citrate dextrose|Acid citrate dextrose
C1977298|T201|COMP|49541-6|LNC|Fasting status|Fasting status
C1977299|T201|COMP|49542-4|LNC|Date and time of pheresis procedure|Date and time of pheresis procedure
C1977301|T201|COMP|49543-2|LNC|Calcidiol+Calciferol|Calcidiol+Calciferol
C1977302|T201|COMP|49544-0|LNC|Newborn screening recommended follow-up|Newborn screening recommended follow-up
C1977304|T201|COMP|49545-7|LNC|JC virus DNA|JC virus DNA
C1977305|T201|COMP|49546-5|LNC|Specimen age|Specimen age
C1977307|T201|COMP|49547-3|LNC|JC virus DNA|JC virus DNA
C1977308|T201|COMP|49548-1|LNC|Date reference lab test sent|Date reference lab test sent
C1977310|T201|COMP|49549-9|LNC|Reference lab test method|Reference lab test method
C1977312|T201|COMP|49550-7|LNC|Leukocytes.CD59 deficient/100 cells|Leukocytes.CD59 deficient/100 cells
C1977314|T201|COMP|49551-5|LNC|Creatine kinase.MB|Creatine kinase.MB
C1977315|T201|COMP|49552-3|LNC|Epinephrine+Norepinephrine|Epinephrine+Norepinephrine
C1977316|T201|COMP|49562-2|LNC|Holoprosencephaly gene targeted mutation analysis|Holoprosencephaly gene targeted mutation analysis
C1977318|T201|COMP|49563-0|LNC|Troponin I.cardiac|Troponin I.cardiac
C1977319|T201|COMP|49564-8|LNC|Epstein Barr virus band pattern|Epstein Barr virus band pattern
C1977330|T201|COMP|49572-1|LNC|Second trimester triple maternal screen|Second trimester triple maternal screen
C1977331|T201|COMP|49573-9|LNC|HIV genotype|HIV genotype
C1977334|T201|COMP|49575-4|LNC|Sphingomyelin/Surfactant.total|Sphingomyelin/Surfactant.total
C1977336|T201|COMP|49576-2|LNC|Phosphatidylethanolamine/Surfactants.total|Phosphatidylethanolamine/Surfactants.total
C1977338|T201|COMP|49585-3|LNC|Alpha-1-Fetoprotein multiple of the median cutoff|Alpha-1-Fetoprotein multiple of the median cutoff
C1977342|T201|COMP|49587-9|LNC|Protein.abnormal band|Protein.abnormal band
C1977345|T201|COMP|49589-5|LNC|Bacterial susceptibility panel|Bacterial susceptibility panel
C1977346|T201|COMP|49590-3|LNC|Calcidiol & Calciferol panel|Calcidiol & Calciferol panel
C1977348|T201|COMP|49591-1|LNC|Calcidiol & Calciferol|Calcidiol & Calciferol
C1977350|T201|COMP|49592-9|LNC|Satratoxin Ab.IgM|Satratoxin Ab.IgM
C1977352|T201|COMP|49593-7|LNC|Trichothecene Ab.IgA|Trichothecene Ab.IgA
C1977354|T201|COMP|49594-5|LNC|Trichothecene Ab.IgG|Trichothecene Ab.IgG
C1977356|T201|COMP|49595-2|LNC|Trichothecene Ab.IgM|Trichothecene Ab.IgM
C1977358|T201|COMP|49596-0|LNC|Uroporphyrinogen decarboxylase|Uroporphyrinogen decarboxylase
C1977359|T201|COMP|49597-8|LNC|Trichothecene Ab.IgE|Trichothecene Ab.IgE
C1977361|T201|COMP|49598-6|LNC|Natalizumab Ab|Natalizumab Ab
C1977363|T201|COMP|49599-4|LNC|Granulocytes.CD55|Granulocytes.CD55
C1977365|T201|COMP|49600-0|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977366|T201|COMP|49601-8|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977367|T201|COMP|49602-6|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977368|T201|COMP|49603-4|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977369|T201|COMP|49604-2|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977370|T201|COMP|49605-9|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977371|T201|COMP|49606-7|LNC|Hepatitis B virus DNA|Hepatitis B virus DNA
C1977372|T201|COMP|49607-5|LNC|Hepatitis C virus genotype|Hepatitis C virus genotype
C1977373|T201|COMP|49608-3|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977374|T201|COMP|49609-1|LNC|Vibrio sp DNA|Vibrio sp DNA
C1977376|T201|COMP|49610-9|LNC|Streptococcus pyogenes DNA|Streptococcus pyogenes DNA
C1977378|T201|COMP|49611-7|LNC|Streptococcus pneumoniae DNA|Streptococcus pneumoniae DNA
C1977380|T201|COMP|49612-5|LNC|Salmonella sp DNA|Salmonella sp DNA
C1977382|T201|COMP|49613-3|LNC|Enterococcus sp DNA|Enterococcus sp DNA
C1977383|T201|COMP|49614-1|LNC|Campylobacter sp DNA|Campylobacter sp DNA
C1977385|T201|COMP|49615-8|LNC|Borrelia sp DNA|Borrelia sp DNA
C1977387|T201|COMP|49616-6|LNC|Legionella sp DNA|Legionella sp DNA
C1977388|T201|COMP|49617-4|LNC|Bacterial carbapenem resistance blaKPC gene|Bacterial carbapenem resistance blaKPC gene
C1977390|T201|COMP|49618-2|LNC|Atazanavir+Ritonavir|Atazanavir+Ritonavir
C1977392|T201|COMP|49619-0|LNC|Indinavir+Ritonavir|Indinavir+Ritonavir
C1977394|T201|COMP|49620-8|LNC|lamiVUDine or Emtricitabine|lamiVUDine or Emtricitabine
C1977396|T201|COMP|49621-6|LNC|Saquinavir+Ritonavir|Saquinavir+Ritonavir
C1977398|T201|COMP|49622-4|LNC|Tipranavir+Ritonavir|Tipranavir+Ritonavir
C1977400|T201|COMP|49623-2|LNC|Amprenavir or Fosamprenavir|Amprenavir or Fosamprenavir
C1977402|T201|COMP|49624-0|LNC|Cholesterol.in VLDL 1+2|Cholesterol.in VLDL 1+2
C1977404|T201|COMP|49625-7|LNC|Granulocytes.CD59|Granulocytes.CD59
C1977406|T201|COMP|49646-3|LNC|SCA2 gene allele 2.CAG repeats|SCA2 gene allele 2.CAG repeats
C1977407|T201|COMP|49647-1|LNC|MJD gene allele 1.CAG repeats|MJD gene allele 1.CAG repeats
C1977408|T201|COMP|49648-9|LNC|MJD gene allele 2.CAG repeats|MJD gene allele 2.CAG repeats
C1977409|T201|COMP|49649-7|LNC|CACNA1A gene allele 1.CAG repeats|CACNA1A gene allele 1.CAG repeats
C1977411|T201|COMP|49650-5|LNC|CACNA1A gene allele 2.CAG repeats|CACNA1A gene allele 2.CAG repeats
C1977413|T201|COMP|49651-3|LNC|SCA7 gene allele 1.CAG repeats|SCA7 gene allele 1.CAG repeats
C1977415|T201|COMP|49652-1|LNC|SCA7 gene allele 2.CAG repeats|SCA7 gene allele 2.CAG repeats
C1977417|T201|COMP|49653-9|LNC|TPMT gene.c.719A>G|TPMT gene.c.719A>G
C1977419|T201|COMP|49654-7|LNC|TPMT gene.c.238G>C|TPMT gene.c.238G>C
C1977421|T201|COMP|49655-4|LNC|TPMT gene.c.460G>A|TPMT gene.c.460G>A
C1977423|T201|COMP|49656-2|LNC|HIV protease gene mutations|HIV protease gene mutations
C1977429|T201|COMP|49659-6|LNC|HIV reverse transcriptase susceptibility panel|HIV reverse transcriptase susceptibility panel
C1977431|T201|COMP|49660-4|LNC|HIV susceptibility panel|HIV susceptibility panel
C1977433|T201|COMP|49661-2|LNC|HIV protease gene mutations|HIV protease gene mutations
C1977436|T201|COMP|49664-6|LNC|HIV reverse transcriptase susceptibility panel|HIV reverse transcriptase susceptibility panel
C1977437|T201|COMP|49665-3|LNC|HIV susceptibility panel|HIV susceptibility panel
C1977439|T201|COMP|49666-1|LNC|Darunavir|Darunavir
C1977440|T201|COMP|49667-9|LNC|Tipranavir|Tipranavir
C1977441|T201|COMP|49668-7|LNC|Atazanavir|Atazanavir
C1977442|T201|COMP|49669-5|LNC|Emtricitabine|Emtricitabine
C1977443|T201|COMP|49670-3|LNC|Uranium.depleted panel|Uranium.depleted panel
C1977445|T201|COMP|49671-1|LNC|Neisseria meningitidis DNA|Neisseria meningitidis DNA
C1977447|T201|COMP|49672-9|LNC|Streptococcus pneumoniae DNA|Streptococcus pneumoniae DNA
C1977455|T201|COMP|49678-6|LNC|CPT2 gene targeted mutation analysis|CPT2 gene targeted mutation analysis
C1977457|T201|COMP|49679-4|LNC|Cells.CD36/100 cells|Cells.CD36/100 cells
C1977458|T201|COMP|49680-2|LNC|Cells.CD36/100 cells|Cells.CD36/100 cells
C1977459|T201|COMP|49681-0|LNC|Cells.CD36/100 cells|Cells.CD36/100 cells
C1977461|T201|COMP|49683-6|LNC|HER2 gene copy number/Chromosome 17 copy number|HER2 gene copy number/Chromosome 17 copy number
C1977463|T201|COMP|49684-4|LNC|CPT2 gene.p.Arg503Cys|CPT2 gene.p.Arg503Cys
C1977465|T201|COMP|49685-1|LNC|CPT2 gene.p.R549DC|CPT2 gene.p.R549DC
C1977467|T201|COMP|49686-9|LNC|CPT2 gene.p.Arg631Cys|CPT2 gene.p.Arg631Cys
C1977469|T201|COMP|49687-7|LNC|Trichoderma viride Ab.IgG|Trichoderma viride Ab.IgG
C1977470|T201|COMP|49701-6|LNC|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1977471|T201|COMP|49702-4|LNC|Nateglinide|Nateglinide
C1977472|T201|COMP|49704-0|LNC|SH3TC2 gene targeted mutation analysis|SH3TC2 gene targeted mutation analysis
C1977474|T201|COMP|49705-7|LNC|LMNA gene targeted mutation analysis|LMNA gene targeted mutation analysis
C1977475|T201|COMP|49706-5|LNC|ARSA gene targeted mutation analysis|ARSA gene targeted mutation analysis
C1977477|T201|COMP|49707-3|LNC|KCNQ2 gene targeted mutation analysis|KCNQ2 gene targeted mutation analysis
C1977479|T201|COMP|49708-1|LNC|TTR gene targeted mutation analysis|TTR gene targeted mutation analysis
C1977480|T201|COMP|49718-0|LNC|HIV 1 p24 Ag|HIV 1 p24 Ag
C1977481|T201|COMP|49719-8|LNC|Poa pratensis Ab.IgG|Poa pratensis Ab.IgG
C1977482|T201|COMP|49720-6|LNC|Festuca elatior Ab.IgG|Festuca elatior Ab.IgG
C1977483|T201|COMP|49721-4|LNC|Haemophilus influenzae type|Haemophilus influenzae type
C1977485|T201|COMP|49722-2|LNC|Neisseria meningitidis type|Neisseria meningitidis type
C1977487|T201|COMP|49723-0|LNC|Camellia sinensis Ab.IgG|Camellia sinensis Ab.IgG
C1977488|T201|COMP|49724-8|LNC|Aldolase|Aldolase
C1977489|T201|COMP|49725-5|LNC|Melatonin|Melatonin
C1977490|T201|COMP|49742-0|LNC|Plasmodium vivax Ab.IgG|Plasmodium vivax Ab.IgG
C1977492|T201|COMP|49743-8|LNC|Plasmodium falciparum Ab.IgG|Plasmodium falciparum Ab.IgG
C1977494|T201|COMP|49744-6|LNC|Plasmodium ovale Ab.IgG|Plasmodium ovale Ab.IgG
C1977496|T201|COMP|49745-3|LNC|Dolichovespula maculata Ab.IgG|Dolichovespula maculata Ab.IgG
C1977497|T201|COMP|49746-1|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C1977498|T201|COMP|49747-9|LNC|Cocaine+Benzoylecgonine|Cocaine+Benzoylecgonine
C1977499|T201|COMP|49748-7|LNC|Lipoprotein.alpha|Lipoprotein.alpha
C1977500|T201|COMP|49749-5|LNC|6-Monoacetylmorphine.free|6-Monoacetylmorphine.free
C1977501|T201|COMP|49750-3|LNC|Dihydrocodeine.free+Hydrocodol.free|Dihydrocodeine.free+Hydrocodol.free
C1977502|T201|COMP|49751-1|LNC|Norbuprenorphine|Norbuprenorphine
C1977503|T201|COMP|49752-9|LNC|Buprenorphine|Buprenorphine
C1977504|T201|COMP|49753-7|LNC|Norbuprenorphine|Norbuprenorphine
C1977505|T201|COMP|49754-5|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C1977506|T201|COMP|49755-2|LNC|Crystals|Crystals
C1977507|T201|COMP|49756-0|LNC|Norethindrone|Norethindrone
C1977508|T201|COMP|49757-8|LNC|Minocycline|Minocycline
C1977509|T201|COMP|49758-6|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C1977510|T201|COMP|49759-4|LNC|Adenosine deaminase|Adenosine deaminase
C1977511|T201|COMP|49760-2|LNC|Adenosine deaminase|Adenosine deaminase
C1977512|T201|COMP|49761-0|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C1977513|T201|COMP|49762-8|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C1977514|T201|COMP|49763-6|LNC|Bilirubin|Bilirubin
C1977515|T201|COMP|49764-4|LNC|Calcium|Calcium
C1977516|T201|COMP|49765-1|LNC|Calcium|Calcium
C1977517|T201|COMP|49766-9|LNC|Chymotrypsin|Chymotrypsin
C1977518|T201|COMP|49775-0|LNC|Hepatitis D virus Ab.IgG|Hepatitis D virus Ab.IgG
C1977519|T201|COMP|49776-8|LNC|Hepatitis E virus Ab|Hepatitis E virus Ab
C1977520|T201|COMP|49777-6|LNC|Hepatitis G virus Ab|Hepatitis G virus Ab
C1977521|T201|COMP|49778-4|LNC|Immune complex|Immune complex
C1977522|T201|COMP|49779-2|LNC|Ketones|Ketones
C1977523|T201|COMP|49780-0|LNC|Leishmania sp DNA|Leishmania sp DNA
C1977524|T201|COMP|49781-8|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C1977525|T201|COMP|49868-3|LNC|Ibuprofen Ab.IgE|Ibuprofen Ab.IgE
C1977527|T201|COMP|49869-1|LNC|Camel dander Ab.IgE|Camel dander Ab.IgE
C1977529|T201|COMP|49870-9|LNC|Coagulation factor VII Ag actual/Normal|Coagulation factor VII Ag actual/Normal
C1977531|T201|COMP|49871-7|LNC|Codeine Ab.IgE|Codeine Ab.IgE
C1977533|T201|COMP|49872-5|LNC|FH gene targeted mutation analysis|FH gene targeted mutation analysis
C1977535|T201|COMP|49873-3|LNC|POU3F4 gene targeted mutation analysis|POU3F4 gene targeted mutation analysis
C1977537|T201|COMP|49874-1|LNC|ABCB4 gene targeted mutation analysis|ABCB4 gene targeted mutation analysis
C1977539|T201|COMP|49875-8|LNC|Juniperus californica Ab.IgE|Juniperus californica Ab.IgE
C1977541|T201|COMP|50002-5|LNC|Hydrogen/Expired gas^1.5H post XXX challenge|Hydrogen/Expired gas^1.5H post XXX challenge
C1977542|T201|COMP|50003-3|LNC|Hydrogen/Expired gas^2H post XXX challenge|Hydrogen/Expired gas^2H post XXX challenge
C1977543|T201|COMP|50004-1|LNC|Hydrogen/Expired gas^3H post XXX challenge|Hydrogen/Expired gas^3H post XXX challenge
C1977544|T201|COMP|50005-8|LNC|Methaqualone|Methaqualone
C1977545|T201|COMP|50006-6|LNC|Human antimouse Ab|Human antimouse Ab
C1977546|T201|COMP|50007-4|LNC|Cytology report|Cytology report
C1977547|T201|COMP|50008-2|LNC|Mixing studies|Mixing studies
C1977549|T201|COMP|50009-0|LNC|Fetal lung maturity panel|Fetal lung maturity panel
C1977551|T201|COMP|50314-4|LNC|Cytokeratin 19 Ag|Cytokeratin 19 Ag
C1977553|T201|COMP|50315-1|LNC|Cytokeratin 5 Ag|Cytokeratin 5 Ag
C1977555|T201|COMP|50316-9|LNC|Galectin 3 Ag|Galectin 3 Ag
C1977557|T201|COMP|50317-7|LNC|CD235a Ag|CD235a Ag
C1977559|T201|COMP|50318-5|LNC|Granzyme B Ag|Granzyme B Ag
C1977561|T201|COMP|50319-3|LNC|HBME-1 Ag|HBME-1 Ag
C1977562|T201|COMP|50320-1|LNC|Helicobacter pylori Ag|Helicobacter pylori Ag
C1977563|T201|COMP|50321-9|LNC|Hepatocyte Ag|Hepatocyte Ag
C1977565|T201|COMP|50322-7|LNC|MLH-1 Ag|MLH-1 Ag
C1977567|T201|COMP|50734-3|LNC|Serotonin release.heparin.porcine interpretation|Serotonin release.heparin.porcine interpretation
C1977571|T201|COMP|50736-8|LNC|Serotonin release.heparin.unfractionated panel|Serotonin release.heparin.unfractionated panel
C1977573|T201|COMP|50737-6|LNC|Serotonin release.heparin.porcine panel|Serotonin release.heparin.porcine panel
C1977581|T201|COMP|50903-4|LNC|Selenium|Selenium
C1977582|T201|COMP|50904-2|LNC|Selenium|Selenium
C1977583|T201|COMP|50905-9|LNC|Silicon|Silicon
C1977584|T201|COMP|50906-7|LNC|Silicon|Silicon
C1977585|T201|COMP|50907-5|LNC|Silicon|Silicon
C1977586|T201|COMP|50908-3|LNC|Silver|Silver
C1977587|T201|COMP|50909-1|LNC|Silver|Silver
C1977588|T201|COMP|50910-9|LNC|Silver|Silver
C1977589|T201|COMP|50911-7|LNC|Sodium|Sodium
C1977599|T201|COMP|50992-7|LNC|IgM|IgM
C1977600|T201|COMP|50993-5|LNC|Laxatives|Laxatives
C1977601|T201|COMP|50994-3|LNC|CMT demyelinating gene targeted mutation analysis|CMT demyelinating gene targeted mutation analysis
C1977602|T201|COMP|49782-6|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C1977603|T201|COMP|49783-4|LNC|Onchocerca sp Ab.IgG4|Onchocerca sp Ab.IgG4
C1977605|T201|COMP|49784-2|LNC|Onchocerca sp Ab.IgG|Onchocerca sp Ab.IgG
C1977606|T201|COMP|49785-9|LNC|Onchocerca sp Ab.IgG2|Onchocerca sp Ab.IgG2
C1977608|T201|COMP|49786-7|LNC|Onchocerca sp Ab.IgG3|Onchocerca sp Ab.IgG3
C1977610|T201|COMP|49787-5|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C1977611|T201|COMP|49788-3|LNC|Potassium|Potassium
C1977612|T201|COMP|49789-1|LNC|Potassium|Potassium
C1977613|T201|COMP|49798-2|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C1977614|T201|COMP|49799-0|LNC|Treponema pallidum DNA|Treponema pallidum DNA
C1977615|T201|COMP|49800-6|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1977616|T201|COMP|49801-4|LNC|Trypanosoma cruzi DNA|Trypanosoma cruzi DNA
C1977618|T201|COMP|49802-2|LNC|Urea|Urea
C1977619|T201|COMP|49803-0|LNC|Streptococcus pneumoniae 1 Ab^1st specimen|Streptococcus pneumoniae 1 Ab^1st specimen
C1977620|T201|COMP|49804-8|LNC|Streptococcus pneumoniae 19 Ab^1st specimen|Streptococcus pneumoniae 19 Ab^1st specimen
C1977621|T201|COMP|49805-5|LNC|Streptococcus pneumoniae 23 Ab^1st specimen|Streptococcus pneumoniae 23 Ab^1st specimen
C1977622|T201|COMP|49806-3|LNC|Streptococcus pneumoniae 1 Ab^2nd specimen|Streptococcus pneumoniae 1 Ab^2nd specimen
C1977623|T201|COMP|49807-1|LNC|Streptococcus pneumoniae 19 Ab^2nd specimen|Streptococcus pneumoniae 19 Ab^2nd specimen
C1977624|T201|COMP|49808-9|LNC|Streptococcus pneumoniae 23 Ab^2nd specimen|Streptococcus pneumoniae 23 Ab^2nd specimen
C1977625|T201|COMP|49809-7|LNC|2-Ethyl-3-Hydroxypropionate/Creatinine|2-Ethyl-3-Hydroxypropionate/Creatinine
C1977626|T201|COMP|49810-5|LNC|2-Hydroxy-3-Methylvalerate/Creatinine|2-Hydroxy-3-Methylvalerate/Creatinine
C1977627|T201|COMP|49811-3|LNC|2-Hydroxyadipate/Creatinine|2-Hydroxyadipate/Creatinine
C1977628|T201|COMP|49812-1|LNC|2-Hydroxyglutarate/Creatinine|2-Hydroxyglutarate/Creatinine
C1977629|T201|COMP|49813-9|LNC|2-Hydroxyisocaproate/Creatinine|2-Hydroxyisocaproate/Creatinine
C1977630|T201|COMP|49814-7|LNC|2-Hydroxyisovalerate/Creatinine|2-Hydroxyisovalerate/Creatinine
C1977631|T201|COMP|49815-4|LNC|2-Methyl-3-Hydroxybutyrate/Creatinine|2-Methyl-3-Hydroxybutyrate/Creatinine
C1977632|T201|COMP|49816-2|LNC|2-Oxo,3-Methylvalerate/Creatinine|2-Oxo,3-Methylvalerate/Creatinine
C1977633|T201|COMP|49817-0|LNC|2-Oxoisocaproate/Creatinine|2-Oxoisocaproate/Creatinine
C1977634|T201|COMP|49818-8|LNC|2-Oxoisovalerate/Creatinine|2-Oxoisovalerate/Creatinine
C1977635|T201|COMP|49819-6|LNC|3-Hydroxy,3-Methylglutarate/Creatinine|3-Hydroxy,3-Methylglutarate/Creatinine
C1977636|T201|COMP|49820-4|LNC|3-Hydroxyadipate/Creatinine|3-Hydroxyadipate/Creatinine
C1977637|T201|COMP|49821-2|LNC|3-Hydroxyglutarate/Creatinine|3-Hydroxyglutarate/Creatinine
C1977638|T201|COMP|49822-0|LNC|3-Hydroxyisobutyrate/Creatinine|3-Hydroxyisobutyrate/Creatinine
C1977639|T201|COMP|49823-8|LNC|3-Hydroxyisovalerate/Creatinine|3-Hydroxyisovalerate/Creatinine
C1977640|T201|COMP|49824-6|LNC|3-Hydroxypropionate/Creatinine|3-Hydroxypropionate/Creatinine
C1977641|T201|COMP|49825-3|LNC|16-Alpha hydroxyestrone|16-Alpha hydroxyestrone
C1977642|T201|COMP|49826-1|LNC|2-Hydroxyestrone|2-Hydroxyestrone
C1977643|T201|COMP|49827-9|LNC|2-Hydroxyestrone/16-Alpha hydroxyestrone|2-Hydroxyestrone/16-Alpha hydroxyestrone
C1977645|T201|COMP|49828-7|LNC|2-Hydroxyestrone & 16-Alpha hydroxyestrone panel|2-Hydroxyestrone & 16-Alpha hydroxyestrone panel
C1977647|T201|COMP|49829-5|LNC|Norcodeine|Norcodeine
C1977648|T201|COMP|49830-3|LNC|Norcodeine|Norcodeine
C1977649|T201|COMP|49831-1|LNC|Normorphine|Normorphine
C1977650|T201|COMP|49832-9|LNC|Specimen drawn^1st specimen|Specimen drawn^1st specimen
C1977651|T201|COMP|49833-7|LNC|Specimen drawn^2nd specimen|Specimen drawn^2nd specimen
C1977652|T201|COMP|49834-5|LNC|Leucine|Leucine
C1977653|T201|COMP|49835-2|LNC|Cells.CD19+IgD+/100 cells|Cells.CD19+IgD+/100 cells
C1977655|T201|COMP|49851-9|LNC|Cholinesterase|Cholinesterase
C1977656|T201|COMP|49852-7|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C1977657|T201|COMP|49860-0|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C1977658|T201|COMP|49861-8|LNC|Toxocara canis Ab|Toxocara canis Ab
C1977659|T201|COMP|49862-6|LNC|G6PC gene targeted mutation analysis|G6PC gene targeted mutation analysis
C1977661|T201|COMP|49863-4|LNC|Aspergillus sp DNA|Aspergillus sp DNA
C1977663|T201|COMP|49864-2|LNC|Novocaine Ab.IgE|Novocaine Ab.IgE
C1977665|T201|COMP|49865-9|LNC|Coagulation factor VIII activity actual/Normal|Coagulation factor VIII activity actual/Normal
C1977666|T201|COMP|49866-7|LNC|Neuropeptide Y|Neuropeptide Y
C1977667|T201|COMP|49867-5|LNC|Endothelin I|Endothelin I
C1977669|T201|COMP|49986-3|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C1977670|T201|COMP|49987-1|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C1977671|T201|COMP|49988-9|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C1977672|T201|COMP|49989-7|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C1977673|T201|COMP|49990-5|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C1977674|T201|COMP|49991-3|LNC|Borrelia burgdorferi 18_20kD Ab.IgG|Borrelia burgdorferi 18_20kD Ab.IgG
C1977676|T201|COMP|49992-1|LNC|Borrelia burgdorferi 18_20kD Ab.IgG|Borrelia burgdorferi 18_20kD Ab.IgG
C1977677|T201|COMP|49993-9|LNC|Borrelia burgdorferi 18_20kD Ab.IgM|Borrelia burgdorferi 18_20kD Ab.IgM
C1977679|T201|COMP|49994-7|LNC|Borrelia burgdorferi 18_20kD Ab.IgM|Borrelia burgdorferi 18_20kD Ab.IgM
C1977680|T201|COMP|50123-9|LNC|3-Hydroxypalmitoylcarnitine (C16-OH)|3-Hydroxypalmitoylcarnitine (C16-OH)
C1977681|T201|COMP|50124-7|LNC|3-Hydroxypalmitoylcarnitine (C16-OH)|3-Hydroxypalmitoylcarnitine (C16-OH)
C1977682|T201|COMP|50125-4|LNC|3-Hydroxypalmitoylcarnitine (C16-OH)|3-Hydroxypalmitoylcarnitine (C16-OH)
C1977683|T201|COMP|50126-2|LNC|3-Hydroxypalmitoylcarnitine (C16-OH)|3-Hydroxypalmitoylcarnitine (C16-OH)
C1977684|T201|COMP|50127-0|LNC|3-Hydroxypalmitoylcarnitine (C16-OH)/Creatinine|3-Hydroxypalmitoylcarnitine (C16-OH)/Creatinine
C1977686|T201|COMP|50128-8|LNC|3-Hydroxypropionate|3-Hydroxypropionate
C1977687|T201|COMP|50129-6|LNC|3-Hydroxypropionate|3-Hydroxypropionate
C1977688|T201|COMP|50130-4|LNC|3-Hydroxystearoylcarnitine (C18-OH)|3-Hydroxystearoylcarnitine (C18-OH)
C1977689|T201|COMP|50131-2|LNC|3-Hydroxystearoylcarnitine (C18-OH)|3-Hydroxystearoylcarnitine (C18-OH)
C1977690|T201|COMP|50202-1|LNC|Iron^5th specimen|Iron^5th specimen
C1977691|T201|COMP|50203-9|LNC|Iron^6th specimen|Iron^6th specimen
C1977692|T201|COMP|50204-7|LNC|Iron^7th specimen|Iron^7th specimen
C1977693|T201|COMP|50205-4|LNC|Iron^8th specimen|Iron^8th specimen
C1977694|T201|COMP|50206-2|LNC|Glucose^1st specimen|Glucose^1st specimen
C1977695|T201|COMP|50207-0|LNC|Glucose^7th specimen|Glucose^7th specimen
C1977696|T201|COMP|50208-8|LNC|Glucose^10th specimen|Glucose^10th specimen
C1977697|T201|COMP|50209-6|LNC|Albumin^supine|Albumin^supine
C1977698|T201|COMP|50775-6|LNC|Cancer Ag 125|Cancer Ag 125
C1977699|T201|COMP|50776-4|LNC|Cancer Ag 15-3|Cancer Ag 15-3
C1977700|T201|COMP|50777-2|LNC|Cancer Ag 15-3|Cancer Ag 15-3
C1977701|T201|COMP|50778-0|LNC|Cancer Ag 15-3|Cancer Ag 15-3
C1977702|T201|COMP|50779-8|LNC|Cancer Ag 19-9|Cancer Ag 19-9
C1977703|T201|COMP|50780-6|LNC|Cancer Ag 19-9|Cancer Ag 19-9
C1977704|T201|COMP|50781-4|LNC|Cancer Ag 19-9|Cancer Ag 19-9
C1977705|T201|COMP|50782-2|LNC|Cancer Ag 27-29|Cancer Ag 27-29
C1977706|T201|COMP|51265-7|LNC|Cells.CD19/100 cells|Cells.CD19/100 cells
C1977707|T201|COMP|51266-5|LNC|Cells.CD23/100 cells|Cells.CD23/100 cells
C1977708|T201|COMP|51267-3|LNC|Cells.CD23/100 cells|Cells.CD23/100 cells
C1977709|T201|COMP|51268-1|LNC|Cells.CD23/100 cells|Cells.CD23/100 cells
C1977710|T201|COMP|51269-9|LNC|Cells.CD23/100 cells|Cells.CD23/100 cells
C1977711|T201|COMP|51270-7|LNC|Cells.CD25/100 cells|Cells.CD25/100 cells
C1977712|T201|COMP|51271-5|LNC|Cells.CD25/100 cells|Cells.CD25/100 cells
C1977713|T201|COMP|51272-3|LNC|Cells.CD25+CD19+/100 cells|Cells.CD25+CD19+/100 cells
C1977714|T201|COMP|51273-1|LNC|Cells.CD3/100 cells|Cells.CD3/100 cells
C1977717|T201|COMP|51339-0|LNC|Cells.CD45/100 cells|Cells.CD45/100 cells
C1977718|T201|COMP|51340-8|LNC|Cells.CD45/100 cells|Cells.CD45/100 cells
C1977719|T201|COMP|51341-6|LNC|Cells.CD5+CD19+/100 cells|Cells.CD5+CD19+/100 cells
C1977720|T201|COMP|51342-4|LNC|Cells.CD5+CD19+/100 cells|Cells.CD5+CD19+/100 cells
C1977721|T201|COMP|51343-2|LNC|Cells.CD55/100 cells|Cells.CD55/100 cells
C1977722|T201|COMP|51344-0|LNC|Cells.CD55/100 cells|Cells.CD55/100 cells
C1977723|T201|COMP|51345-7|LNC|Cells.CD56+CD57+/100 cells|Cells.CD56+CD57+/100 cells
C1977725|T201|COMP|51346-5|LNC|Cells.CD56+CD57+/100 cells|Cells.CD56+CD57+/100 cells
C1977728|T201|COMP|51413-3|LNC|Butyrylcarnitine+Isobutyrylcarnitine (C4)|Butyrylcarnitine+Isobutyrylcarnitine (C4)
C1977732|T201|COMP|51415-8|LNC|Methylmalonylcarnitine+Succinylcarnitine (C4-DC)|Methylmalonylcarnitine+Succinylcarnitine (C4-DC)
C1977734|T201|COMP|51416-6|LNC|Tiglylcarnitine (C5:1)|Tiglylcarnitine (C5:1)
C1977735|T201|COMP|51417-4|LNC|Coproporphyrin/Porphyrins.total|Coproporphyrin/Porphyrins.total
C1977737|T201|COMP|51418-2|LNC|Domperidone|Domperidone
C1977738|T201|COMP|51419-0|LNC|Sodium^^corrected for glucose|Sodium^^corrected for glucose
C1977739|T201|COMP|49876-6|LNC|Alpha hydroxytriazolam|Alpha hydroxytriazolam
C1977740|T201|COMP|49877-4|LNC|Hepatitis B virus codon 173|Hepatitis B virus codon 173
C1977742|T201|COMP|49878-2|LNC|Hepatitis B virus codon 180|Hepatitis B virus codon 180
C1977744|T201|COMP|49879-0|LNC|Hepatitis B virus codon 181|Hepatitis B virus codon 181
C1977746|T201|COMP|49880-8|LNC|Hepatitis B virus codon 204|Hepatitis B virus codon 204
C1977748|T201|COMP|49881-6|LNC|Hepatitis B virus codon 236|Hepatitis B virus codon 236
C1977750|T201|COMP|49882-4|LNC|Hepatitis B virus codon 80|Hepatitis B virus codon 80
C1977752|T201|COMP|49883-2|LNC|Hepatitis B virus resistance panel|Hepatitis B virus resistance panel
C1977761|T201|COMP|49890-7|LNC|HIV 1 RNA|HIV 1 RNA
C1977762|T201|COMP|49891-5|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C1977763|T201|COMP|49892-3|LNC|Somatotropin^1st specimen post XXX challenge|Somatotropin^1st specimen post XXX challenge
C1977764|T201|COMP|49893-1|LNC|Somatotropin^7th specimen post XXX challenge|Somatotropin^7th specimen post XXX challenge
C1977765|T201|COMP|49894-9|LNC|Somatotropin^9th specimen post XXX challenge|Somatotropin^9th specimen post XXX challenge
C1977766|T201|COMP|49895-6|LNC|Somatotropin^10th specimen post XXX challenge|Somatotropin^10th specimen post XXX challenge
C1977768|T201|COMP|49897-2|LNC|Insulin^pre XXX challenge|Insulin^pre XXX challenge
C1977769|T201|COMP|49898-0|LNC|Metabolic syndrome|Metabolic syndrome
C1977770|T201|COMP|49899-8|LNC|Setomelanomma rostrata Ab.IgE/IgE.total|Setomelanomma rostrata Ab.IgE/IgE.total
C1977771|T201|COMP|49900-4|LNC|Heptacarboxylporphyrin I|Heptacarboxylporphyrin I
C1977772|T201|COMP|49901-2|LNC|Heptacarboxylporphyrin III|Heptacarboxylporphyrin III
C1977773|T201|COMP|49902-0|LNC|Hexanoylglycine/Creatinine|Hexanoylglycine/Creatinine
C1977774|T201|COMP|49903-8|LNC|Hippurate/Creatinine|Hippurate/Creatinine
C1977775|T201|COMP|49904-6|LNC|Histoplasma capsulatum M Ab|Histoplasma capsulatum M Ab
C1977776|T201|COMP|49905-3|LNC|HIV 1 Ab|HIV 1 Ab
C1977777|T201|COMP|49906-1|LNC|Hydroxydecanedioate/Creatinine|Hydroxydecanedioate/Creatinine
C1977778|T201|COMP|49907-9|LNC|IgA Ag|IgA Ag
C1977780|T201|COMP|49909-5|LNC|Interleukin 10|Interleukin 10
C1977781|T201|COMP|49910-3|LNC|Isocitrate/Creatinine|Isocitrate/Creatinine
C1977782|T201|COMP|49911-1|LNC|Isovalerylglycine/Creatinine|Isovalerylglycine/Creatinine
C1977783|T201|COMP|49912-9|LNC|Japanese encephalitis virus Ab|Japanese encephalitis virus Ab
C1977784|T201|COMP|49913-7|LNC|Legionella pneumophila Ab.IgG|Legionella pneumophila Ab.IgG
C1977785|T201|COMP|49914-5|LNC|Legionella pneumophila 1+2+3+4+5+6 Ab.IgM|Legionella pneumophila 1+2+3+4+5+6 Ab.IgM
C1977787|T201|COMP|49915-2|LNC|Legionella sp Ab.IgG|Legionella sp Ab.IgG
C1977789|T201|COMP|49916-0|LNC|Liquidambar styraciflua Ab.IgE/IgE.total|Liquidambar styraciflua Ab.IgE/IgE.total
C1977791|T201|COMP|49918-6|LNC|Heptacarboxylporphyrin II|Heptacarboxylporphyrin II
C1977793|T201|COMP|49919-4|LNC|Interleukin 6|Interleukin 6
C1977794|T201|COMP|49920-2|LNC|Isopropyl ether|Isopropyl ether
C1977802|T201|COMP|49925-1|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C1977803|T201|COMP|49926-9|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C1977804|T201|COMP|49927-7|LNC|Amylase.fld/Amylase.serum|Amylase.fld/Amylase.serum
C1977807|T201|COMP|49928-5|LNC|Leukocytes|Leukocytes
C1977808|T201|COMP|49929-3|LNC|Protein.plr fld/Protein.serum|Protein.plr fld/Protein.serum
C1977813|T201|COMP|49931-9|LNC|3-Hydroxysebacate.unsaturated/Creatinine|3-Hydroxysebacate.unsaturated/Creatinine
C1977815|T201|COMP|49932-7|LNC|3-Hydroxysuberate.unsaturated/Creatinine|3-Hydroxysuberate.unsaturated/Creatinine
C1977817|T201|COMP|49933-5|LNC|Adipate.unsaturated/Creatinine|Adipate.unsaturated/Creatinine
C1977819|T201|COMP|49934-3|LNC|Adipolactone/Creatinine|Adipolactone/Creatinine
C1977824|T201|COMP|49937-6|LNC|Calcium/Oxalate|Calcium/Oxalate
C1977825|T201|COMP|49938-4|LNC|Citrate synthase|Citrate synthase
C1977826|T201|COMP|49954-1|LNC|Somatotropin^4 AM specimen|Somatotropin^4 AM specimen
C1977827|T201|COMP|49955-8|LNC|Somatotropin^4.30 AM specimen|Somatotropin^4.30 AM specimen
C1977828|T201|COMP|49956-6|LNC|Somatotropin^5 AM specimen|Somatotropin^5 AM specimen
C1977829|T201|COMP|49957-4|LNC|Somatotropin^5.30 AM specimen|Somatotropin^5.30 AM specimen
C1977830|T201|COMP|49958-2|LNC|Somatotropin^6 AM specimen|Somatotropin^6 AM specimen
C1977831|T201|COMP|49959-0|LNC|Specific gravity^^adjusted to pH 7.4|Specific gravity^^adjusted to pH 7.4
C1977832|T201|COMP|49960-8|LNC|Suberate.unsaturated/Creatinine|Suberate.unsaturated/Creatinine
C1977834|T201|COMP|49961-6|LNC|Urate renal clearance|Urate renal clearance
C1977835|T201|COMP|49962-4|LNC|Urate renal clearance/1.73 sq M|Urate renal clearance/1.73 sq M
C1977837|T201|COMP|49963-2|LNC|Fibrillarin Ab|Fibrillarin Ab
C1977839|T201|COMP|49964-0|LNC|Siderocytes|Siderocytes
C1977840|T201|COMP|49965-7|LNC|HIV 1 Ab/HIV 2 Ab|HIV 1 Ab/HIV 2 Ab
C1977842|T201|COMP|49966-5|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C1977843|T201|COMP|49967-3|LNC|Charcoal|Charcoal
C1977844|T201|COMP|49968-1|LNC|Cortisol^1H post 250 ug corticotropin IM|Cortisol^1H post 250 ug corticotropin IM
C1977845|T201|COMP|49969-9|LNC|Cortisol^30M post 250 ug corticotropin IM|Cortisol^30M post 250 ug corticotropin IM
C1977846|T201|COMP|49970-7|LNC|Collection time^4th specimen|Collection time^4th specimen
C1977847|T201|COMP|49971-5|LNC|Collection time^3rd specimen|Collection time^3rd specimen
C1977848|T201|COMP|49972-3|LNC|Collection time^2nd specimen|Collection time^2nd specimen
C1977849|T201|COMP|49973-1|LNC|Borrelia burgdorferi 31kD Ab.IgG|Borrelia burgdorferi 31kD Ab.IgG
C1977850|T201|COMP|49974-9|LNC|Borrelia burgdorferi 31kD Ab.IgM|Borrelia burgdorferi 31kD Ab.IgM
C1977851|T201|COMP|49975-6|LNC|Borrelia burgdorferi 34kD Ab.IgG|Borrelia burgdorferi 34kD Ab.IgG
C1977852|T201|COMP|49976-4|LNC|Borrelia burgdorferi 34kD Ab.IgM|Borrelia burgdorferi 34kD Ab.IgM
C1977853|T201|COMP|49977-2|LNC|Borrelia burgdorferi 35kD Ab.IgG|Borrelia burgdorferi 35kD Ab.IgG
C1977855|T201|COMP|49978-0|LNC|Borrelia burgdorferi 35kD Ab.IgG|Borrelia burgdorferi 35kD Ab.IgG
C1977856|T201|COMP|49979-8|LNC|Borrelia burgdorferi 35kD Ab.IgM|Borrelia burgdorferi 35kD Ab.IgM
C1977858|T201|COMP|49980-6|LNC|Borrelia burgdorferi 35kD Ab.IgM|Borrelia burgdorferi 35kD Ab.IgM
C1977859|T201|COMP|49981-4|LNC|Borrelia burgdorferi 37kD Ab.IgG|Borrelia burgdorferi 37kD Ab.IgG
C1977861|T201|COMP|49982-2|LNC|Borrelia burgdorferi 37kD Ab.IgG|Borrelia burgdorferi 37kD Ab.IgG
C1977862|T201|COMP|49983-0|LNC|Borrelia burgdorferi 37kD Ab.IgM|Borrelia burgdorferi 37kD Ab.IgM
C1977864|T201|COMP|49984-8|LNC|Borrelia burgdorferi 37kD Ab.IgM|Borrelia burgdorferi 37kD Ab.IgM
C1977865|T201|COMP|49985-5|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C1977866|T201|COMP|49995-4|LNC|Borrelia burgdorferi 83_93kD Ab.IgG|Borrelia burgdorferi 83_93kD Ab.IgG
C1977868|T201|COMP|49996-2|LNC|Borrelia burgdorferi 83_93kD Ab.IgG|Borrelia burgdorferi 83_93kD Ab.IgG
C1977869|T201|COMP|49997-0|LNC|Borrelia burgdorferi 83_93kD Ab.IgM|Borrelia burgdorferi 83_93kD Ab.IgM
C1977871|T201|COMP|49998-8|LNC|Borrelia burgdorferi 83_93kD Ab.IgM|Borrelia burgdorferi 83_93kD Ab.IgM
C1977872|T201|COMP|49999-6|LNC|Platelet aggregation.collagen induced|Platelet aggregation.collagen induced
C1977873|T201|COMP|50000-9|LNC|Hydrogen/Expired gas^30M post XXX challenge|Hydrogen/Expired gas^30M post XXX challenge
C1977874|T201|COMP|50001-7|LNC|Hydrogen/Expired gas^1H post XXX challenge|Hydrogen/Expired gas^1H post XXX challenge
C1977875|T201|COMP|50010-8|LNC|Transfusion end time|Transfusion end time
C1977877|T201|COMP|50011-6|LNC|Transfusion start time|Transfusion start time
C1977879|T201|COMP|50012-4|LNC|Indirect antiglobulin test.poly specific reagent|Indirect antiglobulin test.poly specific reagent
C1977880|T201|COMP|50013-2|LNC|Hydrogen/Expired gas^2.5H post XXX challenge|Hydrogen/Expired gas^2.5H post XXX challenge
C1977881|T201|COMP|50014-0|LNC|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript
C1977883|T201|COMP|50015-7|LNC|West Nile virus Ag|West Nile virus Ag
C1977884|T201|COMP|50016-5|LNC|Sugar|Sugar
C1977885|T201|COMP|50017-3|LNC|Hemoglobin.gastrointestinal|Hemoglobin.gastrointestinal
C1977887|T201|COMP|50018-1|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C1977888|T201|COMP|50019-9|LNC|HLA-DP+DQ+DR|HLA-DP+DQ+DR
C1977890|T201|COMP|50020-7|LNC|Microdeletion syndromes|Microdeletion syndromes
C1977891|T201|COMP|50021-5|LNC|oxyCODONE|oxyCODONE
C1977892|T201|COMP|50022-3|LNC|Ethanol+Methanol+Isopropyl alcohol+Acetone|Ethanol+Methanol+Isopropyl alcohol+Acetone
C1977893|T201|COMP|50023-1|LNC|Hepatitis C virus RNA panel|Hepatitis C virus RNA panel
C1977895|T201|COMP|50024-9|LNC|Virus identified|Virus identified
C1977896|T201|COMP|50050-4|LNC|Hemicystine/Amino acids.total|Hemicystine/Amino acids.total
C1977897|T201|COMP|50051-2|LNC|Hemicystine/Amino acids.total|Hemicystine/Amino acids.total
C1977898|T201|COMP|50052-0|LNC|Hemicystine/Amino acids.total|Hemicystine/Amino acids.total
C1977899|T201|COMP|50053-8|LNC|Hemicystine/Amino acids.total|Hemicystine/Amino acids.total
C1977900|T201|COMP|50054-6|LNC|Hemicystine/Creatinine|Hemicystine/Creatinine
C1977902|T201|COMP|50055-3|LNC|Iohexol renal clearance|Iohexol renal clearance
C1977904|T201|COMP|50056-1|LNC|Nutritional risk index|Nutritional risk index
C1977906|T201|COMP|50057-9|LNC|Fractional excretion of phosphate|Fractional excretion of phosphate
C1977908|T201|COMP|50058-7|LNC|Phosphate renal clearance|Phosphate renal clearance
C1977909|T201|COMP|50059-5|LNC|Protein fractions.oligoclonal bands/Protein.total|Protein fractions.oligoclonal bands/Protein.total
C1977911|T201|COMP|50060-3|LNC|Fatty acids.very long chain.C24:0/Creatinine|Fatty acids.very long chain.C24:0/Creatinine
C1977913|T201|COMP|50061-1|LNC|Tetradecanedioate/Creatinine|Tetradecanedioate/Creatinine
C1977915|T201|COMP|50062-9|LNC|Tetradecenedioate/Creatinine|Tetradecenedioate/Creatinine
C1977917|T201|COMP|50063-7|LNC|Urea renal clearance/1.73 sq M|Urea renal clearance/1.73 sq M
C1977920|T201|COMP|50065-2|LNC|1-Methylhistidine|1-Methylhistidine
C1977921|T201|COMP|50066-0|LNC|1-Methylhistidine|1-Methylhistidine
C1977922|T201|COMP|50067-8|LNC|11-Hydroxyandrostenedione|11-Hydroxyandrostenedione
C1977926|T201|COMP|50071-0|LNC|11-Deoxycortisol|11-Deoxycortisol
C1977927|T201|COMP|50072-8|LNC|11-Deoxycortisol^pre 250 ug corticotropin|11-Deoxycortisol^pre 250 ug corticotropin
C1977928|T201|COMP|50073-6|LNC|11-Deoxycortisol^30M post 250 ug corticotropin|11-Deoxycortisol^30M post 250 ug corticotropin
C1977929|T201|COMP|50074-4|LNC|11-Deoxycortisol^45M post 250 ug corticotropin|11-Deoxycortisol^45M post 250 ug corticotropin
C1977930|T201|COMP|50075-1|LNC|11-Deoxycortisol^1H post 250 ug corticotropin|11-Deoxycortisol^1H post 250 ug corticotropin
C1977931|T201|COMP|50076-9|LNC|17-Ketosteroids^post dose dexamethasone|17-Ketosteroids^post dose dexamethasone
C1977932|T201|COMP|50077-7|LNC|17-Ketosteroids^2D post dose dexamethasone|17-Ketosteroids^2D post dose dexamethasone
C1977933|T201|COMP|50078-5|LNC|17-Hydroxypregnenolone^pre 250 ug corticotropin|17-Hydroxypregnenolone^pre 250 ug corticotropin
C1977936|T201|COMP|50081-9|LNC|18-Hydroxydeoxycorticosterone|18-Hydroxydeoxycorticosterone
C1977937|T201|COMP|50082-7|LNC|18-Hydroxycorticosterone|18-Hydroxycorticosterone
C1977938|T201|COMP|50083-5|LNC|Alpha aminoadipate|Alpha aminoadipate
C1977939|T201|COMP|50084-3|LNC|Alpha aminoadipate|Alpha aminoadipate
C1977940|T201|COMP|50085-0|LNC|2-Methyl-3-Hydroxyvalerate/Creatinine|2-Methyl-3-Hydroxyvalerate/Creatinine
C1977942|T201|COMP|50086-8|LNC|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)
C1977944|T201|COMP|50087-6|LNC|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)
C1977945|T201|COMP|50088-4|LNC|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)
C1977946|T201|COMP|50089-2|LNC|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)
C1977947|T201|COMP|50090-0|LNC|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)|2-Methyl-3-Hydroxybutyrylcarnitine (C5-OH)
C1977950|T201|COMP|50092-6|LNC|2-Methylcitrate|2-Methylcitrate
C1977951|T201|COMP|50093-4|LNC|21-Deoxycortisol|21-Deoxycortisol
C1977952|T201|COMP|50094-2|LNC|21-Deoxycortisol^45M post 250 ug corticotropin|21-Deoxycortisol^45M post 250 ug corticotropin
C1977953|T201|COMP|50095-9|LNC|21-Deoxycortisol^pre 250 ug corticotropin|21-Deoxycortisol^pre 250 ug corticotropin
C1977954|T201|COMP|50096-7|LNC|21-Deoxycortisol^30M post 250 ug corticotropin|21-Deoxycortisol^30M post 250 ug corticotropin
C1977955|T201|COMP|50097-5|LNC|21-Deoxycortisol^1H post 250 ug corticotropin|21-Deoxycortisol^1H post 250 ug corticotropin
C1977956|T201|COMP|50098-3|LNC|3-Hydroxyvalerate|3-Hydroxyvalerate
C1977957|T201|COMP|50099-1|LNC|Beta hydroxybutyrate/Acetoacetate|Beta hydroxybutyrate/Acetoacetate
C1977959|T201|COMP|50100-7|LNC|Beta hydroxybutyrate/Acetoacetate|Beta hydroxybutyrate/Acetoacetate
C1977960|T201|COMP|50101-5|LNC|3-Hydroxybutyrylcarnitine (C4-OH)|3-Hydroxybutyrylcarnitine (C4-OH)
C1977961|T201|COMP|50102-3|LNC|3-Hydroxybutyrylcarnitine (C4-OH)|3-Hydroxybutyrylcarnitine (C4-OH)
C1977962|T201|COMP|50103-1|LNC|3-Hydroxybutyrylcarnitine (C4-OH)|3-Hydroxybutyrylcarnitine (C4-OH)
C1977963|T201|COMP|50104-9|LNC|3-Hydroxyisovalerylcarnitine (C5-OH)|3-Hydroxyisovalerylcarnitine (C5-OH)
C1977964|T201|COMP|50105-6|LNC|3-Hydroxyisovalerylcarnitine (C5-OH)|3-Hydroxyisovalerylcarnitine (C5-OH)
C1977965|T201|COMP|50106-4|LNC|3-Hydroxyisovalerylcarnitine (C5-OH)|3-Hydroxyisovalerylcarnitine (C5-OH)
C1977966|T201|COMP|50107-2|LNC|3-Hydroxyisovalerylcarnitine (C5-OH)|3-Hydroxyisovalerylcarnitine (C5-OH)
C1977967|T201|COMP|50108-0|LNC|3-Hydroxylinoleoylcarnitine (C18:2-OH)|3-Hydroxylinoleoylcarnitine (C18:2-OH)
C1977968|T201|COMP|50109-8|LNC|3-Hydroxylinoleoylcarnitine (C18:2-OH)|3-Hydroxylinoleoylcarnitine (C18:2-OH)
C1977969|T201|COMP|50110-6|LNC|3-Hydroxylinoleoylcarnitine (C18:2-OH)|3-Hydroxylinoleoylcarnitine (C18:2-OH)
C1977970|T201|COMP|50111-4|LNC|3-Hydroxylinoleoylcarnitine (C18:2-OH)|3-Hydroxylinoleoylcarnitine (C18:2-OH)
C1977971|T201|COMP|50112-2|LNC|3-Hydroxylinoleoylcarnitine (C18:2-OH)/Creatinine|3-Hydroxylinoleoylcarnitine (C18:2-OH)/Creatinine
C1977973|T201|COMP|50113-0|LNC|3-Hydroxyoleoylcarnitine (C18:1-OH)|3-Hydroxyoleoylcarnitine (C18:1-OH)
C1977974|T201|COMP|50114-8|LNC|3-Hydroxyoleoylcarnitine (C18:1-OH)|3-Hydroxyoleoylcarnitine (C18:1-OH)
C1977975|T201|COMP|50115-5|LNC|3-Hydroxyoleoylcarnitine (C18:1-OH)|3-Hydroxyoleoylcarnitine (C18:1-OH)
C1977976|T201|COMP|50116-3|LNC|3-Hydroxyoleoylcarnitine (C18:1-OH)|3-Hydroxyoleoylcarnitine (C18:1-OH)
C1977977|T201|COMP|50117-1|LNC|3-Hydroxyoleoylcarnitine (C18:1-OH)/Creatinine|3-Hydroxyoleoylcarnitine (C18:1-OH)/Creatinine
C1977979|T201|COMP|50118-9|LNC|3-Hydroxypalmitoleylcarnitine (C16:1-OH)|3-Hydroxypalmitoleylcarnitine (C16:1-OH)
C1977980|T201|COMP|50119-7|LNC|3-Hydroxypalmitoleylcarnitine (C16:1-OH)|3-Hydroxypalmitoleylcarnitine (C16:1-OH)
C1977981|T201|COMP|50120-5|LNC|3-Hydroxypalmitoleylcarnitine (C16:1-OH)|3-Hydroxypalmitoleylcarnitine (C16:1-OH)
C1977982|T201|COMP|50121-3|LNC|3-Hydroxypalmitoleylcarnitine (C16:1-OH)|3-Hydroxypalmitoleylcarnitine (C16:1-OH)
C1977985|T201|COMP|50132-0|LNC|3-Hydroxystearoylcarnitine (C18-OH)|3-Hydroxystearoylcarnitine (C18-OH)
C1977986|T201|COMP|50133-8|LNC|3-Hydroxystearoylcarnitine (C18-OH)|3-Hydroxystearoylcarnitine (C18-OH)
C1977987|T201|COMP|50134-6|LNC|3-Hydroxystearoylcarnitine (C18-OH)/Creatinine|3-Hydroxystearoylcarnitine (C18-OH)/Creatinine
C1977989|T201|COMP|50135-3|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C1977990|T201|COMP|50136-1|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C1977991|T201|COMP|50137-9|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C1977992|T201|COMP|50138-7|LNC|3-Methoxy-4-Hydroxyphenylglycol/Creatinine|3-Methoxy-4-Hydroxyphenylglycol/Creatinine
C1977994|T201|COMP|50139-5|LNC|3-Methoxytyramine|3-Methoxytyramine
C1977995|T201|COMP|50140-3|LNC|3-Methoxytyramine|3-Methoxytyramine
C1977996|T201|COMP|50141-1|LNC|3-O-Methyldopa|3-O-Methyldopa
C1977997|T201|COMP|50142-9|LNC|3-O-Methyldopa|3-O-Methyldopa
C1977998|T201|COMP|50143-7|LNC|3-O-Methyldopa|3-O-Methyldopa
C1977999|T201|COMP|50144-5|LNC|3-O-Methyldopa/Creatinine|3-O-Methyldopa/Creatinine
C1978001|T201|COMP|50145-2|LNC|3-Dechloroethylifosfamide^pre dose ifosfamide|3-Dechloroethylifosfamide^pre dose ifosfamide
C1978002|T201|COMP|50146-0|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C1978003|T201|COMP|50147-8|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C1978004|T201|COMP|50148-6|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C1978005|T201|COMP|50149-4|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C1978006|T201|COMP|50150-2|LNC|5-Hydroxytryptophan|5-Hydroxytryptophan
C1978007|T201|COMP|50151-0|LNC|5-Hydroxytryptophan|5-Hydroxytryptophan
C1978008|T201|COMP|50152-8|LNC|5-Hydroxytryptophan/Creatinine|5-Hydroxytryptophan/Creatinine
C1978010|T201|COMP|50153-6|LNC|5-Methyltetrahydrofolate|5-Methyltetrahydrofolate
C1978011|T201|COMP|50154-4|LNC|Acetoacetate|Acetoacetate
C1978012|T201|COMP|50155-1|LNC|Acetylcarnitine (C2)|Acetylcarnitine (C2)
C1978013|T201|COMP|50156-9|LNC|Acetylcarnitine (C2)|Acetylcarnitine (C2)
C1978014|T201|COMP|50157-7|LNC|Acetylcarnitine (C2)|Acetylcarnitine (C2)
C1978015|T201|COMP|50158-5|LNC|Acetylcarnitine (C2)|Acetylcarnitine (C2)
C1978016|T201|COMP|50159-3|LNC|Acetylcarnitine (C2)/Creatinine|Acetylcarnitine (C2)/Creatinine
C1978018|T201|COMP|50160-1|LNC|Amino acids|Amino acids
C1978019|T201|COMP|50161-9|LNC|Organic acids pattern|Organic acids pattern
C1978020|T201|COMP|50162-7|LNC|Acylcarnitine|Acylcarnitine
C1978021|T201|COMP|50163-5|LNC|Acylcarnitine|Acylcarnitine
C1978022|T201|COMP|50164-3|LNC|Acylcarnitine pattern|Acylcarnitine pattern
C1978023|T201|COMP|50165-0|LNC|Adenine phosphoribosyltransferase|Adenine phosphoribosyltransferase
C1978024|T201|COMP|50166-8|LNC|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)
C1978026|T201|COMP|50167-6|LNC|Alanine|Alanine
C1978027|T201|COMP|50168-4|LNC|Alanine aminotransferase|Alanine aminotransferase
C1978028|T201|COMP|50169-2|LNC|Aldosterone^post XXX challenge|Aldosterone^post XXX challenge
C1978029|T201|COMP|50170-0|LNC|Aldosterone^pre XXX challenge|Aldosterone^pre XXX challenge
C1978030|T201|COMP|50171-8|LNC|Aldosterone^pre 250 ug corticotropin IM|Aldosterone^pre 250 ug corticotropin IM
C1978031|T201|COMP|50172-6|LNC|Aldosterone^30M post 250 ug corticotropin IM|Aldosterone^30M post 250 ug corticotropin IM
C1978032|T201|COMP|50173-4|LNC|Aldosterone^1H post 250 ug corticotropin IM|Aldosterone^1H post 250 ug corticotropin IM
C1978034|T201|COMP|50196-5|LNC|Occult blood panel|Occult blood panel
C1978035|T201|COMP|50197-3|LNC|aPTT panel|aPTT panel
C1978037|T201|COMP|50198-1|LNC|Iron^1st specimen|Iron^1st specimen
C1978038|T201|COMP|50199-9|LNC|Iron^2nd specimen|Iron^2nd specimen
C1978039|T201|COMP|50200-5|LNC|Iron^3rd specimen|Iron^3rd specimen
C1978040|T201|COMP|50201-3|LNC|Iron^4th specimen|Iron^4th specimen
C1978041|T201|COMP|50210-4|LNC|Glomerular filtration rate/1.73 sq M.predicted|Glomerular filtration rate/1.73 sq M.predicted
C1978045|T201|COMP|50212-0|LNC|Glucose^2nd specimen|Glucose^2nd specimen
C1978046|T201|COMP|50213-8|LNC|Glucose^3rd specimen|Glucose^3rd specimen
C1978047|T201|COMP|50214-6|LNC|Glucose^4th specimen|Glucose^4th specimen
C1978048|T201|COMP|50215-3|LNC|Glucose^5th specimen|Glucose^5th specimen
C1978049|T201|COMP|50216-1|LNC|Glucose^6th specimen|Glucose^6th specimen
C1978050|T201|COMP|50217-9|LNC|Glucose^8th specimen|Glucose^8th specimen
C1978051|T201|COMP|50218-7|LNC|Glucose^9th specimen|Glucose^9th specimen
C1978052|T201|COMP|50219-5|LNC|Respiratory pathogens DNA & RNA 12a panel|Respiratory pathogens DNA & RNA 12a panel
C1978054|T201|COMP|50220-3|LNC|Collection interval from baseline|Collection interval from baseline
C1978056|T201|COMP|50221-1|LNC|Bacteria|Bacteria
C1978057|T201|COMP|50222-9|LNC|Broad casts|Broad casts
C1978058|T201|COMP|50223-7|LNC|Cholesterol crystals|Cholesterol crystals
C1978059|T201|COMP|50224-5|LNC|Epithelial casts|Epithelial casts
C1978060|T201|COMP|50225-2|LNC|Epithelial cells.non-squamous|Epithelial cells.non-squamous
C1978061|T201|COMP|50226-0|LNC|Erythrocyte clumps|Erythrocyte clumps
C1978063|T201|COMP|50228-6|LNC|Oval fat bodies (globules)|Oval fat bodies (globules)
C1978064|T201|COMP|50229-4|LNC|Fatty casts|Fatty casts
C1978065|T201|COMP|50230-2|LNC|Granular casts|Granular casts
C1978066|T201|COMP|50231-0|LNC|Hyaline casts|Hyaline casts
C1978067|T201|COMP|50232-8|LNC|Leucine crystals|Leucine crystals
C1978068|T201|COMP|50233-6|LNC|Leukocyte clumps|Leukocyte clumps
C1978069|T201|COMP|50234-4|LNC|Mixed cellular casts|Mixed cellular casts
C1978070|T201|COMP|50235-1|LNC|Mucus|Mucus
C1978071|T201|COMP|50236-9|LNC|Phosphate crystals.amorphous|Phosphate crystals.amorphous
C1978072|T201|COMP|50237-7|LNC|Trichomonas sp|Trichomonas sp
C1978073|T201|COMP|50238-5|LNC|Tyrosine crystals|Tyrosine crystals
C1978074|T201|COMP|50239-3|LNC|Urate crystals.amorphous|Urate crystals.amorphous
C1978075|T201|COMP|50240-1|LNC|Yeast.budding|Yeast.budding
C1978076|T201|COMP|50241-9|LNC|17-Ketosteroids^post high dose dexamethasone|17-Ketosteroids^post high dose dexamethasone
C1978077|T201|COMP|50242-7|LNC|17-Ketosteroids^2D post high dose dexamethasone|17-Ketosteroids^2D post high dose dexamethasone
C1978078|T201|COMP|50243-5|LNC|17-Ketosteroids^post dose dexamethasone|17-Ketosteroids^post dose dexamethasone
C1978079|T201|COMP|50244-3|LNC|17-Ketosteroids^2D post dose dexamethasone|17-Ketosteroids^2D post dose dexamethasone
C1978082|T201|COMP|50247-6|LNC|17-Hydroxycorticosteroids^post dose dexamethasone|17-Hydroxycorticosteroids^post dose dexamethasone
C1978085|T201|COMP|50250-0|LNC|21-Deoxycortisol|21-Deoxycortisol
C1978086|T201|COMP|50251-8|LNC|3-Hydroxybutyrylcarnitine (C4-OH)/Creatinine|3-Hydroxybutyrylcarnitine (C4-OH)/Creatinine
C1978088|T201|COMP|50252-6|LNC|3-Hydroxyisovalerylcarnitine (C5-OH)/Creatinine|3-Hydroxyisovalerylcarnitine (C5-OH)/Creatinine
C1978090|T201|COMP|50253-4|LNC|Fatty acids.nonesterified^1st specimen post CFst|Fatty acids.nonesterified^1st specimen post CFst
C1978091|T201|COMP|50254-2|LNC|Fatty acids.nonesterified^2nd specimen post CFst|Fatty acids.nonesterified^2nd specimen post CFst
C1978092|T201|COMP|50255-9|LNC|Fatty acids.nonesterified^3rd specimen post CFst|Fatty acids.nonesterified^3rd specimen post CFst
C1978093|T201|COMP|50256-7|LNC|Fatty acids.nonesterified^4th specimen post CFst|Fatty acids.nonesterified^4th specimen post CFst
C1978094|T201|COMP|50257-5|LNC|Fatty acids.nonesterified^5th specimen post CFst|Fatty acids.nonesterified^5th specimen post CFst
C1978095|T201|COMP|50258-3|LNC|Aldosterone^post 25 mg captopril PO|Aldosterone^post 25 mg captopril PO
C1978096|T201|COMP|50259-1|LNC|Aldosterone^pre 25 mg captopril PO|Aldosterone^pre 25 mg captopril PO
C1978097|T201|COMP|50260-9|LNC|Prekeratocytes|Prekeratocytes
C1978101|T201|COMP|50262-5|LNC|Reticulocytes panel|Reticulocytes panel
C1978103|T201|COMP|50263-3|LNC|17-Ketosteroids^post high dose dexamethasone|17-Ketosteroids^post high dose dexamethasone
C1978104|T201|COMP|50264-1|LNC|17-Ketosteroids^2D post high dose dexamethasone|17-Ketosteroids^2D post high dose dexamethasone
C1978105|T201|COMP|50265-8|LNC|2-Dechloroethylifosfamide^pre dose ifosfamide|2-Dechloroethylifosfamide^pre dose ifosfamide
C1978106|T201|COMP|50266-6|LNC|2-Dechloroethylifosfamide^1D post dose ifosfamide|2-Dechloroethylifosfamide^1D post dose ifosfamide
C1978107|T201|COMP|50267-4|LNC|2-Dechloroethylifosfamide^2D post dose ifosfamide|2-Dechloroethylifosfamide^2D post dose ifosfamide
C1978108|T201|COMP|50268-2|LNC|2-Dechloroethylifosfamide^3D post dose ifosfamide|2-Dechloroethylifosfamide^3D post dose ifosfamide
C1978109|T201|COMP|50269-0|LNC|2-Dechloroethylifosfamide^4D post dose ifosfamide|2-Dechloroethylifosfamide^4D post dose ifosfamide
C1978110|T201|COMP|50270-8|LNC|2-Dechloroethylifosfamide^5D post dose ifosfamide|2-Dechloroethylifosfamide^5D post dose ifosfamide
C1978111|T201|COMP|50271-6|LNC|2-Dechloroethylifosfamide^3H post dose ifosfamide|2-Dechloroethylifosfamide^3H post dose ifosfamide
C1978112|T201|COMP|50272-4|LNC|2-Dechloroethylifosfamide^6H post dose ifosfamide|2-Dechloroethylifosfamide^6H post dose ifosfamide
C1978113|T201|COMP|50273-2|LNC|3-Hydroxymyristoleylcarnitine (C14:1-OH)|3-Hydroxymyristoleylcarnitine (C14:1-OH)
C1978115|T201|COMP|50274-0|LNC|3-Hydroxymyristoleylcarnitine (C14:1-OH)|3-Hydroxymyristoleylcarnitine (C14:1-OH)
C1978116|T201|COMP|50275-7|LNC|3-Hydroxymyristoleylcarnitine (C14:1-OH)|3-Hydroxymyristoleylcarnitine (C14:1-OH)
C1978117|T201|COMP|50276-5|LNC|3-Hydroxymyristoleylcarnitine (C14:1-OH)|3-Hydroxymyristoleylcarnitine (C14:1-OH)
C1978118|T201|COMP|50277-3|LNC|3-Hydroxymyristoleylcarnitine (C14:1-OH)|3-Hydroxymyristoleylcarnitine (C14:1-OH)
C1978121|T201|COMP|50279-9|LNC|3-Hydroxytetradecanoylcarnitine (C14-OH)|3-Hydroxytetradecanoylcarnitine (C14-OH)
C1978122|T201|COMP|50280-7|LNC|3-Hydroxytetradecanoylcarnitine (C14-OH)|3-Hydroxytetradecanoylcarnitine (C14-OH)
C1978123|T201|COMP|50281-5|LNC|3-Hydroxytetradecanoylcarnitine (C14-OH)|3-Hydroxytetradecanoylcarnitine (C14-OH)
C1978124|T201|COMP|50282-3|LNC|3-Hydroxytetradecanoylcarnitine (C14-OH)|3-Hydroxytetradecanoylcarnitine (C14-OH)
C1978125|T201|COMP|50283-1|LNC|3-Hydroxytetradecanoylcarnitine|3-Hydroxytetradecanoylcarnitine
C1978128|T201|COMP|50285-6|LNC|3-Dechloroethylifosfamide^1D post dose ifosfamide|3-Dechloroethylifosfamide^1D post dose ifosfamide
C1978129|T201|COMP|50286-4|LNC|3-Dechloroethylifosfamide^2D post dose ifosfamide|3-Dechloroethylifosfamide^2D post dose ifosfamide
C1978130|T201|COMP|50287-2|LNC|3-Dechloroethylifosfamide^3D post dose ifosfamide|3-Dechloroethylifosfamide^3D post dose ifosfamide
C1978131|T201|COMP|50288-0|LNC|3-Dechloroethylifosfamide^4D post dose ifosfamide|3-Dechloroethylifosfamide^4D post dose ifosfamide
C1978132|T201|COMP|50289-8|LNC|3-Dechloroethylifosfamide^6D post dose ifosfamide|3-Dechloroethylifosfamide^6D post dose ifosfamide
C1978133|T201|COMP|50290-6|LNC|3-Dechloroethylifosfamide^3H post dose ifosfamide|3-Dechloroethylifosfamide^3H post dose ifosfamide
C1978134|T201|COMP|50291-4|LNC|3-Dechloroethylifosfamide^6H post dose ifosfamide|3-Dechloroethylifosfamide^6H post dose ifosfamide
C1978135|T201|COMP|50292-2|LNC|4-Hydroxyifosfamide^pre dose ifosfamide|4-Hydroxyifosfamide^pre dose ifosfamide
C1978136|T201|COMP|50293-0|LNC|4-Hydroxyifosfamide^1D post dose ifosfamide|4-Hydroxyifosfamide^1D post dose ifosfamide
C1978137|T201|COMP|50294-8|LNC|4-Hydroxyifosfamide^2D post dose ifosfamide|4-Hydroxyifosfamide^2D post dose ifosfamide
C1978138|T201|COMP|50295-5|LNC|4-Hydroxyifosfamide^3D post dose ifosfamide|4-Hydroxyifosfamide^3D post dose ifosfamide
C1978139|T201|COMP|50296-3|LNC|4-Hydroxyifosfamide^4D post dose ifosfamide|4-Hydroxyifosfamide^4D post dose ifosfamide
C1978140|T201|COMP|50297-1|LNC|4-Hydroxyifosfamide^5D post dose ifosfamide|4-Hydroxyifosfamide^5D post dose ifosfamide
C1978141|T201|COMP|50298-9|LNC|4-Hydroxyifosfamide^3H post dose ifosfamide|4-Hydroxyifosfamide^3H post dose ifosfamide
C1978142|T201|COMP|50299-7|LNC|4-Hydroxyifosfamide^6H post dose ifosfamide|4-Hydroxyifosfamide^6H post dose ifosfamide
C1978143|T201|COMP|50300-3|LNC|6-Hydroxyheptanoate|6-Hydroxyheptanoate
C1978145|T201|COMP|50301-1|LNC|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)
C1978146|T201|COMP|50302-9|LNC|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)
C1978147|T201|COMP|50303-7|LNC|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)
C1978148|T201|COMP|50304-5|LNC|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)|Adipoylcarnitine+Methylglutarylcarnitine (C6-DC)
C1978151|T201|COMP|50306-0|LNC|Allantoine|Allantoine
C1978153|T201|COMP|50307-8|LNC|BCL10 Ag|BCL10 Ag
C1978155|T201|COMP|50308-6|LNC|Caldesmon Ag|Caldesmon Ag
C1978157|T201|COMP|50309-4|LNC|CD138 Ag|CD138 Ag
C1978158|T201|COMP|50310-2|LNC|CD7 Ag|CD7 Ag
C1978159|T201|COMP|50311-0|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1978160|T201|COMP|50312-8|LNC|Clusterin Ag|Clusterin Ag
C1978162|T201|COMP|50313-6|LNC|Cyclospora sp identified|Cyclospora sp identified
C1978163|T201|COMP|50323-5|LNC|MSH-2 Ag|MSH-2 Ag
C1978165|T201|COMP|50324-3|LNC|MSH-6 Ag|MSH-6 Ag
C1978167|T201|COMP|50325-0|LNC|MUM-1 Ag|MUM-1 Ag
C1978169|T201|COMP|50326-8|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C1978170|T201|COMP|50327-6|LNC|Neu-N Ag|Neu-N Ag
C1978172|T201|COMP|50328-4|LNC|PMS-2 Ag|PMS-2 Ag
C1978174|T201|COMP|50329-2|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C1978175|T201|COMP|50330-0|LNC|SLC6A4 gene targeted mutation analysis|SLC6A4 gene targeted mutation analysis
C1978177|T201|COMP|50331-8|LNC|WT-1 Ag|WT-1 Ag
C1978179|T201|COMP|50332-6|LNC|Hexadecanedioate/Creatinine|Hexadecanedioate/Creatinine
C1978180|T201|COMP|50333-4|LNC|Tetradecanedioate/Creatinine|Tetradecanedioate/Creatinine
C1978181|T201|COMP|50334-2|LNC|Acylglycines panel|Acylglycines panel
C1978183|T201|COMP|50335-9|LNC|Alpha-beta crystallin Ag|Alpha-beta crystallin Ag
C1978185|T201|COMP|50336-7|LNC|Beta cortolone/Cortisol|Beta cortolone/Cortisol
C1978187|T201|COMP|50337-5|LNC|carBAMazepine free & total & 10,11-Epoxide panel|carBAMazepine free & total & 10,11-Epoxide panel
C1978189|T201|COMP|50338-3|LNC|Cannabinoids|Cannabinoids
C1978190|T201|COMP|50339-1|LNC|Cholesterol|Cholesterol
C1978191|T201|COMP|50340-9|LNC|Eosinophils|Eosinophils
C1978192|T201|COMP|50341-7|LNC|Eosinophils|Eosinophils
C1978193|T201|COMP|50342-5|LNC|Ependymal+Choroid plexus cells/100 leukocytes|Ependymal+Choroid plexus cells/100 leukocytes
C1978195|T201|COMP|50343-3|LNC|Ethanol|Ethanol
C1978196|T201|COMP|50344-1|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1978197|T201|COMP|50345-8|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1978198|T201|COMP|50346-6|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1978199|T201|COMP|50347-4|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1978200|T201|COMP|50348-2|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1978201|T201|COMP|50349-0|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C1978202|T201|COMP|50350-8|LNC|Mustard Ab.IgE/IgE.total|Mustard Ab.IgE/IgE.total
C1978203|T201|COMP|50351-6|LNC|Casuarina equisetifolia Ab.IgE/IgE.total|Casuarina equisetifolia Ab.IgE/IgE.total
C1978204|T201|COMP|50352-4|LNC|Papain Ab.IgE/IgE.total|Papain Ab.IgE/IgE.total
C1978205|T201|COMP|50353-2|LNC|Parrot feather Ab.IgE/IgE.total|Parrot feather Ab.IgE/IgE.total
C1978206|T201|COMP|50354-0|LNC|Paspalum notatum Ab.IgE/IgE.total|Paspalum notatum Ab.IgE/IgE.total
C1978207|T201|COMP|50355-7|LNC|Perca spp Ab.IgE/IgE.total|Perca spp Ab.IgE/IgE.total
C1978208|T201|COMP|50356-5|LNC|Phalaris arundinacea Ab.IgE/IgE.total|Phalaris arundinacea Ab.IgE/IgE.total
C1978209|T201|COMP|50357-3|LNC|Phenolphthalein|Phenolphthalein
C1978210|T201|COMP|50358-1|LNC|Phenylacetate/Creatinine|Phenylacetate/Creatinine
C1978211|T201|COMP|50359-9|LNC|Phenyllactate/Creatinine|Phenyllactate/Creatinine
C1978212|T201|COMP|50360-7|LNC|Phenylpropionylglycine/Creatinine|Phenylpropionylglycine/Creatinine
C1978213|T201|COMP|50361-5|LNC|Phenylpyruvate/Creatinine|Phenylpyruvate/Creatinine
C1978214|T201|COMP|50362-3|LNC|Phoma betae Ab.IgE/IgE.total|Phoma betae Ab.IgE/IgE.total
C1978215|T201|COMP|50363-1|LNC|Pigweed common Ab.IgE/IgE.total|Pigweed common Ab.IgE/IgE.total
C1978216|T201|COMP|50364-9|LNC|Piper nigrum Ab.IgE/IgE.total|Piper nigrum Ab.IgE/IgE.total
C1978217|T201|COMP|50365-6|LNC|Platelet glycoprotein IIb-IIIa Ab|Platelet glycoprotein IIb-IIIa Ab
C1978218|T201|COMP|50366-4|LNC|Prolactin.monomeric/Prolactin.total|Prolactin.monomeric/Prolactin.total
C1978220|T201|COMP|50367-2|LNC|Propionylglycine/Creatinine|Propionylglycine/Creatinine
C1978221|T201|COMP|50368-0|LNC|Protoporphyrin|Protoporphyrin
C1978222|T201|COMP|50369-8|LNC|Quercus alba Ab.IgE/IgE.total|Quercus alba Ab.IgE/IgE.total
C1978223|T201|COMP|50370-6|LNC|Syagrus romanzoffianum Ab.IgE/IgE.total|Syagrus romanzoffianum Ab.IgE/IgE.total
C1978224|T201|COMP|50371-4|LNC|Protoporphyrin|Protoporphyrin
C1978225|T201|COMP|50372-2|LNC|Protoporphyrin|Protoporphyrin
C1978226|T201|COMP|50373-0|LNC|Eosinophils.band form/100 cells|Eosinophils.band form/100 cells
C1978228|T201|COMP|50374-8|LNC|Myelocytes.eosinophilic/100 cells|Myelocytes.eosinophilic/100 cells
C1978230|T201|COMP|50375-5|LNC|Nucleated cells|Nucleated cells
C1978237|T201|COMP|50379-7|LNC|Creatinine dialysis fluid clearance/1.73 sq M|Creatinine dialysis fluid clearance/1.73 sq M
C1978242|T201|COMP|50382-1|LNC|Glutathione reductase|Glutathione reductase
C1978243|T201|COMP|50383-9|LNC|Glomerular filtration rate.predicted|Glomerular filtration rate.predicted
C1978244|T201|COMP|50384-7|LNC|Glomerular filtration rate/1.73 sq M.predicted|Glomerular filtration rate/1.73 sq M.predicted
C1978245|T201|COMP|50385-4|LNC|Alpha-1-Microglobulin.placental|Alpha-1-Microglobulin.placental
C1978247|T201|COMP|50386-2|LNC|Parakeet+Parrot droppings Ab.IgE/IgE.total|Parakeet+Parrot droppings Ab.IgE/IgE.total
C1978249|T201|COMP|50387-0|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1978250|T201|COMP|50388-8|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1978252|T201|COMP|50390-4|LNC|Coagulation factor II circulating inhibitor|Coagulation factor II circulating inhibitor
C1978254|T201|COMP|50391-2|LNC|Coagulation surface induced circulating inhibitor|Coagulation surface induced circulating inhibitor
C1978256|T201|COMP|50392-0|LNC|3-Keto n-Valerate|3-Keto n-Valerate
C1978258|T201|COMP|50393-8|LNC|3-Keto n-Valerate/Creatinine|3-Keto n-Valerate/Creatinine
C1978260|T201|COMP|50394-6|LNC|Adenine phosphoribosyltransferase|Adenine phosphoribosyltransferase
C1978261|T201|COMP|50395-3|LNC|Adenosine deaminase|Adenosine deaminase
C1978262|T201|COMP|50396-1|LNC|Molecular diagnostic major findings for display|Molecular diagnostic major findings for display
C1978264|T201|COMP|50397-9|LNC|Molecular diagnostic overall interpretation|Molecular diagnostic overall interpretation
C1978266|T201|COMP|50398-7|LNC|Narrative diagnostic report|Narrative diagnostic report
C1978268|T201|COMP|50399-5|LNC|Clinical genetic report summary panel|Clinical genetic report summary panel
C1978271|T201|COMP|50401-9|LNC|Blood group antibody titered|Blood group antibody titered
C1978274|T201|COMP|50404-3|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C1978276|T201|COMP|50405-0|LNC|Patient symptoms^post transfusion reaction|Patient symptoms^post transfusion reaction
C1978277|T201|COMP|50406-8|LNC|Cannabinoids|Cannabinoids
C1978278|T201|COMP|50407-6|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C1978279|T201|COMP|50408-4|LNC|Protein.abnormal band/Protein.total|Protein.abnormal band/Protein.total
C1978281|T201|COMP|50409-2|LNC|Cholesterol.in HDL 2+3|Cholesterol.in HDL 2+3
C1978285|T201|COMP|50411-8|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1978286|T201|COMP|50412-6|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1978287|T201|COMP|50413-4|LNC|Corticotropin^pre 1 mg dexamethasone PO overnight|Corticotropin^pre 1 mg dexamethasone PO overnight
C1978289|T201|COMP|50415-9|LNC|Cortisol^pre 2 mg dexamethasone PO overnight|Cortisol^pre 2 mg dexamethasone PO overnight
C1978290|T201|COMP|50416-7|LNC|Cortisol^post 2 mg dexamethasone PO overnight|Cortisol^post 2 mg dexamethasone PO overnight
C1978291|T201|COMP|50417-5|LNC|Corticotropin^pre 2 mg dexamethasone PO overnight|Corticotropin^pre 2 mg dexamethasone PO overnight
C1978295|T201|COMP|50421-7|LNC|Cortisol^pre 100 ug CRH IV|Cortisol^pre 100 ug CRH IV
C1978296|T201|COMP|50422-5|LNC|Cortisol^20M post 100 ug CRH IV|Cortisol^20M post 100 ug CRH IV
C1978297|T201|COMP|50423-3|LNC|Cortisol^40M post 100 ug CRH IV|Cortisol^40M post 100 ug CRH IV
C1978298|T201|COMP|50424-1|LNC|Cortisol^1H post 100 ug CRH IV|Cortisol^1H post 100 ug CRH IV
C1978299|T201|COMP|50425-8|LNC|Corticotropin^pre 100 ug CRH IV|Corticotropin^pre 100 ug CRH IV
C1978300|T201|COMP|50426-6|LNC|Corticotropin^20M post 100 ug CRH IV|Corticotropin^20M post 100 ug CRH IV
C1978301|T201|COMP|50427-4|LNC|Corticotropin^40M post 100 ug CRH IV|Corticotropin^40M post 100 ug CRH IV
C1978302|T201|COMP|50428-2|LNC|Corticotropin^1H post 100 ug CRH IV|Corticotropin^1H post 100 ug CRH IV
C1978303|T201|COMP|50429-0|LNC|Cortisol^9 AM specimen|Cortisol^9 AM specimen
C1978304|T201|COMP|50430-8|LNC|Cortisol^3 PM specimen|Cortisol^3 PM specimen
C1978305|T201|COMP|50431-6|LNC|Cortisol^6 PM specimen|Cortisol^6 PM specimen
C1978306|T201|COMP|50432-4|LNC|Cortisol^9 PM specimen|Cortisol^9 PM specimen
C1978307|T201|COMP|50433-2|LNC|Cortisol^3 AM specimen|Cortisol^3 AM specimen
C1978308|T201|COMP|50434-0|LNC|Cortisol^6 AM specimen|Cortisol^6 AM specimen
C1978309|T201|COMP|50435-7|LNC|Corticotropin^9 AM specimen|Corticotropin^9 AM specimen
C1978310|T201|COMP|50436-5|LNC|Corticotropin^3 PM specimen|Corticotropin^3 PM specimen
C1978311|T201|COMP|50437-3|LNC|Corticotropin^6 PM specimen|Corticotropin^6 PM specimen
C1978312|T201|COMP|50438-1|LNC|Corticotropin^9 PM specimen|Corticotropin^9 PM specimen
C1978313|T201|COMP|50439-9|LNC|Corticotropin^3 AM specimen|Corticotropin^3 AM specimen
C1978314|T201|COMP|50440-7|LNC|Corticotropin^6 AM specimen|Corticotropin^6 AM specimen
C1978315|T201|COMP|50441-5|LNC|Cortisol^30M pre dose insulin IV|Cortisol^30M pre dose insulin IV
C1978316|T201|COMP|50442-3|LNC|Cortisol^20M post dose insulin IV|Cortisol^20M post dose insulin IV
C1978317|T201|COMP|50443-1|LNC|Somatotropin^30M pre dose arginine|Somatotropin^30M pre dose arginine
C1978318|T201|COMP|50444-9|LNC|Somatotropin^20M post dose arginine|Somatotropin^20M post dose arginine
C1978319|T201|COMP|50445-6|LNC|Corticotropin^1st specimen|Corticotropin^1st specimen
C1978320|T201|COMP|50446-4|LNC|Corticotropin^2nd specimen|Corticotropin^2nd specimen
C1978321|T201|COMP|50447-2|LNC|Corticotropin^3rd specimen|Corticotropin^3rd specimen
C1978322|T201|COMP|50448-0|LNC|Corticotropin^4th specimen|Corticotropin^4th specimen
C1978323|T201|COMP|50449-8|LNC|Corticotropin^5th specimen|Corticotropin^5th specimen
C1978324|T201|COMP|50450-6|LNC|Corticotropin^6th specimen|Corticotropin^6th specimen
C1978325|T201|COMP|50451-4|LNC|Corticotropin^7th specimen|Corticotropin^7th specimen
C1978326|T201|COMP|50452-2|LNC|Corticotropin^8th specimen|Corticotropin^8th specimen
C1978327|T201|COMP|50453-0|LNC|Cortisol^1st specimen|Cortisol^1st specimen
C1978328|T201|COMP|50454-8|LNC|Cortisol^2nd specimen|Cortisol^2nd specimen
C1978329|T201|COMP|50455-5|LNC|Cortisol^3rd specimen|Cortisol^3rd specimen
C1978330|T201|COMP|50456-3|LNC|Cortisol^4th specimen|Cortisol^4th specimen
C1978331|T201|COMP|50457-1|LNC|Cortisol^5th specimen|Cortisol^5th specimen
C1978332|T201|COMP|50458-9|LNC|Cortisol^6th specimen|Cortisol^6th specimen
C1978333|T201|COMP|50459-7|LNC|Cortisol^7th specimen|Cortisol^7th specimen
C1978334|T201|COMP|50460-5|LNC|Cortisol^8th specimen|Cortisol^8th specimen
C1978335|T201|COMP|50461-3|LNC|C peptide^1st specimen|C peptide^1st specimen
C1978336|T201|COMP|50462-1|LNC|C peptide^2nd specimen|C peptide^2nd specimen
C1978337|T201|COMP|50463-9|LNC|C peptide^3rd specimen|C peptide^3rd specimen
C1978338|T201|COMP|50464-7|LNC|C peptide^4th specimen|C peptide^4th specimen
C1978339|T201|COMP|50465-4|LNC|C peptide^5th specimen|C peptide^5th specimen
C1978340|T201|COMP|50466-2|LNC|C peptide^6th specimen|C peptide^6th specimen
C1978341|T201|COMP|50467-0|LNC|C peptide^7th specimen|C peptide^7th specimen
C1978342|T201|COMP|50468-8|LNC|C peptide^8th specimen|C peptide^8th specimen
C1978343|T201|COMP|50469-6|LNC|Calcitonin^1st specimen|Calcitonin^1st specimen
C1978344|T201|COMP|50470-4|LNC|Calcitonin^2nd specimen|Calcitonin^2nd specimen
C1978345|T201|COMP|50471-2|LNC|Calcitonin^3rd specimen|Calcitonin^3rd specimen
C1978346|T201|COMP|50472-0|LNC|Calcitonin^4th specimen|Calcitonin^4th specimen
C1978347|T201|COMP|50473-8|LNC|Calcitonin^5th specimen|Calcitonin^5th specimen
C1978348|T201|COMP|50474-6|LNC|Calcitonin^6th specimen|Calcitonin^6th specimen
C1978349|T201|COMP|50475-3|LNC|Calcitonin^7th specimen|Calcitonin^7th specimen
C1978350|T201|COMP|50476-1|LNC|Calcitonin^8th specimen|Calcitonin^8th specimen
C1978351|T201|COMP|50477-9|LNC|Follitropin^1st specimen|Follitropin^1st specimen
C1978352|T201|COMP|50478-7|LNC|Follitropin^2nd specimen|Follitropin^2nd specimen
C1978353|T201|COMP|50479-5|LNC|Follitropin^3rd specimen|Follitropin^3rd specimen
C1978354|T201|COMP|50480-3|LNC|Follitropin^4th specimen|Follitropin^4th specimen
C1978355|T201|COMP|50481-1|LNC|Follitropin^5th specimen|Follitropin^5th specimen
C1978356|T201|COMP|50482-9|LNC|Follitropin^6th specimen|Follitropin^6th specimen
C1978357|T201|COMP|50483-7|LNC|Follitropin^7th specimen|Follitropin^7th specimen
C1978358|T201|COMP|50484-5|LNC|Follitropin^8th specimen|Follitropin^8th specimen
C1978359|T201|COMP|50485-2|LNC|Gastrin^1st specimen|Gastrin^1st specimen
C1978360|T201|COMP|50486-0|LNC|Gastrin^2nd specimen|Gastrin^2nd specimen
C1978361|T201|COMP|50487-8|LNC|Gastrin^3rd specimen|Gastrin^3rd specimen
C1978362|T201|COMP|50488-6|LNC|Gastrin^4th specimen|Gastrin^4th specimen
C1978363|T201|COMP|50489-4|LNC|Gastrin^5th specimen|Gastrin^5th specimen
C1978364|T201|COMP|50490-2|LNC|Gastrin^6th specimen|Gastrin^6th specimen
C1978365|T201|COMP|50491-0|LNC|Gastrin^7th specimen|Gastrin^7th specimen
C1978366|T201|COMP|50492-8|LNC|Gastrin^8th specimen|Gastrin^8th specimen
C1978367|T201|COMP|50493-6|LNC|Somatotropin^1st specimen|Somatotropin^1st specimen
C1978368|T201|COMP|50494-4|LNC|Somatotropin^2nd specimen|Somatotropin^2nd specimen
C1978369|T201|COMP|50495-1|LNC|Somatotropin^3rd specimen|Somatotropin^3rd specimen
C1978370|T201|COMP|50496-9|LNC|Somatotropin^4th specimen|Somatotropin^4th specimen
C1978371|T201|COMP|50497-7|LNC|Somatotropin^5th specimen|Somatotropin^5th specimen
C1978372|T201|COMP|50498-5|LNC|Somatotropin^6th specimen|Somatotropin^6th specimen
C1978373|T201|COMP|50499-3|LNC|Somatotropin^7th specimen|Somatotropin^7th specimen
C1978374|T201|COMP|50500-8|LNC|Somatotropin^8th specimen|Somatotropin^8th specimen
C1978375|T201|COMP|50501-6|LNC|Insulin^1st specimen|Insulin^1st specimen
C1978376|T201|COMP|50502-4|LNC|Insulin^2nd specimen|Insulin^2nd specimen
C1978377|T201|COMP|50503-2|LNC|Insulin^3rd specimen|Insulin^3rd specimen
C1978378|T201|COMP|50504-0|LNC|Insulin^4th specimen|Insulin^4th specimen
C1978379|T201|COMP|50505-7|LNC|Insulin^5th specimen|Insulin^5th specimen
C1978380|T201|COMP|50506-5|LNC|Insulin^6th specimen|Insulin^6th specimen
C1978381|T201|COMP|50507-3|LNC|Insulin^7th specimen|Insulin^7th specimen
C1978382|T201|COMP|50508-1|LNC|Insulin^8th specimen|Insulin^8th specimen
C1978383|T201|COMP|50509-9|LNC|Lutropin^1st specimen|Lutropin^1st specimen
C1978384|T201|COMP|50510-7|LNC|Lutropin^2nd specimen|Lutropin^2nd specimen
C1978385|T201|COMP|50511-5|LNC|Lutropin^3rd specimen|Lutropin^3rd specimen
C1978386|T201|COMP|50512-3|LNC|Lutropin^4th specimen|Lutropin^4th specimen
C1978387|T201|COMP|50513-1|LNC|Lutropin^5th specimen|Lutropin^5th specimen
C1978388|T201|COMP|50514-9|LNC|Lutropin^6th specimen|Lutropin^6th specimen
C1978389|T201|COMP|50515-6|LNC|Lutropin^7th specimen|Lutropin^7th specimen
C1978390|T201|COMP|50516-4|LNC|Lutropin^8th specimen|Lutropin^8th specimen
C1978391|T201|COMP|50517-2|LNC|Prolactin^1st specimen|Prolactin^1st specimen
C1978392|T201|COMP|51110-5|LNC|Blasts.CD2/100 blasts|Blasts.CD2/100 blasts
C1978393|T201|COMP|51111-3|LNC|Blasts.CD2/100 blasts|Blasts.CD2/100 blasts
C1978394|T201|COMP|51112-1|LNC|Blasts.CD2|Blasts.CD2
C1978395|T201|COMP|51113-9|LNC|Blasts.CD2|Blasts.CD2
C1978396|T201|COMP|51114-7|LNC|Blasts.CD2|Blasts.CD2
C1978397|T201|COMP|51115-4|LNC|Blasts.CD20/100 blasts|Blasts.CD20/100 blasts
C1978398|T201|COMP|51116-2|LNC|Blasts.CD20/100 blasts|Blasts.CD20/100 blasts
C1978399|T201|COMP|51117-0|LNC|Blasts.CD21/100 blasts|Blasts.CD21/100 blasts
C1978401|T201|COMP|51118-8|LNC|Blasts.cytoplasmic CD22/100 blasts|Blasts.cytoplasmic CD22/100 blasts
C1978403|T201|COMP|51119-6|LNC|Blasts.cytoplasmic CD22/100 blasts|Blasts.cytoplasmic CD22/100 blasts
C1978404|T201|COMP|51120-4|LNC|Blasts.cytoplasmic CD22/100 blasts|Blasts.cytoplasmic CD22/100 blasts
C1978405|T201|COMP|51121-2|LNC|Blasts.cytoplasmic CD22|Blasts.cytoplasmic CD22
C1978407|T201|COMP|51122-0|LNC|Blasts.cytoplasmic CD22|Blasts.cytoplasmic CD22
C1978408|T201|COMP|51123-8|LNC|Blasts.cytoplasmic CD22|Blasts.cytoplasmic CD22
C1978409|T201|COMP|51124-6|LNC|Blasts.CD22/100 blasts|Blasts.CD22/100 blasts
C1978411|T201|COMP|51125-3|LNC|Blasts.CD22/100 blasts|Blasts.CD22/100 blasts
C1978412|T201|COMP|51126-1|LNC|Blasts.CD22/100 blasts|Blasts.CD22/100 blasts
C1978413|T201|COMP|51127-9|LNC|Blasts.CD22|Blasts.CD22
C1978415|T201|COMP|51128-7|LNC|Blasts.CD22|Blasts.CD22
C1978416|T201|COMP|51129-5|LNC|Blasts.CD22|Blasts.CD22
C1978417|T201|COMP|51130-3|LNC|Blasts.CD23/100 blasts|Blasts.CD23/100 blasts
C1978419|T201|COMP|51131-1|LNC|Blasts.CD23/100 blasts|Blasts.CD23/100 blasts
C1978420|T201|COMP|51132-9|LNC|Blasts.CD23/100 blasts|Blasts.CD23/100 blasts
C1978421|T201|COMP|51133-7|LNC|Blasts.CD24/100 blasts|Blasts.CD24/100 blasts
C1978423|T201|COMP|51134-5|LNC|Blasts.CD25/100 blasts|Blasts.CD25/100 blasts
C1978425|T201|COMP|51135-2|LNC|Blasts.CD25/100 blasts|Blasts.CD25/100 blasts
C1978426|T201|COMP|51136-0|LNC|Blasts.CD25/100 blasts|Blasts.CD25/100 blasts
C1978427|T201|COMP|51137-8|LNC|Blasts.cytoplasmic CD3/100 blasts|Blasts.cytoplasmic CD3/100 blasts
C1978429|T201|COMP|51138-6|LNC|Blasts.cytoplasmic CD3/100 blasts|Blasts.cytoplasmic CD3/100 blasts
C1978430|T201|COMP|51139-4|LNC|Blasts.cytoplasmic CD3/100 blasts|Blasts.cytoplasmic CD3/100 blasts
C1978431|T201|COMP|51140-2|LNC|Blasts.cytoplasmic CD3|Blasts.cytoplasmic CD3
C1978433|T201|COMP|51141-0|LNC|Blasts.cytoplasmic CD3|Blasts.cytoplasmic CD3
C1978434|T201|COMP|51385-3|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C1978435|T201|COMP|51386-1|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C1978450|T201|COMP|51396-0|LNC|Cells.CD65w/100 cells|Cells.CD65w/100 cells
C1978452|T201|COMP|51397-8|LNC|Cells.CD65w/100 cells|Cells.CD65w/100 cells
C1978453|T201|COMP|51398-6|LNC|Cells.CD65w/100 cells|Cells.CD65w/100 cells
C1978454|T201|COMP|51399-4|LNC|Cells.CD65w/100 cells|Cells.CD65w/100 cells
C1978455|T201|COMP|50531-3|LNC|Parathyrin.intact^7th specimen|Parathyrin.intact^7th specimen
C1978456|T201|COMP|50532-1|LNC|Parathyrin.intact^8th specimen|Parathyrin.intact^8th specimen
C1978457|T201|COMP|50533-9|LNC|Thyrotropin^1st specimen|Thyrotropin^1st specimen
C1978458|T201|COMP|50534-7|LNC|Thyrotropin^2nd specimen|Thyrotropin^2nd specimen
C1978459|T201|COMP|50535-4|LNC|Thyrotropin^3rd specimen|Thyrotropin^3rd specimen
C1978460|T201|COMP|50536-2|LNC|Thyrotropin^4th specimen|Thyrotropin^4th specimen
C1978461|T201|COMP|50537-0|LNC|Thyrotropin^5th specimen|Thyrotropin^5th specimen
C1978462|T201|COMP|50538-8|LNC|Thyrotropin^6th specimen|Thyrotropin^6th specimen
C1978463|T201|COMP|50539-6|LNC|Thyrotropin^7th specimen|Thyrotropin^7th specimen
C1978464|T201|COMP|50540-4|LNC|Thyrotropin^8th specimen|Thyrotropin^8th specimen
C1978465|T201|COMP|50541-2|LNC|Thyrotropin^20M post dose TRH|Thyrotropin^20M post dose TRH
C1978466|T201|COMP|50542-0|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C1978467|T201|COMP|50543-8|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C1978468|T201|COMP|50544-6|LNC|Everolimus|Everolimus
C1978469|T201|COMP|50545-3|LNC|Bacterial susceptibility panel|Bacterial susceptibility panel
C1978470|T201|COMP|50546-1|LNC|Bacterial susceptibility panel|Bacterial susceptibility panel
C1978471|T201|COMP|50547-9|LNC|Eastern equine encephalitis virus RNA|Eastern equine encephalitis virus RNA
C1978472|T201|COMP|50548-7|LNC|Respiratory virus DNA+RNA|Respiratory virus DNA+RNA
C1978474|T201|COMP|50549-5|LNC|Cytomegalovirus+Epstein Barr virus DNA|Cytomegalovirus+Epstein Barr virus DNA
C1978476|T201|COMP|50550-3|LNC|Malondialdehyde.free|Malondialdehyde.free
C1978478|T201|COMP|50551-1|LNC|Bilirubin|Bilirubin
C1978479|T201|COMP|50552-9|LNC|Clarity|Clarity
C1978480|T201|COMP|50553-7|LNC|Color|Color
C1978481|T201|COMP|50554-5|LNC|Urinalysis microscopic panel|Urinalysis microscopic panel
C1978482|T201|COMP|50555-2|LNC|Glucose|Glucose
C1978483|T201|COMP|50556-0|LNC|Urinalysis dipstick panel|Urinalysis dipstick panel
C1978484|T201|COMP|50557-8|LNC|Ketones|Ketones
C1978485|T201|COMP|50558-6|LNC|Nitrite|Nitrite
C1978486|T201|COMP|50559-4|LNC|Hemoglobin|Hemoglobin
C1978488|T201|COMP|50561-0|LNC|Protein|Protein
C1978489|T201|COMP|50562-8|LNC|Specific gravity|Specific gravity
C1978490|T201|COMP|50563-6|LNC|Urobilinogen|Urobilinogen
C1978491|T201|COMP|50564-4|LNC|Urinalysis panel|Urinalysis panel
C1978520|T201|COMP|50579-2|LNC|Gastric analysis panel|Gastric analysis panel
C1978524|T201|COMP|50581-8|LNC|Adenosine monophosphate.cyclic stimulation panel|Adenosine monophosphate.cyclic stimulation panel
C1978526|T201|COMP|50582-6|LNC|Glucose tolerance gestational panel|Glucose tolerance gestational panel
C1978528|T201|COMP|50583-4|LNC|Glucose screen gestational panel|Glucose screen gestational panel
C1978530|T201|COMP|50584-2|LNC|Lactose challenge panel|Lactose challenge panel
C1978532|T201|COMP|50585-9|LNC|Triple bolus stimulation panel|Triple bolus stimulation panel
C1978534|T201|COMP|50586-7|LNC|Glucose tolerance 3H panel|Glucose tolerance 3H panel
C1978536|T201|COMP|50587-5|LNC|Glucose tolerance 4H panel|Glucose tolerance 4H panel
C1978538|T201|COMP|50588-3|LNC|Glucose tolerance 5H panel|Glucose tolerance 5H panel
C1978540|T201|COMP|50589-1|LNC|Glucose tolerance 6H panel|Glucose tolerance 6H panel
C1978542|T201|COMP|50590-9|LNC|Adenine phosphoribosyltransferase|Adenine phosphoribosyltransferase
C1978543|T201|COMP|50591-7|LNC|Adenosine deaminase|Adenosine deaminase
C1978544|T201|COMP|50592-5|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C1978545|T201|COMP|50593-3|LNC|3-Hydroxybenzoylecgonine|3-Hydroxybenzoylecgonine
C1978546|T201|COMP|50594-1|LNC|3-Hydroxybenzoylecgonine|3-Hydroxybenzoylecgonine
C1978547|T201|COMP|50595-8|LNC|Pathologist interpretation|Pathologist interpretation
C1978548|T201|COMP|50596-6|LNC|HPA-1a|HPA-1a
C1978549|T201|COMP|50597-4|LNC|HPA-2|HPA-2
C1978551|T201|COMP|50598-2|LNC|HPA-15|HPA-15
C1978553|T201|COMP|50599-0|LNC|HPA-1|HPA-1
C1978554|T201|COMP|50600-6|LNC|HPA-3|HPA-3
C1978556|T201|COMP|50601-4|LNC|HPA-4|HPA-4
C1978558|T201|COMP|50602-2|LNC|HPA-5|HPA-5
C1978559|T201|COMP|50603-0|LNC|HPA-6|HPA-6
C1978561|T201|COMP|50604-8|LNC|HPA panel|HPA panel
C1978562|T201|COMP|50605-5|LNC|Hydrogen/Expired gas^pre XXX challenge|Hydrogen/Expired gas^pre XXX challenge
C1978563|T201|COMP|50606-3|LNC|Hydrogen/Expired gas^4H post XXX challenge|Hydrogen/Expired gas^4H post XXX challenge
C1978564|T201|COMP|50607-1|LNC|Neisseria meningitidis serogroups Ag panel|Neisseria meningitidis serogroups Ag panel
C1978566|T201|COMP|50608-9|LNC|Glucose tolerance 3H gestational panel|Glucose tolerance 3H gestational panel
C1978568|T201|COMP|50609-7|LNC|Nitroblue tetrazolium test|Nitroblue tetrazolium test
C1978570|T201|COMP|50611-3|LNC|Felbamate|Felbamate
C1978571|T201|COMP|50612-1|LNC|Chlamydophila pneumoniae Ab.IgA & IgG & IgM|Chlamydophila pneumoniae Ab.IgA & IgG & IgM
C1978573|T201|COMP|50613-9|LNC|Hydrogen/Expired gas^3.5H post XXX challenge|Hydrogen/Expired gas^3.5H post XXX challenge
C1978574|T201|COMP|50614-7|LNC|Hydrogen/Expired gas^4.5H post XXX challenge|Hydrogen/Expired gas^4.5H post XXX challenge
C1978575|T201|COMP|50615-4|LNC|Hydrogen/Expired gas^5H post XXX challenge|Hydrogen/Expired gas^5H post XXX challenge
C1978576|T201|COMP|50616-2|LNC|Hydrogen/Expired gas^5.5H post XXX challenge|Hydrogen/Expired gas^5.5H post XXX challenge
C1978577|T201|COMP|50617-0|LNC|Hydrogen/Expired gas^6H post XXX challenge|Hydrogen/Expired gas^6H post XXX challenge
C1978578|T201|COMP|50618-8|LNC|Phosphatidylcholine.saturated/Surfactant.total|Phosphatidylcholine.saturated/Surfactant.total
C1978580|T201|COMP|50619-6|LNC|Karyotype|Karyotype
C1978581|T201|COMP|50620-4|LNC|Opiates cutoff|Opiates cutoff
C1978582|T201|COMP|50621-2|LNC|HTT gene targeted mutation analysis|HTT gene targeted mutation analysis
C1978583|T201|COMP|50622-0|LNC|Allergen.miscellaneous Ab.IgG|Allergen.miscellaneous Ab.IgG
C1978585|T201|COMP|50623-8|LNC|AS gene targeted mutation analysis|AS gene targeted mutation analysis
C1978586|T201|COMP|50624-6|LNC|HIV 1 RNA panel|HIV 1 RNA panel
C1978588|T201|COMP|50625-3|LNC|Ova & parasites identified|Ova & parasites identified
C1978589|T201|COMP|50626-1|LNC|DMD gene targeted mutation analysis|DMD gene targeted mutation analysis
C1978590|T201|COMP|50627-9|LNC|Immunoglobulin heavy chain gene rearrangements|Immunoglobulin heavy chain gene rearrangements
C1978591|T201|COMP|50628-7|LNC|Heptacarboxylporphyrin/Creatinine|Heptacarboxylporphyrin/Creatinine
C1978592|T201|COMP|50629-5|LNC|Liver kidney microsomal Ab.IgG|Liver kidney microsomal Ab.IgG
C1978593|T201|COMP|50630-3|LNC|Gentamicin|Gentamicin
C1978594|T201|COMP|50631-1|LNC|Cefepime|Cefepime
C1978595|T201|COMP|50632-9|LNC|Cefotaxime|Cefotaxime
C1978596|T201|COMP|50633-7|LNC|cefTRIAXone|cefTRIAXone
C1978597|T201|COMP|50634-5|LNC|Populus balsamifera Ab.IgE|Populus balsamifera Ab.IgE
C1978599|T201|COMP|50635-2|LNC|Cupressus macrocarpa Ab.IgE|Cupressus macrocarpa Ab.IgE
C1978601|T201|COMP|50636-0|LNC|Macrocheira kaempferi Ab.IgE|Macrocheira kaempferi Ab.IgE
C1978603|T201|COMP|50637-8|LNC|Coagulation factor XIII inhibitor|Coagulation factor XIII inhibitor
C1978604|T201|COMP|50638-6|LNC|Bixa orellana seed Ab.IgE|Bixa orellana seed Ab.IgE
C1978606|T201|COMP|50639-4|LNC|Harmonia axyridis Ab.IgE|Harmonia axyridis Ab.IgE
C1978608|T201|COMP|50640-2|LNC|Cells.CD3+CD57+|Cells.CD3+CD57+
C1978610|T201|COMP|50641-0|LNC|Cells.CD3+CD8+CD57+|Cells.CD3+CD8+CD57+
C1978612|T201|COMP|50642-8|LNC|Human papilloma virus 6+11+42+43+44 DNA|Human papilloma virus 6+11+42+43+44 DNA
C1978613|T201|COMP|50643-6|LNC|Pregnanetriolone|Pregnanetriolone
C1978614|T201|COMP|50644-4|LNC|Tetrahydrocorticosterone/Creatinine|Tetrahydrocorticosterone/Creatinine
C1978616|T201|COMP|50645-1|LNC|Tetrahydrocortisol/Creatinine|Tetrahydrocortisol/Creatinine
C1978618|T201|COMP|50646-9|LNC|Latex recombinant (rHev b) 1 Ab.IgE|Latex recombinant (rHev b) 1 Ab.IgE
C1978620|T201|COMP|50647-7|LNC|Latex recombinant (rHev b) 11 Ab.IgE|Latex recombinant (rHev b) 11 Ab.IgE
C1978622|T201|COMP|50648-5|LNC|Latex recombinant (rHev b) 6.01 Ab.IgE|Latex recombinant (rHev b) 6.01 Ab.IgE
C1978624|T201|COMP|50649-3|LNC|Latex recombinant (rHev b) 6.02 Ab.IgE|Latex recombinant (rHev b) 6.02 Ab.IgE
C1978626|T201|COMP|50650-1|LNC|Lupinus albus seed Ab.IgE|Lupinus albus seed Ab.IgE
C1978635|T201|COMP|50658-4|LNC|Basophils.band form/100 leukocytes|Basophils.band form/100 leukocytes
C1978637|T201|COMP|50659-2|LNC|Chromosome analysis.interphase|Chromosome analysis.interphase
C1978639|T201|COMP|50660-0|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C1978640|T201|COMP|50661-8|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C1978641|T201|COMP|50662-6|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C1978642|T201|COMP|50663-4|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C1978643|T201|COMP|50664-2|LNC|Cells.CD19+Kappa+|Cells.CD19+Kappa+
C1978644|T201|COMP|50665-9|LNC|Cells.CD19+Lambda+|Cells.CD19+Lambda+
C1978645|T201|COMP|50666-7|LNC|Nuclear matrix protein 22|Nuclear matrix protein 22
C1978646|T201|COMP|50667-5|LNC|Glucose tolerance|Glucose tolerance
C1978648|T201|COMP|50669-1|LNC|Transfuse antithrombin|Transfuse antithrombin
C1978650|T201|COMP|50670-9|LNC|Erythrocyte agglutination|Erythrocyte agglutination
C1978651|T201|COMP|50671-7|LNC|Corticotropin releasing hormone|Corticotropin releasing hormone
C1978652|T201|COMP|50672-5|LNC|Leukocyte toxic vacuoles|Leukocyte toxic vacuoles
C1978654|T201|COMP|50673-3|LNC|Insulin XXX challenge panel|Insulin XXX challenge panel
C1978656|T201|COMP|50674-1|LNC|Spherocytes|Spherocytes
C1978657|T201|COMP|50675-8|LNC|Calcium-phosphorus product|Calcium-phosphorus product
C1978658|T201|COMP|50676-6|LNC|Calcium-phosphorus product panel|Calcium-phosphorus product panel
C1978660|T201|COMP|50677-4|LNC|Semen analysis post vasectomy panel|Semen analysis post vasectomy panel
C1978662|T201|COMP|50678-2|LNC|Spondylocladium sp Ab.IgE.Rast Class|Spondylocladium sp Ab.IgE.Rast Class
C1978665|T201|COMP|50680-8|LNC|Paecilomyces variottii Ab.IgE|Paecilomyces variottii Ab.IgE
C1978667|T201|COMP|50681-6|LNC|Thyroxine binding protein pattern|Thyroxine binding protein pattern
C1978669|T201|COMP|50682-4|LNC|PRKCG gene.CAG repeats|PRKCG gene.CAG repeats
C1978673|T201|COMP|50684-0|LNC|Chromosome analysis.interphase|Chromosome analysis.interphase
C1978674|T201|COMP|50685-7|LNC|Somatotropin|Somatotropin
C1978675|T201|COMP|50686-5|LNC|11-Dehydro thromboxane beta 2/Creatinine|11-Dehydro thromboxane beta 2/Creatinine
C1978677|T201|COMP|50687-3|LNC|Plasmodium sp Ag|Plasmodium sp Ag
C1978678|T201|COMP|50688-1|LNC|Plasmodium sp lactate dehydrogenase|Plasmodium sp lactate dehydrogenase
C1978680|T201|COMP|50689-9|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1978681|T201|COMP|50690-7|LNC|Reagin Ab|Reagin Ab
C1978682|T201|COMP|50691-5|LNC|Coxsackievirus A9+B1+B2+B3+B4+B5+B6 Ab|Coxsackievirus A9+B1+B2+B3+B4+B5+B6 Ab
C1978684|T201|COMP|50692-3|LNC|Parainfluenza virus 1+2+3 Ab|Parainfluenza virus 1+2+3 Ab
C1978685|T201|COMP|50693-1|LNC|Influenza virus A+B Ab|Influenza virus A+B Ab
C1978688|T201|COMP|50704-6|LNC|Influenza virus A nucleoprotein RNA|Influenza virus A nucleoprotein RNA
C1978690|T201|COMP|50705-3|LNC|Influenza virus A non-structural protein RNA|Influenza virus A non-structural protein RNA
C1978692|T201|COMP|50706-1|LNC|Influenza virus A polymerase A RNA|Influenza virus A polymerase A RNA
C1978694|T201|COMP|50707-9|LNC|Influenza virus A polymerase B1 cDNA|Influenza virus A polymerase B1 cDNA
C1978696|T201|COMP|50708-7|LNC|Influenza virus A polymerase B2 RNA|Influenza virus A polymerase B2 RNA
C1978698|T201|COMP|50709-5|LNC|Influenza virus B Ab|Influenza virus B Ab
C1978699|T201|COMP|50710-3|LNC|Influenza virus susceptibility panel|Influenza virus susceptibility panel
C1978701|T201|COMP|50711-1|LNC|Influenza virus A polymerase RNA|Influenza virus A polymerase RNA
C1978707|T201|COMP|50714-5|LNC|Rumex obtusifolius Ab.IgE|Rumex obtusifolius Ab.IgE
C1978711|T201|COMP|50716-0|LNC|11-Deoxycortisol^7th specimen post XXX challenge|11-Deoxycortisol^7th specimen post XXX challenge
C1978712|T201|COMP|50717-8|LNC|11-Deoxycortisol^6th specimen post XXX challenge|11-Deoxycortisol^6th specimen post XXX challenge
C1978713|T201|COMP|50718-6|LNC|11-Deoxycortisol^5th specimen post XXX challenge|11-Deoxycortisol^5th specimen post XXX challenge
C1978714|T201|COMP|50719-4|LNC|11-Deoxycortisol^4th specimen post XXX challenge|11-Deoxycortisol^4th specimen post XXX challenge
C1978715|T201|COMP|50720-2|LNC|11-Deoxycortisol^3rd specimen post XXX challenge|11-Deoxycortisol^3rd specimen post XXX challenge
C1978716|T201|COMP|50721-0|LNC|11-Deoxycortisol^1st specimen post XXX challenge|11-Deoxycortisol^1st specimen post XXX challenge
C1978717|T201|COMP|50722-8|LNC|VKORC1 gene targeted mutation analysis|VKORC1 gene targeted mutation analysis
C1978719|T201|COMP|50723-6|LNC|Cells.CD38+Lambda+|Cells.CD38+Lambda+
C1978720|T201|COMP|50724-4|LNC|Lymphoblasts/100 leukocytes|Lymphoblasts/100 leukocytes
C1978721|T201|COMP|50725-1|LNC|Monoblasts/100 leukocytes|Monoblasts/100 leukocytes
C1978722|T201|COMP|50726-9|LNC|Reticulum cell/100 cells|Reticulum cell/100 cells
C1978728|T201|COMP|50729-3|LNC|Serotonin release 100 U/mL heparin.porcine|Serotonin release 100 U/mL heparin.porcine
C1978730|T201|COMP|50730-1|LNC|Serotonin release 0.1 U/mL heparin.porcine|Serotonin release 0.1 U/mL heparin.porcine
C1978736|T201|COMP|50733-5|LNC|Serotonin release interpretation|Serotonin release interpretation
C1978748|T201|COMP|50746-7|LNC|Hirudin|Hirudin
C1978749|T201|COMP|50747-5|LNC|Platelet factor 4 Ag|Platelet factor 4 Ag
C1978750|T201|COMP|50748-3|LNC|Alpha-2-Macroglobulin/Creatinine|Alpha-2-Macroglobulin/Creatinine
C1978752|T201|COMP|50749-1|LNC|Protein|Protein
C1978753|T201|COMP|50750-9|LNC|F13A1 gene.p.Val34Leu|F13A1 gene.p.Val34Leu
C1978755|T201|COMP|50751-7|LNC|Glucose^15M post 0.1 U/kg insulin|Glucose^15M post 0.1 U/kg insulin
C1978756|T201|COMP|50752-5|LNC|Cortisol^15M post dose insulin IV|Cortisol^15M post dose insulin IV
C1978757|T201|COMP|50753-3|LNC|Somatotropin^15M post dose insulin IV|Somatotropin^15M post dose insulin IV
C1978758|T201|COMP|50754-1|LNC|Coagulation surface induced|Coagulation surface induced
C1978760|T201|COMP|50756-6|LNC|Creatine kinase|Creatine kinase
C1978761|T201|COMP|50757-4|LNC|Creatine kinase.total/Creatine kinase.MB|Creatine kinase.total/Creatine kinase.MB
C1978762|T201|COMP|50758-2|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C1978763|T201|COMP|50759-0|LNC|Beta-N-acetylhexosaminidase.A|Beta-N-acetylhexosaminidase.A
C1978765|T201|COMP|50761-6|LNC|A Ab.IgG|A Ab.IgG
C1978767|T201|COMP|50762-4|LNC|A Ab.IgM|A Ab.IgM
C1978769|T201|COMP|50763-2|LNC|B Ab.IgM|B Ab.IgM
C1978771|T201|COMP|50764-0|LNC|B Ab.IgG|B Ab.IgG
C1978773|T201|COMP|50765-7|LNC|Hemoglobin Hasharon/Hemoglobin.total|Hemoglobin Hasharon/Hemoglobin.total
C1978775|T201|COMP|50766-5|LNC|Fungus identified ^^^8|Fungus identified ^^^8
C1978776|T201|COMP|50767-3|LNC|Ganglioside GD1a Ab.IgG/Ganglioside GD1a Ab.IgM|Ganglioside GD1a Ab.IgG/Ganglioside GD1a Ab.IgM
C1978778|T201|COMP|50768-1|LNC|Ganglioside GD1b Ab.IgG/Ganglioside GD1b Ab.IgM|Ganglioside GD1b Ab.IgG/Ganglioside GD1b Ab.IgM
C1978782|T201|COMP|50770-7|LNC|Ganglioside GM1 Ab.IgG/Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgG/Ganglioside GM1 Ab.IgM
C1978784|T201|COMP|50771-5|LNC|Ganglioside GM2 Ab.IgG/Ganglioside GM2 Ab.IgM|Ganglioside GM2 Ab.IgG/Ganglioside GM2 Ab.IgM
C1978786|T201|COMP|50772-3|LNC|Ganglioside GQ1b Ab.IgG/Ganglioside GQ1b Ab.IgM|Ganglioside GQ1b Ab.IgG/Ganglioside GQ1b Ab.IgM
C1978788|T201|COMP|50773-1|LNC|ABO & Rh group^post transfusion reaction|ABO & Rh group^post transfusion reaction
C1978789|T201|COMP|50774-9|LNC|Nucleated cells|Nucleated cells
C1978790|T201|COMP|50783-0|LNC|Cells.CD15 actual/normal|Cells.CD15 actual/normal
C1978792|T201|COMP|50784-8|LNC|Cells.CD16 actual/normal|Cells.CD16 actual/normal
C1978794|T201|COMP|50785-5|LNC|Cells.CD18 actual/normal|Cells.CD18 actual/normal
C1978799|T201|COMP|50788-9|LNC|Cytokeratin cells/100 cells|Cytokeratin cells/100 cells
C1978801|T201|COMP|50789-7|LNC|Cytokeratin cells|Cytokeratin cells
C1978803|T201|COMP|50790-5|LNC|HIV 1 RNA tropism|HIV 1 RNA tropism
C1978805|T201|COMP|50791-3|LNC|Hemoglobin pattern|Hemoglobin pattern
C1978806|T201|COMP|50963-8|LNC|XXX blood group Ab.IgM|XXX blood group Ab.IgM
C1978808|T201|COMP|50964-6|LNC|Liley Zone|Liley Zone
C1978810|T201|COMP|50965-3|LNC|Gamma hydroxybutyrate cutoff|Gamma hydroxybutyrate cutoff
C1978812|T201|COMP|50966-1|LNC|Flunitrazepam|Flunitrazepam
C1978813|T201|COMP|50967-9|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C1978814|T201|COMP|50968-7|LNC|HLA Ab|HLA Ab
C1978815|T201|COMP|50969-5|LNC|Epstein Barr virus early diffuse Ab.IgG|Epstein Barr virus early diffuse Ab.IgG
C1978817|T201|COMP|50970-3|LNC|XXX blood group Ab|XXX blood group Ab
C1978819|T201|COMP|51461-2|LNC|Listeria sp Ab|Listeria sp Ab
C1978820|T201|COMP|51462-0|LNC|Onchocerca sp Ab.IgG2|Onchocerca sp Ab.IgG2
C1978821|T201|COMP|51463-8|LNC|Onchocerca sp Ab.IgG3|Onchocerca sp Ab.IgG3
C1978822|T201|COMP|51464-6|LNC|Onchocerca sp Ab.IgG4|Onchocerca sp Ab.IgG4
C1978823|T201|COMP|51465-3|LNC|Paragonimus sp Ab|Paragonimus sp Ab
C1978824|T201|COMP|51466-1|LNC|Parainfluenza virus 1+2+3 Ab|Parainfluenza virus 1+2+3 Ab
C1978825|T201|COMP|51467-9|LNC|Plasmodium falciparum Ab.IgG|Plasmodium falciparum Ab.IgG
C1978826|T201|COMP|51468-7|LNC|Plasmodium ovale Ab.IgG|Plasmodium ovale Ab.IgG
C1978827|T201|COMP|50792-1|LNC|Protein.monoclonal band 3/Protein.total|Protein.monoclonal band 3/Protein.total
C1978829|T201|COMP|50793-9|LNC|Protein.monoclonal band 4/Protein.total|Protein.monoclonal band 4/Protein.total
C1978831|T201|COMP|50794-7|LNC|Osmotic fragility.beginning hemolysis|Osmotic fragility.beginning hemolysis
C1978833|T201|COMP|50795-4|LNC|Osmotic fragility.full hemolysis|Osmotic fragility.full hemolysis
C1978835|T201|COMP|50796-2|LNC|Protein.monoclonal band 3|Protein.monoclonal band 3
C1978837|T201|COMP|50797-0|LNC|Protein.monoclonal band 4|Protein.monoclonal band 4
C1978839|T201|COMP|50798-8|LNC|17-Ketogenic steroids|17-Ketogenic steroids
C1978840|T201|COMP|50799-6|LNC|7-Dehydrocholesterol|7-Dehydrocholesterol
C1978841|T201|COMP|50800-2|LNC|Acetone|Acetone
C1978842|T201|COMP|50801-0|LNC|Aluminum|Aluminum
C1978843|T201|COMP|50802-8|LNC|Amikacin^peak|Amikacin^peak
C1978844|T201|COMP|50803-6|LNC|Amikacin^trough|Amikacin^trough
C1978845|T201|COMP|50804-4|LNC|Amitriptyline|Amitriptyline
C1978846|T201|COMP|50805-1|LNC|Amitriptyline|Amitriptyline
C1978847|T201|COMP|50806-9|LNC|Antimony|Antimony
C1978848|T201|COMP|50807-7|LNC|Antimony|Antimony
C1978849|T201|COMP|50808-5|LNC|Antimony|Antimony
C1978850|T201|COMP|50809-3|LNC|Antimony|Antimony
C1978851|T201|COMP|50810-1|LNC|Antimony|Antimony
C1978852|T201|COMP|50811-9|LNC|Antimony|Antimony
C1978853|T201|COMP|50812-7|LNC|Arsenic|Arsenic
C1978854|T201|COMP|50813-5|LNC|Arsenic|Arsenic
C1978855|T201|COMP|50814-3|LNC|Arsenic.inorganic|Arsenic.inorganic
C1978856|T201|COMP|50815-0|LNC|Arsenic.inorganic|Arsenic.inorganic
C1978857|T201|COMP|50816-8|LNC|Arsenic.organic|Arsenic.organic
C1978858|T201|COMP|50817-6|LNC|Arsenic/Creatinine|Arsenic/Creatinine
C1978859|T201|COMP|50818-4|LNC|Barium|Barium
C1978860|T201|COMP|50819-2|LNC|Barium|Barium
C1978861|T201|COMP|50820-0|LNC|Base excess|Base excess
C1978862|T201|COMP|50821-8|LNC|Beryllium|Beryllium
C1978863|T201|COMP|50822-6|LNC|Beryllium|Beryllium
C1978864|T201|COMP|50823-4|LNC|Beryllium|Beryllium
C1978865|T201|COMP|50824-2|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C1978866|T201|COMP|50825-9|LNC|Bile acid|Bile acid
C1978867|T201|COMP|50826-7|LNC|Bismuth|Bismuth
C1978868|T201|COMP|50827-5|LNC|Boron|Boron
C1978869|T201|COMP|50828-3|LNC|Boron|Boron
C1978870|T201|COMP|50829-1|LNC|Boron|Boron
C1978871|T201|COMP|50830-9|LNC|Boron|Boron
C1978872|T201|COMP|50831-7|LNC|Boron/Creatinine|Boron/Creatinine
C1978873|T201|COMP|50832-5|LNC|Boron/Creatinine|Boron/Creatinine
C1978874|T201|COMP|50833-3|LNC|Cadmium|Cadmium
C1978875|T201|COMP|50834-1|LNC|Cadmium|Cadmium
C1978876|T201|COMP|50835-8|LNC|Cadmium/Creatinine|Cadmium/Creatinine
C1978877|T201|COMP|50836-6|LNC|Calcium|Calcium
C1978878|T201|COMP|50837-4|LNC|Calcium.ionized|Calcium.ionized
C1978879|T201|COMP|50838-2|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C1978880|T201|COMP|50839-0|LNC|Calcium/Creatinine|Calcium/Creatinine
C1978881|T201|COMP|50840-8|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C1978882|T201|COMP|50841-6|LNC|Chromium|Chromium
C1978883|T201|COMP|50842-4|LNC|Chromium|Chromium
C1978884|T201|COMP|50843-2|LNC|clonazePAM|clonazePAM
C1978885|T201|COMP|50844-0|LNC|cloZAPine|cloZAPine
C1978886|T201|COMP|50845-7|LNC|Cobalt|Cobalt
C1978887|T201|COMP|50846-5|LNC|Cobalt|Cobalt
C1978888|T201|COMP|50847-3|LNC|Cobalt|Cobalt
C1978889|T201|COMP|50848-1|LNC|Cortisol|Cortisol
C1978890|T201|COMP|50849-9|LNC|Diazepam+Nordiazepam|Diazepam+Nordiazepam
C1978891|T201|COMP|50850-7|LNC|Fluoride/Creatinine|Fluoride/Creatinine
C1978892|T201|COMP|50851-5|LNC|Germanium|Germanium
C1978893|T201|COMP|50852-3|LNC|Gold|Gold
C1978894|T201|COMP|50853-1|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C1978895|T201|COMP|50854-9|LNC|Heptaporphyrin|Heptaporphyrin
C1978896|T201|COMP|50855-6|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C1978897|T201|COMP|50856-4|LNC|Hexaporphyrin|Hexaporphyrin
C1978898|T201|COMP|50857-2|LNC|Histamine|Histamine
C1978899|T201|COMP|50858-0|LNC|Hydrogen ion|Hydrogen ion
C1978900|T201|COMP|50859-8|LNC|Hydrogen ion|Hydrogen ion
C1978901|T201|COMP|50860-6|LNC|Hydrogen ion|Hydrogen ion
C1978902|T201|COMP|50861-4|LNC|Hydrogen ion|Hydrogen ion
C1978903|T201|COMP|50862-2|LNC|Hydrogen ion|Hydrogen ion
C1978904|T201|COMP|50863-0|LNC|Hydrogen ion|Hydrogen ion
C1978905|T201|COMP|50864-8|LNC|Hydrogen ion|Hydrogen ion
C1978906|T201|COMP|50865-5|LNC|Hydrogen ion|Hydrogen ion
C1978907|T201|COMP|50866-3|LNC|Indicans/Creatinine|Indicans/Creatinine
C1978908|T201|COMP|50867-1|LNC|Insulin|Insulin
C1978909|T201|COMP|50868-9|LNC|Iodine|Iodine
C1978910|T201|COMP|50869-7|LNC|Iron|Iron
C1978911|T201|COMP|50870-5|LNC|Isopropanol|Isopropanol
C1978912|T201|COMP|50871-3|LNC|Lead|Lead
C1978913|T201|COMP|50872-1|LNC|Lithium|Lithium
C1978914|T201|COMP|50873-9|LNC|Magnesium/Creatinine|Magnesium/Creatinine
C1978915|T201|COMP|50874-7|LNC|Manganese|Manganese
C1978916|T201|COMP|50875-4|LNC|Manganese|Manganese
C1978917|T201|COMP|50876-2|LNC|Mercury|Mercury
C1978918|T201|COMP|50877-0|LNC|Mercury|Mercury
C1978919|T201|COMP|50878-8|LNC|Mercury|Mercury
C1978920|T201|COMP|50879-6|LNC|Methyl ethyl ketone|Methyl ethyl ketone
C1978921|T201|COMP|50880-4|LNC|Methyl ethyl ketone|Methyl ethyl ketone
C1978922|T201|COMP|50881-2|LNC|Molybdenum|Molybdenum
C1978923|T201|COMP|50882-0|LNC|Molybdenum|Molybdenum
C1978924|T201|COMP|50883-8|LNC|Molybdenum|Molybdenum
C1978925|T201|COMP|50884-6|LNC|Molybdenum|Molybdenum
C1978926|T201|COMP|50885-3|LNC|Naproxen|Naproxen
C1978927|T201|COMP|50886-1|LNC|Nickel|Nickel
C1978928|T201|COMP|50887-9|LNC|Nickel|Nickel
C1978929|T201|COMP|50888-7|LNC|Nitrogen|Nitrogen
C1978930|T201|COMP|50889-5|LNC|Nitrogen|Nitrogen
C1978931|T201|COMP|50890-3|LNC|Norclozapine|Norclozapine
C1978932|T201|COMP|50891-1|LNC|OLANZapine|OLANZapine
C1978933|T201|COMP|50892-9|LNC|Palladium|Palladium
C1978934|T201|COMP|50893-7|LNC|Paraquat|Paraquat
C1978935|T201|COMP|50894-5|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C1978939|T201|COMP|50898-6|LNC|Phosphate|Phosphate
C1978940|T201|COMP|50899-4|LNC|Platinum|Platinum
C1978941|T201|COMP|50900-0|LNC|Platinum|Platinum
C1978942|T201|COMP|50901-8|LNC|Porphyrins|Porphyrins
C1978943|T201|COMP|50902-6|LNC|Potassium|Potassium
C1978944|T201|COMP|50912-5|LNC|Sodium|Sodium
C1978945|T201|COMP|50913-3|LNC|Strontium|Strontium
C1978946|T201|COMP|50914-1|LNC|Strontium|Strontium
C1978947|T201|COMP|50915-8|LNC|Strontium|Strontium
C1978948|T201|COMP|50916-6|LNC|Sucrose|Sucrose
C1978949|T201|COMP|50917-4|LNC|Thallium|Thallium
C1978950|T201|COMP|50918-2|LNC|Thallium|Thallium
C1978951|T201|COMP|50919-0|LNC|Thorium|Thorium
C1978952|T201|COMP|50920-8|LNC|Thorium|Thorium
C1978953|T201|COMP|50921-6|LNC|Tin|Tin
C1978954|T201|COMP|50922-4|LNC|Tin|Tin
C1978955|T201|COMP|50923-2|LNC|Tin|Tin
C1978956|T201|COMP|50924-0|LNC|Titanium|Titanium
C1978957|T201|COMP|50925-7|LNC|Titanium|Titanium
C1978958|T201|COMP|50926-5|LNC|Titanium|Titanium
C1978959|T201|COMP|50927-3|LNC|Tobramycin|Tobramycin
C1978960|T201|COMP|50928-1|LNC|Uranium|Uranium
C1978961|T201|COMP|50929-9|LNC|Uranium|Uranium
C1978962|T201|COMP|50930-7|LNC|Uranium|Uranium
C1978963|T201|COMP|50931-5|LNC|Uroporphyrin 1 isomer|Uroporphyrin 1 isomer
C1978964|T201|COMP|50932-3|LNC|Uroporphyrin/Porphyrins.total|Uroporphyrin/Porphyrins.total
C1978965|T201|COMP|50933-1|LNC|Vanadium|Vanadium
C1978966|T201|COMP|50934-9|LNC|Vanadium|Vanadium
C1978967|T201|COMP|50935-6|LNC|Vanadium|Vanadium
C1978968|T201|COMP|50936-4|LNC|Vanadium|Vanadium
C1978969|T201|COMP|50937-2|LNC|Vanadium|Vanadium
C1978970|T201|COMP|50938-0|LNC|Vancomycin|Vancomycin
C1978971|T201|COMP|50939-8|LNC|Zinc|Zinc
C1978972|T201|COMP|50940-6|LNC|Zinc/Creatinine|Zinc/Creatinine
C1978973|T201|COMP|50941-4|LNC|Mycobacterium sp|Mycobacterium sp
C1978974|T201|COMP|50942-2|LNC|Acarboxyprothrombin|Acarboxyprothrombin
C1978980|T201|COMP|50947-1|LNC|Platelet aggregation.collagen induced^190 ug/mL|Platelet aggregation.collagen induced^190 ug/mL
C1978981|T201|COMP|50948-9|LNC|Vanillylmandelate & Creatinine|Vanillylmandelate & Creatinine
C1978983|T201|COMP|50949-7|LNC|Albumin|Albumin
C1978984|T201|COMP|50950-5|LNC|Phosphoethanolamine Ab.IgA|Phosphoethanolamine Ab.IgA
C1978986|T201|COMP|50951-3|LNC|Phosphoserine Ab.IgA|Phosphoserine Ab.IgA
C1978988|T201|COMP|50952-1|LNC|Phosphoserine Ab.IgG|Phosphoserine Ab.IgG
C1978990|T201|COMP|50953-9|LNC|Phosphoethanolamine Ab.IgM|Phosphoethanolamine Ab.IgM
C1978992|T201|COMP|50954-7|LNC|Phosphoethanolamine Ab.IgG|Phosphoethanolamine Ab.IgG
C1978994|T201|COMP|50955-4|LNC|Phosphoserine Ab.IgM|Phosphoserine Ab.IgM
C1978996|T201|COMP|50956-2|LNC|HLA-B*57:01|HLA-B*57:01
C1978997|T201|COMP|50957-0|LNC|Manual differential performed|Manual differential performed
C1979001|T201|COMP|50959-6|LNC|Indirect antiglobulin test.XXX reagent|Indirect antiglobulin test.XXX reagent
C1979002|T201|COMP|50960-4|LNC|Rabbit Ab|Rabbit Ab
C1979004|T201|COMP|50961-2|LNC|Rabbit Ab|Rabbit Ab
C1979005|T201|COMP|50962-0|LNC|XXX blood group Ab.IgG|XXX blood group Ab.IgG
C1979007|T201|COMP|50971-1|LNC|Cytology report|Cytology report
C1979008|T201|COMP|50972-9|LNC|Cells.CD138|Cells.CD138
C1979009|T201|COMP|50973-7|LNC|Cells.CD38+CD138+|Cells.CD38+CD138+
C1979011|T201|COMP|50974-5|LNC|Cells.CD38+CD138+/100 cells|Cells.CD38+CD138+/100 cells
C1979013|T201|COMP|50975-2|LNC|Cells.TCR alpha beta|Cells.TCR alpha beta
C1979014|T201|COMP|50976-0|LNC|Cells.TCR gamma delta|Cells.TCR gamma delta
C1979015|T201|COMP|50977-8|LNC|Echovirus 5 Ab|Echovirus 5 Ab
C1979017|T201|COMP|50978-6|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C1979018|T201|COMP|50979-4|LNC|CBir1 Ab|CBir1 Ab
C1979020|T201|COMP|50980-2|LNC|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1979022|T201|COMP|50982-8|LNC|Horowitz index|Horowitz index
C1979024|T201|COMP|50983-6|LNC|Horowitz index|Horowitz index
C1979025|T201|COMP|50984-4|LNC|Horowitz index|Horowitz index
C1979026|T201|COMP|50985-1|LNC|Horowitz index|Horowitz index
C1979027|T201|COMP|50986-9|LNC|Horowitz index|Horowitz index
C1979029|T201|COMP|50995-0|LNC|BRCA1+BRCA2 gene targeted mutation analysis|BRCA1+BRCA2 gene targeted mutation analysis
C1979031|T201|COMP|50996-8|LNC|HBB gene targeted mutation analysis|HBB gene targeted mutation analysis
C1979032|T201|COMP|50997-6|LNC|Complement C8.functional|Complement C8.functional
C1979034|T201|COMP|50998-4|LNC|CFTR gene mutations tested for|CFTR gene mutations tested for
C1979035|T201|COMP|50999-2|LNC|Leishmania donovani Ab.IgG & IgM|Leishmania donovani Ab.IgG & IgM
C1979037|T201|COMP|51000-8|LNC|Leishmania tropica Ab.IgG & IgM|Leishmania tropica Ab.IgG & IgM
C1979039|T201|COMP|51001-6|LNC|Iodide|Iodide
C1979040|T201|COMP|51002-4|LNC|Lipoprotein midband A|Lipoprotein midband A
C1979042|T201|COMP|51003-2|LNC|Lipoprotein midband B|Lipoprotein midband B
C1979044|T201|COMP|51004-0|LNC|Lipoprotein midband C|Lipoprotein midband C
C1979046|T201|COMP|51005-7|LNC|Testosterone.free+weakly bound|Testosterone.free+weakly bound
C1979047|T201|COMP|51006-5|LNC|Direct antiglobulin test.XXX reagent|Direct antiglobulin test.XXX reagent
C1979050|T201|COMP|51008-1|LNC|Triticum aestivum native (nTri a) 19 Ab.IgE|Triticum aestivum native (nTri a) 19 Ab.IgE
C1979052|T201|COMP|51009-9|LNC|Cells.CD3-CD16+CD56+CD244+/100 cells|Cells.CD3-CD16+CD56+CD244+/100 cells
C1979054|T201|COMP|51010-7|LNC|Cells.CD3-CD16+CD56+CD244+/100 cells|Cells.CD3-CD16+CD56+CD244+/100 cells
C1979055|T201|COMP|51011-5|LNC|Cells.CD3-CD16+CD56+CD244+/100 cells|Cells.CD3-CD16+CD56+CD244+/100 cells
C1979056|T201|COMP|51012-3|LNC|Cells.BCLXL/100 cells|Cells.BCLXL/100 cells
C1979058|T201|COMP|51013-1|LNC|Blasts.CD1/100 blasts|Blasts.CD1/100 blasts
C1979060|T201|COMP|51014-9|LNC|Blasts.CD1/100 blasts|Blasts.CD1/100 blasts
C1979061|T201|COMP|51015-6|LNC|Blasts.CD1/100 blasts|Blasts.CD1/100 blasts
C1979062|T201|COMP|51016-4|LNC|Blasts.CD1|Blasts.CD1
C1979064|T201|COMP|51017-2|LNC|Blasts.CD1|Blasts.CD1
C1979065|T201|COMP|51018-0|LNC|Blasts.CD10/100 blasts|Blasts.CD10/100 blasts
C1979066|T201|COMP|51019-8|LNC|Blasts.CD10/100 blasts|Blasts.CD10/100 blasts
C1979067|T201|COMP|51020-6|LNC|Blasts.CD10|Blasts.CD10
C1979068|T201|COMP|51021-4|LNC|Blasts.CD10|Blasts.CD10
C1979069|T201|COMP|51022-2|LNC|Blasts.cytoplasmic CD117/100 cells|Blasts.cytoplasmic CD117/100 cells
C1979071|T201|COMP|51023-0|LNC|Blasts.cytoplasmic CD117/100 cells|Blasts.cytoplasmic CD117/100 cells
C1979072|T201|COMP|51024-8|LNC|Blasts.cytoplasmic CD117/100 cells|Blasts.cytoplasmic CD117/100 cells
C1979073|T201|COMP|51025-5|LNC|Blasts.CD117/100 blasts|Blasts.CD117/100 blasts
C1979075|T201|COMP|51026-3|LNC|Blasts.CD117/100 blasts|Blasts.CD117/100 blasts
C1979076|T201|COMP|51027-1|LNC|Blasts.CD117/100 blasts|Blasts.CD117/100 blasts
C1979077|T201|COMP|51028-9|LNC|Blasts.CD117|Blasts.CD117
C1979079|T201|COMP|51029-7|LNC|Blasts.CD117|Blasts.CD117
C1979080|T201|COMP|51030-5|LNC|Blasts.CD117|Blasts.CD117
C1979081|T201|COMP|51031-3|LNC|Blasts.CD11a/100 blasts|Blasts.CD11a/100 blasts
C1979083|T201|COMP|51032-1|LNC|Blasts.CD11a/100 blasts|Blasts.CD11a/100 blasts
C1979084|T201|COMP|51033-9|LNC|Blasts.CD11a/100 blasts|Blasts.CD11a/100 blasts
C1979085|T201|COMP|51034-7|LNC|Blasts.CD11a|Blasts.CD11a
C1979087|T201|COMP|51035-4|LNC|Blasts.CD11a|Blasts.CD11a
C1979088|T201|COMP|51036-2|LNC|Blasts.CD11a|Blasts.CD11a
C1979089|T201|COMP|51037-0|LNC|Blasts.CD11b/100 blasts|Blasts.CD11b/100 blasts
C1979091|T201|COMP|51038-8|LNC|Blasts.CD11b/100 blasts|Blasts.CD11b/100 blasts
C1979092|T201|COMP|51039-6|LNC|Blasts.CD11b/100 blasts|Blasts.CD11b/100 blasts
C1979093|T201|COMP|51040-4|LNC|Blasts.CD11c/100 blasts|Blasts.CD11c/100 blasts
C1979095|T201|COMP|51041-2|LNC|Blasts.CD11c/100 blasts|Blasts.CD11c/100 blasts
C1979096|T201|COMP|51042-0|LNC|Blasts.CD11c/100 blasts|Blasts.CD11c/100 blasts
C1979097|T201|COMP|51043-8|LNC|Blasts.CD123/100 blasts|Blasts.CD123/100 blasts
C1979099|T201|COMP|51044-6|LNC|Blasts.CD123/100 blasts|Blasts.CD123/100 blasts
C1979100|T201|COMP|51045-3|LNC|Blasts.CD123/100 blasts|Blasts.CD123/100 blasts
C1979101|T201|COMP|51046-1|LNC|Blasts.CD123|Blasts.CD123
C1979103|T201|COMP|51047-9|LNC|Blasts.CD123|Blasts.CD123
C1979104|T201|COMP|51234-3|LNC|Cells.CD11c+CD19+/100 cells|Cells.CD11c+CD19+/100 cells
C1979105|T201|COMP|51235-0|LNC|Cells.CD13/100 cells|Cells.CD13/100 cells
C1979106|T201|COMP|51236-8|LNC|Cells.CD13/100 cells|Cells.CD13/100 cells
C1979107|T201|COMP|51237-6|LNC|Cells.CD13/100 cells|Cells.CD13/100 cells
C1979108|T201|COMP|51238-4|LNC|Cells.CD13/100 cells|Cells.CD13/100 cells
C1979109|T201|COMP|51239-2|LNC|Cells.CD13+CD33+/100 cells|Cells.CD13+CD33+/100 cells
C1979110|T201|COMP|51240-0|LNC|Cells.CD13+CD33+/100 cells|Cells.CD13+CD33+/100 cells
C1979111|T201|COMP|51241-8|LNC|Cells.CD13+CD33+HLA-DR+/100 cells|Cells.CD13+CD33+HLA-DR+/100 cells
C1979113|T201|COMP|51242-6|LNC|Cells.CD13+CD33+HLA-DR+/100 cells|Cells.CD13+CD33+HLA-DR+/100 cells
C1979114|T201|COMP|51243-4|LNC|Cells.CD13+CD33+HLA-DR+/100 cells|Cells.CD13+CD33+HLA-DR+/100 cells
C1979115|T201|COMP|51244-2|LNC|Cells.CD13+CD33+HLA-DR+/100 cells|Cells.CD13+CD33+HLA-DR+/100 cells
C1979116|T201|COMP|51245-9|LNC|Cells.CD13+CD33+HLA-DR+/100 cells|Cells.CD13+CD33+HLA-DR+/100 cells
C1979117|T201|COMP|51246-7|LNC|Cells.CD138/100 cells|Cells.CD138/100 cells
C1979118|T201|COMP|51048-7|LNC|Blasts.CD123|Blasts.CD123
C1979119|T201|COMP|51049-5|LNC|Blasts.CD126/100 blasts|Blasts.CD126/100 blasts
C1979121|T201|COMP|51050-3|LNC|Blasts.CD126/100 blasts|Blasts.CD126/100 blasts
C1979122|T201|COMP|51051-1|LNC|Blasts.CD126/100 blasts|Blasts.CD126/100 blasts
C1979123|T201|COMP|51052-9|LNC|Blasts.CD126|Blasts.CD126
C1979125|T201|COMP|51053-7|LNC|Blasts.CD126|Blasts.CD126
C1979126|T201|COMP|51054-5|LNC|Blasts.CD126|Blasts.CD126
C1979127|T201|COMP|51055-2|LNC|Blasts.CD127/100 blasts|Blasts.CD127/100 blasts
C1979129|T201|COMP|51056-0|LNC|Blasts.CD127/100 blasts|Blasts.CD127/100 blasts
C1979130|T201|COMP|51057-8|LNC|Blasts.CD127/100 blasts|Blasts.CD127/100 blasts
C1979131|T201|COMP|51058-6|LNC|Blasts.CD127|Blasts.CD127
C1979133|T201|COMP|51059-4|LNC|Blasts.CD127|Blasts.CD127
C1979134|T201|COMP|51060-2|LNC|Blasts.CD127|Blasts.CD127
C1979135|T201|COMP|51061-0|LNC|Blasts.cytoplasmic CD13/100 blasts|Blasts.cytoplasmic CD13/100 blasts
C1979137|T201|COMP|51062-8|LNC|Blasts.cytoplasmic CD13/100 blasts|Blasts.cytoplasmic CD13/100 blasts
C1979138|T201|COMP|51063-6|LNC|Blasts.cytoplasmic CD13/100 blasts|Blasts.cytoplasmic CD13/100 blasts
C1979139|T201|COMP|51064-4|LNC|Blasts.CD13/100 blasts|Blasts.CD13/100 blasts
C1979140|T201|COMP|51065-1|LNC|Blasts.CD13/100 blasts|Blasts.CD13/100 blasts
C1979141|T201|COMP|51066-9|LNC|Blasts.CD13|Blasts.CD13
C1979142|T201|COMP|51067-7|LNC|Blasts.CD13|Blasts.CD13
C1979143|T201|COMP|51068-5|LNC|Blasts.CD13|Blasts.CD13
C1979144|T201|COMP|51069-3|LNC|Blasts.CD135/100 blasts|Blasts.CD135/100 blasts
C1979146|T201|COMP|51070-1|LNC|Blasts.CD135/100 blasts|Blasts.CD135/100 blasts
C1979147|T201|COMP|51071-9|LNC|Blasts.CD135/100 blasts|Blasts.CD135/100 blasts
C1979148|T201|COMP|51072-7|LNC|Blasts.CD135|Blasts.CD135
C1979150|T201|COMP|51073-5|LNC|Blasts.CD135|Blasts.CD135
C1979151|T201|COMP|51074-3|LNC|Blasts.CD135|Blasts.CD135
C1979152|T201|COMP|51075-0|LNC|Blasts.CD14/100 blasts|Blasts.CD14/100 blasts
C1979153|T201|COMP|51076-8|LNC|Blasts.CD14/100 blasts|Blasts.CD14/100 blasts
C1979154|T201|COMP|51077-6|LNC|Blasts.CD14|Blasts.CD14
C1979155|T201|COMP|51078-4|LNC|Blasts.CD14|Blasts.CD14
C1979156|T201|COMP|51079-2|LNC|Blasts.CD14|Blasts.CD14
C1979157|T201|COMP|51080-0|LNC|Blasts.CD15/100 blasts|Blasts.CD15/100 blasts
C1979159|T201|COMP|51081-8|LNC|Blasts.CD15/100 blasts|Blasts.CD15/100 blasts
C1979160|T201|COMP|51082-6|LNC|Blasts.CD15/100 blasts|Blasts.CD15/100 blasts
C1979161|T201|COMP|51083-4|LNC|Blasts.CD15|Blasts.CD15
C1979163|T201|COMP|51084-2|LNC|Blasts.CD15|Blasts.CD15
C1979164|T201|COMP|51085-9|LNC|Blasts.CD15|Blasts.CD15
C1979165|T201|COMP|51086-7|LNC|Blasts.CD16/100 blasts|Blasts.CD16/100 blasts
C1979167|T201|COMP|51087-5|LNC|Blasts.CD16/100 blasts|Blasts.CD16/100 blasts
C1979168|T201|COMP|51088-3|LNC|Blasts.CD16/100 blasts|Blasts.CD16/100 blasts
C1979169|T201|COMP|51089-1|LNC|Blasts.cytoplasmic CD179a/100 blasts|Blasts.cytoplasmic CD179a/100 blasts
C1979171|T201|COMP|51090-9|LNC|Blasts.cytoplasmic CD179a/100 blasts|Blasts.cytoplasmic CD179a/100 blasts
C1979172|T201|COMP|51091-7|LNC|Blasts.cytoplasmic CD179a/100 blasts|Blasts.cytoplasmic CD179a/100 blasts
C1979173|T201|COMP|51092-5|LNC|Blasts.cytoplasmic CD179a|Blasts.cytoplasmic CD179a
C1979175|T201|COMP|51093-3|LNC|Blasts.cytoplasmic CD179a|Blasts.cytoplasmic CD179a
C1979176|T201|COMP|51094-1|LNC|Blasts.cytoplasmic CD179a|Blasts.cytoplasmic CD179a
C1979177|T201|COMP|51095-8|LNC|Blasts.CD179a/100 blasts|Blasts.CD179a/100 blasts
C1979179|T201|COMP|51096-6|LNC|Blasts.CD179a/100 blasts|Blasts.CD179a/100 blasts
C1979180|T201|COMP|51097-4|LNC|Blasts.CD179a/100 blasts|Blasts.CD179a/100 blasts
C1979181|T201|COMP|51098-2|LNC|Blasts.CD179a|Blasts.CD179a
C1979183|T201|COMP|51099-0|LNC|Blasts.CD179a|Blasts.CD179a
C1979184|T201|COMP|51100-6|LNC|Blasts.CD179a|Blasts.CD179a
C1979185|T201|COMP|51101-4|LNC|Blasts.CD19/100 blasts|Blasts.CD19/100 blasts
C1979186|T201|COMP|51102-2|LNC|Blasts.CD19/100 blasts|Blasts.CD19/100 blasts
C1979187|T201|COMP|51103-0|LNC|Blasts.CD19|Blasts.CD19
C1979188|T201|COMP|51104-8|LNC|Blasts.CD19|Blasts.CD19
C1979189|T201|COMP|51105-5|LNC|Blasts.CD19|Blasts.CD19
C1979190|T201|COMP|51106-3|LNC|Blasts.CD1a/100 blasts|Blasts.CD1a/100 blasts
C1979192|T201|COMP|51107-1|LNC|Blasts.CD1a/100 blasts|Blasts.CD1a/100 blasts
C1979193|T201|COMP|51108-9|LNC|Blasts.CD1a/100 blasts|Blasts.CD1a/100 blasts
C1979194|T201|COMP|51109-7|LNC|Blasts.cytoplasmic CD2/100 blasts|Blasts.cytoplasmic CD2/100 blasts
C1979196|T201|COMP|51142-8|LNC|Blasts.cytoplasmic CD3|Blasts.cytoplasmic CD3
C1979197|T201|COMP|51143-6|LNC|Blasts.CD3/100 blasts|Blasts.CD3/100 blasts
C1979199|T201|COMP|51144-4|LNC|Blasts.CD3/100 blasts|Blasts.CD3/100 blasts
C1979200|T201|COMP|51145-1|LNC|Blasts.CD3/100 blasts|Blasts.CD3/100 blasts
C1979201|T201|COMP|51146-9|LNC|Blasts.CD3|Blasts.CD3
C1979203|T201|COMP|51147-7|LNC|Blasts.CD3|Blasts.CD3
C1979204|T201|COMP|51148-5|LNC|Blasts.CD3|Blasts.CD3
C1979205|T201|COMP|51149-3|LNC|Blasts.CD3+CD16+CD56+/100 blasts|Blasts.CD3+CD16+CD56+/100 blasts
C1979207|T201|COMP|51150-1|LNC|Blasts.CD3+CD16+CD56+/100 blasts|Blasts.CD3+CD16+CD56+/100 blasts
C1979208|T201|COMP|51151-9|LNC|Blasts.CD3+CD16+CD56+/100 blasts|Blasts.CD3+CD16+CD56+/100 blasts
C1979209|T201|COMP|51152-7|LNC|Blasts.CD30/100 blasts|Blasts.CD30/100 blasts
C1979211|T201|COMP|51153-5|LNC|Blasts.CD30/100 blasts|Blasts.CD30/100 blasts
C1979212|T201|COMP|51154-3|LNC|Blasts.CD30/100 blasts|Blasts.CD30/100 blasts
C1979213|T201|COMP|51155-0|LNC|Blasts.CD33/100 blasts|Blasts.CD33/100 blasts
C1979214|T201|COMP|51156-8|LNC|Blasts.CD33/100 blasts|Blasts.CD33/100 blasts
C1979215|T201|COMP|51157-6|LNC|Blasts.CD33|Blasts.CD33
C1979216|T201|COMP|51158-4|LNC|Blasts.CD33|Blasts.CD33
C1979217|T201|COMP|51159-2|LNC|Blasts.CD33|Blasts.CD33
C1979218|T201|COMP|51160-0|LNC|Blasts.CD33+CD34+/100 blasts|Blasts.CD33+CD34+/100 blasts
C1979220|T201|COMP|51161-8|LNC|Blasts.cytoplasmic CD34/100 blasts|Blasts.cytoplasmic CD34/100 blasts
C1979222|T201|COMP|51162-6|LNC|Blasts.CD34/100 blasts|Blasts.CD34/100 blasts
C1979223|T201|COMP|51163-4|LNC|Blasts.CD34/100 blasts|Blasts.CD34/100 blasts
C1979224|T201|COMP|51164-2|LNC|Blasts.CD34|Blasts.CD34
C1979225|T201|COMP|51165-9|LNC|Blasts.CD34|Blasts.CD34
C1979226|T201|COMP|51166-7|LNC|Blasts.CD34|Blasts.CD34
C1979227|T201|COMP|51167-5|LNC|Blasts.CD34+CD117+/100 blasts|Blasts.CD34+CD117+/100 blasts
C1979229|T201|COMP|51168-3|LNC|Blasts.CD34+CD117+/100 blasts|Blasts.CD34+CD117+/100 blasts
C1979230|T201|COMP|51169-1|LNC|Blasts.CD34+CD117+/100 blasts|Blasts.CD34+CD117+/100 blasts
C1979231|T201|COMP|51170-9|LNC|Blasts.CD34+CD117+|Blasts.CD34+CD117+
C1979233|T201|COMP|51171-7|LNC|Blasts.CD34+CD117+|Blasts.CD34+CD117+
C1979234|T201|COMP|51172-5|LNC|Blasts.CD34+CD117+|Blasts.CD34+CD117+
C1979235|T201|COMP|51173-3|LNC|Blasts.CD36/100 blasts|Blasts.CD36/100 blasts
C1979237|T201|COMP|51174-1|LNC|Blasts.CD36/100 blasts|Blasts.CD36/100 blasts
C1979238|T201|COMP|51175-8|LNC|Blasts.CD36/100 blasts|Blasts.CD36/100 blasts
C1979239|T201|COMP|51176-6|LNC|Blasts.CD36|Blasts.CD36
C1979241|T201|COMP|51177-4|LNC|Blasts.CD36|Blasts.CD36
C1979242|T201|COMP|51178-2|LNC|Blasts.CD36|Blasts.CD36
C1979243|T201|COMP|51179-0|LNC|Blasts.CD36+CD235a+/100 blasts|Blasts.CD36+CD235a+/100 blasts
C1979245|T201|COMP|51180-8|LNC|Blasts.CD36+CD235a+/100 blasts|Blasts.CD36+CD235a+/100 blasts
C1979246|T201|COMP|51181-6|LNC|Blasts.CD1|Blasts.CD1
C1979247|T201|COMP|51182-4|LNC|Blasts.CD10|Blasts.CD10
C1979248|T201|COMP|51183-2|LNC|CD117 Ag|CD117 Ag
C1979249|T201|COMP|51184-0|LNC|CD117 Ag|CD117 Ag
C1979250|T201|COMP|51185-7|LNC|CD117 Ag|CD117 Ag
C1979251|T201|COMP|51186-5|LNC|CD15 Ag|CD15 Ag
C1979252|T201|COMP|51187-3|LNC|CD15 Ag|CD15 Ag
C1979253|T201|COMP|51188-1|LNC|CD15 Ag|CD15 Ag
C1979254|T201|COMP|51189-9|LNC|4-Hydroxybupivacaine|4-Hydroxybupivacaine
C1979255|T201|COMP|51190-7|LNC|Albumin|Albumin
C1979256|T201|COMP|51191-5|LNC|Antimony|Antimony
C1979257|T201|COMP|51192-3|LNC|Barium|Barium
C1979258|T201|COMP|51193-1|LNC|Cadmium|Cadmium
C1979259|T201|COMP|51194-9|LNC|Cobalt|Cobalt
C1979260|T201|COMP|51195-6|LNC|Desbutylbupivacaine|Desbutylbupivacaine
C1979261|T201|COMP|51196-4|LNC|Hemoglobin A1/Hemoglobin.total|Hemoglobin A1/Hemoglobin.total
C1979262|T201|COMP|51197-2|LNC|Iron|Iron
C1979263|T201|COMP|51198-0|LNC|Manganese|Manganese
C1979264|T201|COMP|51199-8|LNC|Molybdenum|Molybdenum
C1979265|T201|COMP|51200-4|LNC|Nickel|Nickel
C1979266|T201|COMP|51201-2|LNC|Palladium|Palladium
C1979267|T201|COMP|51202-0|LNC|Platinum|Platinum
C1979268|T201|COMP|51203-8|LNC|Ropivacaine|Ropivacaine
C1979269|T201|COMP|51204-6|LNC|Silicon|Silicon
C1979270|T201|COMP|51205-3|LNC|Sodium|Sodium
C1979271|T201|COMP|51206-1|LNC|Strontium|Strontium
C1979272|T201|COMP|51207-9|LNC|Thallium|Thallium
C1979273|T201|COMP|51208-7|LNC|Tin|Tin
C1979274|T201|COMP|51209-5|LNC|Tin|Tin
C1979275|T201|COMP|51210-3|LNC|Titanium|Titanium
C1979276|T201|COMP|51211-1|LNC|Uranium|Uranium
C1979277|T201|COMP|51212-9|LNC|Vanadium|Vanadium
C1979278|T201|COMP|51213-7|LNC|Acetaminophen crystals|Acetaminophen crystals
C1979279|T201|COMP|51214-5|LNC|Cells.CD10/100 cells|Cells.CD10/100 cells
C1979280|T201|COMP|51215-2|LNC|Cells.CD10/100 cells|Cells.CD10/100 cells
C1979281|T201|COMP|51216-0|LNC|Cells.CD10/100 cells|Cells.CD10/100 cells
C1979282|T201|COMP|51217-8|LNC|Cells.CD10/100 cells|Cells.CD10/100 cells
C1979283|T201|COMP|51218-6|LNC|Cells.CD10+CD19+/100 cells|Cells.CD10+CD19+/100 cells
C1979284|T201|COMP|51219-4|LNC|Cells.CD10+CD19+/100 cells|Cells.CD10+CD19+/100 cells
C1979285|T201|COMP|51220-2|LNC|Cells.CD103/100 cells|Cells.CD103/100 cells
C1979286|T201|COMP|51221-0|LNC|Cells.CD103/100 cells|Cells.CD103/100 cells
C1979287|T201|COMP|51222-8|LNC|Cells.CD105/100 cells|Cells.CD105/100 cells
C1979288|T201|COMP|51223-6|LNC|Cells.CD105/100 cells|Cells.CD105/100 cells
C1979289|T201|COMP|51224-4|LNC|Cells.CD105/100 cells|Cells.CD105/100 cells
C1979290|T201|COMP|51225-1|LNC|Cells.CD105/100 cells|Cells.CD105/100 cells
C1979291|T201|COMP|51226-9|LNC|Cells.CD117/100 cells|Cells.CD117/100 cells
C1979292|T201|COMP|51227-7|LNC|Cells.CD11b/100 cells|Cells.CD11b/100 cells
C1979293|T201|COMP|51228-5|LNC|Cells.CD11b/100 cells|Cells.CD11b/100 cells
C1979294|T201|COMP|51229-3|LNC|Cells.CD11b/100 cells|Cells.CD11b/100 cells
C1979295|T201|COMP|51230-1|LNC|Cells.CD11b/100 cells|Cells.CD11b/100 cells
C1979296|T201|COMP|51231-9|LNC|Cells.CD11c/100 cells|Cells.CD11c/100 cells
C1979297|T201|COMP|51232-7|LNC|Cells.CD11c/100 cells|Cells.CD11c/100 cells
C1979298|T201|COMP|51233-5|LNC|Cells.CD11c+CD19+/100 cells|Cells.CD11c+CD19+/100 cells
C1979299|T201|COMP|51247-5|LNC|Cells.CD14/100 cells|Cells.CD14/100 cells
C1979300|T201|COMP|51248-3|LNC|Cells.CD14/100 cells|Cells.CD14/100 cells
C1979301|T201|COMP|51249-1|LNC|Cells.CD15/100 cells|Cells.CD15/100 cells
C1979302|T201|COMP|51250-9|LNC|Cells.CD15/100 cells|Cells.CD15/100 cells
C1979303|T201|COMP|51251-7|LNC|Cells.CD15/100 cells|Cells.CD15/100 cells
C1979304|T201|COMP|51252-5|LNC|Cells.CD15/100 cells|Cells.CD15/100 cells
C1979305|T201|COMP|51253-3|LNC|Cells.CD16+CD56+/100 cells|Cells.CD16+CD56+/100 cells
C1979306|T201|COMP|51254-1|LNC|Cells.CD16+CD56+/100 cells|Cells.CD16+CD56+/100 cells
C1979307|T201|COMP|51255-8|LNC|Cells.CD16+CD56+/100 cells|Cells.CD16+CD56+/100 cells
C1979308|T201|COMP|51256-6|LNC|Cells.CD16+CD57+/100 cells|Cells.CD16+CD57+/100 cells
C1979309|T201|COMP|51257-4|LNC|Cells.CD16+CD57+/100 cells|Cells.CD16+CD57+/100 cells
C1979310|T201|COMP|51258-2|LNC|Cells.CD16+CD57+/100 cells|Cells.CD16+CD57+/100 cells
C1979311|T201|COMP|51259-0|LNC|Cells.CD16+CD57+/100 cells|Cells.CD16+CD57+/100 cells
C1979312|T201|COMP|51260-8|LNC|Cells.CD16b/100 cells|Cells.CD16b/100 cells
C1979313|T201|COMP|51261-6|LNC|Cells.CD16b/100 cells|Cells.CD16b/100 cells
C1979314|T201|COMP|51262-4|LNC|Cells.CD16b/100 cells|Cells.CD16b/100 cells
C1979315|T201|COMP|51263-2|LNC|Cells.CD16b/100 cells|Cells.CD16b/100 cells
C1979316|T201|COMP|51264-0|LNC|Cells.CD19/100 cells|Cells.CD19/100 cells
C1979317|T201|COMP|51274-9|LNC|Cells.CD3+CD16+/100 cells|Cells.CD3+CD16+/100 cells
C1979318|T201|COMP|51275-6|LNC|Cells.CD3+CD16+/100 cells|Cells.CD3+CD16+/100 cells
C1979319|T201|COMP|51276-4|LNC|Cells.CD3+CD16+/100 cells|Cells.CD3+CD16+/100 cells
C1979320|T201|COMP|51277-2|LNC|Cells.CD3+CD16+/100 cells|Cells.CD3+CD16+/100 cells
C1979321|T201|COMP|51278-0|LNC|Cells.CD3+CD56+/100 cells|Cells.CD3+CD56+/100 cells
C1979322|T201|COMP|51279-8|LNC|Cells.CD3+CD56+/100 cells|Cells.CD3+CD56+/100 cells
C1979323|T201|COMP|51280-6|LNC|Cells.CD3+CD56+/100 cells|Cells.CD3+CD56+/100 cells
C1979324|T201|COMP|51281-4|LNC|Cells.CD3+CD56+/100 cells|Cells.CD3+CD56+/100 cells
C1979326|T201|COMP|51283-0|LNC|Cells.CD3+CD57+/100 cells|Cells.CD3+CD57+/100 cells
C1979327|T201|COMP|51284-8|LNC|Cells.CD3+CD57+/100 cells|Cells.CD3+CD57+/100 cells
C1979328|T201|COMP|51285-5|LNC|Cells.CD3+CD57+/100 cells|Cells.CD3+CD57+/100 cells
C1979329|T201|COMP|51286-3|LNC|Cells.CD3+CD57+/100 cells|Cells.CD3+CD57+/100 cells
C1979330|T201|COMP|51287-1|LNC|Cells.CD30/100 cells|Cells.CD30/100 cells
C1979331|T201|COMP|51288-9|LNC|Cells.CD30/100 cells|Cells.CD30/100 cells
C1979332|T201|COMP|51289-7|LNC|Cells.CD30/100 cells|Cells.CD30/100 cells
C1979333|T201|COMP|51290-5|LNC|Cells.CD30/100 cells|Cells.CD30/100 cells
C1979334|T201|COMP|51291-3|LNC|Cells.CD33/100 cells|Cells.CD33/100 cells
C1979335|T201|COMP|51292-1|LNC|Cells.CD33/100 cells|Cells.CD33/100 cells
C1979336|T201|COMP|51293-9|LNC|Cells.CD33/100 cells|Cells.CD33/100 cells
C1979337|T201|COMP|51294-7|LNC|Cells.CD33/100 cells|Cells.CD33/100 cells
C1979338|T201|COMP|51295-4|LNC|Cells.CD36/100 cells|Cells.CD36/100 cells
C1979339|T201|COMP|51296-2|LNC|Cells.CD38/100 cells|Cells.CD38/100 cells
C1979340|T201|COMP|51297-0|LNC|Cells.CD38/100 cells|Cells.CD38/100 cells
C1979341|T201|COMP|51298-8|LNC|Cells.CD38/100 cells|Cells.CD38/100 cells
C1979342|T201|COMP|51299-6|LNC|Cells.CD38/100 cells|Cells.CD38/100 cells
C1979343|T201|COMP|51300-2|LNC|Cells.CD3+CD4+/100 cells|Cells.CD3+CD4+/100 cells
C1979344|T201|COMP|51301-0|LNC|Cells.CD4/100 cells|Cells.CD4/100 cells
C1979345|T201|COMP|51302-8|LNC|Cells.CD4+CD7-/100 cells|Cells.CD4+CD7-/100 cells
C1979347|T201|COMP|51303-6|LNC|Cells.CD4+CD7-/100 cells|Cells.CD4+CD7-/100 cells
C1979348|T201|COMP|51304-4|LNC|Cells.CD4+CD7-/100 cells|Cells.CD4+CD7-/100 cells
C1979349|T201|COMP|51305-1|LNC|Cells.CD4+CD7-/100 cells|Cells.CD4+CD7-/100 cells
C1979350|T201|COMP|51306-9|LNC|Cells.CD4+CD7-/100 cells|Cells.CD4+CD7-/100 cells
C1979351|T201|COMP|51307-7|LNC|Cells.CD4+CD7-CD26-/100 cells|Cells.CD4+CD7-CD26-/100 cells
C1979353|T201|COMP|51308-5|LNC|Cells.CD4+CD7-CD26-/100 cells|Cells.CD4+CD7-CD26-/100 cells
C1979354|T201|COMP|51309-3|LNC|Cells.CD4+CD7-CD26-/100 cells|Cells.CD4+CD7-CD26-/100 cells
C1979355|T201|COMP|51310-1|LNC|Cells.CD4+CD7-CD26-/100 cells|Cells.CD4+CD7-CD26-/100 cells
C1979356|T201|COMP|51311-9|LNC|Cells.CD4+CD7-CD26-/100 cells|Cells.CD4+CD7-CD26-/100 cells
C1979357|T201|COMP|51312-7|LNC|Cells.CD4+CD7-CD49d-/100 cells|Cells.CD4+CD7-CD49d-/100 cells
C1979359|T201|COMP|51313-5|LNC|Cells.CD4+CD7-CD49d-/100 cells|Cells.CD4+CD7-CD49d-/100 cells
C1979360|T201|COMP|51314-3|LNC|Cells.CD4+CD7-CD49d-/100 cells|Cells.CD4+CD7-CD49d-/100 cells
C1979361|T201|COMP|51315-0|LNC|Cells.CD4+CD7-CD49d-/100 cells|Cells.CD4+CD7-CD49d-/100 cells
C1979362|T201|COMP|51316-8|LNC|Cells.CD4+CD7-CD49d-/100 cells|Cells.CD4+CD7-CD49d-/100 cells
C1979363|T201|COMP|51317-6|LNC|Cells.CD41/100 cells|Cells.CD41/100 cells
C1979364|T201|COMP|51318-4|LNC|Cells.CD41/100 cells|Cells.CD41/100 cells
C1979365|T201|COMP|51319-2|LNC|Cells.CD41/100 cells|Cells.CD41/100 cells
C1979366|T201|COMP|51320-0|LNC|Cells.CD41/100 cells|Cells.CD41/100 cells
C1979367|T201|COMP|51321-8|LNC|Cells.CD42/100 cells|Cells.CD42/100 cells
C1979368|T201|COMP|51322-6|LNC|Cells.CD42/100 cells|Cells.CD42/100 cells
C1979369|T201|COMP|51323-4|LNC|Cells.CD42/100 cells|Cells.CD42/100 cells
C1979370|T201|COMP|51324-2|LNC|Cells.CD42/100 cells|Cells.CD42/100 cells
C1979371|T201|COMP|51325-9|LNC|Cells.CD42b/100 cells|Cells.CD42b/100 cells
C1979372|T201|COMP|51326-7|LNC|Cells.CD42b/100 cells|Cells.CD42b/100 cells
C1979373|T201|COMP|51327-5|LNC|Cells.CD42b/100 cells|Cells.CD42b/100 cells
C1979374|T201|COMP|51328-3|LNC|Cells.CD42b/100 cells|Cells.CD42b/100 cells
C1979375|T201|COMP|51329-1|LNC|Cells.CD43/100 cells|Cells.CD43/100 cells
C1979376|T201|COMP|51330-9|LNC|Cells.CD43/100 cells|Cells.CD43/100 cells
C1979377|T201|COMP|51331-7|LNC|Cells.CD43/100 cells|Cells.CD43/100 cells
C1979378|T201|COMP|51332-5|LNC|Cells.CD43/100 cells|Cells.CD43/100 cells
C1979379|T201|COMP|51333-3|LNC|Cells.CD19+CD43+/100 cells|Cells.CD19+CD43+/100 cells
C1979381|T201|COMP|51334-1|LNC|Cells.CD19+CD43+/100 cells|Cells.CD19+CD43+/100 cells
C1979382|T201|COMP|51335-8|LNC|Cells.CD19+CD43+/100 cells|Cells.CD19+CD43+/100 cells
C1979383|T201|COMP|51336-6|LNC|Cells.CD19+CD43+/100 cells|Cells.CD19+CD43+/100 cells
C1979384|T201|COMP|51337-4|LNC|Cells.CD19+CD43+/100 cells|Cells.CD19+CD43+/100 cells
C1979385|T201|COMP|51338-2|LNC|Cells.CD45/100 cells|Cells.CD45/100 cells
C1979386|T201|COMP|51347-3|LNC|Cells.CD56+CD57+/100 cells|Cells.CD56+CD57+/100 cells
C1979387|T201|COMP|51348-1|LNC|Cells.CD56+CD57+/100 cells|Cells.CD56+CD57+/100 cells
C1979388|T201|COMP|51349-9|LNC|Cells.CD56+CD57+/100 cells|Cells.CD56+CD57+/100 cells
C1979389|T201|COMP|51350-7|LNC|Cells.CD57/100 cells|Cells.CD57/100 cells
C1979390|T201|COMP|51351-5|LNC|Cells.CD57/100 cells|Cells.CD57/100 cells
C1979391|T201|COMP|51352-3|LNC|Cells.CD19+CD58+/100 cells|Cells.CD19+CD58+/100 cells
C1979393|T201|COMP|51353-1|LNC|Cells.CD19+CD58+/100 cells|Cells.CD19+CD58+/100 cells
C1979394|T201|COMP|51354-9|LNC|Cells.CD19+CD58+/100 cells|Cells.CD19+CD58+/100 cells
C1979395|T201|COMP|51355-6|LNC|Cells.CD19+CD58+/100 cells|Cells.CD19+CD58+/100 cells
C1979396|T201|COMP|51356-4|LNC|Cells.CD19+CD58+/100 cells|Cells.CD19+CD58+/100 cells
C1979397|T201|COMP|51357-2|LNC|Cells.CD59/100 cells|Cells.CD59/100 cells
C1979398|T201|COMP|51358-0|LNC|Cells.CD59/100 cells|Cells.CD59/100 cells
C1979399|T201|COMP|51359-8|LNC|Cells.CD61/100 cells|Cells.CD61/100 cells
C1979400|T201|COMP|51360-6|LNC|Cells.CD61/100 cells|Cells.CD61/100 cells
C1979401|T201|COMP|51361-4|LNC|Cells.CD61/100 cells|Cells.CD61/100 cells
C1979402|T201|COMP|51362-2|LNC|Cells.CD61/100 cells|Cells.CD61/100 cells
C1979403|T201|COMP|51363-0|LNC|Cells.CD64/100 cells|Cells.CD64/100 cells
C1979404|T201|COMP|51364-8|LNC|Cells.CD64/100 cells|Cells.CD64/100 cells
C1979405|T201|COMP|51365-5|LNC|Cells.CD64/100 cells|Cells.CD64/100 cells
C1979406|T201|COMP|51366-3|LNC|Cells.CD64/100 cells|Cells.CD64/100 cells
C1979407|T201|COMP|51367-1|LNC|Cells.CD79a/100 cells|Cells.CD79a/100 cells
C1979408|T201|COMP|51368-9|LNC|Cells.CD79a/100 cells|Cells.CD79a/100 cells
C1979409|T201|COMP|51369-7|LNC|Cells.CD79b/100 cells|Cells.CD79b/100 cells
C1979411|T201|COMP|51370-5|LNC|Cells.CD8+HLA-DR+/100 cells|Cells.CD8+HLA-DR+/100 cells
C1979412|T201|COMP|51371-3|LNC|Cells.CD8+HLA-DR+/100 cells|Cells.CD8+HLA-DR+/100 cells
C1979413|T201|COMP|51372-1|LNC|Cells.CD8+HLA-DR+/100 cells|Cells.CD8+HLA-DR+/100 cells
C1979414|T201|COMP|51373-9|LNC|Cells.CD8+HLA-DR+/100 cells|Cells.CD8+HLA-DR+/100 cells
C1979415|T201|COMP|51374-7|LNC|Cells.CD9/100 cells|Cells.CD9/100 cells
C1979416|T201|COMP|51375-4|LNC|Cells.CD9/100 cells|Cells.CD9/100 cells
C1979417|T201|COMP|51376-2|LNC|Cells.CD9/100 cells|Cells.CD9/100 cells
C1979418|T201|COMP|51377-0|LNC|Cells.CD9/100 cells|Cells.CD9/100 cells
C1979419|T201|COMP|51378-8|LNC|Cells.HLA-DR+/100 cells|Cells.HLA-DR+/100 cells
C1979420|T201|COMP|51379-6|LNC|Cells.HLA-DR+/100 cells|Cells.HLA-DR+/100 cells
C1979421|T201|COMP|51380-4|LNC|Cells.HLA-DR+/100 cells|Cells.HLA-DR+/100 cells
C1979422|T201|COMP|51381-2|LNC|Cells.HLA-DR+/100 cells|Cells.HLA-DR+/100 cells
C1979423|T201|COMP|51382-0|LNC|Erythrocytes|Erythrocytes
C1979424|T201|COMP|51383-8|LNC|Leukocytes other|Leukocytes other
C1979425|T201|COMP|51384-6|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C1979426|T201|COMP|51400-0|LNC|Cells.CD65w/100 cells|Cells.CD65w/100 cells
C1979427|T201|COMP|51401-8|LNC|Cells.CD81/100 cells|Cells.CD81/100 cells
C1979429|T201|COMP|51402-6|LNC|Cells.CD81/100 cells|Cells.CD81/100 cells
C1979430|T201|COMP|51403-4|LNC|Cells.CD81/100 cells|Cells.CD81/100 cells
C1979431|T201|COMP|51404-2|LNC|Cells.CD81/100 cells|Cells.CD81/100 cells
C1979432|T201|COMP|51405-9|LNC|Cells.CD81/100 cells|Cells.CD81/100 cells
C1979433|T201|COMP|51406-7|LNC|Immunoglobulin light chains.free|Immunoglobulin light chains.free
C1979438|T201|COMP|51409-1|LNC|Fosamprenavir+Ritonavir|Fosamprenavir+Ritonavir
C1979440|T201|COMP|51410-9|LNC|Environmental stressors panel|Environmental stressors panel
C1979442|T201|COMP|51411-7|LNC|Environmental stressors panel|Environmental stressors panel
C1979443|T201|COMP|51420-8|LNC|17-Hydroxyprogesterone^pre or post XXX challenge|17-Hydroxyprogesterone^pre or post XXX challenge
C1979444|T201|COMP|51421-6|LNC|Testosterone^pre or post XXX challenge|Testosterone^pre or post XXX challenge
C1979445|T201|COMP|51422-4|LNC|Aldosterone^pre or post XXX challenge|Aldosterone^pre or post XXX challenge
C1979446|T201|COMP|51423-2|LNC|Corticotropin^pre or post XXX challenge|Corticotropin^pre or post XXX challenge
C1979447|T201|COMP|51424-0|LNC|Cortisol^pre or post XXX challenge|Cortisol^pre or post XXX challenge
C1979448|T201|COMP|51425-7|LNC|EPINEPHrine^pre or post XXX challenge|EPINEPHrine^pre or post XXX challenge
C1979449|T201|COMP|51426-5|LNC|Glucose^pre or post XXX challenge|Glucose^pre or post XXX challenge
C1979450|T201|COMP|51427-3|LNC|Insulin^pre or post XXX challenge|Insulin^pre or post XXX challenge
C1979451|T201|COMP|51428-1|LNC|Lactate^pre or post XXX challenge|Lactate^pre or post XXX challenge
C1979452|T201|COMP|51429-9|LNC|Norepinephrine^pre or post XXX challenge|Norepinephrine^pre or post XXX challenge
C1979453|T201|COMP|51430-7|LNC|Calcitonin^pre or post XXX challenge|Calcitonin^pre or post XXX challenge
C1979454|T201|COMP|51431-5|LNC|Gastrin^pre or post XXX challenge|Gastrin^pre or post XXX challenge
C1979455|T201|COMP|51432-3|LNC|Prolactin^pre or post XXX challenge|Prolactin^pre or post XXX challenge
C1979456|T201|COMP|51433-1|LNC|Renin^pre or post XXX challenge|Renin^pre or post XXX challenge
C1979457|T201|COMP|51434-9|LNC|Somatotropin^pre or post XXX challenge|Somatotropin^pre or post XXX challenge
C1979458|T201|COMP|51435-6|LNC|Protein.monoclonal band 1|Protein.monoclonal band 1
C1979460|T201|COMP|51436-4|LNC|Protein.monoclonal|Protein.monoclonal
C1979461|T201|COMP|51437-2|LNC|Protein.monoclonal band 2|Protein.monoclonal band 2
C1979462|T201|COMP|51438-0|LNC|Protein.monoclonal band 2|Protein.monoclonal band 2
C1979463|T201|COMP|51439-8|LNC|Protein.monoclonal band 3|Protein.monoclonal band 3
C1979464|T201|COMP|51440-6|LNC|Protein.monoclonal band 3|Protein.monoclonal band 3
C1979465|T201|COMP|51441-4|LNC|Macroprolactin/Prolactin|Macroprolactin/Prolactin
C1979466|T201|COMP|51442-2|LNC|Domperidone|Domperidone
C1979467|T201|COMP|51443-0|LNC|Cells.CD117|Cells.CD117
C1979468|T201|COMP|51444-8|LNC|Cells.CD19+CD38+|Cells.CD19+CD38+
C1979469|T201|COMP|51445-5|LNC|Cells.CD41a|Cells.CD41a
C1979470|T201|COMP|51446-3|LNC|Cells.CD64|Cells.CD64
C1979471|T201|COMP|51447-1|LNC|Cells.CD79a|Cells.CD79a
C1979472|T201|COMP|51448-9|LNC|Dihydrocodeine+Hydrocodol|Dihydrocodeine+Hydrocodol
C1979473|T201|COMP|51449-7|LNC|Paragonimus sp Ab|Paragonimus sp Ab
C1979474|T201|COMP|51450-5|LNC|Paragonimus sp Ab|Paragonimus sp Ab
C1979475|T201|COMP|51451-3|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C1979476|T201|COMP|51452-1|LNC|Coccidioides immitis Ab|Coccidioides immitis Ab
C1979477|T201|COMP|51453-9|LNC|Coxsackievirus A9+B1+B2+B3+B4+B5+B6 Ab|Coxsackievirus A9+B1+B2+B3+B4+B5+B6 Ab
C1979478|T201|COMP|51454-7|LNC|Epstein Barr virus early diffuse Ab|Epstein Barr virus early diffuse Ab
C1979479|T201|COMP|51455-4|LNC|Filaria Ab.IgG1|Filaria Ab.IgG1
C1979480|T201|COMP|51456-2|LNC|Filaria Ab.IgG2|Filaria Ab.IgG2
C1979481|T201|COMP|51457-0|LNC|Filaria Ab.IgG3|Filaria Ab.IgG3
C1979482|T201|COMP|51458-8|LNC|Hepatitis D virus Ab.IgG|Hepatitis D virus Ab.IgG
C1979483|T201|COMP|51459-6|LNC|Hepatitis E virus Ab|Hepatitis E virus Ab
C1979484|T201|COMP|51460-4|LNC|Influenza virus A H16 Ab|Influenza virus A H16 Ab
C1979485|T201|COMP|51469-5|LNC|Plasmodium vivax Ab.IgG|Plasmodium vivax Ab.IgG
C1979486|T201|COMP|51470-3|LNC|Satratoxin Ab.IgM|Satratoxin Ab.IgM
C1979487|T201|COMP|51471-1|LNC|Sporothrix schenckii Ab|Sporothrix schenckii Ab
C1979490|T201|COMP|51474-5|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1979491|T201|COMP|51475-2|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C1979492|T201|COMP|51476-0|LNC|ABCB4 gene targeted mutation analysis|ABCB4 gene targeted mutation analysis
C1979493|T201|COMP|51477-8|LNC|Coccidioides sp Ab.IgM|Coccidioides sp Ab.IgM
C1979494|T201|COMP|51478-6|LNC|Mucus|Mucus
C1979495|T201|COMP|51479-4|LNC|Spermatozoa|Spermatozoa
C1979496|T201|COMP|51480-2|LNC|Bacteria|Bacteria
C1979497|T201|COMP|51481-0|LNC|Yeast|Yeast
C1979498|T201|COMP|51482-8|LNC|Crystals|Crystals
C1979499|T201|COMP|51483-6|LNC|Casts|Casts
C1979500|T201|COMP|51484-4|LNC|Hyaline casts|Hyaline casts
C1979501|T201|COMP|51485-1|LNC|Epithelial cells.non-squamous|Epithelial cells.non-squamous
C1979502|T201|COMP|51486-9|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C1979503|T201|COMP|51487-7|LNC|Leukocytes|Leukocytes
C2003845|T201|COMP|51282-2|LNC|Cells.CD3+CD57+/100 cells|Cells.CD3+CD57+/100 cells
C2004100|T201|COMP|22683-7|LNC|Phenylalanine/Creatinine|Phenylalanine/Creatinine
C2004114|T201|COMP|24167-9|LNC|Rat Ab.IgE|Rat Ab.IgE
C2004115|T201|COMP|13191-2|LNC|Rheumatoid factor|Rheumatoid factor
C2359798|T201|COMP|51501-5|LNC|Estradiol^2nd specimen post XXX challenge|Estradiol^2nd specimen post XXX challenge
C2359799|T201|COMP|51502-3|LNC|Estradiol^6th specimen post XXX challenge|Estradiol^6th specimen post XXX challenge
C2359800|T201|COMP|51503-1|LNC|Penicillin G procaine|Penicillin G procaine
C2359801|T201|COMP|51504-9|LNC|Penicillin G benzathine|Penicillin G benzathine
C2359802|T201|COMP|51505-6|LNC|Creatine kinase.BB|Creatine kinase.BB
C2359807|T201|COMP|51524-7|LNC|Betula verrucosa recombinant (rBet v) 2+4 Ab.IgE|Betula verrucosa recombinant (rBet v) 2+4 Ab.IgE
C2359817|T201|COMP|51530-4|LNC|Lactalbumin alpha Ab.IgG|Lactalbumin alpha Ab.IgG
C2359818|T201|COMP|51531-2|LNC|Beta lactoglobulin Ab.IgG|Beta lactoglobulin Ab.IgG
C2359869|T201|COMP|51498-4|LNC|Estradiol^3rd specimen post XXX challenge|Estradiol^3rd specimen post XXX challenge
C2359870|T201|COMP|51499-2|LNC|Estradiol^1st specimen post XXX challenge|Estradiol^1st specimen post XXX challenge
C2359871|T201|COMP|51500-7|LNC|Estradiol^7th specimen post XXX challenge|Estradiol^7th specimen post XXX challenge
C2359873|T201|COMP|51869-6|LNC|Washed packed erythrocytes given|Washed packed erythrocytes given
C2359875|T201|COMP|51870-4|LNC|Frozen erythrocytes given|Frozen erythrocytes given
C2359877|T201|COMP|51871-2|LNC|Direct antiglobulin test.poly specific reagent|Direct antiglobulin test.poly specific reagent
C2359879|T201|COMP|51872-0|LNC|Transfuse platelet concentrate units|Transfuse platelet concentrate units
C2359881|T201|COMP|51873-8|LNC|Platelet concentrate units given|Platelet concentrate units given
C2359883|T201|COMP|51874-6|LNC|Varicella zoster virus immune globulin ordered|Varicella zoster virus immune globulin ordered
C2359885|T201|COMP|51625-2|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C2359887|T201|COMP|51627-8|LNC|Lymphocytes|Lymphocytes
C2359888|T201|COMP|51628-6|LNC|Morphology|Morphology
C2359889|T201|COMP|51629-4|LNC|Macroblasts/100 cells|Macroblasts/100 cells
C2359891|T201|COMP|51630-2|LNC|Schistocytes/1000 erythrocytes|Schistocytes/1000 erythrocytes
C2359893|T201|COMP|51631-0|LNC|Platelet distribution width|Platelet distribution width
C2359894|T201|COMP|51632-8|LNC|Platelets.reticulated|Platelets.reticulated
C2359896|T201|COMP|51633-6|LNC|Platelets.reticulated/100 platelets|Platelets.reticulated/100 platelets
C2359898|T201|COMP|51634-4|LNC|Reticulocytes.mid|Reticulocytes.mid
C2359899|T201|COMP|51635-1|LNC|Reticulocytes.mature|Reticulocytes.mature
C2359900|T201|COMP|51636-9|LNC|Reticulocytes.immature|Reticulocytes.immature
C2359901|T201|COMP|51637-7|LNC|Plateletocrit|Plateletocrit
C2359903|T201|COMP|51638-5|LNC|Erythrocyte aggregates|Erythrocyte aggregates
C2359905|T201|COMP|51795-3|LNC|Complement C1 esterase inhibitor bound Ab|Complement C1 esterase inhibitor bound Ab
C2359906|T201|COMP|51796-1|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C2359907|T201|COMP|51797-9|LNC|CV2 Ab|CV2 Ab
C2359908|T201|COMP|51798-7|LNC|Hepatitis E virus Ab.IgM|Hepatitis E virus Ab.IgM
C2359909|T201|COMP|51799-5|LNC|Adenosine deaminase|Adenosine deaminase
C2359910|T201|COMP|51800-1|LNC|Homogentisate|Homogentisate
C2359911|T201|COMP|51801-9|LNC|Myeloperoxidase Ab|Myeloperoxidase Ab
C2359912|T201|COMP|51802-7|LNC|Phosphatidylserine Ab.IgM|Phosphatidylserine Ab.IgM
C2359913|T201|COMP|51803-5|LNC|Fibrillarin Ab|Fibrillarin Ab
C2359914|T201|COMP|51804-3|LNC|Rickettsia conorii Ab.IgG|Rickettsia conorii Ab.IgG
C2359915|T201|COMP|51805-0|LNC|Rickettsia conorii Ab.IgM|Rickettsia conorii Ab.IgM
C2359916|T201|COMP|51806-8|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C2359917|T201|COMP|51807-6|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C2359918|T201|COMP|51808-4|LNC|Chlamydophila psittaci Ab.IgG|Chlamydophila psittaci Ab.IgG
C2359983|T201|COMP|53158-2|LNC|Homocitrulline|Homocitrulline
C2359984|T201|COMP|53159-0|LNC|Tryptophan|Tryptophan
C2359985|T201|COMP|53160-8|LNC|Propionylcarnitine (C3)|Propionylcarnitine (C3)
C2359986|T201|COMP|53161-6|LNC|Propionylcarnitine (C3)/Methionine|Propionylcarnitine (C3)/Methionine
C2359988|T201|COMP|53162-4|LNC|Propionylcarnitine (C3)/Carnitine.free (C0)|Propionylcarnitine (C3)/Carnitine.free (C0)
C2359990|T201|COMP|53163-2|LNC|Propionylcarnitine (C3)/Acetylcarnitine (C2)|Propionylcarnitine (C3)/Acetylcarnitine (C2)
C2359992|T201|COMP|53164-0|LNC|Propionylcarnitine (C3)/Palmitoylcarnitine (C16)|Propionylcarnitine (C3)/Palmitoylcarnitine (C16)
C2359994|T201|COMP|53165-7|LNC|Formiminoglutamate|Formiminoglutamate
C2359996|T201|COMP|53166-5|LNC|Butyrylcarnitine+Isobutyrylcarnitine (C4)|Butyrylcarnitine+Isobutyrylcarnitine (C4)
C2360003|T201|COMP|53170-7|LNC|Tiglylcarnitine (C5:1)|Tiglylcarnitine (C5:1)
C2360015|T201|COMP|51932-2|LNC|Saquinavir^trough|Saquinavir^trough
C2360016|T201|COMP|51933-0|LNC|Secale cereale Ab.IgG|Secale cereale Ab.IgG
C2360018|T201|COMP|51935-5|LNC|Trypsinogen I.free|Trypsinogen I.free
C2360019|T201|COMP|51936-3|LNC|Yeast bakers Ab.IgG|Yeast bakers Ab.IgG
C2360020|T201|COMP|51937-1|LNC|HLA-A+B+Bw+DR|HLA-A+B+Bw+DR
C2360022|T201|COMP|51938-9|LNC|HLA-A+B+Bw+DR|HLA-A+B+Bw+DR
C2360023|T201|COMP|51939-7|LNC|Escherichia coli shiga-like toxin 2|Escherichia coli shiga-like toxin 2
C2360070|T201|COMP|51488-5|LNC|Cortisol^6th specimen post XXX challenge|Cortisol^6th specimen post XXX challenge
C2360071|T201|COMP|51489-3|LNC|Cortisol^7th specimen post XXX challenge|Cortisol^7th specimen post XXX challenge
C2360072|T201|COMP|51490-1|LNC|Cortisol^5th specimen post XXX challenge|Cortisol^5th specimen post XXX challenge
C2360073|T201|COMP|51491-9|LNC|Cortisol^4th specimen post XXX challenge|Cortisol^4th specimen post XXX challenge
C2360074|T201|COMP|51492-7|LNC|Cortisol^3rd specimen post XXX challenge|Cortisol^3rd specimen post XXX challenge
C2360075|T201|COMP|51493-5|LNC|Cortisol^2nd specimen post XXX challenge|Cortisol^2nd specimen post XXX challenge
C2360076|T201|COMP|51494-3|LNC|Cortisol^1st specimen post XXX challenge|Cortisol^1st specimen post XXX challenge
C2360077|T201|COMP|51495-0|LNC|Cortisol^baseline|Cortisol^baseline
C2360078|T201|COMP|51496-8|LNC|Estradiol^4th specimen post XXX challenge|Estradiol^4th specimen post XXX challenge
C2360079|T201|COMP|51497-6|LNC|Estradiol^5th specimen post XXX challenge|Estradiol^5th specimen post XXX challenge
C2360080|T201|COMP|51506-4|LNC|Creatine kinase.MB|Creatine kinase.MB
C2360081|T201|COMP|51507-2|LNC|Creatine kinase.MM|Creatine kinase.MM
C2360089|T201|COMP|51901-7|LNC|Avena sativa Ab.IgG|Avena sativa Ab.IgG
C2360090|T201|COMP|51902-5|LNC|Cadmium|Cadmium
C2360091|T201|COMP|51903-3|LNC|Chromium|Chromium
C2360092|T201|COMP|51904-1|LNC|Citrus sinensis Ab.IgG|Citrus sinensis Ab.IgG
C2360093|T201|COMP|51905-8|LNC|Collection end time|Collection end time
C2360094|T201|COMP|51906-6|LNC|Collection start time|Collection start time
C2360095|T201|COMP|51907-4|LNC|Efavirenz^trough|Efavirenz^trough
C2360098|T201|COMP|52124-5|LNC|Osmotic fragility^0.90% sodium chloride|Osmotic fragility^0.90% sodium chloride
C2360100|T201|COMP|52126-0|LNC|Acid glycerol lysis|Acid glycerol lysis
C2360102|T201|COMP|52127-8|LNC|Megaloblasts/100 cells|Megaloblasts/100 cells
C2360104|T201|COMP|52128-6|LNC|Cefotaxime|Cefotaxime
C2360117|T201|COMP|52928-9|LNC|Molybdenum/Creatinine|Molybdenum/Creatinine
C2360118|T201|COMP|52929-7|LNC|Mercury/Creatinine|Mercury/Creatinine
C2360119|T201|COMP|52930-5|LNC|Manganese/Creatinine|Manganese/Creatinine
C2360120|T201|COMP|52931-3|LNC|Lead/Creatinine|Lead/Creatinine
C2360121|T201|COMP|52932-1|LNC|Copper/Creatinine|Copper/Creatinine
C2360122|T201|COMP|52933-9|LNC|Cobalt/Creatinine|Cobalt/Creatinine
C2360123|T201|COMP|52934-7|LNC|Chromium/Creatinine|Chromium/Creatinine
C2360124|T201|COMP|52935-4|LNC|Beryllium/Creatinine|Beryllium/Creatinine
C2360170|T201|COMP|51532-0|LNC|Casein Ab.IgG|Casein Ab.IgG
C2360171|T201|COMP|51533-8|LNC|Dermatophagoides pteronyssinus Ab.IgG|Dermatophagoides pteronyssinus Ab.IgG
C2360172|T201|COMP|51534-6|LNC|Dermatophagoides farinae Ab.IgG|Dermatophagoides farinae Ab.IgG
C2360173|T201|COMP|51535-3|LNC|Phleum pratense Ab.IgG|Phleum pratense Ab.IgG
C2360174|T201|COMP|51536-1|LNC|Egg white Ab.IgG|Egg white Ab.IgG
C2360175|T201|COMP|51537-9|LNC|Betula verrucosa Ab.IgG|Betula verrucosa Ab.IgG
C2360176|T201|COMP|51538-7|LNC|Cladosporium herbarum Ab.IgG|Cladosporium herbarum Ab.IgG
C2360177|T201|COMP|51539-5|LNC|Candida albicans Ab.IgG|Candida albicans Ab.IgG
C2360178|T201|COMP|51540-3|LNC|Alternaria alternata Ab.IgG|Alternaria alternata Ab.IgG
C2360179|T201|COMP|51541-1|LNC|Stachybotrys chartarum Ab.IgG|Stachybotrys chartarum Ab.IgG
C2360180|T201|COMP|51542-9|LNC|Aspergillus versicolor Ab.IgG|Aspergillus versicolor Ab.IgG
C2360181|T201|COMP|51543-7|LNC|Cladosporium cladosporioides Ab.IgG|Cladosporium cladosporioides Ab.IgG
C2360182|T201|COMP|51544-5|LNC|Penicillium sp Ab.IgG|Penicillium sp Ab.IgG
C2360183|T201|COMP|51545-2|LNC|Budgerigar droppings Ab.IgG|Budgerigar droppings Ab.IgG
C2360185|T201|COMP|51546-0|LNC|Chicken feather Ab.IgG|Chicken feather Ab.IgG
C2360186|T201|COMP|51547-8|LNC|Canary feather Ab.IgG|Canary feather Ab.IgG
C2360188|T201|COMP|51548-6|LNC|Parrot feather Ab.IgG|Parrot feather Ab.IgG
C2360190|T201|COMP|51549-4|LNC|Pigeon feather Ab.IgG|Pigeon feather Ab.IgG
C2360194|T201|COMP|51551-0|LNC|Chinchilla epithelium Ab.IgE.RAST class|Chinchilla epithelium Ab.IgE.RAST class
C2360196|T201|COMP|51552-8|LNC|Fox epithelium Ab.IgE.RAST class|Fox epithelium Ab.IgE.RAST class
C2360198|T201|COMP|51553-6|LNC|Mace Ab.IgE.RAST class|Mace Ab.IgE.RAST class
C2360200|T201|COMP|51554-4|LNC|Merluccius merluccius Ab.IgE.RAST class|Merluccius merluccius Ab.IgE.RAST class
C2360222|T201|COMP|51565-0|LNC|Ficus sp Ab.IgE.RAST class|Ficus sp Ab.IgE.RAST class
C2360224|T201|COMP|51566-8|LNC|Amylase Ab.IgE.RAST class|Amylase Ab.IgE.RAST class
C2360226|T201|COMP|51567-6|LNC|Trichosporon pullulans Ab.IgE.RAST class|Trichosporon pullulans Ab.IgE.RAST class
C2360246|T201|COMP|51577-5|LNC|Elaeis guineensis Ab.IgE.RAST class|Elaeis guineensis Ab.IgE.RAST class
C2360248|T201|COMP|51578-3|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C2360249|T201|COMP|51579-1|LNC|Normoblasts/100 cells|Normoblasts/100 cells
C2360251|T201|COMP|51580-9|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C2360252|T201|COMP|51581-7|LNC|Other cells/100 cells|Other cells/100 cells
C2360254|T201|COMP|51582-5|LNC|Anisochromasia|Anisochromasia
C2360255|T201|COMP|51583-3|LNC|Anulocytes|Anulocytes
C2360257|T201|COMP|51584-1|LNC|Granulocytes.immature|Granulocytes.immature
C2360258|T201|COMP|51585-8|LNC|Other cells|Other cells
C2360259|T201|COMP|51586-6|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C2360260|T201|COMP|51587-4|LNC|Plasmodium sp|Plasmodium sp
C2360261|T201|COMP|51588-2|LNC|Granulocytes|Granulocytes
C2360262|T201|COMP|51589-0|LNC|Dyserythropoiesis|Dyserythropoiesis
C2360263|T201|COMP|51590-8|LNC|Chloride|Chloride
C2360264|T201|COMP|51591-6|LNC|Cholesterol|Cholesterol
C2360265|T201|COMP|51592-4|LNC|Creatinine|Creatinine
C2360266|T201|COMP|51593-2|LNC|Fructose|Fructose
C2360267|T201|COMP|51594-0|LNC|Galactose|Galactose
C2360268|T201|COMP|51595-7|LNC|Glucose|Glucose
C2360269|T201|COMP|51596-5|LNC|Glucose|Glucose
C2360270|T201|COMP|51597-3|LNC|Glucose^1H post 75 g glucose PO|Glucose^1H post 75 g glucose PO
C2360271|T201|COMP|51598-1|LNC|Lactose|Lactose
C2360272|T201|COMP|51599-9|LNC|Methotrexate^12H post dose|Methotrexate^12H post dose
C2360273|T201|COMP|51600-5|LNC|Methotrexate^24H post dose|Methotrexate^24H post dose
C2360274|T201|COMP|51601-3|LNC|Methotrexate^4H post dose|Methotrexate^4H post dose
C2360275|T201|COMP|51602-1|LNC|Methotrexate^72H post dose|Methotrexate^72H post dose
C2360276|T201|COMP|51603-9|LNC|Cytochrome b5 reductase|Cytochrome b5 reductase
C2360277|T201|COMP|51604-7|LNC|Phosphate|Phosphate
C2360278|T201|COMP|51605-4|LNC|Triglyceride|Triglyceride
C2360279|T201|COMP|51606-2|LNC|Xylose^3H post dose xylose PO|Xylose^3H post dose xylose PO
C2360280|T201|COMP|51607-0|LNC|Xylose^3H post XXX challenge|Xylose^3H post XXX challenge
C2360281|T201|COMP|51608-8|LNC|Xylose^30M post dose xylose PO|Xylose^30M post dose xylose PO
C2360282|T201|COMP|51609-6|LNC|Xylose^30M post XXX challenge|Xylose^30M post XXX challenge
C2360283|T201|COMP|51610-4|LNC|Calcium|Calcium
C2360284|T201|COMP|51611-2|LNC|Methotrexate^48H post dose|Methotrexate^48H post dose
C2360285|T201|COMP|51612-0|LNC|Sucrose|Sucrose
C2360286|T201|COMP|51613-8|LNC|Hemoglobin J/Hemoglobin.total|Hemoglobin J/Hemoglobin.total
C2360288|T201|COMP|51614-6|LNC|Hemoglobin M/Hemoglobin.total|Hemoglobin M/Hemoglobin.total
C2360290|T201|COMP|51615-3|LNC|Hemoglobin A2+C/Hemoglobin.total|Hemoglobin A2+C/Hemoglobin.total
C2360292|T201|COMP|51616-1|LNC|Hemoglobin A2+E/Hemoglobin.total|Hemoglobin A2+E/Hemoglobin.total
C2360294|T201|COMP|51617-9|LNC|Color|Color
C2360295|T201|COMP|51618-7|LNC|Potassium^pre dialysis|Potassium^pre dialysis
C2360296|T201|COMP|51619-5|LNC|Creatinine^pre dialysis|Creatinine^pre dialysis
C2360297|T201|COMP|51620-3|LNC|Creatinine^post dialysis|Creatinine^post dialysis
C2360298|T201|COMP|51621-1|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C2360299|T201|COMP|51622-9|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C2360300|T201|COMP|51623-7|LNC|Spermatozoa^post vasectomy|Spermatozoa^post vasectomy
C2360301|T201|COMP|51624-5|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C2360302|T201|COMP|51639-3|LNC|Acanthocytes/1000 erythrocytes|Acanthocytes/1000 erythrocytes
C2360304|T201|COMP|51640-1|LNC|Platelet anisocytosis|Platelet anisocytosis
C2360305|T201|COMP|51641-9|LNC|Mean sphered cell volume|Mean sphered cell volume
C2360309|T201|COMP|51643-5|LNC|Reticulocytes.high light scatter|Reticulocytes.high light scatter
C2360311|T201|COMP|51644-3|LNC|Megakaryocytic nuclei|Megakaryocytic nuclei
C2360313|T201|COMP|51645-0|LNC|Micromegakaryocytes|Micromegakaryocytes
C2360314|T201|COMP|51646-8|LNC|Rabies virus RNA|Rabies virus RNA
C2360316|T201|COMP|51647-6|LNC|Rabies virus RNA|Rabies virus RNA
C2360317|T201|COMP|51648-4|LNC|Monocytoid cells/100 leukocytes|Monocytoid cells/100 leukocytes
C2360319|T201|COMP|51649-2|LNC|Hepatitis C virus c100p+5-1-1 Ab|Hepatitis C virus c100p+5-1-1 Ab
C2360320|T201|COMP|51650-0|LNC|HLA-B|HLA-B
C2360321|T201|COMP|51651-8|LNC|IgE Ab|IgE Ab
C2360322|T201|COMP|51652-6|LNC|SLC14A1 gene targeted mutation analysis|SLC14A1 gene targeted mutation analysis
C2360324|T201|COMP|51653-4|LNC|Hepatitis E virus Ab|Hepatitis E virus Ab
C2360325|T201|COMP|51654-2|LNC|Hepatitis D virus Ab|Hepatitis D virus Ab
C2360326|T201|COMP|51655-9|LNC|Hepatitis C virus RNA|Hepatitis C virus RNA
C2360327|T201|COMP|51656-7|LNC|Hepatitis C virus Ab Signal/Cutoff|Hepatitis C virus Ab Signal/Cutoff
C2360328|T201|COMP|51657-5|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C2360329|T201|COMP|51658-3|LNC|Hepatitis B virus core Ab.IgM|Hepatitis B virus core Ab.IgM
C2360330|T201|COMP|51659-1|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C2360331|T201|COMP|51660-9|LNC|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C2360332|T201|COMP|51661-7|LNC|Hepatitis A virus Ab|Hepatitis A virus Ab
C2360333|T201|COMP|51662-5|LNC|Core respiratory allergens panel|Core respiratory allergens panel
C2360335|T201|COMP|51663-3|LNC|Alphavirus RNA|Alphavirus RNA
C2360337|T201|COMP|51664-1|LNC|Chikungunya virus RNA|Chikungunya virus RNA
C2360339|T201|COMP|51665-8|LNC|Flavivirus RNA|Flavivirus RNA
C2360341|T201|COMP|51666-6|LNC|Japanese encephalitis virus RNA|Japanese encephalitis virus RNA
C2360342|T201|COMP|51667-4|LNC|Lymphocytic choriomeningitis virus RNA|Lymphocytic choriomeningitis virus RNA
C2360346|T201|COMP|51669-0|LNC|Parechovirus A RNA|Parechovirus A RNA
C2360348|T201|COMP|51670-8|LNC|17-Hydroxypregnenolone^baseline|17-Hydroxypregnenolone^baseline
C2360349|T201|COMP|51671-6|LNC|Brucella sp Ab|Brucella sp Ab
C2360360|T201|COMP|51682-3|LNC|Pregnenolone^3rd specimen post XXX challenge|Pregnenolone^3rd specimen post XXX challenge
C2360361|T201|COMP|51683-1|LNC|Pregnenolone^baseline|Pregnenolone^baseline
C2360362|T201|COMP|51684-9|LNC|Pregnenolone^6th specimen post XXX challenge|Pregnenolone^6th specimen post XXX challenge
C2360363|T201|COMP|51685-6|LNC|Pregnenolone^1st specimen post XXX challenge|Pregnenolone^1st specimen post XXX challenge
C2360364|T201|COMP|51686-4|LNC|Pregnenolone^2nd specimen post XXX challenge|Pregnenolone^2nd specimen post XXX challenge
C2360365|T201|COMP|51687-2|LNC|Pregnenolone^7th specimen post XXX challenge|Pregnenolone^7th specimen post XXX challenge
C2360366|T201|COMP|51688-0|LNC|Pregnenolone^4th specimen post XXX challenge|Pregnenolone^4th specimen post XXX challenge
C2360367|T201|COMP|51689-8|LNC|Pregnenolone^5th specimen post XXX challenge|Pregnenolone^5th specimen post XXX challenge
C2360368|T201|COMP|51690-6|LNC|Amphetamines|Amphetamines
C2360369|T201|COMP|51691-4|LNC|Opiates|Opiates
C2360370|T201|COMP|51692-2|LNC|Phencyclidine|Phencyclidine
C2360371|T201|COMP|51693-0|LNC|Albumin|Albumin
C2360372|T201|COMP|51694-8|LNC|Carumonam|Carumonam
C2360373|T201|COMP|51695-5|LNC|Chloride|Chloride
C2360374|T201|COMP|51696-3|LNC|Corticotropin^afternoon specimen|Corticotropin^afternoon specimen
C2360375|T201|COMP|51697-1|LNC|CV2 Ab|CV2 Ab
C2360376|T201|COMP|51698-9|LNC|Dapsone|Dapsone
C2360377|T201|COMP|51699-7|LNC|Endomysium Ab.IgG|Endomysium Ab.IgG
C2360379|T201|COMP|51701-1|LNC|Ganglioside Ab.IgG|Ganglioside Ab.IgG
C2360381|T201|COMP|51702-9|LNC|Ganglioside Ab.IgM|Ganglioside Ab.IgM
C2360383|T201|COMP|51703-7|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C2360384|T201|COMP|51704-5|LNC|Herpes virus 6 Ab|Herpes virus 6 Ab
C2360385|T201|COMP|51705-2|LNC|Homogentisate|Homogentisate
C2360386|T201|COMP|51706-0|LNC|Hyaluronate|Hyaluronate
C2360387|T201|COMP|51707-8|LNC|Inner Ear 68kD Ab|Inner Ear 68kD Ab
C2360388|T201|COMP|51708-6|LNC|Intercellular substance Ab|Intercellular substance Ab
C2360389|T201|COMP|51709-4|LNC|Leishmania sp identified|Leishmania sp identified
C2360390|T201|COMP|51710-2|LNC|Leishmania sp identified|Leishmania sp identified
C2360391|T201|COMP|51711-0|LNC|Leishmania sp Ab|Leishmania sp Ab
C2360392|T201|COMP|51712-8|LNC|Ma+Ta Ab|Ma+Ta Ab
C2360393|T201|COMP|51713-6|LNC|Metamyelocytes/100 leukocytes|Metamyelocytes/100 leukocytes
C2360395|T201|COMP|51715-1|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C2360396|T201|COMP|51716-9|LNC|Muscle specific receptor tyrosine kinase Ab|Muscle specific receptor tyrosine kinase Ab
C2360397|T201|COMP|51717-7|LNC|Normoblasts.orthochromic/100 cells|Normoblasts.orthochromic/100 cells
C2360398|T201|COMP|51718-5|LNC|Normoblasts.polychromatophilic/100 cells|Normoblasts.polychromatophilic/100 cells
C2360399|T201|COMP|51719-3|LNC|Paromomycin|Paromomycin
C2360400|T201|COMP|51720-1|LNC|Potassium|Potassium
C2360401|T201|COMP|51721-9|LNC|Purkinje cells Ab|Purkinje cells Ab
C2360402|T201|COMP|51722-7|LNC|Reticulin Ab|Reticulin Ab
C2360403|T201|COMP|51723-5|LNC|Fungus|Fungus
C2360404|T201|COMP|51724-3|LNC|Cefuroxime|Cefuroxime
C2360412|T201|COMP|51729-2|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C2360413|T201|COMP|51730-0|LNC|Herpes virus 6 Ab.IgG & IgM|Herpes virus 6 Ab.IgG & IgM
C2360414|T201|COMP|51731-8|LNC|Oxygen saturation|Oxygen saturation
C2360415|T201|COMP|51732-6|LNC|Oxygen saturation|Oxygen saturation
C2360416|T201|COMP|51733-4|LNC|Oxygen saturation|Oxygen saturation
C2360417|T201|COMP|51734-2|LNC|Chlamydia trachomatis L2 Ab.IgA & IgG & IgM|Chlamydia trachomatis L2 Ab.IgA & IgG & IgM
C2360419|T201|COMP|51735-9|LNC|Urea nitrogen renal clearance|Urea nitrogen renal clearance
C2360420|T201|COMP|51736-7|LNC|oxyMORphone.free|oxyMORphone.free
C2360421|T201|COMP|51737-5|LNC|HYDROmorphone.free|HYDROmorphone.free
C2360422|T201|COMP|51738-3|LNC|HYDROcodone.free|HYDROcodone.free
C2360423|T201|COMP|51739-1|LNC|Codeine.free|Codeine.free
C2360424|T201|COMP|51740-9|LNC|6-Monoacetylmorphine.free|6-Monoacetylmorphine.free
C2360425|T201|COMP|51741-7|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C2360426|T201|COMP|51742-5|LNC|Borrelia burgdorferi 49736 Ab.IgM|Borrelia burgdorferi 49736 Ab.IgM
C2360428|T201|COMP|51743-3|LNC|Borrelia burgdorferi 49736 Ab.IgG|Borrelia burgdorferi 49736 Ab.IgG
C2360430|T201|COMP|51744-1|LNC|Borrelia burgdorferi 49736 Ab.IgA|Borrelia burgdorferi 49736 Ab.IgA
C2360432|T201|COMP|51745-8|LNC|Borrelia burgdorferi G39_40 Ab.IgG|Borrelia burgdorferi G39_40 Ab.IgG
C2360434|T201|COMP|51746-6|LNC|Borrelia burgdorferi 49736 Ab.IgG|Borrelia burgdorferi 49736 Ab.IgG
C2360435|T201|COMP|51747-4|LNC|Borrelia burgdorferi Ab.IgA & IgG & IgM|Borrelia burgdorferi Ab.IgA & IgG & IgM
C2360437|T201|COMP|51748-2|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C2360438|T201|COMP|51749-0|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C2360439|T201|COMP|51750-8|LNC|Pyruvate|Pyruvate
C2360440|T201|COMP|51751-6|LNC|Pyruvate|Pyruvate
C2360443|T201|COMP|51753-2|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C2360444|T201|COMP|51754-0|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C2360445|T201|COMP|51755-7|LNC|Cells.CD3+CD4-CD8-CD45+/100 cells|Cells.CD3+CD4-CD8-CD45+/100 cells
C2360447|T201|COMP|51756-5|LNC|ATP7B gene targeted mutation analysis|ATP7B gene targeted mutation analysis
C2360448|T201|COMP|51757-3|LNC|POMT1 gene targeted mutation analysis|POMT1 gene targeted mutation analysis
C2360450|T201|COMP|51758-1|LNC|POMT2 gene targeted mutation analysis|POMT2 gene targeted mutation analysis
C2360452|T201|COMP|51759-9|LNC|RAI1 gene targeted mutation analysis|RAI1 gene targeted mutation analysis
C2360454|T201|COMP|51760-7|LNC|Ehrlichia chaffeensis Ab.IgG+IgM|Ehrlichia chaffeensis Ab.IgG+IgM
C2360456|T201|COMP|51761-5|LNC|Giardia lamblia Ab.IgA & IgG & IgM|Giardia lamblia Ab.IgA & IgG & IgM
C2360458|T201|COMP|51762-3|LNC|Helicobacter pylori Ab.IgA & IgG & IgM|Helicobacter pylori Ab.IgA & IgG & IgM
C2360460|T201|COMP|51763-1|LNC|Muscle specific receptor tyrosine kinase Ab|Muscle specific receptor tyrosine kinase Ab
C2360461|T201|COMP|51764-9|LNC|Trypanosoma cruzi Ab.IgG & IgM|Trypanosoma cruzi Ab.IgG & IgM
C2360463|T201|COMP|51765-6|LNC|Dihydrocodeine+Hydrocodol|Dihydrocodeine+Hydrocodol
C2360464|T201|COMP|51766-4|LNC|Glucose^2.5H post dose fructose PO|Glucose^2.5H post dose fructose PO
C2360465|T201|COMP|51767-2|LNC|Glucose^1.5H post dose fructose PO|Glucose^1.5H post dose fructose PO
C2360466|T201|COMP|51768-0|LNC|Glucose^3H post dose fructose PO|Glucose^3H post dose fructose PO
C2360467|T201|COMP|51769-8|LNC|Glucose^2H post dose fructose PO|Glucose^2H post dose fructose PO
C2360468|T201|COMP|51770-6|LNC|Leukocytes|Leukocytes
C2360469|T201|COMP|51771-4|LNC|Histoplasma capsulatum DNA|Histoplasma capsulatum DNA
C2360470|T201|COMP|51772-2|LNC|F9 gene mutations tested for|F9 gene mutations tested for
C2360472|T201|COMP|51773-0|LNC|HEXA gene targeted mutation analysis|HEXA gene targeted mutation analysis
C2360473|T201|COMP|51774-8|LNC|Cefuroxime|Cefuroxime
C2360474|T201|COMP|51775-5|LNC|Chromatin Ab|Chromatin Ab
C2360475|T201|COMP|51776-3|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2360476|T201|COMP|51777-1|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C2360477|T201|COMP|51778-9|LNC|YY1 gene targeted mutation analysis|YY1 gene targeted mutation analysis
C2360479|T201|COMP|51779-7|LNC|CFH gene targeted mutation analysis|CFH gene targeted mutation analysis
C2360481|T201|COMP|51780-5|LNC|HIV 1 RNA|HIV 1 RNA
C2360482|T201|COMP|51781-3|LNC|Carbon dioxide|Carbon dioxide
C2360483|T201|COMP|51782-1|LNC|Drugs of abuse 7 & Alcohol & Tricyclics panel|Drugs of abuse 7 & Alcohol & Tricyclics panel
C2360485|T201|COMP|51783-9|LNC|Reagin Ab|Reagin Ab
C2360486|T201|COMP|51784-7|LNC|Lot number|Lot number
C2360487|T201|COMP|51785-4|LNC|Dengue virus Ab.IgG & IgM|Dengue virus Ab.IgG & IgM
C2360489|T201|COMP|51786-2|LNC|HIV 2 Ab Signal/Cutoff|HIV 2 Ab Signal/Cutoff
C2360491|T201|COMP|51787-0|LNC|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C2360492|T201|COMP|51788-8|LNC|Coccidioides sp Ab|Coccidioides sp Ab
C2360493|T201|COMP|51789-6|LNC|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C2360494|T201|COMP|51790-4|LNC|Erythrocyte casts|Erythrocyte casts
C2360495|T201|COMP|51791-2|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C2360496|T201|COMP|51792-0|LNC|Citrate/Creatinine|Citrate/Creatinine
C2360497|T201|COMP|51793-8|LNC|Xylose^1H post 5 g xylose PO|Xylose^1H post 5 g xylose PO
C2360498|T201|COMP|51794-6|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C2360499|T201|COMP|51809-2|LNC|Chlamydophila psittaci Ab.IgM|Chlamydophila psittaci Ab.IgM
C2360500|T201|COMP|51810-0|LNC|Coxiella burnetii phase 1 Ab.IgG|Coxiella burnetii phase 1 Ab.IgG
C2360501|T201|COMP|51811-8|LNC|Coxiella burnetii phase 1 Ab.IgM|Coxiella burnetii phase 1 Ab.IgM
C2360502|T201|COMP|51812-6|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C2360503|T201|COMP|51813-4|LNC|Coxiella burnetii phase 2 Ab.IgM|Coxiella burnetii phase 2 Ab.IgM
C2360504|T201|COMP|51814-2|LNC|Legionella pneumophila Ab.IgM|Legionella pneumophila Ab.IgM
C2360505|T201|COMP|51815-9|LNC|Leptospira sp Ab.IgG|Leptospira sp Ab.IgG
C2360506|T201|COMP|51816-7|LNC|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C2360507|T201|COMP|51817-5|LNC|Coxsackievirus B Ab.IgG|Coxsackievirus B Ab.IgG
C2360508|T201|COMP|51818-3|LNC|Coxsackievirus B Ab.IgM|Coxsackievirus B Ab.IgM
C2360509|T201|COMP|51819-1|LNC|Leptospira sp Ab.IgM|Leptospira sp Ab.IgM
C2360510|T201|COMP|51820-9|LNC|Listeria monocytogenes Ab.IgG|Listeria monocytogenes Ab.IgG
C2360511|T201|COMP|51821-7|LNC|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C2360512|T201|COMP|51822-5|LNC|Adenovirus Ab.IgG|Adenovirus Ab.IgG
C2360513|T201|COMP|51823-3|LNC|Adenovirus Ab.IgM|Adenovirus Ab.IgM
C2360514|T201|COMP|51824-1|LNC|Hepatitis C virus Ab.IgM|Hepatitis C virus Ab.IgM
C2360516|T201|COMP|51825-8|LNC|Bordetella parapertussis Ab|Bordetella parapertussis Ab
C2360517|T201|COMP|51826-6|LNC|Herpes virus 8 Ab.IgG|Herpes virus 8 Ab.IgG
C2360518|T201|COMP|51827-4|LNC|Trypanosoma cruzi Ab.IgM|Trypanosoma cruzi Ab.IgM
C2360520|T201|COMP|51829-0|LNC|Lactate|Lactate
C2360521|T201|COMP|51830-8|LNC|Prolymphocytes/100 leukocytes|Prolymphocytes/100 leukocytes
C2360522|T201|COMP|51831-6|LNC|Beta-2 transferrin|Beta-2 transferrin
C2360523|T201|COMP|51832-4|LNC|Brucella abortus Ab|Brucella abortus Ab
C2360524|T201|COMP|51833-2|LNC|14-3-3 protein|14-3-3 protein
C2360525|T201|COMP|51834-0|LNC|Tryptase|Tryptase
C2360526|T201|COMP|51835-7|LNC|Angiotensin converting enzyme|Angiotensin converting enzyme
C2360527|T201|COMP|51836-5|LNC|Angiotensin II^upright|Angiotensin II^upright
C2360528|T201|COMP|51837-3|LNC|Bordetella parapertussis Ab.IgG|Bordetella parapertussis Ab.IgG
C2360530|T201|COMP|51838-1|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C2360531|T201|COMP|51839-9|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C2360532|T201|COMP|51840-7|LNC|Echovirus Ab.IgG|Echovirus Ab.IgG
C2360534|T201|COMP|51841-5|LNC|Echovirus Ab.IgM|Echovirus Ab.IgM
C2360536|T201|COMP|51842-3|LNC|Plasmodium falciparum Ab.IgM|Plasmodium falciparum Ab.IgM
C2360538|T201|COMP|51843-1|LNC|Malonate/Creatinine|Malonate/Creatinine
C2360539|T201|COMP|51844-9|LNC|Cortisol|Cortisol
C2360555|T201|COMP|51856-3|LNC|Staphylococcus aureus TSST-1 Ab.IgE|Staphylococcus aureus TSST-1 Ab.IgE
C2360557|T201|COMP|51857-1|LNC|Malassezia sp Ab.IgE|Malassezia sp Ab.IgE
C2360561|T201|COMP|51859-7|LNC|Pigeon serum proteins+feathers+droppings Ab.IgG|Pigeon serum proteins+feathers+droppings Ab.IgG
C2360563|T201|COMP|51860-5|LNC|Parrot serum proteins+feathers+droppings Ab.IgG|Parrot serum proteins+feathers+droppings Ab.IgG
C2360569|T201|COMP|51863-9|LNC|Staphylococcus aureus TSST-1 Ab.IgE.RAST class|Staphylococcus aureus TSST-1 Ab.IgE.RAST class
C2360571|T201|COMP|51864-7|LNC|Malassezia sp Ab.IgE.RAST class|Malassezia sp Ab.IgE.RAST class
C2360573|T201|COMP|51865-4|LNC|Plasmodium sp Ag|Plasmodium sp Ag
C2360574|T201|COMP|51866-2|LNC|HIV 1 Ab+Ag|HIV 1 Ab+Ag
C2360576|T201|COMP|51867-0|LNC|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript
C2360578|T201|COMP|51876-1|LNC|Whole blood units given|Whole blood units given
C2360579|T201|COMP|51877-9|LNC|Transfuse fresh frozen plasma units|Transfuse fresh frozen plasma units
C2360581|T201|COMP|51878-7|LNC|Fresh frozen plasma units given|Fresh frozen plasma units given
C2360582|T201|COMP|51879-5|LNC|Transfuse packed erythrocytes units|Transfuse packed erythrocytes units
C2360584|T201|COMP|51880-3|LNC|Packed erythrocytes units given|Packed erythrocytes units given
C2360585|T201|COMP|51881-1|LNC|Transfuse cryoprecipitate units|Transfuse cryoprecipitate units
C2360586|T201|COMP|51882-9|LNC|Cryoprecipitate units given|Cryoprecipitate units given
C2360587|T201|COMP|51883-7|LNC|Transfuse whole blood units|Transfuse whole blood units
C2360588|T201|COMP|51884-5|LNC|Transfuse pooled platelets units|Transfuse pooled platelets units
C2360590|T201|COMP|51885-2|LNC|Transfuse whole blood autologous units|Transfuse whole blood autologous units
C2360591|T201|COMP|51886-0|LNC|Autologous whole blood units given|Autologous whole blood units given
C2360592|T201|COMP|51887-8|LNC|Transfuse Rh immune globulin units|Transfuse Rh immune globulin units
C2360593|T201|COMP|51888-6|LNC|Rh immune globulin units given|Rh immune globulin units given
C2360594|T201|COMP|51889-4|LNC|Transfuse factor VIII units|Transfuse factor VIII units
C2360652|T201|COMP|51890-2|LNC|Factor VIII units given|Factor VIII units given
C2360653|T201|COMP|51891-0|LNC|Transfuse factor IX units|Transfuse factor IX units
C2360654|T201|COMP|51892-8|LNC|ABO group|ABO group
C2360655|T201|COMP|51893-6|LNC|Transfuse cryoprecipitate poor plasma units|Transfuse cryoprecipitate poor plasma units
C2360656|T201|COMP|51894-4|LNC|Fresh frozen plasma given|Fresh frozen plasma given
C2360657|T201|COMP|51895-1|LNC|Lot number|Lot number
C2360663|T201|COMP|51908-2|LNC|Efavirenz^peak|Efavirenz^peak
C2360664|T201|COMP|51909-0|LNC|Ependymal cells/100 cells|Ependymal cells/100 cells
C2360666|T201|COMP|51910-8|LNC|Erythrocytes|Erythrocytes
C2360669|T201|COMP|51913-2|LNC|Hepatitis A virus Ab.IgG+IgM|Hepatitis A virus Ab.IgG+IgM
C2360671|T201|COMP|51914-0|LNC|Hepatitis B virus core Ab.IgG+IgM|Hepatitis B virus core Ab.IgG+IgM
C2360673|T201|COMP|51915-7|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C2360674|T201|COMP|51916-5|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C2360675|T201|COMP|51917-3|LNC|Hordeum vulgare Ab.IgG|Hordeum vulgare Ab.IgG
C2360676|T201|COMP|51918-1|LNC|Indinavir^trough|Indinavir^trough
C2360677|T201|COMP|51919-9|LNC|Lactuca sativa Ab.IgG|Lactuca sativa Ab.IgG
C2360678|T201|COMP|51920-7|LNC|Legionella sp Ab^2nd specimen|Legionella sp Ab^2nd specimen
C2360679|T201|COMP|51921-5|LNC|Lopinavir^trough|Lopinavir^trough
C2360680|T201|COMP|51922-3|LNC|Malt Ab.IgG|Malt Ab.IgG
C2360681|T201|COMP|51923-1|LNC|Nelfinavir^peak|Nelfinavir^peak
C2360682|T201|COMP|51924-9|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C2360683|T201|COMP|51925-6|LNC|Nevirapine^peak|Nevirapine^peak
C2360684|T201|COMP|51926-4|LNC|Nucleated cells|Nucleated cells
C2360685|T201|COMP|51927-2|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C2360686|T201|COMP|51928-0|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C2360687|T201|COMP|51929-8|LNC|Ritonavir^peak|Ritonavir^peak
C2360688|T201|COMP|51930-6|LNC|Ritonavir^trough|Ritonavir^trough
C2360689|T201|COMP|51931-4|LNC|Rubella virus Ab|Rubella virus Ab
C2360690|T201|COMP|51940-5|LNC|Escherichia coli shiga-like toxin 1|Escherichia coli shiga-like toxin 1
C2360708|T201|COMP|51949-6|LNC|History of trisomy 21|History of trisomy 21
C2360709|T201|COMP|51950-4|LNC|Calcium^post dialysis|Calcium^post dialysis
C2360710|T201|COMP|51951-2|LNC|UGT1A1 gene allele 1|UGT1A1 gene allele 1
C2360712|T201|COMP|51952-0|LNC|UGT1A1 gene allele 2|UGT1A1 gene allele 2
C2360714|T201|COMP|51953-8|LNC|Collection date|Collection date
C2360715|T201|COMP|51954-6|LNC|oxyCODONE.free|oxyCODONE.free
C2360716|T201|COMP|51955-3|LNC|Dihydrocodeine.free+Hydrocodol.free|Dihydrocodeine.free+Hydrocodol.free
C2360717|T201|COMP|51956-1|LNC|DNA region analysis test coverage panel|DNA region analysis test coverage panel
C2360719|T201|COMP|51957-9|LNC|Placer DNA analysis test identifier|Placer DNA analysis test identifier
C2360721|T201|COMP|51958-7|LNC|Transcript reference sequence identifier|Transcript reference sequence identifier
C2360723|T201|COMP|51959-5|LNC|DNA region of interest|DNA region of interest
C2360725|T201|COMP|51960-3|LNC|DNA marker results panel|DNA marker results panel
C2360727|T201|COMP|51961-1|LNC|Drug efficacy sequence variation interpretation|Drug efficacy sequence variation interpretation
C2360729|T201|COMP|51962-9|LNC|Pharmacogenetic DNA analysis panel|Pharmacogenetic DNA analysis panel
C2360731|T201|COMP|51963-7|LNC|Medication assessed|Medication assessed
C2360733|T201|COMP|51964-5|LNC|Drug efficacy analysis overall interpretation|Drug efficacy analysis overall interpretation
C2360735|T201|COMP|51965-2|LNC|Pharmacogenetic analysis report|Pharmacogenetic analysis report
C2360737|T201|COMP|51966-0|LNC|Genetic disease DNA analysis panel|Genetic disease DNA analysis panel
C2360739|T201|COMP|51967-8|LNC|Genetic disease assessed|Genetic disease assessed
C2360741|T201|COMP|51968-6|LNC|Genetic disease analysis overall interpretation|Genetic disease analysis overall interpretation
C2360743|T201|COMP|51969-4|LNC|Genetic analysis summary report|Genetic analysis summary report
C2360745|T201|COMP|51970-2|LNC|Individual allele identifier|Individual allele identifier
C2360747|T201|COMP|51971-0|LNC|Gene product metabolic activity interpretation|Gene product metabolic activity interpretation
C2360749|T201|COMP|51972-8|LNC|Gas panel|Gas panel
C2360750|T201|COMP|51973-6|LNC|Gas panel|Gas panel
C2360751|T201|COMP|51974-4|LNC|Gas panel|Gas panel
C2360752|T201|COMP|51975-1|LNC|Individual allele results panel|Individual allele results panel
C2360754|T201|COMP|51976-9|LNC|Bacillus anthracis capsule Ag|Bacillus anthracis capsule Ag
C2360756|T201|COMP|51977-7|LNC|Chromium|Chromium
C2360757|T201|COMP|51978-5|LNC|Coxsackievirus A Ab|Coxsackievirus A Ab
C2360758|T201|COMP|51979-3|LNC|Donepezil|Donepezil
C2360759|T201|COMP|51980-1|LNC|Glomerular basement membrane Ab|Glomerular basement membrane Ab
C2360760|T201|COMP|51981-9|LNC|HER2|HER2
C2360761|T201|COMP|51982-7|LNC|lamoTRIgine|lamoTRIgine
C2360762|T201|COMP|51983-5|LNC|Levodopa|Levodopa
C2360763|T201|COMP|51984-3|LNC|Meperidine+Normeperidine|Meperidine+Normeperidine
C2360765|T201|COMP|51985-0|LNC|Modafinil|Modafinil
C2360766|T201|COMP|51986-8|LNC|niCARdipine|niCARdipine
C2360767|T201|COMP|51987-6|LNC|Ubiquinone 10|Ubiquinone 10
C2360768|T201|COMP|51988-4|LNC|Ureaplasma urealyticum DNA|Ureaplasma urealyticum DNA
C2360770|T201|COMP|51989-2|LNC|Vasoactive intestinal peptide|Vasoactive intestinal peptide
C2360771|T201|COMP|51990-0|LNC|Basic metabolic panel|Basic metabolic panel
C2360772|T201|COMP|51991-8|LNC|Reference lab test panel|Reference lab test panel
C2360774|T201|COMP|51992-6|LNC|Heavy metals panel|Heavy metals panel
C2360775|T201|COMP|51993-4|LNC|Metanephrine & Normetanephrine panel|Metanephrine & Normetanephrine panel
C2360776|T201|COMP|51994-2|LNC|Homovanillate/Creatinine|Homovanillate/Creatinine
C2360857|T201|COMP|52107-0|LNC|Bacterial capsule|Bacterial capsule
C2360858|T201|COMP|52108-8|LNC|C little o super little b Ab|C little o super little b Ab
C2360860|T201|COMP|52109-6|LNC|C little o super little a Ab|C little o super little a Ab
C2360862|T201|COMP|52110-4|LNC|Blood product unit 4 expiration|Blood product unit 4 expiration
C2360864|T201|COMP|52111-2|LNC|Blood product unit 3 expiration|Blood product unit 3 expiration
C2360866|T201|COMP|52112-0|LNC|Blood product unit 2 expiration|Blood product unit 2 expiration
C2360868|T201|COMP|52113-8|LNC|Blood product unit 1 expiration|Blood product unit 1 expiration
C2360870|T201|COMP|52114-6|LNC|Direct antiglobulin test.IgG specific reagent|Direct antiglobulin test.IgG specific reagent
C2360871|T201|COMP|52115-3|LNC|D Ab|D Ab
C2360872|T201|COMP|52116-1|LNC|Date blood product unit received|Date blood product unit received
C2360874|T201|COMP|52117-9|LNC|B little x Ab|B little x Ab
C2360876|T201|COMP|52118-7|LNC|Pooled platelets units available|Pooled platelets units available
C2360878|T201|COMP|52119-5|LNC|Apheresis available|Apheresis available
C2360881|T201|COMP|52121-1|LNC|Biopsy|Biopsy
C2361130|T201|COMP|53101-2|LNC|Kynurenate|Kynurenate
C2361131|T201|COMP|53102-0|LNC|Decanoylcarnitine (C10)|Decanoylcarnitine (C10)
C2361132|T201|COMP|53103-8|LNC|Decenoylcarnitine (C10:1)|Decenoylcarnitine (C10:1)
C2361133|T201|COMP|53104-6|LNC|Dodecenoylcarnitine (C12:1)|Dodecenoylcarnitine (C12:1)
C2361134|T201|COMP|53105-3|LNC|3-Hydroxybutyrylcarnitine (C4-OH)|3-Hydroxybutyrylcarnitine (C4-OH)
C2361135|T201|COMP|53106-1|LNC|Butyrylcarnitine (C4)|Butyrylcarnitine (C4)
C2361136|T201|COMP|53107-9|LNC|Kynurenate/Creatinine|Kynurenate/Creatinine
C2361138|T201|COMP|53108-7|LNC|Decenoylcarnitine (C10:1)/Creatinine|Decenoylcarnitine (C10:1)/Creatinine
C2361144|T201|COMP|53040-2|LNC|Drug metabolism sequence variation interpretation|Drug metabolism sequence variation interpretation
C2361146|T201|COMP|53041-0|LNC|DNA region of interest panel|DNA region of interest panel
C2361148|T201|COMP|53042-8|LNC|DNA marker assessed panel|DNA marker assessed panel
C2361150|T201|COMP|53043-6|LNC|DNA marker analysis test coverage panel|DNA marker analysis test coverage panel
C2361152|T201|COMP|52749-9|LNC|Etravirine|Etravirine
C2361153|T201|COMP|52750-7|LNC|Activated protein C resistance|Activated protein C resistance
C2361154|T201|COMP|52751-5|LNC|Coagulation surface induced.factor sensitive|Coagulation surface induced.factor sensitive
C2361160|T201|COMP|52755-6|LNC|Coagulation surface induced.lupus sensitive|Coagulation surface induced.lupus sensitive
C2361162|T201|COMP|52757-2|LNC|SERPINE1 gene.c.-675 4G+5G|SERPINE1 gene.c.-675 4G+5G
C2361164|T201|COMP|52758-0|LNC|SERPINE1 gene.c.-844A>G|SERPINE1 gene.c.-844A>G
C2361166|T201|COMP|52759-8|LNC|Prekallikrein activity actual/Normal|Prekallikrein activity actual/Normal
C2361177|T201|COMP|52765-5|LNC|Thromboelastography without activation panel|Thromboelastography without activation panel
C2361181|T201|COMP|52768-9|LNC|Clot formation|Clot formation
C2361200|T201|COMP|52778-8|LNC|Maximum clot firmness|Maximum clot firmness
C2361212|T201|COMP|52784-6|LNC|Maximum lysis|Maximum lysis
C2361222|T201|COMP|52789-5|LNC|Clotting time|Clotting time
C2361225|T201|COMP|52792-9|LNC|Rh|Rh
C2361226|T201|COMP|52793-7|LNC|ABO group|ABO group
C2361227|T201|COMP|52794-5|LNC|Ova & parasites identified^3rd specimen|Ova & parasites identified^3rd specimen
C2361228|T201|COMP|52795-2|LNC|Ova & parasites identified^2nd specimen|Ova & parasites identified^2nd specimen
C2361231|T201|COMP|52812-5|LNC|Appearance|Appearance
C2361232|T201|COMP|52813-3|LNC|Appearance|Appearance
C2361233|T201|COMP|52814-1|LNC|Appearance|Appearance
C2361234|T201|COMP|52815-8|LNC|Nucleated cells|Nucleated cells
C2361235|T201|COMP|52816-6|LNC|Nucleated cells|Nucleated cells
C2361236|T201|COMP|52817-4|LNC|Nucleated cells|Nucleated cells
C2361237|T201|COMP|52818-2|LNC|Nucleated cells|Nucleated cells
C2361238|T201|COMP|52819-0|LNC|Nucleated cells|Nucleated cells
C2361239|T201|COMP|52820-8|LNC|Appearance|Appearance
C2361240|T201|COMP|52821-6|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C2361241|T201|COMP|52822-4|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C2361242|T201|COMP|52823-2|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C2361243|T201|COMP|52824-0|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C2361244|T201|COMP|52825-7|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C2361299|T201|COMP|52873-7|LNC|Cells.CD1a/100 cells|Cells.CD1a/100 cells
C2361300|T201|COMP|52874-5|LNC|Cells.CD1a/100 cells|Cells.CD1a/100 cells
C2361301|T201|COMP|52875-2|LNC|Cells.CD1a/100 cells|Cells.CD1a/100 cells
C2361302|T201|COMP|52876-0|LNC|Cells.CD1a/100 cells|Cells.CD1a/100 cells
C2361303|T201|COMP|52877-8|LNC|Cells.cytoplasmic CD22/100 cells|Cells.cytoplasmic CD22/100 cells
C2361304|T201|COMP|52878-6|LNC|Cells.cytoplasmic CD22/100 cells|Cells.cytoplasmic CD22/100 cells
C2361305|T201|COMP|52879-4|LNC|Cells.cytoplasmic CD22/100 cells|Cells.cytoplasmic CD22/100 cells
C2361306|T201|COMP|52880-2|LNC|Cells.cytoplasmic CD22/100 cells|Cells.cytoplasmic CD22/100 cells
C2361307|T201|COMP|52881-0|LNC|Cells.cytoplasmic CD22/100 cells|Cells.cytoplasmic CD22/100 cells
C2361308|T201|COMP|52882-8|LNC|Cells.cytoplasmic CD3/100 cells|Cells.cytoplasmic CD3/100 cells
C2361309|T201|COMP|52883-6|LNC|Cells.cytoplasmic CD3/100 cells|Cells.cytoplasmic CD3/100 cells
C2361310|T201|COMP|52884-4|LNC|Cells.cytoplasmic CD3/100 cells|Cells.cytoplasmic CD3/100 cells
C2361311|T201|COMP|52885-1|LNC|Cells.cytoplasmic CD3/100 cells|Cells.cytoplasmic CD3/100 cells
C2361312|T201|COMP|52886-9|LNC|Tellurium|Tellurium
C2361313|T201|COMP|52887-7|LNC|Bismuth|Bismuth
C2361314|T201|COMP|53005-5|LNC|Fibrillarin Ab|Fibrillarin Ab
C2361315|T201|COMP|53006-3|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C2361316|T201|COMP|53007-1|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C2361317|T201|COMP|53008-9|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C2361318|T201|COMP|53009-7|LNC|Ribosomal Ab|Ribosomal Ab
C2361319|T201|COMP|53010-5|LNC|Signal recognition particle Ab|Signal recognition particle Ab
C2361320|T201|COMP|53011-3|LNC|Signal recognition particle Ab|Signal recognition particle Ab
C2361321|T201|COMP|53315-8|LNC|Urinalysis microscopic panel|Urinalysis microscopic panel
C2361322|T201|COMP|53316-6|LNC|Leukocytes|Leukocytes
C2361323|T201|COMP|53317-4|LNC|Leukocyte clumps|Leukocyte clumps
C2361324|T201|COMP|53318-2|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C2361325|T201|COMP|53319-0|LNC|Crystals|Crystals
C2361326|T201|COMP|53320-8|LNC|Casts|Casts
C2361327|T201|COMP|53321-6|LNC|Mucus|Mucus
C2361328|T201|COMP|53322-4|LNC|Crystals|Crystals
C2361350|T201|COMP|52888-5|LNC|Silicon|Silicon
C2361351|T201|COMP|52889-3|LNC|Selenium|Selenium
C2361352|T201|COMP|52890-1|LNC|Lead|Lead
C2361353|T201|COMP|52891-9|LNC|Chromium|Chromium
C2361354|T201|COMP|52892-7|LNC|Aluminum|Aluminum
C2361355|T201|COMP|52893-5|LNC|Vanadium|Vanadium
C2361356|T201|COMP|52894-3|LNC|Titanium|Titanium
C2361357|T201|COMP|52895-0|LNC|Tellurium|Tellurium
C2361358|T201|COMP|52896-8|LNC|Silver|Silver
C2361359|T201|COMP|52897-6|LNC|Platinum|Platinum
C2361360|T201|COMP|52898-4|LNC|Bismuth|Bismuth
C2361361|T201|COMP|52899-2|LNC|Beryllium|Beryllium
C2361362|T201|COMP|52900-8|LNC|Vanadium/Creatinine|Vanadium/Creatinine
C2361363|T201|COMP|52901-6|LNC|Vanadium/Creatinine|Vanadium/Creatinine
C2361364|T201|COMP|52902-4|LNC|Uranium/Creatinine|Uranium/Creatinine
C2361365|T201|COMP|52903-2|LNC|Uranium/Creatinine|Uranium/Creatinine
C2361366|T201|COMP|52904-0|LNC|Silver/Creatinine|Silver/Creatinine
C2361367|T201|COMP|52905-7|LNC|Silver/Creatinine|Silver/Creatinine
C2361368|T201|COMP|52906-5|LNC|Bismuth/Creatinine|Bismuth/Creatinine
C2361369|T201|COMP|52907-3|LNC|Bismuth/Creatinine|Bismuth/Creatinine
C2361370|T201|COMP|52908-1|LNC|Selenium|Selenium
C2361371|T201|COMP|52909-9|LNC|Platinum|Platinum
C2361372|T201|COMP|52910-7|LNC|Zinc|Zinc
C2361373|T201|COMP|52911-5|LNC|Magnesium|Magnesium
C2361374|T201|COMP|52912-3|LNC|Copper|Copper
C2361375|T201|COMP|52913-1|LNC|Selenium|Selenium
C2361376|T201|COMP|52914-9|LNC|Boron|Boron
C2361377|T201|COMP|52915-6|LNC|Aluminum|Aluminum
C2361378|T201|COMP|52916-4|LNC|Tin/Creatinine|Tin/Creatinine
C2361379|T201|COMP|52917-2|LNC|Tin/Creatinine|Tin/Creatinine
C2361380|T201|COMP|52918-0|LNC|Thallium/Creatinine|Thallium/Creatinine
C2361381|T201|COMP|52919-8|LNC|Tellurium/Creatinine|Tellurium/Creatinine
C2361382|T201|COMP|52920-6|LNC|Tellurium/Creatinine|Tellurium/Creatinine
C2361383|T201|COMP|52921-4|LNC|Strontium/Creatinine|Strontium/Creatinine
C2361384|T201|COMP|52922-2|LNC|Strontium/Creatinine|Strontium/Creatinine
C2361385|T201|COMP|52923-0|LNC|Selenium/Creatinine|Selenium/Creatinine
C2361386|T201|COMP|52924-8|LNC|Platinum/Creatinine|Platinum/Creatinine
C2361388|T201|COMP|52925-5|LNC|Platinum/Creatinine|Platinum/Creatinine
C2361389|T201|COMP|52926-3|LNC|Nickel/Creatinine|Nickel/Creatinine
C2361390|T201|COMP|52927-1|LNC|Molybdenum/Creatinine|Molybdenum/Creatinine
C2361391|T201|COMP|52936-2|LNC|Beryllium/Creatinine|Beryllium/Creatinine
C2361392|T201|COMP|52937-0|LNC|Barium/Creatinine|Barium/Creatinine
C2361393|T201|COMP|52938-8|LNC|Barium/Creatinine|Barium/Creatinine
C2361394|T201|COMP|52939-6|LNC|Arsenic.inorganic/Creatinine|Arsenic.inorganic/Creatinine
C2361395|T201|COMP|52940-4|LNC|Arsenic.inorganic/Creatinine|Arsenic.inorganic/Creatinine
C2361396|T201|COMP|52941-2|LNC|Antimony/Creatinine|Antimony/Creatinine
C2361397|T201|COMP|52942-0|LNC|Antimony/Creatinine|Antimony/Creatinine
C2361398|T201|COMP|52943-8|LNC|Aluminum/Creatinine|Aluminum/Creatinine
C2361399|T201|COMP|53250-7|LNC|Influenza virus A RNA|Influenza virus A RNA
C2361400|T201|COMP|53251-5|LNC|Influenza virus B RNA|Influenza virus B RNA
C2361401|T201|COMP|53252-3|LNC|Parainfluenza virus 1 RNA|Parainfluenza virus 1 RNA
C2361402|T201|COMP|53253-1|LNC|Parainfluenza virus 2 RNA|Parainfluenza virus 2 RNA
C2361403|T201|COMP|53254-9|LNC|Parainfluenza virus 3 RNA|Parainfluenza virus 3 RNA
C2361404|T201|COMP|53255-6|LNC|Mycoplasma pneumoniae DNA|Mycoplasma pneumoniae DNA
C2361405|T201|COMP|53391-9|LNC|Trichothecene Ab.IgM|Trichothecene Ab.IgM
C2361406|T201|COMP|53392-7|LNC|Proline/Phenylalanine|Proline/Phenylalanine
C2361410|T201|COMP|53394-3|LNC|5-Oxoproline+Pipecolate/Phenylalanine|5-Oxoproline+Pipecolate/Phenylalanine
C2361412|T201|COMP|53395-0|LNC|Asparagine+Ornithine/Serine|Asparagine+Ornithine/Serine
C2361414|T201|COMP|53396-8|LNC|Asparagine+Ornithine/Phenylalanine|Asparagine+Ornithine/Phenylalanine
C2361418|T201|COMP|53398-4|LNC|Arginine/Phenylalanine|Arginine/Phenylalanine
C2361420|T201|COMP|53399-2|LNC|Citrulline/Tyrosine|Citrulline/Tyrosine
C2361422|T201|COMP|53400-8|LNC|Stearoylcarnitine (C18)/Propionylcarnitine (C3)|Stearoylcarnitine (C18)/Propionylcarnitine (C3)
C2361430|T201|COMP|52944-6|LNC|Aluminum/Creatinine|Aluminum/Creatinine
C2361431|T201|COMP|52945-3|LNC|LORazepam|LORazepam
C2361432|T201|COMP|52946-1|LNC|diazePAM|diazePAM
C2361433|T201|COMP|52947-9|LNC|Dextromethorphan|Dextromethorphan
C2361434|T201|COMP|52948-7|LNC|cloBAZam|cloBAZam
C2361435|T201|COMP|52949-5|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2361436|T201|COMP|52950-3|LNC|Barbital|Barbital
C2361437|T201|COMP|52951-1|LNC|Phencyclidine|Phencyclidine
C2361438|T201|COMP|52952-9|LNC|Opiates|Opiates
C2361439|T201|COMP|52953-7|LNC|Cocaine|Cocaine
C2361440|T201|COMP|52954-5|LNC|Cannabinoids|Cannabinoids
C2361441|T201|COMP|52955-2|LNC|Benzodiazepines|Benzodiazepines
C2361442|T201|COMP|52956-0|LNC|Barbiturates|Barbiturates
C2361443|T201|COMP|52957-8|LNC|Amphetamine|Amphetamine
C2361444|T201|COMP|52958-6|LNC|Methadone|Methadone
C2361445|T201|COMP|52959-4|LNC|cloBAZam|cloBAZam
C2361446|T201|COMP|52960-2|LNC|cloNIDine|cloNIDine
C2361447|T201|COMP|52961-0|LNC|Paraquat|Paraquat
C2361448|T201|COMP|52962-8|LNC|Tobramycin|Tobramycin
C2361449|T201|COMP|52963-6|LNC|Flurazepam|Flurazepam
C2361450|T201|COMP|52964-4|LNC|cloBAZam|cloBAZam
C2361451|T201|COMP|52965-1|LNC|clonazePAM|clonazePAM
C2361452|T201|COMP|52966-9|LNC|Bacteria identified|Bacteria identified
C2361453|T201|COMP|52967-7|LNC|Bacteria identified|Bacteria identified
C2361454|T201|COMP|52968-5|LNC|Streptococcus agalactiae|Streptococcus agalactiae
C2361456|T201|COMP|52970-1|LNC|CV2 Ab|CV2 Ab
C2361457|T201|COMP|52971-9|LNC|Immune complex|Immune complex
C2361459|T201|COMP|52973-5|LNC|Bacteria identified|Bacteria identified
C2361460|T201|COMP|52974-3|LNC|Influenza virus B Ab|Influenza virus B Ab
C2361461|T201|COMP|52975-0|LNC|Respiratory syncytial virus Ab|Respiratory syncytial virus Ab
C2361462|T201|COMP|52976-8|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C2361463|T201|COMP|52977-6|LNC|Herpes simplex virus Ab|Herpes simplex virus Ab
C2361464|T201|COMP|52978-4|LNC|Varicella zoster virus Ab|Varicella zoster virus Ab
C2361465|T201|COMP|52979-2|LNC|Trichinella spiralis Ab.IgG|Trichinella spiralis Ab.IgG
C2361466|T201|COMP|52980-0|LNC|Plasmodium sp Ab.IgG|Plasmodium sp Ab.IgG
C2361468|T201|COMP|52981-8|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C2361469|T201|COMP|52982-6|LNC|Echinococcus sp Ab.IgG1|Echinococcus sp Ab.IgG1
C2361471|T201|COMP|52983-4|LNC|Echinococcus sp Ab.IgG4|Echinococcus sp Ab.IgG4
C2361473|T201|COMP|52984-2|LNC|Cytomegalovirus Ab.IgG avidity|Cytomegalovirus Ab.IgG avidity
C2361474|T201|COMP|52985-9|LNC|Leishmania sp Ab.IgG|Leishmania sp Ab.IgG
C2361475|T201|COMP|52986-7|LNC|Rubella virus Ab.IgG avidity|Rubella virus Ab.IgG avidity
C2361476|T201|COMP|52987-5|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C2361477|T201|COMP|52988-3|LNC|Leptospira sp DNA|Leptospira sp DNA
C2361478|T201|COMP|52989-1|LNC|Leptospira sp DNA|Leptospira sp DNA
C2361479|T201|COMP|52990-9|LNC|Leptospira sp DNA|Leptospira sp DNA
C2361480|T201|COMP|52991-7|LNC|Cells.cytoplasmic CD79a/100 cells|Cells.cytoplasmic CD79a/100 cells
C2361482|T201|COMP|52992-5|LNC|Cells.cytoplasmic CD79a/100 cells|Cells.cytoplasmic CD79a/100 cells
C2361483|T201|COMP|52993-3|LNC|Cells.cytoplasmic CD79a/100 cells|Cells.cytoplasmic CD79a/100 cells
C2361484|T201|COMP|52994-1|LNC|Cells.cytoplasmic CD79a/100 cells|Cells.cytoplasmic CD79a/100 cells
C2361485|T201|COMP|52995-8|LNC|Cells.cytoplasmic CD79a/100 cells|Cells.cytoplasmic CD79a/100 cells
C2361489|T201|COMP|52999-0|LNC|Leukocytes.disintegrated|Leukocytes.disintegrated
C2361491|T201|COMP|53000-6|LNC|Mitochondria M4 Ab|Mitochondria M4 Ab
C2361492|T201|COMP|53001-4|LNC|Mitochondria M9 Ab|Mitochondria M9 Ab
C2361493|T201|COMP|53002-2|LNC|Nuclear Ab pattern.fine speckled|Nuclear Ab pattern.fine speckled
C2361494|T201|COMP|53003-0|LNC|Mitotic spindle apparatus Ab|Mitotic spindle apparatus Ab
C2361495|T201|COMP|53004-8|LNC|Mitotic spindle apparatus Ab|Mitotic spindle apparatus Ab
C2361496|T201|COMP|53012-1|LNC|Neutrophil cytoplasmic Ab.atypical|Neutrophil cytoplasmic Ab.atypical
C2361497|T201|COMP|53013-9|LNC|Bactericidal permeability increasing protein Ab|Bactericidal permeability increasing protein Ab
C2361498|T201|COMP|53014-7|LNC|Nucleosome Ab|Nucleosome Ab
C2361499|T201|COMP|53015-4|LNC|Nucleosome Ab|Nucleosome Ab
C2361500|T201|COMP|53016-2|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C2361502|T201|COMP|53017-0|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C2361503|T201|COMP|53018-8|LNC|Sjogrens syndrome-A extractable nuclear 60kD Ab|Sjogrens syndrome-A extractable nuclear 60kD Ab
C2361505|T201|COMP|53019-6|LNC|Sjogrens syndrome-A extractable nuclear 60kD Ab|Sjogrens syndrome-A extractable nuclear 60kD Ab
C2361506|T201|COMP|53020-4|LNC|Complement C1q Ab|Complement C1q Ab
C2361507|T201|COMP|53021-2|LNC|Salivary gland Ab|Salivary gland Ab
C2361508|T201|COMP|53022-0|LNC|U1 small nuclear ribonucleoprotein Ab|U1 small nuclear ribonucleoprotein Ab
C2361509|T201|COMP|53023-8|LNC|Tissue transglutaminase Ab|Tissue transglutaminase Ab
C2361510|T201|COMP|53024-6|LNC|Saccharomyces cerevisiae Ab|Saccharomyces cerevisiae Ab
C2361511|T201|COMP|53025-3|LNC|Gliadin Ab|Gliadin Ab
C2361512|T201|COMP|53026-1|LNC|Tissue transglutaminase Ab.IgG|Tissue transglutaminase Ab.IgG
C2361513|T201|COMP|53027-9|LNC|Cyclic citrullinated peptide Ab|Cyclic citrullinated peptide Ab
C2361514|T201|COMP|53028-7|LNC|Cyclic citrullinated peptide Ab|Cyclic citrullinated peptide Ab
C2361515|T201|COMP|53029-5|LNC|Neutrophil cytoplasmic Ab.perinuclear.atypical|Neutrophil cytoplasmic Ab.perinuclear.atypical
C2361516|T201|COMP|53030-3|LNC|Liver kidney microsomal Ab|Liver kidney microsomal Ab
C2361517|T201|COMP|53031-1|LNC|Signal recognition particle Ab|Signal recognition particle Ab
C2361518|T201|COMP|53032-9|LNC|U1 small nuclear ribonucleoprotein 70kD Ab|U1 small nuclear ribonucleoprotein 70kD Ab
C2361522|T201|COMP|53034-5|LNC|Allelic state|Allelic state
C2361524|T201|COMP|53035-2|LNC|DNA marker assessed|DNA marker assessed
C2361526|T201|COMP|53036-0|LNC|Filler DNA analysis test identifier|Filler DNA analysis test identifier
C2361528|T201|COMP|53037-8|LNC|Genetic disease sequence variation interpretation|Genetic disease sequence variation interpretation
C2361530|T201|COMP|53044-4|LNC|DNA marker identified panel|DNA marker identified panel
C2361532|T201|COMP|53045-1|LNC|Reference sequence alteration|Reference sequence alteration
C2361534|T201|COMP|53046-9|LNC|Beta globulin+Gamma globulin|Beta globulin+Gamma globulin
C2361535|T201|COMP|53047-7|LNC|Chromogranin A|Chromogranin A
C2361536|T201|COMP|53048-5|LNC|Ferritin|Ferritin
C2361537|T201|COMP|53049-3|LNC|Glucose^pre-meal|Glucose^pre-meal
C2361538|T201|COMP|53050-1|LNC|Glucose|Glucose
C2361539|T201|COMP|53051-9|LNC|Beta globulin+Gamma globulin/Protein.total|Beta globulin+Gamma globulin/Protein.total
C2361540|T201|COMP|53052-7|LNC|Collagen crosslinked C-telopeptide|Collagen crosslinked C-telopeptide
C2361541|T201|COMP|53053-5|LNC|Carnitine|Carnitine
C2361542|T201|COMP|53054-3|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C2361543|T201|COMP|53055-0|LNC|Creatine|Creatine
C2361544|T201|COMP|53056-8|LNC|Decanoylcarnitine (C10)|Decanoylcarnitine (C10)
C2361545|T201|COMP|53057-6|LNC|Decenoylcarnitine (C10:1)|Decenoylcarnitine (C10:1)
C2361546|T201|COMP|53058-4|LNC|Dodecanoylcarnitine (C12)|Dodecanoylcarnitine (C12)
C2361547|T201|COMP|53059-2|LNC|Dodecenoylcarnitine (C12:1)|Dodecenoylcarnitine (C12:1)
C2361548|T201|COMP|53060-0|LNC|Butyrylcarnitine (C4)|Butyrylcarnitine (C4)
C2361549|T201|COMP|53061-8|LNC|Ketones|Ketones
C2361550|T201|COMP|53062-6|LNC|Argininosuccinate|Argininosuccinate
C2361551|T201|COMP|53063-4|LNC|Beta alanine|Beta alanine
C2361552|T201|COMP|53064-2|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C2361553|T201|COMP|53065-9|LNC|Butyrylcarnitine (C4)|Butyrylcarnitine (C4)
C2361554|T201|COMP|53066-7|LNC|Cystathionine|Cystathionine
C2361555|T201|COMP|53067-5|LNC|Argininosuccinate|Argininosuccinate
C2361556|T201|COMP|53068-3|LNC|Beta alanine|Beta alanine
C2361557|T201|COMP|53069-1|LNC|Cystathionine|Cystathionine
C2361558|T201|COMP|53070-9|LNC|Butyrylcarnitine (C4)|Butyrylcarnitine (C4)
C2361559|T201|COMP|53071-7|LNC|Carnitine|Carnitine
C2361560|T201|COMP|53072-5|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C2361561|T201|COMP|53073-3|LNC|Ceruloplasmin|Ceruloplasmin
C2361562|T201|COMP|53074-1|LNC|Creatine|Creatine
C2361563|T201|COMP|53075-8|LNC|Decanoylcarnitine (C10)|Decanoylcarnitine (C10)
C2361564|T201|COMP|53076-6|LNC|Decenoylcarnitine (C10:1)|Decenoylcarnitine (C10:1)
C2361565|T201|COMP|53077-4|LNC|Levodopa|Levodopa
C2361566|T201|COMP|53078-2|LNC|Dodecanoylcarnitine (C12)|Dodecanoylcarnitine (C12)
C2361567|T201|COMP|53079-0|LNC|Dodecenoylcarnitine (C12:1)|Dodecenoylcarnitine (C12:1)
C2361568|T201|COMP|53080-8|LNC|Cystine|Cystine
C2361569|T201|COMP|53081-6|LNC|Ammonia|Ammonia
C2361570|T201|COMP|53082-4|LNC|Cholesterol|Cholesterol
C2361571|T201|COMP|53083-2|LNC|Bilirubin.glucuronidated|Bilirubin.glucuronidated
C2361572|T201|COMP|53084-0|LNC|Glucose|Glucose
C2361573|T201|COMP|53085-7|LNC|Base excess|Base excess
C2361574|T201|COMP|53086-5|LNC|Bicarbonate|Bicarbonate
C2361575|T201|COMP|53087-3|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C2361576|T201|COMP|53088-1|LNC|Calcium.ionized|Calcium.ionized
C2361577|T201|COMP|53089-9|LNC|Carbon dioxide|Carbon dioxide
C2361578|T201|COMP|53090-7|LNC|Carbon dioxide|Carbon dioxide
C2361579|T201|COMP|53091-5|LNC|Nitrogen.nonprotein|Nitrogen.nonprotein
C2361580|T201|COMP|53092-3|LNC|Collagen crosslinked C-telopeptide|Collagen crosslinked C-telopeptide
C2361581|T201|COMP|53093-1|LNC|Glucose^post XXX challenge|Glucose^post XXX challenge
C2361582|T201|COMP|53094-9|LNC|Glucose^post meal|Glucose^post meal
C2361583|T201|COMP|53095-6|LNC|Carnitine.free (C0)/Carnitine.total|Carnitine.free (C0)/Carnitine.total
C2361584|T201|COMP|53096-4|LNC|Carnitine.free (C0)/Carnitine.total|Carnitine.free (C0)/Carnitine.total
C2361585|T201|COMP|53097-2|LNC|3-O-Methyldopa|3-O-Methyldopa
C2361586|T201|COMP|53098-0|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C2361587|T201|COMP|53099-8|LNC|Chloride|Chloride
C2361588|T201|COMP|53100-4|LNC|Calcium|Calcium
C2361589|T201|COMP|53109-5|LNC|Docosenoate/Creatinine|Docosenoate/Creatinine
C2361591|T201|COMP|53110-3|LNC|5-Hydroxytryptophan/Creatinine|5-Hydroxytryptophan/Creatinine
C2361592|T201|COMP|53111-1|LNC|Butyrylcarnitine (C4)/Creatinine|Butyrylcarnitine (C4)/Creatinine
C2361594|T201|COMP|53112-9|LNC|Carnitine.free (C0)/Carnitine.total|Carnitine.free (C0)/Carnitine.total
C2361595|T201|COMP|53113-7|LNC|Spermatids/100 spermatozoa|Spermatids/100 spermatozoa
C2361597|T201|COMP|53114-5|LNC|Glucose^post CFst|Glucose^post CFst
C2361598|T201|COMP|53115-2|LNC|Granulocytes.immature|Granulocytes.immature
C2361599|T201|COMP|53116-0|LNC|Base deficit|Base deficit
C2361600|T201|COMP|53117-8|LNC|Hemoglobin.thermolabile|Hemoglobin.thermolabile
C2361601|T201|COMP|53118-6|LNC|Sulfonamide crystals|Sulfonamide crystals
C2361602|T201|COMP|53119-4|LNC|Tyrosine crystals|Tyrosine crystals
C2361603|T201|COMP|53120-2|LNC|Creatinine|Creatinine
C2361604|T201|COMP|53121-0|LNC|Protein|Protein
C2361605|T201|COMP|53122-8|LNC|Sodium|Sodium
C2361606|T201|COMP|53123-6|LNC|Potassium|Potassium
C2361607|T201|COMP|53124-4|LNC|Calcium|Calcium
C2361608|T201|COMP|53125-1|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C2361609|T201|COMP|53126-9|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C2361610|T201|COMP|53127-7|LNC|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C2361611|T201|COMP|53128-5|LNC|Bacterial casts|Bacterial casts
C2361612|T201|COMP|53129-3|LNC|Sodium urate crystals|Sodium urate crystals
C2361613|T201|COMP|53130-1|LNC|Ammonium urate crystals|Ammonium urate crystals
C2361614|T201|COMP|53131-9|LNC|Calcium oxalate crystals|Calcium oxalate crystals
C2361615|T201|COMP|53132-7|LNC|Epithelial cells.non-squamous|Epithelial cells.non-squamous
C2361616|T201|COMP|53133-5|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C2361617|T201|COMP|53134-3|LNC|Amylase isoenzymes|Amylase isoenzymes
C2361618|T201|COMP|53135-0|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C2361619|T201|COMP|53136-8|LNC|Organic acids pattern|Organic acids pattern
C2361620|T201|COMP|53137-6|LNC|Urea|Urea
C2361621|T201|COMP|53138-4|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C2361622|T201|COMP|53139-2|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C2361623|T201|COMP|53140-0|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C2361624|T201|COMP|53141-8|LNC|17-Hydroxyprogesterone^30M post XXX challenge|17-Hydroxyprogesterone^30M post XXX challenge
C2361625|T201|COMP|53142-6|LNC|Nitrogen|Nitrogen
C2361626|T201|COMP|53143-4|LNC|Hydrogen ion|Hydrogen ion
C2361627|T201|COMP|53144-2|LNC|Somatotropin^75M post XXX challenge|Somatotropin^75M post XXX challenge
C2361628|T201|COMP|53145-9|LNC|Lutropin^45M post XXX challenge|Lutropin^45M post XXX challenge
C2361629|T201|COMP|53146-7|LNC|Follitropin^45M post XXX challenge|Follitropin^45M post XXX challenge
C2361630|T201|COMP|53147-5|LNC|Follitropin^2H post XXX challenge|Follitropin^2H post XXX challenge
C2361631|T201|COMP|53148-3|LNC|DNA double strand Ab|DNA double strand Ab
C2361632|T201|COMP|53149-1|LNC|Iron/Creatinine|Iron/Creatinine
C2361633|T201|COMP|53150-9|LNC|Alanine+Beta Alanine+Sarcosine|Alanine+Beta Alanine+Sarcosine
C2361635|T201|COMP|53151-7|LNC|Valine/Phenylalanine|Valine/Phenylalanine
C2361637|T201|COMP|53152-5|LNC|Alloisoleucine+Isoleucine+Leucine+Hydroxyproline|Alloisoleucine+Isoleucine+Leucine+Hydroxyproline
C2361643|T201|COMP|53155-8|LNC|Asparagine+Ornithine|Asparagine+Ornithine
C2361645|T201|COMP|53156-6|LNC|Methionine/Phenylalanine|Methionine/Phenylalanine
C2361647|T201|COMP|53157-4|LNC|Citrulline/Phenylalanine|Citrulline/Phenylalanine
C2361649|T201|COMP|53173-1|LNC|3-Hydroxyhexanoylcarnitine (C6-OH)|3-Hydroxyhexanoylcarnitine (C6-OH)
C2361650|T201|COMP|53174-9|LNC|Octenoylcarnitine (C8:1)|Octenoylcarnitine (C8:1)
C2361651|T201|COMP|53175-6|LNC|Octanoylcarnitine (C8)|Octanoylcarnitine (C8)
C2361652|T201|COMP|53176-4|LNC|Octanoylcarnitine (C8)/Acetylcarnitine (C2)|Octanoylcarnitine (C8)/Acetylcarnitine (C2)
C2361654|T201|COMP|53177-2|LNC|Octanoylcarnitine (C8)/Decanoylcarnitine (C10)|Octanoylcarnitine (C8)/Decanoylcarnitine (C10)
C2361660|T201|COMP|53180-6|LNC|Decadienoylcarnitine (C10:2)|Decadienoylcarnitine (C10:2)
C2361664|T201|COMP|53182-2|LNC|3-Hydroxydecenoylcarnitine (C10:1-OH)|3-Hydroxydecenoylcarnitine (C10:1-OH)
C2361673|T201|COMP|53187-1|LNC|Methylglutarylcarnitine (C6-DC)|Methylglutarylcarnitine (C6-DC)
C2361675|T201|COMP|53188-9|LNC|3-Hydroxydodecenoylcarnitine (C12:1-OH)|3-Hydroxydodecenoylcarnitine (C12:1-OH)
C2361677|T201|COMP|53189-7|LNC|3-Hydroxydodecanoylcarnitine (C12-OH)|3-Hydroxydodecanoylcarnitine (C12-OH)
C2361678|T201|COMP|53190-5|LNC|Tetradecadienoylcarnitine (C14:2)|Tetradecadienoylcarnitine (C14:2)
C2361679|T201|COMP|53191-3|LNC|Tetradecenoylcarnitine (C14:1)|Tetradecenoylcarnitine (C14:1)
C2361680|T201|COMP|53192-1|LNC|Tetradecanoylcarnitine (C14)|Tetradecanoylcarnitine (C14)
C2361687|T201|COMP|53196-2|LNC|3-Hydroxytetradecadienoylcarnitine (C14:2-OH)|3-Hydroxytetradecadienoylcarnitine (C14:2-OH)
C2361689|T201|COMP|53197-0|LNC|3-Hydroxytetradecenoylcarnitine (C14:1-OH)|3-Hydroxytetradecenoylcarnitine (C14:1-OH)
C2361690|T201|COMP|53198-8|LNC|Palmitoleylcarnitine (C16:1)|Palmitoleylcarnitine (C16:1)
C2361691|T201|COMP|53199-6|LNC|Palmitoylcarnitine (C16)|Palmitoylcarnitine (C16)
C2361692|T201|COMP|53200-2|LNC|Argininosuccinate/Arginine|Argininosuccinate/Arginine
C2361696|T201|COMP|53202-8|LNC|Oleoylcarnitine (C18:1)|Oleoylcarnitine (C18:1)
C2361697|T201|COMP|53203-6|LNC|Hexenoylcarnitine (C6:1)|Hexenoylcarnitine (C6:1)
C2361699|T201|COMP|53204-4|LNC|Heptanoylcarnitine (C7)|Heptanoylcarnitine (C7)
C2361701|T201|COMP|53205-1|LNC|Phenylacetylcarnitine (PheC2)|Phenylacetylcarnitine (PheC2)
C2361703|T201|COMP|53206-9|LNC|Salicylylcarnitine (Salc)|Salicylylcarnitine (Salc)
C2361705|T201|COMP|53207-7|LNC|Nonanoylcarnitine (C9)|Nonanoylcarnitine (C9)
C2361707|T201|COMP|53208-5|LNC|Decatrienoylcarnitine (C10:3)|Decatrienoylcarnitine (C10:3)
C2361709|T201|COMP|53209-3|LNC|Dehydrosuberylcarnitine (C8:1-DC)|Dehydrosuberylcarnitine (C8:1-DC)
C2361711|T201|COMP|53210-1|LNC|Suberylcarnitine (C8-DC)|Suberylcarnitine (C8-DC)
C2361712|T201|COMP|53211-9|LNC|Dehydrosebacylcarnitine (C10:1-DC)|Dehydrosebacylcarnitine (C10:1-DC)
C2361714|T201|COMP|53212-7|LNC|Sebacylcarnitine (C10-DC)|Sebacylcarnitine (C10-DC)
C2361716|T201|COMP|53213-5|LNC|Dicarboxydodecenoylcarnitine (C12:1-DC)|Dicarboxydodecenoylcarnitine (C12:1-DC)
C2361718|T201|COMP|53214-3|LNC|Dicarboxydodecanoylcarnitine (C12-DC)|Dicarboxydodecanoylcarnitine (C12-DC)
C2361720|T201|COMP|53215-0|LNC|Dicarboxytetradecenoylcarnitine (C14:1-DC)|Dicarboxytetradecenoylcarnitine (C14:1-DC)
C2361722|T201|COMP|53216-8|LNC|Dicarboxytetradecanoylcarnitine (C14-DC)|Dicarboxytetradecanoylcarnitine (C14-DC)
C2361724|T201|COMP|53217-6|LNC|Dicarboxypalmitoleylcarnitine (C16:1-DC)|Dicarboxypalmitoleylcarnitine (C16:1-DC)
C2361726|T201|COMP|54479-1|LNC|Dicarboxypalmitolycarnitine (C16-DC)|Dicarboxypalmitolycarnitine (C16-DC)
C2361726|T201|COMP|53218-4|LNC|Dicarboxypalmitoylcarnitine (C16-DC)|Dicarboxypalmitoylcarnitine (C16-DC)
C2361728|T201|COMP|53219-2|LNC|Dicarboxyoleylcarnitine (C18:1-DC)|Dicarboxyoleylcarnitine (C18:1-DC)
C2361730|T201|COMP|53220-0|LNC|Dicarboxystearoylcarnitine (C18-DC)|Dicarboxystearoylcarnitine (C18-DC)
C2361732|T201|COMP|53221-8|LNC|Coagulation dilute Russell viper venom induced|Coagulation dilute Russell viper venom induced
C2361733|T201|COMP|53222-6|LNC|Coagulation factor XI activated activity|Coagulation factor XI activated activity
C2361734|T201|COMP|53223-4|LNC|Hemoglobin G/Hemoglobin.total|Hemoglobin G/Hemoglobin.total
C2361736|T201|COMP|53224-2|LNC|Hemoglobin M|Hemoglobin M
C2361737|T201|COMP|53225-9|LNC|Leukocytes|Leukocytes
C2361738|T201|COMP|53226-7|LNC|Leukocytes|Leukocytes
C2361739|T201|COMP|53227-5|LNC|Leukocytes|Leukocytes
C2361740|T201|COMP|53229-1|LNC|Prealbumin|Prealbumin
C2361742|T201|COMP|53231-7|LNC|Succinylacetone|Succinylacetone
C2361743|T201|COMP|53232-5|LNC|5-Oxoproline+Pipecolate|5-Oxoproline+Pipecolate
C2361745|T201|COMP|53233-3|LNC|Carnitine.free (C0)/Palmitoylcarnitine (C16)|Carnitine.free (C0)/Palmitoylcarnitine (C16)
C2361747|T201|COMP|53234-1|LNC|Carnitine.free (C0)/Stearoylcarnitine (C18)|Carnitine.free (C0)/Stearoylcarnitine (C18)
C2361753|T201|COMP|53237-4|LNC|Acrylylcarnitine (C3:1)|Acrylylcarnitine (C3:1)
C2361760|T201|COMP|53241-6|LNC|Stearoylcarnitine (C18)|Stearoylcarnitine (C18)
C2361773|T201|COMP|53248-1|LNC|Plasmodium sp lactate dehydrogenase|Plasmodium sp lactate dehydrogenase
C2361774|T201|COMP|53249-9|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C2361775|T201|COMP|53256-4|LNC|Enterovirus RNA|Enterovirus RNA
C2361776|T201|COMP|53257-2|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C2361777|T201|COMP|53258-0|LNC|Beta vulgaris Ab.IgE.RAST class|Beta vulgaris Ab.IgE.RAST class
C2361779|T201|COMP|53259-8|LNC|Glomerular basement membrane Ab|Glomerular basement membrane Ab
C2361780|T201|COMP|53260-6|LNC|Glomerular basement membrane Ab|Glomerular basement membrane Ab
C2361781|T201|COMP|53261-4|LNC|Amino acid newborn screen panel|Amino acid newborn screen panel
C2361783|T201|COMP|53262-2|LNC|Carnitine newborn screen panel|Carnitine newborn screen panel
C2361785|T201|COMP|53263-0|LNC|Urinalysis yeast variants panel|Urinalysis yeast variants panel
C2361787|T201|COMP|53264-8|LNC|Urinalysis yeast variants panel|Urinalysis yeast variants panel
C2361788|T201|COMP|53265-5|LNC|Yeast.hyphae|Yeast.hyphae
C2361789|T201|COMP|53266-3|LNC|Yeast.budding|Yeast.budding
C2361790|T201|COMP|53267-1|LNC|Urinalysis yeast variants panel|Urinalysis yeast variants panel
C2361791|T201|COMP|53268-9|LNC|Yeast.hyphae|Yeast.hyphae
C2361792|T201|COMP|53269-7|LNC|Yeast.budding|Yeast.budding
C2361795|T201|COMP|53271-3|LNC|Epithelial cells.renal|Epithelial cells.renal
C2361796|T201|COMP|53272-1|LNC|Transitional cells|Transitional cells
C2361798|T201|COMP|53274-7|LNC|Epithelial cells.renal|Epithelial cells.renal
C2361799|T201|COMP|53275-4|LNC|Transitional cells|Transitional cells
C2361801|T201|COMP|53277-0|LNC|Urinalysis type of cast panel|Urinalysis type of cast panel
C2361803|T201|COMP|53278-8|LNC|Erythrocyte casts|Erythrocyte casts
C2361804|T201|COMP|53279-6|LNC|Leukocyte casts|Leukocyte casts
C2361805|T201|COMP|53280-4|LNC|Casts type not specified|Casts type not specified
C2361807|T201|COMP|53281-2|LNC|Urinalysis type of cast panel|Urinalysis type of cast panel
C2361808|T201|COMP|53282-0|LNC|Granular casts|Granular casts
C2361809|T201|COMP|53283-8|LNC|Mixed cellular casts|Mixed cellular casts
C2361810|T201|COMP|53284-6|LNC|Broad casts|Broad casts
C2361811|T201|COMP|53285-3|LNC|Erythrocyte casts|Erythrocyte casts
C2361812|T201|COMP|53286-1|LNC|Leukocyte casts|Leukocyte casts
C2361813|T201|COMP|53287-9|LNC|Epithelial casts|Epithelial casts
C2361814|T201|COMP|53288-7|LNC|Fatty casts|Fatty casts
C2361815|T201|COMP|53289-5|LNC|Mixed cellular casts|Mixed cellular casts
C2361816|T201|COMP|53290-3|LNC|Broad casts|Broad casts
C2361817|T201|COMP|53291-1|LNC|Epithelial casts|Epithelial casts
C2361818|T201|COMP|53292-9|LNC|Erythrocytes|Erythrocytes
C2361819|T201|COMP|53293-7|LNC|Urinalysis microscopic panel|Urinalysis microscopic panel
C2361820|T201|COMP|53294-5|LNC|Epithelial cells.non-squamous|Epithelial cells.non-squamous
C2361821|T201|COMP|53295-2|LNC|Urinalysis type of crystal panel|Urinalysis type of crystal panel
C2361823|T201|COMP|53296-0|LNC|Calcium oxalate crystals|Calcium oxalate crystals
C2361824|T201|COMP|53297-8|LNC|Crystals unspecified|Crystals unspecified
C2361826|T201|COMP|53298-6|LNC|Triple phosphate crystals|Triple phosphate crystals
C2361827|T201|COMP|53299-4|LNC|Calcium phosphate crystals|Calcium phosphate crystals
C2361828|T201|COMP|53300-0|LNC|Leucine crystals|Leucine crystals
C2361829|T201|COMP|53301-8|LNC|Urate crystals|Urate crystals
C2361830|T201|COMP|53302-6|LNC|Calcium carbonate crystals|Calcium carbonate crystals
C2361831|T201|COMP|53303-4|LNC|Cystine crystals|Cystine crystals
C2361832|T201|COMP|53304-2|LNC|Tyrosine crystals|Tyrosine crystals
C2361833|T201|COMP|53305-9|LNC|Urinalysis type of crystal panel|Urinalysis type of crystal panel
C2361834|T201|COMP|53306-7|LNC|Calcium oxalate crystals|Calcium oxalate crystals
C2361835|T201|COMP|53307-5|LNC|Crystals unspecified|Crystals unspecified
C2361836|T201|COMP|53308-3|LNC|Triple phosphate crystals|Triple phosphate crystals
C2361837|T201|COMP|53309-1|LNC|Calcium phosphate crystals|Calcium phosphate crystals
C2361838|T201|COMP|53310-9|LNC|Leucine crystals|Leucine crystals
C2361839|T201|COMP|53311-7|LNC|Urate crystals|Urate crystals
C2361840|T201|COMP|53312-5|LNC|Calcium carbonate crystals|Calcium carbonate crystals
C2361841|T201|COMP|53313-3|LNC|Cystine crystals|Cystine crystals
C2361842|T201|COMP|53314-1|LNC|Tyrosine crystals|Tyrosine crystals
C2361843|T201|COMP|53323-2|LNC|Casts type not specified|Casts type not specified
C2361844|T201|COMP|53324-0|LNC|Spermatozoa|Spermatozoa
C2361845|T201|COMP|53325-7|LNC|Urinalysis type of crystal panel|Urinalysis type of crystal panel
C2361846|T201|COMP|53326-5|LNC|Specific gravity|Specific gravity
C2361847|T201|COMP|53327-3|LNC|Bilirubin|Bilirubin
C2361848|T201|COMP|53328-1|LNC|Glucose|Glucose
C2361849|T201|COMP|53329-9|LNC|Crystals.amorphous|Crystals.amorphous
C2361851|T201|COMP|53330-7|LNC|Urinalysis type of cast panel|Urinalysis type of cast panel
C2361852|T201|COMP|53331-5|LNC|Crystals.amorphous|Crystals.amorphous
C2361853|T201|COMP|53332-3|LNC|Crystals.amorphous|Crystals.amorphous
C2361854|T201|COMP|53333-1|LNC|Urinalysis other formed elements panel|Urinalysis other formed elements panel
C2361856|T201|COMP|53334-9|LNC|Crystals unspecified|Crystals unspecified
C2361857|T201|COMP|53335-6|LNC|Casts type not specified|Casts type not specified
C2361858|T201|COMP|53336-4|LNC|17-Hydroxyprogesterone+Androstenedione/Cortisol|17-Hydroxyprogesterone+Androstenedione/Cortisol
C2361860|T201|COMP|53337-2|LNC|17-Hydroxyprogesterone+Androstenedione/Cortisol|17-Hydroxyprogesterone+Androstenedione/Cortisol
C2361861|T201|COMP|53338-0|LNC|11-Deoxycortisol|11-Deoxycortisol
C2361862|T201|COMP|53339-8|LNC|11-Deoxycortisol|11-Deoxycortisol
C2361863|T201|COMP|53340-6|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C2361864|T201|COMP|53341-4|LNC|21-Deoxycortisol|21-Deoxycortisol
C2361865|T201|COMP|53342-2|LNC|21-Deoxycortisol|21-Deoxycortisol
C2361866|T201|COMP|53343-0|LNC|Androstenedione|Androstenedione
C2361867|T201|COMP|53344-8|LNC|Androstenedione|Androstenedione
C2361868|T201|COMP|53345-5|LNC|Cortisol|Cortisol
C2361869|T201|COMP|53346-3|LNC|Cortisol|Cortisol
C2361870|T201|COMP|53347-1|LNC|11-Deoxycorticosterone|11-Deoxycorticosterone
C2361871|T201|COMP|53348-9|LNC|11-Deoxycorticosterone|11-Deoxycorticosterone
C2361872|T201|COMP|53349-7|LNC|Thyroxine.free|Thyroxine.free
C2361873|T201|COMP|53350-5|LNC|Thyroxine.free|Thyroxine.free
C2361874|T201|COMP|53351-3|LNC|Urinalysis other formed elements panel|Urinalysis other formed elements panel
C2361875|T201|COMP|53352-1|LNC|Oval fat bodies (globules)|Oval fat bodies (globules)
C2361876|T201|COMP|53353-9|LNC|Urinalysis other formed elements panel|Urinalysis other formed elements panel
C2361877|T201|COMP|53354-7|LNC|Oval fat bodies (globules)|Oval fat bodies (globules)
C2361878|T201|COMP|53355-4|LNC|Trichomonas sp|Trichomonas sp
C2361880|T201|COMP|53357-0|LNC|Trichomonas sp|Trichomonas sp
C2361881|T201|COMP|53358-8|LNC|Erythrocyte clumps|Erythrocyte clumps
C2361883|T201|COMP|53360-4|LNC|Erythrocyte clumps|Erythrocyte clumps
C2361884|T201|COMP|53361-2|LNC|Bordetella parapertussis Ab.IgG|Bordetella parapertussis Ab.IgG
C2361885|T201|COMP|53362-0|LNC|Borrelia burgdorferi 49736 Ab.IgA|Borrelia burgdorferi 49736 Ab.IgA
C2361886|T201|COMP|53363-8|LNC|Borrelia burgdorferi 49736 Ab.IgG|Borrelia burgdorferi 49736 Ab.IgG
C2361887|T201|COMP|53364-6|LNC|Borrelia burgdorferi 49736 Ab.IgM|Borrelia burgdorferi 49736 Ab.IgM
C2361888|T201|COMP|53367-9|LNC|Coccidioides sp Ab.IgM|Coccidioides sp Ab.IgM
C2361889|T201|COMP|53368-7|LNC|Colorado tick fever virus Ab|Colorado tick fever virus Ab
C2361890|T201|COMP|53369-5|LNC|Echinococcus sp Ab.IgG1|Echinococcus sp Ab.IgG1
C2361891|T201|COMP|53370-3|LNC|Echinococcus sp Ab.IgG4|Echinococcus sp Ab.IgG4
C2361892|T201|COMP|53371-1|LNC|Echovirus Ab.IgG|Echovirus Ab.IgG
C2361893|T201|COMP|53372-9|LNC|Echovirus Ab.IgM|Echovirus Ab.IgM
C2361894|T201|COMP|53373-7|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C2361895|T201|COMP|53374-5|LNC|Francisella tularensis Ab|Francisella tularensis Ab
C2361896|T201|COMP|53376-0|LNC|Hepatitis C virus Ab.IgM|Hepatitis C virus Ab.IgM
C2361897|T201|COMP|53377-8|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C2361898|T201|COMP|53378-6|LNC|Herpes virus 6 Ab|Herpes virus 6 Ab
C2361899|T201|COMP|53379-4|LNC|HIV 1 Ab|HIV 1 Ab
C2361900|T201|COMP|53381-0|LNC|Influenza virus A Ab|Influenza virus A Ab
C2361901|T201|COMP|53382-8|LNC|Plasmodium falciparum Ab.IgM|Plasmodium falciparum Ab.IgM
C2361902|T201|COMP|53383-6|LNC|Plasmodium sp Ab.IgG|Plasmodium sp Ab.IgG
C2361903|T201|COMP|53384-4|LNC|Powassan virus Ab|Powassan virus Ab
C2361904|T201|COMP|53385-1|LNC|Snowshoe hare virus Ab|Snowshoe hare virus Ab
C2361905|T201|COMP|53386-9|LNC|Toxocara canis Ab|Toxocara canis Ab
C2361906|T201|COMP|53387-7|LNC|Trichinella spiralis Ab.IgG|Trichinella spiralis Ab.IgG
C2361907|T201|COMP|53388-5|LNC|Trichothecene Ab.IgA|Trichothecene Ab.IgA
C2361908|T201|COMP|53389-3|LNC|Trichothecene Ab.IgE|Trichothecene Ab.IgE
C2361909|T201|COMP|53390-1|LNC|Trichothecene Ab.IgG|Trichothecene Ab.IgG
C2363247|T201|COMP|779-9|LNC|Poikilocytosis|Poikilocytosis
C2363248|T201|COMP|35260-9|LNC|Histamine|Histamine
C2363249|T201|COMP|35213-8|LNC|Insulin-like growth factor-I|Insulin-like growth factor-I
C2363250|T201|COMP|35214-6|LNC|Iron|Iron
C2363251|T201|COMP|35215-3|LNC|Iron binding capacity|Iron binding capacity
C2363252|T201|COMP|35216-1|LNC|Iron binding capacity.unsaturated|Iron binding capacity.unsaturated
C2363253|T201|COMP|35217-9|LNC|Triglyceride|Triglyceride
C2363254|T201|COMP|35218-7|LNC|Osteocalcin|Osteocalcin
C2363255|T201|COMP|35219-5|LNC|Parathyrin.intact|Parathyrin.intact
C2363256|T201|COMP|35220-3|LNC|Phosphate|Phosphate
C2363257|T201|COMP|35222-9|LNC|Phosphate|Phosphate
C2363258|T201|COMP|35263-3|LNC|Phosphate|Phosphate
C2363259|T201|COMP|35223-7|LNC|Progesterone|Progesterone
C2363260|T201|COMP|35224-5|LNC|Testosterone|Testosterone
C2363261|T201|COMP|35225-2|LNC|Testosterone.free|Testosterone.free
C2363262|T201|COMP|35227-8|LNC|Thyroxine binding globulin|Thyroxine binding globulin
C2363263|T201|COMP|35228-6|LNC|Thyroxine.free|Thyroxine.free
C2363264|T201|COMP|35226-0|LNC|Thyroxine|Thyroxine
C2363265|T201|COMP|35229-4|LNC|Transferrin|Transferrin
C2363266|T201|COMP|35230-2|LNC|Triiodothyronine.free|Triiodothyronine.free
C2363267|T201|COMP|35231-0|LNC|Triiodothyronine|Triiodothyronine
C2363268|T201|COMP|35233-6|LNC|Urate|Urate
C2363269|T201|COMP|42571-0|LNC|Urea|Urea
C2363270|T201|COMP|35235-1|LNC|Urea nitrogen|Urea nitrogen
C2363271|T201|COMP|35236-9|LNC|Urobilinogen|Urobilinogen
C2363272|T201|COMP|3213-6|LNC|Coagulation factor VIII Ag|Coagulation factor VIII Ag
C2363273|T201|COMP|17878-0|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C2363274|T201|COMP|35243-5|LNC|Cholesterol.in HDL 3|Cholesterol.in HDL 3
C2363275|T201|COMP|10398-6|LNC|I Ag|I Ag
C2363284|T201|COMP|40572-0|LNC|Neutrophils.band form|Neutrophils.band form
C2363285|T201|COMP|35221-1|LNC|Phosphate|Phosphate
C2363286|T201|COMP|35232-8|LNC|Urate|Urate
C2363327|T201|COMP|26513-2|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C2363333|T201|COMP|41197-5|LNC|Xylose^30M post dose xylose PO|Xylose^30M post dose xylose PO
C2363338|T201|COMP|31113-4|LNC|Cells.HLA-DR+/100 cells|Cells.HLA-DR+/100 cells
C2363356|T201|COMP|41068-8|LNC|PRF1 gene targeted mutation analysis|PRF1 gene targeted mutation analysis
C2363357|T201|COMP|41061-3|LNC|SDHD gene targeted mutation analysis|SDHD gene targeted mutation analysis
C2363358|T201|COMP|41075-3|LNC|NPHS1 gene targeted mutation analysis|NPHS1 gene targeted mutation analysis
C2363359|T201|COMP|41052-2|LNC|SPAST gene targeted mutation analysis|SPAST gene targeted mutation analysis
C2363360|T201|COMP|41054-8|LNC|SMA@ gene mutation analysis|SMA@ gene mutation analysis
C2363361|T201|COMP|35245-0|LNC|Lactate|Lactate
C2363362|T201|COMP|35253-4|LNC|Urate|Urate
C2363363|T201|COMP|35256-7|LNC|Iron|Iron
C2363364|T201|COMP|35259-1|LNC|Neopterin|Neopterin
C2363372|T201|COMP|41048-0|LNC|TPMT gene targeted mutation analysis|TPMT gene targeted mutation analysis
C2363374|T201|COMP|41094-4|LNC|LAMA2 gene targeted mutation analysis|LAMA2 gene targeted mutation analysis
C2363391|T201|COMP|42569-4|LNC|Potassium|Potassium
C2587195|T201|COMP|10399-4|LNC|I Ag|I Ag
C2598065|T201|COMP|53432-1|LNC|Gamma glutamyl transferase|Gamma glutamyl transferase
C2598066|T201|COMP|53433-9|LNC|Creatine kinase|Creatine kinase
C2598067|T201|COMP|53434-7|LNC|Carnitine palmitoyltransferase 2|Carnitine palmitoyltransferase 2
C2598069|T201|COMP|53435-4|LNC|Argininosuccinate lyase|Argininosuccinate lyase
C2598070|T201|COMP|53436-2|LNC|Carnitine palmitoyltransferase 2|Carnitine palmitoyltransferase 2
C2598071|T201|COMP|53437-0|LNC|Carnitine palmitoyltransferase 1|Carnitine palmitoyltransferase 1
C2598072|T201|COMP|53438-8|LNC|Carnitine palmitoyltransferase 2|Carnitine palmitoyltransferase 2
C2598073|T201|COMP|53926-2|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C2598074|T201|COMP|53927-0|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2598075|T201|COMP|53928-8|LNC|Glucose^20M post 50 g lactose PO|Glucose^20M post 50 g lactose PO
C2598076|T201|COMP|53929-6|LNC|Glucose^40M post 50 g lactose PO|Glucose^40M post 50 g lactose PO
C2598077|T201|COMP|53930-4|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C2598078|T201|COMP|53931-2|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C2598096|T201|COMP|53462-8|LNC|Eicosanoylcarnitine (C20)|Eicosanoylcarnitine (C20)
C2598097|T201|COMP|53463-6|LNC|Beta aminoisobutyrate|Beta aminoisobutyrate
C2598098|T201|COMP|53464-4|LNC|Decadienoylcarnitine (C10:2)|Decadienoylcarnitine (C10:2)
C2598099|T201|COMP|53465-1|LNC|Sebacylcarnitine (C10-DC)|Sebacylcarnitine (C10-DC)
C2598100|T201|COMP|53466-9|LNC|Eicosanoylcarnitine (C20)|Eicosanoylcarnitine (C20)
C2598101|T201|COMP|53467-7|LNC|3-Keto n-Valerate|3-Keto n-Valerate
C2598102|T201|COMP|53468-5|LNC|Anthranilate|Anthranilate
C2598103|T201|COMP|53469-3|LNC|Kynurenate|Kynurenate
C2598404|T201|COMP|53553-4|LNC|Estimated average glucose|Estimated average glucose
C2598405|T201|COMP|53554-2|LNC|Nitrogen|Nitrogen
C2598406|T201|COMP|53555-9|LNC|Specific gravity|Specific gravity
C2598409|T201|COMP|53557-5|LNC|Nucleated cells|Nucleated cells
C2598410|T201|COMP|53558-3|LNC|Bacteria identified|Bacteria identified
C2598411|T201|COMP|53559-1|LNC|Beta-2 transferrin|Beta-2 transferrin
C2598412|T201|COMP|53560-9|LNC|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C2598413|T201|COMP|53561-7|LNC|Lactate dehydrogenase/Creatinine|Lactate dehydrogenase/Creatinine
C2598415|T201|COMP|53562-5|LNC|Rheumatoid factor|Rheumatoid factor
C2598441|T201|COMP|53415-6|LNC|Bilirubin|Bilirubin
C2598442|T201|COMP|53416-4|LNC|Alpha naphthylesterase|Alpha naphthylesterase
C2598443|T201|COMP|53417-2|LNC|Alpha naphthylesterase|Alpha naphthylesterase
C2598451|T201|COMP|53425-5|LNC|Fibroblast growth factor 23 ^pre XXX challenge|Fibroblast growth factor 23 ^pre XXX challenge
C2598459|T201|COMP|53447-9|LNC|Carboxymefloquine|Carboxymefloquine
C2598460|T201|COMP|53448-7|LNC|Cycloguanil|Cycloguanil
C2598461|T201|COMP|53449-5|LNC|Cyclophosphamide|Cyclophosphamide
C2598462|T201|COMP|53450-3|LNC|Cytarabine|Cytarabine
C2598464|T201|COMP|53451-1|LNC|Uracil arabinoside|Uracil arabinoside
C2598466|T201|COMP|53452-9|LNC|Gamma 3 globulin.abnormal band|Gamma 3 globulin.abnormal band
C2598468|T201|COMP|53453-7|LNC|Cyclophosphamide|Cyclophosphamide
C2598469|T201|COMP|53454-5|LNC|Iron^post dose deferoxamine|Iron^post dose deferoxamine
C2598471|T201|COMP|53745-6|LNC|Benzodiazepines panel|Benzodiazepines panel
C2598473|T201|COMP|53746-4|LNC|Barbiturates panel|Barbiturates panel
C2598475|T201|COMP|53747-2|LNC|Cocaine panel|Cocaine panel
C2598478|T201|COMP|53749-8|LNC|Collection time^5th specimen|Collection time^5th specimen
C2598479|T201|COMP|53750-6|LNC|Hydrogen/Expired gas^15M post XXX challenge|Hydrogen/Expired gas^15M post XXX challenge
C2598480|T201|COMP|53751-4|LNC|Hydrogen/Expired gas^2.75H post XXX challenge|Hydrogen/Expired gas^2.75H post XXX challenge
C2598481|T201|COMP|53752-2|LNC|Hydrogen/Expired gas^1.75H post XXX challenge|Hydrogen/Expired gas^1.75H post XXX challenge
C2598482|T201|COMP|53753-0|LNC|Hydrogen/Expired gas^2.25H post XXX challenge|Hydrogen/Expired gas^2.25H post XXX challenge
C2598483|T201|COMP|53754-8|LNC|Hydrogen/Expired gas^45M post XXX challenge|Hydrogen/Expired gas^45M post XXX challenge
C2598484|T201|COMP|53755-5|LNC|Hydrogen/Expired gas^1.25H post XXX challenge|Hydrogen/Expired gas^1.25H post XXX challenge
C2598486|T201|COMP|53758-9|LNC|HLA-DRB1 SBT|HLA-DRB1 SBT
C2598487|T201|COMP|53759-7|LNC|Natural killer cell panel|Natural killer cell panel
C2598489|T201|COMP|53760-5|LNC|Cladosporium sp Ab.IgE|Cladosporium sp Ab.IgE
C2598490|T201|COMP|53958-5|LNC|Choriogonadotropin.tumor marker|Choriogonadotropin.tumor marker
C2598492|T201|COMP|53959-3|LNC|Choriogonadotropin.tumor marker|Choriogonadotropin.tumor marker
C2598493|T201|COMP|53960-1|LNC|Alpha-1-Fetoprotein.tumor marker|Alpha-1-Fetoprotein.tumor marker
C2598495|T201|COMP|53961-9|LNC|Alpha-1-Fetoprotein.tumor marker|Alpha-1-Fetoprotein.tumor marker
C2598496|T201|COMP|53962-7|LNC|Alpha-1-Fetoprotein.tumor marker|Alpha-1-Fetoprotein.tumor marker
C2598497|T201|COMP|53963-5|LNC|Blood|Blood
C2598498|T201|COMP|53964-3|LNC|Leukocytes|Leukocytes
C2598499|T201|COMP|53965-0|LNC|Brickdust deposit|Brickdust deposit
C2598500|T201|COMP|53966-8|LNC|Erythrocytes.dysmorphic G1/100 erythrocytes|Erythrocytes.dysmorphic G1/100 erythrocytes
C2598502|T201|COMP|53967-6|LNC|Erythrocytes.dysmorphic/100 erythrocytes|Erythrocytes.dysmorphic/100 erythrocytes
C2598504|T201|COMP|53968-4|LNC|Erythrocytes.non-dysmorphic|Erythrocytes.non-dysmorphic
C2598505|T201|COMP|53969-2|LNC|Microcytes|Microcytes
C2598506|T201|COMP|53970-0|LNC|Macrocytes|Macrocytes
C2598507|T201|COMP|53971-8|LNC|Spherocytes|Spherocytes
C2598556|T201|COMP|53439-6|LNC|Argininosuccinate lyase|Argininosuccinate lyase
C2598557|T201|COMP|53440-4|LNC|Argininosuccinate synthase|Argininosuccinate synthase
C2598558|T201|COMP|53441-2|LNC|Carnitine palmitoyltransferase 1|Carnitine palmitoyltransferase 1
C2598559|T201|COMP|53442-0|LNC|Carnitine palmitoyltransferase 2|Carnitine palmitoyltransferase 2
C2598560|T201|COMP|53443-8|LNC|Carnitine palmitoyltransferase 2|Carnitine palmitoyltransferase 2
C2598561|T201|COMP|53444-6|LNC|Citrate synthase|Citrate synthase
C2598562|T201|COMP|53445-3|LNC|Carnitine palmitoyltransferase 2/Citrate synthase|Carnitine palmitoyltransferase 2/Citrate synthase
C2598564|T201|COMP|53446-1|LNC|Carnitine palmitoyltransferase 2/Citrate synthase|Carnitine palmitoyltransferase 2/Citrate synthase
C2598565|T201|COMP|53455-2|LNC|Calcium|Calcium
C2598566|T201|COMP|53456-0|LNC|Iron|Iron
C2598567|T201|COMP|53457-8|LNC|Gamma 3 globulin.abnormal band/Protein.total|Gamma 3 globulin.abnormal band/Protein.total
C2598569|T201|COMP|53458-6|LNC|Carbon dioxide|Carbon dioxide
C2598570|T201|COMP|53459-4|LNC|Decadienoylcarnitine (C10:2)|Decadienoylcarnitine (C10:2)
C2598571|T201|COMP|53460-2|LNC|Sebacylcarnitine (C10-DC)|Sebacylcarnitine (C10-DC)
C2598572|T201|COMP|53461-0|LNC|Eicosanoylcarnitine (C20)|Eicosanoylcarnitine (C20)
C2598573|T201|COMP|53470-1|LNC|Kynurenin|Kynurenin
C2598575|T201|COMP|53471-9|LNC|Decadienoylcarnitine (C10:2)|Decadienoylcarnitine (C10:2)
C2598576|T201|COMP|53472-7|LNC|Sebacylcarnitine (C10-DC)|Sebacylcarnitine (C10-DC)
C2598577|T201|COMP|53473-5|LNC|Eicosanoylcarnitine (C20)|Eicosanoylcarnitine (C20)
C2598578|T201|COMP|53474-3|LNC|Glucose^4 AM specimen|Glucose^4 AM specimen
C2598579|T201|COMP|53475-0|LNC|Glucose^pre dose betaxolol|Glucose^pre dose betaxolol
C2598580|T201|COMP|53476-8|LNC|Glucose^2H post dose betaxolol|Glucose^2H post dose betaxolol
C2598581|T201|COMP|53477-6|LNC|Levodopa/Tyrosine|Levodopa/Tyrosine
C2598583|T201|COMP|53478-4|LNC|Anthranilate|Anthranilate
C2598584|T201|COMP|53479-2|LNC|Dihydroxycholestanoate|Dihydroxycholestanoate
C2598585|T201|COMP|53480-0|LNC|Glucose^2.5H post dose betaxolol|Glucose^2.5H post dose betaxolol
C2598586|T201|COMP|53481-8|LNC|Glucose^15M pre dose betaxolol|Glucose^15M pre dose betaxolol
C2598587|T201|COMP|53482-6|LNC|Glucose^3H post dose betaxolol|Glucose^3H post dose betaxolol
C2598588|T201|COMP|53483-4|LNC|Glucose^30M post dose betaxolol|Glucose^30M post dose betaxolol
C2598589|T201|COMP|53484-2|LNC|Glucose^30M pre dose betaxolol|Glucose^30M pre dose betaxolol
C2598590|T201|COMP|53485-9|LNC|Glucose^45M post dose betaxolol|Glucose^45M post dose betaxolol
C2598591|T201|COMP|53486-7|LNC|Glucose^1H post dose betaxolol|Glucose^1H post dose betaxolol
C2598592|T201|COMP|53487-5|LNC|Glucose^1.5H post dose betaxolol|Glucose^1.5H post dose betaxolol
C2598593|T201|COMP|53488-3|LNC|3-O-Methyldopa|3-O-Methyldopa
C2598594|T201|COMP|53489-1|LNC|Kynurenate|Kynurenate
C2598595|T201|COMP|53490-9|LNC|Kynurenin|Kynurenin
C2598596|T201|COMP|53491-7|LNC|Kynurenin|Kynurenin
C2598597|T201|COMP|53492-5|LNC|Decadienoylcarnitine (C10:2)|Decadienoylcarnitine (C10:2)
C2598598|T201|COMP|53493-3|LNC|Sebacylcarnitine (C10-DC)|Sebacylcarnitine (C10-DC)
C2598599|T201|COMP|53494-1|LNC|Eicosanoylcarnitine (C20)|Eicosanoylcarnitine (C20)
C2598600|T201|COMP|53495-8|LNC|Iron^post dose deferoxamine|Iron^post dose deferoxamine
C2598601|T201|COMP|53496-6|LNC|3-Methoxy-4-Hydroxyphenylglycol|3-Methoxy-4-Hydroxyphenylglycol
C2598602|T201|COMP|53497-4|LNC|5-Hydroxytryptophan|5-Hydroxytryptophan
C2598603|T201|COMP|53498-2|LNC|Anthranilate|Anthranilate
C2598604|T201|COMP|53499-0|LNC|Creatinine|Creatinine
C2598605|T201|COMP|53500-5|LNC|Ammonia|Ammonia
C2598606|T201|COMP|53501-3|LNC|Iron|Iron
C2598607|T201|COMP|53502-1|LNC|Calcium|Calcium
C2598608|T201|COMP|53503-9|LNC|Iron|Iron
C2598609|T201|COMP|53504-7|LNC|Decanoylcarnitine (C10)/Creatinine|Decanoylcarnitine (C10)/Creatinine
C2598611|T201|COMP|53505-4|LNC|Asparagine/Amino acids.total|Asparagine/Amino acids.total
C2598613|T201|COMP|53506-2|LNC|Citrulline/Amino acids.total|Citrulline/Amino acids.total
C2598615|T201|COMP|53507-0|LNC|Kynurenin/Creatinine|Kynurenin/Creatinine
C2598617|T201|COMP|53508-8|LNC|Decadienoylcarnitine (C10:2)/Creatinine|Decadienoylcarnitine (C10:2)/Creatinine
C2598618|T201|COMP|53509-6|LNC|Sebacylcarnitine (C10-DC)/Creatinine|Sebacylcarnitine (C10-DC)/Creatinine
C2598620|T201|COMP|53510-4|LNC|Dodecanoylcarnitine (C12)/Creatinine|Dodecanoylcarnitine (C12)/Creatinine
C2598622|T201|COMP|53511-2|LNC|Dodecenoylcarnitine (C12:1)/Creatinine|Dodecenoylcarnitine (C12:1)/Creatinine
C2598624|T201|COMP|53512-0|LNC|Eicosanoylcarnitine (C20)/Creatinine|Eicosanoylcarnitine (C20)/Creatinine
C2598626|T201|COMP|53513-8|LNC|Anthranilate/Creatinine|Anthranilate/Creatinine
C2598628|T201|COMP|53514-6|LNC|Carnitine palmitoyltransferase 2|Carnitine palmitoyltransferase 2
C2598629|T201|COMP|53515-3|LNC|Citrate synthase|Citrate synthase
C2598630|T201|COMP|53516-1|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C2598631|T201|COMP|53517-9|LNC|Erythrocytes|Erythrocytes
C2598632|T201|COMP|53518-7|LNC|Leukocytes|Leukocytes
C2598633|T201|COMP|53519-5|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C2598634|T201|COMP|53520-3|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C2598635|T201|COMP|53521-1|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C2598637|T201|COMP|53523-7|LNC|Vasoactive intestinal peptide|Vasoactive intestinal peptide
C2598640|T201|COMP|53525-2|LNC|Protein|Protein
C2598641|T201|COMP|53526-0|LNC|Triglyceride.in VLDL|Triglyceride.in VLDL
C2598643|T201|COMP|53527-8|LNC|Triglyceride.in HDL 2|Triglyceride.in HDL 2
C2598645|T201|COMP|53528-6|LNC|Triglyceride.in HDL 3|Triglyceride.in HDL 3
C2598647|T201|COMP|53529-4|LNC|Albumin|Albumin
C2598648|T201|COMP|53530-2|LNC|Albumin|Albumin
C2598649|T201|COMP|53531-0|LNC|Albumin|Albumin
C2598650|T201|COMP|53532-8|LNC|Albumin|Albumin
C2598651|T201|COMP|53533-6|LNC|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C2598652|T201|COMP|53534-4|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C2598653|T201|COMP|53535-1|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C2598654|T201|COMP|53536-9|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C2598655|T201|COMP|53537-7|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C2598656|T201|COMP|53538-5|LNC|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C2598657|T201|COMP|53539-3|LNC|Alpha globulin.abnormal band|Alpha globulin.abnormal band
C2598659|T201|COMP|53540-1|LNC|Alpha globulin.abnormal band/Protein.total|Alpha globulin.abnormal band/Protein.total
C2598661|T201|COMP|53541-9|LNC|Epithelial cells|Epithelial cells
C2598662|T201|COMP|53542-7|LNC|Dodeicosanoylcarnitine (C22)|Dodeicosanoylcarnitine (C22)
C2598664|T201|COMP|53543-5|LNC|Dodeicosanoylcarnitine (C22)|Dodeicosanoylcarnitine (C22)
C2598665|T201|COMP|53544-3|LNC|3,4-Dihydroxyphenylacetate|3,4-Dihydroxyphenylacetate
C2598666|T201|COMP|53545-0|LNC|Dodeicosanoylcarnitine (C22)|Dodeicosanoylcarnitine (C22)
C2598667|T201|COMP|53546-8|LNC|Dodeicosanoylcarnitine (C22)|Dodeicosanoylcarnitine (C22)
C2598668|T201|COMP|53547-6|LNC|3,4-Dihydroxyphenylacetate|3,4-Dihydroxyphenylacetate
C2598669|T201|COMP|53548-4|LNC|3,4-Dihydroxyphenylacetate|3,4-Dihydroxyphenylacetate
C2598670|T201|COMP|53549-2|LNC|Dodeicosanoylcarnitine (C22)|Dodeicosanoylcarnitine (C22)
C2598671|T201|COMP|53550-0|LNC|Fructosamine/Protein|Fructosamine/Protein
C2598673|T201|COMP|53551-8|LNC|3,4-Dihydroxyphenylacetate/Creatinine|3,4-Dihydroxyphenylacetate/Creatinine
C2598675|T201|COMP|53552-6|LNC|Dodeicosanoylcarnitine (C22)/Creatinine|Dodeicosanoylcarnitine (C22)/Creatinine
C2598679|T201|COMP|53566-6|LNC|Platelet aggregation.collagen induced^8.0 ug/mL|Platelet aggregation.collagen induced^8.0 ug/mL
C2598682|T201|COMP|53569-0|LNC|Platelet aggregation.ristocetin induced^800 ug/mL|Platelet aggregation.ristocetin induced^800 ug/mL
C2598683|T201|COMP|53570-8|LNC|Coagulation surface induced.lupus insensitive|Coagulation surface induced.lupus insensitive
C2598685|T201|COMP|53571-6|LNC|Yeast identified|Yeast identified
C2598688|T201|COMP|53573-2|LNC|cycloSPORINE^post dose|cycloSPORINE^post dose
C2598689|T201|COMP|53574-0|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C2598690|T201|COMP|53575-7|LNC|VAP panel|VAP panel
C2598694|T201|COMP|53577-3|LNC|Reason for study additional note|Reason for study additional note
C2598700|T201|COMP|53580-7|LNC|Galactosylceramidase|Galactosylceramidase
C2598701|T201|COMP|53581-5|LNC|Angiotensin converting enzyme|Angiotensin converting enzyme
C2598702|T201|COMP|53582-3|LNC|Echovirus Ab|Echovirus Ab
C2598703|T201|COMP|53583-1|LNC|Echovirus Ab.IgM|Echovirus Ab.IgM
C2598704|T201|COMP|53584-9|LNC|Loa loa DNA|Loa loa DNA
C2598706|T201|COMP|53585-6|LNC|Toxocara canis Ab.IgE|Toxocara canis Ab.IgE
C2598708|T201|COMP|53586-4|LNC|HLA-B6|HLA-B6
C2598710|T201|COMP|53587-2|LNC|Beta globulin.abnormal band|Beta globulin.abnormal band
C2598712|T201|COMP|53588-0|LNC|Beta globulin+Gamma globulin.abnormal band|Beta globulin+Gamma globulin.abnormal band
C2598714|T201|COMP|53589-8|LNC|Beta globulin.abnormal band/Protein.total|Beta globulin.abnormal band/Protein.total
C2598716|T201|COMP|53590-6|LNC|Gamma globulin.abnormal band/Protein.total|Gamma globulin.abnormal band/Protein.total
C2598718|T201|COMP|53591-4|LNC|Gamma globulin.abnormal band|Gamma globulin.abnormal band
C2598720|T201|COMP|53592-2|LNC|Gamma 2 globulin.abnormal band|Gamma 2 globulin.abnormal band
C2598722|T201|COMP|53593-0|LNC|Gamma 2 globulin.abnormal band/Protein.total|Gamma 2 globulin.abnormal band/Protein.total
C2598724|T201|COMP|53594-8|LNC|Chitobioside Ab.IgA|Chitobioside Ab.IgA
C2598726|T201|COMP|53595-5|LNC|Homovanillate|Homovanillate
C2598727|T201|COMP|53596-3|LNC|Laminaribioside Ab.IgG|Laminaribioside Ab.IgG
C2598729|T201|COMP|53597-1|LNC|Mannobioside Ab.IgG|Mannobioside Ab.IgG
C2598731|T201|COMP|53598-9|LNC|Irritable bowel disease prognostic panel|Irritable bowel disease prognostic panel
C2598736|T201|COMP|53601-1|LNC|HIV 1 p24 Ag|HIV 1 p24 Ag
C2598737|T201|COMP|53602-9|LNC|Taenia solium larva Ag|Taenia solium larva Ag
C2598739|T201|COMP|53603-7|LNC|Mumps virus RNA|Mumps virus RNA
C2598740|T201|COMP|53604-5|LNC|Brucella sp DNA|Brucella sp DNA
C2598741|T201|COMP|53605-2|LNC|Treponema pallidum DNA|Treponema pallidum DNA
C2598742|T201|COMP|53606-0|LNC|Neisseria meningitidis DNA|Neisseria meningitidis DNA
C2598743|T201|COMP|53607-8|LNC|Haemophilus influenzae B DNA|Haemophilus influenzae B DNA
C2598744|T201|COMP|53608-6|LNC|Rickettsia sp DNA|Rickettsia sp DNA
C2598745|T201|COMP|53609-4|LNC|Parasite identified|Parasite identified
C2598746|T201|COMP|53610-2|LNC|Erythroid cells|Erythroid cells
C2598747|T201|COMP|53611-0|LNC|Toxoplasma gondii|Toxoplasma gondii
C2598748|T201|COMP|53612-8|LNC|Urate|Urate
C2598749|T201|COMP|53613-6|LNC|Benzoylcarnitine (BzCn)|Benzoylcarnitine (BzCn)
C2598750|T201|COMP|53614-4|LNC|Bacteria identified^^^2|Bacteria identified^^^2
C2598751|T201|COMP|53615-1|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C2598752|T201|COMP|53616-9|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C2598753|T201|COMP|53617-7|LNC|Bacteria identified|Bacteria identified
C2598754|T201|COMP|53618-5|LNC|Cells.ZAP70|Cells.ZAP70
C2598755|T201|COMP|53619-3|LNC|Cells.ZAP70|Cells.ZAP70
C2598756|T201|COMP|53620-1|LNC|KRAS gene targeted mutation analysis|KRAS gene targeted mutation analysis
C2598757|T201|COMP|53621-9|LNC|NRAS gene targeted mutation analysis|NRAS gene targeted mutation analysis
C2598760|T201|COMP|53623-5|LNC|HRAS gene targeted mutation analysis|HRAS gene targeted mutation analysis
C2598761|T201|COMP|53624-3|LNC|Carnitine esters|Carnitine esters
C2598762|T201|COMP|53625-0|LNC|Leishmania sp identified|Leishmania sp identified
C2598765|T201|COMP|53627-6|LNC|Chloride|Chloride
C2598766|T201|COMP|53628-4|LNC|20q chromosome deletion|20q chromosome deletion
C2598768|T201|COMP|53776-1|LNC|Hepatitis A virus Ab.IgM & total|Hepatitis A virus Ab.IgM & total
C2598770|T201|COMP|53777-9|LNC|Cortisone.free|Cortisone.free
C2598771|T201|COMP|53778-7|LNC|Arsenic.organic|Arsenic.organic
C2598772|T201|COMP|53779-5|LNC|Arsenic.methylated|Arsenic.methylated
C2598774|T201|COMP|53780-3|LNC|Chromium panel|Chromium panel
C2598776|T201|COMP|53781-1|LNC|Acetaminophen & Propoxyphene panel|Acetaminophen & Propoxyphene panel
C2598778|T201|COMP|53782-9|LNC|HTT gene.CAG repeats|HTT gene.CAG repeats
C2598779|T201|COMP|53783-7|LNC|HTT gene mutation panel|HTT gene mutation panel
C2598781|T201|COMP|53784-5|LNC|Legionella pneumophila 1+2+3+4+5+6 Ab.IgM|Legionella pneumophila 1+2+3+4+5+6 Ab.IgM
C2598784|T201|COMP|53787-8|LNC|Zolpidem|Zolpidem
C2598785|T201|COMP|53788-6|LNC|Sodium urate crystals|Sodium urate crystals
C2598786|T201|COMP|53789-4|LNC|CFTR gene.p.IVS8 polyT 7T/9T variant|CFTR gene.p.IVS8 polyT 7T/9T variant
C2598788|T201|COMP|53790-2|LNC|CILD2 gene targeted mutation analysis|CILD2 gene targeted mutation analysis
C2598790|T201|COMP|53877-7|LNC|NAGS gene targeted mutation analysis|NAGS gene targeted mutation analysis
C2598792|T201|COMP|53878-5|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2598793|T201|COMP|53879-3|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2598794|T201|COMP|53880-1|LNC|Norbuprenorphine|Norbuprenorphine
C2598795|T201|COMP|53881-9|LNC|Norbuprenorphine|Norbuprenorphine
C2598796|T201|COMP|53882-7|LNC|Norvenlafaxine|Norvenlafaxine
C2598797|T201|COMP|53883-5|LNC|OCRL1 gene targeted mutation analysis|OCRL1 gene targeted mutation analysis
C2598799|T201|COMP|53884-3|LNC|OTOF gene targeted mutation analysis|OTOF gene targeted mutation analysis
C2598801|T201|COMP|53629-2|LNC|Alpha cortol|Alpha cortol
C2598802|T201|COMP|53630-0|LNC|Alpha cortol/Creatinine|Alpha cortol/Creatinine
C2598804|T201|COMP|53631-8|LNC|Alpha cortol/Creatinine|Alpha cortol/Creatinine
C2598805|T201|COMP|53632-6|LNC|Breast Cancer Ag 225|Breast Cancer Ag 225
C2598807|T201|COMP|53633-4|LNC|BCL1 Ag|BCL1 Ag
C2598809|T201|COMP|53634-2|LNC|Beta cortol|Beta cortol
C2598810|T201|COMP|53635-9|LNC|Beta cortol/Creatinine|Beta cortol/Creatinine
C2598812|T201|COMP|53636-7|LNC|Beta cortol/Creatinine|Beta cortol/Creatinine
C2598813|T201|COMP|53637-5|LNC|BOB1 Ag|BOB1 Ag
C2598815|T201|COMP|53638-3|LNC|CD45RB Ag|CD45RB Ag
C2598816|T201|COMP|53639-1|LNC|CD52 Ag|CD52 Ag
C2598817|T201|COMP|53640-9|LNC|Chloride/Creatinine|Chloride/Creatinine
C2598818|T201|COMP|53641-7|LNC|OCT2 Ag|OCT2 Ag
C2598820|T201|COMP|53642-5|LNC|Glutathione.reduced/glutathione.oxidized|Glutathione.reduced/glutathione.oxidized
C2598822|T201|COMP|53643-3|LNC|Dichlorodiphenyltrichloroethane|Dichlorodiphenyltrichloroethane
C2598823|T201|COMP|53644-1|LNC|Carbaryl|Carbaryl
C2598824|T201|COMP|53645-8|LNC|Polio virus identified|Polio virus identified
C2598826|T201|COMP|53646-6|LNC|Aldicarb|Aldicarb
C2598827|T201|COMP|53647-4|LNC|Flavin adenine dinucleotide|Flavin adenine dinucleotide
C2598828|T201|COMP|53648-2|LNC|Flavin mononucleotide|Flavin mononucleotide
C2598829|T201|COMP|53649-0|LNC|Parathion|Parathion
C2598830|T201|COMP|53650-8|LNC|Methyl parathion|Methyl parathion
C2598898|T201|COMP|53705-0|LNC|Myasthenia gravis evaluation pediatric panel|Myasthenia gravis evaluation pediatric panel
C2598900|T201|COMP|53706-8|LNC|Myasthenia gravis evaluation adult reflex panel|Myasthenia gravis evaluation adult reflex panel
C2598902|T201|COMP|53707-6|LNC|CV2 Ab.IgG|CV2 Ab.IgG
C2598903|T201|COMP|53708-4|LNC|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C2598904|T201|COMP|53709-2|LNC|Glial nuclear type 1 Ab|Glial nuclear type 1 Ab
C2598906|T201|COMP|53710-0|LNC|Hyperoxaluria panel|Hyperoxaluria panel
C2598908|T201|COMP|53711-8|LNC|Neuronal nuclear type 1 Ab|Neuronal nuclear type 1 Ab
C2598909|T201|COMP|53712-6|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C2598910|T201|COMP|53713-4|LNC|Purkinje cell cytoplasmic type 1 Ab|Purkinje cell cytoplasmic type 1 Ab
C2598912|T201|COMP|53714-2|LNC|Glial nuclear type 1 Ab|Glial nuclear type 1 Ab
C2598913|T201|COMP|53715-9|LNC|Paraneoplastic Ab|Paraneoplastic Ab
C2598914|T201|COMP|53716-7|LNC|levoFLOXacin|levoFLOXacin
C2598915|T201|COMP|53717-5|LNC|Purkinje cell cytoplasmic type 1 Ab|Purkinje cell cytoplasmic type 1 Ab
C2598916|T201|COMP|53718-3|LNC|Acylglycines|Acylglycines
C2598920|T201|COMP|53721-7|LNC|Amino acid marker assessed|Amino acid marker assessed
C2598922|T201|COMP|53722-5|LNC|SLC26A4 gene.p.Glu384Gly|SLC26A4 gene.p.Glu384Gly
C2598924|T201|COMP|53723-3|LNC|SLC26A4 gene.p.Leu236Pro|SLC26A4 gene.p.Leu236Pro
C2598926|T201|COMP|53724-1|LNC|SLC26A4 gene.p.Thr416Pro|SLC26A4 gene.p.Thr416Pro
C2598928|T201|COMP|53725-8|LNC|SLC25A4 gene targeted mutation analysis|SLC25A4 gene targeted mutation analysis
C2598930|T201|COMP|53726-6|LNC|KCNC3 gene targeted mutation analysis|KCNC3 gene targeted mutation analysis
C2598932|T201|COMP|53727-4|LNC|SOS1 gene targeted mutation analysis|SOS1 gene targeted mutation analysis
C2598934|T201|COMP|53728-2|LNC|WS2A gene targeted mutation analysis|WS2A gene targeted mutation analysis
C2598936|T201|COMP|53729-0|LNC|Borrelia burgdorferi 49736 Ab.IgG|Borrelia burgdorferi 49736 Ab.IgG
C2598937|T201|COMP|53730-8|LNC|Borrelia burgdorferi G39_40 Ab.IgG|Borrelia burgdorferi G39_40 Ab.IgG
C2598938|T201|COMP|53731-6|LNC|Posaconazole|Posaconazole
C2598939|T201|COMP|53732-4|LNC|GCK gene targeted mutation analysis|GCK gene targeted mutation analysis
C2598941|T201|COMP|53733-2|LNC|Color|Color
C2598942|T201|COMP|53734-0|LNC|Kynurenine|Kynurenine
C2598943|T201|COMP|53735-7|LNC|Barbiturates.other|Barbiturates.other
C2598945|T201|COMP|53736-5|LNC|Benzodiazepines.other|Benzodiazepines.other
C2598947|T201|COMP|53737-3|LNC|HLA-DQA1*01:02|HLA-DQA1*01:02
C2598949|T201|COMP|53738-1|LNC|HLA-DQB1*2|HLA-DQB1*2
C2598951|T201|COMP|53739-9|LNC|HLA-DQB1*9|HLA-DQB1*9
C2598953|T201|COMP|53740-7|LNC|HLA-DRB1*17|HLA-DRB1*17
C2598955|T201|COMP|53741-5|LNC|HLA-DRB1*7|HLA-DRB1*7
C2598957|T201|COMP|53742-3|LNC|Legionella pneumophila 2+3+4+5+6+8 Ab|Legionella pneumophila 2+3+4+5+6+8 Ab
C2598958|T201|COMP|53743-1|LNC|Cocaine metabolites.other|Cocaine metabolites.other
C2598960|T201|COMP|53761-3|LNC|JAK2 gene.p.Val617Phe mutant/normal|JAK2 gene.p.Val617Phe mutant/normal
C2598962|T201|COMP|53762-1|LNC|Neisseria gonorrhoeae Ab.IgG|Neisseria gonorrhoeae Ab.IgG
C2598964|T201|COMP|53763-9|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C2598965|T201|COMP|53764-7|LNC|Prostate specific Ag panel|Prostate specific Ag panel
C2598967|T201|COMP|53765-4|LNC|Estrogen|Estrogen
C2598968|T201|COMP|53766-2|LNC|Estrogen fraction panel|Estrogen fraction panel
C2598970|T201|COMP|53767-0|LNC|HLA-A+B+C SBT|HLA-A+B+C SBT
C2598971|T201|COMP|53768-8|LNC|Erythrocytes.CD55+CD59 actual/normal|Erythrocytes.CD55+CD59 actual/normal
C2598973|T201|COMP|53769-6|LNC|Erythrocytes.CD55+CD59 deficient actual/normal|Erythrocytes.CD55+CD59 deficient actual/normal
C2598975|T201|COMP|53770-4|LNC|Legionella pneumophila 1+2+3+4+5+6 Ab.IgG|Legionella pneumophila 1+2+3+4+5+6 Ab.IgG
C2598977|T201|COMP|53771-2|LNC|Alpha 2 globulin|Alpha 2 globulin
C2598978|T201|COMP|53772-0|LNC|Beta globulin|Beta globulin
C2598979|T201|COMP|53773-8|LNC|Gamma globulin|Gamma globulin
C2598980|T201|COMP|53774-6|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C2598981|T201|COMP|53775-3|LNC|Hepatitis A virus Ab panel|Hepatitis A virus Ab panel
C2598983|T201|COMP|53791-0|LNC|PTPN11 gene targeted mutation analysis.tier 1|PTPN11 gene targeted mutation analysis.tier 1
C2598985|T201|COMP|53792-8|LNC|PTPN11 gene targeted mutation analysis.tier 3|PTPN11 gene targeted mutation analysis.tier 3
C2598987|T201|COMP|53793-6|LNC|RPS6KA3 gene targeted mutation analysis.tier 1|RPS6KA3 gene targeted mutation analysis.tier 1
C2598989|T201|COMP|53794-4|LNC|RPS6KA3 gene targeted mutation analysis.tier 2|RPS6KA3 gene targeted mutation analysis.tier 2
C2598991|T201|COMP|53795-1|LNC|STK11 gene targeted mutation analysis|STK11 gene targeted mutation analysis
C2598993|T201|COMP|53796-9|LNC|Interferon drug given|Interferon drug given
C2598995|T201|COMP|53797-7|LNC|Neutrophils.immature/100 leukocytes|Neutrophils.immature/100 leukocytes
C2598999|T201|COMP|53799-3|LNC|Major crossmatch|Major crossmatch
C2599000|T201|COMP|53800-9|LNC|Platelets panel|Platelets panel
C2599003|T201|COMP|53802-5|LNC|Arbovirus Ab.IgG|Arbovirus Ab.IgG
C2599004|T201|COMP|53803-3|LNC|Transferrin.carbohydrate deficient panel|Transferrin.carbohydrate deficient panel
C2599006|T201|COMP|53804-1|LNC|Arbovirus Ab.IgG panel|Arbovirus Ab.IgG panel
C2599008|T201|COMP|53805-8|LNC|LDL apheresis procedure|LDL apheresis procedure
C2599010|T201|COMP|53806-6|LNC|LDL apheresis procedure|LDL apheresis procedure
C2599011|T201|COMP|53807-4|LNC|Basement membrane zone BP230 Ab.IgG|Basement membrane zone BP230 Ab.IgG
C2599013|T201|COMP|53808-2|LNC|Oligosaccharides pattern|Oligosaccharides pattern
C2599015|T201|COMP|53810-8|LNC|Lymphocyte proliferation|Lymphocyte proliferation
C2599016|T201|COMP|53811-6|LNC|Triple phosphate|Triple phosphate
C2599017|T201|COMP|53812-4|LNC|Micafungin|Micafungin
C2599019|T201|COMP|53814-0|LNC|Platelet aggregation.arachidonate induced|Platelet aggregation.arachidonate induced
C2599020|T201|COMP|53815-7|LNC|Platelet glycoprotein IIb-IIIa Ab|Platelet glycoprotein IIb-IIIa Ab
C2599021|T201|COMP|53816-5|LNC|Alpha hydroxytriazolam|Alpha hydroxytriazolam
C2599022|T201|COMP|53817-3|LNC|Carnosine|Carnosine
C2599023|T201|COMP|53818-1|LNC|Arbekacin|Arbekacin
C2599024|T201|COMP|53819-9|LNC|Thiopurine methyltransferase|Thiopurine methyltransferase
C2599025|T201|COMP|53820-7|LNC|Cefozopran|Cefozopran
C2599026|T201|COMP|53821-5|LNC|Chloroamphetamine|Chloroamphetamine
C2599028|T201|COMP|53822-3|LNC|Flomoxef|Flomoxef
C2599029|T201|COMP|53823-1|LNC|Panipenem|Panipenem
C2599030|T201|COMP|53824-9|LNC|Paromomycin|Paromomycin
C2599031|T201|COMP|53825-6|LNC|HIV 1+Hepatitis C virus RNA|HIV 1+Hepatitis C virus RNA
C2599034|T201|COMP|53828-0|LNC|cycloSPORINE^trough|cycloSPORINE^trough
C2599035|T201|COMP|53829-8|LNC|Casein Ab.IgG|Casein Ab.IgG
C2599036|T201|COMP|53830-6|LNC|Granulocytes.CD55 deficient/100 cells|Granulocytes.CD55 deficient/100 cells
C2599038|T201|COMP|53831-4|LNC|Granulocytes.CD59 deficient/100 cells|Granulocytes.CD59 deficient/100 cells
C2599040|T201|COMP|53832-2|LNC|Erythrocytes.CD55 deficient/100 erythrocytes|Erythrocytes.CD55 deficient/100 erythrocytes
C2599042|T201|COMP|53833-0|LNC|Myoglobin|Myoglobin
C2599043|T201|COMP|53834-8|LNC|cycloSPORINE^peak|cycloSPORINE^peak
C2599044|T201|COMP|53835-5|LNC|1,5-Anhydroglucitol|1,5-Anhydroglucitol
C2599045|T201|COMP|53836-3|LNC|ABCD1 gene targeted mutation analysis|ABCD1 gene targeted mutation analysis
C2599047|T201|COMP|53837-1|LNC|ACVRL1 gene+ENG gene targeted mutation analysis|ACVRL1 gene+ENG gene targeted mutation analysis
C2599049|T201|COMP|53838-9|LNC|Arsenic.inorganic|Arsenic.inorganic
C2599050|T201|COMP|53839-7|LNC|Arsenic.organic|Arsenic.organic
C2599051|T201|COMP|53840-5|LNC|TGFB3 gene targeted mutation analysis|TGFB3 gene targeted mutation analysis
C2599053|T201|COMP|53841-3|LNC|ATRX gene targeted mutation analysis|ATRX gene targeted mutation analysis
C2599055|T201|COMP|53842-1|LNC|Basement membrane zone BP180 Ab.IgG|Basement membrane zone BP180 Ab.IgG
C2599057|T201|COMP|53843-9|LNC|Basement membrane zone BP230 Ab.IgG|Basement membrane zone BP230 Ab.IgG
C2599059|T201|COMP|53844-7|LNC|BRAF gene targeted mutation analysis|BRAF gene targeted mutation analysis
C2599061|T201|COMP|53845-4|LNC|BTD gene targeted mutation analysis|BTD gene targeted mutation analysis
C2599063|T201|COMP|53846-2|LNC|Buprenorphine|Buprenorphine
C2599064|T201|COMP|53847-0|LNC|CACT gene targeted mutation analysis|CACT gene targeted mutation analysis
C2599066|T201|COMP|53848-8|LNC|Mixed cellular casts|Mixed cellular casts
C2599067|T201|COMP|53849-6|LNC|HTC2 gene targeted mutation analysis|HTC2 gene targeted mutation analysis
C2599069|T201|COMP|53850-4|LNC|HTC2 gene mutations tested for|HTC2 gene mutations tested for
C2599071|T201|COMP|53851-2|LNC|COL10A1 gene targeted mutation analysis|COL10A1 gene targeted mutation analysis
C2599075|T201|COMP|53853-8|LNC|COL4A5 gene targeted mutation analysis|COL4A5 gene targeted mutation analysis
C2599077|T201|COMP|53854-6|LNC|CPS1 gene targeted mutation analysis|CPS1 gene targeted mutation analysis
C2599079|T201|COMP|53855-3|LNC|DNAI1+DNAH5 gene targeted mutation analysis|DNAI1+DNAH5 gene targeted mutation analysis
C2599081|T201|COMP|53856-1|LNC|DYSF gene targeted mutation analysis|DYSF gene targeted mutation analysis
C2599083|T201|COMP|53857-9|LNC|Hemoglobin F|Hemoglobin F
C2599084|T201|COMP|53858-7|LNC|EXT1 gene targeted mutation analysis|EXT1 gene targeted mutation analysis
C2599085|T201|COMP|53859-5|LNC|Fatty acids.very long chain.C22:0|Fatty acids.very long chain.C22:0
C2599086|T201|COMP|53860-3|LNC|Fatty acids.very long chain.C24:0|Fatty acids.very long chain.C24:0
C2599087|T201|COMP|53861-1|LNC|FKTN gene targeted mutation analysis|FKTN gene targeted mutation analysis
C2599089|T201|COMP|53862-9|LNC|FIG4 gene targeted mutation analysis|FIG4 gene targeted mutation analysis
C2599091|T201|COMP|53863-7|LNC|FLNA gene targeted mutation analysis|FLNA gene targeted mutation analysis
C2599093|T201|COMP|53864-5|LNC|GAA gene targeted mutation analysis|GAA gene targeted mutation analysis
C2599095|T201|COMP|53865-2|LNC|Galactomannan Ag|Galactomannan Ag
C2599096|T201|COMP|53866-0|LNC|GCH1 gene targeted mutation analysis|GCH1 gene targeted mutation analysis
C2599098|T201|COMP|53867-8|LNC|GYS2 gene targeted mutation analysis|GYS2 gene targeted mutation analysis
C2599100|T201|COMP|53868-6|LNC|Glucose tetrasaccharide/Creatinine|Glucose tetrasaccharide/Creatinine
C2599102|T201|COMP|53869-4|LNC|HPRT1 gene targeted mutation analysis|HPRT1 gene targeted mutation analysis
C2599104|T201|COMP|53870-2|LNC|HPS1 gene targeted mutation analysis|HPS1 gene targeted mutation analysis
C2599106|T201|COMP|53871-0|LNC|HRAS gene targeted mutation analysis|HRAS gene targeted mutation analysis
C2599107|T201|COMP|53872-8|LNC|Iodine|Iodine
C2599108|T201|COMP|53873-6|LNC|IRF6 gene targeted mutation analysis|IRF6 gene targeted mutation analysis
C2599110|T201|COMP|53874-4|LNC|Jamestown canyon virus RNA|Jamestown canyon virus RNA
C2599111|T201|COMP|53875-1|LNC|LMX1B gene targeted mutation analysis|LMX1B gene targeted mutation analysis
C2599113|T201|COMP|53876-9|LNC|LRRK2 gene targeted mutation analysis|LRRK2 gene targeted mutation analysis
C2599115|T201|COMP|53885-0|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C2599116|T201|COMP|53886-8|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C2599117|T201|COMP|53887-6|LNC|PCCA gene+PCCB gene targeted mutation analysis|PCCA gene+PCCB gene targeted mutation analysis
C2599119|T201|COMP|53888-4|LNC|PHEX gene targeted mutation analysis|PHEX gene targeted mutation analysis
C2599121|T201|COMP|53889-2|LNC|Platelet aggregation.arachidonate induced|Platelet aggregation.arachidonate induced
C2599122|T201|COMP|53890-0|LNC|PLOD1 gene targeted mutation analysis|PLOD1 gene targeted mutation analysis
C2599124|T201|COMP|53891-8|LNC|PNKD gene targeted mutation analysis|PNKD gene targeted mutation analysis
C2599131|T201|COMP|53892-6|LNC|Ribosomal P Ab.IgG|Ribosomal P Ab.IgG
C2599132|T201|COMP|53893-4|LNC|RNA polymerase III Ab|RNA polymerase III Ab
C2599134|T201|COMP|53894-2|LNC|TRAPPC2 gene targeted mutation analysis|TRAPPC2 gene targeted mutation analysis
C2599136|T201|COMP|53895-9|LNC|SH3BP2 gene targeted mutation analysis|SH3BP2 gene targeted mutation analysis
C2599138|T201|COMP|53896-7|LNC|SMC1A gene targeted mutation analysis|SMC1A gene targeted mutation analysis
C2599142|T201|COMP|53898-3|LNC|KIAA0196 gene targeted mutation analysis|KIAA0196 gene targeted mutation analysis
C2599146|T201|COMP|53900-7|LNC|C10orf2 gene targeted mutation analysis|C10orf2 gene targeted mutation analysis
C2599148|T201|COMP|53901-5|LNC|USH2A gene targeted mutation analysis|USH2A gene targeted mutation analysis
C2599150|T201|COMP|53902-3|LNC|Voriconazole|Voriconazole
C2599151|T201|COMP|53903-1|LNC|Collection method|Collection method
C2599156|T201|COMP|53908-0|LNC|Bacteria identified|Bacteria identified
C2599157|T201|COMP|53909-8|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C2599159|T201|COMP|53911-4|LNC|Bacteria identified|Bacteria identified
C2599165|T201|COMP|53917-1|LNC|Streptococcus pneumoniae DNA|Streptococcus pneumoniae DNA
C2599167|T201|COMP|53919-7|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C2599168|T201|COMP|53920-5|LNC|Thyroglobulin|Thyroglobulin
C2599169|T201|COMP|53921-3|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C2599170|T201|COMP|53922-1|LNC|Thyroglobulin|Thyroglobulin
C2599171|T201|COMP|53923-9|LNC|HIV 1 tropism|HIV 1 tropism
C2599172|T201|COMP|53924-7|LNC|Rheumatoid factor|Rheumatoid factor
C2599173|T201|COMP|53925-4|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C2599180|T201|COMP|53935-3|LNC|Clostridium tetani toxoid Ab.IgG|Clostridium tetani toxoid Ab.IgG
C2599181|T201|COMP|53936-1|LNC|Cells.CD3-CD56+|Cells.CD3-CD56+
C2599182|T201|COMP|53937-9|LNC|HLA-B w4+w6|HLA-B w4+w6
C2599184|T201|COMP|53938-7|LNC|HLA-DQB1|HLA-DQB1
C2599186|T201|COMP|53939-5|LNC|CD4 stimulated ATP immune response|CD4 stimulated ATP immune response
C2599188|T201|COMP|53940-3|LNC|CD4 stimulated ATP immune response|CD4 stimulated ATP immune response
C2599189|T201|COMP|53941-1|LNC|Vibrio cholerae toxin Ag|Vibrio cholerae toxin Ag
C2599191|T201|COMP|53942-9|LNC|Vibrio cholerae toxin ctx gene|Vibrio cholerae toxin ctx gene
C2599193|T201|COMP|53943-7|LNC|Bacterial cytolethal distending toxin cdt gene|Bacterial cytolethal distending toxin cdt gene
C2599195|T201|COMP|53944-5|LNC|Escherichia coli enteroinvasive|Escherichia coli enteroinvasive
C2599196|T201|COMP|53945-2|LNC|Escherichia coli adherence pattern|Escherichia coli adherence pattern
C2599198|T201|COMP|53946-0|LNC|Escherichia coli shiga-like toxin identified|Escherichia coli shiga-like toxin identified
C2599202|T201|COMP|53948-6|LNC|Donated egg|Donated egg
C2599204|T201|COMP|53949-4|LNC|HPA 1a-1a+HPA 3b-3b|HPA 1a-1a+HPA 3b-3b
C2599206|T201|COMP|53950-2|LNC|HPA 1a-1a+Glycoprotein IIb-IIIa|HPA 1a-1a+Glycoprotein IIb-IIIa
C2599208|T201|COMP|53951-0|LNC|HPA 1b-1b+HPA 3a-3a|HPA 1b-1b+HPA 3a-3a
C2599210|T201|COMP|53952-8|LNC|HPA 1b-1b+Glycoprotein IIb-IIIa|HPA 1b-1b+Glycoprotein IIb-IIIa
C2599212|T201|COMP|53953-6|LNC|HPA 5a-5a+Glycoprotein Ia-IIa|HPA 5a-5a+Glycoprotein Ia-IIa
C2599214|T201|COMP|53954-4|LNC|HPA 5a-5b+Glycoprotein Ia-IIa|HPA 5a-5b+Glycoprotein Ia-IIa
C2599216|T201|COMP|53955-1|LNC|Escherichia coli O157 identified|Escherichia coli O157 identified
C2599218|T201|COMP|53956-9|LNC|Salmonella typhi|Salmonella typhi
C2599219|T201|COMP|53957-7|LNC|Choriogonadotropin.tumor marker|Choriogonadotropin.tumor marker
C2599220|T201|COMP|53972-6|LNC|Burr cells|Burr cells
C2599221|T201|COMP|53973-4|LNC|Erythrocytes.ghost cells|Erythrocytes.ghost cells
C2599222|T201|COMP|53974-2|LNC|Erythrocyte morphology|Erythrocyte morphology
C2599224|T201|COMP|53975-9|LNC|Drug crystals|Drug crystals
C2599226|T201|COMP|53976-7|LNC|Pseudocasts|Pseudocasts
C2599227|T201|COMP|53977-5|LNC|Dimagnesium phosphate crystals|Dimagnesium phosphate crystals
C2599229|T201|COMP|53978-3|LNC|Epithelial cells.non-squamous|Epithelial cells.non-squamous
C2599230|T201|COMP|53979-1|LNC|Actin Ab|Actin Ab
C2599231|T201|COMP|53980-9|LNC|Actin Ab|Actin Ab
C2599232|T201|COMP|53981-7|LNC|Centromere protein B Ab|Centromere protein B Ab
C2599234|T201|COMP|53982-5|LNC|Centromere protein B Ab|Centromere protein B Ab
C2599235|T201|COMP|53983-3|LNC|Nuclear Ab pattern.homogeneous|Nuclear Ab pattern.homogeneous
C2599236|T201|COMP|53984-1|LNC|Nuclear Ab pattern.fine speckled|Nuclear Ab pattern.fine speckled
C2599237|T201|COMP|53985-8|LNC|Nuclear Ab pattern.coarse speckled|Nuclear Ab pattern.coarse speckled
C2599239|T201|COMP|53986-6|LNC|Nuclear Ab pattern.coarse speckled|Nuclear Ab pattern.coarse speckled
C2599240|T201|COMP|53987-4|LNC|Nuclear Ab pattern.atypic speckled|Nuclear Ab pattern.atypic speckled
C2599242|T201|COMP|53988-2|LNC|Nuclear Ab pattern.atypic speckled|Nuclear Ab pattern.atypic speckled
C2599243|T201|COMP|53989-0|LNC|Nuclear Ab pattern.chromosomal|Nuclear Ab pattern.chromosomal
C2599245|T201|COMP|53990-8|LNC|Nuclear Ab pattern.chromosomal|Nuclear Ab pattern.chromosomal
C2599246|T201|COMP|53991-6|LNC|Nuclear Ab pattern.nucleolar|Nuclear Ab pattern.nucleolar
C2599247|T201|COMP|53992-4|LNC|Nuclear Ab pattern.nucleolar|Nuclear Ab pattern.nucleolar
C2599248|T201|COMP|53993-2|LNC|Nuclear Ab pattern.centrosomal|Nuclear Ab pattern.centrosomal
C2599250|T201|COMP|53994-0|LNC|Nuclear Ab pattern.centrosomal|Nuclear Ab pattern.centrosomal
C2599251|T201|COMP|53995-7|LNC|Nuclear Ab pattern.nuclear matrix|Nuclear Ab pattern.nuclear matrix
C2599253|T201|COMP|53996-5|LNC|Nuclear Ab pattern.nuclear matrix|Nuclear Ab pattern.nuclear matrix
C2599254|T201|COMP|53997-3|LNC|Nuclear Ab pattern.nuclear dots|Nuclear Ab pattern.nuclear dots
C2599256|T201|COMP|53998-1|LNC|Nuclear Ab pattern.nuclear dots|Nuclear Ab pattern.nuclear dots
C2599257|T201|COMP|53999-9|LNC|Nuclear Ab pattern.multiple nuclear dots|Nuclear Ab pattern.multiple nuclear dots
C2599259|T201|COMP|54000-5|LNC|Nuclear Ab pattern.multiple nuclear dots|Nuclear Ab pattern.multiple nuclear dots
C2599260|T201|COMP|54001-3|LNC|Centromere protein F Ab|Centromere protein F Ab
C2599262|T201|COMP|54002-1|LNC|Centromere protein F Ab|Centromere protein F Ab
C2599263|T201|COMP|54003-9|LNC|Human upstream binding factor Ab|Human upstream binding factor Ab
C2599265|T201|COMP|54004-7|LNC|Human upstream binding factor Ab|Human upstream binding factor Ab
C2599266|T201|COMP|54005-4|LNC|Nuclear Ab pattern.nuclear membrane pores|Nuclear Ab pattern.nuclear membrane pores
C2599268|T201|COMP|54006-2|LNC|Nuclear Ab pattern.nuclear membrane pores|Nuclear Ab pattern.nuclear membrane pores
C2599269|T201|COMP|54007-0|LNC|Golgi apparatus Ab|Golgi apparatus Ab
C2599271|T201|COMP|54008-8|LNC|Golgi apparatus Ab|Golgi apparatus Ab
C2599272|T201|COMP|54009-6|LNC|Lysosome Ab|Lysosome Ab
C2599274|T201|COMP|54010-4|LNC|Lysosome Ab|Lysosome Ab
C2599275|T201|COMP|54011-2|LNC|Vimentin Ab|Vimentin Ab
C2599276|T201|COMP|54012-0|LNC|Vimentin Ab|Vimentin Ab
C2599277|T201|COMP|54013-8|LNC|Vinculin Ab|Vinculin Ab
C2599279|T201|COMP|54014-6|LNC|Vinculin Ab|Vinculin Ab
C2599280|T201|COMP|54015-3|LNC|Azurocidin Ab|Azurocidin Ab
C2599282|T201|COMP|54016-1|LNC|Cathepsin G Ab|Cathepsin G Ab
C2599283|T201|COMP|54017-9|LNC|Elastase Ab|Elastase Ab
C2599284|T201|COMP|54018-7|LNC|Lactoferrin Ab|Lactoferrin Ab
C2599285|T201|COMP|54019-5|LNC|Lysozyme Ab|Lysozyme Ab
C2599286|T201|COMP|54020-3|LNC|Actin.filamentous Ab|Actin.filamentous Ab
C2599288|T201|COMP|54021-1|LNC|Actin.filamentous Ab|Actin.filamentous Ab
C2599289|T201|COMP|54022-9|LNC|Mutated citrullinated vimentin Ab|Mutated citrullinated vimentin Ab
C2599291|T201|COMP|54023-7|LNC|U1 small nuclear ribonucleoprotein C Ab|U1 small nuclear ribonucleoprotein C Ab
C2599293|T201|COMP|54024-5|LNC|sp100 Ab|sp100 Ab
C2599295|T201|COMP|54025-2|LNC|Nuclear pore protein gp210 Ab|Nuclear pore protein gp210 Ab
C2599297|T201|COMP|54026-0|LNC|Soluble liver Ab|Soluble liver Ab
C2599299|T201|COMP|54027-8|LNC|Lamin Ab|Lamin Ab
C2599301|T201|COMP|54028-6|LNC|Lamin Ab|Lamin Ab
C2599302|T201|COMP|54029-4|LNC|Soluble liver Ab|Soluble liver Ab
C2599303|T201|COMP|54030-2|LNC|Smith extractable nuclear B Ab|Smith extractable nuclear B Ab
C2599305|T201|COMP|54031-0|LNC|Smith extractable nuclear D Ab|Smith extractable nuclear D Ab
C2599307|T201|COMP|54032-8|LNC|U1 small nuclear ribonucleoprotein A Ab|U1 small nuclear ribonucleoprotein A Ab
C2599309|T201|COMP|54033-6|LNC|Rickettsia spotted fever group Ag|Rickettsia spotted fever group Ag
C2599310|T201|COMP|54034-4|LNC|Anaplasma phagocytophilum Ag|Anaplasma phagocytophilum Ag
C2599312|T201|COMP|54035-1|LNC|Ehrlichia chaffeensis Ag|Ehrlichia chaffeensis Ag
C2599313|T201|COMP|54036-9|LNC|Western equine encephalitis virus RNA|Western equine encephalitis virus RNA
C2599314|T201|COMP|54037-7|LNC|HEDIS 2009 panel|HEDIS 2009 panel
C2599338|T201|COMP|54049-2|LNC|HEDIS 2009-2013 Codes to identify lead (LSC-A)|HEDIS 2009-2013 Codes to identify lead (LSC-A)
C2599374|T201|COMP|54067-4|LNC|Clostridioides difficile toxin genes|Clostridioides difficile toxin genes
C2599376|T201|COMP|54068-2|LNC|Hemoglobin O-Arab/Hemoglobin.total|Hemoglobin O-Arab/Hemoglobin.total
C2599377|T201|COMP|54069-0|LNC|Hemoglobin Barts/Hemoglobin.total|Hemoglobin Barts/Hemoglobin.total
C2599378|T201|COMP|54070-8|LNC|Hemoglobin D/Hemoglobin.total|Hemoglobin D/Hemoglobin.total
C2599379|T201|COMP|54071-6|LNC|Hemoglobin E/Hemoglobin.total|Hemoglobin E/Hemoglobin.total
C2599380|T201|COMP|54072-4|LNC|Hemoglobin A/Hemoglobin.total|Hemoglobin A/Hemoglobin.total
C2599381|T201|COMP|54073-2|LNC|Hemoglobin C/Hemoglobin.total|Hemoglobin C/Hemoglobin.total
C2599382|T201|COMP|54074-0|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C2599383|T201|COMP|54075-7|LNC|Endocrine newborn screening panel (SI units)|Endocrine newborn screening panel (SI units)
C2599385|T201|COMP|54076-5|LNC|Endocrine newborn screening panel|Endocrine newborn screening panel
C2599386|T201|COMP|54077-3|LNC|Thyroid newborn screening panel (SI units)|Thyroid newborn screening panel (SI units)
C2599388|T201|COMP|54078-1|LNC|Cystic fibrosis newborn screening panel|Cystic fibrosis newborn screening panel
C2599390|T201|COMP|54079-9|LNC|Galactosemia newborn screening panel|Galactosemia newborn screening panel
C2599392|T201|COMP|54080-7|LNC|Galactosemia newborn screening panel (SI units)|Galactosemia newborn screening panel (SI units)
C2599393|T201|COMP|54081-5|LNC|Hemoglobinopathies newborn screening panel|Hemoglobinopathies newborn screening panel
C2599395|T201|COMP|54082-3|LNC|Infectious diseases newborn screening panel|Infectious diseases newborn screening panel
C2599397|T201|COMP|54083-1|LNC|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C2599398|T201|COMP|54084-9|LNC|Galactose|Galactose
C2599399|T201|COMP|54085-6|LNC|Galactose|Galactose
C2599400|T201|COMP|54086-4|LNC|HIV 1+2 Ab.IgG|HIV 1+2 Ab.IgG
C2599401|T201|COMP|54087-2|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C2599402|T201|COMP|54088-0|LNC|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C2599403|T201|COMP|54089-8|LNC|Newborn screening panel|Newborn screening panel
C2599404|T201|COMP|54090-6|LNC|Thyroid newborn screening panel|Thyroid newborn screening panel
C2599405|T201|COMP|54091-4|LNC|Rubella virus RNA|Rubella virus RNA
C2599407|T201|COMP|54092-2|LNC|Citrulline/Arginine|Citrulline/Arginine
C2599409|T201|COMP|54093-0|LNC|Pesticides|Pesticides
C2599412|T201|COMP|54095-5|LNC|Chemotherapy effectiveness panel|Chemotherapy effectiveness panel
C2599414|T201|COMP|54096-3|LNC|Identity testing|Identity testing
C2599416|T201|COMP|54097-1|LNC|Organophosphonate nerve agent metabolite panel|Organophosphonate nerve agent metabolite panel
C2599418|T201|COMP|54098-9|LNC|Isopropyl methylphosphonate|Isopropyl methylphosphonate
C2599420|T201|COMP|54099-7|LNC|1,2,2-Trimethylpropyl methylphosphonate|1,2,2-Trimethylpropyl methylphosphonate
C2599422|T201|COMP|54100-3|LNC|Monocyclohexyl methylphosphonate|Monocyclohexyl methylphosphonate
C2599424|T201|COMP|54101-1|LNC|2-Methylpropyl methylphosphonate|2-Methylpropyl methylphosphonate
C2599426|T201|COMP|54102-9|LNC|Monoethyl methylphosphonate|Monoethyl methylphosphonate
C2599428|T201|COMP|54103-7|LNC|Hemoglobin pattern|Hemoglobin pattern
C2599429|T201|COMP|54104-5|LNC|Hemoglobin pattern|Hemoglobin pattern
C2599430|T201|COMP|54105-2|LNC|Hemoglobin pattern|Hemoglobin pattern
C2603365|T201|COMP|16629-8|LNC|Coagulation surface induced|Coagulation surface induced
C2603368|T201|COMP|16321-2|LNC|Acyl carnitine|Acyl carnitine
C2603371|T201|COMP|40573-8|LNC|Lymphocytes.variant|Lymphocytes.variant
C2603373|T201|COMP|35255-9|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C2603374|T201|COMP|35257-5|LNC|Natriuretic peptide.B|Natriuretic peptide.B
C2603375|T201|COMP|35234-4|LNC|Urea nitrogen|Urea nitrogen
C2603376|T201|COMP|604-9|LNC|Bacteria identified|Bacteria identified
C2603377|T201|COMP|17881-4|LNC|Bacteria identified^^^5|Bacteria identified^^^5
C2603378|T201|COMP|17880-6|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C2603379|T201|COMP|17879-8|LNC|Bacteria identified^^^3|Bacteria identified^^^3
C2603387|T201|COMP|35197-3|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C2603388|T201|COMP|35198-1|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C2603389|T201|COMP|35199-9|LNC|Cholesterol.in VLDL|Cholesterol.in VLDL
C2603390|T201|COMP|35200-5|LNC|Cholesterol|Cholesterol
C2603391|T201|COMP|35201-3|LNC|Cobalamins|Cobalamins
C2603393|T201|COMP|35206-2|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C2603394|T201|COMP|35205-4|LNC|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C2603395|T201|COMP|35355-7|LNC|PABPN1 gene targeted mutation analysis|PABPN1 gene targeted mutation analysis
C2603399|T201|COMP|21694-5|LNC|HFE gene targeted mutation analysis|HFE gene targeted mutation analysis
C2603400|T201|COMP|35244-3|LNC|Digoxin|Digoxin
C2607826|T201|COMP|14337-0|LNC|Phenytoin.total/Phenytoin.free|Phenytoin.total/Phenytoin.free
C2607827|T201|COMP|41107-4|LNC|FMR1 gene targeted mutation analysis|FMR1 gene targeted mutation analysis
C2607828|T201|COMP|13599-6|LNC|Promonocytes/100 leukocytes|Promonocytes/100 leukocytes
C2607829|T201|COMP|35209-6|LNC|Ferritin|Ferritin
C2607830|T201|COMP|42568-6|LNC|Fibrinogen|Fibrinogen
C2607831|T201|COMP|35210-4|LNC|Folate|Folate
C2607833|T201|COMP|41104-1|LNC|GBA gene targeted mutation analysis|GBA gene targeted mutation analysis
C2607834|T201|COMP|41101-7|LNC|GJB2 gene targeted mutation analysis|GJB2 gene targeted mutation analysis
C2607835|T201|COMP|41099-3|LNC|GLA gene targeted mutation analysis|GLA gene targeted mutation analysis
C2607836|T201|COMP|35211-2|LNC|Glucose|Glucose
C2607837|T201|COMP|35212-0|LNC|Glucose|Glucose
C2607838|T201|COMP|35184-1|LNC|Glucose^post CFst|Glucose^post CFst
C2607839|T201|COMP|40294-1|LNC|Insulin^pre or post dose glucose|Insulin^pre or post dose glucose
C2607840|T201|COMP|17637-0|LNC|Streptococcus pneumoniae 6b Ab^2nd specimen|Streptococcus pneumoniae 6b Ab^2nd specimen
C2607841|T201|COMP|22554-0|LNC|Streptococcus pneumoniae 7f Ab^2nd specimen|Streptococcus pneumoniae 7f Ab^2nd specimen
C2607842|T201|COMP|17620-6|LNC|Streptococcus pneumoniae 18c Ab^1st specimen|Streptococcus pneumoniae 18c Ab^1st specimen
C2607843|T201|COMP|17621-4|LNC|Streptococcus pneumoniae 18c Ab^2nd specimen|Streptococcus pneumoniae 18c Ab^2nd specimen
C2607844|T201|COMP|22559-9|LNC|Streptococcus pneumoniae 9n Ab^1st specimen|Streptococcus pneumoniae 9n Ab^1st specimen
C2607845|T201|COMP|10852-2|LNC|Fungus identified|Fungus identified
C2607847|T201|COMP|35238-5|LNC|Theophylline|Theophylline
C2607848|T201|COMP|35239-3|LNC|Tobramycin^trough|Tobramycin^trough
C2607849|T201|COMP|35241-9|LNC|Urea nitrogen|Urea nitrogen
C2607853|T201|COMP|41088-6|LNC|MERRF gene targeted mutation analysis|MERRF gene targeted mutation analysis
C2607854|T201|COMP|35252-6|LNC|Magnesium|Magnesium
C2607855|T201|COMP|35249-2|LNC|Magnesium|Magnesium
C2607856|T201|COMP|35250-0|LNC|Magnesium|Magnesium
C2607936|T201|COMP|7357-7|LNC|Poa pratensis Ab.IgE|Poa pratensis Ab.IgE
C2607937|T201|COMP|7540-8|LNC|Avena sativa cultivated Ab.IgE|Avena sativa cultivated Ab.IgE
C2607937|T201|COMP|6191-1|LNC|Avena sativa cultivated Ab.IgE|Avena sativa cultivated Ab.IgE
C2607938|T201|COMP|5439-5|LNC|CD16+CD57+|CD16+CD57+
C2607952|T201|COMP|10962-9|LNC|Artemisia tridentata Ab.IgE|Artemisia tridentata Ab.IgE
C2607952|T201|COMP|7684-4|LNC|Artemisia tridentata Ab.IgE|Artemisia tridentata Ab.IgE
C2607995|T201|COMP|14845-2|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C2706069|T201|COMP|54146-6|LNC|Mycobacterium tuberculosis Ab.IgG|Mycobacterium tuberculosis Ab.IgG
C2706070|T201|COMP|54147-4|LNC|Autoantibodies|Autoantibodies
C2706071|T201|COMP|54148-2|LNC|Autoantibodies|Autoantibodies
C2706072|T201|COMP|54149-0|LNC|Nuclear Ab pattern.homogeneous|Nuclear Ab pattern.homogeneous
C2706073|T201|COMP|54150-8|LNC|Centriole Ab|Centriole Ab
C2706074|T201|COMP|54151-6|LNC|Centriole Ab|Centriole Ab
C2706075|T201|COMP|54152-4|LNC|Nuclear mitotic apparatus Ab|Nuclear mitotic apparatus Ab
C2706076|T201|COMP|54153-2|LNC|Nuclear mitotic apparatus Ab|Nuclear mitotic apparatus Ab
C2706077|T201|COMP|54154-0|LNC|Midbody Ab|Midbody Ab
C2706644|T201|COMP|54443-7|LNC|Echovirus 2 Ab|Echovirus 2 Ab
C2706646|T201|COMP|54444-5|LNC|Echovirus 8 Ab|Echovirus 8 Ab
C2706648|T201|COMP|54445-2|LNC|Fatty acids.very long chain.C22:1n9|Fatty acids.very long chain.C22:1n9
C2706650|T201|COMP|54446-0|LNC|Fatty acids.very long chain.C26:1|Fatty acids.very long chain.C26:1
C2706651|T201|COMP|54447-8|LNC|FLT3 gene targeted mutation analysis|FLT3 gene targeted mutation analysis
C2706652|T201|COMP|54448-6|LNC|NPM1 gene targeted mutation analysis|NPM1 gene targeted mutation analysis
C2706654|T201|COMP|54449-4|LNC|SMN2 gene targeted mutation analysis|SMN2 gene targeted mutation analysis
C2706656|T201|COMP|54450-2|LNC|CYP2C9 & VKORC1 panel|CYP2C9 & VKORC1 panel
C2706659|T201|COMP|54166-4|LNC|Cefoperazone+Sulbactam|Cefoperazone+Sulbactam
C2706660|T201|COMP|54167-2|LNC|Cefoperazone+Sulbactam|Cefoperazone+Sulbactam
C2706661|T201|COMP|54168-0|LNC|Cefoperazone+Sulbactam|Cefoperazone+Sulbactam
C2706662|T201|COMP|54169-8|LNC|Thiamphenicol|Thiamphenicol
C2706663|T201|COMP|54170-6|LNC|Imipenem+EDTA|Imipenem+EDTA
C2706664|T201|COMP|54171-4|LNC|Imipenem+EDTA|Imipenem+EDTA
C2706665|T201|COMP|54172-2|LNC|Imipenem+EDTA|Imipenem+EDTA
C2706666|T201|COMP|54173-0|LNC|Arbekacin|Arbekacin
C2706682|T201|COMP|55289-3|LNC|Sulopenem|Sulopenem
C2706683|T201|COMP|55290-1|LNC|Sulopenem|Sulopenem
C2706684|T201|COMP|55291-9|LNC|Sulopenem|Sulopenem
C2706685|T201|COMP|55292-7|LNC|Linopristin+Flopristin|Linopristin+Flopristin
C2706687|T201|COMP|55529-2|LNC|Clopenthixol|Clopenthixol
C2706688|T201|COMP|55530-0|LNC|Cocaethylene|Cocaethylene
C2706689|T201|COMP|55531-8|LNC|Cyclobenzaprine|Cyclobenzaprine
C2706690|T201|COMP|55532-6|LNC|Diethylpropion|Diethylpropion
C2706691|T201|COMP|55533-4|LNC|dilTIAZem|dilTIAZem
C2706692|T201|COMP|55534-2|LNC|Doxylamine|Doxylamine
C2706693|T201|COMP|55535-9|LNC|ePHEDrine|ePHEDrine
C2706694|T201|COMP|55536-7|LNC|Fenoprofen|Fenoprofen
C2706695|T201|COMP|55537-5|LNC|fentaNYL|fentaNYL
C2706696|T201|COMP|55538-3|LNC|Flupenthixol|Flupenthixol
C2706697|T201|COMP|55539-1|LNC|Flurbiprofen|Flurbiprofen
C2706698|T201|COMP|54362-9|LNC|Bilirubin|Bilirubin
C2706699|T201|COMP|54363-7|LNC|Bilirubin|Bilirubin
C2706700|T201|COMP|54364-5|LNC|Calcium|Calcium
C2706701|T201|COMP|54365-2|LNC|Calcium|Calcium
C2706702|T201|COMP|54366-0|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C2706703|T201|COMP|54367-8|LNC|Calcium.ionized|Calcium.ionized
C2706704|T201|COMP|54368-6|LNC|Catalase|Catalase
C2706705|T201|COMP|54369-4|LNC|Chloride^post dialysis|Chloride^post dialysis
C2706706|T201|COMP|54370-2|LNC|Chloride|Chloride
C2706707|T201|COMP|54371-0|LNC|Cholesterol|Cholesterol
C2706708|T201|COMP|54372-8|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C2706709|T201|COMP|54373-6|LNC|Cholesterol.non-esterified|Cholesterol.non-esterified
C2706710|T201|COMP|54374-4|LNC|Creatinine/body weight|Creatinine/body weight
C2706711|T201|COMP|54375-1|LNC|Creatinine|Creatinine
C2706712|T201|COMP|54376-9|LNC|Cobalamins|Cobalamins
C2706713|T201|COMP|54377-7|LNC|Cobalamins|Cobalamins
C2706714|T201|COMP|54378-5|LNC|Cobalamins|Cobalamins
C2706715|T201|COMP|54379-3|LNC|Cystatin C/Creatinine|Cystatin C/Creatinine
C2706720|T201|COMP|54142-5|LNC|Candida sp DNA|Candida sp DNA
C2706721|T201|COMP|54143-3|LNC|Gardnerella vaginalis DNA|Gardnerella vaginalis DNA
C2706722|T201|COMP|54144-1|LNC|Trichomonas vaginalis DNA|Trichomonas vaginalis DNA
C2706723|T201|COMP|54145-8|LNC|Bacterial vaginosis & vaginitis DNA panel|Bacterial vaginosis & vaginitis DNA panel
C2706724|T201|COMP|54155-7|LNC|Midbody Ab|Midbody Ab
C2706725|T201|COMP|54156-5|LNC|RNA polymerase I Ab|RNA polymerase I Ab
C2706726|T201|COMP|54157-3|LNC|RNA polymerase I Ab|RNA polymerase I Ab
C2706727|T201|COMP|54158-1|LNC|Pancytokeratin Ab|Pancytokeratin Ab
C2706728|T201|COMP|54159-9|LNC|Pancytokeratin Ab|Pancytokeratin Ab
C2706729|T201|COMP|54160-7|LNC|Ki Ab|Ki Ab
C2706730|T201|COMP|54161-5|LNC|Cytoplasmic Ab pattern.PL-7+PL-12|Cytoplasmic Ab pattern.PL-7+PL-12
C2706731|T201|COMP|54162-3|LNC|Cytoplasmic Ab pattern.PL-7+PL-12|Cytoplasmic Ab pattern.PL-7+PL-12
C2706732|T201|COMP|54163-1|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C2706733|T201|COMP|54164-9|LNC|Cytomegalovirus immediate-early Ag|Cytomegalovirus immediate-early Ag
C2706734|T201|COMP|54165-6|LNC|Tumor necrosis factor binding protein|Tumor necrosis factor binding protein
C2706735|T201|COMP|54174-8|LNC|Cefmenoxime|Cefmenoxime
C2706736|T201|COMP|54175-5|LNC|Caspofungin|Caspofungin
C2706737|T201|COMP|54176-3|LNC|Caspofungin|Caspofungin
C2706738|T201|COMP|54177-1|LNC|Clotrimazole|Clotrimazole
C2706739|T201|COMP|54178-9|LNC|Econazole|Econazole
C2706740|T201|COMP|54179-7|LNC|Itraconazole|Itraconazole
C2706741|T201|COMP|54180-5|LNC|Miconazole|Miconazole
C2706742|T201|COMP|54181-3|LNC|Nitroxoline|Nitroxoline
C2706743|T201|COMP|54182-1|LNC|Para aminosalicylate|Para aminosalicylate
C2706744|T201|COMP|54183-9|LNC|Rifabutin|Rifabutin
C2706745|T201|COMP|54184-7|LNC|Thiacetazone|Thiacetazone
C2706746|T201|COMP|54185-4|LNC|Caspofungin|Caspofungin
C2706747|T201|COMP|54186-2|LNC|Posaconazole|Posaconazole
C2706748|T201|COMP|54187-0|LNC|Posaconazole|Posaconazole
C2706749|T201|COMP|54188-8|LNC|Posaconazole|Posaconazole
C2706750|T201|COMP|54189-6|LNC|Posaconazole|Posaconazole
C2706751|T201|COMP|54190-4|LNC|Temocillin|Temocillin
C2706752|T201|COMP|54191-2|LNC|Cefotaxime+Sulbactam|Cefotaxime+Sulbactam
C2706753|T201|COMP|54192-0|LNC|Cefotaxime+Sulbactam|Cefotaxime+Sulbactam
C2706754|T201|COMP|54193-8|LNC|Cefotaxime+Sulbactam|Cefotaxime+Sulbactam
C2706755|T201|COMP|54194-6|LNC|Mezlocillin+Sulbactam|Mezlocillin+Sulbactam
C2706756|T201|COMP|54195-3|LNC|Mezlocillin+Sulbactam|Mezlocillin+Sulbactam
C2706757|T201|COMP|54196-1|LNC|Mezlocillin+Sulbactam|Mezlocillin+Sulbactam
C2706758|T201|COMP|54197-9|LNC|Piperacillin+Sulbactam|Piperacillin+Sulbactam
C2706759|T201|COMP|54198-7|LNC|Piperacillin+Sulbactam|Piperacillin+Sulbactam
C2706760|T201|COMP|54199-5|LNC|Piperacillin+Sulbactam|Piperacillin+Sulbactam
C2706761|T201|COMP|54200-1|LNC|Griseofulvin|Griseofulvin
C2706762|T201|COMP|54201-9|LNC|Griseofulvin|Griseofulvin
C2706763|T201|COMP|54202-7|LNC|Griseofulvin|Griseofulvin
C2706764|T201|COMP|54203-5|LNC|Cefmenoxime|Cefmenoxime
C2706765|T201|COMP|54204-3|LNC|Thiacetazone|Thiacetazone
C2706766|T201|COMP|54205-0|LNC|Legionella pneumophila 7+8+9+10+11+12+13+14 Ab|Legionella pneumophila 7+8+9+10+11+12+13+14 Ab
C2706767|T201|COMP|54206-8|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C2706770|T201|COMP|54209-2|LNC|Hemoglobin C-Harlem/Hemoglobin.total|Hemoglobin C-Harlem/Hemoglobin.total
C2706772|T201|COMP|54210-0|LNC|Hepatitis B virus basal core promoter mutation|Hepatitis B virus basal core promoter mutation
C2706773|T201|COMP|54211-8|LNC|Cortisol^24H post dose dexamethasone|Cortisol^24H post dose dexamethasone
C2706774|T201|COMP|54212-6|LNC|Cortisol^3D post dose dexamethasone|Cortisol^3D post dose dexamethasone
C2706775|T201|COMP|54213-4|LNC|Cortisol^4D post dose corticotropin|Cortisol^4D post dose corticotropin
C2706776|T201|COMP|54214-2|LNC|Cortisol^5D post dose dexamethasone|Cortisol^5D post dose dexamethasone
C2706777|T201|COMP|54215-9|LNC|Cortisol^5H post dose corticotropin|Cortisol^5H post dose corticotropin
C2706780|T201|COMP|54218-3|LNC|Cells.CD3+CD4+/Cells.CD3+CD8+|Cells.CD3+CD4+/Cells.CD3+CD8+
C2706783|T201|COMP|54220-9|LNC|Immune response markers|Immune response markers
C2706784|T201|COMP|54221-7|LNC|Lymphoma markers|Lymphoma markers
C2706785|T201|COMP|54222-5|LNC|Lymphoma - acute screen markers|Lymphoma - acute screen markers
C2706786|T201|COMP|54223-3|LNC|Lymphoma - CLL screen markers|Lymphoma - CLL screen markers
C2706787|T201|COMP|54224-1|LNC|Lymphoma - T-cell markers|Lymphoma - T-cell markers
C2706788|T201|COMP|54225-8|LNC|Immune response panel|Immune response panel
C2706789|T201|COMP|54226-6|LNC|Lymphoma panel|Lymphoma panel
C2706790|T201|COMP|54227-4|LNC|Lymphoma - acute screen panel|Lymphoma - acute screen panel
C2706791|T201|COMP|54228-2|LNC|Lymphoma - CLL screen panel|Lymphoma - CLL screen panel
C2706792|T201|COMP|54229-0|LNC|Lymphoma - T-cell screen panel|Lymphoma - T-cell screen panel
C2706794|T201|COMP|54231-6|LNC|Semen analysis fertility panel|Semen analysis fertility panel
C2706795|T201|COMP|54232-4|LNC|Metabolic panel.large animal|Metabolic panel.large animal
C2706796|T201|COMP|54233-2|LNC|Metabolic panel.small animal|Metabolic panel.small animal
C2706798|T201|COMP|54235-7|LNC|Cortisol challenge panel|Cortisol challenge panel
C2706799|T201|COMP|54236-5|LNC|Cortisol^9 AM 2nd day specimen|Cortisol^9 AM 2nd day specimen
C2706800|T201|COMP|54237-3|LNC|Corticotropin^9 AM 2nd day specimen|Corticotropin^9 AM 2nd day specimen
C2706801|T201|COMP|54238-1|LNC|LDL.oxidized|LDL.oxidized
C2706802|T201|COMP|54239-9|LNC|Cytopathic effect|Cytopathic effect
C2706803|T201|COMP|54240-7|LNC|Influenza virus Ag|Influenza virus Ag
C2706804|T201|COMP|54241-5|LNC|Influenza virus B Ag|Influenza virus B Ag
C2706805|T201|COMP|54242-3|LNC|Influenza virus identified|Influenza virus identified
C2706806|T201|COMP|54243-1|LNC|Influenza virus RNA|Influenza virus RNA
C2706807|T201|COMP|54244-9|LNC|Influenza virus identified|Influenza virus identified
C2706808|T201|COMP|54245-6|LNC|Respiratory virus Ag|Respiratory virus Ag
C2706809|T201|COMP|54246-4|LNC|Protein & Glucose panel|Protein & Glucose panel
C2706810|T201|COMP|54247-2|LNC|Drug screen comment|Drug screen comment
C2706811|T201|COMP|54248-0|LNC|Glucose^10M pre dose glucagon|Glucose^10M pre dose glucagon
C2706812|T201|COMP|54249-8|LNC|Glucose^15M post dose glucagon|Glucose^15M post dose glucagon
C2706813|T201|COMP|54250-6|LNC|Glucose^15M pre dose glucagon|Glucose^15M pre dose glucagon
C2706814|T201|COMP|54251-4|LNC|Glucose^20M post dose glucagon|Glucose^20M post dose glucagon
C2706815|T201|COMP|54252-2|LNC|Glucose^2M post dose glucagon|Glucose^2M post dose glucagon
C2706816|T201|COMP|54253-0|LNC|Glucose^4M post dose glucagon|Glucose^4M post dose glucagon
C2706817|T201|COMP|54254-8|LNC|Glucose^5M pre dose glucagon|Glucose^5M pre dose glucagon
C2706818|T201|COMP|54255-5|LNC|Glucose^6M post dose glucagon|Glucose^6M post dose glucagon
C2706819|T201|COMP|54256-3|LNC|Glucose^8M post dose glucagon|Glucose^8M post dose glucagon
C2706820|T201|COMP|54257-1|LNC|Glucose^pre dose insulin IV|Glucose^pre dose insulin IV
C2706821|T201|COMP|54258-9|LNC|Glucose^2H post dose insulin IV|Glucose^2H post dose insulin IV
C2706822|T201|COMP|54259-7|LNC|Glucose^2.5H post dose insulin IV|Glucose^2.5H post dose insulin IV
C2706823|T201|COMP|54260-5|LNC|Glucose^15M post dose insulin IV|Glucose^15M post dose insulin IV
C2706824|T201|COMP|54261-3|LNC|Glucose^15M pre dose insulin IV|Glucose^15M pre dose insulin IV
C2706825|T201|COMP|54262-1|LNC|Glucose^3H pre dose insulin IV|Glucose^3H pre dose insulin IV
C2706826|T201|COMP|54263-9|LNC|Glucose^30M post dose insulin IV|Glucose^30M post dose insulin IV
C2706827|T201|COMP|54264-7|LNC|Glucose^45M post dose insulin IV|Glucose^45M post dose insulin IV
C2706828|T201|COMP|54265-4|LNC|Glucose^1H post dose insulin IV|Glucose^1H post dose insulin IV
C2706829|T201|COMP|54266-2|LNC|Glucose^1.3H post dose insulin IV|Glucose^1.3H post dose insulin IV
C2706830|T201|COMP|54267-0|LNC|Glucose^1.5H post dose insulin IV|Glucose^1.5H post dose insulin IV
C2706831|T201|COMP|54268-8|LNC|Glucose^pre dose ornithine alpha-ketoglutarate|Glucose^pre dose ornithine alpha-ketoglutarate
C2706841|T201|COMP|54278-7|LNC|Glutarate|Glutarate
C2706842|T201|COMP|54279-5|LNC|Glutarylcarnitine (C5-DC)/Creatinine|Glutarylcarnitine (C5-DC)/Creatinine
C2706844|T201|COMP|54280-3|LNC|Glutarylcarnitine (C5-DC)|Glutarylcarnitine (C5-DC)
C2706845|T201|COMP|54281-1|LNC|Glutarylcarnitine (C5-DC)|Glutarylcarnitine (C5-DC)
C2706846|T201|COMP|54282-9|LNC|Glutarylcarnitine (C5-DC)|Glutarylcarnitine (C5-DC)
C2706847|T201|COMP|54283-7|LNC|Glycerol|Glycerol
C2706848|T201|COMP|54284-5|LNC|Glycerol|Glycerol
C2706849|T201|COMP|54285-2|LNC|Glycerol|Glycerol
C2706850|T201|COMP|54286-0|LNC|Glycolate|Glycolate
C2706851|T201|COMP|54287-8|LNC|Guanidinoacetate|Guanidinoacetate
C2706852|T201|COMP|54288-6|LNC|Guanidinoacetate|Guanidinoacetate
C2706853|T201|COMP|54289-4|LNC|Hemoglobin|Hemoglobin
C2706854|T201|COMP|54290-2|LNC|Heptanoylcarnitine (C7)/Creatinine|Heptanoylcarnitine (C7)/Creatinine
C2706856|T201|COMP|54291-0|LNC|Heptanoylcarnitine (C7)|Heptanoylcarnitine (C7)
C2706857|T201|COMP|54292-8|LNC|Heptanoylcarnitine (C7)|Heptanoylcarnitine (C7)
C2706858|T201|COMP|54293-6|LNC|Heptanoylcarnitine (C7)|Heptanoylcarnitine (C7)
C2706859|T201|COMP|54294-4|LNC|Fatty acids.very long chain.C26:0/Creatinine|Fatty acids.very long chain.C26:0/Creatinine
C2706861|T201|COMP|54295-1|LNC|Hexanoylcarnitine (C6)/Creatinine|Hexanoylcarnitine (C6)/Creatinine
C2706863|T201|COMP|54296-9|LNC|Hexanoylcarnitine (C6)|Hexanoylcarnitine (C6)
C2706864|T201|COMP|54297-7|LNC|Hexanoylcarnitine (C6)|Hexanoylcarnitine (C6)
C2706865|T201|COMP|54298-5|LNC|Hexanoylcarnitine (C6)|Hexanoylcarnitine (C6)
C2706866|T201|COMP|54299-3|LNC|Homocitrulline|Homocitrulline
C2706867|T201|COMP|54301-7|LNC|Homocysteine|Homocysteine
C2706868|T201|COMP|54302-5|LNC|Homocystine|Homocystine
C2706869|T201|COMP|54303-3|LNC|Hydroxylysine|Hydroxylysine
C2706870|T201|COMP|54304-1|LNC|Isobutyrylglycine|Isobutyrylglycine
C2706871|T201|COMP|54305-8|LNC|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)
C2706872|T201|COMP|54306-6|LNC|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)
C2706873|T201|COMP|54307-4|LNC|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)
C2706874|T201|COMP|54308-2|LNC|Isovalerylglycine|Isovalerylglycine
C2706875|T201|COMP|54309-0|LNC|Lactate/Pyruvate|Lactate/Pyruvate
C2706876|T201|COMP|54310-8|LNC|Linoleoylcarnitine (C18:2)/Creatinine|Linoleoylcarnitine (C18:2)/Creatinine
C2706878|T201|COMP|54311-6|LNC|Linoleoylcarnitine (C18:2)|Linoleoylcarnitine (C18:2)
C2706879|T201|COMP|54312-4|LNC|Linoleoylcarnitine (C18:2)|Linoleoylcarnitine (C18:2)
C2706880|T201|COMP|54313-2|LNC|Linoleoylcarnitine (C18:2)|Linoleoylcarnitine (C18:2)
C2706881|T201|COMP|54314-0|LNC|Malonylcarnitine (C3-DC)/Creatinine|Malonylcarnitine (C3-DC)/Creatinine
C2706883|T201|COMP|54315-7|LNC|Methylmalonate|Methylmalonate
C2706884|T201|COMP|54316-5|LNC|Methylmalonylcarnitine (C4-DC)/Creatinine|Methylmalonylcarnitine (C4-DC)/Creatinine
C2706886|T201|COMP|54317-3|LNC|Methylmalonylcarnitine (C4-DC)|Methylmalonylcarnitine (C4-DC)
C2706887|T201|COMP|54318-1|LNC|Methylmalonylcarnitine (C4-DC)|Methylmalonylcarnitine (C4-DC)
C2706888|T201|COMP|54319-9|LNC|Methylmalonylcarnitine (C4-DC)|Methylmalonylcarnitine (C4-DC)
C2706889|T201|COMP|54320-7|LNC|Octanoylcarnitine (C8)/Creatinine|Octanoylcarnitine (C8)/Creatinine
C2706891|T201|COMP|54321-5|LNC|Octanoylcarnitine (C8)|Octanoylcarnitine (C8)
C2706892|T201|COMP|54322-3|LNC|Octanoylcarnitine (C8)|Octanoylcarnitine (C8)
C2706893|T201|COMP|54323-1|LNC|Palmitoylcarnitine (C16)/Creatinine|Palmitoylcarnitine (C16)/Creatinine
C2706895|T201|COMP|54324-9|LNC|Palmitoylcarnitine (C16)|Palmitoylcarnitine (C16)
C2706896|T201|COMP|54325-6|LNC|Palmitoylcarnitine (C16)|Palmitoylcarnitine (C16)
C2706897|T201|COMP|54326-4|LNC|Phosphoethanolamine|Phosphoethanolamine
C2706898|T201|COMP|54327-2|LNC|Pipecolate|Pipecolate
C2706899|T201|COMP|54328-0|LNC|Pipecolate|Pipecolate
C2706900|T201|COMP|54494-0|LNC|Chloride|Chloride
C2706901|T201|COMP|54495-7|LNC|Glucose^post dialysis|Glucose^post dialysis
C2706902|T201|COMP|54496-5|LNC|Glucose^5th specimen post XXX challenge|Glucose^5th specimen post XXX challenge
C2706903|T201|COMP|54497-3|LNC|Glucose^6th specimen post XXX challenge|Glucose^6th specimen post XXX challenge
C2706904|T201|COMP|54498-1|LNC|Glucose^7th specimen post XXX challenge|Glucose^7th specimen post XXX challenge
C2706905|T201|COMP|54499-9|LNC|Glucose^8th specimen post XXX challenge|Glucose^8th specimen post XXX challenge
C2706924|T201|COMP|55621-7|LNC|Bambermycins|Bambermycins
C2706925|T201|COMP|55622-5|LNC|Butirosin|Butirosin
C2706926|T201|COMP|55623-3|LNC|Capreomycin|Capreomycin
C2706927|T201|COMP|55624-1|LNC|Cefacetrile|Cefacetrile
C2706928|T201|COMP|55625-8|LNC|Cefacetrile|Cefacetrile
C2706929|T201|COMP|55626-6|LNC|Cefacetrile|Cefacetrile
C2706930|T201|COMP|55627-4|LNC|Cefacetrile|Cefacetrile
C2706977|T201|COMP|54916-2|LNC|Lophius piscatorius Ab.IgE|Lophius piscatorius Ab.IgE
C2706979|T201|COMP|54917-0|LNC|Lysozyme|Lysozyme
C2706980|T201|COMP|54918-8|LNC|Ma+Ta Ab|Ma+Ta Ab
C2706981|T201|COMP|54919-6|LNC|Magnesium|Magnesium
C2706982|T201|COMP|54920-4|LNC|Myrmecia pilosula Ab.IgE|Myrmecia pilosula Ab.IgE
C2706984|T201|COMP|54921-2|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C2706985|T201|COMP|54922-0|LNC|Phosphate|Phosphate
C2706998|T201|COMP|55178-8|LNC|Calcium phosphate crystals|Calcium phosphate crystals
C2706999|T201|COMP|55179-6|LNC|Sodium urate crystals|Sodium urate crystals
C2707000|T201|COMP|55180-4|LNC|Human epididymis protein 4|Human epididymis protein 4
C2707067|T201|COMP|54329-8|LNC|Propionylcarnitine (C3)/Creatinine|Propionylcarnitine (C3)/Creatinine
C2707069|T201|COMP|54330-6|LNC|Propionylcarnitine (C3)|Propionylcarnitine (C3)
C2707070|T201|COMP|54331-4|LNC|Propionylcarnitine (C3)|Propionylcarnitine (C3)
C2707071|T201|COMP|54332-2|LNC|Propionylglycine|Propionylglycine
C2707072|T201|COMP|54333-0|LNC|Stearoylcarnitine (C18)/Creatinine|Stearoylcarnitine (C18)/Creatinine
C2707074|T201|COMP|54334-8|LNC|Stearoylcarnitine (C18)|Stearoylcarnitine (C18)
C2707075|T201|COMP|54335-5|LNC|Stearoylcarnitine (C18)|Stearoylcarnitine (C18)
C2707076|T201|COMP|54336-3|LNC|Sulfocysteine|Sulfocysteine
C2707077|T201|COMP|54337-1|LNC|Sulfocysteine|Sulfocysteine
C2707078|T201|COMP|54338-9|LNC|Tetradecanoylcarnitine (C14)/Creatinine|Tetradecanoylcarnitine (C14)/Creatinine
C2707080|T201|COMP|54339-7|LNC|Tetradecanoylcarnitine (C14)|Tetradecanoylcarnitine (C14)
C2707081|T201|COMP|54340-5|LNC|Tetradecanoylcarnitine (C14)|Tetradecanoylcarnitine (C14)
C2707082|T201|COMP|54341-3|LNC|Myristoleate/Creatinine|Myristoleate/Creatinine
C2707084|T201|COMP|54342-1|LNC|Tiglylglycine|Tiglylglycine
C2707085|T201|COMP|54343-9|LNC|3-Methoxytyramine/Creatinine|3-Methoxytyramine/Creatinine
C2707086|T201|COMP|54344-7|LNC|3-Methoxytyramine|3-Methoxytyramine
C2707087|T201|COMP|54345-4|LNC|Acetylcarnitine (C2)|Acetylcarnitine (C2)
C2707088|T201|COMP|54346-2|LNC|Albumin|Albumin
C2707089|T201|COMP|54347-0|LNC|Albumin|Albumin
C2707090|T201|COMP|54348-8|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C2707091|T201|COMP|54349-6|LNC|Ammonia|Ammonia
C2707092|T201|COMP|54350-4|LNC|Ascorbate+Dehydroascorbate|Ascorbate+Dehydroascorbate
C2707093|T201|COMP|54351-2|LNC|Ascorbate+Dehydroascorbate|Ascorbate+Dehydroascorbate
C2707094|T201|COMP|54352-0|LNC|Nitrogen|Nitrogen
C2707095|T201|COMP|54353-8|LNC|Beta 1 globulin|Beta 1 globulin
C2707096|T201|COMP|54354-6|LNC|Beta 2 globulin|Beta 2 globulin
C2707099|T201|COMP|54356-1|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C2707100|T201|COMP|54357-9|LNC|Beta 2 globulin+Gamma globulin/Protein.total|Beta 2 globulin+Gamma globulin/Protein.total
C2707101|T201|COMP|54358-7|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C2707102|T201|COMP|54359-5|LNC|Bicarbonate^post dialysis|Bicarbonate^post dialysis
C2707103|T201|COMP|54360-3|LNC|Bicarbonate|Bicarbonate
C2707104|T201|COMP|54361-1|LNC|Bicarbonate|Bicarbonate
C2707105|T201|COMP|54380-1|LNC|Cystatin C|Cystatin C
C2707106|T201|COMP|54381-9|LNC|Cystatin C|Cystatin C
C2707107|T201|COMP|54382-7|LNC|Cytochrome C oxidase|Cytochrome C oxidase
C2707108|T201|COMP|54383-5|LNC|Cytochrome C oxidase|Cytochrome C oxidase
C2707109|T201|COMP|54384-3|LNC|Cytochrome C oxidase|Cytochrome C oxidase
C2707110|T201|COMP|54385-0|LNC|Dehydroascorbate/Ascorbate|Dehydroascorbate/Ascorbate
C2707112|T201|COMP|54386-8|LNC|Dehydroascorbate|Dehydroascorbate
C2707113|T201|COMP|54387-6|LNC|Dihydroxycholestanoate|Dihydroxycholestanoate
C2707114|T201|COMP|54388-4|LNC|Dihydroxycholestanoate|Dihydroxycholestanoate
C2707115|T201|COMP|54389-2|LNC|Dodecanoylcarnitine (C12)|Dodecanoylcarnitine (C12)
C2707116|T201|COMP|54390-0|LNC|Fibroblast growth factor 23.intact|Fibroblast growth factor 23.intact
C2707117|T201|COMP|54391-8|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C2707118|T201|COMP|54392-6|LNC|Glucose^1st specimen post XXX challenge|Glucose^1st specimen post XXX challenge
C2707119|T201|COMP|54393-4|LNC|Glucose^10th specimen post XXX challenge|Glucose^10th specimen post XXX challenge
C2707120|T201|COMP|54394-2|LNC|Glucose^11th specimen post XXX challenge|Glucose^11th specimen post XXX challenge
C2707121|T201|COMP|54395-9|LNC|Glucose^12th specimen post XXX challenge|Glucose^12th specimen post XXX challenge
C2707122|T201|COMP|54396-7|LNC|Glucose^2nd specimen post XXX challenge|Glucose^2nd specimen post XXX challenge
C2707123|T201|COMP|54397-5|LNC|Glucose^3rd specimen post XXX challenge|Glucose^3rd specimen post XXX challenge
C2707124|T201|COMP|54398-3|LNC|Glucose^4th specimen post XXX challenge|Glucose^4th specimen post XXX challenge
C2707125|T201|COMP|54399-1|LNC|Glucose^9th specimen post XXX challenge|Glucose^9th specimen post XXX challenge
C2707126|T201|COMP|54400-7|LNC|Glucose^pre dose glucagon|Glucose^pre dose glucagon
C2707127|T201|COMP|54401-5|LNC|Glucose^10M post dose glucagon|Glucose^10M post dose glucagon
C2707128|T201|COMP|54402-3|LNC|4-Hydroxymidazolam|4-Hydroxymidazolam
C2707129|T201|COMP|54403-1|LNC|Transfuse 5% plasma protein fraction units|Transfuse 5% plasma protein fraction units
C2707130|T201|COMP|54404-9|LNC|Pooled platelet concentrate units given|Pooled platelet concentrate units given
C2707131|T201|COMP|54405-6|LNC|Transfuse pooled cryoprecipitate units|Transfuse pooled cryoprecipitate units
C2707132|T201|COMP|54406-4|LNC|Pooled cryoprecipitate units given|Pooled cryoprecipitate units given
C2707133|T201|COMP|54407-2|LNC|Transfuse pooled fresh frozen plasma units|Transfuse pooled fresh frozen plasma units
C2707134|T201|COMP|54408-0|LNC|Pooled fresh frozen plasma units given|Pooled fresh frozen plasma units given
C2707137|T201|COMP|54411-4|LNC|Rh immune globulin given|Rh immune globulin given
C2707139|T201|COMP|54412-2|LNC|Cryoprecipitate poor plasma units given|Cryoprecipitate poor plasma units given
C2707141|T201|COMP|54413-0|LNC|Transfuse leukocyte-poor plateletpheresis units|Transfuse leukocyte-poor plateletpheresis units
C2707142|T201|COMP|54414-8|LNC|Leukocyte-poor plateletpheresis units given|Leukocyte-poor plateletpheresis units given
C2707143|T201|COMP|54415-5|LNC|Transfuse leukocyte-poor platelets units|Transfuse leukocyte-poor platelets units
C2707144|T201|COMP|54416-3|LNC|Rh|Rh
C2707145|T201|COMP|54417-1|LNC|ABO & Rh group|ABO & Rh group
C2707146|T201|COMP|54418-9|LNC|Transfuse fresh frozen plasma pediatric units|Transfuse fresh frozen plasma pediatric units
C2707148|T201|COMP|54419-7|LNC|Whole blood pediatric units given|Whole blood pediatric units given
C2707150|T201|COMP|54420-5|LNC|Frozen erythrocytes newborn units given|Frozen erythrocytes newborn units given
C2707152|T201|COMP|54421-3|LNC|Transfuse frozen erythrocytes pediatric units|Transfuse frozen erythrocytes pediatric units
C2707154|T201|COMP|54422-1|LNC|Frozen erythrocytes pediatric units given|Frozen erythrocytes pediatric units given
C2707156|T201|COMP|54423-9|LNC|Transfuse plateletpheresis half units|Transfuse plateletpheresis half units
C2707157|T201|COMP|54424-7|LNC|Plateletpheresis half units given|Plateletpheresis half units given
C2707159|T201|COMP|54425-4|LNC|D little u Ag|D little u Ag
C2707160|T201|COMP|54426-2|LNC|Fresh frozen plasma pediatric units given|Fresh frozen plasma pediatric units given
C2707162|T201|COMP|54427-0|LNC|Transfuse frozen erythrocytes newborn units|Transfuse frozen erythrocytes newborn units
C2707163|T201|COMP|54428-8|LNC|Frozen packed erythrocytes given|Frozen packed erythrocytes given
C2707165|T201|COMP|54429-6|LNC|5% plasma protein fraction given|5% plasma protein fraction given
C2707166|T201|COMP|54430-4|LNC|Pooled platelets given|Pooled platelets given
C2707168|T201|COMP|54431-2|LNC|Pooled cryoprecipitate given|Pooled cryoprecipitate given
C2707170|T201|COMP|54432-0|LNC|Pooled fresh frozen plasma given|Pooled fresh frozen plasma given
C2707174|T201|COMP|54434-6|LNC|Lipoprotein.beta.subparticle|Lipoprotein.beta.subparticle
C2707176|T201|COMP|54435-3|LNC|Aspergillus fumigatus Ab|Aspergillus fumigatus Ab
C2707177|T201|COMP|54436-1|LNC|Urate dihydrate/Total|Urate dihydrate/Total
C2707179|T201|COMP|54437-9|LNC|Sodium urate/Total|Sodium urate/Total
C2707180|T201|COMP|54438-7|LNC|Cholesterol/Total|Cholesterol/Total
C2707181|T201|COMP|54439-5|LNC|Calcium bilirubinate/Total|Calcium bilirubinate/Total
C2707182|T201|COMP|54440-3|LNC|Newberyite/Total|Newberyite/Total
C2707183|T201|COMP|54441-1|LNC|Lipoprotein goals|Lipoprotein goals
C2707185|T201|COMP|54442-9|LNC|Carnitine esters/Carnitine.free (C0)|Carnitine esters/Carnitine.free (C0)
C2707186|T201|COMP|54451-0|LNC|CYP2C9 & VKORC1|CYP2C9 & VKORC1
C2707188|T201|COMP|54452-8|LNC|Ferning|Ferning
C2707189|T201|COMP|54453-6|LNC|Test method|Test method
C2707191|T201|COMP|54454-4|LNC|Arsenic fractions panel|Arsenic fractions panel
C2707193|T201|COMP|54455-1|LNC|Blastomyces dermatitidis Ag|Blastomyces dermatitidis Ag
C2707194|T201|COMP|54456-9|LNC|Urea reduction ratio|Urea reduction ratio
C2707195|T201|COMP|54457-7|LNC|Biotinidase|Biotinidase
C2707196|T201|COMP|54458-5|LNC|Granulocyte colony stimulating factor|Granulocyte colony stimulating factor
C2707197|T201|COMP|54459-3|LNC|Dicarboxypalmitoylcarnitine (C16-DC)/Creatinine|Dicarboxypalmitoylcarnitine (C16-DC)/Creatinine
C2707199|T201|COMP|54460-1|LNC|Malonylcarnitine (C3-DC)|Malonylcarnitine (C3-DC)
C2707200|T201|COMP|54461-9|LNC|Malonylcarnitine (C3-DC)|Malonylcarnitine (C3-DC)
C2707201|T201|COMP|54462-7|LNC|Malonylcarnitine (C3-DC)|Malonylcarnitine (C3-DC)
C2707202|T201|COMP|54463-5|LNC|Malonylcarnitine (C3-DC)|Malonylcarnitine (C3-DC)
C2707203|T201|COMP|54464-3|LNC|Albumin/Protein.total|Albumin/Protein.total
C2707204|T201|COMP|54465-0|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C2707205|T201|COMP|54466-8|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C2707206|T201|COMP|54467-6|LNC|Cholesterol.in HDL 2a/Cholesterol.in HDL.total|Cholesterol.in HDL 2a/Cholesterol.in HDL.total
C2707208|T201|COMP|54468-4|LNC|Cholesterol.in HDL 2b/Cholesterol.in HDL.total|Cholesterol.in HDL 2b/Cholesterol.in HDL.total
C2707210|T201|COMP|54469-2|LNC|Cholesterol.in HDL 3a/Cholesterol.in HDL.total|Cholesterol.in HDL 3a/Cholesterol.in HDL.total
C2707212|T201|COMP|54470-0|LNC|Cholesterol.in HDL 3b/Cholesterol.in HDL.total|Cholesterol.in HDL 3b/Cholesterol.in HDL.total
C2707214|T201|COMP|54471-8|LNC|Cholesterol.in HDL 3c/Cholesterol.in HDL.total|Cholesterol.in HDL 3c/Cholesterol.in HDL.total
C2707216|T201|COMP|54472-6|LNC|Amylase.macromolecular/Amylase.total|Amylase.macromolecular/Amylase.total
C2707218|T201|COMP|54473-4|LNC|Pimeloylcarnitine (C7-DC)|Pimeloylcarnitine (C7-DC)
C2707220|T201|COMP|54474-2|LNC|Pimeloylcarnitine (C7-DC)|Pimeloylcarnitine (C7-DC)
C2707221|T201|COMP|54475-9|LNC|Pimeloylcarnitine (C7-DC)|Pimeloylcarnitine (C7-DC)
C2707222|T201|COMP|54476-7|LNC|Pimeloylcarnitine (C7-DC)|Pimeloylcarnitine (C7-DC)
C2707223|T201|COMP|54477-5|LNC|Dicarboxypalmitoylcarnitine (C16-DC)|Dicarboxypalmitoylcarnitine (C16-DC)
C2707224|T201|COMP|54478-3|LNC|Dicarboxypalmitoylcarnitine (C16-DC)|Dicarboxypalmitoylcarnitine (C16-DC)
C2707227|T201|COMP|54480-9|LNC|Dicarboxypalmitoylcarnitine (C16-DC)|Dicarboxypalmitoylcarnitine (C16-DC)
C2707228|T201|COMP|54481-7|LNC|Dicarboxystearoylcarnitine (C18-DC)/Creatinine|Dicarboxystearoylcarnitine (C18-DC)/Creatinine
C2707230|T201|COMP|54482-5|LNC|Dicarboxystearoylcarnitine (C18-DC)|Dicarboxystearoylcarnitine (C18-DC)
C2707231|T201|COMP|54483-3|LNC|Dicarboxystearoylcarnitine (C18-DC)|Dicarboxystearoylcarnitine (C18-DC)
C2707232|T201|COMP|54484-1|LNC|Octadecanedioylcarnitine (C18-DC)|Octadecanedioylcarnitine (C18-DC)
C2707234|T201|COMP|54485-8|LNC|Dicarboxystearoylcarnitine (C18-DC)|Dicarboxystearoylcarnitine (C18-DC)
C2707235|T201|COMP|54486-6|LNC|Glucose|Glucose
C2707236|T201|COMP|54487-4|LNC|Glucose|Glucose
C2707237|T201|COMP|54488-2|LNC|Pimeloylcarnitine (C7-DC)/Creatinine|Pimeloylcarnitine (C7-DC)/Creatinine
C2707239|T201|COMP|54489-0|LNC|Phosphoserine|Phosphoserine
C2707240|T201|COMP|54490-8|LNC|Pipecolate|Pipecolate
C2707241|T201|COMP|54491-6|LNC|Alanine aminotransferase|Alanine aminotransferase
C2707242|T201|COMP|54492-4|LNC|Alanine aminotransferase|Alanine aminotransferase
C2707243|T201|COMP|54493-2|LNC|Allantoine|Allantoine
C2707378|T201|COMP|54908-9|LNC|Cefminox|Cefminox
C2707379|T201|COMP|54909-7|LNC|Culex pipiens Ab.IgE|Culex pipiens Ab.IgE
C2707381|T201|COMP|54910-5|LNC|DNA double strand Ab|DNA double strand Ab
C2707382|T201|COMP|54911-3|LNC|Epinephelus lanceolatus Ab.IgE|Epinephelus lanceolatus Ab.IgE
C2707384|T201|COMP|54912-1|LNC|Fosfomycin Ab.IgE|Fosfomycin Ab.IgE
C2707386|T201|COMP|54913-9|LNC|Gentamicin Ab.IgE|Gentamicin Ab.IgE
C2707388|T201|COMP|54914-7|LNC|Hepatitis C virus core Ag|Hepatitis C virus core Ag
C2707389|T201|COMP|54915-4|LNC|Chlorophora excelsa Ab.IgE|Chlorophora excelsa Ab.IgE
C2707395|T201|COMP|55540-9|LNC|Furosemide|Furosemide
C2707396|T201|COMP|55541-7|LNC|hydroCHLOROthiazide|hydroCHLOROthiazide
C2707397|T201|COMP|55542-5|LNC|Hydroxybupropion|Hydroxybupropion
C2707398|T201|COMP|55543-3|LNC|Hydroxychloroquine|Hydroxychloroquine
C2707521|T201|COMP|55189-5|LNC|Cefotaxime|Cefotaxime
C2707522|T201|COMP|55190-3|LNC|cefTRIAXone|cefTRIAXone
C2707523|T201|COMP|55192-9|LNC|Chromosome analysis.interphase|Chromosome analysis.interphase
C2707524|T201|COMP|55193-7|LNC|Chromosome analysis.interphase|Chromosome analysis.interphase
C2707525|T201|COMP|55449-3|LNC|Fibrin D-dimer|Fibrin D-dimer
C2707526|T201|COMP|55450-1|LNC|Fibrin+Fibrinogen fragments|Fibrin+Fibrinogen fragments
C2707527|T201|COMP|55451-9|LNC|Fibrin+Fibrinogen fragments|Fibrin+Fibrinogen fragments
C2707528|T201|COMP|55452-7|LNC|Fibrinogen|Fibrinogen
C2707529|T201|COMP|55453-5|LNC|Haptoglobin|Haptoglobin
C2707530|T201|COMP|55454-3|LNC|Hemoglobin A1c|Hemoglobin A1c
C2707531|T201|COMP|55455-0|LNC|Hemoglobin F|Hemoglobin F
C2707532|T201|COMP|55458-4|LNC|Interferon.alpha|Interferon.alpha
C2707535|T201|COMP|55614-2|LNC|Amoxicillin+Sulbactam|Amoxicillin+Sulbactam
C2707537|T201|COMP|55615-9|LNC|Amoxicillin+Sulbactam|Amoxicillin+Sulbactam
C2707538|T201|COMP|55616-7|LNC|Amoxicillin+Sulbactam|Amoxicillin+Sulbactam
C2707539|T201|COMP|55617-5|LNC|Antibiotic XXX|Antibiotic XXX
C2707540|T201|COMP|55618-3|LNC|Atovaquone|Atovaquone
C2707541|T201|COMP|55619-1|LNC|Avilamycin|Avilamycin
C2707542|T201|COMP|55620-9|LNC|Bacampicillin|Bacampicillin
C2707629|T201|COMP|54900-6|LNC|IgA|IgA
C2707630|T201|COMP|54901-4|LNC|IgG|IgG
C2707631|T201|COMP|54902-2|LNC|IgM|IgM
C2707634|T201|COMP|54905-5|LNC|Norovirus Genogroup I RNA|Norovirus Genogroup I RNA
C2707636|T201|COMP|54906-3|LNC|Norovirus Genogroup II RNA|Norovirus Genogroup II RNA
C2707638|T201|COMP|54907-1|LNC|Alkaline phosphatase|Alkaline phosphatase
C2707641|T201|COMP|55090-5|LNC|Cells.CD3-CD56+/100 cells|Cells.CD3-CD56+/100 cells
C2707642|T201|COMP|55091-3|LNC|Darunavir|Darunavir
C2707643|T201|COMP|55092-1|LNC|PDGFRA gene rearrangements|PDGFRA gene rearrangements
C2707648|T201|COMP|55095-4|LNC|Adenovirus|Adenovirus
C2707649|T201|COMP|55096-2|LNC|Nocardia sp identified|Nocardia sp identified
C2707650|T201|COMP|55097-0|LNC|Parainfluenza virus 1|Parainfluenza virus 1
C2707651|T201|COMP|55098-8|LNC|Parainfluenza virus 2|Parainfluenza virus 2
C2707652|T201|COMP|55099-6|LNC|Parainfluenza virus 3|Parainfluenza virus 3
C2707653|T201|COMP|55100-2|LNC|Respiratory syncytial virus|Respiratory syncytial virus
C2707654|T201|COMP|55101-0|LNC|Respiratory pathogens panel|Respiratory pathogens panel
C2707659|T201|COMP|55251-3|LNC|HBA2 gene alpha 3.7kb deletion|HBA2 gene alpha 3.7kb deletion
C2707661|T201|COMP|55252-1|LNC|Methoxsalen 0.02 mg per mL given|Methoxsalen 0.02 mg per mL given
C2707663|T201|COMP|55253-9|LNC|Heparin 10000 U per mL given|Heparin 10000 U per mL given
C2707665|T201|COMP|55254-7|LNC|Heparin 5000 U per mL given|Heparin 5000 U per mL given
C2707667|T201|COMP|55255-4|LNC|Pyridinoline panel|Pyridinoline panel
C2707991|T201|COMP|54923-8|LNC|Propyphenazone Ab.IgE|Propyphenazone Ab.IgE
C2707993|T201|COMP|54924-6|LNC|Purkinje cells Ab|Purkinje cells Ab
C2707994|T201|COMP|54925-3|LNC|Selenium|Selenium
C2707997|T201|COMP|54927-9|LNC|Tetranychus urticae Ab.IgE|Tetranychus urticae Ab.IgE
C2707999|T201|COMP|54928-7|LNC|Tinidazole|Tinidazole
C2708000|T201|COMP|54929-5|LNC|Tissue transglutaminase Ab|Tissue transglutaminase Ab
C2708001|T201|COMP|54930-3|LNC|Vicia faba Ab.IgE|Vicia faba Ab.IgE
C2708005|T201|COMP|54932-9|LNC|CEH abrine & ricinine panel|CEH abrine & ricinine panel
C2708007|T201|COMP|54933-7|LNC|Abrine|Abrine
C2708008|T201|COMP|54934-5|LNC|Ricinine|Ricinine
C2708009|T201|COMP|54935-2|LNC|1,2-Dichloroethane|1,2-Dichloroethane
C2708010|T201|COMP|54936-0|LNC|Carbon tetrachloride|Carbon tetrachloride
C2708011|T201|COMP|54937-8|LNC|Chloroform|Chloroform
C2708012|T201|COMP|54938-6|LNC|Ethyl benzene|Ethyl benzene
C2708013|T201|COMP|54939-4|LNC|Meta methylhippurate+Para methylhippurate|Meta methylhippurate+Para methylhippurate
C2708014|T201|COMP|54940-2|LNC|Styrene|Styrene
C2708015|T201|COMP|54941-0|LNC|Tungsten|Tungsten
C2708016|T201|COMP|54942-8|LNC|N-ethyldiethanolamine|N-ethyldiethanolamine
C2708018|T201|COMP|54943-6|LNC|N-methyldiethanolamine|N-methyldiethanolamine
C2708019|T201|COMP|54944-4|LNC|Monofluoroacetate|Monofluoroacetate
C2708020|T201|COMP|54945-1|LNC|Monochloroacetate|Monochloroacetate
C2708273|T201|COMP|55440-2|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C2708274|T201|COMP|55441-0|LNC|Antithrombin Ag|Antithrombin Ag
C2708275|T201|COMP|55442-8|LNC|Antithrombin|Antithrombin
C2708276|T201|COMP|55443-6|LNC|Cardiolipin Ab|Cardiolipin Ab
C2708277|T201|COMP|55444-4|LNC|Cardiolipin Ab.IgA|Cardiolipin Ab.IgA
C2708278|T201|COMP|55445-1|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C2708279|T201|COMP|55446-9|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C2708280|T201|COMP|55447-7|LNC|Coagulation factor VIII Ag|Coagulation factor VIII Ag
C2708281|T201|COMP|55448-5|LNC|Complement total hemolytic CH50|Complement total hemolytic CH50
C2708295|T201|COMP|55116-8|LNC|CEH volatile organic compounds panel|CEH volatile organic compounds panel
C2708297|T201|COMP|55117-6|LNC|CEH trace metals screen panel|CEH trace metals screen panel
C2708299|T201|COMP|55118-4|LNC|CEH trace metals panel|CEH trace metals panel
C2708301|T201|COMP|55119-2|LNC|CEH nitrogen mustard metabolite panel|CEH nitrogen mustard metabolite panel
C2708303|T201|COMP|55120-0|LNC|CEH metabolic toxin panel|CEH metabolic toxin panel
C2708305|T201|COMP|55121-8|LNC|Multiple sclerosis panel|Multiple sclerosis panel
C2708323|T201|COMP|55133-3|LNC|Influenza virus A hemagglutinin cDNA|Influenza virus A hemagglutinin cDNA
C2708324|T201|COMP|55134-1|LNC|Influenza virus A neuraminidase RNA|Influenza virus A neuraminidase RNA
C2708325|T201|COMP|55135-8|LNC|BCR-ABL1 kinase domain targeted mutation analysis|BCR-ABL1 kinase domain targeted mutation analysis
C2708327|T201|COMP|55136-6|LNC|Penicillin.parenteral|Penicillin.parenteral
C2708329|T201|COMP|55137-4|LNC|Penicillin.parenteral|Penicillin.parenteral
C2708331|T201|COMP|55138-2|LNC|Cortisol^post dose dexamethasone PO overnight|Cortisol^post dose dexamethasone PO overnight
C2708332|T201|COMP|55139-0|LNC|SCN5A gene targeted mutation analysis|SCN5A gene targeted mutation analysis
C2708336|T201|COMP|55141-6|LNC|Fc epsilon RI + RII Ab|Fc epsilon RI + RII Ab
C2708338|T201|COMP|55142-4|LNC|Cache valley virus RNA|Cache valley virus RNA
C2708339|T201|COMP|55143-2|LNC|California serogroup virus RNA|California serogroup virus RNA
C2708340|T201|COMP|55144-0|LNC|Powassan virus RNA|Powassan virus RNA
C2708341|T201|COMP|55145-7|LNC|Saint Louis encephalitis virus RNA|Saint Louis encephalitis virus RNA
C2708346|T201|COMP|55148-1|LNC|BCR-ABL1 b2a2+b3a2 fusion transcript|BCR-ABL1 b2a2+b3a2 fusion transcript
C2708347|T201|COMP|55149-9|LNC|BCR-ABL1 e1a2 fusion protein|BCR-ABL1 e1a2 fusion protein
C2708348|T201|COMP|55150-7|LNC|Anaplasma phagocytophilum Ab.IgG & IgM panel|Anaplasma phagocytophilum Ab.IgG & IgM panel
C2708350|T201|COMP|55151-5|LNC|Aldosterone & renin activity panel|Aldosterone & renin activity panel
C2708352|T201|COMP|55152-3|LNC|Amiodarone & Desethylamiodarone panel|Amiodarone & Desethylamiodarone panel
C2708354|T201|COMP|55153-1|LNC|Biotinidase panel|Biotinidase panel
C2708356|T201|COMP|55154-9|LNC|Ethambutol+rifAMPin|Ethambutol+rifAMPin
C2708357|T201|COMP|55155-6|LNC|Flunitrazepam & 7-Aminoflunitrazepam panel|Flunitrazepam & 7-Aminoflunitrazepam panel
C2708359|T201|COMP|55156-4|LNC|Minocycline|Minocycline
C2708360|T201|COMP|55157-2|LNC|Risperidone & 9-Hydroxyrisperidone panel|Risperidone & 9-Hydroxyrisperidone panel
C2708362|T201|COMP|55158-0|LNC|Tigecycline|Tigecycline
C2708363|T201|COMP|55159-8|LNC|Ursodeoxycholate|Ursodeoxycholate
C2708364|T201|COMP|55160-6|LNC|Adenovirus Ab.IgG & IgM panel|Adenovirus Ab.IgG & IgM panel
C2708366|T201|COMP|55161-4|LNC|Bordetella pertussis Ab.IgA & IgG panel|Bordetella pertussis Ab.IgA & IgG panel
C2708368|T201|COMP|55162-2|LNC|HTLV I+II Ab panel|HTLV I+II Ab panel
C2708370|T201|COMP|55163-0|LNC|Streptococcus pyogenes enzyme Ab panel|Streptococcus pyogenes enzyme Ab panel
C2708372|T201|COMP|55164-8|LNC|Paroxysmal nocturnal panel|Paroxysmal nocturnal panel
C2708374|T201|COMP|55165-5|LNC|Echinococcus sp Ab.IgG4|Echinococcus sp Ab.IgG4
C2708375|T201|COMP|55166-3|LNC|Hepatitis G virus E2 Ab|Hepatitis G virus E2 Ab
C2708377|T201|COMP|55167-1|LNC|Mycoplasma sp Ab|Mycoplasma sp Ab
C2708382|T201|COMP|55170-5|LNC|Cytoplasmic Ab|Cytoplasmic Ab
C2708383|T201|COMP|55171-3|LNC|Cytoplasmic Ab pattern|Cytoplasmic Ab pattern
C2708390|T201|COMP|55194-5|LNC|Ciprofloxacin 1.0 ug/mL|Ciprofloxacin 1.0 ug/mL
C2708392|T201|COMP|55195-2|LNC|DHCR7 gene targeted mutation analysis|DHCR7 gene targeted mutation analysis
C2708394|T201|COMP|55196-0|LNC|Terconazole|Terconazole
C2708395|T201|COMP|55197-8|LNC|Transfusion status|Transfusion status
C2708397|T201|COMP|55198-6|LNC|Zygosity|Zygosity
C2708399|T201|COMP|55199-4|LNC|Cells karyotyped.total|Cells karyotyped.total
C2708401|T201|COMP|55200-0|LNC|Carnitine|Carnitine
C2708402|T201|COMP|55201-8|LNC|KIT gene targeted mutation analysis|KIT gene targeted mutation analysis
C2708406|T201|COMP|55204-2|LNC|Macroamylase|Macroamylase
C2708407|T201|COMP|55205-9|LNC|Vasoactive intestinal peptide|Vasoactive intestinal peptide
C2708408|T201|COMP|55206-7|LNC|Platelet mass|Platelet mass
C2708410|T201|COMP|55207-5|LNC|Genetic analysis discrete result panel|Genetic analysis discrete result panel
C2708412|T201|COMP|55208-3|LNC|DNA analysis discrete sequence variation panel|DNA analysis discrete sequence variation panel
C2708434|T201|COMP|55219-0|LNC|Antioxidants|Antioxidants
C2708435|T201|COMP|55220-8|LNC|Asialoglycoprotein receptor Ab|Asialoglycoprotein receptor Ab
C2708437|T201|COMP|55221-6|LNC|Carbohydrates|Carbohydrates
C2708439|T201|COMP|55223-2|LNC|Mycobacterium tuberculosis A60 Ab.IgM|Mycobacterium tuberculosis A60 Ab.IgM
C2708441|T201|COMP|55224-0|LNC|Mycobacterium tuberculosis A60 Ab|Mycobacterium tuberculosis A60 Ab
C2708443|T201|COMP|55225-7|LNC|Aucoumea klaineana Ab.IgE|Aucoumea klaineana Ab.IgE
C2708445|T201|COMP|55226-5|LNC|Pancreatic polypeptide|Pancreatic polypeptide
C2708446|T201|COMP|55227-3|LNC|Entandrophragma cylindricum Ab.IgE|Entandrophragma cylindricum Ab.IgE
C2708451|T201|COMP|55231-5|LNC|Electrolytes panel|Electrolytes panel
C2708452|T201|COMP|55232-3|LNC|Genetic analysis summary panel|Genetic analysis summary panel
C2708454|T201|COMP|55233-1|LNC|Genetic analysis master panel|Genetic analysis master panel
C2708456|T201|COMP|55234-9|LNC|Alpha thalassemia gene panel|Alpha thalassemia gene panel
C2708458|T201|COMP|55235-6|LNC|Abnormal hemoglobin gene panel|Abnormal hemoglobin gene panel
C2708460|T201|COMP|55236-4|LNC|HBA2 gene alpha 4.2kb deletion|HBA2 gene alpha 4.2kb deletion
C2708462|T201|COMP|55237-2|LNC|HBA2 gene.c.427T>C|HBA2 gene.c.427T>C
C2708464|T201|COMP|55238-0|LNC|HBA2 gene.c.429A>T|HBA2 gene.c.429A>T
C2708466|T201|COMP|55239-8|LNC|HBB gene.c.441_442insAC|HBB gene.c.441_442insAC
C2708468|T201|COMP|55240-6|LNC|HBB gene.c.251G>A|HBB gene.c.251G>A
C2708470|T201|COMP|55241-4|LNC|HBB gene.c.19G>A|HBB gene.c.19G>A
C2708472|T201|COMP|55242-2|LNC|HBB gene.c.20A>T|HBB gene.c.20A>T
C2708474|T201|COMP|55243-0|LNC|HBB gene.c.364G>C|HBB gene.c.364G>C
C2708476|T201|COMP|55244-8|LNC|HPFH-6 gene|HPFH-6 gene
C2708478|T201|COMP|55245-5|LNC|HBB gene.c.220G>A|HBB gene.c.220G>A
C2708480|T201|COMP|55246-3|LNC|HBA2 gene.c.84G>C|HBA2 gene.c.84G>C
C2708482|T201|COMP|55247-1|LNC|HBA1 gene.c.223G>C|HBA1 gene.c.223G>C
C2708484|T201|COMP|55248-9|LNC|HBB gene.c.79G>A|HBB gene.c.79G>A
C2708486|T201|COMP|55249-7|LNC|HBA2 gene SEA deletion|HBA2 gene SEA deletion
C2708488|T201|COMP|55250-5|LNC|HBA2 gene THAI+FIL+MED+alpha 20.5 deletion|HBA2 gene THAI+FIL+MED+alpha 20.5 deletion
C2708512|T201|COMP|55293-5|LNC|Linopristin+Flopristin|Linopristin+Flopristin
C2708513|T201|COMP|55294-3|LNC|Linopristin+Flopristin|Linopristin+Flopristin
C2708514|T201|COMP|55295-0|LNC|Protein fractions & Immunoglobulins panel|Protein fractions & Immunoglobulins panel
C2708516|T201|COMP|55296-8|LNC|CAV3 gene targeted mutation analysis|CAV3 gene targeted mutation analysis
C2708518|T201|COMP|55297-6|LNC|FIP1L1+PDGFRA gene rearrangements|FIP1L1+PDGFRA gene rearrangements
C2708520|T201|COMP|55298-4|LNC|Human papilloma virus 6+11+42+43+44 DNA|Human papilloma virus 6+11+42+43+44 DNA
C2708521|T201|COMP|55299-2|LNC|Human papilloma virus 6+11+42+43+44 DNA|Human papilloma virus 6+11+42+43+44 DNA
C2708522|T201|COMP|55300-8|LNC|JAK2 gene exon 12 targeted mutation analysis|JAK2 gene exon 12 targeted mutation analysis
C2708524|T201|COMP|55301-6|LNC|JAK2 gene exon 13 targeted mutation analysis|JAK2 gene exon 13 targeted mutation analysis
C2708526|T201|COMP|55302-4|LNC|Paraneoplastic pemphigus Ab|Paraneoplastic pemphigus Ab
C2708528|T201|COMP|55303-2|LNC|Fungus|Fungus
C2708529|T201|COMP|55304-0|LNC|Fungus|Fungus
C2708530|T201|COMP|55305-7|LNC|Fungus|Fungus
C2708531|T201|COMP|55306-5|LNC|Fungus|Fungus
C2708532|T201|COMP|55307-3|LNC|Fungus|Fungus
C2708533|T201|COMP|55308-1|LNC|Yeast.pseudohyphae|Yeast.pseudohyphae
C2708534|T201|COMP|55309-9|LNC|Yeast.pseudohyphae|Yeast.pseudohyphae
C2708535|T201|COMP|55310-7|LNC|Yeast.pseudohyphae|Yeast.pseudohyphae
C2708536|T201|COMP|55311-5|LNC|Yeast.pseudohyphae|Yeast.pseudohyphae
C2708537|T201|COMP|55312-3|LNC|Yeast.pseudohyphae|Yeast.pseudohyphae
C2708538|T201|COMP|55313-1|LNC|Yeast|Yeast
C2708539|T201|COMP|55314-9|LNC|Yeast|Yeast
C2708540|T201|COMP|55315-6|LNC|Yeast|Yeast
C2708541|T201|COMP|55316-4|LNC|Yeast|Yeast
C2708542|T201|COMP|55317-2|LNC|Yeast|Yeast
C2708543|T201|COMP|55318-0|LNC|Fungus|Fungus
C2708544|T201|COMP|55319-8|LNC|Yeast.pseudohyphae|Yeast.pseudohyphae
C2708545|T201|COMP|55320-6|LNC|Yeast|Yeast
C2708546|T201|COMP|55321-4|LNC|C little w Ab|C little w Ab
C2708547|T201|COMP|55322-2|LNC|F little y super little b Ab|F little y super little b Ab
C2708548|T201|COMP|55323-0|LNC|J little k super little a Ab|J little k super little a Ab
C2708549|T201|COMP|55324-8|LNC|J little k super little b Ab|J little k super little b Ab
C2708550|T201|COMP|55325-5|LNC|J little s super little a Ab|J little s super little a Ab
C2708551|T201|COMP|55326-3|LNC|K little p super little a Ab|K little p super little a Ab
C2708552|T201|COMP|55327-1|LNC|K little p super little b Ab|K little p super little b Ab
C2708553|T201|COMP|55328-9|LNC|L little e super little a Ab|L little e super little a Ab
C2708554|T201|COMP|55329-7|LNC|L little e super little b Ab|L little e super little b Ab
C2708555|T201|COMP|55330-5|LNC|L little u super little a Ab|L little u super little a Ab
C2708556|T201|COMP|55331-3|LNC|L little u super little b Ab|L little u super little b Ab
C2708557|T201|COMP|55332-1|LNC|little c Ab|little c Ab
C2708558|T201|COMP|55333-9|LNC|little f Ab|little f Ab
C2708559|T201|COMP|55334-7|LNC|little k Ab|little k Ab
C2708560|T201|COMP|55335-4|LNC|little s Ab|little s Ab
C2708561|T201|COMP|55336-2|LNC|N Ab|N Ab
C2708562|T201|COMP|55337-0|LNC|P1 Ab|P1 Ab
C2708563|T201|COMP|55338-8|LNC|S little d super little a Ab|S little d super little a Ab
C2708565|T201|COMP|55339-6|LNC|S little d super little a Ab|S little d super little a Ab
C2708566|T201|COMP|55340-4|LNC|V Ab|V Ab
C2708567|T201|COMP|55341-2|LNC|X little g super little a Ab|X little g super little a Ab
C2708568|T201|COMP|55342-0|LNC|S little d super little a Ag|S little d super little a Ag
C2708570|T201|COMP|55343-8|LNC|Anidulafungin|Anidulafungin
C2708572|T201|COMP|55345-3|LNC|VIM gene methylation|VIM gene methylation
C2708574|T201|COMP|55346-1|LNC|Clobazam+Norclobazam|Clobazam+Norclobazam
C2708576|T201|COMP|55347-9|LNC|Coagulation ecarin induced|Coagulation ecarin induced
C2708578|T201|COMP|55348-7|LNC|Cortisol^20M post XXX challenge|Cortisol^20M post XXX challenge
C2708579|T201|COMP|55349-5|LNC|Ethyl glucuronide|Ethyl glucuronide
C2708580|T201|COMP|55350-3|LNC|Fenfluramine|Fenfluramine
C2708581|T201|COMP|55351-1|LNC|Glucose^1.5H post 75 g glucose PO|Glucose^1.5H post 75 g glucose PO
C2708582|T201|COMP|55352-9|LNC|Glucose^45M post 75 g glucose PO|Glucose^45M post 75 g glucose PO
C2708583|T201|COMP|55353-7|LNC|Hirudin|Hirudin
C2708584|T201|COMP|55354-5|LNC|Osmolality^post 4H FFst|Osmolality^post 4H FFst
C2708585|T201|COMP|55355-2|LNC|Osmolality^post 7H FFst|Osmolality^post 7H FFst
C2708586|T201|COMP|55356-0|LNC|Osmolality^post 5H FFst|Osmolality^post 5H FFst
C2708587|T201|COMP|55357-8|LNC|Osmolality^post 3H FFst|Osmolality^post 3H FFst
C2708588|T201|COMP|55358-6|LNC|Osmolality^post 2H FFst|Osmolality^post 2H FFst
C2708589|T201|COMP|55359-4|LNC|Osmolality^post 1H FFst|Osmolality^post 1H FFst
C2708590|T201|COMP|55360-2|LNC|Osmolality^post 6H FFst|Osmolality^post 6H FFst
C2708591|T201|COMP|55361-0|LNC|Osmolality^baseline|Osmolality^baseline
C2708593|T201|COMP|55363-6|LNC|Argatroban|Argatroban
C2708594|T201|COMP|55364-4|LNC|Cells.CD5+CD19+CD38+/100 cells|Cells.CD5+CD19+CD38+/100 cells
C2708596|T201|COMP|55365-1|LNC|Cells.CD138+Kappa+/100 cells|Cells.CD138+Kappa+/100 cells
C2708598|T201|COMP|55366-9|LNC|Cells.CD138+Lambda+/100 cells|Cells.CD138+Lambda+/100 cells
C2708600|T201|COMP|55367-7|LNC|Cholesterol crystals|Cholesterol crystals
C2708601|T201|COMP|55368-5|LNC|Crystals.amorphous|Crystals.amorphous
C2708602|T201|COMP|55369-3|LNC|Dengue virus Ab|Dengue virus Ab
C2708603|T201|COMP|55370-1|LNC|Hemoglobin A2+C+E+O/Hemoglobin.total|Hemoglobin A2+C+E+O/Hemoglobin.total
C2708605|T201|COMP|55371-9|LNC|Hemoglobin A2+E+O/Hemoglobin.total|Hemoglobin A2+E+O/Hemoglobin.total
C2708607|T201|COMP|55372-7|LNC|Hemoglobin Constant Spring/Hemoglobin.total|Hemoglobin Constant Spring/Hemoglobin.total
C2708609|T201|COMP|55373-5|LNC|Hemoglobin D+G/Hemoglobin.total|Hemoglobin D+G/Hemoglobin.total
C2708611|T201|COMP|55374-3|LNC|Hemoglobin N+I/Hemoglobin.total|Hemoglobin N+I/Hemoglobin.total
C2708613|T201|COMP|55375-0|LNC|Megaloblasts|Megaloblasts
C2708614|T201|COMP|55376-8|LNC|Megaloblasts/100 leukocytes|Megaloblasts/100 leukocytes
C2708616|T201|COMP|55377-6|LNC|Mononuclear cells.immature/100 leukocytes|Mononuclear cells.immature/100 leukocytes
C2708618|T201|COMP|55378-4|LNC|Phosphate crystals.amorphous|Phosphate crystals.amorphous
C2708619|T201|COMP|55379-2|LNC|Snowshoe hare virus Ab.IgM|Snowshoe hare virus Ab.IgM
C2708620|T201|COMP|55380-0|LNC|West Nile virus Ab|West Nile virus Ab
C2708621|T201|COMP|55381-8|LNC|Glucose^2.5H post 75 g glucose PO|Glucose^2.5H post 75 g glucose PO
C2708622|T201|COMP|55382-6|LNC|Insulin^5M post XXX challenge|Insulin^5M post XXX challenge
C2708623|T201|COMP|55383-4|LNC|Insulin^10M post XXX challenge|Insulin^10M post XXX challenge
C2708624|T201|COMP|55384-2|LNC|Insulin^3M post XXX challenge|Insulin^3M post XXX challenge
C2708625|T201|COMP|55385-9|LNC|Insulin^15M post XXX challenge|Insulin^15M post XXX challenge
C2708626|T201|COMP|55386-7|LNC|Insulin^2M post XXX challenge|Insulin^2M post XXX challenge
C2708627|T201|COMP|55387-5|LNC|Insulin^45M post XXX challenge|Insulin^45M post XXX challenge
C2708628|T201|COMP|55388-3|LNC|Insulin^4H post XXX challenge|Insulin^4H post XXX challenge
C2708629|T201|COMP|55389-1|LNC|Insulin^5H post XXX challenge|Insulin^5H post XXX challenge
C2708630|T201|COMP|55390-9|LNC|Insulin^6H post XXX challenge|Insulin^6H post XXX challenge
C2708631|T201|COMP|55391-7|LNC|Insulin^4M post XXX challenge|Insulin^4M post XXX challenge
C2708632|T201|COMP|55392-5|LNC|Insulin^1M post XXX challenge|Insulin^1M post XXX challenge
C2708633|T201|COMP|55393-3|LNC|Lead|Lead
C2708634|T201|COMP|55394-1|LNC|Protein & Glucose panel|Protein & Glucose panel
C2708635|T201|COMP|55395-8|LNC|Phospholipid Ab.IgA & IgG & IgM panel|Phospholipid Ab.IgA & IgG & IgM panel
C2708637|T201|COMP|55396-6|LNC|Beta 2 glycoprotein 1 Ab.IgA & IgG panel|Beta 2 glycoprotein 1 Ab.IgA & IgG panel
C2708639|T201|COMP|55397-4|LNC|Short myasthenia gravis panel|Short myasthenia gravis panel
C2708641|T201|COMP|55398-2|LNC|Short Fibrin D-dimer FEU & DDU panel|Short Fibrin D-dimer FEU & DDU panel
C2708647|T201|COMP|55401-4|LNC|Warfarin tracking panel|Warfarin tracking panel
C2708649|T201|COMP|55402-2|LNC|West Nile virus Ab.IgG & IgM panel|West Nile virus Ab.IgG & IgM panel
C2708680|T201|COMP|55419-6|LNC|Home drug screening panel|Home drug screening panel
C2708682|T201|COMP|55420-4|LNC|Hours after meal|Hours after meal
C2708692|T201|COMP|55428-7|LNC|Drug test kit name|Drug test kit name
C2708694|T201|COMP|55429-5|LNC|Short blood count panel|Short blood count panel
C2708697|T201|COMP|55431-1|LNC|Cells.HLA-B27|Cells.HLA-B27
C2708699|T201|COMP|55432-9|LNC|Immature cells|Immature cells
C2708701|T201|COMP|55433-7|LNC|Immature cells/100 leukocytes|Immature cells/100 leukocytes
C2708703|T201|COMP|55434-5|LNC|Insulin^20M post XXX challenge|Insulin^20M post XXX challenge
C2708704|T201|COMP|55435-2|LNC|Mononuclear cells.immature|Mononuclear cells.immature
C2708706|T201|COMP|55436-0|LNC|Myeloblasts/100 leukocytes|Myeloblasts/100 leukocytes
C2708707|T201|COMP|55437-8|LNC|Neoplastic cells/100 leukocytes|Neoplastic cells/100 leukocytes
C2708709|T201|COMP|55438-6|LNC|Dengue virus Ab|Dengue virus Ab
C2708711|T201|COMP|55581-3|LNC|sulfaSALAzine|sulfaSALAzine
C2708712|T201|COMP|55582-1|LNC|Timolol|Timolol
C2708713|T201|COMP|55583-9|LNC|Tranylcypromine|Tranylcypromine
C2708714|T201|COMP|55584-7|LNC|Trimethoprim|Trimethoprim
C2708715|T201|COMP|55585-4|LNC|Tripelennamine|Tripelennamine
C2708716|T201|COMP|55586-2|LNC|Verapamil|Verapamil
C2708717|T201|COMP|55587-0|LNC|Methamphetamine|Methamphetamine
C2708718|T201|COMP|55588-8|LNC|OXcarbazepine+10-Hydroxycarbazepine|OXcarbazepine+10-Hydroxycarbazepine
C2708736|T201|COMP|55459-2|LNC|Prekallikrein|Prekallikrein
C2708737|T201|COMP|55460-0|LNC|Protein C Ag|Protein C Ag
C2708738|T201|COMP|55461-8|LNC|Protein C|Protein C
C2708739|T201|COMP|55462-6|LNC|Thyrotropin|Thyrotropin
C2708740|T201|COMP|55463-4|LNC|Influenza virus A swine origin RNA|Influenza virus A swine origin RNA
C2708742|T201|COMP|55464-2|LNC|Influenza virus A swine origin RNA|Influenza virus A swine origin RNA
C2708743|T201|COMP|55465-9|LNC|Influenza virus A H1 2009 pandemic RNA|Influenza virus A H1 2009 pandemic RNA
C2708745|T201|COMP|55466-7|LNC|Influenza virus A H1 2009 pandemic RNA panel|Influenza virus A H1 2009 pandemic RNA panel
C2708747|T201|COMP|55467-5|LNC|11-Deoxycortisol^baseline|11-Deoxycortisol^baseline
C2708748|T201|COMP|55468-3|LNC|11-Deoxycortisol^1H post dose corticotropin|11-Deoxycortisol^1H post dose corticotropin
C2708750|T201|COMP|55470-9|LNC|17-Hydroxyprogesterone^1H post dose corticotropin|17-Hydroxyprogesterone^1H post dose corticotropin
C2708751|T201|COMP|55471-7|LNC|Aldosterone^1H post dose corticotropin|Aldosterone^1H post dose corticotropin
C2708752|T201|COMP|55472-5|LNC|Cortisol^2.5H post XXX challenge|Cortisol^2.5H post XXX challenge
C2708753|T201|COMP|55473-3|LNC|Cortisol^3H post XXX challenge|Cortisol^3H post XXX challenge
C2708754|T201|COMP|55474-1|LNC|Dehydroepiandrosterone^baseline|Dehydroepiandrosterone^baseline
C2708755|T201|COMP|55475-8|LNC|Dehydroepiandrosterone^1H post dose corticotropin|Dehydroepiandrosterone^1H post dose corticotropin
C2708756|T201|COMP|55476-6|LNC|Estradiol^baseline|Estradiol^baseline
C2708757|T201|COMP|55477-4|LNC|Estradiol^4H post XXX challenge|Estradiol^4H post XXX challenge
C2708758|T201|COMP|55478-2|LNC|Follitropin^4H post XXX challenge|Follitropin^4H post XXX challenge
C2708759|T201|COMP|55479-0|LNC|Insulin^7M post dose glucose IV|Insulin^7M post dose glucose IV
C2708760|T201|COMP|55480-8|LNC|Insulin^5M pre dose glucose|Insulin^5M pre dose glucose
C2708761|T201|COMP|55481-6|LNC|Insulin^10M pre dose glucose|Insulin^10M pre dose glucose
C2708762|T201|COMP|55482-4|LNC|Insulin^4H post dose glucose IV|Insulin^4H post dose glucose IV
C2708763|T201|COMP|55483-2|LNC|Insulin^1.5H post dose glucose IV|Insulin^1.5H post dose glucose IV
C2708764|T201|COMP|55484-0|LNC|Insulin^10M post dose glucose IV|Insulin^10M post dose glucose IV
C2708765|T201|COMP|55485-7|LNC|Insulin^1H post dose glucose IV|Insulin^1H post dose glucose IV
C2708766|T201|COMP|55486-5|LNC|Insulin^1M post dose glucose IV|Insulin^1M post dose glucose IV
C2708767|T201|COMP|55487-3|LNC|Insulin^2.5H post dose glucose IV|Insulin^2.5H post dose glucose IV
C2708768|T201|COMP|55488-1|LNC|Insulin^1H post dose glucagon|Insulin^1H post dose glucagon
C2708769|T201|COMP|55489-9|LNC|Insulin^1.5H post dose glucagon|Insulin^1.5H post dose glucagon
C2708770|T201|COMP|55490-7|LNC|Insulin^45M post dose glucagon|Insulin^45M post dose glucagon
C2708771|T201|COMP|55491-5|LNC|Insulin^2H post dose glucagon|Insulin^2H post dose glucagon
C2708772|T201|COMP|55492-3|LNC|Insulin^30M post dose glucose IV|Insulin^30M post dose glucose IV
C2708773|T201|COMP|55493-1|LNC|Insulin^3H post dose glucose IV|Insulin^3H post dose glucose IV
C2708774|T201|COMP|55494-9|LNC|Insulin^5M post dose glucose IV|Insulin^5M post dose glucose IV
C2708775|T201|COMP|55495-6|LNC|Insulin^45M post dose glucose IV|Insulin^45M post dose glucose IV
C2708776|T201|COMP|55496-4|LNC|Insulin^2H post dose glucose IV|Insulin^2H post dose glucose IV
C2708777|T201|COMP|55497-2|LNC|Insulin^3M post dose glucose IV|Insulin^3M post dose glucose IV
C2708778|T201|COMP|55498-0|LNC|Insulin^7M pre dose glucose|Insulin^7M pre dose glucose
C2708779|T201|COMP|55499-8|LNC|Insulin^15M post dose glucose IV|Insulin^15M post dose glucose IV
C2708780|T201|COMP|55500-3|LNC|Insulin^30M post dose glucagon|Insulin^30M post dose glucagon
C2708781|T201|COMP|55501-1|LNC|Lutropin^4H post XXX challenge|Lutropin^4H post XXX challenge
C2708782|T201|COMP|55502-9|LNC|Prolactin^20M post dose TRH IV|Prolactin^20M post dose TRH IV
C2708783|T201|COMP|55503-7|LNC|Prolactin^40M post dose TRH IV|Prolactin^40M post dose TRH IV
C2708784|T201|COMP|55504-5|LNC|Somatotropin^2H post dose glucagon|Somatotropin^2H post dose glucagon
C2708785|T201|COMP|55505-2|LNC|Somatotropin^30M post dose glucose|Somatotropin^30M post dose glucose
C2708786|T201|COMP|55506-0|LNC|Somatotropin^10M post exercise|Somatotropin^10M post exercise
C2708787|T201|COMP|55507-8|LNC|Somatotropin^2H post dose glucose|Somatotropin^2H post dose glucose
C2708788|T201|COMP|55508-6|LNC|Somatotropin^1H post dose glucose|Somatotropin^1H post dose glucose
C2708789|T201|COMP|55509-4|LNC|Somatotropin^45M post dose cloNIDine|Somatotropin^45M post dose cloNIDine
C2708790|T201|COMP|55510-2|LNC|Somatotropin^1.5H post dose glucose|Somatotropin^1.5H post dose glucose
C2708791|T201|COMP|55511-0|LNC|Somatotropin^3H post dose glucagon|Somatotropin^3H post dose glucagon
C2708792|T201|COMP|55512-8|LNC|Somatotropin^30M post dose glucagon|Somatotropin^30M post dose glucagon
C2708793|T201|COMP|55513-6|LNC|Somatotropin^30M post dose cloNIDine|Somatotropin^30M post dose cloNIDine
C2708794|T201|COMP|55514-4|LNC|Somatotropin^20M post exercise|Somatotropin^20M post exercise
C2708795|T201|COMP|55515-1|LNC|Somatotropin^2.5H post dose glucagon|Somatotropin^2.5H post dose glucagon
C2708796|T201|COMP|55516-9|LNC|Somatotropin^1.5H post dose glucagon|Somatotropin^1.5H post dose glucagon
C2708797|T201|COMP|55517-7|LNC|Somatotropin^1H post dose glucagon|Somatotropin^1H post dose glucagon
C2708799|T201|COMP|55519-3|LNC|Testosterone^baseline|Testosterone^baseline
C2708800|T201|COMP|55520-1|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C2708801|T201|COMP|55521-9|LNC|Acebutolol|Acebutolol
C2708802|T201|COMP|55522-7|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C2708803|T201|COMP|55523-5|LNC|Anileridine|Anileridine
C2708804|T201|COMP|55524-3|LNC|Atropine|Atropine
C2708805|T201|COMP|55525-0|LNC|Benzoylecgonine|Benzoylecgonine
C2708806|T201|COMP|55526-8|LNC|Brompheniramine|Brompheniramine
C2708807|T201|COMP|55527-6|LNC|buPROPion|buPROPion
C2708808|T201|COMP|55528-4|LNC|Chloral hydrate|Chloral hydrate
C2708809|T201|COMP|55544-1|LNC|hydrOXYzine|hydrOXYzine
C2708810|T201|COMP|55545-8|LNC|Indomethacin|Indomethacin
C2708811|T201|COMP|55546-6|LNC|Ketoprofen|Ketoprofen
C2708812|T201|COMP|55547-4|LNC|Labetalol|Labetalol
C2708813|T201|COMP|55548-2|LNC|metFORMIN|metFORMIN
C2708814|T201|COMP|55549-0|LNC|Methocarbamol|Methocarbamol
C2708815|T201|COMP|55550-8|LNC|Methsuximide+Normethsuximide|Methsuximide+Normethsuximide
C2708816|T201|COMP|55551-6|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C2708817|T201|COMP|55552-4|LNC|Methylphenidate|Methylphenidate
C2708818|T201|COMP|55553-2|LNC|Metoprolol|Metoprolol
C2708819|T201|COMP|55554-0|LNC|Mirtazapine|Mirtazapine
C2708820|T201|COMP|55555-7|LNC|Molybdenum|Molybdenum
C2708821|T201|COMP|55556-5|LNC|Nadolol|Nadolol
C2708822|T201|COMP|55557-3|LNC|Nicotine|Nicotine
C2708823|T201|COMP|55558-1|LNC|Nicotine|Nicotine
C2708824|T201|COMP|55559-9|LNC|Norpropoxyphene|Norpropoxyphene
C2708825|T201|COMP|55560-7|LNC|Orphenadrine|Orphenadrine
C2708826|T201|COMP|55561-5|LNC|Oxprenolol|Oxprenolol
C2708827|T201|COMP|55562-3|LNC|Oxyphenbutazone|Oxyphenbutazone
C2708828|T201|COMP|55563-1|LNC|Paraldehyde|Paraldehyde
C2708829|T201|COMP|55564-9|LNC|Pentazocine|Pentazocine
C2708830|T201|COMP|55565-6|LNC|Phenacetin|Phenacetin
C2708831|T201|COMP|55566-4|LNC|Phenelzine|Phenelzine
C2708832|T201|COMP|55567-2|LNC|Pheniramine|Pheniramine
C2708833|T201|COMP|55568-0|LNC|Phenolphthalein|Phenolphthalein
C2708834|T201|COMP|55569-8|LNC|Phentermine|Phentermine
C2708835|T201|COMP|55570-6|LNC|predniSONE|predniSONE
C2708836|T201|COMP|55571-4|LNC|Prilocaine|Prilocaine
C2708837|T201|COMP|55572-2|LNC|Procaine|Procaine
C2708838|T201|COMP|55573-0|LNC|Promethazine|Promethazine
C2708839|T201|COMP|55574-8|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C2708840|T201|COMP|55575-5|LNC|Pseudoephedrine|Pseudoephedrine
C2708841|T201|COMP|55576-3|LNC|QUEtiapine|QUEtiapine
C2708842|T201|COMP|55577-1|LNC|Salicylamide|Salicylamide
C2708843|T201|COMP|55578-9|LNC|Sildenafil citrate|Sildenafil citrate
C2708844|T201|COMP|55579-7|LNC|Sotalol|Sotalol
C2708845|T201|COMP|55580-5|LNC|Sulfapyridine|Sulfapyridine
C2708846|T201|COMP|55589-6|LNC|Budgerigar feather Ab.IgE|Budgerigar feather Ab.IgE
C2708847|T201|COMP|55590-4|LNC|Canary feather Ab.IgE|Canary feather Ab.IgE
C2708848|T201|COMP|55591-2|LNC|Chicken feather Ab.IgE|Chicken feather Ab.IgE
C2708849|T201|COMP|55592-0|LNC|Cockatiel feather Ab.IgE|Cockatiel feather Ab.IgE
C2708850|T201|COMP|55593-8|LNC|Creatinine|Creatinine
C2708851|T201|COMP|55594-6|LNC|Duck feather Ab.IgE|Duck feather Ab.IgE
C2708852|T201|COMP|55595-3|LNC|Finch feather Ab.IgE|Finch feather Ab.IgE
C2708853|T201|COMP|55596-1|LNC|Goose feather Ab.IgE|Goose feather Ab.IgE
C2708854|T201|COMP|55597-9|LNC|J little s super little b Ab|J little s super little b Ab
C2708855|T201|COMP|55598-7|LNC|Leukocytes.disintegrated/100 leukocytes|Leukocytes.disintegrated/100 leukocytes
C2708857|T201|COMP|55599-5|LNC|Leukocytes.disintegrated/100 leukocytes|Leukocytes.disintegrated/100 leukocytes
C2708863|T201|COMP|55605-0|LNC|Parakeet feather Ab.IgE|Parakeet feather Ab.IgE
C2708864|T201|COMP|55606-8|LNC|Parrot feather Ab.IgE|Parrot feather Ab.IgE
C2708865|T201|COMP|55607-6|LNC|Triglyceride/Cholesterol.in HDL|Triglyceride/Cholesterol.in HDL
C2708866|T201|COMP|55608-4|LNC|Turkey feather Ab.IgE|Turkey feather Ab.IgE
C2708867|T201|COMP|55609-2|LNC|Urea|Urea
C2708868|T201|COMP|55610-0|LNC|Follitropin^2nd specimen post XXX challenge|Follitropin^2nd specimen post XXX challenge
C2708869|T201|COMP|55611-8|LNC|Follitropin^1st specimen post XXX challenge|Follitropin^1st specimen post XXX challenge
C2708870|T201|COMP|55612-6|LNC|Follitropin^7th specimen post XXX challenge|Follitropin^7th specimen post XXX challenge
C2708871|T201|COMP|55628-2|LNC|Cefadroxil|Cefadroxil
C2708872|T201|COMP|55629-0|LNC|Cephaloglycin|Cephaloglycin
C2708873|T201|COMP|55630-8|LNC|Cephalothin+Sulbactam|Cephalothin+Sulbactam
C2708875|T201|COMP|55631-6|LNC|Cephalothin+Sulbactam|Cephalothin+Sulbactam
C2708876|T201|COMP|55632-4|LNC|Cephalothin+Sulbactam|Cephalothin+Sulbactam
C2708877|T201|COMP|55633-2|LNC|Cephalothin+Sulbactam|Cephalothin+Sulbactam
C2708878|T201|COMP|55634-0|LNC|Cefamandole+Sulbactam|Cefamandole+Sulbactam
C2708880|T201|COMP|55635-7|LNC|Cefamandole+Sulbactam|Cefamandole+Sulbactam
C2708881|T201|COMP|55636-5|LNC|Cefamandole+Sulbactam|Cefamandole+Sulbactam
C2708882|T201|COMP|55637-3|LNC|Cefamandole+Sulbactam|Cefamandole+Sulbactam
C2708883|T201|COMP|55638-1|LNC|Cephapirin|Cephapirin
C2708884|T201|COMP|55639-9|LNC|Cefatrizine|Cefatrizine
C2708885|T201|COMP|55640-7|LNC|Cefetamet|Cefetamet
C2708886|T201|COMP|55641-5|LNC|Cefmenoxime|Cefmenoxime
C2708887|T201|COMP|55642-3|LNC|Cefonicid|Cefonicid
C2708888|T201|COMP|55643-1|LNC|Ceforanide|Ceforanide
C2708889|T201|COMP|55644-9|LNC|Cefotaxime+Sulbactam|Cefotaxime+Sulbactam
C2708890|T201|COMP|55645-6|LNC|Cefotiam|Cefotiam
C2708891|T201|COMP|55646-4|LNC|Cephradine|Cephradine
C2708892|T201|COMP|55647-2|LNC|Cefsulodin|Cefsulodin
C2708893|T201|COMP|55648-0|LNC|cefTAZidime+Sulbactam|cefTAZidime+Sulbactam
C2708895|T201|COMP|55649-8|LNC|cefTAZidime+Sulbactam|cefTAZidime+Sulbactam
C2708896|T201|COMP|55650-6|LNC|cefTAZidime+Sulbactam|cefTAZidime+Sulbactam
C2708897|T201|COMP|55651-4|LNC|cefTAZidime+Sulbactam|cefTAZidime+Sulbactam
C2708898|T201|COMP|55652-2|LNC|Ceftiofur|Ceftiofur
C2708899|T201|COMP|55653-0|LNC|Cefuroxime.oral|Cefuroxime.oral
C2708900|T201|COMP|55654-8|LNC|Cefuroxime|Cefuroxime
C2708901|T201|COMP|55655-5|LNC|Chlortetracycline|Chlortetracycline
C2708902|T201|COMP|55656-3|LNC|Cinoxacin|Cinoxacin
C2708903|T201|COMP|55657-1|LNC|Clindamycin.high potency|Clindamycin.high potency
C2708905|T201|COMP|55658-9|LNC|Clindamycin.high potency|Clindamycin.high potency
C2708906|T201|COMP|55659-7|LNC|Clindamycin.high potency|Clindamycin.high potency
C2708907|T201|COMP|55660-5|LNC|Clindamycin.high potency|Clindamycin.high potency
C2708908|T201|COMP|55661-3|LNC|Clofazimine|Clofazimine
C2708909|T201|COMP|55662-1|LNC|Clofazimine|Clofazimine
C2708910|T201|COMP|55663-9|LNC|Clotrimazole|Clotrimazole
C2708911|T201|COMP|55664-7|LNC|Cloxacillin|Cloxacillin
C2708912|T201|COMP|55665-4|LNC|Colistimethate|Colistimethate
C2708913|T201|COMP|55666-2|LNC|Cyclacillin|Cyclacillin
C2708914|T201|COMP|55667-0|LNC|cycloSERINE|cycloSERINE
C2708915|T201|COMP|55668-8|LNC|Dicloxacillin|Dicloxacillin
C2708916|T201|COMP|55669-6|LNC|Dibekacin|Dibekacin
C2708917|T201|COMP|55670-4|LNC|Dibekacin|Dibekacin
C2708918|T201|COMP|55671-2|LNC|Dibekacin|Dibekacin
C2708919|T201|COMP|55672-0|LNC|Dibekacin|Dibekacin
C2708920|T201|COMP|55673-8|LNC|Econazole|Econazole
C2708921|T201|COMP|55674-6|LNC|Ethambutol 2.0 ug/mL|Ethambutol 2.0 ug/mL
C2708923|T201|COMP|55675-3|LNC|Flumequine|Flumequine
C2708924|T201|COMP|55676-1|LNC|Flumequine|Flumequine
C2708925|T201|COMP|55677-9|LNC|Flumequine|Flumequine
C2708926|T201|COMP|55678-7|LNC|Flumequine|Flumequine
C2708927|T201|COMP|55679-5|LNC|Framycetin|Framycetin
C2708928|T201|COMP|55680-3|LNC|Isepamicin|Isepamicin
C2708929|T201|COMP|55681-1|LNC|Isoconazole|Isoconazole
C2708930|T201|COMP|55682-9|LNC|Isoconazole|Isoconazole
C2708931|T201|COMP|55683-7|LNC|Isoconazole|Isoconazole
C2708932|T201|COMP|55684-5|LNC|Isoconazole|Isoconazole
C2708933|T201|COMP|55685-2|LNC|Isoniazid 10.0 ug/mL|Isoniazid 10.0 ug/mL
C2708935|T201|COMP|55686-0|LNC|Miconazole|Miconazole
C2708936|T201|COMP|55687-8|LNC|Miocamycin|Miocamycin
C2708937|T201|COMP|55688-6|LNC|Nitroxoline|Nitroxoline
C2708938|T201|COMP|55689-4|LNC|Nystatin|Nystatin
C2708939|T201|COMP|55690-2|LNC|Oleandomycin|Oleandomycin
C2708940|T201|COMP|55691-0|LNC|Ornidazole|Ornidazole
C2708941|T201|COMP|55692-8|LNC|Ornidazole|Ornidazole
C2708942|T201|COMP|55693-6|LNC|Ornidazole|Ornidazole
C2708943|T201|COMP|55694-4|LNC|Ornidazole|Ornidazole
C2708944|T201|COMP|55695-1|LNC|Oxolinate|Oxolinate
C2708946|T201|COMP|55696-9|LNC|Oxolinate|Oxolinate
C2708947|T201|COMP|55697-7|LNC|Oxolinate|Oxolinate
C2708948|T201|COMP|55698-5|LNC|Oxolinate|Oxolinate
C2708949|T201|COMP|55699-3|LNC|Oxytetracycline|Oxytetracycline
C2708950|T201|COMP|55700-9|LNC|Paromomycin|Paromomycin
C2708951|T201|COMP|55701-7|LNC|Paromomycin|Paromomycin
C2708952|T201|COMP|55702-5|LNC|Paromomycin|Paromomycin
C2708953|T201|COMP|55703-3|LNC|Pipemidate|Pipemidate
C2708954|T201|COMP|55704-1|LNC|Piperacillin+Sulbactam|Piperacillin+Sulbactam
C2708955|T201|COMP|55705-8|LNC|Piromidate|Piromidate
C2708957|T201|COMP|55706-6|LNC|Piromidate|Piromidate
C2708958|T201|COMP|55707-4|LNC|Piromidate|Piromidate
C2708959|T201|COMP|55708-2|LNC|Piromidate|Piromidate
C2708960|T201|COMP|55709-0|LNC|Pristinamycin|Pristinamycin
C2708961|T201|COMP|55710-8|LNC|Pyrazinamide|Pyrazinamide
C2708962|T201|COMP|55711-6|LNC|Pyrazinamide 200.0 ug/mL|Pyrazinamide 200.0 ug/mL
C2708964|T201|COMP|55712-4|LNC|rifAMPin 40.0 ug/mL|rifAMPin 40.0 ug/mL
C2708966|T201|COMP|55713-2|LNC|Rosoxacin|Rosoxacin
C2708967|T201|COMP|55714-0|LNC|Sisomicin|Sisomicin
C2708968|T201|COMP|55715-7|LNC|Spiramycin|Spiramycin
C2708969|T201|COMP|55716-5|LNC|Ticarcillin+Sulbactam|Ticarcillin+Sulbactam
C2708971|T201|COMP|55717-3|LNC|Ticarcillin+Sulbactam|Ticarcillin+Sulbactam
C2708972|T201|COMP|55718-1|LNC|Ticarcillin+Sulbactam|Ticarcillin+Sulbactam
C2708973|T201|COMP|55719-9|LNC|Ticarcillin+Sulbactam|Ticarcillin+Sulbactam
C2708974|T201|COMP|55720-7|LNC|Tinidazole|Tinidazole
C2708975|T201|COMP|55721-5|LNC|Tinidazole|Tinidazole
C2708976|T201|COMP|55722-3|LNC|Tinidazole|Tinidazole
C2708977|T201|COMP|55723-1|LNC|Virginiamycin|Virginiamycin
C2708978|T201|COMP|55724-9|LNC|Apolipoprotein A-I & A-II & B & C panel|Apolipoprotein A-I & A-II & B & C panel
C2708982|T201|COMP|55726-4|LNC|Borrelia burgdorferi Ab.IgA & IgG & IgM panel|Borrelia burgdorferi Ab.IgA & IgG & IgM panel
C2708984|T201|COMP|55727-2|LNC|Tissue transglutaminase Ab.IgA & IgG panel|Tissue transglutaminase Ab.IgA & IgG panel
C2708986|T201|COMP|55728-0|LNC|Yersinia sp Ab.IgG & IgM panel|Yersinia sp Ab.IgG & IgM panel
C2708988|T201|COMP|55729-8|LNC|Erythrocytes.fetal/100 erythrocytes|Erythrocytes.fetal/100 erythrocytes
C2708990|T201|COMP|55730-6|LNC|Fetal blood|Fetal blood
C2708991|T201|COMP|55731-4|LNC|Inject Rh immune globulin|Inject Rh immune globulin
C2708992|T201|COMP|55737-1|LNC|Cefotiam hexetil|Cefotiam hexetil
C2708993|T201|COMP|55738-9|LNC|Cefotiam hexetil|Cefotiam hexetil
C2708994|T201|COMP|55739-7|LNC|Cefotiam hexetil|Cefotiam hexetil
C2708995|T201|COMP|55740-5|LNC|Cefotiam hexetil|Cefotiam hexetil
C2709273|T201|COMP|19594-1|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C2713036|T201|COMP|14111-9|LNC|Lymphocytes.CD23/100 lymphocytes|Lymphocytes.CD23/100 lymphocytes
C2713037|T201|COMP|2010-7|LNC|Cancer Ag 19-9|Cancer Ag 19-9
C2713038|T201|COMP|2566-8|LNC|Fatty acids.nonesterified|Fatty acids.nonesterified
C2713039|T201|COMP|2782-1|LNC|Phosphate|Phosphate
C2713040|T201|COMP|5937-8|LNC|Cocaine|Cocaine
C2713041|T201|COMP|5935-2|LNC|Benzoylecgonine|Benzoylecgonine
C2713042|T201|COMP|26922-5|LNC|Cells.CD4+CD45RA+/100 cells|Cells.CD4+CD45RA+/100 cells
C2713043|T201|COMP|6028-5|LNC|Aureobasidium pullulans Ab.IgE|Aureobasidium pullulans Ab.IgE
C2713053|T201|COMP|18433-3|LNC|1,3-Dichlorobenzene|1,3-Dichlorobenzene
C2713054|T201|COMP|1672-5|LNC|17-Ketogenic steroids|17-Ketogenic steroids
C2713055|T201|COMP|6828-8|LNC|Alternaria alternata Ab.IgE|Alternaria alternata Ab.IgE
C2713056|T201|COMP|15531-7|LNC|Alternaria alternata Ab.IgE.RAST class|Alternaria alternata Ab.IgE.RAST class
C2713058|T201|COMP|25307-0|LNC|Alternaria alternata Ab.IgG.RAST class|Alternaria alternata Ab.IgG.RAST class
C2713059|T201|COMP|25497-9|LNC|Acarus siro Ab.IgE.RAST class|Acarus siro Ab.IgE.RAST class
C2713060|T201|COMP|21040-1|LNC|Alpha ketoglutarate/Creatinine|Alpha ketoglutarate/Creatinine
C2713061|T201|COMP|24090-3|LNC|Alpha-N-acetylglucosaminidase|Alpha-N-acetylglucosaminidase
C2713062|T201|COMP|20422-2|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C2713063|T201|COMP|26883-9|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C2713064|T201|COMP|16358-4|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C2713065|T201|COMP|16357-6|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C2713066|T201|COMP|16356-8|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C2713067|T201|COMP|16354-3|LNC|Amino beta guanidinopropionate|Amino beta guanidinopropionate
C2713068|T201|COMP|28611-2|LNC|Amino beta guanidinopropionate/Creatinine|Amino beta guanidinopropionate/Creatinine
C2713069|T201|COMP|16336-0|LNC|Alkaline phosphatase.placental|Alkaline phosphatase.placental
C2713070|T201|COMP|6769-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C2713071|T201|COMP|11567-5|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C2713076|T201|COMP|17223-9|LNC|Cells.CD14/100 cells|Cells.CD14/100 cells
C2713077|T201|COMP|31121-7|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C2713079|T201|COMP|7352-8|LNC|Agrostis stolonifera Ab.IgE|Agrostis stolonifera Ab.IgE
C2713081|T201|COMP|11036-1|LNC|Aldolase|Aldolase
C2713085|T201|COMP|7561-4|LNC|Amaranthus palmeri Ab.IgE|Amaranthus palmeri Ab.IgE
C2713089|T201|COMP|33298-1|LNC|Amdinocillin|Amdinocillin
C2713090|T201|COMP|7730-5|LNC|Platanus occidentalis Ab.IgE|Platanus occidentalis Ab.IgE
C2713091|T201|COMP|14602-7|LNC|Amoxapine+8-Hydroxyamoxapine|Amoxapine+8-Hydroxyamoxapine
C2713092|T201|COMP|6697-7|LNC|Amylase|Amylase
C2713098|T201|COMP|9319-5|LNC|Androstenedione|Androstenedione
C2713099|T201|COMP|19060-3|LNC|Antibodies identified|Antibodies identified
C2713100|T201|COMP|6843-7|LNC|Apis mellifera Ab.IgE|Apis mellifera Ab.IgE
C2713101|T201|COMP|6772-8|LNC|Apolipoprotein B|Apolipoprotein B
C2713102|T201|COMP|6685-2|LNC|Apolipoprotein B/Apolipoprotein A-I|Apolipoprotein B/Apolipoprotein A-I
C2713103|T201|COMP|15116-7|LNC|Arsenic|Arsenic
C2713104|T201|COMP|16004-4|LNC|Artemisia tridentata Ab.IgE.RAST class|Artemisia tridentata Ab.IgE.RAST class
C2713113|T201|COMP|16573-8|LNC|Cerebroside sulfatase|Cerebroside sulfatase
C2713114|T201|COMP|6686-0|LNC|Ascorbate|Ascorbate
C2713115|T201|COMP|22677-9|LNC|Aspartate|Aspartate
C2713116|T201|COMP|21083-1|LNC|Populus tremula Ab.IgE.RAST class|Populus tremula Ab.IgE.RAST class
C2713117|T201|COMP|16010-1|LNC|Atriplex lentiformis Ab.IgE.RAST class|Atriplex lentiformis Ab.IgE.RAST class
C2713118|T201|COMP|7457-5|LNC|Atriplex lentiformis Ab.IgE|Atriplex lentiformis Ab.IgE
C2713119|T201|COMP|21427-0|LNC|Avena sativa Ab.IgE.RAST class|Avena sativa Ab.IgE.RAST class
C2713120|T201|COMP|7541-6|LNC|Avena sativa Ab.IgE|Avena sativa Ab.IgE
C2713121|T201|COMP|22835-3|LNC|Avian pneumovirus Ab|Avian pneumovirus Ab
C2713122|T201|COMP|13504-6|LNC|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C2713123|T201|COMP|27983-6|LNC|Borrelia burgdorferi 41kD Ab|Borrelia burgdorferi 41kD Ab
C2713124|T201|COMP|22957-5|LNC|Burkholderia mallei Ab|Burkholderia mallei Ab
C2713125|T201|COMP|26579-3|LNC|Beta aminoisobutyrate/Creatinine|Beta aminoisobutyrate/Creatinine
C2713126|T201|COMP|2928-0|LNC|Beta fructofuranosidase|Beta fructofuranosidase
C2713127|T201|COMP|14150-7|LNC|Beta glucuronidase|Beta glucuronidase
C2713128|T201|COMP|1948-9|LNC|Beta hydroxybutyrate dehydrogenase|Beta hydroxybutyrate dehydrogenase
C2713129|T201|COMP|17423-5|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C2713130|T201|COMP|6255-4|LNC|Lepidoglyphus destructor Ab.IgE|Lepidoglyphus destructor Ab.IgE
C2713131|T201|COMP|24157-0|LNC|Quercus virginiana Ab.IgE|Quercus virginiana Ab.IgE
C2713132|T201|COMP|7363-5|LNC|Festuca elatior Ab.IgE|Festuca elatior Ab.IgE
C2713133|T201|COMP|30988-0|LNC|Panicum milliaceum Ab.IgE|Panicum milliaceum Ab.IgE
C2713134|T201|COMP|19735-0|LNC|Dactylis glomerata Ab.IgE|Dactylis glomerata Ab.IgE
C2713135|T201|COMP|7582-0|LNC|Carya illinoinensis nut Ab.IgE|Carya illinoinensis nut Ab.IgE
C2713136|T201|COMP|21477-5|LNC|Solanum tuberosum Ab.IgE|Solanum tuberosum Ab.IgE
C2713137|T201|COMP|15282-7|LNC|Secale cereale pollen Ab.IgE|Secale cereale pollen Ab.IgE
C2713139|T201|COMP|6283-6|LNC|Elymus triticoides Ab.IgE|Elymus triticoides Ab.IgE
C2713140|T201|COMP|1009-0|LNC|Direct antiglobulin test.poly specific reagent|Direct antiglobulin test.poly specific reagent
C2713141|T201|COMP|1405-0|LNC|Cortisol^1H post dose U/kg insulin IV|Cortisol^1H post dose U/kg insulin IV
C2713142|T201|COMP|1420-9|LNC|Cortisol^30M post dose U/kg insulin IV|Cortisol^30M post dose U/kg insulin IV
C2713143|T201|COMP|1511-5|LNC|Glucose^1H post dose U/kg insulin IV|Glucose^1H post dose U/kg insulin IV
C2713144|T201|COMP|1529-7|LNC|Glucose^30M post dose U/kg insulin IV|Glucose^30M post dose U/kg insulin IV
C2713145|T201|COMP|23941-8|LNC|Xylose^2H post 25 g xylose PO|Xylose^2H post 25 g xylose PO
C2713146|T201|COMP|2088-3|LNC|Cholesterol.in IDL|Cholesterol.in IDL
C2713147|T201|COMP|2090-9|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C2713148|T201|COMP|2565-0|LNC|Cholesterol|Cholesterol
C2713149|T201|COMP|2803-5|LNC|Phytanate|Phytanate
C2713150|T201|COMP|16744-5|LNC|Nordiazepam|Nordiazepam
C2713151|T201|COMP|4033-7|LNC|Spironolactone|Spironolactone
C2713152|T201|COMP|17345-0|LNC|Neutrophil Ab|Neutrophil Ab
C2713153|T201|COMP|3733-3|LNC|Lysergate diethylamide|Lysergate diethylamide
C2713154|T201|COMP|7666-1|LNC|Rhodotorula spp Ab.IgE|Rhodotorula spp Ab.IgE
C2713155|T201|COMP|15277-7|LNC|Turkey feather Ab.IgE|Turkey feather Ab.IgE
C2713156|T201|COMP|16540-7|LNC|Cannabinoids|Cannabinoids
C2713157|T201|COMP|13222-5|LNC|Chlamydia trachomatis C Ab|Chlamydia trachomatis C Ab
C2713158|T201|COMP|17613-1|LNC|Streptococcus pneumoniae 1 Ab^2nd specimen|Streptococcus pneumoniae 1 Ab^2nd specimen
C2713159|T201|COMP|13163-1|LNC|Streptococcus pneumoniae 12 Ab|Streptococcus pneumoniae 12 Ab
C2713161|T201|COMP|20653-2|LNC|Phenylalanine|Phenylalanine
C2713162|T201|COMP|15830-3|LNC|Zea mays Ab.IgE.RAST class|Zea mays Ab.IgE.RAST class
C2713163|T201|COMP|22852-8|LNC|Babesia caballi Ab|Babesia caballi Ab
C2713164|T201|COMP|21318-1|LNC|Baccharis spp Ab.IgE.RAST class|Baccharis spp Ab.IgE.RAST class
C2713165|T201|COMP|21317-3|LNC|Baccharis spp Ab.IgE|Baccharis spp Ab.IgE
C2713166|T201|COMP|14476-6|LNC|Microorganism identified|Microorganism identified
C2713167|T201|COMP|3373-8|LNC|Barbiturate screen absent|Barbiturate screen absent
C2713168|T201|COMP|27376-3|LNC|C peptide|C peptide
C2713169|T201|COMP|35195-7|LNC|C peptide|C peptide
C2713170|T201|COMP|22165-5|LNC|Caprine arthritis encephalitis virus Ab|Caprine arthritis encephalitis virus Ab
C2713171|T201|COMP|20743-1|LNC|Caprine arthritis encephalitis virus Ab|Caprine arthritis encephalitis virus Ab
C2713172|T201|COMP|9499-5|LNC|Candida sp Ab.IgG|Candida sp Ab.IgG
C2713173|T201|COMP|20744-9|LNC|Caprine arthritis encephalitis virus Ab|Caprine arthritis encephalitis virus Ab
C2713174|T201|COMP|22985-6|LNC|Capripox virus Ab|Capripox virus Ab
C2713175|T201|COMP|9697-4|LNC|carBAMazepine 10,11-Epoxide|carBAMazepine 10,11-Epoxide
C2713176|T201|COMP|9370-8|LNC|Carbon tetrachloride|Carbon tetrachloride
C2713177|T201|COMP|7581-2|LNC|Carya illinoinensis nut basophil bound Ab|Carya illinoinensis nut basophil bound Ab
C2713178|T201|COMP|15920-2|LNC|Carya illinoinensis tree Ab.IgE.RAST class|Carya illinoinensis tree Ab.IgE.RAST class
C2713179|T201|COMP|7406-2|LNC|Carya illinoinensis tree Ab.IgE|Carya illinoinensis tree Ab.IgE
C2713180|T201|COMP|15631-5|LNC|Castanea sativa Ab.IgE.RAST class|Castanea sativa Ab.IgE.RAST class
C2713181|T201|COMP|7219-9|LNC|Castanea sativa Ab.IgE|Castanea sativa Ab.IgE
C2713182|T201|COMP|10532-0|LNC|Noramiodarone|Noramiodarone
C2713183|T201|COMP|25380-7|LNC|Dactylis glomerata Ab.IgE.RAST class|Dactylis glomerata Ab.IgE.RAST class
C2713184|T201|COMP|15056-5|LNC|Deoxypyridinoline|Deoxypyridinoline
C2713190|T201|COMP|7300-7|LNC|Ulmus americana Ab.IgE|Ulmus americana Ab.IgE
C2713191|T201|COMP|7303-1|LNC|Ulmus pumila Ab.IgE|Ulmus pumila Ab.IgE
C2713192|T201|COMP|14395-8|LNC|Urea nitrogen|Urea nitrogen
C2713193|T201|COMP|23556-4|LNC|Vesicular stomatitis virus Ab|Vesicular stomatitis virus Ab
C2713194|T201|COMP|22622-5|LNC|Xylose^1H post 25 g xylose PO|Xylose^1H post 25 g xylose PO
C2713195|T201|COMP|23944-2|LNC|Xylose^1H post 25 g xylose PO|Xylose^1H post 25 g xylose PO
C2713196|T201|COMP|22623-3|LNC|Xylose^2H post 25 g xylose PO|Xylose^2H post 25 g xylose PO
C2713197|T201|COMP|11563-4|LNC|DNA double strand Ab|DNA double strand Ab
C2713198|T201|COMP|9337-7|LNC|IgA subclass 1/IgA.total|IgA subclass 1/IgA.total
C2713202|T201|COMP|13049-2|LNC|von Willebrand factor Ag|von Willebrand factor Ag
C2713203|T201|COMP|6716-5|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C2713203|T201|COMP|8064-8|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C2713204|T201|COMP|8066-3|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C2713204|T201|COMP|6717-3|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C2713205|T201|COMP|15919-4|LNC|Carya illinoinensis nut Ab.IgE.RAST class|Carya illinoinensis nut Ab.IgE.RAST class
C2713206|T201|COMP|14110-1|LNC|Lymphocytes.CD22/100 lymphocytes|Lymphocytes.CD22/100 lymphocytes
C2713207|T201|COMP|13224-1|LNC|Chlamydia trachomatis G+F+K Ab|Chlamydia trachomatis G+F+K Ab
C2713208|T201|COMP|13223-3|LNC|Chlamydia trachomatis B Ab|Chlamydia trachomatis B Ab
C2713211|T201|COMP|25814-5|LNC|Lathyrus sativus Ab.IgE|Lathyrus sativus Ab.IgE
C2713212|T201|COMP|16143-0|LNC|Butane|Butane
C2713213|T201|COMP|13849-5|LNC|Lymphocytes.CD3+CD26+/100 lymphocytes|Lymphocytes.CD3+CD26+/100 lymphocytes
C2713214|T201|COMP|41111-6|LNC|COL5A1 gene targeted mutation analysis|COL5A1 gene targeted mutation analysis
C2713215|T201|COMP|5940-2|LNC|Cocaine|Cocaine
C2713216|T201|COMP|5941-0|LNC|Cocaine|Cocaine
C2713217|T201|COMP|14289-3|LNC|Coproporphyrin|Coproporphyrin
C2713218|T201|COMP|17694-1|LNC|Coproporphyrin|Coproporphyrin
C2713219|T201|COMP|2146-9|LNC|Cortisol.free|Cortisol.free
C2713220|T201|COMP|19426-6|LNC|Dextromethamphetamine|Dextromethamphetamine
C2713221|T201|COMP|32380-8|LNC|Dicloxacillin|Dicloxacillin
C2713222|T201|COMP|21244-9|LNC|Diethylpropion|Diethylpropion
C2713223|T201|COMP|7306-4|LNC|Epicoccum purpurascens Ab.IgE|Epicoccum purpurascens Ab.IgE
C2713230|T201|COMP|25504-2|LNC|Pinus radiata Ab.IgE.RAST class|Pinus radiata Ab.IgE.RAST class
C2713231|T201|COMP|5707-5|LNC|Opiates|Opiates
C2713232|T201|COMP|16079-6|LNC|Juglans california pollen Ab.IgE.RAST class|Juglans california pollen Ab.IgE.RAST class
C2713235|T201|COMP|3375-3|LNC|Barbiturate screen present|Barbiturate screen present
C2713236|T201|COMP|27274-0|LNC|Benzfetamine|Benzfetamine
C2713242|T201|COMP|19046-2|LNC|Bovine serum albumin Ab.IgE.RAST class|Bovine serum albumin Ab.IgE.RAST class
C2713243|T201|COMP|20480-0|LNC|Benzoylecgonine|Benzoylecgonine
C2713245|T201|COMP|6036-8|LNC|Hordeum vulgare Ab.IgE|Hordeum vulgare Ab.IgE
C2713246|T201|COMP|3386-0|LNC|Benzodiazepines negative|Benzodiazepines negative
C2713247|T201|COMP|3388-6|LNC|Benzodiazepines positive|Benzodiazepines positive
C2713248|T201|COMP|7620-8|LNC|Populus nigra Ab.IgE|Populus nigra Ab.IgE
C2713249|T201|COMP|6079-8|LNC|Blatella germanica Ab.IgE|Blatella germanica Ab.IgE
C2713250|T201|COMP|5939-4|LNC|Benzoylecgonine|Benzoylecgonine
C2713251|T201|COMP|14342-0|LNC|Catecholamines/Creatinine|Catecholamines/Creatinine
C2713252|T201|COMP|21149-0|LNC|Cefaclor Ab.IgE|Cefaclor Ab.IgE
C2713253|T201|COMP|3442-1|LNC|ceFAZolin|ceFAZolin
C2713254|T201|COMP|4158-2|LNC|ceFAZolin|ceFAZolin
C2713255|T201|COMP|6646-5|LNC|Cefepime|Cefepime
C2713256|T201|COMP|6648-1|LNC|Cefpirome|Cefpirome
C2713257|T201|COMP|6647-3|LNC|Cefpirome|Cefpirome
C2713258|T201|COMP|9503-4|LNC|Chloral hydrate|Chloral hydrate
C2713259|T201|COMP|9504-2|LNC|Chloral hydrate|Chloral hydrate
C2713260|T201|COMP|5928-1|LNC|Chloride|Chloride
C2713261|T201|COMP|2086-7|LNC|Cholesterol.in HDL|Cholesterol.in HDL
C2713262|T201|COMP|24164-6|LNC|Citrus reticulata Ab.IgE|Citrus reticulata Ab.IgE
C2713263|T201|COMP|33284-1|LNC|Clinafloxacin|Clinafloxacin
C2713264|T201|COMP|4209-3|LNC|clomiPRAMINE|clomiPRAMINE
C2713265|T201|COMP|32607-4|LNC|Clorazepate|Clorazepate
C2713266|T201|COMP|5897-3|LNC|Coagulation dilute Russell viper venom induced|Coagulation dilute Russell viper venom induced
C2713267|T201|COMP|16790-8|LNC|Doxepin+Desmethyldoxepin|Doxepin+Desmethyldoxepin
C2713268|T201|COMP|10537-9|LNC|Doxepin+Nordoxepin|Doxepin+Nordoxepin
C2713269|T201|COMP|13460-1|LNC|Cholesterol.in LDL/Cholesterol.in HDL|Cholesterol.in LDL/Cholesterol.in HDL
C2713270|T201|COMP|2092-5|LNC|Cholesterol.in VLDL|Cholesterol.in VLDL
C2713271|T201|COMP|7390-8|LNC|Corylus avellana Ab.IgE|Corylus avellana Ab.IgE
C2713272|T201|COMP|23847-7|LNC|Cotton fibers Ab.IgE|Cotton fibers Ab.IgE
C2713273|T201|COMP|14400-6|LNC|Creatinine|Creatinine
C2713274|T201|COMP|15867-5|LNC|Cucumis melo spp Ab.IgE.RAST class|Cucumis melo spp Ab.IgE.RAST class
C2713275|T201|COMP|15842-8|LNC|Cucumis melo spp Ab.IgE.RAST class|Cucumis melo spp Ab.IgE.RAST class
C2713276|T201|COMP|24161-2|LNC|Cucumis melo spp Ab.IgE|Cucumis melo spp Ab.IgE
C2713278|T201|COMP|7490-6|LNC|Cucumis melo spp Ab.IgG|Cucumis melo spp Ab.IgG
C2713280|T201|COMP|6104-4|LNC|Echinococcus sp Ab.IgE|Echinococcus sp Ab.IgE
C2713281|T201|COMP|13350-4|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C2713283|T201|COMP|30393-3|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C2713290|T201|COMP|9698-2|LNC|Desmethylclomipramine|Desmethylclomipramine
C2713291|T201|COMP|23312-2|LNC|Nairobi sheep disease virus Ab|Nairobi sheep disease virus Ab
C2713292|T201|COMP|689-0|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C2713293|T201|COMP|22433-7|LNC|Neospora caninum Ab|Neospora caninum Ab
C2713295|T201|COMP|21392-6|LNC|Panicum milliaceum Ab.IgE.RAST class|Panicum milliaceum Ab.IgE.RAST class
C2713296|T201|COMP|22762-9|LNC|Streptococcus pneumoniae 12 Ab.IgG|Streptococcus pneumoniae 12 Ab.IgG
C2713297|T201|COMP|8044-0|LNC|Trypanosoma brucei Ab|Trypanosoma brucei Ab
C2713298|T201|COMP|23516-8|LNC|Trypanosoma equiperdum Ab|Trypanosoma equiperdum Ab
C2718099|T201|COMP|4312-5|LNC|Mesantoin|Mesantoin
C2718100|T201|COMP|17268-4|LNC|Methsuximide+Desmethylmethsuximide|Methsuximide+Desmethylmethsuximide
C2718101|T201|COMP|11554-3|LNC|Magnesium|Magnesium
C2718104|T201|COMP|17298-1|LNC|Mycobacterium tuberculosis rRNA|Mycobacterium tuberculosis rRNA
C2718105|T201|COMP|20820-7|LNC|Escherichia coli K99|Escherichia coli K99
C2718106|T201|COMP|13885-9|LNC|Estrogen/Creatinine|Estrogen/Creatinine
C2718107|T201|COMP|22667-0|LNC|Fatty acids.nonesterified|Fatty acids.nonesterified
C2718108|T201|COMP|26025-7|LNC|Festuca elatior Ab.IgE.RAST class|Festuca elatior Ab.IgE.RAST class
C2718109|T201|COMP|3258-1|LNC|Fibrinogen Ag|Fibrinogen Ag
C2718110|T201|COMP|25347-6|LNC|Filaria Ab.IgG|Filaria Ab.IgG
C2718111|T201|COMP|10538-7|LNC|Fluoxetine+Norfluoxetine|Fluoxetine+Norfluoxetine
C2718112|T201|COMP|7329-6|LNC|Fusarium oxysporum Ab.IgE|Fusarium oxysporum Ab.IgE
C2718124|T201|COMP|16884-9|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C2718125|T201|COMP|16886-4|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C2718126|T201|COMP|16885-6|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C2718127|T201|COMP|16883-1|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C2718129|T201|COMP|28065-1|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C2718130|T201|COMP|12216-8|LNC|Gastrin|Gastrin
C2718131|T201|COMP|6777-7|LNC|Glucose|Glucose
C2718132|T201|COMP|22669-6|LNC|Glutamate|Glutamate
C2718133|T201|COMP|21325-6|LNC|Helminthosporium sp Ab.IgE.RAST class|Helminthosporium sp Ab.IgE.RAST class
C2718134|T201|COMP|4620-1|LNC|Hemoglobin S|Hemoglobin S
C2718135|T201|COMP|4642-5|LNC|Hemopexin|Hemopexin
C2718136|T201|COMP|13125-0|LNC|Hepatitis C virus c33c Ab|Hepatitis C virus c33c Ab
C2718137|T201|COMP|22336-2|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C2718138|T201|COMP|6423-8|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C2718139|T201|COMP|5214-2|LNC|Heterophile Ab|Heterophile Ab
C2718140|T201|COMP|17361-7|LNC|Hexane|Hexane
C2718141|T201|COMP|22673-8|LNC|Homocystine|Homocystine
C2718142|T201|COMP|6146-5|LNC|House dust Ab.IgE|House dust Ab.IgE
C2718143|T201|COMP|4277-0|LNC|HYDROmorphone|HYDROmorphone
C2718144|T201|COMP|20531-0|LNC|Hydroxyalprazolam|Hydroxyalprazolam
C2718145|T201|COMP|25935-8|LNC|Hydroxyproline/Creatinine|Hydroxyproline/Creatinine
C2718146|T201|COMP|11049-4|LNC|Hydroxyproline|Hydroxyproline
C2718147|T201|COMP|6710-8|LNC|Hydroxyproline|Hydroxyproline
C2718148|T201|COMP|20534-4|LNC|Hydroxytriazolam|Hydroxytriazolam
C2718149|T201|COMP|7165-4|LNC|Hymenoclea salsola Ab.IgE|Hymenoclea salsola Ab.IgE
C2718150|T201|COMP|13630-9|LNC|Immune complex|Immune complex
C2718151|T201|COMP|17023-3|LNC|Interleukin 7|Interleukin 7
C2718154|T201|COMP|12392-7|LNC|Itraconazole|Itraconazole
C2718155|T201|COMP|31447-6|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C2718156|T201|COMP|12393-5|LNC|Ketoconazole|Ketoconazole
C2718157|T201|COMP|25713-9|LNC|Linum usitatissimum Ab.IgE.RAST class|Linum usitatissimum Ab.IgE.RAST class
C2718158|T201|COMP|19745-9|LNC|Linum usitatissimum Ab.IgE|Linum usitatissimum Ab.IgE
C2718159|T201|COMP|17077-9|LNC|Lindane|Lindane
C2718160|T201|COMP|21549-1|LNC|Liquidambar styraciflua Ab.IgE.RAST class|Liquidambar styraciflua Ab.IgE.RAST class
C2718163|T201|COMP|7373-4|LNC|Lolium perenne Ab.IgG|Lolium perenne Ab.IgG
C2718165|T201|COMP|3736-6|LNC|Maprotiline|Maprotiline
C2718166|T201|COMP|17245-2|LNC|Meclizine|Meclizine
C2718167|T201|COMP|3751-5|LNC|Mephobarbital|Mephobarbital
C2718168|T201|COMP|22757-9|LNC|Metanephrine|Metanephrine
C2718170|T201|COMP|6798-3|LNC|Metanephrines|Metanephrines
C2718171|T201|COMP|9373-2|LNC|Methanol|Methanol
C2718172|T201|COMP|13647-3|LNC|Methylene chloride|Methylene chloride
C2718173|T201|COMP|27215-3|LNC|Mitochondria M2 Ab.IgG|Mitochondria M2 Ab.IgG
C2718174|T201|COMP|8206-5|LNC|Molybdenum|Molybdenum
C2718175|T201|COMP|9739-4|LNC|Morphine|Morphine
C2718177|T201|COMP|3835-6|LNC|N-ethylnicotinamide|N-ethylnicotinamide
C2718178|T201|COMP|4340-6|LNC|N-ethylnicotinamide|N-ethylnicotinamide
C2718179|T201|COMP|32382-4|LNC|Nitroxoline|Nitroxoline
C2718180|T201|COMP|12373-7|LNC|Norchlordiazepoxide|Norchlordiazepoxide
C2718181|T201|COMP|12376-0|LNC|Norclozapine|Norclozapine
C2718183|T201|COMP|16743-7|LNC|Nordiazepam|Nordiazepam
C2718184|T201|COMP|4354-7|LNC|Nordiazepam|Nordiazepam
C2718185|T201|COMP|4355-4|LNC|Nordoxepin|Nordoxepin
C2718186|T201|COMP|25724-6|LNC|Norsertraline|Norsertraline
C2718187|T201|COMP|20481-8|LNC|Opiates|Opiates
C2718188|T201|COMP|23323-9|LNC|Ovine herpesvirus 2 Ab|Ovine herpesvirus 2 Ab
C2718189|T201|COMP|23331-2|LNC|Ovine progressive pneumonia virus Ab|Ovine progressive pneumonia virus Ab
C2718190|T201|COMP|5712-5|LNC|Pentachlorophenol|Pentachlorophenol
C2718192|T201|COMP|12409-9|LNC|Pentoxyfylline|Pentoxyfylline
C2718193|T201|COMP|23353-6|LNC|Peste des petits ruminants virus Ab|Peste des petits ruminants virus Ab
C2718194|T201|COMP|4400-8|LNC|Phenytoin|Phenytoin
C2718195|T201|COMP|2781-3|LNC|Phosphate|Phosphate
C2718196|T201|COMP|14880-9|LNC|Phosphate|Phosphate
C2718197|T201|COMP|2801-9|LNC|Phospholipid|Phospholipid
C2718198|T201|COMP|24166-1|LNC|Pinus radiata Ab.IgE|Pinus radiata Ab.IgE
C2718199|T201|COMP|7607-5|LNC|Pinus strobus Ab.IgE|Pinus strobus Ab.IgE
C2718200|T201|COMP|32711-4|LNC|Platelet mean volume|Platelet mean volume
C2718201|T201|COMP|16081-2|LNC|Polistes spp Ab.IgE.RAST class|Polistes spp Ab.IgE.RAST class
C2718202|T201|COMP|11205-2|LNC|Polistes spp Ab.IgE|Polistes spp Ab.IgE
C2718203|T201|COMP|7256-1|LNC|Populus fremontii Ab.IgE|Populus fremontii Ab.IgE
C2718208|T201|COMP|23375-9|LNC|Porcine respiratory coronavirus Ab|Porcine respiratory coronavirus Ab
C2718209|T201|COMP|5927-9|LNC|Potassium|Potassium
C2718211|T201|COMP|1616-2|LNC|Prolactin^30M post dose U/kg insulin IV|Prolactin^30M post dose U/kg insulin IV
C2718212|T201|COMP|30463-4|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C2718213|T201|COMP|13598-8|LNC|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C2718214|T201|COMP|3544-4|LNC|Propoxyphene|Propoxyphene
C2718215|T201|COMP|22065-7|LNC|Propoxyphene|Propoxyphene
C2718217|T201|COMP|23928-5|LNC|Protoporphyrin|Protoporphyrin
C2718218|T201|COMP|19689-9|LNC|Psilocybin|Psilocybin
C2718219|T201|COMP|15884-0|LNC|Quercus alba Ab.IgE.RAST class|Quercus alba Ab.IgE.RAST class
C2718220|T201|COMP|6849-4|LNC|Quercus alba Ab.IgE|Quercus alba Ab.IgE
C2718221|T201|COMP|15883-2|LNC|Quercus virginiana Ab.IgE.RAST class|Quercus virginiana Ab.IgE.RAST class
C2718222|T201|COMP|23395-7|LNC|Reticuloendotheliosis virus Ab|Reticuloendotheliosis virus Ab
C2718223|T201|COMP|23394-0|LNC|Reticuloendotheliosis virus Ab|Reticuloendotheliosis virus Ab
C2718224|T201|COMP|16386-5|LNC|Rifabutin|Rifabutin
C2718225|T201|COMP|17615-6|LNC|Streptococcus pneumoniae 12f Ab^1st specimen|Streptococcus pneumoniae 12f Ab^1st specimen
C2718226|T201|COMP|13165-6|LNC|Streptococcus pneumoniae 19 Ab|Streptococcus pneumoniae 19 Ab
C2718227|T201|COMP|26939-9|LNC|Streptococcus pneumoniae 19 Ab|Streptococcus pneumoniae 19 Ab
C2718228|T201|COMP|17623-0|LNC|Streptococcus pneumoniae 19f Ab^2nd specimen|Streptococcus pneumoniae 19f Ab^2nd specimen
C2718229|T201|COMP|29513-9|LNC|Cysticercus Ab|Cysticercus Ab
C2718230|T201|COMP|10550-2|LNC|Temazepam|Temazepam
C2718231|T201|COMP|2993-4|LNC|Testosterone|Testosterone
C2718232|T201|COMP|13017-9|LNC|Perchloroethylene|Perchloroethylene
C2718233|T201|COMP|15648-9|LNC|Theobroma cacao Ab.IgE.RAST class|Theobroma cacao Ab.IgE.RAST class
C2718234|T201|COMP|11162-5|LNC|Theobroma cacao Ab.IgE|Theobroma cacao Ab.IgE
C2718235|T201|COMP|11574-1|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C2718236|T201|COMP|22574-8|LNC|Toxocara canis Ab.IgA|Toxocara canis Ab.IgA
C2718237|T201|COMP|22576-3|LNC|Toxocara canis Ab.IgM|Toxocara canis Ab.IgM
C2718238|T201|COMP|23490-6|LNC|Transmissible gastroenteritis virus Ab|Transmissible gastroenteritis virus Ab
C2718239|T201|COMP|22597-9|LNC|Trichinella spiralis Ab.IgA|Trichinella spiralis Ab.IgA
C2718240|T201|COMP|22598-7|LNC|Trichinella spiralis Ab.IgM|Trichinella spiralis Ab.IgM
C2718241|T201|COMP|7773-5|LNC|Triticum aestivum pollen Ab.IgE|Triticum aestivum pollen Ab.IgE
C2718242|T201|COMP|23525-9|LNC|Trypanosoma evansi Ab|Trypanosoma evansi Ab
C2718243|T201|COMP|24457-4|LNC|Tryptophan|Tryptophan
C2718244|T201|COMP|13166-4|LNC|Streptococcus pneumoniae 23 Ab|Streptococcus pneumoniae 23 Ab
C2718245|T201|COMP|26917-5|LNC|Streptococcus pneumoniae 23 Ab|Streptococcus pneumoniae 23 Ab
C2718246|T201|COMP|17624-8|LNC|Streptococcus pneumoniae 23f Ab^1st specimen|Streptococcus pneumoniae 23f Ab^1st specimen
C2718247|T201|COMP|29333-2|LNC|Saccharomonospora viridis Ab|Saccharomonospora viridis Ab
C2718248|T201|COMP|22508-6|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C2718249|T201|COMP|23430-2|LNC|Salmonella gallinarum Ab|Salmonella gallinarum Ab
C2718250|T201|COMP|7679-4|LNC|Salvia officinalis Ab.IgE|Salvia officinalis Ab.IgE
C2718251|T201|COMP|15695-0|LNC|Sambucus nigra Ab.IgE.RAST class|Sambucus nigra Ab.IgE.RAST class
C2718252|T201|COMP|7299-1|LNC|Sambucus nigra Ab.IgE|Sambucus nigra Ab.IgE
C2718253|T201|COMP|25594-3|LNC|Schistosoma sp Ab.IgG|Schistosoma sp Ab.IgG
C2718254|T201|COMP|6235-6|LNC|Secale cereale Ab.IgE|Secale cereale Ab.IgE
C2718255|T201|COMP|21504-6|LNC|Secale cereale Ab.IgG.RAST class|Secale cereale Ab.IgG.RAST class
C2718256|T201|COMP|15999-6|LNC|Secale cereale pollen Ab.IgE.RAST class|Secale cereale pollen Ab.IgE.RAST class
C2718257|T201|COMP|18375-6|LNC|Serotonin|Serotonin
C2718258|T201|COMP|5926-1|LNC|Sodium|Sodium
C2718259|T201|COMP|21478-3|LNC|Solanum tuberosum Ab.IgE.RAST class|Solanum tuberosum Ab.IgE.RAST class
C2718260|T201|COMP|7630-7|LNC|Solanum tuberosum Ab.IgG|Solanum tuberosum Ab.IgG
C2718261|T201|COMP|15538-2|LNC|Solenopsis invicta Ab.IgE.RAST class|Solenopsis invicta Ab.IgE.RAST class
C2718262|T201|COMP|7085-4|LNC|Solenopsis invicta Ab.IgE|Solenopsis invicta Ab.IgE
C2718264|T201|COMP|4434-7|LNC|Sulfonamide|Sulfonamide
C2718266|T201|COMP|23439-3|LNC|Swine vesicular disease virus Ab|Swine vesicular disease virus Ab
C2718272|T201|COMP|17612-3|LNC|Streptococcus pneumoniae 1 Ab^1st specimen|Streptococcus pneumoniae 1 Ab^1st specimen
C2718274|T201|COMP|22544-1|LNC|Streptococcus pneumoniae 14 Ab^1st specimen|Streptococcus pneumoniae 14 Ab^1st specimen
C2718275|T201|COMP|27388-8|LNC|Streptococcus pneumoniae 26 Ab.IgG|Streptococcus pneumoniae 26 Ab.IgG
C2718276|T201|COMP|17626-3|LNC|Streptococcus pneumoniae 3 Ab^1st specimen|Streptococcus pneumoniae 3 Ab^1st specimen
C2718277|T201|COMP|17628-9|LNC|Streptococcus pneumoniae 3 Ab^2nd specimen|Streptococcus pneumoniae 3 Ab^2nd specimen
C2718278|T201|COMP|17633-9|LNC|Streptococcus pneumoniae 4 Ab^1st specimen|Streptococcus pneumoniae 4 Ab^1st specimen
C2718279|T201|COMP|17634-7|LNC|Streptococcus pneumoniae 4 Ab^2nd specimen|Streptococcus pneumoniae 4 Ab^2nd specimen
C2718280|T201|COMP|27405-0|LNC|Streptococcus pneumoniae 56 Ab.IgG|Streptococcus pneumoniae 56 Ab.IgG
C2718281|T201|COMP|26941-5|LNC|Streptococcus pneumoniae 9 Ab|Streptococcus pneumoniae 9 Ab
C2718307|T201|COMP|55457-6|LNC|Hemoglobin.free|Hemoglobin.free
C2718308|T201|COMP|54300-9|LNC|Homocysteine|Homocysteine
C2718316|T201|COMP|55456-8|LNC|Hemoglobin S|Hemoglobin S
C2733654|T201|COMP|55767-8|LNC|EGFR gene.c.2582T>A|EGFR gene.c.2582T>A
C2733656|T201|COMP|55768-6|LNC|EGFR gene.c.2303G>T|EGFR gene.c.2303G>T
C2733658|T201|COMP|55769-4|LNC|EGFR gene.c.2369C>T|EGFR gene.c.2369C>T
C2733660|T201|COMP|55770-2|LNC|EGFR gene exon 20 insertion|EGFR gene exon 20 insertion
C2733662|T201|COMP|55771-0|LNC|Basophils|Basophils
C2733663|T201|COMP|55772-8|LNC|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C2733664|T201|COMP|55773-6|LNC|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C2733667|T201|COMP|55775-1|LNC|Direct antiglobulin test.IgA specific reagent|Direct antiglobulin test.IgA specific reagent
C2733669|T201|COMP|55776-9|LNC|Direct antiglobulin test.IgG specific reagent|Direct antiglobulin test.IgG specific reagent
C2733670|T201|COMP|55777-7|LNC|Direct antiglobulin test.IgM specific reagent|Direct antiglobulin test.IgM specific reagent
C2733672|T201|COMP|55778-5|LNC|Eosinophils|Eosinophils
C2733673|T201|COMP|55779-3|LNC|Erythrocytes|Erythrocytes
C2733674|T201|COMP|55780-1|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C2733675|T201|COMP|55781-9|LNC|Hematocrit|Hematocrit
C2733676|T201|COMP|55782-7|LNC|Hemoglobin|Hemoglobin
C2733677|T201|COMP|55783-5|LNC|Hemoglobin Barts|Hemoglobin Barts
C2733678|T201|COMP|55784-3|LNC|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C2733681|T201|COMP|55787-6|LNC|Lymphocytes|Lymphocytes
C2733682|T201|COMP|55788-4|LNC|Mononuclear cells|Mononuclear cells
C2733683|T201|COMP|55789-2|LNC|Myelocytes|Myelocytes
C2733684|T201|COMP|55790-0|LNC|Neutrophils.band form|Neutrophils.band form
C2733685|T201|COMP|55791-8|LNC|Neutrophils|Neutrophils
C2733686|T201|COMP|55792-6|LNC|Nucleated cells|Nucleated cells
C2733687|T201|COMP|55793-4|LNC|Nucleated cells|Nucleated cells
C2733688|T201|COMP|55794-2|LNC|Other cells|Other cells
C2733689|T201|COMP|55795-9|LNC|Phosphatidylserine Ab.IgG|Phosphatidylserine Ab.IgG
C2733690|T201|COMP|55796-7|LNC|Phosphatidylserine Ab.IgM|Phosphatidylserine Ab.IgM
C2733693|T201|COMP|55799-1|LNC|Platelet aggregation.ristocetin induced^1125 mg/L|Platelet aggregation.ristocetin induced^1125 mg/L
C2733694|T201|COMP|55800-7|LNC|Platelet aggregation.ristocetin induced^1000 mg/L|Platelet aggregation.ristocetin induced^1000 mg/L
C2733695|T201|COMP|55801-5|LNC|Platelet aggregation.ristocetin induced^500 mg/L|Platelet aggregation.ristocetin induced^500 mg/L
C2733696|T201|COMP|55802-3|LNC|Platelets|Platelets
C2733697|T201|COMP|55803-1|LNC|Promyelocytes|Promyelocytes
C2733698|T201|COMP|55804-9|LNC|Phosphatase.leukocyte|Phosphatase.leukocyte
C2733699|T201|COMP|55805-6|LNC|cycloSPORINE|cycloSPORINE
C2733700|T201|COMP|55806-4|LNC|Mycophenolate|Mycophenolate
C2733701|T201|COMP|55807-2|LNC|Mycophenolate glucuronide|Mycophenolate glucuronide
C2733702|T201|COMP|55808-0|LNC|11-Deoxycorticosterone|11-Deoxycorticosterone
C2733703|T201|COMP|55809-8|LNC|11-Deoxycortisol|11-Deoxycortisol
C2733704|T201|COMP|55810-6|LNC|18-Hydroxycortisol|18-Hydroxycortisol
C2733705|T201|COMP|55811-4|LNC|18-Hydroxycortisol|18-Hydroxycortisol
C2733706|T201|COMP|55812-2|LNC|18-Hydroxycortisol|18-Hydroxycortisol
C2733707|T201|COMP|55813-0|LNC|Alpha aminobutyrate/Amino acids.total|Alpha aminobutyrate/Amino acids.total
C2733709|T201|COMP|55814-8|LNC|Calcidiol|Calcidiol
C2733710|T201|COMP|55815-5|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C2733711|T201|COMP|55816-3|LNC|3,4-Dihydroxyphenylacetate|3,4-Dihydroxyphenylacetate
C2733712|T201|COMP|55817-1|LNC|Amino acids|Amino acids
C2733713|T201|COMP|55818-9|LNC|Organic acids|Organic acids
C2733714|T201|COMP|55819-7|LNC|Adiponectin.high molecular weight|Adiponectin.high molecular weight
C2733716|T201|COMP|55820-5|LNC|Allo-pregnanediol|Allo-pregnanediol
C2733718|T201|COMP|55821-3|LNC|Allo-pregnanediol|Allo-pregnanediol
C2733719|T201|COMP|55822-1|LNC|Allo-tetrahydrodeoxycortisol|Allo-tetrahydrodeoxycortisol
C2733720|T201|COMP|55823-9|LNC|Allo-tetrahydrodeoxycortisol|Allo-tetrahydrodeoxycortisol
C2733721|T201|COMP|55824-7|LNC|Allo-tetrahydrocorticosterone|Allo-tetrahydrocorticosterone
C2733723|T201|COMP|55825-4|LNC|Allo-tetrahydrocorticosterone|Allo-tetrahydrocorticosterone
C2733724|T201|COMP|55826-2|LNC|Allo-tetrahydrocortisol|Allo-tetrahydrocortisol
C2733725|T201|COMP|55827-0|LNC|Acid alpha glucosidase|Acid alpha glucosidase
C2733726|T201|COMP|55828-8|LNC|Aliphatic carboxylate C14-C26.esters|Aliphatic carboxylate C14-C26.esters
C2733727|T201|COMP|55829-6|LNC|Catalase|Catalase
C2733728|T201|COMP|55830-4|LNC|Catecholamines|Catecholamines
C2733729|T201|COMP|55831-2|LNC|Catecholamines|Catecholamines
C2733730|T201|COMP|55832-0|LNC|Cathepsin K|Cathepsin K
C2733731|T201|COMP|55833-8|LNC|Cathepsin L|Cathepsin L
C2733732|T201|COMP|55834-6|LNC|Cathepsin S|Cathepsin S
C2733733|T201|COMP|55835-3|LNC|Vegetable fibers|Vegetable fibers
C2733734|T201|COMP|56009-4|LNC|Platelet aggregation.collagen induced^5 ug/mL|Platelet aggregation.collagen induced^5 ug/mL
C2733735|T201|COMP|56010-2|LNC|Platelet aggregation.ristocetin induced^250 ug/mL|Platelet aggregation.ristocetin induced^250 ug/mL
C2733743|T201|COMP|56180-3|LNC|Aspergillus fumigatus Ab.IgG4|Aspergillus fumigatus Ab.IgG4
C2733744|T201|COMP|56181-1|LNC|Aspergillus niger Ab.IgG4|Aspergillus niger Ab.IgG4
C2733746|T201|COMP|56182-9|LNC|Aspergillus versicolor Ab.IgG4|Aspergillus versicolor Ab.IgG4
C2733748|T201|COMP|56183-7|LNC|Casuarina equisetifolia Ab.IgG4|Casuarina equisetifolia Ab.IgG4
C2733750|T201|COMP|56184-5|LNC|Persea americana Ab.IgG4|Persea americana Ab.IgG4
C2733752|T201|COMP|56185-2|LNC|Paspalum notatum Ab.IgG4|Paspalum notatum Ab.IgG4
C2733754|T201|COMP|56186-0|LNC|Musa spp Ab.IgG4|Musa spp Ab.IgG4
C2733756|T201|COMP|56187-8|LNC|Hordeum vulgare Ab.IgG4|Hordeum vulgare Ab.IgG4
C2733758|T201|COMP|56357-7|LNC|Lolium perenne Ab.IgG4|Lolium perenne Ab.IgG4
C2733760|T201|COMP|56358-5|LNC|Ananas comosus Ab.IgG4|Ananas comosus Ab.IgG4
C2733762|T201|COMP|56359-3|LNC|Bean pinto Ab.IgG4|Bean pinto Ab.IgG4
C2733764|T201|COMP|56360-1|LNC|Pistacia vera Ab.IgG4|Pistacia vera Ab.IgG4
C2733766|T201|COMP|56361-9|LNC|Prunus domestica Ab.IgG4|Prunus domestica Ab.IgG4
C2733768|T201|COMP|56362-7|LNC|Papaver somniferum Ab.IgG4|Papaver somniferum Ab.IgG4
C2733770|T201|COMP|56363-5|LNC|Insulin porcine Ab.IgG4|Insulin porcine Ab.IgG4
C2733772|T201|COMP|56364-3|LNC|Iva axillaris Ab.IgG4|Iva axillaris Ab.IgG4
C2733774|T201|COMP|56687-7|LNC|Pancreatic islet cell Ab.IgG|Pancreatic islet cell Ab.IgG
C2733775|T201|COMP|56688-5|LNC|IgD|IgD
C2733776|T201|COMP|56689-3|LNC|Isoleucine/Creatinine|Isoleucine/Creatinine
C2733777|T201|COMP|56690-1|LNC|Insulin^16H post XXX challenge|Insulin^16H post XXX challenge
C2733778|T201|COMP|56691-9|LNC|Insulin^20H post XXX challenge|Insulin^20H post XXX challenge
C2733779|T201|COMP|56692-7|LNC|Insulin^1D post XXX challenge|Insulin^1D post XXX challenge
C2733780|T201|COMP|56693-5|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C2733781|T201|COMP|56950-9|LNC|Legionella pneumophila Ab.IgG^2nd specimen|Legionella pneumophila Ab.IgG^2nd specimen
C2733782|T201|COMP|56951-7|LNC|Leishmania sp Ab.IgG|Leishmania sp Ab.IgG
C2733783|T201|COMP|56952-5|LNC|Leptospira interrogans Ab|Leptospira interrogans Ab
C2733784|T201|COMP|56953-3|LNC|Leptospira interrogans Ab.IgM|Leptospira interrogans Ab.IgM
C2733786|T201|COMP|56954-1|LNC|Leucine/Creatinine|Leucine/Creatinine
C2733787|T201|COMP|56955-8|LNC|Lysine/Creatinine|Lysine/Creatinine
C2733788|T201|COMP|56956-6|LNC|Magnesium/Creatinine|Magnesium/Creatinine
C2733803|T201|COMP|55836-1|LNC|Chitotriosidase|Chitotriosidase
C2733804|T201|COMP|55837-9|LNC|Chloride|Chloride
C2733805|T201|COMP|55838-7|LNC|Cholesterol/Phospholipid|Cholesterol/Phospholipid
C2733807|T201|COMP|55839-5|LNC|Cholesterol ester transfer protein|Cholesterol ester transfer protein
C2733808|T201|COMP|55840-3|LNC|Cholesterol esters|Cholesterol esters
C2733809|T201|COMP|55841-1|LNC|Corticosterone|Corticosterone
C2733810|T201|COMP|55842-9|LNC|Corticosterone|Corticosterone
C2733811|T201|COMP|55843-7|LNC|Corticosterone|Corticosterone
C2733812|T201|COMP|55844-5|LNC|Cortisol.free|Cortisol.free
C2733813|T201|COMP|55845-2|LNC|Cortisol.free|Cortisol.free
C2733814|T201|COMP|55846-0|LNC|Cryoglobulin.IgA.monoclonal|Cryoglobulin.IgA.monoclonal
C2733816|T201|COMP|55847-8|LNC|Cryoglobulin.IgG.monoclonal|Cryoglobulin.IgG.monoclonal
C2733818|T201|COMP|55848-6|LNC|Cryoglobulin.IgG|Cryoglobulin.IgG
C2733819|T201|COMP|55849-4|LNC|Cryoglobulin.IgM.monoclonal|Cryoglobulin.IgM.monoclonal
C2733821|T201|COMP|55850-2|LNC|Cobalamins|Cobalamins
C2733822|T201|COMP|55851-0|LNC|Androstenediol|Androstenediol
C2733823|T201|COMP|55852-8|LNC|Dicarboxydodecanoylcarnitine (C12-DC)/Creatinine|Dicarboxydodecanoylcarnitine (C12-DC)/Creatinine
C2733825|T201|COMP|55853-6|LNC|Dicarboxydodecanoylcarnitine (C12-DC)|Dicarboxydodecanoylcarnitine (C12-DC)
C2733826|T201|COMP|55854-4|LNC|Dicarboxydodecanoylcarnitine (C12-DC)|Dicarboxydodecanoylcarnitine (C12-DC)
C2733827|T201|COMP|55855-1|LNC|Dicarboxydodecanoylcarnitine (C12-DC)|Dicarboxydodecanoylcarnitine (C12-DC)
C2733828|T201|COMP|55856-9|LNC|Dicarboxydodecanoylcarnitine (C12-DC)|Dicarboxydodecanoylcarnitine (C12-DC)
C2733829|T201|COMP|55857-7|LNC|Estradiol|Estradiol
C2733830|T201|COMP|55858-5|LNC|Estradiol|Estradiol
C2733831|T201|COMP|55859-3|LNC|Folate|Folate
C2733832|T201|COMP|55860-1|LNC|Glucose|Glucose
C2733833|T201|COMP|55861-9|LNC|Glutamate|Glutamate
C2733834|T201|COMP|55862-7|LNC|Glycine|Glycine
C2733835|T201|COMP|55863-5|LNC|Glycolate|Glycolate
C2733836|T201|COMP|55864-3|LNC|Glycolate|Glycolate
C2733837|T201|COMP|55865-0|LNC|Glycolate|Glycolate
C2733838|T201|COMP|55866-8|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C2733839|T201|COMP|55867-6|LNC|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C2733840|T201|COMP|55868-4|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C2733841|T201|COMP|55869-2|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C2733842|T201|COMP|55870-0|LNC|Choriogonadotropin|Choriogonadotropin
C2733843|T201|COMP|55871-8|LNC|Heptanoylcarnitine (C7)|Heptanoylcarnitine (C7)
C2733844|T201|COMP|55872-6|LNC|Dicarboxypalmitoylcarnitine (C16-DC)|Dicarboxypalmitoylcarnitine (C16-DC)
C2733845|T201|COMP|55873-4|LNC|Palmitate/Laurate|Palmitate/Laurate
C2733847|T201|COMP|55874-2|LNC|Histidine|Histidine
C2733848|T201|COMP|55875-9|LNC|Homocitrulline|Homocitrulline
C2733849|T201|COMP|55876-7|LNC|Homocitrulline|Homocitrulline
C2733850|T201|COMP|55877-5|LNC|Homocysteine|Homocysteine
C2733851|T201|COMP|55878-3|LNC|Homocysteine|Homocysteine
C2733852|T201|COMP|55879-1|LNC|Homocystine|Homocystine
C2733853|T201|COMP|55880-9|LNC|Homovanillate|Homovanillate
C2733854|T201|COMP|55881-7|LNC|Hydroxocobalamin|Hydroxocobalamin
C2733855|T201|COMP|55882-5|LNC|Hydroxocobalamin|Hydroxocobalamin
C2733856|T201|COMP|55883-3|LNC|Hydroxocobalamin|Hydroxocobalamin
C2733857|T201|COMP|55884-1|LNC|Hydroxocobalamin|Hydroxocobalamin
C2733858|T201|COMP|55885-8|LNC|Hydroxocobalamin|Hydroxocobalamin
C2733859|T201|COMP|55886-6|LNC|3-Hydroxyanthranilate/Creatinine|3-Hydroxyanthranilate/Creatinine
C2733861|T201|COMP|55887-4|LNC|3-Hydroxyanthranilate|3-Hydroxyanthranilate
C2733863|T201|COMP|55888-2|LNC|3-Hydroxyanthranilate|3-Hydroxyanthranilate
C2733864|T201|COMP|55889-0|LNC|3-Hydroxyanthranilate|3-Hydroxyanthranilate
C2733865|T201|COMP|55890-8|LNC|Hydroxylysine/Amino acids.total|Hydroxylysine/Amino acids.total
C2733867|T201|COMP|55891-6|LNC|Hydroxylysine|Hydroxylysine
C2733873|T201|COMP|55896-5|LNC|Hypoxanthine phosphoribosyltransferase|Hypoxanthine phosphoribosyltransferase
C2733874|T201|COMP|55897-3|LNC|Immunoglobulin light chains.free|Immunoglobulin light chains.free
C2733875|T201|COMP|55898-1|LNC|Immunoglobulin light chains.free|Immunoglobulin light chains.free
C2733876|T201|COMP|55899-9|LNC|Immunoglobulin light chains.free|Immunoglobulin light chains.free
C2733877|T201|COMP|55900-5|LNC|Immunoglobulin light chains.free|Immunoglobulin light chains.free
C2733878|T201|COMP|55901-3|LNC|IgA.monoclonal|IgA.monoclonal
C2733879|T201|COMP|55902-1|LNC|IgA|IgA
C2733880|T201|COMP|55903-9|LNC|IgD.monoclonal|IgD.monoclonal
C2733881|T201|COMP|55904-7|LNC|IgE.monoclonal|IgE.monoclonal
C2733882|T201|COMP|55905-4|LNC|Alpha cortol|Alpha cortol
C2733883|T201|COMP|55914-6|LNC|Beta 1 globulin|Beta 1 globulin
C2733884|T201|COMP|55915-3|LNC|Beta 2 globulin|Beta 2 globulin
C2733885|T201|COMP|55916-1|LNC|Beta galactosidase|Beta galactosidase
C2733886|T201|COMP|55917-9|LNC|Glucosylceramidase|Glucosylceramidase
C2733887|T201|COMP|55918-7|LNC|C peptide^post meal|C peptide^post meal
C2733888|T201|COMP|55919-5|LNC|C peptide^post meal|C peptide^post meal
C2733889|T201|COMP|55920-3|LNC|C peptide|C peptide
C2733890|T201|COMP|55921-1|LNC|IgG.monoclonal|IgG.monoclonal
C2733891|T201|COMP|55922-9|LNC|IgG|IgG
C2733892|T201|COMP|55923-7|LNC|IgG|IgG
C2733893|T201|COMP|55924-5|LNC|IgM.monoclonal|IgM.monoclonal
C2733894|T201|COMP|55925-2|LNC|IgM|IgM
C2733895|T201|COMP|55926-0|LNC|Interleukin 1 receptor alpha chain|Interleukin 1 receptor alpha chain
C2733897|T201|COMP|55927-8|LNC|Interleukin 1 receptor alpha chain.soluble|Interleukin 1 receptor alpha chain.soluble
C2733899|T201|COMP|55928-6|LNC|Iodine/Creatinine|Iodine/Creatinine
C2733900|T201|COMP|55929-4|LNC|Isoleucine|Isoleucine
C2733901|T201|COMP|55930-2|LNC|Isovalerylglycine|Isovalerylglycine
C2733902|T201|COMP|55931-0|LNC|Lactate|Lactate
C2733903|T201|COMP|55932-8|LNC|Lactate|Lactate
C2733904|T201|COMP|55933-6|LNC|Leucine|Leucine
C2733905|T201|COMP|55934-4|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C2733906|T201|COMP|55935-1|LNC|Lysine|Lysine
C2733907|T201|COMP|55936-9|LNC|Lysozyme|Lysozyme
C2733908|T201|COMP|55937-7|LNC|Magnesium^post dialysis|Magnesium^post dialysis
C2733909|T201|COMP|55938-5|LNC|Magnesium|Magnesium
C2733910|T201|COMP|55939-3|LNC|Malondialdehyde|Malondialdehyde
C2733911|T201|COMP|55940-1|LNC|Malonylcarnitine (C3-DC)|Malonylcarnitine (C3-DC)
C2733912|T201|COMP|55941-9|LNC|Mannitol|Mannitol
C2733913|T201|COMP|55942-7|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C2733914|T201|COMP|55943-5|LNC|Methionine|Methionine
C2733915|T201|COMP|55966-6|LNC|Palmitoleylcarnitine (C16:1)|Palmitoleylcarnitine (C16:1)
C2733916|T201|COMP|55967-4|LNC|Palmitoylcarnitine (C16)|Palmitoylcarnitine (C16)
C2733918|T201|COMP|55969-0|LNC|Phenylalanine/Amino acids.total|Phenylalanine/Amino acids.total
C2733919|T201|COMP|55970-8|LNC|Phenylalanine|Phenylalanine
C2733920|T201|COMP|55971-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C2733921|T201|COMP|55972-4|LNC|Phosphate^post dialysis|Phosphate^post dialysis
C2733922|T201|COMP|55973-2|LNC|Phosphate|Phosphate
C2733923|T201|COMP|55974-0|LNC|IgG|IgG
C2733924|T201|COMP|55975-7|LNC|IgG|IgG
C2733957|T201|COMP|56008-6|LNC|Platelet aggregation.collagen induced^1 ug/mL|Platelet aggregation.collagen induced^1 ug/mL
C2733966|T201|COMP|56022-7|LNC|ACE gene targeted mutation analysis|ACE gene targeted mutation analysis
C2733968|T201|COMP|56023-5|LNC|Foot and mouth disease virus RNA|Foot and mouth disease virus RNA
C2733969|T201|COMP|56024-3|LNC|Influenza virus A N1 RNA|Influenza virus A N1 RNA
C2733971|T201|COMP|56025-0|LNC|Ethambutol 8.0 ug/mL|Ethambutol 8.0 ug/mL
C2733973|T201|COMP|56026-8|LNC|Pyrazinamide 300.0 ug/mL|Pyrazinamide 300.0 ug/mL
C2733975|T201|COMP|56027-6|LNC|Platelet aggregation.ristocetin induced^1.0 mg/mL|Platelet aggregation.ristocetin induced^1.0 mg/mL
C2733976|T201|COMP|56028-4|LNC|Cells.CD3-CD56+/100 cells|Cells.CD3-CD56+/100 cells
C2733977|T201|COMP|56029-2|LNC|Cells.CD3-CD56+/100 cells|Cells.CD3-CD56+/100 cells
C2733978|T201|COMP|56030-0|LNC|Karyotype|Karyotype
C2733979|T201|COMP|56031-8|LNC|Doripenem|Doripenem
C2733980|T201|COMP|56032-6|LNC|Lithium|Lithium
C2733981|T201|COMP|56033-4|LNC|Androstenediol|Androstenediol
C2733982|T201|COMP|56034-2|LNC|Hydroxylysine|Hydroxylysine
C2733983|T201|COMP|56035-9|LNC|Apolipoprotein A-I/Cholesterol.in HDL|Apolipoprotein A-I/Cholesterol.in HDL
C2733985|T201|COMP|56036-7|LNC|Apolipoprotein B/Cholesterol.in LDL|Apolipoprotein B/Cholesterol.in LDL
C2733987|T201|COMP|56037-5|LNC|Protein phosphatase 3|Protein phosphatase 3
C2733988|T201|COMP|56038-3|LNC|Lysozyme|Lysozyme
C2733989|T201|COMP|56039-1|LNC|Lysozyme|Lysozyme
C2733990|T201|COMP|56040-9|LNC|Methemoglobin|Methemoglobin
C2733991|T201|COMP|56041-7|LNC|Beta defensin|Beta defensin
C2733993|T201|COMP|56042-5|LNC|Beta defensin|Beta defensin
C2734072|T201|COMP|56119-1|LNC|Cellular material|Cellular material
C2734074|T201|COMP|56120-9|LNC|Amphetamine+Methamphetamine|Amphetamine+Methamphetamine
C2734075|T201|COMP|56121-7|LNC|IgA|IgA
C2734076|T201|COMP|56122-5|LNC|IgG|IgG
C2734077|T201|COMP|56123-3|LNC|IgM|IgM
C2734078|T201|COMP|56124-1|LNC|Glucose^1H post meal|Glucose^1H post meal
C2734079|T201|COMP|56125-8|LNC|Immunoglobulin light chains.free|Immunoglobulin light chains.free
C2734080|T201|COMP|56126-6|LNC|Copper|Copper
C2734081|T201|COMP|56127-4|LNC|CD38 Ag|CD38 Ag
C2734082|T201|COMP|56128-2|LNC|Chikungunya virus Ab.IgG|Chikungunya virus Ab.IgG
C2734084|T201|COMP|56129-0|LNC|Chikungunya virus Ab.IgG|Chikungunya virus Ab.IgG
C2734085|T201|COMP|56130-8|LNC|Chikungunya virus Ab.IgM|Chikungunya virus Ab.IgM
C2734087|T201|COMP|56131-6|LNC|Chikungunya virus Ab.IgM|Chikungunya virus Ab.IgM
C2734088|T201|COMP|56132-4|LNC|Cholesterol.in HDL 2a|Cholesterol.in HDL 2a
C2734089|T201|COMP|56133-2|LNC|Cholesterol.in HDL 2b|Cholesterol.in HDL 2b
C2734090|T201|COMP|56134-0|LNC|Cholesterol.in IDL 1|Cholesterol.in IDL 1
C2734092|T201|COMP|56135-7|LNC|Cholesterol.in IDL 2|Cholesterol.in IDL 2
C2734094|T201|COMP|56136-5|LNC|LDL 1|LDL 1
C2734095|T201|COMP|56137-3|LNC|LDL 2|LDL 2
C2734096|T201|COMP|56138-1|LNC|LDL 3|LDL 3
C2734097|T201|COMP|56139-9|LNC|LDL 4|LDL 4
C2734099|T201|COMP|56141-5|LNC|MPL gene.p.Ser505Asn|MPL gene.p.Ser505Asn
C2734101|T201|COMP|56142-3|LNC|MPL gene.p.Trp515Leu+Trp515Lys|MPL gene.p.Trp515Leu+Trp515Lys
C2734103|T201|COMP|56143-1|LNC|Potassium/Creatinine|Potassium/Creatinine
C2734104|T201|COMP|56144-9|LNC|CHIC2 gene 4q12 deletion|CHIC2 gene 4q12 deletion
C2734106|T201|COMP|56145-6|LNC|Erythrocytes+Granulocytes.CD55+CD59 deficient|Erythrocytes+Granulocytes.CD55+CD59 deficient
C2734108|T201|COMP|56146-4|LNC|Fungal Ab panel|Fungal Ab panel
C2734110|T201|COMP|56147-2|LNC|Parietal cell Ab|Parietal cell Ab
C2734115|T201|COMP|56150-6|LNC|Candida albicans Ab.IgM|Candida albicans Ab.IgM
C2734117|T201|COMP|56151-4|LNC|Candida albicans Ab.IgA|Candida albicans Ab.IgA
C2734119|T201|COMP|56152-2|LNC|Beta 2 glycoprotein 1 Ab.IgA & IgG & IgM panel|Beta 2 glycoprotein 1 Ab.IgA & IgG & IgM panel
C2734121|T201|COMP|56153-0|LNC|Albumin.serum/Albumin.Periton fld|Albumin.serum/Albumin.Periton fld
C2734123|T201|COMP|56154-8|LNC|Protein.abnormal band/Protein.total|Protein.abnormal band/Protein.total
C2734124|T201|COMP|56155-5|LNC|Date reference lab test results received|Date reference lab test results received
C2734127|T201|COMP|56157-1|LNC|HOXB13 gene/IL17BR gene|HOXB13 gene/IL17BR gene
C2734129|T201|COMP|56158-9|LNC|PCSK9 gene targeted mutation analysis|PCSK9 gene targeted mutation analysis
C2734131|T201|COMP|56159-7|LNC|LDLR gene targeted mutation analysis|LDLR gene targeted mutation analysis
C2734133|T201|COMP|56160-5|LNC|Glucose^4H post peritoneal dialysis|Glucose^4H post peritoneal dialysis
C2734134|T201|COMP|56161-3|LNC|Calculus analysis with calculus photography|Calculus analysis with calculus photography
C2734139|T201|COMP|56164-7|LNC|CYP2C9 gene allele 2|CYP2C9 gene allele 2
C2734141|T201|COMP|56165-4|LNC|CYP2C9 gene allele 3|CYP2C9 gene allele 3
C2734143|T201|COMP|56166-2|LNC|Gum arabic Ab.IgG4|Gum arabic Ab.IgG4
C2734145|T201|COMP|56167-0|LNC|Corticotropin Ab.IgG4|Corticotropin Ab.IgG4
C2734147|T201|COMP|56168-8|LNC|Pimenta dioica Ab.IgG4|Pimenta dioica Ab.IgG4
C2734149|T201|COMP|56169-6|LNC|Prunus dulcis Ab.IgG4|Prunus dulcis Ab.IgG4
C2734151|T201|COMP|56170-4|LNC|Alternaria alternata Ab.IgG4|Alternaria alternata Ab.IgG4
C2734152|T201|COMP|56171-2|LNC|Fagus grandifolia Ab.IgG4|Fagus grandifolia Ab.IgG4
C2734154|T201|COMP|56172-0|LNC|Cheese American Ab.IgG4|Cheese American Ab.IgG4
C2734156|T201|COMP|56173-8|LNC|Periplaneta americana Ab.IgG4|Periplaneta americana Ab.IgG4
C2734158|T201|COMP|56174-6|LNC|Ulmus americana Ab.IgG4|Ulmus americana Ab.IgG4
C2734160|T201|COMP|56175-3|LNC|Platanus occidentalis Ab.IgG4|Platanus occidentalis Ab.IgG4
C2734162|T201|COMP|56176-1|LNC|Malus sylvestris Ab.IgG4|Malus sylvestris Ab.IgG4
C2734164|T201|COMP|56177-9|LNC|Prunus armeniaca Ab.IgG4|Prunus armeniaca Ab.IgG4
C2734166|T201|COMP|56178-7|LNC|Cynara scolymus Ab.IgG4|Cynara scolymus Ab.IgG4
C2734168|T201|COMP|56179-5|LNC|Asparagus officinalis Ab.IgG4|Asparagus officinalis Ab.IgG4
C2734170|T201|COMP|56188-6|LNC|Ocimum basilicum Ab.IgG4|Ocimum basilicum Ab.IgG4
C2734172|T201|COMP|56189-4|LNC|Laurus nobilis Ab.IgG4|Laurus nobilis Ab.IgG4
C2734174|T201|COMP|56190-2|LNC|Cynodon dactylon Ab.IgG4|Cynodon dactylon Ab.IgG4
C2734176|T201|COMP|56191-0|LNC|Prunus avium Ab.IgG4|Prunus avium Ab.IgG4
C2734178|T201|COMP|56192-8|LNC|Micropterus salmoides Ab.IgG4|Micropterus salmoides Ab.IgG4
C2734180|T201|COMP|56193-6|LNC|Salix nigra Ab.IgG4|Salix nigra Ab.IgG4
C2734182|T201|COMP|56194-4|LNC|Rubus fruticosus Ab.IgG4|Rubus fruticosus Ab.IgG4
C2734184|T201|COMP|56195-1|LNC|Vigna sinensis Ab.IgG4|Vigna sinensis Ab.IgG4
C2734186|T201|COMP|56196-9|LNC|Vaccinium myrtillus Ab.IgG4|Vaccinium myrtillus Ab.IgG4
C2734188|T201|COMP|56197-7|LNC|Insulin bovine Ab.IgG4|Insulin bovine Ab.IgG4
C2734190|T201|COMP|56198-5|LNC|Bertholletia excelsa Ab.IgG4|Bertholletia excelsa Ab.IgG4
C2734192|T201|COMP|56199-3|LNC|Yeast brewer's Ab.IgG4|Yeast brewer's Ab.IgG4
C2734194|T201|COMP|56200-9|LNC|Brassica oleracea var italica Ab.IgG4|Brassica oleracea var italica Ab.IgG4
C2734196|T201|COMP|56201-7|LNC|Brassica oleracea var gemmifera Ab.IgG4|Brassica oleracea var gemmifera Ab.IgG4
C2734198|T201|COMP|56202-5|LNC|Fagopyrum esculentum Ab.IgG4|Fagopyrum esculentum Ab.IgG4
C2734200|T201|COMP|56203-3|LNC|Brassica oleracea var capitata Ab.IgG4|Brassica oleracea var capitata Ab.IgG4
C2734202|T201|COMP|56204-1|LNC|Candida albicans Ab.IgG4|Candida albicans Ab.IgG4
C2734203|T201|COMP|56205-8|LNC|Amaranthus palmeri Ab.IgG4|Amaranthus palmeri Ab.IgG4
C2734205|T201|COMP|56206-6|LNC|Daucus carota Ab.IgG4|Daucus carota Ab.IgG4
C2734207|T201|COMP|56207-4|LNC|Casein Ab.IgG4|Casein Ab.IgG4
C2734208|T201|COMP|56208-2|LNC|Anacardium occidentale Ab.IgG4|Anacardium occidentale Ab.IgG4
C2734210|T201|COMP|56209-0|LNC|Ricinus communis Ab.IgG4|Ricinus communis Ab.IgG4
C2734212|T201|COMP|56210-8|LNC|Cat dander Ab.IgG4|Cat dander Ab.IgG4
C2734214|T201|COMP|56211-6|LNC|Ictalurus punctatus Ab.IgG4|Ictalurus punctatus Ab.IgG4
C2734216|T201|COMP|56212-4|LNC|Brassica oleracea var botrytis Ab.IgG4|Brassica oleracea var botrytis Ab.IgG4
C2734218|T201|COMP|56213-2|LNC|Apium graveolens Ab.IgG4|Apium graveolens Ab.IgG4
C2734220|T201|COMP|56214-0|LNC|Acremonium sp Ab.IgG4|Acremonium sp Ab.IgG4
C2734222|T201|COMP|56215-7|LNC|Cheese cheddar type Ab.IgG4|Cheese cheddar type Ab.IgG4
C2734224|T201|COMP|56216-5|LNC|Cheese mold type Ab.IgG4|Cheese mold type Ab.IgG4
C2734226|T201|COMP|56217-3|LNC|Cicer arietinus Ab.IgG4|Cicer arietinus Ab.IgG4
C2734228|T201|COMP|56218-1|LNC|Chicken Ab.IgG4|Chicken Ab.IgG4
C2734230|T201|COMP|56219-9|LNC|Cichorium intybus Ab.IgG4|Cichorium intybus Ab.IgG4
C2734232|T201|COMP|56220-7|LNC|Capsicum frutescens Ab.IgG4|Capsicum frutescens Ab.IgG4
C2734234|T201|COMP|56221-5|LNC|Ulmus pumila Ab.IgG4|Ulmus pumila Ab.IgG4
C2734236|T201|COMP|56222-3|LNC|Chocolate Ab.IgG4|Chocolate Ab.IgG4
C2734238|T201|COMP|56231-4|LNC|Zea mays Ab.IgG4|Zea mays Ab.IgG4
C2734240|T201|COMP|56232-2|LNC|Ustilago maydis Ab.IgG4|Ustilago maydis Ab.IgG4
C2734242|T201|COMP|56233-0|LNC|Populus deltoides Ab.IgG4|Populus deltoides Ab.IgG4
C2734244|T201|COMP|56234-8|LNC|Cow milk Ab.IgG4|Cow milk Ab.IgG4
C2734246|T201|COMP|56235-5|LNC|Cancer pagurus Ab.IgG4|Cancer pagurus Ab.IgG4
C2734248|T201|COMP|56236-3|LNC|Vaccinium oxycoccos Ab.IgG4|Vaccinium oxycoccos Ab.IgG4
C2734250|T201|COMP|56237-1|LNC|Astacus astacus Ab.IgG4|Astacus astacus Ab.IgG4
C2734252|T201|COMP|56238-9|LNC|Cucumis sativus Ab.IgG4|Cucumis sativus Ab.IgG4
C2734254|T201|COMP|56239-7|LNC|Curry Ab.IgG4|Curry Ab.IgG4
C2734256|T201|COMP|56240-5|LNC|Loligo sp Ab.IgG4|Loligo sp Ab.IgG4
C2734258|T201|COMP|56241-3|LNC|Dermatophagoides farinae Ab.IgG4|Dermatophagoides farinae Ab.IgG4
C2734259|T201|COMP|56242-1|LNC|Dermatophagoides pteronyssinus Ab.IgG4|Dermatophagoides pteronyssinus Ab.IgG4
C2734260|T201|COMP|56243-9|LNC|Taraxacum vulgare Ab.IgG4|Taraxacum vulgare Ab.IgG4
C2734262|T201|COMP|56244-7|LNC|Phoenix dactylifera Ab.IgG4|Phoenix dactylifera Ab.IgG4
C2734264|T201|COMP|56245-4|LNC|Chrysops flavidus (whole body) Ab.IgG4|Chrysops flavidus (whole body) Ab.IgG4
C2734266|T201|COMP|56246-2|LNC|Anethum graveolens Ab.IgG4|Anethum graveolens Ab.IgG4
C2734268|T201|COMP|56247-0|LNC|Dog epithelium Ab.IgG4|Dog epithelium Ab.IgG4
C2734270|T201|COMP|56248-8|LNC|Dog dander Ab.IgG4|Dog dander Ab.IgG4
C2734272|T201|COMP|56249-6|LNC|Pseudotsuga taxifolia Ab.IgG4|Pseudotsuga taxifolia Ab.IgG4
C2734274|T201|COMP|56250-4|LNC|Duck feather Ab.IgG4|Duck feather Ab.IgG4
C2734276|T201|COMP|56251-2|LNC|Duck meat Ab.IgG4|Duck meat Ab.IgG4
C2734278|T201|COMP|56252-0|LNC|Anguilla anguilla Ab.IgG4|Anguilla anguilla Ab.IgG4
C2734280|T201|COMP|56261-1|LNC|Linum usitatissimum Ab.IgG4|Linum usitatissimum Ab.IgG4
C2734282|T201|COMP|56262-9|LNC|Ctenocephalides sp Ab.IgG4|Ctenocephalides sp Ab.IgG4
C2734284|T201|COMP|56263-7|LNC|Flounder Ab.IgG4|Flounder Ab.IgG4
C2734286|T201|COMP|56264-5|LNC|Glycyphagus domesticus Ab.IgG4|Glycyphagus domesticus Ab.IgG4
C2734288|T201|COMP|56265-2|LNC|Allium sativum Ab.IgG4|Allium sativum Ab.IgG4
C2734290|T201|COMP|56266-0|LNC|Blatella germanica Ab.IgG4|Blatella germanica Ab.IgG4
C2734292|T201|COMP|56267-8|LNC|Zingiber officinale Ab.IgG4|Zingiber officinale Ab.IgG4
C2734294|T201|COMP|56268-6|LNC|Gluten Ab.IgG4|Gluten Ab.IgG4
C2734296|T201|COMP|56269-4|LNC|Goat milk Ab.IgG4|Goat milk Ab.IgG4
C2734298|T201|COMP|56270-2|LNC|Hamster epithelium Ab.IgG4|Hamster epithelium Ab.IgG4
C2734300|T201|COMP|56271-0|LNC|Solidago virgaurea Ab.IgG4|Solidago virgaurea Ab.IgG4
C2734302|T201|COMP|56272-8|LNC|Goose feather Ab.IgG4|Goose feather Ab.IgG4
C2734304|T201|COMP|56273-6|LNC|Vitis vinifera Ab.IgG4|Vitis vinifera Ab.IgG4
C2734306|T201|COMP|56274-4|LNC|Citrus paradisis Ab.IgG4|Citrus paradisis Ab.IgG4
C2734308|T201|COMP|56275-1|LNC|Bean green Ab.IgG4|Bean green Ab.IgG4
C2734310|T201|COMP|56276-9|LNC|Olea europaea Ab.IgG4|Olea europaea Ab.IgG4
C2734312|T201|COMP|56277-7|LNC|Pisum sativum Ab.IgG4|Pisum sativum Ab.IgG4
C2734314|T201|COMP|56278-5|LNC|Pepper green Ab.IgG4|Pepper green Ab.IgG4
C2734316|T201|COMP|56279-3|LNC|Guinea pig epithelium Ab.IgG4|Guinea pig epithelium Ab.IgG4
C2734318|T201|COMP|56280-1|LNC|Melanogrammus aeglefinus Ab.IgG4|Melanogrammus aeglefinus Ab.IgG4
C2734320|T201|COMP|56281-9|LNC|Hippoglossus hippoglossus Ab.IgG4|Hippoglossus hippoglossus Ab.IgG4
C2734322|T201|COMP|56282-7|LNC|Corylus avellana pollen Ab.IgG4|Corylus avellana pollen Ab.IgG4
C2734324|T201|COMP|56283-5|LNC|Corylus avellana Ab.IgG4|Corylus avellana Ab.IgG4
C2734326|T201|COMP|56284-3|LNC|Clupea harengus Ab.IgG4|Clupea harengus Ab.IgG4
C2734328|T201|COMP|56285-0|LNC|Honey Ab.IgG4|Honey Ab.IgG4
C2734330|T201|COMP|56286-8|LNC|Apis mellifera Ab.IgG4|Apis mellifera Ab.IgG4
C2734331|T201|COMP|56287-6|LNC|Cucumis melo spp Ab.IgG4|Cucumis melo spp Ab.IgG4
C2734333|T201|COMP|56288-4|LNC|Humulus lupus Ab.IgG4|Humulus lupus Ab.IgG4
C2734335|T201|COMP|56289-2|LNC|Armoracia rusticana Ab.IgG4|Armoracia rusticana Ab.IgG4
C2734337|T201|COMP|56290-0|LNC|House dust Greer Ab.IgG4|House dust Greer Ab.IgG4
C2734341|T201|COMP|56292-6|LNC|Insulin human Ab.IgG4|Insulin human Ab.IgG4
C2734343|T201|COMP|56293-4|LNC|Cupressus sempervirens Ab.IgG4|Cupressus sempervirens Ab.IgG4
C2734345|T201|COMP|56294-2|LNC|Sorghum halepense Ab.IgG4|Sorghum halepense Ab.IgG4
C2734347|T201|COMP|56295-9|LNC|Karaya gum Ab.IgG4|Karaya gum Ab.IgG4
C2734349|T201|COMP|56296-7|LNC|Poa pratensis Ab.IgG4|Poa pratensis Ab.IgG4
C2734351|T201|COMP|56297-5|LNC|Bean kidney red Ab.IgG4|Bean kidney red Ab.IgG4
C2734353|T201|COMP|56298-3|LNC|Actinidia chinensis Ab.IgG4|Actinidia chinensis Ab.IgG4
C2734355|T201|COMP|56299-1|LNC|Kochia scoparia Ab.IgG4|Kochia scoparia Ab.IgG4
C2734357|T201|COMP|56300-7|LNC|Lepidoglyphus destructor Ab.IgG4|Lepidoglyphus destructor Ab.IgG4
C2734359|T201|COMP|56301-5|LNC|Lactalbumin alpha Ab.IgG4|Lactalbumin alpha Ab.IgG4
C2734360|T201|COMP|56302-3|LNC|Beta lactoglobulin Ab.IgG4|Beta lactoglobulin Ab.IgG4
C2734362|T201|COMP|56303-1|LNC|Chenopodium album Ab.IgG4|Chenopodium album Ab.IgG4
C2734364|T201|COMP|56304-9|LNC|Citrus limon Ab.IgG4|Citrus limon Ab.IgG4
C2734366|T201|COMP|56305-6|LNC|Atriplex lentiformis Ab.IgG4|Atriplex lentiformis Ab.IgG4
C2734368|T201|COMP|56306-4|LNC|Lens esculenta Ab.IgG4|Lens esculenta Ab.IgG4
C2734370|T201|COMP|56318-9|LNC|Alopercurus pratensis Ab.IgG4|Alopercurus pratensis Ab.IgG4
C2734372|T201|COMP|56319-7|LNC|Melaleuca leucadendron Ab.IgG4|Melaleuca leucadendron Ab.IgG4
C2734374|T201|COMP|56320-5|LNC|Prosopis juliflora Ab.IgG4|Prosopis juliflora Ab.IgG4
C2734376|T201|COMP|56321-3|LNC|Panicum milliaceum Ab.IgG4|Panicum milliaceum Ab.IgG4
C2734378|T201|COMP|56322-1|LNC|Aedes communis Ab.IgG4|Aedes communis Ab.IgG4
C2734380|T201|COMP|56323-9|LNC|Juniperus sabinoides Ab.IgG4|Juniperus sabinoides Ab.IgG4
C2734382|T201|COMP|56324-7|LNC|Mucor racemosus Ab.IgG4|Mucor racemosus Ab.IgG4
C2734384|T201|COMP|56325-4|LNC|Artemisia vulgaris Ab.IgG4|Artemisia vulgaris Ab.IgG4
C2734386|T201|COMP|56326-2|LNC|Agaricus hortensis Ab.IgG4|Agaricus hortensis Ab.IgG4
C2734388|T201|COMP|56327-0|LNC|Mytilus edulis Ab.IgG4|Mytilus edulis Ab.IgG4
C2734390|T201|COMP|56328-8|LNC|Mustard Ab.IgG4|Mustard Ab.IgG4
C2734392|T201|COMP|56329-6|LNC|Prunus persica var nucipersica Ab.IgG4|Prunus persica var nucipersica Ab.IgG4
C2734394|T201|COMP|56330-4|LNC|Urtica dioica Ab.IgG4|Urtica dioica Ab.IgG4
C2734398|T201|COMP|56332-0|LNC|Nutmeg Ab.IgG4|Nutmeg Ab.IgG4
C2734400|T201|COMP|56333-8|LNC|Avena sativa Ab.IgG4|Avena sativa Ab.IgG4
C2734402|T201|COMP|56334-6|LNC|Avena sativa cultivated Ab.IgG4|Avena sativa cultivated Ab.IgG4
C2734404|T201|COMP|56335-3|LNC|Abelmoschus esculentus Ab.IgG4|Abelmoschus esculentus Ab.IgG4
C2734406|T201|COMP|56336-1|LNC|Olea europaea pollen Ab.IgG4|Olea europaea pollen Ab.IgG4
C2734408|T201|COMP|56337-9|LNC|Allium cepa Ab.IgG4|Allium cepa Ab.IgG4
C2734410|T201|COMP|56338-7|LNC|Citrus sinensis Ab.IgG4|Citrus sinensis Ab.IgG4
C2734412|T201|COMP|56339-5|LNC|Dactylis glomerata Ab.IgG4|Dactylis glomerata Ab.IgG4
C2734414|T201|COMP|56340-3|LNC|Origanum vulgare Ab.IgG4|Origanum vulgare Ab.IgG4
C2734416|T201|COMP|56341-1|LNC|Chrysanthemum leucanthemum Ab.IgG4|Chrysanthemum leucanthemum Ab.IgG4
C2734418|T201|COMP|56342-9|LNC|Ostrea edulis Ab.IgG4|Ostrea edulis Ab.IgG4
C2734420|T201|COMP|56343-7|LNC|Carica papaya Ab.IgG4|Carica papaya Ab.IgG4
C2734422|T201|COMP|56344-5|LNC|Polistes spp Ab.IgG4|Polistes spp Ab.IgG4
C2734424|T201|COMP|56345-2|LNC|Capsicum annuum Ab.IgG4|Capsicum annuum Ab.IgG4
C2734426|T201|COMP|56346-0|LNC|Cheese parmesan Ab.IgG4|Cheese parmesan Ab.IgG4
C2734428|T201|COMP|56347-8|LNC|Parrot feather Ab.IgG4|Parrot feather Ab.IgG4
C2734430|T201|COMP|56348-6|LNC|Petroselinum crispum Ab.IgG4|Petroselinum crispum Ab.IgG4
C2734432|T201|COMP|56349-4|LNC|Pastinaca sativa Ab.IgG4|Pastinaca sativa Ab.IgG4
C2734434|T201|COMP|56350-2|LNC|Prunus persica Ab.IgG4|Prunus persica Ab.IgG4
C2734436|T201|COMP|56351-0|LNC|Arachis hypogaea Ab.IgG4|Arachis hypogaea Ab.IgG4
C2734438|T201|COMP|56352-8|LNC|Pyrus communis Ab.IgG4|Pyrus communis Ab.IgG4
C2734440|T201|COMP|56353-6|LNC|Carya illinoinensis nut Ab.IgG4|Carya illinoinensis nut Ab.IgG4
C2734442|T201|COMP|56354-4|LNC|Carya illinoinensis tree Ab.IgG4|Carya illinoinensis tree Ab.IgG4
C2734444|T201|COMP|56355-1|LNC|Penicillium notatum Ab.IgG4|Penicillium notatum Ab.IgG4
C2734446|T201|COMP|56356-9|LNC|Perca spp Ab.IgG4|Perca spp Ab.IgG4
C2734448|T201|COMP|56365-0|LNC|Syagrus romanzoffianum Ab.IgG4|Syagrus romanzoffianum Ab.IgG4
C2734450|T201|COMP|56366-8|LNC|Rabbit Ab.IgG4|Rabbit Ab.IgG4
C2734452|T201|COMP|56367-6|LNC|Rabbit epithelium Ab.IgG4|Rabbit epithelium Ab.IgG4
C2734454|T201|COMP|56368-4|LNC|Raphanus sativus Ab.IgG4|Raphanus sativus Ab.IgG4
C2734456|T201|COMP|56369-2|LNC|Franseria acanthicarpa Ab.IgG4|Franseria acanthicarpa Ab.IgG4
C2734458|T201|COMP|56370-0|LNC|Ambrosia trifida Ab.IgG4|Ambrosia trifida Ab.IgG4
C2734460|T201|COMP|56371-8|LNC|Ambrosia elatior Ab.IgG4|Ambrosia elatior Ab.IgG4
C2734462|T201|COMP|56372-6|LNC|Ambrosia psilostachya Ab.IgG4|Ambrosia psilostachya Ab.IgG4
C2734464|T201|COMP|56373-4|LNC|Rubus idaeus Ab.IgG4|Rubus idaeus Ab.IgG4
C2734466|T201|COMP|56374-2|LNC|Rat epithelium Ab.IgG4|Rat epithelium Ab.IgG4
C2734468|T201|COMP|56375-9|LNC|Beet red Ab.IgG4|Beet red Ab.IgG4
C2734470|T201|COMP|56376-7|LNC|Snapper red Ab.IgG4|Snapper red Ab.IgG4
C2734472|T201|COMP|56377-5|LNC|Agrostis stolonifera Ab.IgG4|Agrostis stolonifera Ab.IgG4
C2734474|T201|COMP|56378-3|LNC|Rheum spp Ab.IgG4|Rheum spp Ab.IgG4
C2734476|T201|COMP|56379-1|LNC|Oryza sativa Ab.IgG4|Oryza sativa Ab.IgG4
C2734477|T201|COMP|56380-9|LNC|Salsola kali Ab.IgG4|Salsola kali Ab.IgG4
C2734479|T201|COMP|56381-7|LNC|Secale cereale pollen Ab.IgG4|Secale cereale pollen Ab.IgG4
C2734481|T201|COMP|56382-5|LNC|Carthamus tinctorius Ab.IgG4|Carthamus tinctorius Ab.IgG4
C2734483|T201|COMP|56400-5|LNC|Citrus reticulata Ab.IgG4|Citrus reticulata Ab.IgG4
C2734485|T201|COMP|56401-3|LNC|Camellia sinensis Ab.IgG4|Camellia sinensis Ab.IgG4
C2734487|T201|COMP|56402-1|LNC|Thymus vulgaris Ab.IgG4|Thymus vulgaris Ab.IgG4
C2734489|T201|COMP|56403-9|LNC|Phleum pratense Ab.IgG4|Phleum pratense Ab.IgG4
C2734490|T201|COMP|56404-7|LNC|Nicotiana tabacum Ab.IgG4|Nicotiana tabacum Ab.IgG4
C2734492|T201|COMP|56405-4|LNC|Lycopersicon lycopersicum Ab.IgG4|Lycopersicon lycopersicum Ab.IgG4
C2734494|T201|COMP|56406-2|LNC|Trichoderma viride Ab.IgG4|Trichoderma viride Ab.IgG4
C2734496|T201|COMP|56407-0|LNC|Oncorhynchus mykiss Ab.IgG4|Oncorhynchus mykiss Ab.IgG4
C2734498|T201|COMP|56408-8|LNC|Thunnus albacares Ab.IgG4|Thunnus albacares Ab.IgG4
C2734500|T201|COMP|56409-6|LNC|Turkey Ab.IgG4|Turkey Ab.IgG4
C2734502|T201|COMP|56410-4|LNC|Vanilla planifolia Ab.IgG4|Vanilla planifolia Ab.IgG4
C2734504|T201|COMP|56411-2|LNC|Holcus lanatus Ab.IgG4|Holcus lanatus Ab.IgG4
C2734506|T201|COMP|56412-0|LNC|Venison Ab.IgG4|Venison Ab.IgG4
C2734508|T201|COMP|56429-4|LNC|Solanum tuberosum Ab.IgG4|Solanum tuberosum Ab.IgG4
C2734510|T201|COMP|56430-2|LNC|Whitefish Ab.IgG4|Whitefish Ab.IgG4
C2734512|T201|COMP|56431-0|LNC|Wine Vinegar Ab.IgG4|Wine Vinegar Ab.IgG4
C2734514|T201|COMP|56432-8|LNC|Artemisia absinthium Ab.IgG4|Artemisia absinthium Ab.IgG4
C2734516|T201|COMP|56433-6|LNC|Dolichovespula arenaria Ab.IgG4|Dolichovespula arenaria Ab.IgG4
C2734517|T201|COMP|56434-4|LNC|Vespula spp Ab.IgG4|Vespula spp Ab.IgG4
C2734518|T201|COMP|56435-1|LNC|Yogurt Ab.IgG4|Yogurt Ab.IgG4
C2734520|T201|COMP|56436-9|LNC|Squash zucchini Ab.IgG4|Squash zucchini Ab.IgG4
C2734522|T201|COMP|56437-7|LNC|Chicken feather Ab.IgG4|Chicken feather Ab.IgG4
C2734524|T201|COMP|56438-5|LNC|Beef Ab.IgG4|Beef Ab.IgG4
C2734526|T201|COMP|56439-3|LNC|Scomber japonicus Ab.IgG4|Scomber japonicus Ab.IgG4
C2734528|T201|COMP|56440-1|LNC|Syzygium aromaticum Ab.IgG4|Syzygium aromaticum Ab.IgG4
C2734530|T201|COMP|56441-9|LNC|Latex Ab.IgG4|Latex Ab.IgG4
C2734532|T201|COMP|56442-7|LNC|Pork Ab.IgG4|Pork Ab.IgG4
C2734534|T201|COMP|56443-5|LNC|Secale cereale Ab.IgG4|Secale cereale Ab.IgG4
C2734543|T201|COMP|56448-4|LNC|Chloride|Chloride
C2734544|T201|COMP|56449-2|LNC|Saccharomyces cerevisiae Ab.IgG4|Saccharomyces cerevisiae Ab.IgG4
C2734546|T201|COMP|56450-0|LNC|Piper nigrum Ab.IgG4|Piper nigrum Ab.IgG4
C2734548|T201|COMP|56451-8|LNC|Chymopapain Ab.IgG4|Chymopapain Ab.IgG4
C2734550|T201|COMP|56452-6|LNC|Cottonseed Ab.IgG4|Cottonseed Ab.IgG4
C2734552|T201|COMP|56465-8|LNC|Distichlis spicata Ab.IgG4|Distichlis spicata Ab.IgG4
C2734554|T201|COMP|56466-6|LNC|Xiphias gladius Ab.IgG4|Xiphias gladius Ab.IgG4
C2734556|T201|COMP|56467-4|LNC|Tabanus spp Ab.IgG4|Tabanus spp Ab.IgG4
C2734558|T201|COMP|56468-2|LNC|Cucurbita pepo Ab.IgG4|Cucurbita pepo Ab.IgG4
C2734560|T201|COMP|56469-0|LNC|Cardiac heart disease risk|Cardiac heart disease risk
C2734562|T201|COMP|56470-8|LNC|Blasts|Blasts
C2734565|T201|COMP|56472-4|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C2734566|T201|COMP|56473-2|LNC|Metamyelocytes|Metamyelocytes
C2734567|T201|COMP|56474-0|LNC|Salmonella sp identified|Salmonella sp identified
C2734568|T201|COMP|56475-7|LNC|Salmonella sp antigenic formula|Salmonella sp antigenic formula
C2734570|T201|COMP|56476-5|LNC|Hemoglobin S/Hemoglobin.total|Hemoglobin S/Hemoglobin.total
C2734571|T201|COMP|56477-3|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C2734572|T201|COMP|56478-1|LNC|Ethanol|Ethanol
C2734573|T201|COMP|56479-9|LNC|Superoxide dismutase|Superoxide dismutase
C2734574|T201|COMP|56480-7|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C2734575|T201|COMP|56481-5|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C2734576|T201|COMP|56482-3|LNC|Insulin^baseline|Insulin^baseline
C2734577|T201|COMP|56483-1|LNC|Porphobilinogen|Porphobilinogen
C2734578|T201|COMP|56484-9|LNC|Uroporphyrin|Uroporphyrin
C2734579|T201|COMP|56485-6|LNC|Taenia solium Ab.IgG|Taenia solium Ab.IgG
C2734580|T201|COMP|56486-4|LNC|Taenia solium Ab.IgG|Taenia solium Ab.IgG
C2734581|T201|COMP|56487-2|LNC|Androsterone|Androsterone
C2734582|T201|COMP|56488-0|LNC|Etiocholanolone|Etiocholanolone
C2734583|T201|COMP|56489-8|LNC|Acidity.titratable|Acidity.titratable
C2734584|T201|COMP|56490-6|LNC|Hemoglobin.gastrointestinal.lower^2nd specimen|Hemoglobin.gastrointestinal.lower^2nd specimen
C2734585|T201|COMP|56491-4|LNC|Hemoglobin.gastrointestinal.lower^3rd specimen|Hemoglobin.gastrointestinal.lower^3rd specimen
C2734586|T201|COMP|56492-2|LNC|Insulin^6M post XXX challenge|Insulin^6M post XXX challenge
C2734587|T201|COMP|56493-0|LNC|Lutropin^10M post XXX challenge|Lutropin^10M post XXX challenge
C2734588|T201|COMP|56494-8|LNC|Lutropin^2H post XXX challenge|Lutropin^2H post XXX challenge
C2734589|T201|COMP|56495-5|LNC|Lutropin^3H post XXX challenge|Lutropin^3H post XXX challenge
C2734590|T201|COMP|56496-3|LNC|Prolactin^2H post XXX challenge|Prolactin^2H post XXX challenge
C2734591|T201|COMP|56497-1|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C2734592|T201|COMP|56498-9|LNC|Androstenedione^30M post XXX challenge|Androstenedione^30M post XXX challenge
C2734593|T201|COMP|56499-7|LNC|Somatotropin^45M post XXX challenge|Somatotropin^45M post XXX challenge
C2734594|T201|COMP|56500-2|LNC|Somatotropin^3H post XXX challenge|Somatotropin^3H post XXX challenge
C2734595|T201|COMP|56501-0|LNC|Somatotropin^6H post XXX challenge|Somatotropin^6H post XXX challenge
C2734596|T201|COMP|56502-8|LNC|Somatotropin^7H post XXX challenge|Somatotropin^7H post XXX challenge
C2734597|T201|COMP|56503-6|LNC|Somatotropin^8H post XXX challenge|Somatotropin^8H post XXX challenge
C2734598|T201|COMP|56504-4|LNC|Corticotropin^15M post XXX challenge|Corticotropin^15M post XXX challenge
C2734599|T201|COMP|56505-1|LNC|Corticotropin^45M post XXX challenge|Corticotropin^45M post XXX challenge
C2734600|T201|COMP|56506-9|LNC|Corticotropin^2H post XXX challenge|Corticotropin^2H post XXX challenge
C2734603|T201|COMP|56510-1|LNC|Dehydroepiandrosterone^1H post XXX challenge|Dehydroepiandrosterone^1H post XXX challenge
C2734604|T201|COMP|56511-9|LNC|Calcitonin^2M post XXX challenge|Calcitonin^2M post XXX challenge
C2734605|T201|COMP|56512-7|LNC|Porphyrins|Porphyrins
C2734606|T201|COMP|56513-5|LNC|Hepatitis E virus Ab.IgG|Hepatitis E virus Ab.IgG
C2734607|T201|COMP|56514-3|LNC|Legionella pneumophila Ab.IgG|Legionella pneumophila Ab.IgG
C2734608|T201|COMP|56515-0|LNC|Plasmodium falciparum Ab.IgG|Plasmodium falciparum Ab.IgG
C2734609|T201|COMP|56516-8|LNC|C peptide^6M post XXX challenge|C peptide^6M post XXX challenge
C2734610|T201|COMP|56517-6|LNC|11-Deoxycortisol^2H post XXX challenge|11-Deoxycortisol^2H post XXX challenge
C2734611|T201|COMP|56518-4|LNC|11-Deoxycortisol^15M post XXX challenge|11-Deoxycortisol^15M post XXX challenge
C2734612|T201|COMP|56519-2|LNC|11-Deoxycortisol^30M post XXX challenge|11-Deoxycortisol^30M post XXX challenge
C2734613|T201|COMP|56520-0|LNC|11-Deoxycortisol^45M post XXX challenge|11-Deoxycortisol^45M post XXX challenge
C2734614|T201|COMP|56521-8|LNC|11-Deoxycortisol^1.5H post XXX challenge|11-Deoxycortisol^1.5H post XXX challenge
C2734617|T201|COMP|56525-9|LNC|5-Hydroxytryptophan|5-Hydroxytryptophan
C2734618|T201|COMP|56526-7|LNC|Somatotropin^30M post exercise|Somatotropin^30M post exercise
C2734619|T201|COMP|56527-5|LNC|Vasopressin^1H post XXX challenge|Vasopressin^1H post XXX challenge
C2734620|T201|COMP|56528-3|LNC|Androstenedione^20M post XXX challenge|Androstenedione^20M post XXX challenge
C2734621|T201|COMP|56529-1|LNC|Ma+Ta Ab|Ma+Ta Ab
C2734622|T201|COMP|56530-9|LNC|CV2 Ab|CV2 Ab
C2734623|T201|COMP|56531-7|LNC|Amphiphysin Ab|Amphiphysin Ab
C2734624|T201|COMP|56532-5|LNC|Asialoglycoprotein receptor Ab|Asialoglycoprotein receptor Ab
C2734625|T201|COMP|56533-3|LNC|Insulin Ab.IgG|Insulin Ab.IgG
C2734627|T201|COMP|56534-1|LNC|Calcitonin^15M post XXX challenge|Calcitonin^15M post XXX challenge
C2734628|T201|COMP|56535-8|LNC|8-Dehydrocholesterol|8-Dehydrocholesterol
C2734629|T201|COMP|56536-6|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C2734630|T201|COMP|56537-4|LNC|Tissue transglutaminase Ab.IgG|Tissue transglutaminase Ab.IgG
C2734631|T201|COMP|56538-2|LNC|Beta 2 glycoprotein 1 Ab|Beta 2 glycoprotein 1 Ab
C2734632|T201|COMP|56539-0|LNC|Intrinsic factor Ab|Intrinsic factor Ab
C2734633|T201|COMP|56540-8|LNC|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C2734634|T201|COMP|56541-6|LNC|Ganglioside GD1b Ab.IgG|Ganglioside GD1b Ab.IgG
C2734635|T201|COMP|56542-4|LNC|Ganglioside GD1b Ab.IgM|Ganglioside GD1b Ab.IgM
C2734636|T201|COMP|56543-2|LNC|Ganglioside GM2 Ab.IgG|Ganglioside GM2 Ab.IgG
C2734637|T201|COMP|56544-0|LNC|Ganglioside GM2 Ab.IgM|Ganglioside GM2 Ab.IgM
C2734638|T201|COMP|56545-7|LNC|Ganglioside GQ1b Ab.IgM|Ganglioside GQ1b Ab.IgM
C2734639|T201|COMP|56546-5|LNC|Insulin Ab|Insulin Ab
C2734640|T201|COMP|56547-3|LNC|Tubular basement membrane Ab.IgG|Tubular basement membrane Ab.IgG
C2734641|T201|COMP|56548-1|LNC|U1 small nuclear ribonucleoprotein Ab.IgG|U1 small nuclear ribonucleoprotein Ab.IgG
C2734642|T201|COMP|56549-9|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C2734643|T201|COMP|56550-7|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C2734644|T201|COMP|56551-5|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C2734645|T201|COMP|56552-3|LNC|Dehydroepiandrosterone sulfate^baseline|Dehydroepiandrosterone sulfate^baseline
C2734646|T201|COMP|56553-1|LNC|Albumin|Albumin
C2734647|T201|COMP|56554-9|LNC|Porphyrins|Porphyrins
C2734648|T201|COMP|56555-6|LNC|11-Deoxycorticosterone^baseline|11-Deoxycorticosterone^baseline
C2734649|T201|COMP|56556-4|LNC|11-Deoxycorticosterone^30M post XXX challenge|11-Deoxycorticosterone^30M post XXX challenge
C2734650|T201|COMP|56557-2|LNC|Renin^10M post XXX challenge|Renin^10M post XXX challenge
C2734651|T201|COMP|56558-0|LNC|Aldosterone^10M post XXX challenge|Aldosterone^10M post XXX challenge
C2734652|T201|COMP|56559-8|LNC|Norepinephrine^pre/post XXX challenge|Norepinephrine^pre/post XXX challenge
C2734653|T201|COMP|56560-6|LNC|Somatotropin^4.5H post XXX challenge|Somatotropin^4.5H post XXX challenge
C2734654|T201|COMP|56561-4|LNC|Somatotropin^5.5H post XXX challenge|Somatotropin^5.5H post XXX challenge
C2734655|T201|COMP|56562-2|LNC|Somatotropin^6.5H post XXX challenge|Somatotropin^6.5H post XXX challenge
C2734656|T201|COMP|56563-0|LNC|Somatotropin^7.5H post XXX challenge|Somatotropin^7.5H post XXX challenge
C2734657|T201|COMP|56564-8|LNC|Somatotropin^8H post XXX challenge|Somatotropin^8H post XXX challenge
C2734658|T201|COMP|56565-5|LNC|Somatotropin^9H post XXX challenge|Somatotropin^9H post XXX challenge
C2734659|T201|COMP|56566-3|LNC|Somatotropin^9.5H post XXX challenge|Somatotropin^9.5H post XXX challenge
C2734660|T201|COMP|56567-1|LNC|Somatotropin^10H post XXX challenge|Somatotropin^10H post XXX challenge
C2734661|T201|COMP|56568-9|LNC|Somatotropin^10.5H post XXX challenge|Somatotropin^10.5H post XXX challenge
C2734662|T201|COMP|56569-7|LNC|Somatotropin^11H post XXX challenge|Somatotropin^11H post XXX challenge
C2734663|T201|COMP|56570-5|LNC|Somatotropin^11.5H post XXX challenge|Somatotropin^11.5H post XXX challenge
C2734664|T201|COMP|56571-3|LNC|Somatotropin^post exercise|Somatotropin^post exercise
C2734665|T201|COMP|56572-1|LNC|Somatotropin^20H post XXX challenge|Somatotropin^20H post XXX challenge
C2734666|T201|COMP|56573-9|LNC|Renin^30M post XXX challenge|Renin^30M post XXX challenge
C2734667|T201|COMP|56574-7|LNC|Renin^1H post XXX challenge|Renin^1H post XXX challenge
C2734668|T201|COMP|56575-4|LNC|17-Hydroxyprogesterone^15M post XXX challenge|17-Hydroxyprogesterone^15M post XXX challenge
C2734669|T201|COMP|56892-3|LNC|Cells.CD13+HLA-DR+/100 cells|Cells.CD13+HLA-DR+/100 cells
C2734692|T201|COMP|57018-4|LNC|Hydrogen/Expired gas^3H post dose lactulose|Hydrogen/Expired gas^3H post dose lactulose
C2734693|T201|COMP|57019-2|LNC|Urinalysis dipstick W Reflex Culture panel|Urinalysis dipstick W Reflex Culture panel
C2734695|T201|COMP|57020-0|LNC|Urinalysis dipstick W Reflex Microscopic panel|Urinalysis dipstick W Reflex Microscopic panel
C2734697|T201|COMP|57021-8|LNC|CBC W Auto Differential panel|CBC W Auto Differential panel
C2734699|T201|COMP|57022-6|LNC|CBC W Reflex Manual Differential panel|CBC W Reflex Manual Differential panel
C2734701|T201|COMP|57023-4|LNC|Auto Differential panel|Auto Differential panel
C2734711|T201|COMP|57028-3|LNC|Iron|Iron
C2734712|T201|COMP|57029-1|LNC|Fetal chromosome 13+18+21+X+Y aneuploidy|Fetal chromosome 13+18+21+X+Y aneuploidy
C2734714|T201|COMP|57030-9|LNC|Chromosome 13+18+21+X+Y aneuploidy|Chromosome 13+18+21+X+Y aneuploidy
C2734715|T201|COMP|57031-7|LNC|Herpesviruses 6 DNA panel|Herpesviruses 6 DNA panel
C2734717|T201|COMP|57032-5|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C2734718|T201|COMP|57033-3|LNC|Alternaria alternata Ab|Alternaria alternata Ab
C2734719|T201|COMP|57034-1|LNC|Penicillium sp Ab|Penicillium sp Ab
C2734720|T201|COMP|57035-8|LNC|Cow milk Ab|Cow milk Ab
C2734721|T201|COMP|57036-6|LNC|Phadiatop inhalant allergen Ab.IgE|Phadiatop inhalant allergen Ab.IgE
C2734723|T201|COMP|57037-4|LNC|Chromosome 13+18+21+X+Y aneuploidy|Chromosome 13+18+21+X+Y aneuploidy
C2734742|T201|COMP|56576-2|LNC|17-Hydroxyprogesterone^45M post XXX challenge|17-Hydroxyprogesterone^45M post XXX challenge
C2734743|T201|COMP|56577-0|LNC|Renin^1.5H post XXX challenge|Renin^1.5H post XXX challenge
C2734744|T201|COMP|56578-8|LNC|Aldosterone^1.5H post XXX challenge|Aldosterone^1.5H post XXX challenge
C2734745|T201|COMP|56579-6|LNC|Aldosterone^20M post XXX challenge|Aldosterone^20M post XXX challenge
C2734746|T201|COMP|56580-4|LNC|Renin^20M post XXX challenge|Renin^20M post XXX challenge
C2734747|T201|COMP|56581-2|LNC|Insulin^12M post XXX challenge|Insulin^12M post XXX challenge
C2734748|T201|COMP|56582-0|LNC|C peptide^10M post XXX challenge|C peptide^10M post XXX challenge
C2734749|T201|COMP|56583-8|LNC|C peptide^45M post XXX challenge|C peptide^45M post XXX challenge
C2734750|T201|COMP|56584-6|LNC|C peptide^12M post XXX challenge|C peptide^12M post XXX challenge
C2734751|T201|COMP|56585-3|LNC|Cortisol^45M post XXX challenge|Cortisol^45M post XXX challenge
C2734752|T201|COMP|56586-1|LNC|Dehydroepiandrosterone^15M post XXX challenge|Dehydroepiandrosterone^15M post XXX challenge
C2734753|T201|COMP|56587-9|LNC|Dehydroepiandrosterone^30M post XXX challenge|Dehydroepiandrosterone^30M post XXX challenge
C2734755|T201|COMP|56589-5|LNC|Dehydroepiandrosterone^1.5H post XXX challenge|Dehydroepiandrosterone^1.5H post XXX challenge
C2734756|T201|COMP|56590-3|LNC|Dehydroepiandrosterone^2H post XXX challenge|Dehydroepiandrosterone^2H post XXX challenge
C2734758|T201|COMP|56592-9|LNC|Follitropin^10M post XXX challenge|Follitropin^10M post XXX challenge
C2734759|T201|COMP|56593-7|LNC|Follitropin^3H post XXX challenge|Follitropin^3H post XXX challenge
C2734762|T201|COMP|56608-3|LNC|11-Deoxycorticosterone^15M post XXX challenge|11-Deoxycorticosterone^15M post XXX challenge
C2734763|T201|COMP|56609-1|LNC|11-Deoxycorticosterone^20M post XXX challenge|11-Deoxycorticosterone^20M post XXX challenge
C2734764|T201|COMP|56610-9|LNC|11-Deoxycorticosterone^40M post XXX challenge|11-Deoxycorticosterone^40M post XXX challenge
C2734765|T201|COMP|56611-7|LNC|11-Deoxycorticosterone^1.5H post XXX challenge|11-Deoxycorticosterone^1.5H post XXX challenge
C2734766|T201|COMP|56612-5|LNC|11-Deoxycorticosterone^2H post XXX challenge|11-Deoxycorticosterone^2H post XXX challenge
C2734767|T201|COMP|56613-3|LNC|11-Deoxycorticosterone^2.5H post XXX challenge|11-Deoxycorticosterone^2.5H post XXX challenge
C2734768|T201|COMP|56614-1|LNC|17-Hydroxyprogesterone^10M post XXX challenge|17-Hydroxyprogesterone^10M post XXX challenge
C2734769|T201|COMP|56615-8|LNC|17-Hydroxyprogesterone^20M post XXX challenge|17-Hydroxyprogesterone^20M post XXX challenge
C2734770|T201|COMP|56616-6|LNC|17-Hydroxyprogesterone^1.5H post XXX challenge|17-Hydroxyprogesterone^1.5H post XXX challenge
C2734771|T201|COMP|56617-4|LNC|17-Hydroxyprogesterone^2H post XXX challenge|17-Hydroxyprogesterone^2H post XXX challenge
C2734774|T201|COMP|56620-8|LNC|Elastase Ab|Elastase Ab
C2734775|T201|COMP|56621-6|LNC|Coxsackievirus A9 Ab.IgG|Coxsackievirus A9 Ab.IgG
C2734777|T201|COMP|56622-4|LNC|Echovirus Ab.IgG|Echovirus Ab.IgG
C2734778|T201|COMP|56623-2|LNC|Echovirus Ab.IgM|Echovirus Ab.IgM
C2734779|T201|COMP|56624-0|LNC|Fructose|Fructose
C2734780|T201|COMP|56625-7|LNC|Methylene chloride|Methylene chloride
C2734781|T201|COMP|56626-5|LNC|Tetrachloroethylene|Tetrachloroethylene
C2734782|T201|COMP|56627-3|LNC|Procollagen type III|Procollagen type III
C2734783|T201|COMP|56628-1|LNC|Amikacin|Amikacin
C2734784|T201|COMP|56629-9|LNC|Myelin Ab|Myelin Ab
C2734785|T201|COMP|56630-7|LNC|Brucella sp Ab.IgG|Brucella sp Ab.IgG
C2734786|T201|COMP|56631-5|LNC|Brucella sp Ab.IgM|Brucella sp Ab.IgM
C2734787|T201|COMP|56632-3|LNC|Mitochondria M2 Ab.IgG|Mitochondria M2 Ab.IgG
C2734788|T201|COMP|56633-1|LNC|Myocardium Ab.IgG|Myocardium Ab.IgG
C2734789|T201|COMP|56634-9|LNC|Nuclear Ab.IgG|Nuclear Ab.IgG
C2734790|T201|COMP|56635-6|LNC|Thyroglobulin Ab.IgG|Thyroglobulin Ab.IgG
C2734792|T201|COMP|56636-4|LNC|Bordetella parapertussis Ab.IgM|Bordetella parapertussis Ab.IgM
C2734794|T201|COMP|56637-2|LNC|Mi-2 Ab|Mi-2 Ab
C2734795|T201|COMP|56638-0|LNC|Rheumatoid arthritis nuclear Ab|Rheumatoid arthritis nuclear Ab
C2734796|T201|COMP|56639-8|LNC|Methyl ethyl ketone|Methyl ethyl ketone
C2734797|T201|COMP|56640-6|LNC|Aspartate/Creatinine|Aspartate/Creatinine
C2734798|T201|COMP|56641-4|LNC|Threonine/Creatinine|Threonine/Creatinine
C2734799|T201|COMP|56642-2|LNC|Serine/Creatinine|Serine/Creatinine
C2734800|T201|COMP|56643-0|LNC|Asparagine/Creatinine|Asparagine/Creatinine
C2734801|T201|COMP|56644-8|LNC|Glutamate/Creatinine|Glutamate/Creatinine
C2734802|T201|COMP|56645-5|LNC|Vanillylmandelate/Creatine|Vanillylmandelate/Creatine
C2734803|T201|COMP|56646-3|LNC|Trichloroacetate/Creatinine|Trichloroacetate/Creatinine
C2734804|T201|COMP|56647-1|LNC|Phenol/Creatinine|Phenol/Creatinine
C2734805|T201|COMP|56648-9|LNC|Phenylglyoxylate/Creatinine|Phenylglyoxylate/Creatinine
C2734806|T201|COMP|56649-7|LNC|Hippurate/Creatinine|Hippurate/Creatinine
C2734807|T201|COMP|56655-4|LNC|Bromide/Creatinine|Bromide/Creatinine
C2734809|T201|COMP|56657-0|LNC|Tetrahydrocortisone|Tetrahydrocortisone
C2734810|T201|COMP|56658-8|LNC|Delta aminolevulinate/Creatinine|Delta aminolevulinate/Creatinine
C2734811|T201|COMP|56659-6|LNC|Para aminophenol/Creatinine|Para aminophenol/Creatinine
C2734812|T201|COMP|56660-4|LNC|Methyl formamide/Creatinine|Methyl formamide/Creatinine
C2734814|T201|COMP|56661-2|LNC|Myelin basic protein|Myelin basic protein
C2734815|T201|COMP|56662-0|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C2734816|T201|COMP|56663-8|LNC|5-Hydroxytryptophan|5-Hydroxytryptophan
C2734817|T201|COMP|56664-6|LNC|Methylmalonate/Creatinine|Methylmalonate/Creatinine
C2734818|T201|COMP|56665-3|LNC|Taenia solium Ab.IgG|Taenia solium Ab.IgG
C2734819|T201|COMP|56666-1|LNC|1-Methylhistidine/Creatinine|1-Methylhistidine/Creatinine
C2734820|T201|COMP|56667-9|LNC|3-Methylhistidine/Creatinine|3-Methylhistidine/Creatinine
C2734821|T201|COMP|56668-7|LNC|Alpha aminoadipate/Creatinine|Alpha aminoadipate/Creatinine
C2734822|T201|COMP|56669-5|LNC|Carotene.alpha|Carotene.alpha
C2734823|T201|COMP|56670-3|LNC|Adrenal cortex Ab.IgG|Adrenal cortex Ab.IgG
C2734825|T201|COMP|56671-1|LNC|Alanine/Creatinine|Alanine/Creatinine
C2734826|T201|COMP|56672-9|LNC|Arginine/Creatinine|Arginine/Creatinine
C2734827|T201|COMP|56673-7|LNC|Beta aminoisobutyrate/Creatinine|Beta aminoisobutyrate/Creatinine
C2734828|T201|COMP|56674-5|LNC|Beta alanine/Creatinine|Beta alanine/Creatinine
C2734829|T201|COMP|56675-2|LNC|Carnosine/Creatinine|Carnosine/Creatinine
C2734830|T201|COMP|56676-0|LNC|Citrulline/Creatinine|Citrulline/Creatinine
C2734831|T201|COMP|56677-8|LNC|Cystine/Creatinine|Cystine/Creatinine
C2734832|T201|COMP|56678-6|LNC|Ethanolamine/Creatinine|Ethanolamine/Creatinine
C2734833|T201|COMP|56679-4|LNC|Gamma aminobutyrate/Creatinine|Gamma aminobutyrate/Creatinine
C2734834|T201|COMP|56680-2|LNC|Glutamine/Creatinine|Glutamine/Creatinine
C2734835|T201|COMP|56681-0|LNC|Glycine/Creatinine|Glycine/Creatinine
C2734836|T201|COMP|56682-8|LNC|Homocystine/Creatinine|Homocystine/Creatinine
C2734837|T201|COMP|56683-6|LNC|Histidine/Creatinine|Histidine/Creatinine
C2734838|T201|COMP|56684-4|LNC|Hydroxylysine/Creatinine|Hydroxylysine/Creatinine
C2734839|T201|COMP|56685-1|LNC|Hydroxyproline.free|Hydroxyproline.free
C2734840|T201|COMP|56686-9|LNC|Hydroxyproline.free/Creatinine|Hydroxyproline.free/Creatinine
C2734842|T201|COMP|56694-3|LNC|Chicken droppings Ab|Chicken droppings Ab
C2734844|T201|COMP|56695-0|LNC|Cephalexin Ab.IgE|Cephalexin Ab.IgE
C2734846|T201|COMP|56696-8|LNC|Cloxacillin Ab.IgE|Cloxacillin Ab.IgE
C2734848|T201|COMP|56697-6|LNC|Thiopental Ab.IgE|Thiopental Ab.IgE
C2734850|T201|COMP|56698-4|LNC|Atropine Ab.IgE|Atropine Ab.IgE
C2734852|T201|COMP|56699-2|LNC|Bupivacaine Ab.IgE|Bupivacaine Ab.IgE
C2734854|T201|COMP|56700-8|LNC|Naproxen Ab.IgE|Naproxen Ab.IgE
C2734856|T201|COMP|56701-6|LNC|Diclofenac Ab.IgE|Diclofenac Ab.IgE
C2734858|T201|COMP|56702-4|LNC|Ciprofloxacin Ab.IgE|Ciprofloxacin Ab.IgE
C2734860|T201|COMP|56703-2|LNC|Piroxicam Ab.IgE|Piroxicam Ab.IgE
C2734862|T201|COMP|56704-0|LNC|Droperidol Ab.IgE|Droperidol Ab.IgE
C2734864|T201|COMP|56705-7|LNC|Tobramycin Ab.IgE|Tobramycin Ab.IgE
C2734866|T201|COMP|56706-5|LNC|Doxycycline Ab.IgE|Doxycycline Ab.IgE
C2734868|T201|COMP|56707-3|LNC|Spiramycin Ab.IgE|Spiramycin Ab.IgE
C2734870|T201|COMP|56708-1|LNC|metroNIDAZOLE Ab.IgE|metroNIDAZOLE Ab.IgE
C2734872|T201|COMP|56709-9|LNC|Tartrazine Ab.IgE|Tartrazine Ab.IgE
C2734874|T201|COMP|56710-7|LNC|Clarithromycin Ab.IgE|Clarithromycin Ab.IgE
C2734876|T201|COMP|56711-5|LNC|Sodium benzoate Ab.IgE|Sodium benzoate Ab.IgE
C2734878|T201|COMP|56712-3|LNC|Dexamethasone Ab.IgE|Dexamethasone Ab.IgE
C2734880|T201|COMP|56713-1|LNC|Dog dander+Dog epithelium Ab.IgE|Dog dander+Dog epithelium Ab.IgE
C2734882|T201|COMP|56714-9|LNC|Bacteria identified|Bacteria identified
C2734883|T201|COMP|56715-6|LNC|Bacteria identified|Bacteria identified
C2734884|T201|COMP|56716-4|LNC|Nuclear pore protein gp210 Ab|Nuclear pore protein gp210 Ab
C2734885|T201|COMP|56717-2|LNC|Histone Ab|Histone Ab
C2734886|T201|COMP|56718-0|LNC|Islet cell 512 Ab|Islet cell 512 Ab
C2734887|T201|COMP|56719-8|LNC|Liver cytosol Ab|Liver cytosol Ab
C2734888|T201|COMP|56720-6|LNC|Ma+Ta Ab|Ma+Ta Ab
C2734889|T201|COMP|56721-4|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C2734890|T201|COMP|56722-2|LNC|Soluble liver Ab|Soluble liver Ab
C2734891|T201|COMP|56723-0|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C2734892|T201|COMP|56724-8|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C2734893|T201|COMP|56725-5|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C2734894|T201|COMP|56726-3|LNC|Lolium perenne recombinant profilin Ab.IgE|Lolium perenne recombinant profilin Ab.IgE
C2734896|T201|COMP|56727-1|LNC|Olea europaea recombinant (rOle e) 2 Ab.IgE|Olea europaea recombinant (rOle e) 2 Ab.IgE
C2734898|T201|COMP|56728-9|LNC|Thermoactinomyces vulgaris Ab.IgE|Thermoactinomyces vulgaris Ab.IgE
C2734900|T201|COMP|56729-7|LNC|Cladosporium cladosporioides Ab.IgE|Cladosporium cladosporioides Ab.IgE
C2734902|T201|COMP|56730-5|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C2734903|T201|COMP|56731-3|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C2734904|T201|COMP|56732-1|LNC|Ribosomal P Ab|Ribosomal P Ab
C2734905|T201|COMP|56886-5|LNC|Indirect antiglobulin test.XXX reagent|Indirect antiglobulin test.XXX reagent
C2734906|T201|COMP|56887-3|LNC|Myoglobin|Myoglobin
C2734907|T201|COMP|56888-1|LNC|HIV 1+2 Ab+HIV1 p24 Ag|HIV 1+2 Ab+HIV1 p24 Ag
C2734909|T201|COMP|56889-9|LNC|Cells.CD13+HLA-DR+/100 cells|Cells.CD13+HLA-DR+/100 cells
C2734910|T201|COMP|56890-7|LNC|Cells.CD13+HLA-DR+/100 cells|Cells.CD13+HLA-DR+/100 cells
C2734911|T201|COMP|56891-5|LNC|Cells.CD13+HLA-DR+/100 cells|Cells.CD13+HLA-DR+/100 cells
C2734914|T201|COMP|57382-4|LNC|Sodium|Sodium
C2734915|T201|COMP|57383-2|LNC|Tipranavir|Tipranavir
C2734916|T201|COMP|57385-7|LNC|Urea|Urea
C2734917|T201|COMP|57386-5|LNC|Urate|Urate
C2734918|T201|COMP|57387-3|LNC|Urate|Urate
C2734919|T201|COMP|57388-1|LNC|Urea|Urea
C2734920|T201|COMP|57389-9|LNC|Urea|Urea
C2734921|T201|COMP|57390-7|LNC|Specimen volume|Specimen volume
C2734922|T201|COMP|57391-5|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C2734923|T201|COMP|57392-3|LNC|Urea|Urea
C2734924|T201|COMP|57393-1|LNC|Cells.CD11a/100 cells|Cells.CD11a/100 cells
C2734925|T201|COMP|57394-9|LNC|Cells.CD19+CD34+/100 cells|Cells.CD19+CD34+/100 cells
C2734927|T201|COMP|57395-6|LNC|Cells.CD19+CD38+/100 cells|Cells.CD19+CD38+/100 cells
C2734928|T201|COMP|57396-4|LNC|Cells.CD19+CD56+/100 cells|Cells.CD19+CD56+/100 cells
C2734930|T201|COMP|57397-2|LNC|Cells.CD19+CD20+/100 cells|Cells.CD19+CD20+/100 cells
C2734932|T201|COMP|57667-8|LNC|Protein.monoclonal.beta|Protein.monoclonal.beta
C2734935|T201|COMP|57670-2|LNC|Brucella melitensis Ab.IgG|Brucella melitensis Ab.IgG
C2734937|T201|COMP|57671-0|LNC|Brucella melitensis Ab.IgM|Brucella melitensis Ab.IgM
C2734939|T201|COMP|57672-8|LNC|11-Deoxycortisol^2D post XXX challenge|11-Deoxycortisol^2D post XXX challenge
C2734940|T201|COMP|57673-6|LNC|Coxiella burnetii Ab.IgM^1st specimen|Coxiella burnetii Ab.IgM^1st specimen
C2734945|T201|COMP|57824-5|LNC|Cortisol.free^AM peak specimen|Cortisol.free^AM peak specimen
C2734946|T201|COMP|57825-2|LNC|Cortisol.free^PM trough specimen|Cortisol.free^PM trough specimen
C2734951|T201|COMP|56733-9|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C2734952|T201|COMP|56734-7|LNC|Centromere protein B Ab|Centromere protein B Ab
C2734953|T201|COMP|56735-4|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C2734954|T201|COMP|56736-2|LNC|Purkinje cells Ab|Purkinje cells Ab
C2734955|T201|COMP|56737-0|LNC|Ganglioside GM2 Ab.IgG|Ganglioside GM2 Ab.IgG
C2734956|T201|COMP|56738-8|LNC|Ganglioside GM2 Ab.IgM|Ganglioside GM2 Ab.IgM
C2734957|T201|COMP|56739-6|LNC|Ganglioside GD1b Ab.IgG|Ganglioside GD1b Ab.IgG
C2734958|T201|COMP|56740-4|LNC|Ganglioside GD1b Ab.IgM|Ganglioside GD1b Ab.IgM
C2734959|T201|COMP|56741-2|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C2734960|T201|COMP|56742-0|LNC|Ganglioside GQ1b Ab.IgM|Ganglioside GQ1b Ab.IgM
C2734961|T201|COMP|56743-8|LNC|Mi-2 Ab|Mi-2 Ab
C2734962|T201|COMP|56744-6|LNC|Pl-7 Ab|Pl-7 Ab
C2734963|T201|COMP|56745-3|LNC|Pl-12 Ab|Pl-12 Ab
C2734964|T201|COMP|56746-1|LNC|Allium ampeloprasum Ab.IgE|Allium ampeloprasum Ab.IgE
C2734966|T201|COMP|56747-9|LNC|Azithromycin Ab.IgE|Azithromycin Ab.IgE
C2734968|T201|COMP|56748-7|LNC|Norovirus RNA|Norovirus RNA
C2734970|T201|COMP|56749-5|LNC|Estradiol^30M post XXX challenge|Estradiol^30M post XXX challenge
C2734971|T201|COMP|56750-3|LNC|Estradiol^1H post XXX challenge|Estradiol^1H post XXX challenge
C2734972|T201|COMP|56751-1|LNC|Glucose^2.17H post XXX challenge|Glucose^2.17H post XXX challenge
C2734973|T201|COMP|56752-9|LNC|APOB gene+LDLR gene targeted mutation analysis|APOB gene+LDLR gene targeted mutation analysis
C2734975|T201|COMP|56753-7|LNC|PML Ab|PML Ab
C2734977|T201|COMP|56754-5|LNC|sp100 Ab|sp100 Ab
C2734978|T201|COMP|56755-2|LNC|Aldosterone^100M post XXX challenge|Aldosterone^100M post XXX challenge
C2734979|T201|COMP|56756-0|LNC|Aldosterone^70M post XXX challenge|Aldosterone^70M post XXX challenge
C2734980|T201|COMP|56757-8|LNC|Renin^100M post XXX challenge|Renin^100M post XXX challenge
C2734981|T201|COMP|56758-6|LNC|Renin^70M post XXX challenge|Renin^70M post XXX challenge
C2734982|T201|COMP|56759-4|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2734983|T201|COMP|56760-2|LNC|Liver kidney microsomal Ab|Liver kidney microsomal Ab
C2734984|T201|COMP|56761-0|LNC|Saccharomyces cerevisiae Ab|Saccharomyces cerevisiae Ab
C2734985|T201|COMP|56762-8|LNC|Protein fractions.oligoclonal bands.IgG|Protein fractions.oligoclonal bands.IgG
C2734987|T201|COMP|56763-6|LNC|Protein fractions.oligoclonal bands.IgM|Protein fractions.oligoclonal bands.IgM
C2734989|T201|COMP|56764-4|LNC|Protein fractions.oligoclonal bands.IgG|Protein fractions.oligoclonal bands.IgG
C2734990|T201|COMP|56765-1|LNC|Protein fractions.oligoclonal bands.IgM|Protein fractions.oligoclonal bands.IgM
C2734991|T201|COMP|56766-9|LNC|Protein.monoclonal band 1/Protein.total|Protein.monoclonal band 1/Protein.total
C2734993|T201|COMP|56778-4|LNC|Articaine Ab.IgE|Articaine Ab.IgE
C2734995|T201|COMP|56779-2|LNC|Ascorbate|Ascorbate
C2734996|T201|COMP|56780-0|LNC|CYP21A2 gene mutations tested for|CYP21A2 gene mutations tested for
C2735000|T201|COMP|56782-6|LNC|Amylase.S4/Amylase.total|Amylase.S4/Amylase.total
C2735002|T201|COMP|56783-4|LNC|Trichloroethane|Trichloroethane
C2735003|T201|COMP|56784-2|LNC|Fibrinogen fragments|Fibrinogen fragments
C2735004|T201|COMP|56785-9|LNC|Saccharomyces cerevisiae Ab|Saccharomyces cerevisiae Ab
C2735005|T201|COMP|56786-7|LNC|Beta-2-Microglobulin.tumor marker|Beta-2-Microglobulin.tumor marker
C2735007|T201|COMP|56787-5|LNC|Cytokeratin 19|Cytokeratin 19
C2735008|T201|COMP|56788-3|LNC|Insulin^28H post XXX challenge|Insulin^28H post XXX challenge
C2735009|T201|COMP|56789-1|LNC|Insulin^32H post XXX challenge|Insulin^32H post XXX challenge
C2735010|T201|COMP|56790-9|LNC|Insulin^36H post XXX challenge|Insulin^36H post XXX challenge
C2735011|T201|COMP|56791-7|LNC|Entecavir|Entecavir
C2735012|T201|COMP|56792-5|LNC|Telbivudine|Telbivudine
C2735013|T201|COMP|56793-3|LNC|Tenefovir|Tenefovir
C2735153|T201|COMP|56877-4|LNC|Mepivacaine Ab.IgE|Mepivacaine Ab.IgE
C2735155|T201|COMP|56878-2|LNC|Phenylbutazone Ab.IgE|Phenylbutazone Ab.IgE
C2735157|T201|COMP|56879-0|LNC|Lactose Ab.IgE|Lactose Ab.IgE
C2735159|T201|COMP|56880-8|LNC|TCRB gene+TCRD gene+TCRG gene rearrangements|TCRB gene+TCRD gene+TCRG gene rearrangements
C2735161|T201|COMP|56881-6|LNC|Rickettsia typhi Ab.IgG|Rickettsia typhi Ab.IgG
C2735162|T201|COMP|56882-4|LNC|Parietaria judaica recombinant (rPar j) 2 Ab.IgE|Parietaria judaica recombinant (rPar j) 2 Ab.IgE
C2735164|T201|COMP|56883-2|LNC|BCHE gene targeted mutation analysis|BCHE gene targeted mutation analysis
C2735166|T201|COMP|56884-0|LNC|Somatotropin^160M post exercise|Somatotropin^160M post exercise
C2735167|T201|COMP|56885-7|LNC|Somatotropin^3H post exercise|Somatotropin^3H post exercise
C2735168|T201|COMP|56893-1|LNC|Cells.CD13+HLA-DR+/100 cells|Cells.CD13+HLA-DR+/100 cells
C2735169|T201|COMP|56894-9|LNC|Cells.CD13+HLA-DR+/100 cells|Cells.CD13+HLA-DR+/100 cells
C2735170|T201|COMP|56895-6|LNC|Cells.CD13+HLA-DR+/100 cells|Cells.CD13+HLA-DR+/100 cells
C2735171|T201|COMP|56896-4|LNC|Cells.CD33+CD34+/100 cells|Cells.CD33+CD34+/100 cells
C2735172|T201|COMP|56897-2|LNC|Cells.CD3-CD56+/100 cells|Cells.CD3-CD56+/100 cells
C2735173|T201|COMP|56898-0|LNC|Cells.CD5+FMC7+/100 cells|Cells.CD5+FMC7+/100 cells
C2735175|T201|COMP|56899-8|LNC|Cells.CD5+FMC7+/100 cells|Cells.CD5+FMC7+/100 cells
C2735177|T201|COMP|56901-2|LNC|Amino acid pattern|Amino acid pattern
C2735178|T201|COMP|56902-0|LNC|Amylase/Creatinine|Amylase/Creatinine
C2735179|T201|COMP|56903-8|LNC|Anserine/Creatinine|Anserine/Creatinine
C2735180|T201|COMP|56904-6|LNC|APOE gene mutation analysis|APOE gene mutation analysis
C2735181|T201|COMP|56905-3|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C2735182|T201|COMP|56906-1|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C2735183|T201|COMP|56907-9|LNC|Cells.CD3+CD45+/100 cells|Cells.CD3+CD45+/100 cells
C2735185|T201|COMP|56908-7|LNC|Cells.CD3+CD8+CD45+/100 cells|Cells.CD3+CD8+CD45+/100 cells
C2735187|T201|COMP|56909-5|LNC|Chlamydia sp Ab.IgG|Chlamydia sp Ab.IgG
C2735188|T201|COMP|56910-3|LNC|Chlamydia sp Ab.IgG^1st specimen|Chlamydia sp Ab.IgG^1st specimen
C2735189|T201|COMP|56911-1|LNC|Chlamydia sp Ab.IgG^2nd specimen|Chlamydia sp Ab.IgG^2nd specimen
C2735190|T201|COMP|56912-9|LNC|Cholesterol|Cholesterol
C2735191|T201|COMP|56913-7|LNC|Corticotropin^morning specimen|Corticotropin^morning specimen
C2735192|T201|COMP|56914-5|LNC|Corticotropin^evening specimen|Corticotropin^evening specimen
C2735193|T201|COMP|56915-2|LNC|Coxiella burnetii Ab.IgG|Coxiella burnetii Ab.IgG
C2735194|T201|COMP|56916-0|LNC|Coxiella burnetii Ab.IgM^2nd specimen|Coxiella burnetii Ab.IgM^2nd specimen
C2735195|T201|COMP|56917-8|LNC|Coxiella burnetii Ab.IgM|Coxiella burnetii Ab.IgM
C2735196|T201|COMP|56918-6|LNC|Coxiella burnetii Ab.IgM^1st specimen|Coxiella burnetii Ab.IgM^1st specimen
C2735197|T201|COMP|56919-4|LNC|Coxiella burnetii Ab.IgG^2nd specimen|Coxiella burnetii Ab.IgG^2nd specimen
C2735198|T201|COMP|56920-2|LNC|Coxiella burnetii Ab.IgG^1st specimen|Coxiella burnetii Ab.IgG^1st specimen
C2735199|T201|COMP|56921-0|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C2735200|T201|COMP|56922-8|LNC|Entamoeba histolytica Ab.IgG|Entamoeba histolytica Ab.IgG
C2735201|T201|COMP|56923-6|LNC|Fasciola hepatica Ab|Fasciola hepatica Ab
C2735202|T201|COMP|56924-4|LNC|Fasciola hepatica Ab|Fasciola hepatica Ab
C2735203|T201|COMP|56925-1|LNC|Fractional excretion of phosphate|Fractional excretion of phosphate
C2735204|T201|COMP|56926-9|LNC|Hepatitis C virus c1 Ab|Hepatitis C virus c1 Ab
C2735206|T201|COMP|56927-7|LNC|Hepatitis C virus c2 Ab|Hepatitis C virus c2 Ab
C2735208|T201|COMP|56928-5|LNC|Hepatitis C virus E2 Ab|Hepatitis C virus E2 Ab
C2735210|T201|COMP|56929-3|LNC|Hepatitis C virus NS3 Ab|Hepatitis C virus NS3 Ab
C2735212|T201|COMP|56930-1|LNC|Hepatitis C virus NS4 Ab|Hepatitis C virus NS4 Ab
C2735214|T201|COMP|56931-9|LNC|Hydrogen/Expired gas^pre dose lactulose|Hydrogen/Expired gas^pre dose lactulose
C2735215|T201|COMP|56932-7|LNC|Hydrogen/Expired gas^1H post dose lactulose|Hydrogen/Expired gas^1H post dose lactulose
C2735216|T201|COMP|56933-5|LNC|Hydrogen/Expired gas^2H post dose lactulose|Hydrogen/Expired gas^2H post dose lactulose
C2735217|T201|COMP|56934-3|LNC|Hydrogen/Expired gas^2.5H post dose lactulose|Hydrogen/Expired gas^2.5H post dose lactulose
C2735218|T201|COMP|56935-0|LNC|Hydrogen/Expired gas^3.5H post dose lactulose|Hydrogen/Expired gas^3.5H post dose lactulose
C2735219|T201|COMP|56936-8|LNC|Hydrogen/Expired gas^1.5H post dose lactulose|Hydrogen/Expired gas^1.5H post dose lactulose
C2735220|T201|COMP|56937-6|LNC|Hydrogen/Expired gas^30M post dose glucose|Hydrogen/Expired gas^30M post dose glucose
C2735221|T201|COMP|56938-4|LNC|Hydrogen/Expired gas^30M post dose lactulose|Hydrogen/Expired gas^30M post dose lactulose
C2735222|T201|COMP|56939-2|LNC|Hydroxyproline/Creatinine|Hydroxyproline/Creatinine
C2735223|T201|COMP|56940-0|LNC|Inhibin B|Inhibin B
C2735224|T201|COMP|56941-8|LNC|Insulin^8H post XXX challenge|Insulin^8H post XXX challenge
C2735225|T201|COMP|56942-6|LNC|Insulin^64H post XXX challenge|Insulin^64H post XXX challenge
C2735226|T201|COMP|56943-4|LNC|Insulin^68H post XXX challenge|Insulin^68H post XXX challenge
C2735230|T201|COMP|56944-2|LNC|Insulin^3D post XXX challenge|Insulin^3D post XXX challenge
C2735231|T201|COMP|56945-9|LNC|Insulin^56H post XXX challenge|Insulin^56H post XXX challenge
C2735232|T201|COMP|56946-7|LNC|Insulin^2D post XXX challenge|Insulin^2D post XXX challenge
C2735233|T201|COMP|56947-5|LNC|Insulin^60H post XXX challenge|Insulin^60H post XXX challenge
C2735234|T201|COMP|56948-3|LNC|Insulin^44H post XXX challenge|Insulin^44H post XXX challenge
C2735235|T201|COMP|56949-1|LNC|Insulin^40H post XXX challenge|Insulin^40H post XXX challenge
C2735236|T201|COMP|56957-4|LNC|Methionine/Creatinine|Methionine/Creatinine
C2735237|T201|COMP|56958-2|LNC|Mycoplasma pneumoniae Ab.IgG^1st specimen|Mycoplasma pneumoniae Ab.IgG^1st specimen
C2735238|T201|COMP|56959-0|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C2735239|T201|COMP|56960-8|LNC|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C2735240|T201|COMP|56961-6|LNC|Nicotinamide|Nicotinamide
C2735241|T201|COMP|56962-4|LNC|Ovary Ab.IgG|Ovary Ab.IgG
C2735243|T201|COMP|56964-0|LNC|Phosphate/Creatinine|Phosphate/Creatinine
C2735244|T201|COMP|56965-7|LNC|Phosphate/Creatinine|Phosphate/Creatinine
C2735245|T201|COMP|56966-5|LNC|Phosphoethanolamine/Creatinine|Phosphoethanolamine/Creatinine
C2735246|T201|COMP|56967-3|LNC|Plasmodium falciparum Ab|Plasmodium falciparum Ab
C2735247|T201|COMP|56968-1|LNC|Plasmodium sp Ab|Plasmodium sp Ab
C2735248|T201|COMP|56969-9|LNC|Polistes spp Ab.IgG4|Polistes spp Ab.IgG4
C2735249|T201|COMP|56970-7|LNC|Porphyrins|Porphyrins
C2735250|T201|COMP|56971-5|LNC|Potassium/Creatinine|Potassium/Creatinine
C2735251|T201|COMP|56972-3|LNC|Prolactin^post precipitation|Prolactin^post precipitation
C2735252|T201|COMP|56973-1|LNC|Proline/Creatinine|Proline/Creatinine
C2735253|T201|COMP|56974-9|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C2735254|T201|COMP|56975-6|LNC|Renin^upright+30M post XXX challenge|Renin^upright+30M post XXX challenge
C2735255|T201|COMP|56976-4|LNC|Renin^upright+1H post XXX challenge|Renin^upright+1H post XXX challenge
C2735256|T201|COMP|56977-2|LNC|Rheumatoid arthritis nuclear Ab|Rheumatoid arthritis nuclear Ab
C2735257|T201|COMP|56978-0|LNC|Serotonin|Serotonin
C2735258|T201|COMP|56979-8|LNC|Sodium|Sodium
C2735259|T201|COMP|56980-6|LNC|Sodium/Creatinine|Sodium/Creatinine
C2735260|T201|COMP|56981-4|LNC|Somatotropin^30M post resting|Somatotropin^30M post resting
C2735261|T201|COMP|56982-2|LNC|Somatotropin^90M post resting|Somatotropin^90M post resting
C2735262|T201|COMP|56983-0|LNC|Somatotropin^1H post resting|Somatotropin^1H post resting
C2735263|T201|COMP|56984-8|LNC|Taenia solium larva Ab|Taenia solium larva Ab
C2735264|T201|COMP|56985-5|LNC|Taurine/Creatinine|Taurine/Creatinine
C2735265|T201|COMP|56997-0|LNC|Urea/Creatinine|Urea/Creatinine
C2735266|T201|COMP|56998-8|LNC|Valine/Creatinine|Valine/Creatinine
C2735267|T201|COMP|56999-6|LNC|Vespa crabro Ab.IgG4|Vespa crabro Ab.IgG4
C2735269|T201|COMP|57000-2|LNC|Vespula spp Ab.IgG4|Vespula spp Ab.IgG4
C2735270|T201|COMP|57001-0|LNC|Yersinia sp Ab.IgA|Yersinia sp Ab.IgA
C2735271|T201|COMP|57002-8|LNC|11-Deoxycortisol^4D post XXX challenge|11-Deoxycortisol^4D post XXX challenge
C2735272|T201|COMP|57003-6|LNC|17-Hydroxyprogesterone^4H post XXX challenge|17-Hydroxyprogesterone^4H post XXX challenge
C2735273|T201|COMP|57004-4|LNC|Glucose/Creatinine|Glucose/Creatinine
C2735274|T201|COMP|57005-1|LNC|Glutathione|Glutathione
C2735275|T201|COMP|57006-9|LNC|Hepatitis C virus Ab.IgG|Hepatitis C virus Ab.IgG
C2735276|T201|COMP|57007-7|LNC|Insulin^52H post XXX challenge|Insulin^52H post XXX challenge
C2735277|T201|COMP|57008-5|LNC|Legionella pneumophila Ab.IgG^1st specimen|Legionella pneumophila Ab.IgG^1st specimen
C2735278|T201|COMP|57009-3|LNC|Mycoplasma pneumoniae Ab.IgG^2nd specimen|Mycoplasma pneumoniae Ab.IgG^2nd specimen
C2735279|T201|COMP|57010-1|LNC|Nuclear Ab|Nuclear Ab
C2735280|T201|COMP|57011-9|LNC|Ornithine/Creatinine|Ornithine/Creatinine
C2735281|T201|COMP|57012-7|LNC|Osteoblasts/100 cells|Osteoblasts/100 cells
C2735283|T201|COMP|57013-5|LNC|Phosphoserine/Creatinine|Phosphoserine/Creatinine
C2735284|T201|COMP|57014-3|LNC|Iron/Creatinine|Iron/Creatinine
C2735285|T201|COMP|57015-0|LNC|Lactulose.PO|Lactulose.PO
C2735291|T201|COMP|57038-2|LNC|Chromosome 12 aneuploidy|Chromosome 12 aneuploidy
C2735368|T201|COMP|57084-6|LNC|Fatty acid oxidation newborn screen panel|Fatty acid oxidation newborn screen panel
C2735370|T201|COMP|57085-3|LNC|Organic acid newborn screen panel|Organic acid newborn screen panel
C2735374|T201|COMP|57087-9|LNC|Biotinidase newborn screening panel|Biotinidase newborn screening panel
C2735377|T201|COMP|57089-5|LNC|Eosinophil cationic protein|Eosinophil cationic protein
C2735378|T201|COMP|57090-3|LNC|HLA-DQA1*05:01|HLA-DQA1*05:01
C2735379|T201|COMP|57091-1|LNC|HLA-DQB1*02:01|HLA-DQB1*02:01
C2735380|T201|COMP|57092-9|LNC|IgE|IgE
C2735381|T201|COMP|57093-7|LNC|Cyclic citrullinated peptide Ab.IgA+IgG|Cyclic citrullinated peptide Ab.IgA+IgG
C2735382|T201|COMP|57094-5|LNC|Phenol^^adjusted to specific gravity 1.024|Phenol^^adjusted to specific gravity 1.024
C2735383|T201|COMP|57095-2|LNC|Anidulafungin|Anidulafungin
C2735384|T201|COMP|57096-0|LNC|HPA 1a-1a+HPA 3a-3a|HPA 1a-1a+HPA 3a-3a
C2735423|T201|COMP|57128-1|LNC|Newborn Screening Report summary panel|Newborn Screening Report summary panel
C2735427|T201|COMP|57308-9|LNC|CYP11B1 gene targeted mutation analysis|CYP11B1 gene targeted mutation analysis
C2735429|T201|COMP|57309-7|LNC|PRNP gene targeted mutation analysis|PRNP gene targeted mutation analysis
C2735431|T201|COMP|57310-5|LNC|SRY gene targeted mutation analysis|SRY gene targeted mutation analysis
C2735433|T201|COMP|57311-3|LNC|CYP11B1 gene mutations tested for|CYP11B1 gene mutations tested for
C2735435|T201|COMP|57312-1|LNC|PRNP gene mutations tested for|PRNP gene mutations tested for
C2735437|T201|COMP|57313-9|LNC|Pyrazole Ab.IgE|Pyrazole Ab.IgE
C2735439|T201|COMP|57314-7|LNC|SRY gene mutations tested for|SRY gene mutations tested for
C2735441|T201|COMP|57315-4|LNC|Sulphonamide Ab.IgE|Sulphonamide Ab.IgE
C2735443|T201|COMP|57316-2|LNC|Tropomyosin Ab.IgE|Tropomyosin Ab.IgE
C2735445|T201|COMP|57317-0|LNC|Chromosome 13+18+21+X+Y aneuploidy|Chromosome 13+18+21+X+Y aneuploidy
C2735446|T201|COMP|57318-8|LNC|Chromosome 13+18+21+X+Y aneuploidy|Chromosome 13+18+21+X+Y aneuploidy
C2735449|T201|COMP|57320-4|LNC|Trypanosoma cruzi Ab|Trypanosoma cruzi Ab
C2735451|T201|COMP|57487-1|LNC|11-Ketoetiocholanolone^pre dose dexamethasone|11-Ketoetiocholanolone^pre dose dexamethasone
C2735452|T201|COMP|57488-9|LNC|11-Ketoetiocholanolone^pre dose dexamethasone|11-Ketoetiocholanolone^pre dose dexamethasone
C2735453|T201|COMP|57489-7|LNC|11-Ketoetiocholanolone^2D post dose dexamethasone|11-Ketoetiocholanolone^2D post dose dexamethasone
C2735454|T201|COMP|57490-5|LNC|11-Ketoetiocholanolone^2D post dose dexamethasone|11-Ketoetiocholanolone^2D post dose dexamethasone
C2735455|T201|COMP|57491-3|LNC|11-Deoxycorticosterone^pre 250 ug corticotropin|11-Deoxycorticosterone^pre 250 ug corticotropin
C2735456|T201|COMP|57770-0|LNC|Toxoplasma gondii Ab.IgG & IgM panel|Toxoplasma gondii Ab.IgG & IgM panel
C2735458|T201|COMP|57771-8|LNC|Paraneoplastic Ab|Paraneoplastic Ab
C2735459|T201|COMP|57772-6|LNC|Metanephrine.free & Normetanephrine.free panel|Metanephrine.free & Normetanephrine.free panel
C2735461|T201|COMP|57773-4|LNC|Colorado tick fever virus Ab.IgG & IgM|Colorado tick fever virus Ab.IgG & IgM
C2735463|T201|COMP|57774-2|LNC|Colorado tick fever virus Ab.IgG & IgM panel|Colorado tick fever virus Ab.IgG & IgM panel
C2735464|T201|COMP|57775-9|LNC|Valproate.free & Valproate panel|Valproate.free & Valproate panel
C2735466|T201|COMP|57776-7|LNC|Gliadin peptide Ab.IgA & IgG panel|Gliadin peptide Ab.IgA & IgG panel
C2735468|T201|COMP|57934-2|LNC|Chikungunya virus Ab.IgM|Chikungunya virus Ab.IgM
C2735469|T201|COMP|57936-7|LNC|Cholesterol.in HDL 2a|Cholesterol.in HDL 2a
C2735470|T201|COMP|57937-5|LNC|Cholesterol.in HDL 3a|Cholesterol.in HDL 3a
C2735471|T201|COMP|57938-3|LNC|LDL 5|LDL 5
C2735473|T201|COMP|57939-1|LNC|Chromium|Chromium
C2735478|T201|COMP|58092-8|LNC|Acylcarnitine newborn screen panel|Acylcarnitine newborn screen panel
C2735492|T201|COMP|57130-7|LNC|Newborn screening report - overall interpretation|Newborn screening report - overall interpretation
C2735494|T201|COMP|57131-5|LNC|Newborn conditions with positive markers|Newborn conditions with positive markers
C2735496|T201|COMP|57132-3|LNC|CYP2C19 gene targeted mutation analysis|CYP2C19 gene targeted mutation analysis
C2735526|T201|COMP|57374-1|LNC|Oxalate|Oxalate
C2735527|T201|COMP|57375-8|LNC|Oxalate|Oxalate
C2735528|T201|COMP|57376-6|LNC|C peptide^baseline|C peptide^baseline
C2735529|T201|COMP|57377-4|LNC|Pyruvate^5M post XXX challenge|Pyruvate^5M post XXX challenge
C2735530|T201|COMP|57378-2|LNC|Porphyrins/Creatinine|Porphyrins/Creatinine
C2735531|T201|COMP|57379-0|LNC|Potassium|Potassium
C2735532|T201|COMP|57380-8|LNC|Potassium|Potassium
C2735533|T201|COMP|57398-0|LNC|Cells.CD22+CD19+/100 cells|Cells.CD22+CD19+/100 cells
C2735534|T201|COMP|57399-8|LNC|Cells.CD19+CD23+/100 cells|Cells.CD19+CD23+/100 cells
C2735535|T201|COMP|57400-4|LNC|Cells.CD34/100 cells|Cells.CD34/100 cells
C2735536|T201|COMP|57401-2|LNC|Cells.CD4+CD8+/100 cells|Cells.CD4+CD8+/100 cells
C2735537|T201|COMP|57402-0|LNC|Cells.CD42a/100 cells|Cells.CD42a/100 cells
C2735538|T201|COMP|57403-8|LNC|Cells.CD45RA/100 cells|Cells.CD45RA/100 cells
C2735539|T201|COMP|57404-6|LNC|Cells.CD45RO/100 cells|Cells.CD45RO/100 cells
C2735540|T201|COMP|57405-3|LNC|Cells.CD8+CD56+/100 cells|Cells.CD8+CD56+/100 cells
C2735541|T201|COMP|57554-8|LNC|18-Hydroxycorticosterone^pre dose corticotropin|18-Hydroxycorticosterone^pre dose corticotropin
C2735544|T201|COMP|57557-1|LNC|18-Hydroxycortisol^pre dose corticotropin|18-Hydroxycortisol^pre dose corticotropin
C2735545|T201|COMP|57700-7|LNC|Hearing loss newborn screening comment-discussion|Hearing loss newborn screening comment-discussion
C2735549|T201|COMP|57702-3|LNC|Infectious diseases|Infectious diseases
C2735566|T201|COMP|57711-4|LNC|Unique bar code number|Unique bar code number
C2735573|T201|COMP|57180-2|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C2735576|T201|COMP|57182-8|LNC|HIV 1 RNA tropism|HIV 1 RNA tropism
C2735714|T201|COMP|57287-5|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C2735715|T201|COMP|57288-3|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C2735716|T201|COMP|57289-1|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2735717|T201|COMP|57290-9|LNC|HLA-A|HLA-A
C2735718|T201|COMP|57291-7|LNC|HLA-B|HLA-B
C2735719|T201|COMP|57292-5|LNC|HLA-B57*01|HLA-B57*01
C2735721|T201|COMP|57293-3|LNC|HLA-DRB1|HLA-DRB1
C2735722|T201|COMP|57294-1|LNC|HLA-DRB3|HLA-DRB3
C2735723|T201|COMP|57295-8|LNC|HLA-DRB4|HLA-DRB4
C2735724|T201|COMP|57296-6|LNC|HLA-DRB5|HLA-DRB5
C2735725|T201|COMP|57297-4|LNC|HLA-Cw|HLA-Cw
C2735726|T201|COMP|57299-0|LNC|HLA-DQB1|HLA-DQB1
C2735727|T201|COMP|57300-6|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C2735728|T201|COMP|57301-4|LNC|Benzoylecgonine|Benzoylecgonine
C2735729|T201|COMP|57302-2|LNC|Temazepam|Temazepam
C2735730|T201|COMP|57303-0|LNC|7-Aminonitrazepam|7-Aminonitrazepam
C2735731|T201|COMP|57304-8|LNC|Codeine|Codeine
C2735732|T201|COMP|57305-5|LNC|Tropomyosin Ab.IgE|Tropomyosin Ab.IgE
C2735735|T201|COMP|57321-2|LNC|Herpes simplex virus 2 Ab.IgG^2nd specimen|Herpes simplex virus 2 Ab.IgG^2nd specimen
C2735736|T201|COMP|57322-0|LNC|Varicella zoster virus Ab.IgM^1st specimen|Varicella zoster virus Ab.IgM^1st specimen
C2735737|T201|COMP|57334-5|LNC|Calcium|Calcium
C2735738|T201|COMP|57335-2|LNC|Calcium|Calcium
C2735739|T201|COMP|57336-0|LNC|Beta hydroxybutyrate^1H post XXX challenge|Beta hydroxybutyrate^1H post XXX challenge
C2735740|T201|COMP|57337-8|LNC|Citrate|Citrate
C2735741|T201|COMP|57338-6|LNC|Citrate|Citrate
C2735742|T201|COMP|57339-4|LNC|Citrate|Citrate
C2735743|T201|COMP|57340-2|LNC|Chloride|Chloride
C2735744|T201|COMP|57341-0|LNC|Chloride|Chloride
C2735745|T201|COMP|57342-8|LNC|Chloride|Chloride
C2735746|T201|COMP|57344-4|LNC|Creatinine|Creatinine
C2735747|T201|COMP|57345-1|LNC|Creatinine^overnight|Creatinine^overnight
C2735748|T201|COMP|57346-9|LNC|Creatinine|Creatinine
C2735749|T201|COMP|57347-7|LNC|Copper|Copper
C2735750|T201|COMP|57348-5|LNC|Phosphate|Phosphate
C2735751|T201|COMP|57349-3|LNC|Phosphate|Phosphate
C2735752|T201|COMP|57350-1|LNC|Glucose^1M post XXX challenge|Glucose^1M post XXX challenge
C2735753|T201|COMP|57353-5|LNC|Insulin^5M post XXX challenge|Insulin^5M post XXX challenge
C2735754|T201|COMP|57355-0|LNC|Potassium|Potassium
C2735755|T201|COMP|57356-8|LNC|Lactate^1M post XXX challenge|Lactate^1M post XXX challenge
C2735756|T201|COMP|57357-6|LNC|Lactate^10M post XXX challenge|Lactate^10M post XXX challenge
C2735757|T201|COMP|57358-4|LNC|Lactate^2H post XXX challenge|Lactate^2H post XXX challenge
C2735758|T201|COMP|57359-2|LNC|Lactate^3H post XXX challenge|Lactate^3H post XXX challenge
C2735759|T201|COMP|57360-0|LNC|Lactate^20M post XXX challenge|Lactate^20M post XXX challenge
C2735760|T201|COMP|57361-8|LNC|Lactate^3M post XXX challenge|Lactate^3M post XXX challenge
C2735761|T201|COMP|57362-6|LNC|Lactate^30M post XXX challenge|Lactate^30M post XXX challenge
C2735762|T201|COMP|57363-4|LNC|Lactate^5M post XXX challenge|Lactate^5M post XXX challenge
C2735763|T201|COMP|57364-2|LNC|Lactate^1H post XXX challenge|Lactate^1H post XXX challenge
C2735764|T201|COMP|57365-9|LNC|Lactate^1.5H post XXX challenge|Lactate^1.5H post XXX challenge
C2735765|T201|COMP|57367-5|LNC|Magnesium|Magnesium
C2735766|T201|COMP|57368-3|LNC|Magnesium|Magnesium
C2735767|T201|COMP|57369-1|LNC|Albumin|Albumin
C2735768|T201|COMP|57370-9|LNC|Sodium|Sodium
C2735769|T201|COMP|57371-7|LNC|Enolase.neuron specific|Enolase.neuron specific
C2735770|T201|COMP|57372-5|LNC|Osmolality|Osmolality
C2735771|T201|COMP|57373-3|LNC|Oxalate|Oxalate
C2735772|T201|COMP|57407-9|LNC|Cells.CD8+CD45RA+/100 cells|Cells.CD8+CD45RA+/100 cells
C2735774|T201|COMP|57408-7|LNC|Cells.CD8+CD45RO+/100 cells|Cells.CD8+CD45RO+/100 cells
C2735776|T201|COMP|57409-5|LNC|Cells.CD3+TCR alpha beta+/100 cells|Cells.CD3+TCR alpha beta+/100 cells
C2735777|T201|COMP|57410-3|LNC|Actin.filamentous Ab|Actin.filamentous Ab
C2735778|T201|COMP|57411-1|LNC|Desmoglein 1 Ab|Desmoglein 1 Ab
C2735779|T201|COMP|57412-9|LNC|Desmoglein 3 Ab|Desmoglein 3 Ab
C2735780|T201|COMP|57413-7|LNC|Mitochondria Ab|Mitochondria Ab
C2735781|T201|COMP|57414-5|LNC|Reticulin Ab|Reticulin Ab
C2735782|T201|COMP|57415-2|LNC|Saccharomyces cerevisiae Ab.IgA|Saccharomyces cerevisiae Ab.IgA
C2735783|T201|COMP|57416-0|LNC|Thyrotropin receptor Ab|Thyrotropin receptor Ab
C2735784|T201|COMP|57417-8|LNC|Cells.CD18/100 cells|Cells.CD18/100 cells
C2735785|T201|COMP|57418-6|LNC|Cells.CD20/100 cells|Cells.CD20/100 cells
C2735786|T201|COMP|57419-4|LNC|Cells.CD21/100 cells|Cells.CD21/100 cells
C2735787|T201|COMP|57420-2|LNC|Cells.CD27/100 cells|Cells.CD27/100 cells
C2735788|T201|COMP|57421-0|LNC|Cells.CD34/100 cells|Cells.CD34/100 cells
C2735789|T201|COMP|57422-8|LNC|Cells.CD40/100 cells|Cells.CD40/100 cells
C2735790|T201|COMP|57423-6|LNC|Cells.CD5/100 cells|Cells.CD5/100 cells
C2735791|T201|COMP|57424-4|LNC|Cells.CD56/100 cells|Cells.CD56/100 cells
C2735792|T201|COMP|57425-1|LNC|Cells.CD7/100 cells|Cells.CD7/100 cells
C2735793|T201|COMP|57426-9|LNC|Cells.CD71/100 cells|Cells.CD71/100 cells
C2735794|T201|COMP|57427-7|LNC|Cells.CD10+FMC7+/100 cells|Cells.CD10+FMC7+/100 cells
C2735796|T201|COMP|57428-5|LNC|Cells.FMC7/100 cells|Cells.FMC7/100 cells
C2735797|T201|COMP|57429-3|LNC|Cells.CD3+TCR gamma delta+/100 cells|Cells.CD3+TCR gamma delta+/100 cells
C2735798|T201|COMP|57430-1|LNC|Cells.CD235a/100 cells|Cells.CD235a/100 cells
C2735799|T201|COMP|57431-9|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C2735800|T201|COMP|57432-7|LNC|Cells.CD19+Kappa+/100 cells|Cells.CD19+Kappa+/100 cells
C2735801|T201|COMP|57433-5|LNC|Cells.CD19+Lambda+/100 cells|Cells.CD19+Lambda+/100 cells
C2735802|T201|COMP|57434-3|LNC|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C2735803|T201|COMP|57435-0|LNC|Cells.myeloperoxidase|Cells.myeloperoxidase
C2735804|T201|COMP|57436-8|LNC|Muscle specific receptor tyrosine kinase Ab|Muscle specific receptor tyrosine kinase Ab
C2735805|T201|COMP|57437-6|LNC|Cells.CD56+CD138+/100 cells|Cells.CD56+CD138+/100 cells
C2735807|T201|COMP|57438-4|LNC|Cells.CD56-CD138+/100 cells|Cells.CD56-CD138+/100 cells
C2735809|T201|COMP|57439-2|LNC|Cells.terminal deoxyribonucleotidyl transferase|Cells.terminal deoxyribonucleotidyl transferase
C2735810|T201|COMP|57440-0|LNC|Platelet Ab|Platelet Ab
C2735811|T201|COMP|57441-8|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C2735812|T201|COMP|57442-6|LNC|Specimen volume^post concentration|Specimen volume^post concentration
C2735817|T201|COMP|57447-5|LNC|Nuclear Ab|Nuclear Ab
C2735818|T201|COMP|57448-3|LNC|Nuclear Ab pattern|Nuclear Ab pattern
C2735819|T201|COMP|57449-1|LNC|Tubular basement membrane Ab|Tubular basement membrane Ab
C2735820|T201|COMP|57450-9|LNC|Soluble liver Ab|Soluble liver Ab
C2735821|T201|COMP|57451-7|LNC|CV2 Ab|CV2 Ab
C2735822|T201|COMP|57452-5|LNC|Ma+Ta Ab|Ma+Ta Ab
C2735823|T201|COMP|57453-3|LNC|Chromosome 18 aneuploidy|Chromosome 18 aneuploidy
C2735825|T201|COMP|57454-1|LNC|Chromosome 13 aneuploidy|Chromosome 13 aneuploidy
C2735827|T201|COMP|57455-8|LNC|Taenia solium Ab.IgG|Taenia solium Ab.IgG
C2735828|T201|COMP|57456-6|LNC|Spermatozoa.progressive^post concentration|Spermatozoa.progressive^post concentration
C2735829|T201|COMP|57457-4|LNC|Interpretation|Interpretation
C2735830|T201|COMP|57458-2|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2735835|T201|COMP|57462-4|LNC|Normetanephrine.free|Normetanephrine.free
C2735836|T201|COMP|57463-2|LNC|Cortisol^12th specimen|Cortisol^12th specimen
C2735837|T201|COMP|57464-0|LNC|Cortisol^11th specimen|Cortisol^11th specimen
C2735838|T201|COMP|57465-7|LNC|Cortisol^10th specimen|Cortisol^10th specimen
C2735839|T201|COMP|57466-5|LNC|Cortisol^9th specimen|Cortisol^9th specimen
C2735840|T201|COMP|57467-3|LNC|Calcitriol^pre dose calcium|Calcitriol^pre dose calcium
C2735841|T201|COMP|57468-1|LNC|Calcitriol^pre dose calcium|Calcitriol^pre dose calcium
C2735842|T201|COMP|57469-9|LNC|Calcitriol^2H post dose calcium|Calcitriol^2H post dose calcium
C2735843|T201|COMP|57470-7|LNC|Calcitriol^2H post dose calcium|Calcitriol^2H post dose calcium
C2735844|T201|COMP|57471-5|LNC|Calcitriol^3H post dose calcium|Calcitriol^3H post dose calcium
C2735845|T201|COMP|57472-3|LNC|Calcitriol^3H post dose calcium|Calcitriol^3H post dose calcium
C2735846|T201|COMP|57473-1|LNC|Calcitriol^1H post dose calcium|Calcitriol^1H post dose calcium
C2735847|T201|COMP|57474-9|LNC|Calcitriol^1H post dose calcium|Calcitriol^1H post dose calcium
C2735848|T201|COMP|57475-6|LNC|11-Ketoandrosterone^pre high dose dexamethasone|11-Ketoandrosterone^pre high dose dexamethasone
C2735849|T201|COMP|57476-4|LNC|11-Ketoandrosterone^pre high dose dexamethasone|11-Ketoandrosterone^pre high dose dexamethasone
C2735852|T201|COMP|57479-8|LNC|11-Ketoandrosterone^pre dose dexamethasone|11-Ketoandrosterone^pre dose dexamethasone
C2735853|T201|COMP|57480-6|LNC|11-Ketoandrosterone^pre dose dexamethasone|11-Ketoandrosterone^pre dose dexamethasone
C2735854|T201|COMP|57481-4|LNC|11-Ketoandrosterone^2D post dose dexamethasone|11-Ketoandrosterone^2D post dose dexamethasone
C2735855|T201|COMP|57482-2|LNC|11-Ketoandrosterone^2D post dose dexamethasone|11-Ketoandrosterone^2D post dose dexamethasone
C2735861|T201|COMP|57494-7|LNC|11-Deoxycortisol^pre dose dexamethasone|11-Deoxycortisol^pre dose dexamethasone
C2735862|T201|COMP|57495-4|LNC|11-Deoxycortisol^pre dose dexamethasone|11-Deoxycortisol^pre dose dexamethasone
C2735863|T201|COMP|57496-2|LNC|11-Deoxycortisol^1D post dose dexamethasone|11-Deoxycortisol^1D post dose dexamethasone
C2735864|T201|COMP|57497-0|LNC|11-Deoxycortisol^1D post dose dexamethasone|11-Deoxycortisol^1D post dose dexamethasone
C2735865|T201|COMP|57498-8|LNC|11-Deoxycortisol^2D post dose dexamethasone|11-Deoxycortisol^2D post dose dexamethasone
C2735866|T201|COMP|57499-6|LNC|11-Deoxycortisol^2D post dose dexamethasone|11-Deoxycortisol^2D post dose dexamethasone
C2735867|T201|COMP|57500-1|LNC|11-Deoxycortisol^pre dose metyraPONE|11-Deoxycortisol^pre dose metyraPONE
C2735868|T201|COMP|57501-9|LNC|11-Deoxycortisol^pre dose metyraPONE|11-Deoxycortisol^pre dose metyraPONE
C2735869|T201|COMP|57502-7|LNC|11-Deoxycortisol^1D post dose metyraPONE|11-Deoxycortisol^1D post dose metyraPONE
C2735870|T201|COMP|57503-5|LNC|11-Deoxycortisol^1D post dose metyraPONE|11-Deoxycortisol^1D post dose metyraPONE
C2735871|T201|COMP|57504-3|LNC|11-Deoxycortisol^2D post dose metyraPONE|11-Deoxycortisol^2D post dose metyraPONE
C2735872|T201|COMP|57505-0|LNC|11-Deoxycortisol^2D post dose metyraPONE|11-Deoxycortisol^2D post dose metyraPONE
C2735873|T201|COMP|57506-8|LNC|11-Deoxycortisol^pre 250 ug corticotropin|11-Deoxycortisol^pre 250 ug corticotropin
C2735874|T201|COMP|57507-6|LNC|11-Deoxycortisol^45M post 250 ug corticotropin|11-Deoxycortisol^45M post 250 ug corticotropin
C2735879|T201|COMP|57512-6|LNC|11-Hydroxyandrosterone^pre dose dexamethasone|11-Hydroxyandrosterone^pre dose dexamethasone
C2735880|T201|COMP|57513-4|LNC|11-Hydroxyandrosterone^pre dose dexamethasone|11-Hydroxyandrosterone^pre dose dexamethasone
C2735881|T201|COMP|57514-2|LNC|11-Hydroxyandrosterone^2D post dose dexamethasone|11-Hydroxyandrosterone^2D post dose dexamethasone
C2735882|T201|COMP|57515-9|LNC|11-Hydroxyandrosterone^2D post dose dexamethasone|11-Hydroxyandrosterone^2D post dose dexamethasone
C2735887|T201|COMP|57520-9|LNC|11-Hydroxyetiocholanolone^pre dose dexamethasone|11-Hydroxyetiocholanolone^pre dose dexamethasone
C2735888|T201|COMP|57521-7|LNC|11-Hydroxyetiocholanolone^pre dose dexamethasone|11-Hydroxyetiocholanolone^pre dose dexamethasone
C2735891|T201|COMP|57524-1|LNC|17-Ketogenic steroids^pre dose dexamethasone|17-Ketogenic steroids^pre dose dexamethasone
C2735892|T201|COMP|57525-8|LNC|17-Ketogenic steroids^2D post dose dexamethasone|17-Ketogenic steroids^2D post dose dexamethasone
C2735895|T201|COMP|57528-2|LNC|17-Hydroxycorticosteroids^pre dose dexamethasone|17-Hydroxycorticosteroids^pre dose dexamethasone
C2735897|T201|COMP|57530-8|LNC|17-Hydroxypregnenolone^pre dose dexamethasone|17-Hydroxypregnenolone^pre dose dexamethasone
C2735898|T201|COMP|57531-6|LNC|17-Hydroxypregnenolone^1D post dose dexamethasone|17-Hydroxypregnenolone^1D post dose dexamethasone
C2735899|T201|COMP|57532-4|LNC|17-Hydroxypregnenolone^2D post dose dexamethasone|17-Hydroxypregnenolone^2D post dose dexamethasone
C2735912|T201|COMP|57545-6|LNC|17-Hydroxyprogesterone^pre dose dexamethasone|17-Hydroxyprogesterone^pre dose dexamethasone
C2735913|T201|COMP|57558-9|LNC|18-Hydroxycortisol^30M post dose corticotropin|18-Hydroxycortisol^30M post dose corticotropin
C2735914|T201|COMP|57559-7|LNC|18-Hydroxycortisol^1H post dose corticotropin|18-Hydroxycortisol^1H post dose corticotropin
C2735915|T201|COMP|57560-5|LNC|21-Deoxycorticosterone^pre dose corticotropin|21-Deoxycorticosterone^pre dose corticotropin
C2735918|T201|COMP|57562-1|LNC|21-Deoxycorticosterone^1H post dose corticotropin|21-Deoxycorticosterone^1H post dose corticotropin
C2735919|T201|COMP|57563-9|LNC|21-Deoxycortisol^pre dose dexamethasone|21-Deoxycortisol^pre dose dexamethasone
C2735920|T201|COMP|57564-7|LNC|21-Deoxycortisol^1D post dose dexamethasone|21-Deoxycortisol^1D post dose dexamethasone
C2735921|T201|COMP|57565-4|LNC|21-Deoxycortisol^2D post dose dexamethasone|21-Deoxycortisol^2D post dose dexamethasone
C2735922|T201|COMP|57566-2|LNC|Calcidiol^pre dose calcium|Calcidiol^pre dose calcium
C2735923|T201|COMP|57567-0|LNC|Calcidiol^2H post dose calcium|Calcidiol^2H post dose calcium
C2735924|T201|COMP|57568-8|LNC|Calcidiol^3H post dose calcium|Calcidiol^3H post dose calcium
C2735925|T201|COMP|57569-6|LNC|Calcidiol^1H post dose calcium|Calcidiol^1H post dose calcium
C2735928|T201|COMP|57630-6|LNC|Alpha cortolone^pre high dose dexamethasone|Alpha cortolone^pre high dose dexamethasone
C2735929|T201|COMP|57631-4|LNC|Alpha cortolone^2D post high dose dexamethasone|Alpha cortolone^2D post high dose dexamethasone
C2735930|T201|COMP|57632-2|LNC|Alpha cortolone^2D post high dose dexamethasone|Alpha cortolone^2D post high dose dexamethasone
C2735931|T201|COMP|57633-0|LNC|Alpha cortolone^pre dose dexamethasone|Alpha cortolone^pre dose dexamethasone
C2735932|T201|COMP|57634-8|LNC|Alpha cortolone^pre dose dexamethasone|Alpha cortolone^pre dose dexamethasone
C2735933|T201|COMP|57635-5|LNC|Alpha cortolone^2D post dose dexamethasone|Alpha cortolone^2D post dose dexamethasone
C2735934|T201|COMP|57636-3|LNC|Alpha cortolone^2D post dose dexamethasone|Alpha cortolone^2D post dose dexamethasone
C2735935|T201|COMP|57637-1|LNC|Androsterone^pre high dose dexamethasone|Androsterone^pre high dose dexamethasone
C2735936|T201|COMP|57638-9|LNC|Androsterone^pre high dose dexamethasone|Androsterone^pre high dose dexamethasone
C2735986|T201|COMP|57576-1|LNC|Androstanolone^pre dose corticotropin|Androstanolone^pre dose corticotropin
C2735987|T201|COMP|57577-9|LNC|Androstanolone^30M post dose corticotropin|Androstanolone^30M post dose corticotropin
C2735988|T201|COMP|57578-7|LNC|Androstanolone^1H post dose corticotropin|Androstanolone^1H post dose corticotropin
C2735989|T201|COMP|57579-5|LNC|Aldosterone^post 25 mg captopril PO|Aldosterone^post 25 mg captopril PO
C2735990|T201|COMP|57580-3|LNC|Aldosterone^post XXX challenge|Aldosterone^post XXX challenge
C2735991|T201|COMP|57582-9|LNC|Aldosterone^pre 25 mg captopril PO|Aldosterone^pre 25 mg captopril PO
C2735992|T201|COMP|57583-7|LNC|Aldosterone^2H post 25 mg captopril PO|Aldosterone^2H post 25 mg captopril PO
C2735993|T201|COMP|57584-5|LNC|Aldosterone^3H post 25 mg captopril PO|Aldosterone^3H post 25 mg captopril PO
C2735994|T201|COMP|57585-2|LNC|Aldosterone^3H post 25 mg captopril PO|Aldosterone^3H post 25 mg captopril PO
C2735995|T201|COMP|57586-0|LNC|Aldosterone^1H post 25 mg captopril PO|Aldosterone^1H post 25 mg captopril PO
C2735996|T201|COMP|57587-8|LNC|Aldosterone^2H post XXX challenge|Aldosterone^2H post XXX challenge
C2735997|T201|COMP|57588-6|LNC|Aldosterone^15M post XXX challenge|Aldosterone^15M post XXX challenge
C2735998|T201|COMP|57589-4|LNC|Aldosterone^15M post XXX challenge|Aldosterone^15M post XXX challenge
C2735999|T201|COMP|57590-2|LNC|Aldosterone^3H post XXX challenge|Aldosterone^3H post XXX challenge
C2736000|T201|COMP|57591-0|LNC|Aldosterone^3H post XXX challenge|Aldosterone^3H post XXX challenge
C2736001|T201|COMP|57592-8|LNC|Aldosterone^30M post XXX challenge|Aldosterone^30M post XXX challenge
C2736002|T201|COMP|57595-1|LNC|Aldosterone^1H post XXX challenge|Aldosterone^1H post XXX challenge
C2736003|T201|COMP|57596-9|LNC|Aldosterone^pre 250 ug corticotropin IM|Aldosterone^pre 250 ug corticotropin IM
C2736024|T201|COMP|57617-3|LNC|5-Alpha tetrahydrocortisol^pre dose dexamethasone|5-Alpha tetrahydrocortisol^pre dose dexamethasone
C2736025|T201|COMP|57618-1|LNC|5-Alpha tetrahydrocortisol^pre dose dexamethasone|5-Alpha tetrahydrocortisol^pre dose dexamethasone
C2736028|T201|COMP|57621-5|LNC|Alpha cortol^pre high dose dexamethasone|Alpha cortol^pre high dose dexamethasone
C2736029|T201|COMP|57622-3|LNC|Alpha cortol^pre high dose dexamethasone|Alpha cortol^pre high dose dexamethasone
C2736030|T201|COMP|57623-1|LNC|Alpha cortol^2D post high dose dexamethasone|Alpha cortol^2D post high dose dexamethasone
C2736031|T201|COMP|57624-9|LNC|Alpha cortol^2D post high dose dexamethasone|Alpha cortol^2D post high dose dexamethasone
C2736032|T201|COMP|57625-6|LNC|Alpha cortol^pre dose dexamethasone|Alpha cortol^pre dose dexamethasone
C2736033|T201|COMP|57626-4|LNC|Alpha cortol^pre dose dexamethasone|Alpha cortol^pre dose dexamethasone
C2736034|T201|COMP|57627-2|LNC|Alpha cortol^2D post dose dexamethasone|Alpha cortol^2D post dose dexamethasone
C2736035|T201|COMP|57628-0|LNC|Alpha cortol^2D post dose dexamethasone|Alpha cortol^2D post dose dexamethasone
C2736036|T201|COMP|57629-8|LNC|Alpha cortolone^pre high dose dexamethasone|Alpha cortolone^pre high dose dexamethasone
C2736037|T201|COMP|57794-0|LNC|Newborn screening test results panel|Newborn screening test results panel
C2736039|T201|COMP|57796-5|LNC|Reducing substances|Reducing substances
C2736040|T201|COMP|57797-3|LNC|Glucose|Glucose
C2736041|T201|COMP|57798-1|LNC|Progesterone^20M post XXX challenge|Progesterone^20M post XXX challenge
C2736042|T201|COMP|57800-5|LNC|Oxygen content|Oxygen content
C2736045|T201|COMP|57802-1|LNC|Chromosome analysis.interphase|Chromosome analysis.interphase
C2736046|T201|COMP|57803-9|LNC|Occult blood panel|Occult blood panel
C2736053|T201|COMP|57639-7|LNC|Androsterone^2D post high dose dexamethasone|Androsterone^2D post high dose dexamethasone
C2736054|T201|COMP|57640-5|LNC|Androsterone^2D post high dose dexamethasone|Androsterone^2D post high dose dexamethasone
C2736055|T201|COMP|57641-3|LNC|Androsterone^pre dose dexamethasone|Androsterone^pre dose dexamethasone
C2736056|T201|COMP|57642-1|LNC|Androsterone^pre dose dexamethasone|Androsterone^pre dose dexamethasone
C2736057|T201|COMP|57643-9|LNC|Androsterone^2D post dose dexamethasone|Androsterone^2D post dose dexamethasone
C2736058|T201|COMP|57644-7|LNC|Androsterone^2D post dose dexamethasone|Androsterone^2D post dose dexamethasone
C2736059|T201|COMP|57646-2|LNC|C peptide^190M post XXX challenge|C peptide^190M post XXX challenge
C2736060|T201|COMP|57647-0|LNC|C peptide^3.3H post XXX challenge|C peptide^3.3H post XXX challenge
C2736061|T201|COMP|57651-2|LNC|C peptide^1.3H post XXX challenge|C peptide^1.3H post XXX challenge
C2736076|T201|COMP|57660-3|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C2736077|T201|COMP|57661-1|LNC|Tubular basement membrane Ab|Tubular basement membrane Ab
C2736078|T201|COMP|57662-9|LNC|U1 small nuclear ribonucleoprotein Ab|U1 small nuclear ribonucleoprotein Ab
C2736079|T201|COMP|57663-7|LNC|Norepinephrine^post XXX challenge|Norepinephrine^post XXX challenge
C2736080|T201|COMP|57664-5|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2736081|T201|COMP|57665-2|LNC|Protein fractions.oligoclonal bands.IgG|Protein fractions.oligoclonal bands.IgG
C2736082|T201|COMP|57666-0|LNC|Protein fractions.oligoclonal bands.IgM|Protein fractions.oligoclonal bands.IgM
C2736083|T201|COMP|57674-4|LNC|Coxiella burnetii Ab.IgM^2nd specimen|Coxiella burnetii Ab.IgM^2nd specimen
C2736084|T201|COMP|57675-1|LNC|Legionella pneumophila Ab.IgG^1st specimen|Legionella pneumophila Ab.IgG^1st specimen
C2736085|T201|COMP|57676-9|LNC|Legionella pneumophila Ab.IgG^2nd specimen|Legionella pneumophila Ab.IgG^2nd specimen
C2736086|T201|COMP|57677-7|LNC|Mycoplasma pneumoniae Ab.IgG^1st specimen|Mycoplasma pneumoniae Ab.IgG^1st specimen
C2736087|T201|COMP|57678-5|LNC|Mycoplasma pneumoniae Ab.IgG^2nd specimen|Mycoplasma pneumoniae Ab.IgG^2nd specimen
C2736088|T201|COMP|57679-3|LNC|Chlamydia sp Ab.IgG^1st specimen|Chlamydia sp Ab.IgG^1st specimen
C2736089|T201|COMP|57680-1|LNC|Chlamydia sp Ab.IgG^2nd specimen|Chlamydia sp Ab.IgG^2nd specimen
C2736090|T201|COMP|57681-9|LNC|Coxiella burnetii Ab.IgG^1st specimen|Coxiella burnetii Ab.IgG^1st specimen
C2736091|T201|COMP|57682-7|LNC|Coxiella burnetii Ab.IgG^2nd specimen|Coxiella burnetii Ab.IgG^2nd specimen
C2736092|T201|COMP|57683-5|LNC|Plasmodium falciparum Ab.IgM|Plasmodium falciparum Ab.IgM
C2736093|T201|COMP|57684-3|LNC|Cortisol^11th specimen|Cortisol^11th specimen
C2736094|T201|COMP|57685-0|LNC|Cortisol^2nd specimen|Cortisol^2nd specimen
C2736095|T201|COMP|57686-8|LNC|Cortisol^12th specimen|Cortisol^12th specimen
C2736096|T201|COMP|57687-6|LNC|Cortisol^1st specimen|Cortisol^1st specimen
C2736097|T201|COMP|57688-4|LNC|Cortisol^3rd specimen|Cortisol^3rd specimen
C2736098|T201|COMP|57689-2|LNC|Cortisol^4th specimen|Cortisol^4th specimen
C2736099|T201|COMP|57690-0|LNC|Cortisol^10th specimen|Cortisol^10th specimen
C2736100|T201|COMP|57691-8|LNC|Cortisol^9th specimen|Cortisol^9th specimen
C2736101|T201|COMP|57692-6|LNC|Cortisol^5th specimen|Cortisol^5th specimen
C2736102|T201|COMP|57693-4|LNC|Cortisol^6th specimen|Cortisol^6th specimen
C2736103|T201|COMP|57694-2|LNC|Cortisol^7th specimen|Cortisol^7th specimen
C2736104|T201|COMP|57695-9|LNC|Cortisol^8th specimen|Cortisol^8th specimen
C2736106|T201|COMP|57697-5|LNC|Protein Z Ag|Protein Z Ag
C2736108|T201|COMP|57698-3|LNC|Lipid panel with direct LDL|Lipid panel with direct LDL
C2736117|T201|COMP|57716-3|LNC|State printed on filter paper card|State printed on filter paper card
C2736120|T201|COMP|57717-1|LNC|Newborn screen card data panel|Newborn screen card data panel
C2736122|T201|COMP|57718-9|LNC|Sample condition|Sample condition
C2736126|T201|COMP|57720-5|LNC|Newborn conditions with equivocal markers|Newborn conditions with equivocal markers
C2736128|T201|COMP|57721-3|LNC|Reason for lab test|Reason for lab test
C2736132|T201|COMP|57723-9|LNC|Unique bar code number|Unique bar code number
C2736134|T201|COMP|57724-7|LNC|Newborn screening short narrative summary|Newborn screening short narrative summary
C2736136|T201|COMP|57725-4|LNC|Corticotropin^20M post XXX challenge|Corticotropin^20M post XXX challenge
C2736137|T201|COMP|57726-2|LNC|Creatinine|Creatinine
C2736138|T201|COMP|57727-0|LNC|Norolanzapine|Norolanzapine
C2736140|T201|COMP|57728-8|LNC|Lactate^40M post XXX challenge|Lactate^40M post XXX challenge
C2736141|T201|COMP|57729-6|LNC|Lactate^6M post XXX challenge|Lactate^6M post XXX challenge
C2736142|T201|COMP|57731-2|LNC|Osmolality^2nd specimen|Osmolality^2nd specimen
C2736143|T201|COMP|57732-0|LNC|Osmolality^3rd specimen|Osmolality^3rd specimen
C2736144|T201|COMP|57733-8|LNC|Beta-trace protein|Beta-trace protein
C2736145|T201|COMP|57734-6|LNC|Ketones|Ketones
C2736146|T201|COMP|57735-3|LNC|Protein|Protein
C2736147|T201|COMP|57736-1|LNC|Cells.CD154/100 cells|Cells.CD154/100 cells
C2736149|T201|COMP|57737-9|LNC|Basement membrane Ab|Basement membrane Ab
C2736150|T201|COMP|57738-7|LNC|Basement membrane zone BP180 Ab|Basement membrane zone BP180 Ab
C2736151|T201|COMP|57739-5|LNC|Centromere Ab|Centromere Ab
C2736152|T201|COMP|57740-3|LNC|Cells.CD3+HLA-DR+/100 cells|Cells.CD3+HLA-DR+/100 cells
C2736153|T201|COMP|57741-1|LNC|Lymphocyte proliferation.OKT3 stimulation|Lymphocyte proliferation.OKT3 stimulation
C2736155|T201|COMP|57742-9|LNC|Phadiatop Infant Ab.IgE|Phadiatop Infant Ab.IgE
C2736157|T201|COMP|57743-7|LNC|ABO group|ABO group
C2736158|T201|COMP|57744-5|LNC|Striated muscle Ab|Striated muscle Ab
C2736159|T201|COMP|57745-2|LNC|Adrenal Ab|Adrenal Ab
C2736160|T201|COMP|57746-0|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C2736161|T201|COMP|57747-8|LNC|Erythrocytes|Erythrocytes
C2736162|T201|COMP|57748-6|LNC|Liver cytosol Ab|Liver cytosol Ab
C2736163|T201|COMP|57749-4|LNC|Amphiphysin Ab|Amphiphysin Ab
C2736164|T201|COMP|57750-2|LNC|Amphiphysin Ab|Amphiphysin Ab
C2736165|T201|COMP|57751-0|LNC|Hemoglobin|Hemoglobin
C2736166|T201|COMP|57752-8|LNC|Urea^overnight|Urea^overnight
C2736167|T201|COMP|57753-6|LNC|IKBKG gene targeted mutation analysis|IKBKG gene targeted mutation analysis
C2736169|T201|COMP|57754-4|LNC|TNFRSF13B gene mutations tested for|TNFRSF13B gene mutations tested for
C2736171|T201|COMP|57755-1|LNC|WAS gene mutations tested for|WAS gene mutations tested for
C2736173|T201|COMP|57756-9|LNC|Procollagen type III.N-terminal propeptide|Procollagen type III.N-terminal propeptide
C2736175|T201|COMP|57757-7|LNC|IKBKG gene mutations tested for|IKBKG gene mutations tested for
C2736177|T201|COMP|57758-5|LNC|TNFRSF13B gene targeted mutation analysis|TNFRSF13B gene targeted mutation analysis
C2736179|T201|COMP|57759-3|LNC|WAS gene targeted mutation analysis|WAS gene targeted mutation analysis
C2736181|T201|COMP|57760-1|LNC|Coagulation factor XIII inhibitor|Coagulation factor XIII inhibitor
C2736182|T201|COMP|57761-9|LNC|Platelet factor 4 heparin complex induced Ab|Platelet factor 4 heparin complex induced Ab
C2736183|T201|COMP|57762-7|LNC|Cells.CD55+CD59|Cells.CD55+CD59
C2736186|T201|COMP|57764-3|LNC|Microscopic exam|Microscopic exam
C2736187|T201|COMP|57765-0|LNC|Disaccharidases panel|Disaccharidases panel
C2736189|T201|COMP|57766-8|LNC|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C2736190|T201|COMP|57767-6|LNC|Trimipramine & Nortrimipramine panel|Trimipramine & Nortrimipramine panel
C2736192|T201|COMP|57768-4|LNC|Campylobacter jejuni+Campylobacter coli Ag|Campylobacter jejuni+Campylobacter coli Ag
C2736194|T201|COMP|57769-2|LNC|Salmonella typhi O Vi Ab|Salmonella typhi O Vi Ab
C2736196|T201|COMP|57777-5|LNC|Myeloperoxidase Ab & Proteinase 3 panel|Myeloperoxidase Ab & Proteinase 3 panel
C2736198|T201|COMP|57778-3|LNC|Immunoglobulin light chains.free panel|Immunoglobulin light chains.free panel
C2736200|T201|COMP|57779-1|LNC|Disaccharidases|Disaccharidases
C2736201|T201|COMP|57780-9|LNC|Thyroglobulin & Thyrogobulin Ab panel|Thyroglobulin & Thyrogobulin Ab panel
C2736203|T201|COMP|57781-7|LNC|Chromosome breakage|Chromosome breakage
C2736204|T201|COMP|57782-5|LNC|CBC W Ordered Manual Differential panel|CBC W Ordered Manual Differential panel
C2736210|T201|COMP|57787-4|LNC|Dehydroepiandrosterone^pre dose dexamethasone|Dehydroepiandrosterone^pre dose dexamethasone
C2736211|T201|COMP|57788-2|LNC|Dehydroepiandrosterone^pre dose dexamethasone|Dehydroepiandrosterone^pre dose dexamethasone
C2736212|T201|COMP|57789-0|LNC|Dehydroepiandrosterone^2D post dose dexamethasone|Dehydroepiandrosterone^2D post dose dexamethasone
C2736213|T201|COMP|57790-8|LNC|Dehydroepiandrosterone^2D post dose dexamethasone|Dehydroepiandrosterone^2D post dose dexamethasone
C2736214|T201|COMP|57791-6|LNC|Organic acidemia conditions suspected|Organic acidemia conditions suspected
C2736216|T201|COMP|57792-4|LNC|Fatty acid oxidation conditions suspected|Fatty acid oxidation conditions suspected
C2736218|T201|COMP|57793-2|LNC|Amino acidemia disorder suspected|Amino acidemia disorder suspected
C2736246|T201|COMP|57820-3|LNC|HEDIS 2010 panel|HEDIS 2010 panel
C2736259|T201|COMP|57835-1|LNC|Appearance|Appearance
C2736260|T201|COMP|57837-7|LNC|Beta-1 transferrin|Beta-1 transferrin
C2736263|T201|COMP|57839-3|LNC|Activated clotting time|Activated clotting time
C2736264|T201|COMP|57841-9|LNC|Erythrocytes|Erythrocytes
C2736265|T201|COMP|57842-7|LNC|Erythrocytes|Erythrocytes
C2736266|T201|COMP|57843-5|LNC|Erythrocytes|Erythrocytes
C2736267|T201|COMP|57844-3|LNC|Imatinib mesylate|Imatinib mesylate
C2736268|T201|COMP|57845-0|LNC|Leukocytes|Leukocytes
C2736269|T201|COMP|57846-8|LNC|Leukocytes|Leukocytes
C2736270|T201|COMP|57847-6|LNC|Leukocytes|Leukocytes
C2736271|T201|COMP|57848-4|LNC|Maltose|Maltose
C2736275|T201|COMP|57853-4|LNC|Snowshoe hare virus Ab.IgG|Snowshoe hare virus Ab.IgG
C2736277|T201|COMP|57854-2|LNC|Thyrotropin^5M post XXX challenge|Thyrotropin^5M post XXX challenge
C2736278|T201|COMP|57855-9|LNC|Atenolol|Atenolol
C2736279|T201|COMP|57856-7|LNC|Carisoprodol|Carisoprodol
C2736280|T201|COMP|57857-5|LNC|Chlorpheniramine|Chlorpheniramine
C2736281|T201|COMP|57858-3|LNC|Normaprotiline|Normaprotiline
C2736282|T201|COMP|57859-1|LNC|Dextromethorphan|Dextromethorphan
C2736283|T201|COMP|57860-9|LNC|Diethylamine|Diethylamine
C2736284|T201|COMP|57861-7|LNC|HYDROcodone|HYDROcodone
C2736285|T201|COMP|57862-5|LNC|Hydrocortisone|Hydrocortisone
C2736286|T201|COMP|57863-3|LNC|HYDROmorphone|HYDROmorphone
C2736287|T201|COMP|57864-1|LNC|Meperidine|Meperidine
C2736288|T201|COMP|57865-8|LNC|oxyCODONE|oxyCODONE
C2736289|T201|COMP|57866-6|LNC|PENTobarbital|PENTobarbital
C2736290|T201|COMP|57867-4|LNC|Pericyazine|Pericyazine
C2736291|T201|COMP|57868-2|LNC|Perphenazine|Perphenazine
C2736292|T201|COMP|57869-0|LNC|Phencyclidine|Phencyclidine
C2736293|T201|COMP|57870-8|LNC|Phenylpropanolamine|Phenylpropanolamine
C2736294|T201|COMP|57871-6|LNC|quiNINE|quiNINE
C2736295|T201|COMP|57872-4|LNC|Strychnine|Strychnine
C2736296|T201|COMP|57873-2|LNC|Thiothixene|Thiothixene
C2736297|T201|COMP|57874-0|LNC|Cucumis melo cantalupensis basophil bound Ab|Cucumis melo cantalupensis basophil bound Ab
C2736299|T201|COMP|57875-7|LNC|Cucumis melo cantalupensis Ab.IgG4|Cucumis melo cantalupensis Ab.IgG4
C2736301|T201|COMP|57876-5|LNC|Cucumis melo spp Ab.IgG4|Cucumis melo spp Ab.IgG4
C2736302|T201|COMP|57877-3|LNC|Cucumis melo cantalupensis Ab.IgG.RAST class|Cucumis melo cantalupensis Ab.IgG.RAST class
C2736304|T201|COMP|57878-1|LNC|Cucumis melo spp Ab.IgG.RAST class|Cucumis melo spp Ab.IgG.RAST class
C2736305|T201|COMP|57879-9|LNC|Cucumis melo cantalupensis Ab.IgG|Cucumis melo cantalupensis Ab.IgG
C2736307|T201|COMP|57881-5|LNC|Cucumis melo cantalupensis Ab.IgE.RAST class|Cucumis melo cantalupensis Ab.IgE.RAST class
C2736309|T201|COMP|57883-1|LNC|Cucumis melo cantalupensis Ab.IgE|Cucumis melo cantalupensis Ab.IgE
C2736311|T201|COMP|57885-6|LNC|Cucumis melo spp basophil bound Ab|Cucumis melo spp basophil bound Ab
C2736312|T201|COMP|57886-4|LNC|Pregnanediol^pre high dose dexamethasone|Pregnanediol^pre high dose dexamethasone
C2736313|T201|COMP|57887-2|LNC|Pregnanediol^pre high dose dexamethasone|Pregnanediol^pre high dose dexamethasone
C2736314|T201|COMP|57888-0|LNC|Pregnanediol^2D post high dose dexamethasone|Pregnanediol^2D post high dose dexamethasone
C2736315|T201|COMP|57889-8|LNC|Pregnanediol^2D post high dose dexamethasone|Pregnanediol^2D post high dose dexamethasone
C2736316|T201|COMP|57890-6|LNC|Pregnanediol^pre dose dexamethasone|Pregnanediol^pre dose dexamethasone
C2736317|T201|COMP|57891-4|LNC|Pregnanediol^pre dose dexamethasone|Pregnanediol^pre dose dexamethasone
C2736318|T201|COMP|57892-2|LNC|Pregnanediol^2D post dose dexamethasone|Pregnanediol^2D post dose dexamethasone
C2736319|T201|COMP|57893-0|LNC|Pregnanediol^2D post dose dexamethasone|Pregnanediol^2D post dose dexamethasone
C2736320|T201|COMP|57894-8|LNC|C peptide^100M post XXX challenge|C peptide^100M post XXX challenge
C2736327|T201|COMP|57898-9|LNC|Cocaine|Cocaine
C2736328|T201|COMP|57899-7|LNC|Triiodothyronine/Triiodothyronine.reverse|Triiodothyronine/Triiodothyronine.reverse
C2736330|T201|COMP|57900-3|LNC|Specimen age|Specimen age
C2736331|T201|COMP|57901-1|LNC|Clostridioides difficile glutamate dehydrogenase|Clostridioides difficile glutamate dehydrogenase
C2736333|T201|COMP|57902-9|LNC|B little g super little a Ab|B little g super little a Ab
C2736335|T201|COMP|57903-7|LNC|B little g super little a Ab|B little g super little a Ab
C2736336|T201|COMP|57904-5|LNC|B little g super little a Ag|B little g super little a Ag
C2736338|T201|COMP|57905-2|LNC|Hemoglobin.gastrointestinal.lower^1st specimen|Hemoglobin.gastrointestinal.lower^1st specimen
C2736339|T201|COMP|57907-8|LNC|Atazanavir+Ritonavir|Atazanavir+Ritonavir
C2736340|T201|COMP|57908-6|LNC|AIRE gene targeted mutation analysis|AIRE gene targeted mutation analysis
C2736342|T201|COMP|57909-4|LNC|ADNFLE gene targeted mutation analysis|ADNFLE gene targeted mutation analysis
C2736344|T201|COMP|57910-2|LNC|Bartonella quintana DNA|Bartonella quintana DNA
C2736345|T201|COMP|57911-0|LNC|Basement membrane zone BP230 Ab|Basement membrane zone BP230 Ab
C2736346|T201|COMP|57916-9|LNC|Borrelia burgdorferi C6 Ab|Borrelia burgdorferi C6 Ab
C2736347|T201|COMP|57917-7|LNC|Budgerigar droppings Ab.IgG|Budgerigar droppings Ab.IgG
C2736348|T201|COMP|57918-5|LNC|CACNA1S+SCN4A gene targeted mutation analysis|CACNA1S+SCN4A gene targeted mutation analysis
C2736350|T201|COMP|57919-3|LNC|Calcium|Calcium
C2736351|T201|COMP|57920-1|LNC|Carbon dioxide|Carbon dioxide
C2736352|T201|COMP|57921-9|LNC|Carbon dioxide|Carbon dioxide
C2736353|T201|COMP|57922-7|LNC|Carbon dioxide|Carbon dioxide
C2736354|T201|COMP|57923-5|LNC|Carbon dioxide|Carbon dioxide
C2736355|T201|COMP|57924-3|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C2736356|T201|COMP|57927-6|LNC|CDKN2A+CDK4 gene targeted mutation analysis|CDKN2A+CDK4 gene targeted mutation analysis
C2736358|T201|COMP|57930-0|LNC|CFTR gene.p.Asp1152His|CFTR gene.p.Asp1152His
C2736360|T201|COMP|57931-8|LNC|CFTR+PRSS1+SPINK1 gene targeted mutation analysis|CFTR+PRSS1+SPINK1 gene targeted mutation analysis
C2736362|T201|COMP|57942-5|LNC|Cladosporium sp Ab.IgG4|Cladosporium sp Ab.IgG4
C2736364|T201|COMP|57943-3|LNC|Clenbuterol|Clenbuterol
C2736365|T201|COMP|57944-1|LNC|Cobalt|Cobalt
C2736366|T201|COMP|57945-8|LNC|Cocaethylene|Cocaethylene
C2736367|T201|COMP|57946-6|LNC|Coccidioides immitis Ab.IgG|Coccidioides immitis Ab.IgG
C2736368|T201|COMP|57948-2|LNC|Collagen crosslinked C-telopeptide|Collagen crosslinked C-telopeptide
C2736369|T201|COMP|57949-0|LNC|Complement C4c|Complement C4c
C2736370|T201|COMP|57951-6|LNC|CPVT1 gene targeted mutation analysis|CPVT1 gene targeted mutation analysis
C2736372|T201|COMP|57953-2|LNC|Ethisterone|Ethisterone
C2736373|T201|COMP|57954-0|LNC|Darunavir|Darunavir
C2736374|T201|COMP|57955-7|LNC|Darunavir+Ritonavir|Darunavir+Ritonavir
C2736375|T201|COMP|57956-5|LNC|DesoxymethylTESTOSTERone|DesoxymethylTESTOSTERone
C2736377|T201|COMP|57957-3|LNC|Difenacoum|Difenacoum
C2736378|T201|COMP|57958-1|LNC|DPYD2A gene targeted mutation analysis|DPYD2A gene targeted mutation analysis
C2736380|T201|COMP|57959-9|LNC|Drostanolone|Drostanolone
C2736381|T201|COMP|57960-7|LNC|Erythrocytes|Erythrocytes
C2736382|T201|COMP|57961-5|LNC|Etravirine|Etravirine
C2736383|T201|COMP|57962-3|LNC|FECH gene targeted mutation analysis|FECH gene targeted mutation analysis
C2736385|T201|COMP|57963-1|LNC|FLCN gene targeted mutation analysis|FLCN gene targeted mutation analysis
C2736387|T201|COMP|57964-9|LNC|Formebolone metabolite|Formebolone metabolite
C2736389|T201|COMP|57965-6|LNC|Fosamprenavir+Ritonavir|Fosamprenavir+Ritonavir
C2736390|T201|COMP|57966-4|LNC|Furazabol metabolite|Furazabol metabolite
C2736392|T201|COMP|57967-2|LNC|Galactitol|Galactitol
C2736393|T201|COMP|57968-0|LNC|Ganglioside GD1a Ab.IgG|Ganglioside GD1a Ab.IgG
C2736394|T201|COMP|57969-8|LNC|Ganglioside GD1a Ab.IgM|Ganglioside GD1a Ab.IgM
C2736395|T201|COMP|57970-6|LNC|Glucose^3H post 75 g glucose PO|Glucose^3H post 75 g glucose PO
C2736396|T201|COMP|57971-4|LNC|Glucose^4th specimen post dose lactose|Glucose^4th specimen post dose lactose
C2736397|T201|COMP|57972-2|LNC|Glucose^5th specimen post dose lactose|Glucose^5th specimen post dose lactose
C2736398|T201|COMP|57973-0|LNC|Histoplasma capsulatum Ab.IgM|Histoplasma capsulatum Ab.IgM
C2736399|T201|COMP|57974-8|LNC|HIV 1 Ab|HIV 1 Ab
C2736400|T201|COMP|57975-5|LNC|HIV 1+O+2 Ab|HIV 1+O+2 Ab
C2736401|T201|COMP|57976-3|LNC|HIV 2 gp140 Ab|HIV 2 gp140 Ab
C2736403|T201|COMP|57977-1|LNC|HIV 2 p16 Ab|HIV 2 p16 Ab
C2736405|T201|COMP|57978-9|LNC|HIV 2 p34 Ab|HIV 2 p34 Ab
C2736407|T201|COMP|57979-7|LNC|HLA-B*15:02|HLA-B*15:02
C2736408|T201|COMP|57980-5|LNC|HLA-B51|HLA-B51
C2736409|T201|COMP|57981-3|LNC|HYDROcodone|HYDROcodone
C2736410|T201|COMP|57982-1|LNC|HYDROmorphone|HYDROmorphone
C2736411|T201|COMP|57983-9|LNC|IDUA gene targeted mutation analysis|IDUA gene targeted mutation analysis
C2736413|T201|COMP|57984-7|LNC|Indinavir+Ritonavir|Indinavir+Ritonavir
C2736414|T201|COMP|57985-4|LNC|Influenza virus A H2 RNA|Influenza virus A H2 RNA
C2736417|T201|COMP|57988-8|LNC|Iron|Iron
C2736418|T201|COMP|57990-4|LNC|KRIT1 gene targeted mutation analysis|KRIT1 gene targeted mutation analysis
C2736420|T201|COMP|57992-0|LNC|Legionella pneumophila 1+3+4+5+6+8 Ab|Legionella pneumophila 1+3+4+5+6+8 Ab
C2736421|T201|COMP|57994-6|LNC|Leucine/Alanine|Leucine/Alanine
C2736423|T201|COMP|57995-3|LNC|Leucine/Phenylalanine|Leucine/Phenylalanine
C2736425|T201|COMP|57996-1|LNC|Leucine+Isoleucine|Leucine+Isoleucine
C2736426|T201|COMP|57997-9|LNC|Lopinavir+Ritonavir|Lopinavir+Ritonavir
C2736427|T201|COMP|57998-7|LNC|Magnesium|Magnesium
C2736428|T201|COMP|57999-5|LNC|Manganese|Manganese
C2736429|T201|COMP|58001-9|LNC|Matrix metallopeptidase 9|Matrix metallopeptidase 9
C2736431|T201|COMP|58002-7|LNC|Mestanolone metabolite|Mestanolone metabolite
C2736433|T201|COMP|58003-5|LNC|Methylandrostenediol|Methylandrostenediol
C2736434|T201|COMP|58004-3|LNC|Methasterone|Methasterone
C2736436|T201|COMP|58005-0|LNC|Methylnortestosterone|Methylnortestosterone
C2736437|T201|COMP|58006-8|LNC|Mibolerone|Mibolerone
C2736438|T201|COMP|58008-4|LNC|Morus alba Ab.IgG.RAST class|Morus alba Ab.IgG.RAST class
C2736440|T201|COMP|58009-2|LNC|MPL gene.p.Trp515|MPL gene.p.Trp515
C2736444|T201|COMP|58011-8|LNC|Myelin Ab.IgG|Myelin Ab.IgG
C2736445|T201|COMP|58012-6|LNC|Natalizumab Ab|Natalizumab Ab
C2736446|T201|COMP|58013-4|LNC|Norclomipramine|Norclomipramine
C2736447|T201|COMP|58014-2|LNC|Nordoxepin|Nordoxepin
C2736448|T201|COMP|58015-9|LNC|Nortrimipramine|Nortrimipramine
C2736449|T201|COMP|58016-7|LNC|Octreotide|Octreotide
C2736450|T201|COMP|58018-3|LNC|Oxabolone|Oxabolone
C2736452|T201|COMP|58019-1|LNC|Phosphate|Phosphate
C2736453|T201|COMP|58020-9|LNC|PKD2 gene targeted mutation analysis|PKD2 gene targeted mutation analysis
C2736455|T201|COMP|58021-7|LNC|Populus deltoides Ab.IgG.RAST class|Populus deltoides Ab.IgG.RAST class
C2736457|T201|COMP|58022-5|LNC|Prostanozol|Prostanozol
C2736459|T201|COMP|58023-3|LNC|Rabies virus Ab.IgG|Rabies virus Ab.IgG
C2736460|T201|COMP|58024-1|LNC|Saquinavir+Ritonavir|Saquinavir+Ritonavir
C2736461|T201|COMP|58026-6|LNC|Selenium|Selenium
C2736462|T201|COMP|58027-4|LNC|Testolactone|Testolactone
C2736463|T201|COMP|58028-2|LNC|Tetrahydrogestrinone|Tetrahydrogestrinone
C2736464|T201|COMP|58029-0|LNC|Tipranavir+Ritonavir|Tipranavir+Ritonavir
C2736465|T201|COMP|58030-8|LNC|Tranylcypromine|Tranylcypromine
C2736466|T201|COMP|58031-6|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C2736467|T201|COMP|58032-4|LNC|Ulmus americana Ab.IgG|Ulmus americana Ab.IgG
C2736468|T201|COMP|58035-7|LNC|Vaccinium myrtillus Ab.IgG|Vaccinium myrtillus Ab.IgG
C2736469|T201|COMP|58036-5|LNC|Xanthine/Total|Xanthine/Total
C2736470|T201|COMP|58037-3|LNC|Zinc|Zinc
C2736471|T201|COMP|58038-1|LNC|Gestrinone|Gestrinone
C2736472|T201|COMP|58039-9|LNC|HLA-B SBT|HLA-B SBT
C2736473|T201|COMP|58041-5|LNC|Norclostebol|Norclostebol
C2736474|T201|COMP|58042-3|LNC|Phencyclidine|Phencyclidine
C2736475|T201|COMP|58044-9|LNC|RYR1 gene targeted mutation analysis|RYR1 gene targeted mutation analysis
C2736477|T201|COMP|58045-6|LNC|SCN4A gene targeted mutation analysis|SCN4A gene targeted mutation analysis
C2736479|T201|COMP|58046-4|LNC|Strongyloides stercoralis Ab|Strongyloides stercoralis Ab
C2736480|T201|COMP|58047-2|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C2736486|T201|COMP|58053-0|LNC|C little h super little a Ag|C little h super little a Ag
C2736488|T201|COMP|58054-8|LNC|C little h super little a Ab|C little h super little a Ab
C2736490|T201|COMP|58055-5|LNC|C little o super little a Ag|C little o super little a Ag
C2736492|T201|COMP|58056-3|LNC|C little o super little b Ag|C little o super little b Ag
C2736494|T201|COMP|58057-1|LNC|C little s super little a Ab|C little s super little a Ab
C2736496|T201|COMP|58058-9|LNC|C little s super little a Ag|C little s super little a Ag
C2736498|T201|COMP|58059-7|LNC|D little o super little b Ab|D little o super little b Ab
C2736500|T201|COMP|58060-5|LNC|D little o super little b Ag|D little o super little b Ag
C2736502|T201|COMP|58061-3|LNC|G little o super little a Ab|G little o super little a Ab
C2736504|T201|COMP|58062-1|LNC|I little n super little b Ag|I little n super little b Ag
C2736506|T201|COMP|58063-9|LNC|I little n super little b Ab|I little n super little b Ab
C2736508|T201|COMP|58064-7|LNC|J little r super little a Ag|J little r super little a Ag
C2736510|T201|COMP|58065-4|LNC|J little r super little a Ab|J little r super little a Ab
C2736512|T201|COMP|58066-2|LNC|K little n super little a Ag|K little n super little a Ag
C2736514|T201|COMP|58067-0|LNC|K little n super little a Ab|K little n super little a Ab
C2736516|T201|COMP|58068-8|LNC|K little n super little b Ab|K little n super little b Ab
C2736518|T201|COMP|58069-6|LNC|K little n super little b Ag|K little n super little b Ag
C2736520|T201|COMP|58070-4|LNC|M little c C super little a Ab|M little c C super little a Ab
C2736522|T201|COMP|58071-2|LNC|R little g super little a Ag|R little g super little a Ag
C2736524|T201|COMP|58072-0|LNC|R little g super little a Ab|R little g super little a Ab
C2736526|T201|COMP|58073-8|LNC|W little r super little a Ag|W little r super little a Ag
C2736528|T201|COMP|58074-6|LNC|W little r super little a Ab|W little r super little a Ab
C2736530|T201|COMP|58075-3|LNC|Y little k super little a Ag|Y little k super little a Ag
C2736532|T201|COMP|58076-1|LNC|Y little k super little a Ab|Y little k super little a Ab
C2736534|T201|COMP|58077-9|LNC|Urinalysis complete W Reflex Culture panel|Urinalysis complete W Reflex Culture panel
C2736536|T201|COMP|58078-7|LNC|IH Ab|IH Ab
C2736538|T201|COMP|58079-5|LNC|JMH Ab|JMH Ab
C2736540|T201|COMP|58080-3|LNC|Penicillin.parenteral|Penicillin.parenteral
C2736541|T201|COMP|58081-1|LNC|Vel Ab|Vel Ab
C2736543|T201|COMP|58082-9|LNC|Vel Ag|Vel Ag
C2736571|T201|COMP|58083-7|LNC|Vw Ag|Vw Ag
C2736573|T201|COMP|58084-5|LNC|Vw Ab|Vw Ab
C2736575|T201|COMP|58085-2|LNC|Penicillin.parenteral|Penicillin.parenteral
C2736576|T201|COMP|58086-0|LNC|NOS Ab|NOS Ab
C2736577|T201|COMP|58087-8|LNC|NOS Ab|NOS Ab
C2736578|T201|COMP|58088-6|LNC|Acylcarnitine|Acylcarnitine
C2736579|T201|COMP|58089-4|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C2738953|T201|COMP|56307-2|LNC|Lactuca sativa Ab.IgG4|Lactuca sativa Ab.IgG4
C2738954|T201|COMP|56308-0|LNC|Phaseolus limensis Ab.IgG4|Phaseolus limensis Ab.IgG4
C2738955|T201|COMP|56309-8|LNC|Citrus aurantifolia Ab.IgG4|Citrus aurantifolia Ab.IgG4
C2738956|T201|COMP|56310-6|LNC|Homarus gammarus Ab.IgG4|Homarus gammarus Ab.IgG4
C2738957|T201|COMP|56311-4|LNC|Locust tree Ab.IgG4|Locust tree Ab.IgG4
C2738958|T201|COMP|56312-2|LNC|Malt Ab.IgG4|Malt Ab.IgG4
C2738959|T201|COMP|56313-0|LNC|Mangifera indica Ab.IgG4|Mangifera indica Ab.IgG4
C2738960|T201|COMP|56314-8|LNC|Maple syrup Ab.IgG4|Maple syrup Ab.IgG4
C2738961|T201|COMP|56315-5|LNC|Acer negundo Ab.IgG4|Acer negundo Ab.IgG4
C2738962|T201|COMP|56316-3|LNC|Iva ciliata Ab.IgG4|Iva ciliata Ab.IgG4
C2738963|T201|COMP|56317-1|LNC|Festuca elatior Ab.IgG4|Festuca elatior Ab.IgG4
C2738964|T201|COMP|57323-8|LNC|Varicella zoster virus Ab.IgM^2nd specimen|Varicella zoster virus Ab.IgM^2nd specimen
C2738965|T201|COMP|57324-6|LNC|Influenza virus A Ab.IgG^1st specimen|Influenza virus A Ab.IgG^1st specimen
C2738966|T201|COMP|57325-3|LNC|Influenza virus A Ab.IgG^2nd specimen|Influenza virus A Ab.IgG^2nd specimen
C2738967|T201|COMP|57326-1|LNC|Influenza virus A Ab.IgM^1st specimen|Influenza virus A Ab.IgM^1st specimen
C2738968|T201|COMP|57327-9|LNC|Influenza virus A Ab.IgM^2nd specimen|Influenza virus A Ab.IgM^2nd specimen
C2738969|T201|COMP|57328-7|LNC|Influenza virus B Ab.IgM^1st specimen|Influenza virus B Ab.IgM^1st specimen
C2738970|T201|COMP|57329-5|LNC|Influenza virus B Ab.IgM^2nd specimen|Influenza virus B Ab.IgM^2nd specimen
C2738971|T201|COMP|57330-3|LNC|Corticotropin^40M post XXX challenge|Corticotropin^40M post XXX challenge
C2738972|T201|COMP|57332-9|LNC|Urate|Urate
C2738973|T201|COMP|57333-7|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C2739408|T201|COMP|55944-3|LNC|Neopterin|Neopterin
C2739409|T201|COMP|55945-0|LNC|Neopterin|Neopterin
C2739410|T201|COMP|55946-8|LNC|Neopterin|Neopterin
C2739411|T201|COMP|55947-6|LNC|Nitrite|Nitrite
C2739412|T201|COMP|55948-4|LNC|Nitrite|Nitrite
C2739413|T201|COMP|55949-2|LNC|Dicarboxystearoylcarnitine (C18-DC)|Dicarboxystearoylcarnitine (C18-DC)
C2739414|T201|COMP|55950-0|LNC|Octanoylcarnitine (C8)|Octanoylcarnitine (C8)
C2739415|T201|COMP|55951-8|LNC|Octenoylcarnitine (C8:1)/Creatinine|Octenoylcarnitine (C8:1)/Creatinine
C2739417|T201|COMP|55952-6|LNC|Octenoylcarnitine (C8:1)|Octenoylcarnitine (C8:1)
C2739418|T201|COMP|55953-4|LNC|Octenoylcarnitine (C8:1)|Octenoylcarnitine (C8:1)
C2739419|T201|COMP|55954-2|LNC|Octenoylcarnitine (C8:1)|Octenoylcarnitine (C8:1)
C2739420|T201|COMP|55955-9|LNC|Oleoylcarnitine (C18:1)/Creatinine|Oleoylcarnitine (C18:1)/Creatinine
C2739422|T201|COMP|55956-7|LNC|Oleoylcarnitine (C18:1)|Oleoylcarnitine (C18:1)
C2739423|T201|COMP|55957-5|LNC|Oleoylcarnitine (C18:1)|Oleoylcarnitine (C18:1)
C2739424|T201|COMP|55958-3|LNC|Oleoylcarnitine (C18:1)|Oleoylcarnitine (C18:1)
C2739425|T201|COMP|55959-1|LNC|Ornithine/Amino acids.total|Ornithine/Amino acids.total
C2739427|T201|COMP|55960-9|LNC|Osmolality|Osmolality
C2739428|T201|COMP|55961-7|LNC|Oxalate|Oxalate
C2739429|T201|COMP|55962-5|LNC|Oxygen content|Oxygen content
C2739430|T201|COMP|55963-3|LNC|Palmitoleylcarnitine (C16:1)/Creatinine|Palmitoleylcarnitine (C16:1)/Creatinine
C2739432|T201|COMP|55964-1|LNC|Palmitoleylcarnitine (C16:1)|Palmitoleylcarnitine (C16:1)
C2739433|T201|COMP|55965-8|LNC|Palmitoleylcarnitine (C16:1)|Palmitoleylcarnitine (C16:1)
C2739434|T201|COMP|56453-4|LNC|Cow dander Ab.IgG4|Cow dander Ab.IgG4
C2739435|T201|COMP|56454-2|LNC|Cuminum cyminum Ab.IgG4|Cuminum cyminum Ab.IgG4
C2739436|T201|COMP|56455-9|LNC|Gelatin Ab.IgG4|Gelatin Ab.IgG4
C2739438|T201|COMP|56456-7|LNC|Horse dander Ab.IgG4|Horse dander Ab.IgG4
C2739440|T201|COMP|56457-5|LNC|Lamb Ab.IgG4|Lamb Ab.IgG4
C2739441|T201|COMP|56458-3|LNC|Acacia longifolia Ab.IgG4|Acacia longifolia Ab.IgG4
C2739442|T201|COMP|56459-1|LNC|Ustilago avenae Ab.IgG4|Ustilago avenae Ab.IgG4
C2739443|T201|COMP|56460-9|LNC|Schinus molle Ab.IgG4|Schinus molle Ab.IgG4
C2739444|T201|COMP|56461-7|LNC|Alnus rubra Ab.IgG4|Alnus rubra Ab.IgG4
C2739445|T201|COMP|56462-5|LNC|Pepper red Ab.IgG4|Pepper red Ab.IgG4
C2739447|T201|COMP|56463-3|LNC|Pigweed rough Ab.IgG4|Pigweed rough Ab.IgG4
C2739448|T201|COMP|56464-1|LNC|Salvia officinalis Ab.IgG4|Salvia officinalis Ab.IgG4
C2739449|T201|COMP|56594-5|LNC|Thyrotropin^3H post XXX challenge|Thyrotropin^3H post XXX challenge
C2739450|T201|COMP|56595-2|LNC|Latex recombinant (rHev b) 3 Ab.IgE|Latex recombinant (rHev b) 3 Ab.IgE
C2739452|T201|COMP|56596-0|LNC|Latex recombinant (rHev b) 5 Ab.IgE|Latex recombinant (rHev b) 5 Ab.IgE
C2739454|T201|COMP|56597-8|LNC|Latex recombinant (rHev b) 8 Ab.IgE|Latex recombinant (rHev b) 8 Ab.IgE
C2739456|T201|COMP|56598-6|LNC|Epstein Barr virus early Ab.IgM|Epstein Barr virus early Ab.IgM
C2739457|T201|COMP|56599-4|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C2739458|T201|COMP|56600-0|LNC|Vespa crabro Ab.IgG|Vespa crabro Ab.IgG
C2739459|T201|COMP|56601-8|LNC|Hyaluronate|Hyaluronate
C2739462|T201|COMP|56767-7|LNC|Protein.monoclonal.beta|Protein.monoclonal.beta
C2739463|T201|COMP|56768-5|LNC|Protein.monoclonal.beta/Protein.total|Protein.monoclonal.beta/Protein.total
C2739465|T201|COMP|56769-3|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C2739466|T201|COMP|56770-1|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C2739467|T201|COMP|56771-9|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C2739468|T201|COMP|56772-7|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C2739469|T201|COMP|56773-5|LNC|Cells.CD1a/100 cells|Cells.CD1a/100 cells
C2739470|T201|COMP|56774-3|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C2739471|T201|COMP|56775-0|LNC|Cells.CD3-CD16+CD56+|Cells.CD3-CD16+CD56+
C2739472|T201|COMP|56776-8|LNC|Amylase.S3+S4/Amylase.total|Amylase.S3+S4/Amylase.total
C2739474|T201|COMP|56777-6|LNC|Lipoprotein.pre-beta/Lipoprotein.beta|Lipoprotein.pre-beta/Lipoprotein.beta
C2739476|T201|COMP|56986-3|LNC|Thyroxine.free^1H post XXX challenge|Thyroxine.free^1H post XXX challenge
C2739477|T201|COMP|56987-1|LNC|Thyroxine.free^40M post XXX challenge|Thyroxine.free^40M post XXX challenge
C2739478|T201|COMP|56988-9|LNC|Thyroxine.free^1.5H post XXX challenge|Thyroxine.free^1.5H post XXX challenge
C2739479|T201|COMP|56989-7|LNC|Thyroxine.free^20M post XXX challenge|Thyroxine.free^20M post XXX challenge
C2739480|T201|COMP|56990-5|LNC|Toxoplasma gondii Ab.IgG avidity|Toxoplasma gondii Ab.IgG avidity
C2739481|T201|COMP|56991-3|LNC|Toxoplasma gondii Ab.IgG avidity|Toxoplasma gondii Ab.IgG avidity
C2739482|T201|COMP|56992-1|LNC|Trichinella sp Ab.IgG|Trichinella sp Ab.IgG
C2739483|T201|COMP|56993-9|LNC|Tryptophan/Creatinine|Tryptophan/Creatinine
C2739484|T201|COMP|56994-7|LNC|Tyrosine/Creatinine|Tyrosine/Creatinine
C2739485|T201|COMP|56995-4|LNC|Urea|Urea
C2739486|T201|COMP|56996-2|LNC|Urea/Creatinine|Urea/Creatinine
C2739487|T201|COMP|57406-1|LNC|Cells.CD8+CD57+/100 cells|Cells.CD8+CD57+/100 cells
C2739488|T201|COMP|57546-4|LNC|17-Hydroxyprogesterone^pre dose dexamethasone|17-Hydroxyprogesterone^pre dose dexamethasone
C2739489|T201|COMP|57547-2|LNC|17-Hydroxyprogesterone^1D post dose dexamethasone|17-Hydroxyprogesterone^1D post dose dexamethasone
C2739490|T201|COMP|57548-0|LNC|17-Hydroxyprogesterone^1D post dose dexamethasone|17-Hydroxyprogesterone^1D post dose dexamethasone
C2739491|T201|COMP|57549-8|LNC|17-Hydroxyprogesterone^2D post dose dexamethasone|17-Hydroxyprogesterone^2D post dose dexamethasone
C2739492|T201|COMP|57550-6|LNC|17-Hydroxyprogesterone^2D post dose dexamethasone|17-Hydroxyprogesterone^2D post dose dexamethasone
C2739497|T201|COMP|56223-1|LNC|Cinnamomum spp Ab.IgG4|Cinnamomum spp Ab.IgG4
C2739498|T201|COMP|56224-9|LNC|Cladosporium herbarum Ab.IgG4|Cladosporium herbarum Ab.IgG4
C2739499|T201|COMP|56225-6|LNC|Ruditapes spp Ab.IgG4|Ruditapes spp Ab.IgG4
C2739500|T201|COMP|56226-4|LNC|Xanthium commune Ab.IgG4|Xanthium commune Ab.IgG4
C2739501|T201|COMP|56227-2|LNC|Cocos nucifera Ab.IgG4|Cocos nucifera Ab.IgG4
C2739502|T201|COMP|56228-0|LNC|Gadus morhua Ab.IgG4|Gadus morhua Ab.IgG4
C2739503|T201|COMP|56229-8|LNC|Coffea spp Ab.IgG4|Coffea spp Ab.IgG4
C2739504|T201|COMP|56230-6|LNC|Phragmites communis Ab.IgG4|Phragmites communis Ab.IgG4
C2739505|T201|COMP|56383-3|LNC|Salmo salar Ab.IgG4|Salmo salar Ab.IgG4
C2739506|T201|COMP|56384-1|LNC|Sardina pilchardus Ab.IgG4|Sardina pilchardus Ab.IgG4
C2739507|T201|COMP|56385-8|LNC|Pecten spp Ab.IgG4|Pecten spp Ab.IgG4
C2739508|T201|COMP|56386-6|LNC|Sesamum indicum Ab.IgG4|Sesamum indicum Ab.IgG4
C2739509|T201|COMP|56387-4|LNC|Rumex acetosella Ab.IgG4|Rumex acetosella Ab.IgG4
C2739510|T201|COMP|56388-2|LNC|Pandalus borealis Ab.IgG4|Pandalus borealis Ab.IgG4
C2739511|T201|COMP|56389-0|LNC|Solea solea Ab.IgG4|Solea solea Ab.IgG4
C2739512|T201|COMP|56390-8|LNC|Glycine max Ab.IgG4|Glycine max Ab.IgG4
C2739513|T201|COMP|56391-6|LNC|Spinacia oleracea Ab.IgG4|Spinacia oleracea Ab.IgG4
C2739514|T201|COMP|56392-4|LNC|Pigweed spiny Ab.IgG4|Pigweed spiny Ab.IgG4
C2739515|T201|COMP|56393-2|LNC|Fragaria vesca Ab.IgG4|Fragaria vesca Ab.IgG4
C2739516|T201|COMP|56394-0|LNC|Saccharum officinarum Ab.IgG4|Saccharum officinarum Ab.IgG4
C2739517|T201|COMP|56395-7|LNC|Helianthus annuus seed Ab.IgG4|Helianthus annuus seed Ab.IgG4
C2739518|T201|COMP|56396-5|LNC|Castanea sativa Ab.IgG4|Castanea sativa Ab.IgG4
C2739519|T201|COMP|56397-3|LNC|Ipomoea batatas Ab.IgG4|Ipomoea batatas Ab.IgG4
C2739520|T201|COMP|56398-1|LNC|Anthoxanthum odoratum Ab.IgG4|Anthoxanthum odoratum Ab.IgG4
C2739521|T201|COMP|56399-9|LNC|Cheese swiss Ab.IgG4|Cheese swiss Ab.IgG4
C2739522|T201|COMP|55906-2|LNC|Alpha cortolone|Alpha cortolone
C2739523|T201|COMP|55907-0|LNC|Alpha cortolone|Alpha cortolone
C2739524|T201|COMP|55908-8|LNC|Alpha galactosidase A|Alpha galactosidase A
C2739525|T201|COMP|55909-6|LNC|Alpha-L-iduronidase|Alpha-L-iduronidase
C2739526|T201|COMP|55910-4|LNC|Alpha mannosidase|Alpha mannosidase
C2739527|T201|COMP|55911-2|LNC|Arginine|Arginine
C2739528|T201|COMP|55912-0|LNC|Arylsulfatase|Arylsulfatase
C2739529|T201|COMP|55913-8|LNC|Aspartate|Aspartate
C2739537|T201|COMP|56253-8|LNC|Egg white Ab.IgG4|Egg white Ab.IgG4
C2739538|T201|COMP|56254-6|LNC|Egg yolk Ab.IgG4|Egg yolk Ab.IgG4
C2739539|T201|COMP|56255-3|LNC|Egg whole Ab.IgG4|Egg whole Ab.IgG4
C2739540|T201|COMP|56256-1|LNC|Solanum melongena Ab.IgG4|Solanum melongena Ab.IgG4
C2739541|T201|COMP|56257-9|LNC|Plantago lanceolata Ab.IgG4|Plantago lanceolata Ab.IgG4
C2739542|T201|COMP|56258-7|LNC|Eucalyptus spp Ab.IgG4|Eucalyptus spp Ab.IgG4
C2739544|T201|COMP|56260-3|LNC|Solenopsis invicta Ab.IgG4|Solenopsis invicta Ab.IgG4
C2739545|T201|COMP|56413-8|LNC|Quercus virginiana Ab.IgG4|Quercus virginiana Ab.IgG4
C2739546|T201|COMP|56414-6|LNC|Juglans spp Ab.IgG4|Juglans spp Ab.IgG4
C2739547|T201|COMP|56415-3|LNC|Citrullus lanatus Ab.IgG4|Citrullus lanatus Ab.IgG4
C2739548|T201|COMP|56416-1|LNC|Acnida tamariscina Ab.IgG4|Acnida tamariscina Ab.IgG4
C2739549|T201|COMP|56417-9|LNC|Triticum aestivum Ab.IgG4|Triticum aestivum Ab.IgG4
C2739550|T201|COMP|56418-7|LNC|Triticum aestivum pollen Ab.IgG4|Triticum aestivum pollen Ab.IgG4
C2739551|T201|COMP|56419-5|LNC|Cow whey Ab.IgG4|Cow whey Ab.IgG4
C2739552|T201|COMP|56420-3|LNC|Fraxinus americana Ab.IgG4|Fraxinus americana Ab.IgG4
C2739553|T201|COMP|56421-1|LNC|Bean white Ab.IgG4|Bean white Ab.IgG4
C2739554|T201|COMP|56422-9|LNC|Betula populifolia Ab.IgG4|Betula populifolia Ab.IgG4
C2739555|T201|COMP|56423-7|LNC|Carya tomentosa Ab.IgG4|Carya tomentosa Ab.IgG4
C2739556|T201|COMP|56424-5|LNC|Dolichovespula maculata Ab.IgG4|Dolichovespula maculata Ab.IgG4
C2739557|T201|COMP|56425-2|LNC|Morus alba Ab.IgG4|Morus alba Ab.IgG4
C2739558|T201|COMP|56426-0|LNC|Quercus alba Ab.IgG4|Quercus alba Ab.IgG4
C2739559|T201|COMP|56427-8|LNC|Pinus strobus Ab.IgG4|Pinus strobus Ab.IgG4
C2739560|T201|COMP|56428-6|LNC|Populus alba Ab.IgG4|Populus alba Ab.IgG4
C2739561|T201|COMP|55764-5|LNC|EGFR gene exon 19 deletion|EGFR gene exon 19 deletion
C2739562|T201|COMP|55765-2|LNC|EGFR gene.c.2156G>C+2155G>A+2155G>T|EGFR gene.c.2156G>C+2155G>A+2155G>T
C2739563|T201|COMP|55766-0|LNC|EGFR gene.c.2573T>G|EGFR gene.c.2573T>G
C2739805|T201|COMP|35203-9|LNC|Creatinine|Creatinine
C2741668|T201|COMP|57298-2|LNC|HLA-DRB1|HLA-DRB1
C2741675|T201|COMP|56156-3|LNC|Candida albicans Ab.IgA & IgG & IgM panel|Candida albicans Ab.IgA & IgG & IgM panel
C2745875|T201|COMP|56652-1|LNC|Arsenic/Creatinine|Arsenic/Creatinine
C2745876|T201|COMP|56651-3|LNC|Cadmium/Creatinine|Cadmium/Creatinine
C2745893|T201|COMP|56650-5|LNC|Chromium/Creatinine|Chromium/Creatinine
C2745898|T201|COMP|56653-9|LNC|Mercury/Creatinine|Mercury/Creatinine
C2745899|T201|COMP|56654-7|LNC|Nickel/Creatinine|Nickel/Creatinine
C2923066|T201|COMP|58737-8|LNC|Parvovirus B19 Ab.IgG & IgM|Parvovirus B19 Ab.IgG & IgM
C2923067|T201|COMP|58738-6|LNC|Drugs of abuse|Drugs of abuse
C2923068|T201|COMP|58739-4|LNC|Haemophilus influenzae serotype|Haemophilus influenzae serotype
C2923073|T201|COMP|58752-7|LNC|Triticum aestivum recombinant (rTri a) 19 Ab.IgE|Triticum aestivum recombinant (rTri a) 19 Ab.IgE
C2923075|T201|COMP|58753-5|LNC|Corylus avellana recombinant (rCor a) 8 Ab.IgE|Corylus avellana recombinant (rCor a) 8 Ab.IgE
C2923077|T201|COMP|58754-3|LNC|Olea europaea native (nOle e) 1 Ab.IgE|Olea europaea native (nOle e) 1 Ab.IgE
C2923079|T201|COMP|58755-0|LNC|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C2923080|T201|COMP|58756-8|LNC|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C2923081|T201|COMP|58757-6|LNC|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C2923082|T201|COMP|58758-4|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C2923083|T201|COMP|58759-2|LNC|Echovirus Ab|Echovirus Ab
C2923084|T201|COMP|58760-0|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C2923085|T201|COMP|58761-8|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C2923086|T201|COMP|58762-6|LNC|Coxiella burnetii phase 2 Ab.IgG|Coxiella burnetii phase 2 Ab.IgG
C2923087|T201|COMP|58763-4|LNC|IgA|IgA
C2923088|T201|COMP|58764-2|LNC|IgM|IgM
C2923089|T201|COMP|58765-9|LNC|Histone Ab|Histone Ab
C2923090|T201|COMP|58768-3|LNC|Gamma glutamyl transferase|Gamma glutamyl transferase
C2923091|T201|COMP|58769-1|LNC|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C2923093|T201|COMP|58770-9|LNC|Clostridium tetani toxoid Ab.IgG|Clostridium tetani toxoid Ab.IgG
C2923094|T201|COMP|58771-7|LNC|Bactericidal permeability increasing protein Ab|Bactericidal permeability increasing protein Ab
C2923095|T201|COMP|58772-5|LNC|Dog recombinant (rCan f) 2 Ab.IgE|Dog recombinant (rCan f) 2 Ab.IgE
C2923097|T201|COMP|58773-3|LNC|Dog recombinant (rCan f) 1 Ab.IgE|Dog recombinant (rCan f) 1 Ab.IgE
C2923101|T201|COMP|58775-8|LNC|Prunus persica recombinant (rPru p) 4 Ab.IgE|Prunus persica recombinant (rPru p) 4 Ab.IgE
C2923103|T201|COMP|58776-6|LNC|Prunus persica recombinant (rPru p) 1 Ab.IgE|Prunus persica recombinant (rPru p) 1 Ab.IgE
C2923105|T201|COMP|58777-4|LNC|Arachis hypogaea recombinant (rAra h) 3 Ab.IgE|Arachis hypogaea recombinant (rAra h) 3 Ab.IgE
C2923107|T201|COMP|58778-2|LNC|Arachis hypogaea recombinant (rAra h) 2 Ab.IgE|Arachis hypogaea recombinant (rAra h) 2 Ab.IgE
C2923109|T201|COMP|58779-0|LNC|Arachis hypogaea recombinant (rAra h) 1 Ab.IgE|Arachis hypogaea recombinant (rAra h) 1 Ab.IgE
C2923111|T201|COMP|58780-8|LNC|Coxsackievirus B Ab.IgG|Coxsackievirus B Ab.IgG
C2923112|T201|COMP|58781-6|LNC|Calcium|Calcium
C2923113|T201|COMP|58782-4|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C2923114|T201|COMP|58783-2|LNC|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C2923115|T201|COMP|58784-0|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C2923116|T201|COMP|58785-7|LNC|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C2923117|T201|COMP|58786-5|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C2923118|T201|COMP|58787-3|LNC|Corynebacterium diphtheriae Ab.IgG|Corynebacterium diphtheriae Ab.IgG
C2923119|T201|COMP|58788-1|LNC|Campylobacter jejuni Ab.IgM|Campylobacter jejuni Ab.IgM
C2923120|T201|COMP|58789-9|LNC|Campylobacter jejuni Ab.IgG|Campylobacter jejuni Ab.IgG
C2923121|T201|COMP|58790-7|LNC|Coxsackievirus B Ab.IgM|Coxsackievirus B Ab.IgM
C2923122|T201|COMP|58791-5|LNC|Coxsackievirus A9 Ab.IgM|Coxsackievirus A9 Ab.IgM
C2923124|T201|COMP|58792-3|LNC|Coxsackievirus A9 Ab.IgG|Coxsackievirus A9 Ab.IgG
C2923125|T201|COMP|58793-1|LNC|Phytonadione|Phytonadione
C2923126|T201|COMP|58794-9|LNC|5-Hydroxytryptophan|5-Hydroxytryptophan
C2923127|T201|COMP|58795-6|LNC|Glomerular basement membrane Ab.IgG|Glomerular basement membrane Ab.IgG
C2923128|T201|COMP|58796-4|LNC|Glomerular basement membrane Ab.IgG|Glomerular basement membrane Ab.IgG
C2923129|T201|COMP|58797-2|LNC|Yersinia enterocolitica Ab|Yersinia enterocolitica Ab
C2923130|T201|COMP|58798-0|LNC|Legionella pneumophila 2 Ab.IgM|Legionella pneumophila 2 Ab.IgM
C2923131|T201|COMP|58799-8|LNC|Legionella pneumophila 1 Ab.IgG|Legionella pneumophila 1 Ab.IgG
C2923132|T201|COMP|58800-4|LNC|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C2923133|T201|COMP|58801-2|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C2923134|T201|COMP|58802-0|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C2923135|T201|COMP|58803-8|LNC|Acetone/Creatinine|Acetone/Creatinine
C2923137|T201|COMP|58804-6|LNC|Polistes dominulus Ab.IgE|Polistes dominulus Ab.IgE
C2923139|T201|COMP|58805-3|LNC|Leukocytes|Leukocytes
C2923140|T201|COMP|58806-1|LNC|Brucella sp Ab|Brucella sp Ab
C2923141|T201|COMP|58807-9|LNC|Conalbumin native (nGal d) 3 Ab.IgE|Conalbumin native (nGal d) 3 Ab.IgE
C2923143|T201|COMP|58808-7|LNC|Aspergillus sp Ab|Aspergillus sp Ab
C2923144|T201|COMP|58809-5|LNC|Rickettsia conorii Ab.IgG|Rickettsia conorii Ab.IgG
C2923145|T201|COMP|58810-3|LNC|Testosterone^2nd specimen|Testosterone^2nd specimen
C2923146|T201|COMP|58811-1|LNC|Renin^post XXX challenge|Renin^post XXX challenge
C2923147|T201|COMP|58822-8|LNC|Cortisol^22nd specimen|Cortisol^22nd specimen
C2923148|T201|COMP|58823-6|LNC|Cortisol^20th specimen|Cortisol^20th specimen
C2923149|T201|COMP|58824-4|LNC|Cortisol^19th specimen|Cortisol^19th specimen
C2923150|T201|COMP|58825-1|LNC|Cortisol^18th specimen|Cortisol^18th specimen
C2923151|T201|COMP|58826-9|LNC|Cortisol^17th specimen|Cortisol^17th specimen
C2923152|T201|COMP|58827-7|LNC|Cortisol^16th specimen|Cortisol^16th specimen
C2923153|T201|COMP|58828-5|LNC|Cortisol^14th specimen|Cortisol^14th specimen
C2923154|T201|COMP|58829-3|LNC|Cortisol^15th specimen|Cortisol^15th specimen
C2923155|T201|COMP|58830-1|LNC|Cortisol^13th specimen|Cortisol^13th specimen
C2923156|T201|COMP|58831-9|LNC|Urea|Urea
C2923158|T201|COMP|58833-5|LNC|Thyrotropin^20M pre XXX challenge|Thyrotropin^20M pre XXX challenge
C2923159|T201|COMP|58834-3|LNC|Thyrotropin^15M pre XXX challenge|Thyrotropin^15M pre XXX challenge
C2923160|T201|COMP|58835-0|LNC|Testosterone^baseline|Testosterone^baseline
C2923161|T201|COMP|58836-8|LNC|Thyroxine.free^3H post XXX challenge|Thyroxine.free^3H post XXX challenge
C2923162|T201|COMP|58837-6|LNC|Thyroxine.free^2H post XXX challenge|Thyroxine.free^2H post XXX challenge
C2923163|T201|COMP|58838-4|LNC|Thyroxine.free^baseline|Thyroxine.free^baseline
C2923164|T201|COMP|58839-2|LNC|Triiodothyronine.free^3H post XXX challenge|Triiodothyronine.free^3H post XXX challenge
C2923165|T201|COMP|58846-7|LNC|Somatotropin^18th specimen|Somatotropin^18th specimen
C2923166|T201|COMP|58847-5|LNC|Somatotropin^17th specimen|Somatotropin^17th specimen
C2923167|T201|COMP|58848-3|LNC|Somatotropin^16th specimen|Somatotropin^16th specimen
C2923168|T201|COMP|58849-1|LNC|Somatotropin^15th specimen|Somatotropin^15th specimen
C2923169|T201|COMP|58850-9|LNC|Somatotropin^14th specimen|Somatotropin^14th specimen
C2923170|T201|COMP|58851-7|LNC|Testosterone^3D post XXX challenge|Testosterone^3D post XXX challenge
C2923171|T201|COMP|58852-5|LNC|Osmolality^post 1.5H FFst|Osmolality^post 1.5H FFst
C2923172|T201|COMP|58853-3|LNC|Osmolality^post 30M FFst|Osmolality^post 30M FFst
C2923173|T201|COMP|58854-1|LNC|Estradiol^4D post XXX challenge|Estradiol^4D post XXX challenge
C2923174|T201|COMP|58855-8|LNC|Somatotropin^13th specimen|Somatotropin^13th specimen
C2923175|T201|COMP|58856-6|LNC|Somatotropin^10th specimen|Somatotropin^10th specimen
C2923176|T201|COMP|58857-4|LNC|Somatotropin^9th specimen|Somatotropin^9th specimen
C2923177|T201|COMP|58858-2|LNC|Parathyrin.intact^post XXX challenge|Parathyrin.intact^post XXX challenge
C2923178|T201|COMP|58859-0|LNC|Homocyst(e)ine^post XXX challenge|Homocyst(e)ine^post XXX challenge
C2923179|T201|COMP|58860-8|LNC|Somatotropin^48th specimen|Somatotropin^48th specimen
C2923180|T201|COMP|58861-6|LNC|Somatotropin^47th specimen|Somatotropin^47th specimen
C2923181|T201|COMP|58862-4|LNC|Somatotropin^46th specimen|Somatotropin^46th specimen
C2923182|T201|COMP|58863-2|LNC|Somatotropin^45th specimen|Somatotropin^45th specimen
C2923183|T201|COMP|58864-0|LNC|Somatotropin^44th specimen|Somatotropin^44th specimen
C2923184|T201|COMP|58865-7|LNC|Somatotropin^43rd specimen|Somatotropin^43rd specimen
C2923185|T201|COMP|58866-5|LNC|Somatotropin^42nd specimen|Somatotropin^42nd specimen
C2923186|T201|COMP|58867-3|LNC|Somatotropin^41st specimen|Somatotropin^41st specimen
C2923187|T201|COMP|58868-1|LNC|Somatotropin^40th specimen|Somatotropin^40th specimen
C2923188|T201|COMP|58869-9|LNC|Somatotropin^39th specimen|Somatotropin^39th specimen
C2923189|T201|COMP|58870-7|LNC|Somatotropin^38th specimen|Somatotropin^38th specimen
C2923190|T201|COMP|58871-5|LNC|Somatotropin^37th specimen|Somatotropin^37th specimen
C2923191|T201|COMP|58872-3|LNC|Somatotropin^36th specimen|Somatotropin^36th specimen
C2923192|T201|COMP|58873-1|LNC|Somatotropin^35th specimen|Somatotropin^35th specimen
C2923193|T201|COMP|58874-9|LNC|Somatotropin^33rd specimen|Somatotropin^33rd specimen
C2923194|T201|COMP|58882-2|LNC|Somatotropin^23rd specimen|Somatotropin^23rd specimen
C2923195|T201|COMP|58883-0|LNC|Somatotropin^22nd specimen|Somatotropin^22nd specimen
C2923196|T201|COMP|58884-8|LNC|Somatotropin^21st specimen|Somatotropin^21st specimen
C2923197|T201|COMP|58885-5|LNC|Urea|Urea
C2923198|T201|COMP|58886-3|LNC|Pyruvate^30M post XXX challenge|Pyruvate^30M post XXX challenge
C2923199|T201|COMP|58887-1|LNC|Pyruvate^15M post XXX challenge|Pyruvate^15M post XXX challenge
C2923200|T201|COMP|58888-9|LNC|Pyruvate^10M post XXX challenge|Pyruvate^10M post XXX challenge
C2923201|T201|COMP|58889-7|LNC|Pyruvate^3M post XXX challenge|Pyruvate^3M post XXX challenge
C2923202|T201|COMP|58890-5|LNC|Pyruvate^1M post XXX challenge|Pyruvate^1M post XXX challenge
C2923203|T201|COMP|58891-3|LNC|Calcitonin^1M post XXX challenge|Calcitonin^1M post XXX challenge
C2923204|T201|COMP|58892-1|LNC|Calcitonin^baseline|Calcitonin^baseline
C2923205|T201|COMP|58893-9|LNC|Vasopressin^1.5H post XXX challenge|Vasopressin^1.5H post XXX challenge
C2923206|T201|COMP|58894-7|LNC|Vasopressin^baseline|Vasopressin^baseline
C2923207|T201|COMP|58895-4|LNC|Pyruvate^post exercise|Pyruvate^post exercise
C2923208|T201|COMP|58896-2|LNC|C peptide^post XXX challenge|C peptide^post XXX challenge
C2923209|T201|COMP|58897-0|LNC|Methyl ethyl ketone/Creatinine|Methyl ethyl ketone/Creatinine
C2923211|T201|COMP|58898-8|LNC|Renin^4H post XXX challenge|Renin^4H post XXX challenge
C2923212|T201|COMP|58899-6|LNC|Aldosterone^4H post XXX challenge|Aldosterone^4H post XXX challenge
C2923213|T201|COMP|58900-2|LNC|HIV 1+2 Ab+HIV1 p24 Ag|HIV 1+2 Ab+HIV1 p24 Ag
C2923214|T201|COMP|58901-0|LNC|Spermatozoa.progressive|Spermatozoa.progressive
C2923215|T201|COMP|58902-8|LNC|F12 gene mutations tested for|F12 gene mutations tested for
C2923217|T201|COMP|58903-6|LNC|Neomycin Ab.IgE|Neomycin Ab.IgE
C2923219|T201|COMP|58907-7|LNC|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C2923220|T201|COMP|58908-5|LNC|11-Deoxycortisol^40M post XXX challenge|11-Deoxycortisol^40M post XXX challenge
C2923221|T201|COMP|58909-3|LNC|11-Deoxycortisol^20M post XXX challenge|11-Deoxycortisol^20M post XXX challenge
C2923222|T201|COMP|58910-1|LNC|11-Deoxycortisol^2.5H post XXX challenge|11-Deoxycortisol^2.5H post XXX challenge
C2923223|T201|COMP|58911-9|LNC|Chicken droppings Ab.IgG|Chicken droppings Ab.IgG
C2923225|T201|COMP|58912-7|LNC|Pigeon feather Ab.IgG|Pigeon feather Ab.IgG
C2923226|T201|COMP|58913-5|LNC|Parrot feather Ab.IgG|Parrot feather Ab.IgG
C2923227|T201|COMP|58914-3|LNC|Aspergillus niger Ab.IgG|Aspergillus niger Ab.IgG
C2923228|T201|COMP|58915-0|LNC|Parakeet feather Ab.IgG|Parakeet feather Ab.IgG
C2923230|T201|COMP|58916-8|LNC|Canary feather Ab.IgG|Canary feather Ab.IgG
C2923231|T201|COMP|58917-6|LNC|Androstanolone^1H post XXX challenge|Androstanolone^1H post XXX challenge
C2923232|T201|COMP|58918-4|LNC|Androstanolone^30M post XXX challenge|Androstanolone^30M post XXX challenge
C2923233|T201|COMP|58919-2|LNC|Androstenedione^1.5H post XXX challenge|Androstenedione^1.5H post XXX challenge
C2923234|T201|COMP|58920-0|LNC|Cells.CD4+CD45RO+/Cells.CD3+CD4+|Cells.CD4+CD45RO+/Cells.CD3+CD4+
C2923236|T201|COMP|58921-8|LNC|Glutamine+Histidine|Glutamine+Histidine
C2923238|T201|COMP|58922-6|LNC|Vasopressin^2H post XXX challenge|Vasopressin^2H post XXX challenge
C2923239|T201|COMP|58923-4|LNC|Lolium perenne Ab.IgG|Lolium perenne Ab.IgG
C2923240|T201|COMP|58924-2|LNC|LCT gene mutations tested for|LCT gene mutations tested for
C2923242|T201|COMP|58925-9|LNC|Dextromethamphetamine|Dextromethamphetamine
C2923243|T201|COMP|58927-5|LNC|Glutamine+Histidine/Creatinine|Glutamine+Histidine/Creatinine
C2923245|T201|COMP|58928-3|LNC|HLA-DQA1*03:01|HLA-DQA1*03:01
C2923247|T201|COMP|58929-1|LNC|HLA-DQB1*03:02|HLA-DQB1*03:02
C2923249|T201|COMP|58930-9|LNC|Glutamine+Histidine|Glutamine+Histidine
C2923250|T201|COMP|58931-7|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C2923251|T201|COMP|58932-5|LNC|Protoporphyrin|Protoporphyrin
C2923252|T201|COMP|58933-3|LNC|Endothelial cell Ab|Endothelial cell Ab
C2923254|T201|COMP|58935-8|LNC|Yersinia pseudotuberculosis Ab|Yersinia pseudotuberculosis Ab
C2923255|T201|COMP|58936-6|LNC|Hepatitis E virus Ab|Hepatitis E virus Ab
C2923256|T201|COMP|58937-4|LNC|F12 gene targeted mutation analysis|F12 gene targeted mutation analysis
C2923258|T201|COMP|58938-2|LNC|LCT gene targeted mutation analysis|LCT gene targeted mutation analysis
C2923260|T201|COMP|58939-0|LNC|Cells.CD34|Cells.CD34
C2923261|T201|COMP|58940-8|LNC|Bacteria identified|Bacteria identified
C2923262|T201|COMP|58941-6|LNC|Bilirubin|Bilirubin
C2923267|T201|COMP|58946-5|LNC|Lutropin^pre XXX challenge|Lutropin^pre XXX challenge
C2923268|T201|COMP|58947-3|LNC|Follitropin^pre XXX challenge|Follitropin^pre XXX challenge
C2923269|T201|COMP|58958-0|LNC|Fusarium oxysporum Ab.IgG|Fusarium oxysporum Ab.IgG
C2923273|T201|COMP|58961-4|LNC|Ganglioside GT1b Ab.IgM|Ganglioside GT1b Ab.IgM
C2923275|T201|COMP|58962-2|LNC|Ganglioside GT1b Ab.IgG|Ganglioside GT1b Ab.IgG
C2923277|T201|COMP|58963-0|LNC|Ganglioside GT1a Ab.IgM|Ganglioside GT1a Ab.IgM
C2923279|T201|COMP|58964-8|LNC|Ganglioside GT1a Ab.IgG|Ganglioside GT1a Ab.IgG
C2923281|T201|COMP|58965-5|LNC|Ganglioside GM4 Ab.IgM|Ganglioside GM4 Ab.IgM
C2923283|T201|COMP|58966-3|LNC|Ganglioside GM4 Ab.IgG|Ganglioside GM4 Ab.IgG
C2923285|T201|COMP|58967-1|LNC|Ganglioside GM3 Ab.IgM|Ganglioside GM3 Ab.IgM
C2923287|T201|COMP|58968-9|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C2923288|T201|COMP|58969-7|LNC|Ganglioside GD1a Ab.IgG|Ganglioside GD1a Ab.IgG
C2923289|T201|COMP|58970-5|LNC|Ganglioside GD1a Ab.IgM|Ganglioside GD1a Ab.IgM
C2923290|T201|COMP|58971-3|LNC|Ganglioside GD1b Ab.IgG|Ganglioside GD1b Ab.IgG
C2923291|T201|COMP|58972-1|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C2923292|T201|COMP|58973-9|LNC|Ganglioside GM2 Ab.IgG|Ganglioside GM2 Ab.IgG
C2923293|T201|COMP|58974-7|LNC|Ganglioside GM2 Ab.IgM|Ganglioside GM2 Ab.IgM
C2923294|T201|COMP|58975-4|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C2923295|T201|COMP|58976-2|LNC|Ganglioside GQ1b Ab.IgM|Ganglioside GQ1b Ab.IgM
C2923296|T201|COMP|58977-0|LNC|Ganglioside GD1b Ab.IgM|Ganglioside GD1b Ab.IgM
C2923297|T201|COMP|58978-8|LNC|Ganglioside GD3 Ab.IgM|Ganglioside GD3 Ab.IgM
C2923299|T201|COMP|58979-6|LNC|Ganglioside GD3 Ab.IgG|Ganglioside GD3 Ab.IgG
C2923301|T201|COMP|58980-4|LNC|Ganglioside GD2 Ab.IgM|Ganglioside GD2 Ab.IgM
C2923303|T201|COMP|58981-2|LNC|Phleum pratense recombinant (rPhl p) 5b Ab.IgE|Phleum pratense recombinant (rPhl p) 5b Ab.IgE
C2923305|T201|COMP|58982-0|LNC|Quercus ilex Ab.IgE|Quercus ilex Ab.IgE
C2923309|T201|COMP|58984-6|LNC|Bromelin MUXF3 Ab.IgE|Bromelin MUXF3 Ab.IgE
C2923311|T201|COMP|58985-3|LNC|11-Deoxycortisol^pre XXX challenge|11-Deoxycortisol^pre XXX challenge
C2923314|T201|COMP|58987-9|LNC|ITGB3 gene targeted mutation analysis|ITGB3 gene targeted mutation analysis
C2923316|T201|COMP|58988-7|LNC|FGB gene targeted mutation analysis|FGB gene targeted mutation analysis
C2923318|T201|COMP|58989-5|LNC|Specimen volume|Specimen volume
C2923319|T201|COMP|58990-3|LNC|Urate|Urate
C2923320|T201|COMP|58991-1|LNC|Urea|Urea
C2923321|T201|COMP|58992-9|LNC|Protein|Protein
C2923322|T201|COMP|58993-7|LNC|Phosphate|Phosphate
C2923323|T201|COMP|58994-5|LNC|Sodium|Sodium
C2923324|T201|COMP|58995-2|LNC|Magnesium|Magnesium
C2923325|T201|COMP|58996-0|LNC|Potassium|Potassium
C2923326|T201|COMP|58997-8|LNC|Glucose|Glucose
C2923327|T201|COMP|58998-6|LNC|Creatinine|Creatinine
C2923328|T201|COMP|58999-4|LNC|Chloride|Chloride
C2923329|T201|COMP|59000-0|LNC|Calcium|Calcium
C2923330|T201|COMP|59001-8|LNC|Amylase|Amylase
C2923331|T201|COMP|59002-6|LNC|Paliperidone|Paliperidone
C2923332|T201|COMP|59003-4|LNC|Lactoferrin Ab|Lactoferrin Ab
C2923333|T201|COMP|59004-2|LNC|Lactate^baseline|Lactate^baseline
C2923334|T201|COMP|59005-9|LNC|Lactate^1M post XXX challenge|Lactate^1M post XXX challenge
C2923335|T201|COMP|59006-7|LNC|Lactate^3M post XXX challenge|Lactate^3M post XXX challenge
C2923336|T201|COMP|59007-5|LNC|Lactate^5M post XXX challenge|Lactate^5M post XXX challenge
C2923338|T201|COMP|59009-1|LNC|Fractional excretion of urea|Fractional excretion of urea
C2923340|T201|COMP|59010-9|LNC|Fractional excretion of potassium|Fractional excretion of potassium
C2923341|T201|COMP|59011-7|LNC|Lactate^10M post XXX challenge|Lactate^10M post XXX challenge
C2923342|T201|COMP|59012-5|LNC|Lactate^15M post XXX challenge|Lactate^15M post XXX challenge
C2923343|T201|COMP|59013-3|LNC|Lactate^30M post XXX challenge|Lactate^30M post XXX challenge
C2923344|T201|COMP|59014-1|LNC|Sjogrens syndrome-A extractable nuclear 60kD Ab|Sjogrens syndrome-A extractable nuclear 60kD Ab
C2923345|T201|COMP|59044-8|LNC|ACE gene mutations tested for|ACE gene mutations tested for
C2923347|T201|COMP|59045-5|LNC|ITGB3 gene mutations tested for|ITGB3 gene mutations tested for
C2923349|T201|COMP|59046-3|LNC|FGB gene mutations tested for|FGB gene mutations tested for
C2923351|T201|COMP|59047-1|LNC|F5 gene.p.His1299Arg|F5 gene.p.His1299Arg
C2923353|T201|COMP|59048-9|LNC|Lactate/Pyruvate|Lactate/Pyruvate
C2923354|T201|COMP|59049-7|LNC|Coccidioides sp Ab.IgG & IgM panel|Coccidioides sp Ab.IgG & IgM panel
C2923356|T201|COMP|59050-5|LNC|Chromosome analysis.interphase|Chromosome analysis.interphase
C2923357|T201|COMP|59051-3|LNC|Bacteria identified^^^4|Bacteria identified^^^4
C2923358|T201|COMP|59052-1|LNC|HIV 1+Hepatitis C virus RNA+Hepatitis B virus DNA|HIV 1+Hepatitis C virus RNA+Hepatitis B virus DNA
C2923360|T201|COMP|59053-9|LNC|Glucagon^5th specimen post CFst|Glucagon^5th specimen post CFst
C2923361|T201|COMP|59054-7|LNC|Glucagon^4th specimen post CFst|Glucagon^4th specimen post CFst
C2923362|T201|COMP|59055-4|LNC|Glucagon^3rd specimen post CFst|Glucagon^3rd specimen post CFst
C2923363|T201|COMP|59056-2|LNC|Glucagon^2nd specimen post CFst|Glucagon^2nd specimen post CFst
C2923364|T201|COMP|59057-0|LNC|Glucagon^1st specimen post CFst|Glucagon^1st specimen post CFst
C2923365|T201|COMP|59058-8|LNC|Cow whey Ab.IgG|Cow whey Ab.IgG
C2923367|T201|COMP|59059-6|LNC|Inflammatory bowel disease Ab 7 panel|Inflammatory bowel disease Ab 7 panel
C2923369|T201|COMP|59060-4|LNC|Inflammatory bowel disease Ab 7|Inflammatory bowel disease Ab 7
C2923371|T201|COMP|59061-2|LNC|Adulterants|Adulterants
C2923373|T201|COMP|59062-0|LNC|Lipoprofile panel|Lipoprofile panel
C2923375|T201|COMP|59063-8|LNC|Lymphocyte proliferation panel|Lymphocyte proliferation panel
C2923377|T201|COMP|59064-6|LNC|PAX6 gene targeted mutation analysis|PAX6 gene targeted mutation analysis
C2923379|T201|COMP|59065-3|LNC|Chlamydophila psittaci|Chlamydophila psittaci
C2923380|T201|COMP|59066-1|LNC|sp100 Ab|sp100 Ab
C2923381|T201|COMP|59067-9|LNC|ALAS2 gene targeted mutation analysis|ALAS2 gene targeted mutation analysis
C2923383|T201|COMP|59068-7|LNC|RPS19 gene targeted mutation analysis|RPS19 gene targeted mutation analysis
C2923385|T201|COMP|59069-5|LNC|Nuclear Ab|Nuclear Ab
C2923386|T201|COMP|59070-3|LNC|Paraquat|Paraquat
C2923387|T201|COMP|59071-1|LNC|Tropheryma whippelii Ab|Tropheryma whippelii Ab
C2923389|T201|COMP|59072-9|LNC|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C2923494|T201|COMP|59134-7|LNC|ePHEDrine|ePHEDrine
C2923495|T201|COMP|59135-4|LNC|Benzylpiperazine|Benzylpiperazine
C2923497|T201|COMP|59136-2|LNC|Cells.CD11c+CD103+/100 cells|Cells.CD11c+CD103+/100 cells
C2923499|T201|COMP|59137-0|LNC|Cells.CD5+CD23+/100 cells|Cells.CD5+CD23+/100 cells
C2923500|T201|COMP|59138-8|LNC|Cells.CD7+CD34+/100 cells|Cells.CD7+CD34+/100 cells
C2923502|T201|COMP|59139-6|LNC|Cells.CD19+CD34+/100 cells|Cells.CD19+CD34+/100 cells
C2923503|T201|COMP|59140-4|LNC|Cells.CD13+CD34+/100 cells|Cells.CD13+CD34+/100 cells
C2923505|T201|COMP|59141-2|LNC|Cells.CD11c-CD103+/100 cells|Cells.CD11c-CD103+/100 cells
C2923507|T201|COMP|59150-3|LNC|Enterococcus species.vancomycin resistant|Enterococcus species.vancomycin resistant
C2923508|T201|COMP|59151-1|LNC|Enterococcus species.vancomycin resistant|Enterococcus species.vancomycin resistant
C2923509|T201|COMP|59152-9|LNC|Enterococcus species.vancomycin resistant DNA|Enterococcus species.vancomycin resistant DNA
C2923511|T201|COMP|59164-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C2923512|T201|COMP|59165-1|LNC|Carbon dioxide|Carbon dioxide
C2923513|T201|COMP|59166-9|LNC|Bilirubin|Bilirubin
C2923514|T201|COMP|59167-7|LNC|Phosphate|Phosphate
C2923515|T201|COMP|59168-5|LNC|Urea|Urea
C2923516|T201|COMP|59169-3|LNC|buPROPion|buPROPion
C2923517|T201|COMP|59170-1|LNC|Citalopram|Citalopram
C2923518|T201|COMP|59171-9|LNC|Norclozapine|Norclozapine
C2923519|T201|COMP|59172-7|LNC|Methotrimeprazine metabolite|Methotrimeprazine metabolite
C2923521|T201|COMP|59323-6|LNC|Rufinamide|Rufinamide
C2923522|T201|COMP|59324-4|LNC|Salvinorin A|Salvinorin A
C2923523|T201|COMP|59290-7|LNC|Iloperidone|Iloperidone
C2923524|T201|COMP|59291-5|LNC|Levamisole|Levamisole
C2923525|T201|COMP|59292-3|LNC|Levamisole|Levamisole
C2923526|T201|COMP|59293-1|LNC|Levamisole|Levamisole
C2923527|T201|COMP|59294-9|LNC|Levamisole|Levamisole
C2923528|T201|COMP|59295-6|LNC|Levamisole|Levamisole
C2923529|T201|COMP|59296-4|LNC|Lacosamide|Lacosamide
C2923530|T201|COMP|59297-2|LNC|Lacosamide|Lacosamide
C2923531|T201|COMP|59298-0|LNC|Lacosamide|Lacosamide
C2923532|T201|COMP|59299-8|LNC|Desloratadine|Desloratadine
C2923533|T201|COMP|59571-0|LNC|Triglyceride|Triglyceride
C2923534|T201|COMP|59572-8|LNC|Triglyceride|Triglyceride
C2923535|T201|COMP|59573-6|LNC|Cannabinoids|Cannabinoids
C2923539|T201|COMP|59577-7|LNC|Glucagon^7th specimen post CFst|Glucagon^7th specimen post CFst
C2923540|T201|COMP|59578-5|LNC|Glucagon^6th specimen post CFst|Glucagon^6th specimen post CFst
C2923541|T201|COMP|59579-3|LNC|Coxsackievirus A24 Ab.IgM|Coxsackievirus A24 Ab.IgM
C2923543|T201|COMP|59580-1|LNC|Coxsackievirus A16 Ab.IgM|Coxsackievirus A16 Ab.IgM
C2923545|T201|COMP|59325-1|LNC|Salvinorin B|Salvinorin B
C2923546|T201|COMP|59326-9|LNC|Salvinorin A|Salvinorin A
C2923547|T201|COMP|59327-7|LNC|Salvinorin B|Salvinorin B
C2923548|T201|COMP|59328-5|LNC|Salvinorin A|Salvinorin A
C2923549|T201|COMP|59329-3|LNC|Salvinorin B|Salvinorin B
C2923550|T201|COMP|59330-1|LNC|Norsibutramine|Norsibutramine
C2923552|T201|COMP|59801-1|LNC|Protein.monoclonal band 3/Protein.total|Protein.monoclonal band 3/Protein.total
C2923553|T201|COMP|59802-9|LNC|Protein.monoclonal band 4/Protein.total|Protein.monoclonal band 4/Protein.total
C2923554|T201|COMP|59803-7|LNC|Cortisol^30M post XXX challenge|Cortisol^30M post XXX challenge
C2923555|T201|COMP|59804-5|LNC|Cortisol^1H post XXX challenge|Cortisol^1H post XXX challenge
C2923556|T201|COMP|59805-2|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C2923558|T201|COMP|59807-8|LNC|Phosphatidylglycerol|Phosphatidylglycerol
C2923559|T201|COMP|59808-6|LNC|Lymphocytes.large granular|Lymphocytes.large granular
C2923560|T201|COMP|59809-4|LNC|Lymphoma cells|Lymphoma cells
C2923561|T201|COMP|59812-8|LNC|Glucose^11 AM specimen|Glucose^11 AM specimen
C2923562|T201|COMP|59813-6|LNC|Glucose^7 AM specimen|Glucose^7 AM specimen
C2923563|T201|COMP|59814-4|LNC|Glucose^7 AM specimen|Glucose^7 AM specimen
C2923564|T201|COMP|59174-3|LNC|QUEtiapine|QUEtiapine
C2923565|T201|COMP|59175-0|LNC|QUEtiapine metabolite|QUEtiapine metabolite
C2923567|T201|COMP|59176-8|LNC|Zopiclone|Zopiclone
C2923568|T201|COMP|59178-4|LNC|Chloride|Chloride
C2923569|T201|COMP|59179-2|LNC|Insulin^post CFst|Insulin^post CFst
C2923570|T201|COMP|59180-0|LNC|Monoethylglycinexylidide|Monoethylglycinexylidide
C2923571|T201|COMP|59181-8|LNC|Interferon.beta given|Interferon.beta given
C2923573|T201|COMP|59182-6|LNC|C reactive protein|C reactive protein
C2923574|T201|COMP|59183-4|LNC|Epstein Barr virus early diffuse Ab.IgG|Epstein Barr virus early diffuse Ab.IgG
C2923575|T201|COMP|59185-9|LNC|Hemoglobin H inclusion bodies|Hemoglobin H inclusion bodies
C2923577|T201|COMP|59186-7|LNC|Cyanide|Cyanide
C2923578|T201|COMP|59187-5|LNC|Urea renal clearance/1.73 sq M|Urea renal clearance/1.73 sq M
C2923579|T201|COMP|59188-3|LNC|Alkaline phosphatase.placental|Alkaline phosphatase.placental
C2923580|T201|COMP|59189-1|LNC|Methyl ethyl ketone/Creatinine|Methyl ethyl ketone/Creatinine
C2923581|T201|COMP|59190-9|LNC|2-Hydroxycaproate/Creatinine|2-Hydroxycaproate/Creatinine
C2923583|T201|COMP|59191-7|LNC|2-Ketobutyrate/Creatinine|2-Ketobutyrate/Creatinine
C2923585|T201|COMP|59192-5|LNC|3-Methyl crotonate/Creatinine|3-Methyl crotonate/Creatinine
C2923587|T201|COMP|59193-3|LNC|Deoxyuridine/Creatinine|Deoxyuridine/Creatinine
C2923590|T201|COMP|59195-8|LNC|3-Hydroxydodecenoylcarnitine (C12:1-OH)|3-Hydroxydodecenoylcarnitine (C12:1-OH)
C2923592|T201|COMP|59197-4|LNC|Propionylcarnitine (C3)/Palmitoylcarnitine (C16)|Propionylcarnitine (C3)/Palmitoylcarnitine (C16)
C2923593|T201|COMP|59198-2|LNC|Propionylcarnitine (C3)/Acetylcarnitine (C2)|Propionylcarnitine (C3)/Acetylcarnitine (C2)
C2923594|T201|COMP|59199-0|LNC|Deoxyadenosine/Creatinine|Deoxyadenosine/Creatinine
C2923596|T201|COMP|59200-6|LNC|Octanoylcarnitine (C8)/Acetylcarnitine (C2)|Octanoylcarnitine (C8)/Acetylcarnitine (C2)
C2923597|T201|COMP|59201-4|LNC|Deoxyguanosine/Creatinine|Deoxyguanosine/Creatinine
C2923599|T201|COMP|59202-2|LNC|Deoxyinosine/Creatinine|Deoxyinosine/Creatinine
C2923601|T201|COMP|59203-0|LNC|Adenine/Creatinine|Adenine/Creatinine
C2923603|T201|COMP|59205-5|LNC|Gamma tocopherol|Gamma tocopherol
C2923605|T201|COMP|59207-1|LNC|Dicarboxyoleylcarnitine (C18:1-DC)|Dicarboxyoleylcarnitine (C18:1-DC)
C2923606|T201|COMP|59208-9|LNC|Octanoylcarnitine (C8)/Decanoylcarnitine (C10)|Octanoylcarnitine (C8)/Decanoylcarnitine (C10)
C2923607|T201|COMP|59209-7|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C2923608|T201|COMP|59210-5|LNC|Inosine/Creatinine|Inosine/Creatinine
C2923610|T201|COMP|59211-3|LNC|Transcobalamin I+Transcobalamin III|Transcobalamin I+Transcobalamin III
C2923612|T201|COMP|59212-1|LNC|Alloisoleucine|Alloisoleucine
C2923613|T201|COMP|59213-9|LNC|Alloisoleucine|Alloisoleucine
C2923614|T201|COMP|59214-7|LNC|Succinyladenosine/Creatinine|Succinyladenosine/Creatinine
C2923616|T201|COMP|59215-4|LNC|Thymidine/Creatinine|Thymidine/Creatinine
C2923618|T201|COMP|59216-2|LNC|Uridine/Creatinine|Uridine/Creatinine
C2923620|T201|COMP|59217-0|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C2923621|T201|COMP|59218-8|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C2923622|T201|COMP|59219-6|LNC|Testosterone|Testosterone
C2923623|T201|COMP|59220-4|LNC|Chromogranin A|Chromogranin A
C2923624|T201|COMP|59221-2|LNC|Prostate specific Ag|Prostate specific Ag
C2923625|T201|COMP|59222-0|LNC|Squamous cell carcinoma Ag|Squamous cell carcinoma Ag
C2923626|T201|COMP|59223-8|LNC|Prostate specific Ag|Prostate specific Ag
C2923627|T201|COMP|59224-6|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C2923628|T201|COMP|59225-3|LNC|Squamous cell carcinoma Ag|Squamous cell carcinoma Ag
C2923629|T201|COMP|59226-1|LNC|Chromogranin A|Chromogranin A
C2923630|T201|COMP|59227-9|LNC|Chromogranin A|Chromogranin A
C2923631|T201|COMP|59228-7|LNC|Squamous cell carcinoma Ag|Squamous cell carcinoma Ag
C2923632|T201|COMP|59229-5|LNC|Testosterone|Testosterone
C2923633|T201|COMP|59230-3|LNC|Prostate specific Ag|Prostate specific Ag
C2923634|T201|COMP|59231-1|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C2923635|T201|COMP|59232-9|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C2923636|T201|COMP|59233-7|LNC|Testosterone|Testosterone
C2923637|T201|COMP|59234-5|LNC|Reducing substances|Reducing substances
C2923642|T201|COMP|59239-4|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C2923643|T201|COMP|59240-2|LNC|Testosterone|Testosterone
C2923644|T201|COMP|59241-0|LNC|Chromogranin A|Chromogranin A
C2923645|T201|COMP|59242-8|LNC|Reducing substances|Reducing substances
C2923646|T201|COMP|59244-4|LNC|Arylsulfatase C|Arylsulfatase C
C2923647|T201|COMP|59245-1|LNC|Alanine glyoxylate aminotransferase|Alanine glyoxylate aminotransferase
C2923648|T201|COMP|59247-7|LNC|Tetrahydrobiopterin|Tetrahydrobiopterin
C2923649|T201|COMP|59248-5|LNC|Cholesterol esterase|Cholesterol esterase
C2923650|T201|COMP|59249-3|LNC|Acylcarnitine/Acylcarnitine+Carnitine Free (C0)|Acylcarnitine/Acylcarnitine+Carnitine Free (C0)
C2923652|T201|COMP|59250-1|LNC|Tocopherols/Cholesterol|Tocopherols/Cholesterol
C2923654|T201|COMP|59251-9|LNC|N-carbamoyl beta alanine/Creatinine|N-carbamoyl beta alanine/Creatinine
C2923656|T201|COMP|59252-7|LNC|Homocysteine cysteine disulfide|Homocysteine cysteine disulfide
C2923657|T201|COMP|59253-5|LNC|Homocysteine cysteine disulfide|Homocysteine cysteine disulfide
C2923658|T201|COMP|59254-3|LNC|Acylcarnitine/Acylcarnitine+Carnitine Free (C0)|Acylcarnitine/Acylcarnitine+Carnitine Free (C0)
C2923660|T201|COMP|59256-8|LNC|Cytologist|Cytologist
C2923661|T201|COMP|59257-6|LNC|Cell count & Differential panel|Cell count & Differential panel
C2923664|T201|COMP|59260-0|LNC|Hemoglobin|Hemoglobin
C2923665|T201|COMP|59261-8|LNC|Hemoglobin A1c/Hemoglobin.total|Hemoglobin A1c/Hemoglobin.total
C2923666|T201|COMP|59262-6|LNC|Leukocyte esterase|Leukocyte esterase
C2923667|T201|COMP|59263-4|LNC|Human papilloma virus 16 DNA|Human papilloma virus 16 DNA
C2923669|T201|COMP|59264-2|LNC|Human papilloma virus 18 DNA|Human papilloma virus 18 DNA
C2923671|T201|COMP|59274-1|LNC|Oxygen content|Oxygen content
C2923672|T201|COMP|59275-8|LNC|Oxygen capacity|Oxygen capacity
C2923674|T201|COMP|59276-6|LNC|Calcium hydrogen phosphate dihydrate crystals|Calcium hydrogen phosphate dihydrate crystals
C2923675|T201|COMP|59277-4|LNC|Cystine crystals|Cystine crystals
C2923676|T201|COMP|59278-2|LNC|Calcium oxalate dihydrate crystals|Calcium oxalate dihydrate crystals
C2923677|T201|COMP|59279-0|LNC|Urate crystals|Urate crystals
C2923678|T201|COMP|59280-8|LNC|Urate dihydrate crystals|Urate dihydrate crystals
C2923686|T201|COMP|59285-7|LNC|Benzylpiperazine|Benzylpiperazine
C2923687|T201|COMP|59286-5|LNC|Benzylpiperazine|Benzylpiperazine
C2923688|T201|COMP|59287-3|LNC|Benzylpiperazine|Benzylpiperazine
C2923689|T201|COMP|59288-1|LNC|Bisphenol A|Bisphenol A
C2923690|T201|COMP|59289-9|LNC|Iloperidone|Iloperidone
C2923691|T201|COMP|59300-4|LNC|Desloratadine|Desloratadine
C2923692|T201|COMP|59301-2|LNC|Desloratadine|Desloratadine
C2923693|T201|COMP|59302-0|LNC|Memantine|Memantine
C2923694|T201|COMP|59303-8|LNC|Memantine|Memantine
C2923695|T201|COMP|59304-6|LNC|Memantine|Memantine
C2923696|T201|COMP|59305-3|LNC|Memantine|Memantine
C2923697|T201|COMP|59306-1|LNC|Memantine|Memantine
C2923698|T201|COMP|59307-9|LNC|Metaxalone|Metaxalone
C2923699|T201|COMP|59308-7|LNC|Metaxalone|Metaxalone
C2923700|T201|COMP|59309-5|LNC|Metaxalone|Metaxalone
C2923701|T201|COMP|59310-3|LNC|Milnacipran|Milnacipran
C2923702|T201|COMP|59311-1|LNC|Milnacipran|Milnacipran
C2923703|T201|COMP|59312-9|LNC|Milnacipran|Milnacipran
C2923704|T201|COMP|59313-7|LNC|Ramelteon M-II|Ramelteon M-II
C2923706|T201|COMP|59314-5|LNC|Ramelteon|Ramelteon
C2923707|T201|COMP|59315-2|LNC|Ramelteon M-II|Ramelteon M-II
C2923708|T201|COMP|59316-0|LNC|Ramelteon|Ramelteon
C2923709|T201|COMP|59317-8|LNC|Ramelteon M-II|Ramelteon M-II
C2923710|T201|COMP|59318-6|LNC|Ramelteon|Ramelteon
C2923711|T201|COMP|59319-4|LNC|Ramelteon M-II|Ramelteon M-II
C2923712|T201|COMP|59320-2|LNC|Ramelteon|Ramelteon
C2923713|T201|COMP|59321-0|LNC|Ramelteon M-II|Ramelteon M-II
C2923714|T201|COMP|59322-8|LNC|Ramelteon|Ramelteon
C2923715|T201|COMP|59331-9|LNC|Dinorsibutramine|Dinorsibutramine
C2923717|T201|COMP|59332-7|LNC|Sibutramine|Sibutramine
C2923718|T201|COMP|59333-5|LNC|Norsibutramine|Norsibutramine
C2923719|T201|COMP|59334-3|LNC|Dinorsibutramine|Dinorsibutramine
C2923720|T201|COMP|59335-0|LNC|Sibutramine|Sibutramine
C2923721|T201|COMP|59336-8|LNC|Norsibutramine|Norsibutramine
C2923722|T201|COMP|59337-6|LNC|Dinorsibutramine|Dinorsibutramine
C2923723|T201|COMP|59338-4|LNC|Sibutramine|Sibutramine
C2923724|T201|COMP|59339-2|LNC|Stiripentol|Stiripentol
C2923725|T201|COMP|59340-0|LNC|Stiripentol|Stiripentol
C2923726|T201|COMP|59341-8|LNC|Stiripentol|Stiripentol
C2923727|T201|COMP|59342-6|LNC|Tadalafil|Tadalafil
C2923728|T201|COMP|59343-4|LNC|Tadalafil|Tadalafil
C2923729|T201|COMP|59344-2|LNC|Tadalafil|Tadalafil
C2923730|T201|COMP|59345-9|LNC|Endoxifen|Endoxifen
C2923731|T201|COMP|59346-7|LNC|4-Hydroxy-Tamoxifen|4-Hydroxy-Tamoxifen
C2923732|T201|COMP|59347-5|LNC|Tamoxifen|Tamoxifen
C2923733|T201|COMP|59348-3|LNC|Nortamoxifen|Nortamoxifen
C2923735|T201|COMP|59349-1|LNC|Endoxifen|Endoxifen
C2923736|T201|COMP|59350-9|LNC|4-Hydroxy-Tamoxifen|4-Hydroxy-Tamoxifen
C2923737|T201|COMP|59351-7|LNC|Nortamoxifen|Nortamoxifen
C2923738|T201|COMP|59352-5|LNC|Tapentadol|Tapentadol
C2923739|T201|COMP|59353-3|LNC|Tapentadol|Tapentadol
C2923740|T201|COMP|59354-1|LNC|Tapentadol|Tapentadol
C2923741|T201|COMP|59355-8|LNC|Tapentadol|Tapentadol
C2923742|T201|COMP|59356-6|LNC|Desethylvardenafil|Desethylvardenafil
C2923744|T201|COMP|59357-4|LNC|Vardenafil|Vardenafil
C2923745|T201|COMP|59358-2|LNC|Desethylvardenafil|Desethylvardenafil
C2923746|T201|COMP|59709-6|LNC|Midazolam|Midazolam
C2923747|T201|COMP|59710-4|LNC|Midazolam|Midazolam
C2923748|T201|COMP|59711-2|LNC|Midazolam|Midazolam
C2923749|T201|COMP|59712-0|LNC|Midazolam|Midazolam
C2923750|T201|COMP|59713-8|LNC|Midazolam|Midazolam
C2923751|T201|COMP|59714-6|LNC|Nitrous oxide|Nitrous oxide
C2923752|T201|COMP|59715-3|LNC|Nitrous oxide|Nitrous oxide
C2923753|T201|COMP|59716-1|LNC|Nordiazepam|Nordiazepam
C2923754|T201|COMP|59717-9|LNC|Nordiazepam|Nordiazepam
C2923755|T201|COMP|59718-7|LNC|Nordiazepam|Nordiazepam
C2923756|T201|COMP|59719-5|LNC|Nordiazepam|Nordiazepam
C2923757|T201|COMP|59720-3|LNC|Nordiazepam|Nordiazepam
C2923758|T201|COMP|59721-1|LNC|Nordiazepam|Nordiazepam
C2923759|T201|COMP|59722-9|LNC|Nordiazepam|Nordiazepam
C2923760|T201|COMP|59359-0|LNC|Vardenafil|Vardenafil
C2923761|T201|COMP|59360-8|LNC|Desethylvardenafil|Desethylvardenafil
C2923762|T201|COMP|59361-6|LNC|Vardenafil|Vardenafil
C2923764|T201|COMP|59363-2|LNC|Leptospira interrogans serovar Manhao Ab|Leptospira interrogans serovar Manhao Ab
C2923766|T201|COMP|59364-0|LNC|Leptospira interrogans serovar Pyrogenes Ab|Leptospira interrogans serovar Pyrogenes Ab
C2923768|T201|COMP|59365-7|LNC|Leptospira interrogans serovar Mini Ab|Leptospira interrogans serovar Mini Ab
C2923770|T201|COMP|59366-5|LNC|Leptospira interrogans serovar Sejroe Ab|Leptospira interrogans serovar Sejroe Ab
C2923772|T201|COMP|59367-3|LNC|Leptospira interrogans serovar Tarassovi Ab|Leptospira interrogans serovar Tarassovi Ab
C2923774|T201|COMP|59368-1|LNC|Leptospira interrogans serovar Bataviae Ab|Leptospira interrogans serovar Bataviae Ab
C2923775|T201|COMP|59369-9|LNC|Leptospira interrogans serovar Hebdomadis Ab|Leptospira interrogans serovar Hebdomadis Ab
C2923776|T201|COMP|59370-7|LNC|Leptospira interrogans serovar Australis Ab|Leptospira interrogans serovar Australis Ab
C2923777|T201|COMP|59371-5|LNC|Leptospira interrogans serovar Autumnalis Ab|Leptospira interrogans serovar Autumnalis Ab
C2923778|T201|COMP|59372-3|LNC|Leptospira interrogans serovar Ballum Ab|Leptospira interrogans serovar Ballum Ab
C2923786|T201|COMP|59376-4|LNC|3-Keto, 2-Methylvalerate/Creatinine|3-Keto, 2-Methylvalerate/Creatinine
C2923788|T201|COMP|59377-2|LNC|2-Methylacetoacetate/Creatinine|2-Methylacetoacetate/Creatinine
C2923790|T201|COMP|59378-0|LNC|Amikacin^post dialysis|Amikacin^post dialysis
C2923791|T201|COMP|59379-8|LNC|Gentamicin^post dialysis|Gentamicin^post dialysis
C2923792|T201|COMP|59380-6|LNC|Tobramycin^post dialysis|Tobramycin^post dialysis
C2923793|T201|COMP|59381-4|LNC|Vancomycin^post dialysis|Vancomycin^post dialysis
C2923794|T201|COMP|59382-2|LNC|Aspergillus versicolor Ab.IgG|Aspergillus versicolor Ab.IgG
C2923795|T201|COMP|59383-0|LNC|Hydroxyproline/Creatinine|Hydroxyproline/Creatinine
C2923796|T201|COMP|59400-2|LNC|RNA Ab|RNA Ab
C2923797|T201|COMP|59401-0|LNC|Echovirus Ab.IgG|Echovirus Ab.IgG
C2923798|T201|COMP|59402-8|LNC|Mi-1+Mi-2 Ab|Mi-1+Mi-2 Ab
C2923800|T201|COMP|59403-6|LNC|Ku Ab|Ku Ab
C2923801|T201|COMP|59404-4|LNC|Oxygen capacity|Oxygen capacity
C2923816|T201|COMP|59419-2|LNC|HIV 1 RNA|HIV 1 RNA
C2923819|T201|COMP|59421-8|LNC|Neisseria meningitidis serogroups A+B+C+w135+Y Ag|Neisseria meningitidis serogroups A+B+C+w135+Y Ag
C2923821|T201|COMP|59422-6|LNC|Leptospira interrogans serovar Javanica Ab|Leptospira interrogans serovar Javanica Ab
C2923822|T201|COMP|59423-4|LNC|Influenza virus A hemagglutinin type RNA|Influenza virus A hemagglutinin type RNA
C2923824|T201|COMP|59424-2|LNC|Influenza virus A hemagglutinin type RNA|Influenza virus A hemagglutinin type RNA
C2923840|T201|COMP|59462-2|LNC|Clinical biochemist review|Clinical biochemist review
C2923842|T201|COMP|59463-0|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C2923843|T201|COMP|59464-8|LNC|Microbiologist review|Microbiologist review
C2923845|T201|COMP|59465-5|LNC|Pathologist review|Pathologist review
C2923846|T201|COMP|59466-3|LNC|Hematologist review|Hematologist review
C2923849|T201|COMP|59468-9|LNC|Erythrocyte mean corpuscular hemoglobin|Erythrocyte mean corpuscular hemoglobin
C2923851|T201|COMP|59561-1|LNC|Propofol glucuronide|Propofol glucuronide
C2923853|T201|COMP|59562-9|LNC|DNA index|DNA index
C2923856|T201|COMP|59563-7|LNC|Protein.monoclonal band 4|Protein.monoclonal band 4
C2923857|T201|COMP|59564-5|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C2923858|T201|COMP|59565-2|LNC|Netilmicin^trough|Netilmicin^trough
C2923859|T201|COMP|59566-0|LNC|Netilmicin|Netilmicin
C2923860|T201|COMP|59567-8|LNC|Netilmicin^peak|Netilmicin^peak
C2923861|T201|COMP|59568-6|LNC|Orotate|Orotate
C2923862|T201|COMP|59569-4|LNC|Calcitonin^post XXX challenge|Calcitonin^post XXX challenge
C2923863|T201|COMP|59570-2|LNC|Urea nitrogen|Urea nitrogen
C2923864|T201|COMP|59581-9|LNC|Coxsackievirus A7 Ab.IgM|Coxsackievirus A7 Ab.IgM
C2923866|T201|COMP|59582-7|LNC|Coxsackievirus A24 Ab.IgG|Coxsackievirus A24 Ab.IgG
C2923868|T201|COMP|59583-5|LNC|Coxsackievirus A16 Ab.IgG|Coxsackievirus A16 Ab.IgG
C2923870|T201|COMP|59584-3|LNC|Coxsackievirus A7 Ab.IgG|Coxsackievirus A7 Ab.IgG
C2923872|T201|COMP|59585-0|LNC|GSTP1 gene+APC gene methylation|GSTP1 gene+APC gene methylation
C2923874|T201|COMP|59587-6|LNC|Homovanillate|Homovanillate
C2923875|T201|COMP|59588-4|LNC|1-Hydroxymidazolam|1-Hydroxymidazolam
C2923876|T201|COMP|59589-2|LNC|1-Hydroxymidazolam|1-Hydroxymidazolam
C2923877|T201|COMP|59590-0|LNC|1-Hydroxymidazolam|1-Hydroxymidazolam
C2923878|T201|COMP|59591-8|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2923879|T201|COMP|59592-6|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2923880|T201|COMP|59593-4|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2923881|T201|COMP|59594-2|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2923882|T201|COMP|59595-9|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2923883|T201|COMP|59596-7|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2923884|T201|COMP|59597-5|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2923885|T201|COMP|59598-3|LNC|acetaZOLAMIDE|acetaZOLAMIDE
C2923886|T201|COMP|59599-1|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2923887|T201|COMP|59600-7|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2923888|T201|COMP|59601-5|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2923889|T201|COMP|59602-3|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2923890|T201|COMP|59603-1|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2923891|T201|COMP|59604-9|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2923892|T201|COMP|59605-6|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2923893|T201|COMP|59606-4|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2923894|T201|COMP|59607-2|LNC|ALPRAZolam|ALPRAZolam
C2923895|T201|COMP|59608-0|LNC|ALPRAZolam|ALPRAZolam
C2923896|T201|COMP|59609-8|LNC|ALPRAZolam|ALPRAZolam
C2923897|T201|COMP|59610-6|LNC|ALPRAZolam|ALPRAZolam
C2923898|T201|COMP|59611-4|LNC|ALPRAZolam|ALPRAZolam
C2923899|T201|COMP|59612-2|LNC|ALPRAZolam|ALPRAZolam
C2923900|T201|COMP|59613-0|LNC|ALPRAZolam|ALPRAZolam
C2923901|T201|COMP|59614-8|LNC|ALPRAZolam|ALPRAZolam
C2923902|T201|COMP|59615-5|LNC|ALPRAZolam|ALPRAZolam
C2923903|T201|COMP|59616-3|LNC|Benzoylecgonine|Benzoylecgonine
C2923904|T201|COMP|59617-1|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2923905|T201|COMP|59618-9|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2923906|T201|COMP|59619-7|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2923907|T201|COMP|59620-5|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2923908|T201|COMP|59621-3|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2923909|T201|COMP|59622-1|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2923910|T201|COMP|59623-9|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2923911|T201|COMP|59624-7|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2923912|T201|COMP|59625-4|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2923913|T201|COMP|59626-2|LNC|cloBAZam|cloBAZam
C2923914|T201|COMP|59627-0|LNC|cloBAZam|cloBAZam
C2923915|T201|COMP|59628-8|LNC|cloBAZam|cloBAZam
C2923916|T201|COMP|59629-6|LNC|cloBAZam|cloBAZam
C2923917|T201|COMP|59630-4|LNC|cloBAZam|cloBAZam
C2923918|T201|COMP|59631-2|LNC|cloBAZam|cloBAZam
C2923919|T201|COMP|59632-0|LNC|cloBAZam|cloBAZam
C2923920|T201|COMP|59633-8|LNC|cloBAZam|cloBAZam
C2923921|T201|COMP|59634-6|LNC|cloBAZam|cloBAZam
C2923922|T201|COMP|59635-3|LNC|cloBAZam|cloBAZam
C2923923|T201|COMP|59636-1|LNC|clonazePAM|clonazePAM
C2923924|T201|COMP|59637-9|LNC|clonazePAM|clonazePAM
C2923925|T201|COMP|59638-7|LNC|clonazePAM|clonazePAM
C2923926|T201|COMP|59639-5|LNC|clonazePAM|clonazePAM
C2923927|T201|COMP|59640-3|LNC|clonazePAM|clonazePAM
C2923928|T201|COMP|59641-1|LNC|clonazePAM|clonazePAM
C2923929|T201|COMP|59642-9|LNC|clonazePAM|clonazePAM
C2923930|T201|COMP|59643-7|LNC|Cocaethylene|Cocaethylene
C2923931|T201|COMP|59644-5|LNC|Cocaine|Cocaine
C2923932|T201|COMP|59645-2|LNC|Cotinine|Cotinine
C2923933|T201|COMP|59646-0|LNC|Cotinine|Cotinine
C2923934|T201|COMP|59647-8|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2923935|T201|COMP|59648-6|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2923936|T201|COMP|59649-4|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2923937|T201|COMP|59650-2|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2923938|T201|COMP|59651-0|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2923939|T201|COMP|59659-3|LNC|diazePAM|diazePAM
C2923940|T201|COMP|59660-1|LNC|diazePAM|diazePAM
C2923941|T201|COMP|59661-9|LNC|diazePAM|diazePAM
C2923942|T201|COMP|59662-7|LNC|Diclofenac|Diclofenac
C2923943|T201|COMP|59663-5|LNC|Diclofenac|Diclofenac
C2923944|T201|COMP|59664-3|LNC|Estazolam|Estazolam
C2923945|T201|COMP|59665-0|LNC|Estazolam|Estazolam
C2923946|T201|COMP|59666-8|LNC|Estazolam|Estazolam
C2923947|T201|COMP|59667-6|LNC|Estazolam|Estazolam
C2923948|T201|COMP|59668-4|LNC|Estazolam|Estazolam
C2923949|T201|COMP|59669-2|LNC|Estazolam|Estazolam
C2923950|T201|COMP|59670-0|LNC|Estazolam|Estazolam
C2923951|T201|COMP|59671-8|LNC|Estazolam|Estazolam
C2923952|T201|COMP|59672-6|LNC|Estazolam|Estazolam
C2923953|T201|COMP|59683-3|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C2923954|T201|COMP|59684-1|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C2923955|T201|COMP|59685-8|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C2923956|T201|COMP|59686-6|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C2923957|T201|COMP|59687-4|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C2923958|T201|COMP|59688-2|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C2923959|T201|COMP|59689-0|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C2923960|T201|COMP|59690-8|LNC|Hydroxytriazolam|Hydroxytriazolam
C2923961|T201|COMP|59691-6|LNC|Hydroxytriazolam|Hydroxytriazolam
C2923962|T201|COMP|59692-4|LNC|Hydroxytriazolam|Hydroxytriazolam
C2923963|T201|COMP|59693-2|LNC|Hydroxytriazolam|Hydroxytriazolam
C2923964|T201|COMP|59694-0|LNC|Hydroxytriazolam|Hydroxytriazolam
C2923965|T201|COMP|59695-7|LNC|Hydroxytriazolam|Hydroxytriazolam
C2923966|T201|COMP|59696-5|LNC|Hydroxytriazolam|Hydroxytriazolam
C2923967|T201|COMP|59699-9|LNC|LORazepam|LORazepam
C2923968|T201|COMP|59700-5|LNC|LORazepam|LORazepam
C2923969|T201|COMP|59701-3|LNC|LORazepam|LORazepam
C2923970|T201|COMP|59702-1|LNC|LORazepam|LORazepam
C2923971|T201|COMP|59703-9|LNC|LORazepam|LORazepam
C2923972|T201|COMP|59704-7|LNC|LORazepam|LORazepam
C2923973|T201|COMP|59705-4|LNC|Methadone|Methadone
C2923974|T201|COMP|59706-2|LNC|MethylePHEDrine|MethylePHEDrine
C2923975|T201|COMP|59707-0|LNC|Midazolam|Midazolam
C2923976|T201|COMP|59708-8|LNC|Midazolam|Midazolam
C2923977|T201|COMP|59723-7|LNC|Nordiazepam|Nordiazepam
C2923978|T201|COMP|59724-5|LNC|Cathine|Cathine
C2923979|T201|COMP|59725-2|LNC|Oxazepam|Oxazepam
C2923980|T201|COMP|59726-0|LNC|Oxazepam|Oxazepam
C2923981|T201|COMP|59727-8|LNC|Oxazepam|Oxazepam
C2923982|T201|COMP|59728-6|LNC|Oxazepam|Oxazepam
C2923983|T201|COMP|59729-4|LNC|Oxazepam|Oxazepam
C2923984|T201|COMP|59730-2|LNC|Oxazepam|Oxazepam
C2923985|T201|COMP|59731-0|LNC|Oxazepam|Oxazepam
C2923986|T201|COMP|59732-8|LNC|Oxazepam|Oxazepam
C2923987|T201|COMP|59733-6|LNC|Potassium|Potassium
C2923988|T201|COMP|59734-4|LNC|Propoxyphene|Propoxyphene
C2923989|T201|COMP|59735-1|LNC|Salicylamide|Salicylamide
C2923990|T201|COMP|59736-9|LNC|Salicylamide|Salicylamide
C2923991|T201|COMP|59737-7|LNC|Selenium|Selenium
C2923992|T201|COMP|59738-5|LNC|Silver|Silver
C2923993|T201|COMP|59739-3|LNC|Silver|Silver
C2923994|T201|COMP|59740-1|LNC|Silver|Silver
C2923995|T201|COMP|59741-9|LNC|Silver|Silver
C2923996|T201|COMP|59742-7|LNC|sulfADIAZINE|sulfADIAZINE
C2923997|T201|COMP|59743-5|LNC|SUMAtriptan|SUMAtriptan
C2923998|T201|COMP|59744-3|LNC|SUMAtriptan|SUMAtriptan
C2923999|T201|COMP|59745-0|LNC|Temazepam|Temazepam
C2924000|T201|COMP|59746-8|LNC|Temazepam|Temazepam
C2924001|T201|COMP|59747-6|LNC|Temazepam|Temazepam
C2924002|T201|COMP|59748-4|LNC|Temazepam|Temazepam
C2924003|T201|COMP|59749-2|LNC|Temazepam|Temazepam
C2924004|T201|COMP|59750-0|LNC|Temazepam|Temazepam
C2924005|T201|COMP|59751-8|LNC|Temazepam|Temazepam
C2924006|T201|COMP|59752-6|LNC|Temazepam|Temazepam
C2924007|T201|COMP|59753-4|LNC|Titanium|Titanium
C2924008|T201|COMP|59754-2|LNC|Titanium|Titanium
C2924009|T201|COMP|59755-9|LNC|Titanium|Titanium
C2924010|T201|COMP|59756-7|LNC|Titanium|Titanium
C2924011|T201|COMP|59757-5|LNC|tiZANidine|tiZANidine
C2924012|T201|COMP|59758-3|LNC|Triazolam|Triazolam
C2924013|T201|COMP|59759-1|LNC|Triazolam|Triazolam
C2924014|T201|COMP|59760-9|LNC|Triazolam|Triazolam
C2924015|T201|COMP|59761-7|LNC|Triazolam|Triazolam
C2924016|T201|COMP|59762-5|LNC|Triazolam|Triazolam
C2924017|T201|COMP|59763-3|LNC|Triazolam|Triazolam
C2924018|T201|COMP|59764-1|LNC|Triazolam|Triazolam
C2924019|T201|COMP|59765-8|LNC|Tungsten|Tungsten
C2924020|T201|COMP|59766-6|LNC|Tungsten|Tungsten
C2924021|T201|COMP|59767-4|LNC|Ziprasidone|Ziprasidone
C2924048|T201|COMP|59786-4|LNC|Urea/Creatinine|Urea/Creatinine
C2924049|T201|COMP|59787-2|LNC|Catecholamines|Catecholamines
C2924052|T201|COMP|59790-6|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C2924053|T201|COMP|59791-4|LNC|Glucose^30M post XXX challenge|Glucose^30M post XXX challenge
C2924054|T201|COMP|59792-2|LNC|Glucose^1H post XXX challenge|Glucose^1H post XXX challenge
C2924055|T201|COMP|59793-0|LNC|Glucose^1.5H post XXX challenge|Glucose^1.5H post XXX challenge
C2924056|T201|COMP|59794-8|LNC|Glucose^2H post XXX challenge|Glucose^2H post XXX challenge
C2924057|T201|COMP|59795-5|LNC|Glucose^3H post XXX challenge|Glucose^3H post XXX challenge
C2924058|T201|COMP|59796-3|LNC|Glucose^4H post XXX challenge|Glucose^4H post XXX challenge
C2924059|T201|COMP|59797-1|LNC|Glucose^5H post XXX challenge|Glucose^5H post XXX challenge
C2924060|T201|COMP|59798-9|LNC|Ganciclovir^peak|Ganciclovir^peak
C2924061|T201|COMP|59799-7|LNC|Ganciclovir^trough|Ganciclovir^trough
C2924062|T201|COMP|59800-3|LNC|Protein.monoclonal band 2/Protein.total|Protein.monoclonal band 2/Protein.total
C2924063|T201|COMP|59815-1|LNC|Glucose^3 PM specimen|Glucose^3 PM specimen
C2924064|T201|COMP|59816-9|LNC|Neutrophils.immature/100 leukocytes|Neutrophils.immature/100 leukocytes
C2924065|T201|COMP|59817-7|LNC|Uroporphyrin 1 isomer/Creatinine|Uroporphyrin 1 isomer/Creatinine
C2924066|T201|COMP|59818-5|LNC|Uroporphyrin 3 isomer/Creatinine|Uroporphyrin 3 isomer/Creatinine
C2924067|T201|COMP|59819-3|LNC|Pentacarboxylporphyrins/Creatinine|Pentacarboxylporphyrins/Creatinine
C2924068|T201|COMP|59820-1|LNC|Coproporphyrin 1/Creatinine|Coproporphyrin 1/Creatinine
C2924069|T201|COMP|59821-9|LNC|Coproporphyrin 3/Creatinine|Coproporphyrin 3/Creatinine
C2924070|T201|COMP|59822-7|LNC|Tacrolimus^4H post dose|Tacrolimus^4H post dose
C2924071|T201|COMP|59823-5|LNC|Tacrolimus^2H post dose|Tacrolimus^2H post dose
C2924072|T201|COMP|59824-3|LNC|Cyanide|Cyanide
C2924073|T201|COMP|59825-0|LNC|Phenols|Phenols
C2924074|T201|COMP|59826-8|LNC|Creatinine|Creatinine
C2924075|T201|COMP|59827-6|LNC|Bilirubin|Bilirubin
C2924076|T201|COMP|59828-4|LNC|Bilirubin|Bilirubin
C2924077|T201|COMP|59829-2|LNC|Leukocytes|Leukocytes
C2924078|T201|COMP|59830-0|LNC|Erythrocytes|Erythrocytes
C2924079|T201|COMP|59831-8|LNC|Gastrin^baseline|Gastrin^baseline
C2924080|T201|COMP|59832-6|LNC|Gastrin^1st specimen post XXX challenge|Gastrin^1st specimen post XXX challenge
C2924081|T201|COMP|59833-4|LNC|Antibiotic XXX|Antibiotic XXX
C2924082|T201|COMP|59834-2|LNC|Creatinine reduction ratio|Creatinine reduction ratio
C2924083|T201|COMP|59835-9|LNC|Parathyrin.intact|Parathyrin.intact
C2924084|T201|COMP|59836-7|LNC|Mycoplasma sp+Ureaplasma urealyticum DNA|Mycoplasma sp+Ureaplasma urealyticum DNA
C2924086|T201|COMP|59837-5|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C2924087|T201|COMP|59838-3|LNC|Cytomegalovirus Ab|Cytomegalovirus Ab
C2924088|T201|COMP|59839-1|LNC|Urate crystals|Urate crystals
C2924090|T201|COMP|59841-7|LNC|Vendor name|Vendor name
C2924096|T201|COMP|59844-1|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C2925364|T201|COMP|55362-8|LNC|Thyrotropin^pre XXX challenge|Thyrotropin^pre XXX challenge
C2925529|T201|COMP|56522-6|LNC|17-Hydroxypregnenolone^30M post XXX challenge|17-Hydroxypregnenolone^30M post XXX challenge
C2925635|T201|COMP|57366-7|LNC|Lactate^pre XXX challenge|Lactate^pre XXX challenge
C2925636|T201|COMP|57950-8|LNC|Cow whey Ab.IgE/IgE.total|Cow whey Ab.IgE/IgE.total
C2925637|T201|COMP|57952-4|LNC|Cucumis melo spp Ab.IgE/IgE.total|Cucumis melo spp Ab.IgE/IgE.total
C2925638|T201|COMP|56606-7|LNC|11-Deoxycorticosterone^pre XXX challenge|11-Deoxycorticosterone^pre XXX challenge
C2925651|T201|COMP|58812-9|LNC|Renin^3rd specimen|Renin^3rd specimen
C2925652|T201|COMP|58813-7|LNC|Renin^2nd specimen|Renin^2nd specimen
C2925653|T201|COMP|58814-5|LNC|17-Hydroxyprogesterone^3rd specimen|17-Hydroxyprogesterone^3rd specimen
C2925654|T201|COMP|58815-2|LNC|17-Hydroxyprogesterone^2nd specimen|17-Hydroxyprogesterone^2nd specimen
C2925655|T201|COMP|58816-0|LNC|C peptide^2nd specimen|C peptide^2nd specimen
C2925656|T201|COMP|58817-8|LNC|Estradiol^3rd specimen|Estradiol^3rd specimen
C2925657|T201|COMP|58818-6|LNC|Estrogen^2nd specimen|Estrogen^2nd specimen
C2925658|T201|COMP|58819-4|LNC|Cortisol^21st specimen|Cortisol^21st specimen
C2925659|T201|COMP|58820-2|LNC|Cortisol^24th specimen|Cortisol^24th specimen
C2925660|T201|COMP|58821-0|LNC|Cortisol^23rd specimen|Cortisol^23rd specimen
C2925661|T201|COMP|59017-4|LNC|HLA-DPB1|HLA-DPB1
C2925662|T201|COMP|59018-2|LNC|HLA-DPA1|HLA-DPA1
C2925663|T201|COMP|59034-9|LNC|Ganglioside GD2 Ab.IgG|Ganglioside GD2 Ab.IgG
C2925664|T201|COMP|59035-6|LNC|Cells.CD54/100 cells|Cells.CD54/100 cells
C2925665|T201|COMP|59036-4|LNC|Triglyceride|Triglyceride
C2925666|T201|COMP|59037-2|LNC|Phosphate|Phosphate
C2925667|T201|COMP|59038-0|LNC|Cholesterol|Cholesterol
C2925668|T201|COMP|59039-8|LNC|Amylase|Amylase
C2925669|T201|COMP|59040-6|LNC|Cancer Ag 125|Cancer Ag 125
C2925670|T201|COMP|59041-4|LNC|BRCA1+BRCA2 gene mutations tested for|BRCA1+BRCA2 gene mutations tested for
C2925672|T201|COMP|59042-2|LNC|Cells.TCR gamma delta/100 cells|Cells.TCR gamma delta/100 cells
C2925673|T201|COMP|59043-0|LNC|Somatotropin^34th specimen|Somatotropin^34th specimen
C2925674|T201|COMP|59673-4|LNC|fentaNYL|fentaNYL
C2925675|T201|COMP|59674-2|LNC|Flurazepam|Flurazepam
C2925676|T201|COMP|59675-9|LNC|Flurazepam|Flurazepam
C2925677|T201|COMP|59676-7|LNC|Flurazepam|Flurazepam
C2925678|T201|COMP|59677-5|LNC|Flurazepam|Flurazepam
C2925679|T201|COMP|59678-3|LNC|Flurazepam|Flurazepam
C2925680|T201|COMP|59679-1|LNC|Flurazepam|Flurazepam
C2925681|T201|COMP|59680-9|LNC|Gabapentin|Gabapentin
C2925682|T201|COMP|59681-7|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C2925683|T201|COMP|59682-5|LNC|Hydroxyethylflurazepam|Hydroxyethylflurazepam
C2925684|T201|COMP|57912-8|LNC|Bean green Ab.IgE/IgE.total|Bean green Ab.IgE/IgE.total
C2925685|T201|COMP|57913-6|LNC|Bean white Ab.IgE/IgE.total|Bean white Ab.IgE/IgE.total
C2925686|T201|COMP|57914-4|LNC|Beta lactoglobulin Ab.IgE/IgE.total|Beta lactoglobulin Ab.IgE/IgE.total
C2925687|T201|COMP|57915-1|LNC|Bombus terrestris Ab.IgE/IgE.total|Bombus terrestris Ab.IgE/IgE.total
C2925688|T201|COMP|58388-0|LNC|Normeperidine|Normeperidine
C2925689|T201|COMP|58389-8|LNC|Normeperidine|Normeperidine
C2925692|T201|COMP|58391-4|LNC|Codeine/Creatinine|Codeine/Creatinine
C2925694|T201|COMP|58392-2|LNC|Morphine/Creatinine|Morphine/Creatinine
C2925696|T201|COMP|58393-0|LNC|HYDROcodone/Creatinine|HYDROcodone/Creatinine
C2925698|T201|COMP|58394-8|LNC|HYDROmorphone/Creatinine|HYDROmorphone/Creatinine
C2925700|T201|COMP|58395-5|LNC|oxyCODONE/Creatinine|oxyCODONE/Creatinine
C2925702|T201|COMP|58396-3|LNC|oxyMORphone/Creatinine|oxyMORphone/Creatinine
C2925704|T201|COMP|58397-1|LNC|Phencyclidine/Creatinine|Phencyclidine/Creatinine
C2925714|T201|COMP|58751-9|LNC|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C2925715|T201|COMP|58948-1|LNC|Somatotropin^pre XXX challenge|Somatotropin^pre XXX challenge
C2925716|T201|COMP|58949-9|LNC|Somatotropin^12th specimen|Somatotropin^12th specimen
C2925717|T201|COMP|58950-7|LNC|Somatotropin^11th specimen|Somatotropin^11th specimen
C2925718|T201|COMP|58951-5|LNC|Creatinine^2nd specimen|Creatinine^2nd specimen
C2925719|T201|COMP|58952-3|LNC|Testosterone free & total panel|Testosterone free & total panel
C2925720|T201|COMP|58953-1|LNC|Meperidine & Normeperidine panel|Meperidine & Normeperidine panel
C2925721|T201|COMP|58954-9|LNC|Deoxypyridinoline/Pyridinoline|Deoxypyridinoline/Pyridinoline
C2925722|T201|COMP|58955-6|LNC|Pyridinoline & Deoxypyridinoline|Pyridinoline & Deoxypyridinoline
C2925724|T201|COMP|58957-2|LNC|Heparin given|Heparin given
C2925726|T201|COMP|59153-7|LNC|Cortisol^5H post XXX challenge|Cortisol^5H post XXX challenge
C2925727|T201|COMP|59154-5|LNC|Base deficit|Base deficit
C2925728|T201|COMP|59155-2|LNC|17-Hydroxyprogesterone^20M post XXX challenge|17-Hydroxyprogesterone^20M post XXX challenge
C2925729|T201|COMP|59156-0|LNC|Glucose|Glucose
C2925730|T201|COMP|59157-8|LNC|Glucose^pre dose lactose PO|Glucose^pre dose lactose PO
C2925731|T201|COMP|59158-6|LNC|Ketones|Ketones
C2925732|T201|COMP|59159-4|LNC|Albumin/Creatinine|Albumin/Creatinine
C2925733|T201|COMP|59160-2|LNC|Cannabinoids|Cannabinoids
C2925734|T201|COMP|59161-0|LNC|Phosphate|Phosphate
C2925735|T201|COMP|59162-8|LNC|Potassium|Potassium
C2925736|T201|COMP|59163-6|LNC|Sodium|Sodium
C2925737|T201|COMP|57581-1|LNC|Aldosterone^pre XXX challenge|Aldosterone^pre XXX challenge
C2925944|T201|COMP|58484-7|LNC|Estradiol^8th specimen post XXX challenge|Estradiol^8th specimen post XXX challenge
C2925945|T201|COMP|58485-4|LNC|Estradiol^baseline|Estradiol^baseline
C2925946|T201|COMP|58486-2|LNC|Estradiol^7th specimen post XXX challenge|Estradiol^7th specimen post XXX challenge
C2925947|T201|COMP|58487-0|LNC|Estradiol^6th specimen post XXX challenge|Estradiol^6th specimen post XXX challenge
C2925948|T201|COMP|58488-8|LNC|Estradiol^5th specimen post XXX challenge|Estradiol^5th specimen post XXX challenge
C2925949|T201|COMP|58489-6|LNC|Estradiol^4th specimen post XXX challenge|Estradiol^4th specimen post XXX challenge
C2925950|T201|COMP|58490-4|LNC|Estradiol^3rd specimen post XXX challenge|Estradiol^3rd specimen post XXX challenge
C2925951|T201|COMP|58491-2|LNC|Estradiol^2nd specimen post XXX challenge|Estradiol^2nd specimen post XXX challenge
C2925952|T201|COMP|58492-0|LNC|Estradiol^1st specimen post XXX challenge|Estradiol^1st specimen post XXX challenge
C2925953|T201|COMP|58493-8|LNC|Coagulation factor VIII Ab|Coagulation factor VIII Ab
C2925954|T201|COMP|58494-6|LNC|C peptide^1.5H post dose glucose|C peptide^1.5H post dose glucose
C2925955|T201|COMP|58495-3|LNC|C peptide^10M post 1 mg glucagon IV|C peptide^10M post 1 mg glucagon IV
C2925956|T201|COMP|57925-0|LNC|Castanea sativa Ab.IgE/IgE.total|Castanea sativa Ab.IgE/IgE.total
C2925957|T201|COMP|57932-6|LNC|Cheese cheddar type Ab.IgE/IgE.total|Cheese cheddar type Ab.IgE/IgE.total
C2925958|T201|COMP|57933-4|LNC|Cheese mold type Ab.IgE/IgE.total|Cheese mold type Ab.IgE/IgE.total
C2925959|T201|COMP|57935-9|LNC|Chocolate Ab.IgE/IgE.total|Chocolate Ab.IgE/IgE.total
C2925960|T201|COMP|57940-9|LNC|Citrullus lanatus Ab.IgE/IgE.total|Citrullus lanatus Ab.IgE/IgE.total
C2925961|T201|COMP|57941-7|LNC|Citrus aurantifolia Ab.IgE/IgE.total|Citrus aurantifolia Ab.IgE/IgE.total
C2925962|T201|COMP|57947-4|LNC|Coffee bean Ab.IgE.RAST class|Coffee bean Ab.IgE.RAST class
C2925964|T201|COMP|57987-0|LNC|Ipomoea batatas Ab.IgE/IgE.total|Ipomoea batatas Ab.IgE/IgE.total
C2925965|T201|COMP|57991-2|LNC|Lactalbumin Ab.IgE/IgE.total|Lactalbumin Ab.IgE/IgE.total
C2925967|T201|COMP|57993-8|LNC|Lepidoglyphus destructor Ab.IgE/IgE.total|Lepidoglyphus destructor Ab.IgE/IgE.total
C2925968|T201|COMP|58000-1|LNC|Maple sugar Ab.IgE/IgE.total|Maple sugar Ab.IgE/IgE.total
C2925969|T201|COMP|58017-5|LNC|Olea europaea pollen Ab.IgE/IgE.total|Olea europaea pollen Ab.IgE/IgE.total
C2925970|T201|COMP|58025-8|LNC|Secale cereale pollen Ab.IgE/IgE.total|Secale cereale pollen Ab.IgE/IgE.total
C2925971|T201|COMP|58033-2|LNC|Urtica dioica Ab.IgE/IgE.total|Urtica dioica Ab.IgE/IgE.total
C2925972|T201|COMP|58034-0|LNC|Ustilago cynodontis Ab.IgE/IgE.total|Ustilago cynodontis Ab.IgE/IgE.total
C2925973|T201|COMP|58043-1|LNC|Platanus occidentalis Ab.IgE/IgE.total|Platanus occidentalis Ab.IgE/IgE.total
C2925974|T201|COMP|58449-0|LNC|Erythrocyte clumps|Erythrocyte clumps
C2925975|T201|COMP|58450-8|LNC|Bilirubin|Bilirubin
C2925976|T201|COMP|58451-6|LNC|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C2925977|T201|COMP|58452-4|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C2925978|T201|COMP|58453-2|LNC|Hemoglobin.gastrointestinal.lower|Hemoglobin.gastrointestinal.lower
C2925979|T201|COMP|58454-0|LNC|Subtelomere analysis|Subtelomere analysis
C2925980|T201|COMP|58455-7|LNC|Taenia solium Ab|Taenia solium Ab
C2925981|T201|COMP|58456-5|LNC|Bladder cells|Bladder cells
C2925982|T201|COMP|58457-3|LNC|Sulfites|Sulfites
C2925983|T201|COMP|58458-1|LNC|Mitochondria Ab pattern|Mitochondria Ab pattern
C2925985|T201|COMP|58459-9|LNC|Ganglioside GT1b Ab|Ganglioside GT1b Ab
C2925986|T201|COMP|58460-7|LNC|Endothelial cell Ab|Endothelial cell Ab
C2925987|T201|COMP|58461-5|LNC|Intestinal goblet cell Ab|Intestinal goblet cell Ab
C2925988|T201|COMP|58462-3|LNC|Complement functional activity|Complement functional activity
C2925993|T201|COMP|58732-9|LNC|Porphyrin fractions panel|Porphyrin fractions panel
C2925994|T201|COMP|58733-7|LNC|Mycoplasma pneumoniae Ab.IgG & IgM panel|Mycoplasma pneumoniae Ab.IgG & IgM panel
C2925995|T201|COMP|58734-5|LNC|Collection date|Collection date
C2925996|T201|COMP|58735-2|LNC|Alpha-1-fetoprotein panel|Alpha-1-fetoprotein panel
C2925997|T201|COMP|58736-0|LNC|Manganese panel|Manganese panel
C2925998|T201|COMP|58875-6|LNC|Somatotropin^32nd specimen|Somatotropin^32nd specimen
C2925999|T201|COMP|58876-4|LNC|Somatotropin^31st specimen|Somatotropin^31st specimen
C2926000|T201|COMP|58877-2|LNC|Somatotropin^30th specimen|Somatotropin^30th specimen
C2926001|T201|COMP|58878-0|LNC|Somatotropin^29th specimen|Somatotropin^29th specimen
C2926002|T201|COMP|58879-8|LNC|Somatotropin^28th specimen|Somatotropin^28th specimen
C2926003|T201|COMP|58880-6|LNC|Somatotropin^27th specimen|Somatotropin^27th specimen
C2926004|T201|COMP|58881-4|LNC|Somatotropin^26th specimen|Somatotropin^26th specimen
C2926005|T201|COMP|59019-0|LNC|HLA-DQA1|HLA-DQA1
C2926006|T201|COMP|59024-0|LNC|Renin^supine+30M post XXX challenge|Renin^supine+30M post XXX challenge
C2926007|T201|COMP|59025-7|LNC|Neutrophil Ab|Neutrophil Ab
C2926008|T201|COMP|59026-5|LNC|U1 small nuclear ribonucleoprotein 70kD Ab|U1 small nuclear ribonucleoprotein 70kD Ab
C2926009|T201|COMP|59027-3|LNC|Asialoganglioside GM1 Ab.IgM|Asialoganglioside GM1 Ab.IgM
C2926010|T201|COMP|59028-1|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C2926011|T201|COMP|59029-9|LNC|HLA-DRB1*15:01|HLA-DRB1*15:01
C2926012|T201|COMP|59030-7|LNC|Cells.CD45+CD103+/100 cells|Cells.CD45+CD103+/100 cells
C2926014|T201|COMP|59031-5|LNC|Cells.CD25+C69+/100 cells|Cells.CD25+C69+/100 cells
C2926016|T201|COMP|59032-3|LNC|Lactate|Lactate
C2926017|T201|COMP|59033-1|LNC|Ganglioside GM3 Ab.IgG|Ganglioside GM3 Ab.IgG
C2926027|T201|COMP|58540-6|LNC|Corticotropin^11th specimen post XXX challenge|Corticotropin^11th specimen post XXX challenge
C2926028|T201|COMP|58541-4|LNC|Corticotropin^11th specimen post XXX challenge|Corticotropin^11th specimen post XXX challenge
C2926029|T201|COMP|58542-2|LNC|Corticotropin^12 AM specimen|Corticotropin^12 AM specimen
C2926030|T201|COMP|58543-0|LNC|Corticotropin^12 PM specimen|Corticotropin^12 PM specimen
C2926031|T201|COMP|58544-8|LNC|Corticotropin^12th specimen post XXX challenge|Corticotropin^12th specimen post XXX challenge
C2926032|T201|COMP|58545-5|LNC|Corticotropin^12th specimen post XXX challenge|Corticotropin^12th specimen post XXX challenge
C2926033|T201|COMP|58546-3|LNC|Corticotropin^15M post 1 ug/kg CRH IV|Corticotropin^15M post 1 ug/kg CRH IV
C2926034|T201|COMP|58685-9|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C2926035|T201|COMP|58686-7|LNC|C peptide^2H post dose glucose|C peptide^2H post dose glucose
C2926036|T201|COMP|58687-5|LNC|Corticotropin^9th specimen post XXX challenge|Corticotropin^9th specimen post XXX challenge
C2926037|T201|COMP|58688-3|LNC|Cortisol^11th specimen post XXX challenge|Cortisol^11th specimen post XXX challenge
C2926038|T201|COMP|58689-1|LNC|Cortisol^11th specimen post XXX challenge|Cortisol^11th specimen post XXX challenge
C2926039|T201|COMP|58690-9|LNC|Cortisol^12th specimen post XXX challenge|Cortisol^12th specimen post XXX challenge
C2926040|T201|COMP|58691-7|LNC|Cortisol^12th specimen post XXX challenge|Cortisol^12th specimen post XXX challenge
C2926041|T201|COMP|58692-5|LNC|Cortisol^5th specimen post XXX challenge|Cortisol^5th specimen post XXX challenge
C2926042|T201|COMP|58693-3|LNC|Cortisol^6th specimen post XXX challenge|Cortisol^6th specimen post XXX challenge
C2926043|T201|COMP|58694-1|LNC|Cortisol^7th specimen post XXX challenge|Cortisol^7th specimen post XXX challenge
C2926044|T201|COMP|58695-8|LNC|Cortisol^8th specimen post XXX challenge|Cortisol^8th specimen post XXX challenge
C2926045|T201|COMP|58696-6|LNC|Cortisol^8th specimen post XXX challenge|Cortisol^8th specimen post XXX challenge
C2926046|T201|COMP|58697-4|LNC|Cortisol^9th specimen post XXX challenge|Cortisol^9th specimen post XXX challenge
C2926047|T201|COMP|58698-2|LNC|Cortisol^9th specimen post XXX challenge|Cortisol^9th specimen post XXX challenge
C2926048|T201|COMP|58840-0|LNC|Triiodothyronine.free^baseline|Triiodothyronine.free^baseline
C2926049|T201|COMP|58841-8|LNC|C peptide^5M post XXX challenge|C peptide^5M post XXX challenge
C2926050|T201|COMP|58842-6|LNC|Somatotropin^25th specimen|Somatotropin^25th specimen
C2926051|T201|COMP|58843-4|LNC|Somatotropin^24th specimen|Somatotropin^24th specimen
C2926052|T201|COMP|58844-2|LNC|Somatotropin^20th specimen|Somatotropin^20th specimen
C2926053|T201|COMP|58845-9|LNC|Somatotropin^19th specimen|Somatotropin^19th specimen
C2926109|T201|COMP|58348-4|LNC|MethylePHEDrine|MethylePHEDrine
C2926111|T201|COMP|58350-0|LNC|Plasma cells.immature/100 cells|Plasma cells.immature/100 cells
C2926112|T201|COMP|58351-8|LNC|Connective tissue growth factor|Connective tissue growth factor
C2926113|T201|COMP|58352-6|LNC|Connective tissue growth factor|Connective tissue growth factor
C2926114|T201|COMP|58355-9|LNC|Plasma cells.immature|Plasma cells.immature
C2926115|T201|COMP|58356-7|LNC|Ethanol/Creatinine|Ethanol/Creatinine
C2926117|T201|COMP|58358-3|LNC|Methamphetamine/Creatinine|Methamphetamine/Creatinine
C2926119|T201|COMP|58359-1|LNC|Buprenorphine+Norbuprenorphine|Buprenorphine+Norbuprenorphine
C2926120|T201|COMP|58360-9|LNC|Buprenorphine/Creatinine|Buprenorphine/Creatinine
C2926122|T201|COMP|58361-7|LNC|Norbuprenorphine/Creatinine|Norbuprenorphine/Creatinine
C2926124|T201|COMP|58362-5|LNC|Norbuprenorphine|Norbuprenorphine
C2926125|T201|COMP|58363-3|LNC|Alpha hydroxyalprazolam/Creatinine|Alpha hydroxyalprazolam/Creatinine
C2926127|T201|COMP|58364-1|LNC|7-Aminoclonazepam/Creatinine|7-Aminoclonazepam/Creatinine
C2926129|T201|COMP|58365-8|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2926130|T201|COMP|58366-6|LNC|LORazepam/Creatinine|LORazepam/Creatinine
C2926132|T201|COMP|58367-4|LNC|Nordiazepam/Creatinine|Nordiazepam/Creatinine
C2926134|T201|COMP|58368-2|LNC|Oxazepam/Creatinine|Oxazepam/Creatinine
C2926136|T201|COMP|58369-0|LNC|Temazepam/Creatinine|Temazepam/Creatinine
C2926138|T201|COMP|58370-8|LNC|Carisoprodol+Meprobamate|Carisoprodol+Meprobamate
C2926139|T201|COMP|58371-6|LNC|Carisoprodol/Creatinine|Carisoprodol/Creatinine
C2926141|T201|COMP|58372-4|LNC|Meprobamate/Creatinine|Meprobamate/Creatinine
C2926143|T201|COMP|58373-2|LNC|Meprobamate|Meprobamate
C2926144|T201|COMP|58374-0|LNC|Meprobamate|Meprobamate
C2926145|T201|COMP|58375-7|LNC|Ethyl glucuronide|Ethyl glucuronide
C2926146|T201|COMP|58376-5|LNC|Ethyl glucuronide/Creatinine|Ethyl glucuronide/Creatinine
C2926148|T201|COMP|58377-3|LNC|Ethyl glucuronide|Ethyl glucuronide
C2926149|T201|COMP|58378-1|LNC|Ethyl glucuronide|Ethyl glucuronide
C2926150|T201|COMP|58379-9|LNC|Fentanyl+Norfentanyl|Fentanyl+Norfentanyl
C2926151|T201|COMP|58380-7|LNC|fentaNYL/Creatinine|fentaNYL/Creatinine
C2926153|T201|COMP|58381-5|LNC|fentaNYL|fentaNYL
C2926154|T201|COMP|58382-3|LNC|Norfentanyl/Creatinine|Norfentanyl/Creatinine
C2926156|T201|COMP|58383-1|LNC|Norfentanyl|Norfentanyl
C2926157|T201|COMP|58384-9|LNC|6-Monoacetylmorphine/Creatinine|6-Monoacetylmorphine/Creatinine
C2926159|T201|COMP|58385-6|LNC|Meperidine+Normeperidine|Meperidine+Normeperidine
C2926160|T201|COMP|58386-4|LNC|Meperidine/Creatinine|Meperidine/Creatinine
C2926162|T201|COMP|58387-2|LNC|Normeperidine/Creatinine|Normeperidine/Creatinine
C2926164|T201|COMP|58398-9|LNC|Propoxyphene/Creatinine|Propoxyphene/Creatinine
C2926166|T201|COMP|58399-7|LNC|Norpropoxyphene/Creatinine|Norpropoxyphene/Creatinine
C2926168|T201|COMP|58400-3|LNC|Specimen pH acceptable|Specimen pH acceptable
C2926169|T201|COMP|58401-1|LNC|Tapentadol|Tapentadol
C2926170|T201|COMP|58402-9|LNC|Tapentadol|Tapentadol
C2926171|T201|COMP|58403-7|LNC|Tricyclic antidepressants/Creatinine|Tricyclic antidepressants/Creatinine
C2926173|T201|COMP|58404-5|LNC|traMADol/Creatinine|traMADol/Creatinine
C2926175|T201|COMP|58405-2|LNC|Hepatitis B virus surface Ab Signal/Cutoff|Hepatitis B virus surface Ab Signal/Cutoff
C2926176|T201|COMP|58406-0|LNC|Platelet morphology panel|Platelet morphology panel
C2926177|T201|COMP|58407-8|LNC|Leukocyte morphology panel|Leukocyte morphology panel
C2926178|T201|COMP|58408-6|LNC|Erythrocyte morphology panel|Erythrocyte morphology panel
C2926179|T201|COMP|58409-4|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C2926180|T201|COMP|58410-2|LNC|Complete blood count (hemogram) panel|Complete blood count (hemogram) panel
C2926181|T201|COMP|58411-0|LNC|Clinical research drug XXX|Clinical research drug XXX
C2926182|T201|COMP|58412-8|LNC|Cefepime|Cefepime
C2926183|T201|COMP|58413-6|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C2926184|T201|COMP|58414-4|LNC|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C2926185|T201|COMP|58415-1|LNC|BRAF gene.p.Val600Glu|BRAF gene.p.Val600Glu
C2926186|T201|COMP|58416-9|LNC|MLH1 gene methylation|MLH1 gene methylation
C2926187|T201|COMP|58417-7|LNC|dilTIAZem|dilTIAZem
C2926188|T201|COMP|58418-5|LNC|Micafungin|Micafungin
C2926189|T201|COMP|58419-3|LNC|Caspofungin|Caspofungin
C2926190|T201|COMP|58420-1|LNC|Anidulafungin|Anidulafungin
C2926193|T201|COMP|58423-5|LNC|Ethyl sulfate/Creatinine|Ethyl sulfate/Creatinine
C2926195|T201|COMP|58424-3|LNC|Ethyl sulfate|Ethyl sulfate
C2926196|T201|COMP|58425-0|LNC|Ethyl sulfate|Ethyl sulfate
C2926197|T201|COMP|58426-8|LNC|Carisoprodol|Carisoprodol
C2926198|T201|COMP|58427-6|LNC|Carisoprodol|Carisoprodol
C2926199|T201|COMP|58428-4|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C2926200|T201|COMP|58429-2|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C2926201|T201|COMP|58430-0|LNC|oxyCODONE+Oxymorphone|oxyCODONE+Oxymorphone
C2926202|T201|COMP|58431-8|LNC|Microalbumin panel|Microalbumin panel
C2926203|T201|COMP|58432-6|LNC|Casts panel|Casts panel
C2926204|T201|COMP|58433-4|LNC|Crystals panel|Crystals panel
C2926205|T201|COMP|58434-2|LNC|Cells panel|Cells panel
C2926206|T201|COMP|58435-9|LNC|Microorganisms panel|Microorganisms panel
C2926207|T201|COMP|58436-7|LNC|Casts|Casts
C2926208|T201|COMP|58437-5|LNC|Microorganisms seen|Microorganisms seen
C2926209|T201|COMP|58438-3|LNC|Cells|Cells
C2926210|T201|COMP|58439-1|LNC|Clinical research drug XXX|Clinical research drug XXX
C2926211|T201|COMP|58440-9|LNC|Classical swine fever virus E2 Ab|Classical swine fever virus E2 Ab
C2926212|T201|COMP|58441-7|LNC|Other elements|Other elements
C2926213|T201|COMP|58442-5|LNC|Other elements|Other elements
C2926214|T201|COMP|58443-3|LNC|Other cells|Other cells
C2926215|T201|COMP|58444-1|LNC|Erythrocytes.dysmorphic|Erythrocytes.dysmorphic
C2926216|T201|COMP|58445-8|LNC|Manual differential comment|Manual differential comment
C2926218|T201|COMP|58447-4|LNC|Microalbumin/Creatinine ratio panel|Microalbumin/Creatinine ratio panel
C2926219|T201|COMP|58448-2|LNC|Albumin ug/min|Albumin ug/min
C2926220|T201|COMP|58463-1|LNC|Tau protein/Protein.total|Tau protein/Protein.total
C2926222|T201|COMP|58464-9|LNC|Campesterol|Campesterol
C2926223|T201|COMP|58465-6|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C2926224|T201|COMP|58466-4|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C2926225|T201|COMP|58467-2|LNC|Gasterophilus intestinalis Ab.IgG4|Gasterophilus intestinalis Ab.IgG4
C2926227|T201|COMP|58468-0|LNC|Pimpinella anisum Ab.IgG4|Pimpinella anisum Ab.IgG4
C2926229|T201|COMP|58470-6|LNC|Nucleated cells|Nucleated cells
C2926230|T201|COMP|58471-4|LNC|Erythrocytes.pitted/Erythrocytes.total|Erythrocytes.pitted/Erythrocytes.total
C2926232|T201|COMP|58473-0|LNC|Haemophilus influenzae serotype DNA|Haemophilus influenzae serotype DNA
C2926237|T201|COMP|58478-9|LNC|Bombus sp Ab.IgG|Bombus sp Ab.IgG
C2926238|T201|COMP|58479-7|LNC|Fatty acids.nonesterified^7th specimen post CFst|Fatty acids.nonesterified^7th specimen post CFst
C2926239|T201|COMP|58480-5|LNC|Fatty acids.nonesterified^6th specimen post CFst|Fatty acids.nonesterified^6th specimen post CFst
C2926240|T201|COMP|58481-3|LNC|Protein C Ag/Coagulation factor IX Ag|Protein C Ag/Coagulation factor IX Ag
C2926242|T201|COMP|58482-1|LNC|Protein S Ag/Coagulation factor IX Ag|Protein S Ag/Coagulation factor IX Ag
C2926244|T201|COMP|58483-9|LNC|BRAF gene targeted mutation analysis|BRAF gene targeted mutation analysis
C2926245|T201|COMP|58496-1|LNC|C peptide^10th specimen post XXX challenge|C peptide^10th specimen post XXX challenge
C2926246|T201|COMP|58497-9|LNC|C peptide^11th specimen post XXX challenge|C peptide^11th specimen post XXX challenge
C2926247|T201|COMP|58498-7|LNC|C peptide^12th specimen post XXX challenge|C peptide^12th specimen post XXX challenge
C2926248|T201|COMP|58499-5|LNC|C peptide^15M post 1 mg glucagon IV|C peptide^15M post 1 mg glucagon IV
C2926249|T201|COMP|58500-0|LNC|C peptide^15M post dose glucose|C peptide^15M post dose glucose
C2926250|T201|COMP|58501-8|LNC|C peptide^15M pre XXX challenge|C peptide^15M pre XXX challenge
C2926251|T201|COMP|58502-6|LNC|C peptide^15M pre XXX challenge|C peptide^15M pre XXX challenge
C2926252|T201|COMP|58503-4|LNC|C peptide^1H post dose glucose|C peptide^1H post dose glucose
C2926253|T201|COMP|58504-2|LNC|C peptide^1st specimen post XXX challenge|C peptide^1st specimen post XXX challenge
C2926254|T201|COMP|58505-9|LNC|C peptide^2.5H post dose glucose|C peptide^2.5H post dose glucose
C2926255|T201|COMP|58506-7|LNC|C peptide^2.5H post dose glucose|C peptide^2.5H post dose glucose
C2926256|T201|COMP|58507-5|LNC|C peptide^2M post 1 mg glucagon IV|C peptide^2M post 1 mg glucagon IV
C2926257|T201|COMP|58508-3|LNC|C peptide^3.5H post dose glucose|C peptide^3.5H post dose glucose
C2926258|T201|COMP|58509-1|LNC|C peptide^3.5H post dose glucose|C peptide^3.5H post dose glucose
C2926259|T201|COMP|58510-9|LNC|C peptide^30M post dose glucose|C peptide^30M post dose glucose
C2926260|T201|COMP|58511-7|LNC|C peptide^3H post dose glucose|C peptide^3H post dose glucose
C2926261|T201|COMP|58512-5|LNC|C peptide^4.5H post dose glucose|C peptide^4.5H post dose glucose
C2926262|T201|COMP|58513-3|LNC|C peptide^4.5H post dose glucose|C peptide^4.5H post dose glucose
C2926263|T201|COMP|58514-1|LNC|C peptide^45M post dose glucose|C peptide^45M post dose glucose
C2926264|T201|COMP|58515-8|LNC|C peptide^45M post dose glucose|C peptide^45M post dose glucose
C2926265|T201|COMP|58516-6|LNC|C peptide^4H post dose glucose|C peptide^4H post dose glucose
C2926266|T201|COMP|58517-4|LNC|C peptide^4H post dose glucose|C peptide^4H post dose glucose
C2926267|T201|COMP|58518-2|LNC|C peptide^5H post dose glucose|C peptide^5H post dose glucose
C2926268|T201|COMP|58519-0|LNC|C peptide^5H post dose glucose|C peptide^5H post dose glucose
C2926269|T201|COMP|58520-8|LNC|C peptide^5M post 1 mg glucagon IV|C peptide^5M post 1 mg glucagon IV
C2926270|T201|COMP|58521-6|LNC|C peptide^9th specimen post XXX challenge|C peptide^9th specimen post XXX challenge
C2926271|T201|COMP|58522-4|LNC|C peptide^pre dose glucose|C peptide^pre dose glucose
C2926272|T201|COMP|58523-2|LNC|Corticosterone^30M post 250 ug corticotropin|Corticosterone^30M post 250 ug corticotropin
C2926273|T201|COMP|58524-0|LNC|Corticosterone^1H post 250 ug corticotropin|Corticosterone^1H post 250 ug corticotropin
C2926274|T201|COMP|58525-7|LNC|Corticosterone^pre 250 ug corticotropin|Corticosterone^pre 250 ug corticotropin
C2926275|T201|COMP|58526-5|LNC|Corticotropin^1.5H post dose glucagon|Corticotropin^1.5H post dose glucagon
C2926276|T201|COMP|58527-3|LNC|Corticotropin^1.5H post dose glucagon|Corticotropin^1.5H post dose glucagon
C2926277|T201|COMP|58528-1|LNC|Corticotropin^1.5H post dose glucose|Corticotropin^1.5H post dose glucose
C2926278|T201|COMP|58529-9|LNC|Corticotropin^1.5H post dose glucose|Corticotropin^1.5H post dose glucose
C2926279|T201|COMP|58530-7|LNC|Corticotropin^1.5H post 1 ug/kg CRH IV|Corticotropin^1.5H post 1 ug/kg CRH IV
C2926280|T201|COMP|58531-5|LNC|Corticotropin^1.5H post dose insulin IV|Corticotropin^1.5H post dose insulin IV
C2926281|T201|COMP|58532-3|LNC|Corticotropin^10 AM specimen|Corticotropin^10 AM specimen
C2926282|T201|COMP|58533-1|LNC|Corticotropin^10 AM specimen|Corticotropin^10 AM specimen
C2926283|T201|COMP|58534-9|LNC|Corticotropin^10 PM specimen|Corticotropin^10 PM specimen
C2926284|T201|COMP|58535-6|LNC|Corticotropin^10 PM specimen|Corticotropin^10 PM specimen
C2926285|T201|COMP|58536-4|LNC|Corticotropin^105M post dose insulin IV|Corticotropin^105M post dose insulin IV
C2926286|T201|COMP|58537-2|LNC|Corticotropin^105M post dose insulin IV|Corticotropin^105M post dose insulin IV
C2926287|T201|COMP|58538-0|LNC|Corticotropin^10th specimen post XXX challenge|Corticotropin^10th specimen post XXX challenge
C2926288|T201|COMP|58539-8|LNC|Corticotropin^10th specimen post XXX challenge|Corticotropin^10th specimen post XXX challenge
C2926289|T201|COMP|58547-1|LNC|Corticotropin^15M post dose insulin IV|Corticotropin^15M post dose insulin IV
C2926290|T201|COMP|58548-9|LNC|Corticotropin^15M post dose insulin IV|Corticotropin^15M post dose insulin IV
C2926291|T201|COMP|58549-7|LNC|Corticotropin^15M post XXX challenge|Corticotropin^15M post XXX challenge
C2926292|T201|COMP|58550-5|LNC|Corticotropin^15M pre 1 ug/kg CRH IV|Corticotropin^15M pre 1 ug/kg CRH IV
C2926293|T201|COMP|58551-3|LNC|Corticotropin^15M pre dose insulin IV|Corticotropin^15M pre dose insulin IV
C2926294|T201|COMP|58552-1|LNC|Corticotropin^15M pre dose insulin IV|Corticotropin^15M pre dose insulin IV
C2926295|T201|COMP|58553-9|LNC|Corticotropin^1H post 1 ug/kg CRH IV|Corticotropin^1H post 1 ug/kg CRH IV
C2926296|T201|COMP|58554-7|LNC|Corticotropin^1H post dose glucagon|Corticotropin^1H post dose glucagon
C2926297|T201|COMP|58555-4|LNC|Corticotropin^1H post dose glucagon|Corticotropin^1H post dose glucagon
C2926298|T201|COMP|58556-2|LNC|Corticotropin^1H post dose glucose|Corticotropin^1H post dose glucose
C2926299|T201|COMP|58557-0|LNC|Corticotropin^1H post dose glucose|Corticotropin^1H post dose glucose
C2926300|T201|COMP|58558-8|LNC|Corticotropin^1H post dose insulin IV|Corticotropin^1H post dose insulin IV
C2926301|T201|COMP|58559-6|LNC|Corticotropin^1H post XXX challenge|Corticotropin^1H post XXX challenge
C2926302|T201|COMP|58560-4|LNC|Corticotropin^1st specimen post XXX challenge|Corticotropin^1st specimen post XXX challenge
C2926303|T201|COMP|58561-2|LNC|Corticotropin^2 PM specimen|Corticotropin^2 PM specimen
C2926304|T201|COMP|58562-0|LNC|Corticotropin^2 PM specimen|Corticotropin^2 PM specimen
C2926305|T201|COMP|58563-8|LNC|Corticotropin^2.5H post dose glucagon|Corticotropin^2.5H post dose glucagon
C2926306|T201|COMP|58564-6|LNC|Corticotropin^2.5H post dose glucagon|Corticotropin^2.5H post dose glucagon
C2926307|T201|COMP|58565-3|LNC|Corticotropin^2.5H post dose insulin IV|Corticotropin^2.5H post dose insulin IV
C2926308|T201|COMP|58566-1|LNC|Corticotropin^2.5H post dose insulin IV|Corticotropin^2.5H post dose insulin IV
C2926309|T201|COMP|58567-9|LNC|Corticotropin^2.5H post dose glucose|Corticotropin^2.5H post dose glucose
C2926310|T201|COMP|58568-7|LNC|Corticotropin^2.5H post dose glucose|Corticotropin^2.5H post dose glucose
C2926311|T201|COMP|58569-5|LNC|Corticotropin^1D post dose metyraPONE|Corticotropin^1D post dose metyraPONE
C2926312|T201|COMP|58570-3|LNC|Corticotropin^1D post dose metyraPONE|Corticotropin^1D post dose metyraPONE
C2926313|T201|COMP|58571-1|LNC|Corticotropin^2H post 1 ug/kg CRH IV|Corticotropin^2H post 1 ug/kg CRH IV
C2926314|T201|COMP|58572-9|LNC|Corticotropin^2H post dose glucagon|Corticotropin^2H post dose glucagon
C2926315|T201|COMP|58573-7|LNC|Corticotropin^2H post dose glucagon|Corticotropin^2H post dose glucagon
C2926316|T201|COMP|58574-5|LNC|Corticotropin^2H post dose glucose|Corticotropin^2H post dose glucose
C2926317|T201|COMP|58575-2|LNC|Corticotropin^2H post dose glucose|Corticotropin^2H post dose glucose
C2926318|T201|COMP|58576-0|LNC|Corticotropin^2H post dose insulin IV|Corticotropin^2H post dose insulin IV
C2926319|T201|COMP|58577-8|LNC|Corticotropin^2H post dose insulin IV|Corticotropin^2H post dose insulin IV
C2926320|T201|COMP|58578-6|LNC|Corticotropin^2H post XXX challenge|Corticotropin^2H post XXX challenge
C2926321|T201|COMP|58579-4|LNC|Corticotropin^2nd specimen post XXX challenge|Corticotropin^2nd specimen post XXX challenge
C2926322|T201|COMP|58580-2|LNC|Corticotropin^30M post 1 ug/kg CRH IV|Corticotropin^30M post 1 ug/kg CRH IV
C2926323|T201|COMP|58581-0|LNC|Corticotropin^30M post dose glucagon|Corticotropin^30M post dose glucagon
C2926324|T201|COMP|58582-8|LNC|Corticotropin^30M post dose glucagon|Corticotropin^30M post dose glucagon
C2926325|T201|COMP|58583-6|LNC|Corticotropin^30M post dose glucose|Corticotropin^30M post dose glucose
C2926326|T201|COMP|58584-4|LNC|Corticotropin^30M post dose glucose|Corticotropin^30M post dose glucose
C2926327|T201|COMP|58585-1|LNC|Corticotropin^30M post dose insulin IV|Corticotropin^30M post dose insulin IV
C2926328|T201|COMP|58586-9|LNC|Corticotropin^30M post XXX challenge|Corticotropin^30M post XXX challenge
C2926329|T201|COMP|58587-7|LNC|Corticotropin^30M pre 1 ug/kg CRH IV|Corticotropin^30M pre 1 ug/kg CRH IV
C2926330|T201|COMP|58588-5|LNC|Corticotropin^30M pre 1 ug/kg CRH IV|Corticotropin^30M pre 1 ug/kg CRH IV
C2926331|T201|COMP|58589-3|LNC|Corticotropin^30M pre dose glucagon|Corticotropin^30M pre dose glucagon
C2926332|T201|COMP|58590-1|LNC|Corticotropin^30M pre dose glucagon|Corticotropin^30M pre dose glucagon
C2926333|T201|COMP|58591-9|LNC|Corticotropin^30M pre dose insulin IV|Corticotropin^30M pre dose insulin IV
C2926334|T201|COMP|58592-7|LNC|Corticotropin^30M pre XXX challenge|Corticotropin^30M pre XXX challenge
C2926335|T201|COMP|58593-5|LNC|Corticotropin^30M pre XXX challenge|Corticotropin^30M pre XXX challenge
C2926336|T201|COMP|58594-3|LNC|Corticotropin^3H post dose glucagon|Corticotropin^3H post dose glucagon
C2926337|T201|COMP|58595-0|LNC|Corticotropin^3H post dose glucagon|Corticotropin^3H post dose glucagon
C2926338|T201|COMP|58596-8|LNC|Corticotropin^3H post dose glucose|Corticotropin^3H post dose glucose
C2926339|T201|COMP|58597-6|LNC|Corticotropin^3H post dose glucose|Corticotropin^3H post dose glucose
C2926340|T201|COMP|58598-4|LNC|Corticotropin^3H post dose insulin IV|Corticotropin^3H post dose insulin IV
C2926341|T201|COMP|58599-2|LNC|Corticotropin^3H post dose insulin IV|Corticotropin^3H post dose insulin IV
C2926342|T201|COMP|58600-8|LNC|Corticotropin^3H post XXX challenge|Corticotropin^3H post XXX challenge
C2926343|T201|COMP|58601-6|LNC|Corticotropin^3H post XXX challenge|Corticotropin^3H post XXX challenge
C2926344|T201|COMP|58602-4|LNC|Corticotropin^3rd specimen post XXX challenge|Corticotropin^3rd specimen post XXX challenge
C2926345|T201|COMP|58603-2|LNC|Corticotropin^4 AM specimen|Corticotropin^4 AM specimen
C2926346|T201|COMP|58604-0|LNC|Corticotropin^4 PM specimen|Corticotropin^4 PM specimen
C2926347|T201|COMP|58605-7|LNC|Corticotropin^45M post 1 ug/kg CRH IV|Corticotropin^45M post 1 ug/kg CRH IV
C2926348|T201|COMP|58606-5|LNC|Corticotropin^45M post dose insulin IV|Corticotropin^45M post dose insulin IV
C2926349|T201|COMP|58607-3|LNC|Corticotropin^2D post dose metyraPONE|Corticotropin^2D post dose metyraPONE
C2926350|T201|COMP|58608-1|LNC|Corticotropin^4th specimen post XXX challenge|Corticotropin^4th specimen post XXX challenge
C2926351|T201|COMP|58609-9|LNC|Corticotropin^5th specimen post XXX challenge|Corticotropin^5th specimen post XXX challenge
C2926352|T201|COMP|58610-7|LNC|Corticotropin^6 PM specimen|Corticotropin^6 PM specimen
C2926353|T201|COMP|58611-5|LNC|Corticotropin^6th specimen post XXX challenge|Corticotropin^6th specimen post XXX challenge
C2926354|T201|COMP|58612-3|LNC|Corticotropin^75M post dose insulin IV|Corticotropin^75M post dose insulin IV
C2926355|T201|COMP|58613-1|LNC|Corticotropin^75M post dose insulin IV|Corticotropin^75M post dose insulin IV
C2926356|T201|COMP|58614-9|LNC|Corticotropin^7th specimen post XXX challenge|Corticotropin^7th specimen post XXX challenge
C2926357|T201|COMP|58615-6|LNC|Corticotropin^8 AM specimen|Corticotropin^8 AM specimen
C2926358|T201|COMP|58616-4|LNC|Corticotropin^8 PM specimen|Corticotropin^8 PM specimen
C2926359|T201|COMP|58617-2|LNC|Corticotropin^8th specimen post XXX challenge|Corticotropin^8th specimen post XXX challenge
C2926360|T201|COMP|58618-0|LNC|Corticotropin^post dose dexamethasone|Corticotropin^post dose dexamethasone
C2926361|T201|COMP|58619-8|LNC|Corticotropin^pre 1 ug/kg CRH IV|Corticotropin^pre 1 ug/kg CRH IV
C2926362|T201|COMP|58620-6|LNC|Corticotropin^pre dose dexamethasone|Corticotropin^pre dose dexamethasone
C2926363|T201|COMP|58621-4|LNC|Corticotropin^pre dose dexamethasone|Corticotropin^pre dose dexamethasone
C2926364|T201|COMP|58622-2|LNC|Corticotropin^pre dose glucagon|Corticotropin^pre dose glucagon
C2926365|T201|COMP|58623-0|LNC|Corticotropin^pre dose glucagon|Corticotropin^pre dose glucagon
C2926366|T201|COMP|58624-8|LNC|Corticotropin^pre dose glucose|Corticotropin^pre dose glucose
C2926367|T201|COMP|58625-5|LNC|Corticotropin^pre dose glucose|Corticotropin^pre dose glucose
C2926368|T201|COMP|58626-3|LNC|Corticotropin^pre dose insulin IV|Corticotropin^pre dose insulin IV
C2926369|T201|COMP|58627-1|LNC|Corticotropin^pre dose metyraPONE|Corticotropin^pre dose metyraPONE
C2926370|T201|COMP|58628-9|LNC|Corticotropin^pre dose metyraPONE|Corticotropin^pre dose metyraPONE
C2926371|T201|COMP|58629-7|LNC|Corticotropin^pre XXX challenge|Corticotropin^pre XXX challenge
C2926372|T201|COMP|58630-5|LNC|Corticotropin^pre XXX challenge|Corticotropin^pre XXX challenge
C2926373|T201|COMP|58631-3|LNC|Cortisol^1.5H post 1 ug/kg CRH IV|Cortisol^1.5H post 1 ug/kg CRH IV
C2926374|T201|COMP|58632-1|LNC|Cortisol^1.5H post 1 ug/kg CRH IV|Cortisol^1.5H post 1 ug/kg CRH IV
C2926375|T201|COMP|58633-9|LNC|Cortisol^10 AM specimen|Cortisol^10 AM specimen
C2926376|T201|COMP|58634-7|LNC|Cortisol^10 AM specimen|Cortisol^10 AM specimen
C2926377|T201|COMP|58635-4|LNC|Cortisol^10 PM specimen|Cortisol^10 PM specimen
C2926378|T201|COMP|58636-2|LNC|Cortisol^10 PM specimen|Cortisol^10 PM specimen
C2926379|T201|COMP|58637-0|LNC|Cortisol^10th specimen post XXX challenge|Cortisol^10th specimen post XXX challenge
C2926380|T201|COMP|58638-8|LNC|Cortisol^10th specimen post XXX challenge|Cortisol^10th specimen post XXX challenge
C2926381|T201|COMP|58639-6|LNC|Cortisol^10th specimen post XXX challenge|Cortisol^10th specimen post XXX challenge
C2926382|T201|COMP|58640-4|LNC|Cortisol^11th specimen post XXX challenge|Cortisol^11th specimen post XXX challenge
C2926383|T201|COMP|58641-2|LNC|Cortisol^11th specimen post XXX challenge|Cortisol^11th specimen post XXX challenge
C2926384|T201|COMP|58642-0|LNC|Cortisol^12 AM specimen|Cortisol^12 AM specimen
C2926385|T201|COMP|58643-8|LNC|Cortisol^12 AM specimen|Cortisol^12 AM specimen
C2926386|T201|COMP|58644-6|LNC|Cortisol^12 PM specimen|Cortisol^12 PM specimen
C2926387|T201|COMP|58645-3|LNC|Cortisol^12 PM specimen|Cortisol^12 PM specimen
C2926388|T201|COMP|59142-0|LNC|Cells.CD11c-CD25+/100 cells|Cells.CD11c-CD25+/100 cells
C2926390|T201|COMP|59143-8|LNC|Cells.CD19+CD38+/100 cells|Cells.CD19+CD38+/100 cells
C2926391|T201|COMP|59144-6|LNC|Cells.CD5+CD23+/100 cells|Cells.CD5+CD23+/100 cells
C2926393|T201|COMP|59145-3|LNC|Cells.CD11c+CD103+|Cells.CD11c+CD103+
C2926394|T201|COMP|59146-1|LNC|Cells.CD11c+CD25+|Cells.CD11c+CD25+
C2926395|T201|COMP|59147-9|LNC|Cells.CD19+CD38+|Cells.CD19+CD38+
C2926396|T201|COMP|59148-7|LNC|Calcium^post dialysis|Calcium^post dialysis
C2926397|T201|COMP|59149-5|LNC|Creatine kinase.macromolecular|Creatine kinase.macromolecular
C2926398|T201|COMP|59265-9|LNC|8-Hydroxydeoxyguanosine/Creatinine|8-Hydroxydeoxyguanosine/Creatinine
C2926400|T201|COMP|59266-7|LNC|Maternal cell contamination|Maternal cell contamination
C2926401|T201|COMP|59267-5|LNC|Karyotype|Karyotype
C2926407|T201|COMP|59384-8|LNC|Acetaminophen|Acetaminophen
C2926408|T201|COMP|59387-1|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C2926409|T201|COMP|59388-9|LNC|Taenia solium larva DNA|Taenia solium larva DNA
C2926410|T201|COMP|59389-7|LNC|Androstanolone^1.5H post XXX challenge|Androstanolone^1.5H post XXX challenge
C2926411|T201|COMP|59390-5|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C2926412|T201|COMP|59391-3|LNC|Prunus persica recombinant (rPru p) 3 Ab.IgE|Prunus persica recombinant (rPru p) 3 Ab.IgE
C2926414|T201|COMP|59392-1|LNC|Hydroxyproline|Hydroxyproline
C2926415|T201|COMP|59393-9|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C2926416|T201|COMP|59394-7|LNC|Glomerular basement membrane Ab|Glomerular basement membrane Ab
C2926417|T201|COMP|59395-4|LNC|Latex recombinant (rHev b) 9 Ab.IgE|Latex recombinant (rHev b) 9 Ab.IgE
C2926419|T201|COMP|59396-2|LNC|Echovirus Ab.IgM|Echovirus Ab.IgM
C2926420|T201|COMP|59397-0|LNC|Echovirus Ab.IgG|Echovirus Ab.IgG
C2926421|T201|COMP|59398-8|LNC|Ascorbate|Ascorbate
C2926422|T201|COMP|59399-6|LNC|PM-1 Ab|PM-1 Ab
C2926423|T201|COMP|59652-8|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2926424|T201|COMP|59653-6|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2926425|T201|COMP|59654-4|LNC|diazePAM|diazePAM
C2926426|T201|COMP|59655-1|LNC|diazePAM|diazePAM
C2926427|T201|COMP|59656-9|LNC|diazePAM|diazePAM
C2926428|T201|COMP|59657-7|LNC|diazePAM|diazePAM
C2926429|T201|COMP|59658-5|LNC|diazePAM|diazePAM
C2926430|T201|COMP|58646-1|LNC|Cortisol^12th specimen post XXX challenge|Cortisol^12th specimen post XXX challenge
C2926431|T201|COMP|58647-9|LNC|Cortisol^12th specimen post XXX challenge|Cortisol^12th specimen post XXX challenge
C2926432|T201|COMP|58648-7|LNC|Cortisol^15M post 1 ug/kg CRH IV|Cortisol^15M post 1 ug/kg CRH IV
C2926433|T201|COMP|58649-5|LNC|Cortisol^15M post 1 ug/kg CRH IV|Cortisol^15M post 1 ug/kg CRH IV
C2926434|T201|COMP|58650-3|LNC|Cortisol^15M pre 1 ug/kg CRH IV|Cortisol^15M pre 1 ug/kg CRH IV
C2926435|T201|COMP|58651-1|LNC|Cortisol^15M pre 1 ug/kg CRH IV|Cortisol^15M pre 1 ug/kg CRH IV
C2926436|T201|COMP|58652-9|LNC|Cortisol^1H post 1 ug/kg CRH IV|Cortisol^1H post 1 ug/kg CRH IV
C2926437|T201|COMP|58653-7|LNC|Cortisol^1H post 1 ug/kg CRH IV|Cortisol^1H post 1 ug/kg CRH IV
C2926438|T201|COMP|58654-5|LNC|Cortisol^1st specimen post XXX challenge|Cortisol^1st specimen post XXX challenge
C2926439|T201|COMP|58655-2|LNC|Cortisol^2 PM specimen|Cortisol^2 PM specimen
C2926440|T201|COMP|58656-0|LNC|Cortisol^2 PM specimen|Cortisol^2 PM specimen
C2926441|T201|COMP|58657-8|LNC|Cortisol^2H post 1 ug/kg CRH IV|Cortisol^2H post 1 ug/kg CRH IV
C2926442|T201|COMP|58658-6|LNC|Cortisol^2H post 1 ug/kg CRH IV|Cortisol^2H post 1 ug/kg CRH IV
C2926443|T201|COMP|58659-4|LNC|Cortisol^2H post 1 ug/kg CRH IV|Cortisol^2H post 1 ug/kg CRH IV
C2926444|T201|COMP|58660-2|LNC|Cortisol^2nd specimen post XXX challenge|Cortisol^2nd specimen post XXX challenge
C2926445|T201|COMP|58661-0|LNC|Cortisol^30M pre 1 ug/kg CRH IV|Cortisol^30M pre 1 ug/kg CRH IV
C2926446|T201|COMP|58662-8|LNC|Cortisol^30M pre 1 ug/kg CRH IV|Cortisol^30M pre 1 ug/kg CRH IV
C2926447|T201|COMP|58663-6|LNC|Cortisol^30M pre 1 ug/kg CRH IV|Cortisol^30M pre 1 ug/kg CRH IV
C2926448|T201|COMP|58664-4|LNC|Cortisol^30M pre 1 ug/kg CRH IV|Cortisol^30M pre 1 ug/kg CRH IV
C2926449|T201|COMP|58665-1|LNC|Cortisol^3rd specimen post XXX challenge|Cortisol^3rd specimen post XXX challenge
C2926450|T201|COMP|58666-9|LNC|Cortisol^4 AM specimen|Cortisol^4 AM specimen
C2926451|T201|COMP|58667-7|LNC|Cortisol^4 AM specimen|Cortisol^4 AM specimen
C2926452|T201|COMP|58668-5|LNC|Cortisol^4 PM specimen|Cortisol^4 PM specimen
C2926453|T201|COMP|58669-3|LNC|Cortisol^4 PM specimen|Cortisol^4 PM specimen
C2926454|T201|COMP|58670-1|LNC|Cortisol^45M post 1 ug/kg CRH IV|Cortisol^45M post 1 ug/kg CRH IV
C2926455|T201|COMP|58671-9|LNC|Cortisol^45M post 1 ug/kg CRH IV|Cortisol^45M post 1 ug/kg CRH IV
C2926456|T201|COMP|58672-7|LNC|Cortisol^45M post 1 ug/kg CRH IV|Cortisol^45M post 1 ug/kg CRH IV
C2926457|T201|COMP|58673-5|LNC|Cortisol^4th specimen post XXX challenge|Cortisol^4th specimen post XXX challenge
C2926458|T201|COMP|58674-3|LNC|Cortisol^8 AM specimen|Cortisol^8 AM specimen
C2926459|T201|COMP|58675-0|LNC|Cortisol^8 AM specimen|Cortisol^8 AM specimen
C2926460|T201|COMP|58676-8|LNC|Cortisol^8 PM specimen|Cortisol^8 PM specimen
C2926461|T201|COMP|58677-6|LNC|Cortisol^8 PM specimen|Cortisol^8 PM specimen
C2926462|T201|COMP|58678-4|LNC|Cortisol^pre 1 ug/kg CRH IV|Cortisol^pre 1 ug/kg CRH IV
C2926463|T201|COMP|58679-2|LNC|Cortisol^pre 1 ug/kg CRH IV|Cortisol^pre 1 ug/kg CRH IV
C2926465|T201|COMP|58681-8|LNC|Temperature|Temperature
C2926466|T201|COMP|58682-6|LNC|Sulfatides|Sulfatides
C2926467|T201|COMP|58683-4|LNC|Complement C5|Complement C5
C2926468|T201|COMP|58684-2|LNC|Uroporphyrin 1 isomer/Creatinine|Uroporphyrin 1 isomer/Creatinine
C2926470|T201|COMP|58705-5|LNC|cefTAZidime|cefTAZidime
C2926471|T201|COMP|58706-3|LNC|OmpC Ab.IgA|OmpC Ab.IgA
C2926472|T201|COMP|58707-1|LNC|Ephedrine+Pseudoephedrine|Ephedrine+Pseudoephedrine
C2926473|T201|COMP|58708-9|LNC|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C2926474|T201|COMP|58709-7|LNC|Gliadin peptide Ab.IgA|Gliadin peptide Ab.IgA
C2926475|T201|COMP|58710-5|LNC|Gliadin peptide Ab.IgG|Gliadin peptide Ab.IgG
C2926476|T201|COMP|58711-3|LNC|Doripenem|Doripenem
C2926477|T201|COMP|58712-1|LNC|Quinupristin+Dalfopristin|Quinupristin+Dalfopristin
C2926479|T201|COMP|58714-7|LNC|Oxidants|Oxidants
C2926480|T201|COMP|58715-4|LNC|Adulterants panel|Adulterants panel
C2926481|T201|COMP|58716-2|LNC|Testosterone.free+weakly bound & total panel|Testosterone.free+weakly bound & total panel
C2926600|T201|COMP|58357-5|LNC|Amphetamine/Creatinine|Amphetamine/Creatinine
C2926608|T201|COMP|59020-8|LNC|HLA-DRB5|HLA-DRB5
C2926609|T201|COMP|59021-6|LNC|HLA-DRB4|HLA-DRB4
C2926620|T201|COMP|59177-6|LNC|Beta-2-Microglobulin/Creatinine|Beta-2-Microglobulin/Creatinine
C2926622|T201|COMP|40611-6|LNC|Blasts|Blasts
C2966435|T201|COMP|57906-0|LNC|9p21 chromosome deletion|9p21 chromosome deletion
C2966439|T201|COMP|59023-2|LNC|Adenosine deaminase|Adenosine deaminase
C2966440|T201|COMP|59386-3|LNC|Starch|Starch
C2966441|T201|COMP|58353-4|LNC|Human antihuman Ab|Human antihuman Ab
C2966442|T201|COMP|58354-2|LNC|Human antihuman Ab|Human antihuman Ab
C2966443|T201|COMP|59385-5|LNC|Nitrogen|Nitrogen
C2966611|T201|COMP|60437-1|LNC|Cells.CD5+CD23+|Cells.CD5+CD23+
C2966612|T201|COMP|60438-9|LNC|Diamine oxidase|Diamine oxidase
C2966613|T201|COMP|60439-7|LNC|Lymphocytes.large granular/100 leukocytes|Lymphocytes.large granular/100 leukocytes
C2966614|T201|COMP|60440-5|LNC|Oseltamivir|Oseltamivir
C2966615|T201|COMP|60441-3|LNC|Oseltamivir+Zanamivir|Oseltamivir+Zanamivir
C2966616|T201|COMP|60442-1|LNC|HEDIS 2011 panel|HEDIS 2011 panel
C2966618|T201|COMP|58766-7|LNC|Epithelial cells|Epithelial cells
C2966619|T201|COMP|58767-5|LNC|Erythrocytes|Erythrocytes
C2966620|T201|COMP|59015-8|LNC|Carbohydrates|Carbohydrates
C2966621|T201|COMP|59016-6|LNC|Water|Water
C2966631|T201|COMP|59957-1|LNC|Promazine|Promazine
C2966632|T201|COMP|59958-9|LNC|Promazine|Promazine
C2966633|T201|COMP|59959-7|LNC|Promazine|Promazine
C2966634|T201|COMP|59960-5|LNC|Propoxyphene|Propoxyphene
C2966635|T201|COMP|59961-3|LNC|Propoxyphene|Propoxyphene
C2966636|T201|COMP|59962-1|LNC|Propranolol|Propranolol
C2966637|T201|COMP|59963-9|LNC|QUEtiapine|QUEtiapine
C2966638|T201|COMP|59964-7|LNC|QUEtiapine|QUEtiapine
C2966639|T201|COMP|59965-4|LNC|quiNINE|quiNINE
C2966640|T201|COMP|59966-2|LNC|quiNINE|quiNINE
C2966641|T201|COMP|59967-0|LNC|quiNINE|quiNINE
C2966642|T201|COMP|60201-1|LNC|Salicylates|Salicylates
C2966643|T201|COMP|60204-5|LNC|Trimethadione|Trimethadione
C2966644|T201|COMP|60205-2|LNC|Trimethadione|Trimethadione
C2966645|T201|COMP|60206-0|LNC|Tripelennamine|Tripelennamine
C2966646|T201|COMP|60207-8|LNC|Vanadium|Vanadium
C2966647|T201|COMP|60208-6|LNC|Venlafaxine|Venlafaxine
C2966648|T201|COMP|60209-4|LNC|Venlafaxine|Venlafaxine
C2966649|T201|COMP|60210-2|LNC|Venlafaxine|Venlafaxine
C2966650|T201|COMP|60211-0|LNC|Zolazepam|Zolazepam
C2966651|T201|COMP|60376-1|LNC|Vitis vinifera Ab.IgG|Vitis vinifera Ab.IgG
C2966652|T201|COMP|60377-9|LNC|Citrus paradisis Ab.IgG|Citrus paradisis Ab.IgG
C2966653|T201|COMP|60378-7|LNC|Melanogrammus aeglefinus Ab.IgG|Melanogrammus aeglefinus Ab.IgG
C2966654|T201|COMP|60379-5|LNC|Hippoglossus hippoglossus Ab.IgG|Hippoglossus hippoglossus Ab.IgG
C2966655|T201|COMP|60380-3|LNC|Lamb Ab.IgG|Lamb Ab.IgG
C2966656|T201|COMP|60381-1|LNC|Citrus limon Ab.IgG|Citrus limon Ab.IgG
C2966657|T201|COMP|60382-9|LNC|Citrus aurantifolia Ab.IgG|Citrus aurantifolia Ab.IgG
C2966658|T201|COMP|60383-7|LNC|Homarus gammarus Ab.IgG|Homarus gammarus Ab.IgG
C2966659|T201|COMP|60384-5|LNC|Mustard Ab.IgG|Mustard Ab.IgG
C2966660|T201|COMP|60385-2|LNC|Nutmeg Ab.IgG|Nutmeg Ab.IgG
C2966661|T201|COMP|60386-0|LNC|Olive green Ab.IgG|Olive green Ab.IgG
C2966662|T201|COMP|60387-8|LNC|Origanum vulgare Ab.IgG|Origanum vulgare Ab.IgG
C2966663|T201|COMP|60388-6|LNC|Ostrea edulis Ab.IgG|Ostrea edulis Ab.IgG
C2966664|T201|COMP|60389-4|LNC|Pisum sativum Ab.IgG|Pisum sativum Ab.IgG
C2966665|T201|COMP|60390-2|LNC|Prunus persica Ab.IgG|Prunus persica Ab.IgG
C2966666|T201|COMP|60391-0|LNC|Pyrus communis Ab.IgG|Pyrus communis Ab.IgG
C2966667|T201|COMP|60392-8|LNC|Piper nigrum Ab.IgG|Piper nigrum Ab.IgG
C2966668|T201|COMP|60393-6|LNC|Pepper green Ab.IgG|Pepper green Ab.IgG
C2966669|T201|COMP|60394-4|LNC|Ananas comosus Ab.IgG|Ananas comosus Ab.IgG
C2966672|T201|COMP|60517-0|LNC|Iron/Transferrin|Iron/Transferrin
C2966673|T201|COMP|60518-8|LNC|Creatinine|Creatinine
C2966674|T201|COMP|60520-4|LNC|Eosinophils|Eosinophils
C2966675|T201|COMP|60521-2|LNC|Babesia microti Ab.IgG+IgM|Babesia microti Ab.IgG+IgM
C2966677|T201|COMP|60522-0|LNC|Borrelia hermsii Ab.IgG+IgM|Borrelia hermsii Ab.IgG+IgM
C2966679|T201|COMP|60523-8|LNC|Carbromal|Carbromal
C2966680|T201|COMP|60524-6|LNC|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C2966682|T201|COMP|59273-3|LNC|Cortisol^post 6 mg dexamethasone PO overnight|Cortisol^post 6 mg dexamethasone PO overnight
C2966683|T201|COMP|59470-5|LNC|Calcium.ionized|Calcium.ionized
C2966684|T201|COMP|59471-3|LNC|Calcium.ionized|Calcium.ionized
C2966685|T201|COMP|59472-1|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C2966686|T201|COMP|59473-9|LNC|Calcium.ionized^^adjusted to pH 7.4|Calcium.ionized^^adjusted to pH 7.4
C2966756|T201|COMP|60341-5|LNC|Sodium urate crystals|Sodium urate crystals
C2966757|T201|COMP|60342-3|LNC|Borrelia burgdorferi Ab.IgG panel|Borrelia burgdorferi Ab.IgG panel
C2966758|T201|COMP|60343-1|LNC|Borrelia burgdorferi Ab.IgM panel|Borrelia burgdorferi Ab.IgM panel
C2966759|T201|COMP|60344-9|LNC|Lipoprotein (little a)/Lipoprotein.total|Lipoprotein (little a)/Lipoprotein.total
C2966761|T201|COMP|60345-6|LNC|Viable CD34 cells/100 cells|Viable CD34 cells/100 cells
C2966763|T201|COMP|60346-4|LNC|Viable CD34 cells/100 cells.CD34|Viable CD34 cells/100 cells.CD34
C2966765|T201|COMP|60347-2|LNC|Viable CD34 cells|Viable CD34 cells
C2966766|T201|COMP|60459-5|LNC|Complement C6.functional|Complement C6.functional
C2966767|T201|COMP|60461-1|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C2966768|T201|COMP|60462-9|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C2966769|T201|COMP|60463-7|LNC|Insulin Ab|Insulin Ab
C2966770|T201|COMP|60464-5|LNC|Monosodium glutamate Ab.IgE.RAST class|Monosodium glutamate Ab.IgE.RAST class
C2966772|T201|COMP|61101-2|LNC|Influenza virus A neuraminidase RNA|Influenza virus A neuraminidase RNA
C2966773|T201|COMP|61102-0|LNC|Influenza virus A & B Ag|Influenza virus A & B Ag
C2966774|T201|COMP|61103-8|LNC|Prochlorperazine|Prochlorperazine
C2966775|T201|COMP|61104-6|LNC|Prochlorperazine|Prochlorperazine
C2966776|T201|COMP|61105-3|LNC|Prochlorperazine|Prochlorperazine
C2966777|T201|COMP|61106-1|LNC|16p11.2 chromosome region deletion+duplication|16p11.2 chromosome region deletion+duplication
C2966778|T201|COMP|61107-9|LNC|SLC25A13 gene targeted mutation analysis|SLC25A13 gene targeted mutation analysis
C2966782|T201|COMP|61256-4|LNC|Dactylis glomerata Ab.IgE/IgE.total|Dactylis glomerata Ab.IgE/IgE.total
C2966783|T201|COMP|61257-2|LNC|Dermatophagoides microceras Ab.IgE/IgE.total|Dermatophagoides microceras Ab.IgE/IgE.total
C2966784|T201|COMP|61258-0|LNC|Dermatophagoides pteronyssinus Ab.IgE/IgE.total|Dermatophagoides pteronyssinus Ab.IgE/IgE.total
C2966785|T201|COMP|61259-8|LNC|Dolichovespula maculata Ab.IgE/IgE.total|Dolichovespula maculata Ab.IgE/IgE.total
C2966786|T201|COMP|61260-6|LNC|Erythromycin Ab.IgE/IgE.total|Erythromycin Ab.IgE/IgE.total
C2966787|T201|COMP|61261-4|LNC|Eucalyptus spp Ab.IgE/IgE.total|Eucalyptus spp Ab.IgE/IgE.total
C2966788|T201|COMP|61262-2|LNC|Fagopyrum esculentum Ab.IgE/IgE.total|Fagopyrum esculentum Ab.IgE/IgE.total
C2966789|T201|COMP|61263-0|LNC|Fagus grandifolia Ab.IgE/IgE.total|Fagus grandifolia Ab.IgE/IgE.total
C2966790|T201|COMP|61264-8|LNC|Festuca elatior Ab.IgE/IgE.total|Festuca elatior Ab.IgE/IgE.total
C2966791|T201|COMP|61265-5|LNC|Foeniculum vulgare seed Ab.IgE/IgE.total|Foeniculum vulgare seed Ab.IgE/IgE.total
C2966792|T201|COMP|61266-3|LNC|Fragaria vesca Ab.IgE/IgE.total|Fragaria vesca Ab.IgE/IgE.total
C2966793|T201|COMP|61267-1|LNC|Franseria acanthicarpa Ab.IgE/IgE.total|Franseria acanthicarpa Ab.IgE/IgE.total
C2966794|T201|COMP|61268-9|LNC|Gadus morhua Ab.IgG/IgE.total|Gadus morhua Ab.IgG/IgE.total
C2966795|T201|COMP|61269-7|LNC|Gelatin Ab.IgE/IgE.total|Gelatin Ab.IgE/IgE.total
C2966796|T201|COMP|61393-5|LNC|Human papilloma virus 6 DNA|Human papilloma virus 6 DNA
C2966797|T201|COMP|61394-3|LNC|Human papilloma virus 11 DNA|Human papilloma virus 11 DNA
C2966798|T201|COMP|61395-0|LNC|Human papilloma virus 42 DNA|Human papilloma virus 42 DNA
C2966799|T201|COMP|61396-8|LNC|Human papilloma virus 56 DNA|Human papilloma virus 56 DNA
C2966800|T201|COMP|61397-6|LNC|Enterococcus faecium DNA|Enterococcus faecium DNA
C2966801|T201|COMP|61398-4|LNC|Escherichia coli DNA|Escherichia coli DNA
C2966802|T201|COMP|61399-2|LNC|Klebsiella pneumoniae DNA|Klebsiella pneumoniae DNA
C2966803|T201|COMP|62360-3|LNC|Cells analyzed|Cells analyzed
C2966804|T201|COMP|62361-1|LNC|Cells counted|Cells counted
C2966805|T201|COMP|62362-9|LNC|Colonies counted|Colonies counted
C2966806|T201|COMP|62363-7|LNC|Mosaicism detected|Mosaicism detected
C2966807|T201|COMP|62364-5|LNC|Test performance information|Test performance information
C2966808|T201|COMP|62365-2|LNC|Diagnostic impression|Diagnostic impression
C2966809|T201|COMP|62366-0|LNC|Recommended follow-up|Recommended follow-up
C2966810|T201|COMP|59697-3|LNC|Iodide|Iodide
C2966813|T201|COMP|60013-0|LNC|Cortisol^40M post XXX challenge|Cortisol^40M post XXX challenge
C2966814|T201|COMP|60014-8|LNC|Corticotropin^baseline|Corticotropin^baseline
C2966815|T201|COMP|60015-5|LNC|Corticotropin^5M post XXX challenge|Corticotropin^5M post XXX challenge
C2966816|T201|COMP|60016-3|LNC|Corticotropin^1.5H post XXX challenge|Corticotropin^1.5H post XXX challenge
C2966817|T201|COMP|60172-4|LNC|Strontium|Strontium
C2966818|T201|COMP|60173-2|LNC|Strontium|Strontium
C2966819|T201|COMP|60174-0|LNC|Strontium|Strontium
C2966820|T201|COMP|60175-7|LNC|Sulfamethizole|Sulfamethizole
C2966821|T201|COMP|60176-5|LNC|Sulfamethizole|Sulfamethizole
C2966822|T201|COMP|60177-3|LNC|Sulfamethizole|Sulfamethizole
C2966823|T201|COMP|60178-1|LNC|Tellurium|Tellurium
C2966824|T201|COMP|60179-9|LNC|Tellurium|Tellurium
C2966825|T201|COMP|60180-7|LNC|Tellurium|Tellurium
C2966826|T201|COMP|60181-5|LNC|Tellurium|Tellurium
C2966827|T201|COMP|60182-3|LNC|Temephos|Temephos
C2966828|T201|COMP|60183-1|LNC|Terazosin|Terazosin
C2966829|T201|COMP|60184-9|LNC|Terazosin|Terazosin
C2966830|T201|COMP|60185-6|LNC|Thallium|Thallium
C2966831|T201|COMP|60186-4|LNC|Thiethylperazine|Thiethylperazine
C2966832|T201|COMP|60187-2|LNC|Thiethylperazine|Thiethylperazine
C2966833|T201|COMP|60188-0|LNC|Thiethylperazine|Thiethylperazine
C2966834|T201|COMP|60189-8|LNC|Tin|Tin
C2966835|T201|COMP|60190-6|LNC|Tin|Tin
C2966836|T201|COMP|60191-4|LNC|Tin|Tin
C2966837|T201|COMP|60192-2|LNC|Topiramate|Topiramate
C2966838|T201|COMP|60193-0|LNC|Topiramate|Topiramate
C2966839|T201|COMP|60435-5|LNC|Cells.CD10+CD19+|Cells.CD10+CD19+
C2966840|T201|COMP|60436-3|LNC|Cells.CD19+CD25+|Cells.CD19+CD25+
C2966842|T201|COMP|60445-4|LNC|HEDIS 2011 Codes to identify exclusions (CHL-D)|HEDIS 2011 Codes to identify exclusions (CHL-D)
C2966848|T201|COMP|60080-9|LNC|Germanium|Germanium
C2966849|T201|COMP|60081-7|LNC|Germanium|Germanium
C2966850|T201|COMP|60082-5|LNC|Gold|Gold
C2966851|T201|COMP|60083-3|LNC|Hydroxybupropion|Hydroxybupropion
C2966852|T201|COMP|60084-1|LNC|Hydroxybupropion|Hydroxybupropion
C2966853|T201|COMP|60085-8|LNC|Hydroxybupropion|Hydroxybupropion
C2966854|T201|COMP|60086-6|LNC|Hydroxybupropion|Hydroxybupropion
C2966855|T201|COMP|60087-4|LNC|Hyoscyamine|Hyoscyamine
C2966856|T201|COMP|60088-2|LNC|Hyoscyamine|Hyoscyamine
C2966857|T201|COMP|60089-0|LNC|Indium|Indium
C2966858|T201|COMP|60309-2|LNC|Imipramine|Imipramine
C2966859|T201|COMP|60310-0|LNC|Indomethacin|Indomethacin
C2966860|T201|COMP|60311-8|LNC|Ketoprofen|Ketoprofen
C2966861|T201|COMP|60312-6|LNC|lamoTRIgine|lamoTRIgine
C2966862|T201|COMP|60313-4|LNC|Maprotiline|Maprotiline
C2966863|T201|COMP|60314-2|LNC|Mefenamate|Mefenamate
C2966864|T201|COMP|60315-9|LNC|Mesoridazine|Mesoridazine
C2966865|T201|COMP|60316-7|LNC|Methaqualone|Methaqualone
C2966866|T201|COMP|60317-5|LNC|Methotrimeprazine|Methotrimeprazine
C2966867|T201|COMP|60318-3|LNC|Mexiletine|Mexiletine
C2966868|T201|COMP|60476-9|LNC|Stage|Stage
C2966877|T201|COMP|60485-0|LNC|Interferon.gamma|Interferon.gamma
C2966891|T201|COMP|62203-5|LNC|t(10;11)(p12;q23)(MLLT10,MLL) fusion transcript|t(10;11)(p12;q23)(MLLT10,MLL) fusion transcript
C2969742|T201|COMP|59810-2|LNC|Caffeine^trough|Caffeine^trough
C2969743|T201|COMP|59811-0|LNC|Caffeine^peak|Caffeine^peak
C2969745|T201|COMP|59846-6|LNC|Salmonella sp identified|Salmonella sp identified
C2969748|T201|COMP|59849-0|LNC|Lactate^post exercise|Lactate^post exercise
C2969749|T201|COMP|59850-8|LNC|Wuchereria bancrofti Ag|Wuchereria bancrofti Ag
C2969762|T201|COMP|59864-9|LNC|Acetone|Acetone
C2969763|T201|COMP|59865-6|LNC|Amobarbital|Amobarbital
C2969764|T201|COMP|59866-4|LNC|Amobarbital|Amobarbital
C2969765|T201|COMP|60020-5|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2969766|T201|COMP|60021-3|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2969767|T201|COMP|60022-1|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2969768|T201|COMP|60023-9|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2969769|T201|COMP|60024-7|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2969770|T201|COMP|60025-4|LNC|Urobilinogen|Urobilinogen
C2969771|T201|COMP|60026-2|LNC|Leukocyte esterase|Leukocyte esterase
C2969772|T201|COMP|60027-0|LNC|Specific gravity|Specific gravity
C2969773|T201|COMP|60028-8|LNC|West Nile Virus Ab.IgG avidity|West Nile Virus Ab.IgG avidity
C2969774|T201|COMP|60029-6|LNC|West Nile Virus Ab.IgG avidity|West Nile Virus Ab.IgG avidity
C2969775|T201|COMP|60030-4|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C2969776|T201|COMP|60032-0|LNC|Bacteria identified|Bacteria identified
C2969777|T201|COMP|60033-8|LNC|PIK3CA gene targeted mutation analysis|PIK3CA gene targeted mutation analysis
C2969779|T201|COMP|60034-6|LNC|PIK3CA gene targeted mutation analysis|PIK3CA gene targeted mutation analysis
C2969780|T201|COMP|60035-3|LNC|10-Hydroxycarbazepine|10-Hydroxycarbazepine
C2969781|T201|COMP|60214-4|LNC|ZOLMitriptan|ZOLMitriptan
C2969782|T201|COMP|60215-1|LNC|ZOLMitriptan|ZOLMitriptan
C2969783|T201|COMP|60216-9|LNC|Zomepirac|Zomepirac
C2969784|T201|COMP|60217-7|LNC|Chloride|Chloride
C2969785|T201|COMP|60218-5|LNC|Potassium|Potassium
C2969786|T201|COMP|60219-3|LNC|Ubiquinone 10/Protein|Ubiquinone 10/Protein
C2969788|T201|COMP|60220-1|LNC|Sodium|Sodium
C2969789|T201|COMP|60221-9|LNC|Intrinsic factor Ab.IgG|Intrinsic factor Ab.IgG
C2969790|T201|COMP|60224-3|LNC|Beta-trace protein|Beta-trace protein
C2969791|T201|COMP|60225-0|LNC|Hydrogen/Expired gas^3H post dose fructose PO|Hydrogen/Expired gas^3H post dose fructose PO
C2969792|T201|COMP|60226-8|LNC|Hydrogen/Expired gas^2.5H post dose fructose PO|Hydrogen/Expired gas^2.5H post dose fructose PO
C2969793|T201|COMP|60227-6|LNC|Hydrogen/Expired gas^2H post dose fructose PO|Hydrogen/Expired gas^2H post dose fructose PO
C2969794|T201|COMP|60228-4|LNC|Hydrogen/Expired gas^1.5H post dose fructose PO|Hydrogen/Expired gas^1.5H post dose fructose PO
C2969795|T201|COMP|60229-2|LNC|Hydrogen/Expired gas^1H post dose fructose PO|Hydrogen/Expired gas^1H post dose fructose PO
C2969796|T201|COMP|60230-0|LNC|Hydrogen/Expired gas^30M post dose fructose PO|Hydrogen/Expired gas^30M post dose fructose PO
C2969797|T201|COMP|60231-8|LNC|Hydrogen/Expired gas^pre dose fructose PO|Hydrogen/Expired gas^pre dose fructose PO
C2969798|T201|COMP|60232-6|LNC|Hydrogen/Expired gas^2.75H post dose lactose PO|Hydrogen/Expired gas^2.75H post dose lactose PO
C2969799|T201|COMP|60233-4|LNC|Hydrogen/Expired gas^2.25H post dose lactose PO|Hydrogen/Expired gas^2.25H post dose lactose PO
C2969800|T201|COMP|60234-2|LNC|Hydrogen/Expired gas^1.75H post dose lactose PO|Hydrogen/Expired gas^1.75H post dose lactose PO
C2969801|T201|COMP|59867-2|LNC|Amoxapine|Amoxapine
C2969802|T201|COMP|59868-0|LNC|Amoxapine|Amoxapine
C2969803|T201|COMP|59869-8|LNC|Benztropine|Benztropine
C2969804|T201|COMP|59870-6|LNC|Benztropine|Benztropine
C2969805|T201|COMP|59871-4|LNC|Benztropine|Benztropine
C2969806|T201|COMP|59872-2|LNC|Bromazepam|Bromazepam
C2969807|T201|COMP|59873-0|LNC|Bromazepam|Bromazepam
C2969808|T201|COMP|59874-8|LNC|Brompheniramine|Brompheniramine
C2969809|T201|COMP|59875-5|LNC|Brompheniramine|Brompheniramine
C2969810|T201|COMP|59876-3|LNC|carBAMazepine|carBAMazepine
C2969811|T201|COMP|59877-1|LNC|Chloral hydrate|Chloral hydrate
C2969812|T201|COMP|59878-9|LNC|Chloral hydrate|Chloral hydrate
C2969813|T201|COMP|59879-7|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2969814|T201|COMP|59880-5|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2969815|T201|COMP|59881-3|LNC|Chlorpheniramine|Chlorpheniramine
C2969816|T201|COMP|59882-1|LNC|Chlorpheniramine|Chlorpheniramine
C2969817|T201|COMP|59883-9|LNC|Chlorpheniramine|Chlorpheniramine
C2969818|T201|COMP|59884-7|LNC|chlorproMAZINE|chlorproMAZINE
C2969819|T201|COMP|59885-4|LNC|chlorproMAZINE|chlorproMAZINE
C2969820|T201|COMP|59886-2|LNC|Citalopram|Citalopram
C2969821|T201|COMP|59887-0|LNC|Citalopram|Citalopram
C2969822|T201|COMP|59888-8|LNC|cloBAZam|cloBAZam
C2969823|T201|COMP|59889-6|LNC|clomiPRAMINE|clomiPRAMINE
C2969824|T201|COMP|59890-4|LNC|cloZAPine|cloZAPine
C2969825|T201|COMP|59891-2|LNC|Cotinine|Cotinine
C2969826|T201|COMP|59892-0|LNC|Cotinine|Cotinine
C2969827|T201|COMP|59893-8|LNC|Desipramine|Desipramine
C2969828|T201|COMP|59894-6|LNC|Dextromethorphan|Dextromethorphan
C2969829|T201|COMP|59895-3|LNC|Dextromethorphan|Dextromethorphan
C2969830|T201|COMP|59896-1|LNC|Dextromethorphan|Dextromethorphan
C2969831|T201|COMP|59897-9|LNC|Disopyramide|Disopyramide
C2969832|T201|COMP|59898-7|LNC|Disopyramide|Disopyramide
C2969833|T201|COMP|59899-5|LNC|Ethylene glycol|Ethylene glycol
C2969834|T201|COMP|59900-1|LNC|Fenoprofen|Fenoprofen
C2969835|T201|COMP|59901-9|LNC|Fenoprofen|Fenoprofen
C2969836|T201|COMP|59902-7|LNC|FLUoxetine|FLUoxetine
C2969837|T201|COMP|59903-5|LNC|FLUoxetine|FLUoxetine
C2969838|T201|COMP|59904-3|LNC|fluPHENAZine|fluPHENAZine
C2969839|T201|COMP|59905-0|LNC|fluPHENAZine|fluPHENAZine
C2969840|T201|COMP|59906-8|LNC|fluvoxaMINE|fluvoxaMINE
C2969841|T201|COMP|59907-6|LNC|fluvoxaMINE|fluvoxaMINE
C2969842|T201|COMP|59908-4|LNC|hydrOXYzine|hydrOXYzine
C2969843|T201|COMP|59909-2|LNC|hydrOXYzine|hydrOXYzine
C2969844|T201|COMP|59910-0|LNC|Ibuprofen|Ibuprofen
C2969845|T201|COMP|59911-8|LNC|Ibuprofen|Ibuprofen
C2969846|T201|COMP|59912-6|LNC|Imipramine|Imipramine
C2969847|T201|COMP|59913-4|LNC|Imipramine|Imipramine
C2969848|T201|COMP|59914-2|LNC|Indomethacin|Indomethacin
C2969849|T201|COMP|59915-9|LNC|Indomethacin|Indomethacin
C2969850|T201|COMP|59916-7|LNC|Isopropanol|Isopropanol
C2969851|T201|COMP|59917-5|LNC|Ketoprofen|Ketoprofen
C2969852|T201|COMP|59918-3|LNC|Ketoprofen|Ketoprofen
C2969853|T201|COMP|59919-1|LNC|lamoTRIgine|lamoTRIgine
C2969854|T201|COMP|59920-9|LNC|lamoTRIgine|lamoTRIgine
C2969855|T201|COMP|59921-7|LNC|Mefenamate|Mefenamate
C2969856|T201|COMP|59922-5|LNC|Mefenamate|Mefenamate
C2969857|T201|COMP|59923-3|LNC|Mefenamate|Mefenamate
C2969858|T201|COMP|59924-1|LNC|Meperidine|Meperidine
C2969859|T201|COMP|59925-8|LNC|Mesoridazine|Mesoridazine
C2969860|T201|COMP|59926-6|LNC|Mesoridazine|Mesoridazine
C2969861|T201|COMP|59927-4|LNC|Methanol|Methanol
C2969862|T201|COMP|59928-2|LNC|Methaqualone|Methaqualone
C2969863|T201|COMP|59929-0|LNC|Methaqualone|Methaqualone
C2969864|T201|COMP|59930-8|LNC|Methotrimeprazine|Methotrimeprazine
C2969865|T201|COMP|59931-6|LNC|Methotrimeprazine|Methotrimeprazine
C2969866|T201|COMP|59932-4|LNC|Mexiletine|Mexiletine
C2969867|T201|COMP|59933-2|LNC|Mexiletine|Mexiletine
C2969868|T201|COMP|59934-0|LNC|Naproxen|Naproxen
C2969869|T201|COMP|59935-7|LNC|Naproxen|Naproxen
C2969870|T201|COMP|59936-5|LNC|Nicotine|Nicotine
C2969871|T201|COMP|59937-3|LNC|Nicotine|Nicotine
C2969872|T201|COMP|59938-1|LNC|Norclobazam|Norclobazam
C2969873|T201|COMP|59939-9|LNC|Norclobazam|Norclobazam
C2969874|T201|COMP|59940-7|LNC|Norclomipramine|Norclomipramine
C2969875|T201|COMP|59941-5|LNC|Norclomipramine|Norclomipramine
C2969876|T201|COMP|59942-3|LNC|Nordoxepin|Nordoxepin
C2969877|T201|COMP|59943-1|LNC|Nordoxepin|Nordoxepin
C2969878|T201|COMP|59944-9|LNC|Normeperidine|Normeperidine
C2969879|T201|COMP|59945-6|LNC|Nortriptyline|Nortriptyline
C2969880|T201|COMP|59946-4|LNC|OLANZapine|OLANZapine
C2969881|T201|COMP|59947-2|LNC|OXcarbazepine|OXcarbazepine
C2969882|T201|COMP|59948-0|LNC|OXcarbazepine|OXcarbazepine
C2969883|T201|COMP|59949-8|LNC|PARoxetine|PARoxetine
C2969884|T201|COMP|59950-6|LNC|PARoxetine|PARoxetine
C2969885|T201|COMP|59951-4|LNC|Pentazocine|Pentazocine
C2969886|T201|COMP|59952-2|LNC|Pentazocine|Pentazocine
C2969887|T201|COMP|59953-0|LNC|Perphenazine|Perphenazine
C2969888|T201|COMP|59954-8|LNC|Perphenazine|Perphenazine
C2969889|T201|COMP|59955-5|LNC|Perphenazine|Perphenazine
C2969890|T201|COMP|59956-3|LNC|Phencyclidine|Phencyclidine
C2969891|T201|COMP|59968-8|LNC|Strychnine|Strychnine
C2969892|T201|COMP|59969-6|LNC|Strychnine|Strychnine
C2969893|T201|COMP|59970-4|LNC|Strychnine|Strychnine
C2969894|T201|COMP|59971-2|LNC|Sulfamethoxazole|Sulfamethoxazole
C2969895|T201|COMP|59972-0|LNC|Sulfamethoxazole|Sulfamethoxazole
C2969896|T201|COMP|59973-8|LNC|Thiocyanate|Thiocyanate
C2969897|T201|COMP|59974-6|LNC|Thiocyanate|Thiocyanate
C2969898|T201|COMP|59975-3|LNC|traZODone|traZODone
C2969899|T201|COMP|59976-1|LNC|traZODone|traZODone
C2969900|T201|COMP|59977-9|LNC|Venlafaxine|Venlafaxine
C2969901|T201|COMP|59978-7|LNC|Venlafaxine|Venlafaxine
C2969902|T201|COMP|59979-5|LNC|Warfarin|Warfarin
C2969903|T201|COMP|59980-3|LNC|Warfarin|Warfarin
C2969904|T201|COMP|59981-1|LNC|Zopiclone|Zopiclone
C2969905|T201|COMP|59982-9|LNC|Zopiclone|Zopiclone
C2969911|T201|COMP|59988-6|LNC|Testosterone^8th specimen post XXX challenge|Testosterone^8th specimen post XXX challenge
C2969912|T201|COMP|59989-4|LNC|Testosterone^7th specimen post XXX challenge|Testosterone^7th specimen post XXX challenge
C2969913|T201|COMP|59990-2|LNC|Testosterone^6th specimen post XXX challenge|Testosterone^6th specimen post XXX challenge
C2969914|T201|COMP|59991-0|LNC|Testosterone^5th specimen post XXX challenge|Testosterone^5th specimen post XXX challenge
C2969915|T201|COMP|59992-8|LNC|Testosterone^4th specimen post XXX challenge|Testosterone^4th specimen post XXX challenge
C2969916|T201|COMP|59993-6|LNC|Testosterone^3rd specimen post XXX challenge|Testosterone^3rd specimen post XXX challenge
C2969917|T201|COMP|59994-4|LNC|Testosterone^2nd specimen post XXX challenge|Testosterone^2nd specimen post XXX challenge
C2969918|T201|COMP|59995-1|LNC|Testosterone^1st specimen post XXX challenge|Testosterone^1st specimen post XXX challenge
C2969934|T201|COMP|60017-1|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2969935|T201|COMP|60018-9|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2969936|T201|COMP|60019-7|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C2969937|T201|COMP|60036-1|LNC|1-Naphthol|1-Naphthol
C2969938|T201|COMP|60037-9|LNC|1-Naphthol|1-Naphthol
C2969939|T201|COMP|60038-7|LNC|1-Naphthol|1-Naphthol
C2969940|T201|COMP|60039-5|LNC|Acebutolol|Acebutolol
C2969941|T201|COMP|60040-3|LNC|Acebutolol|Acebutolol
C2969942|T201|COMP|60041-1|LNC|Acebutolol|Acebutolol
C2969943|T201|COMP|60042-9|LNC|N-acetylprocainamide|N-acetylprocainamide
C2969944|T201|COMP|60043-7|LNC|Acepromazine|Acepromazine
C2969945|T201|COMP|60044-5|LNC|Acepromazine|Acepromazine
C2969946|T201|COMP|60045-2|LNC|Acetaldehyde|Acetaldehyde
C2969947|T201|COMP|60046-0|LNC|Acetaldehyde|Acetaldehyde
C2969948|T201|COMP|60047-8|LNC|Acetaldehyde|Acetaldehyde
C2969949|T201|COMP|60048-6|LNC|Acetaminophen|Acetaminophen
C2969950|T201|COMP|60049-4|LNC|Acetaminophen|Acetaminophen
C2969951|T201|COMP|60050-2|LNC|Acetaminophen|Acetaminophen
C2969952|T201|COMP|60051-0|LNC|Acetophenazine|Acetophenazine
C2969953|T201|COMP|60052-8|LNC|Alphapinene|Alphapinene
C2969954|T201|COMP|60053-6|LNC|aMILoride|aMILoride
C2969955|T201|COMP|60054-4|LNC|Amiodarone|Amiodarone
C2969956|T201|COMP|60055-1|LNC|Astemizole|Astemizole
C2969957|T201|COMP|60056-9|LNC|Astemizole|Astemizole
C2969958|T201|COMP|60057-7|LNC|Bismuth|Bismuth
C2969959|T201|COMP|60058-5|LNC|Bismuth|Bismuth
C2969960|T201|COMP|60059-3|LNC|Bismuth|Bismuth
C2969961|T201|COMP|60060-1|LNC|Boron|Boron
C2969962|T201|COMP|60061-9|LNC|buPROPion|buPROPion
C2969963|T201|COMP|60062-7|LNC|buPROPion|buPROPion
C2969964|T201|COMP|60063-5|LNC|buPROPion|buPROPion
C2969965|T201|COMP|60064-3|LNC|buPROPion|buPROPion
C2969966|T201|COMP|60065-0|LNC|Cobalt|Cobalt
C2969967|T201|COMP|60066-8|LNC|Cobalt|Cobalt
C2969968|T201|COMP|60067-6|LNC|Cobalt|Cobalt
C2969969|T201|COMP|60068-4|LNC|Colchicine|Colchicine
C2969970|T201|COMP|60069-2|LNC|Dantrolene|Dantrolene
C2969971|T201|COMP|60070-0|LNC|Dichlorvos|Dichlorvos
C2969972|T201|COMP|60071-8|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C2969973|T201|COMP|60072-6|LNC|Fexofenadine|Fexofenadine
C2969974|T201|COMP|60073-4|LNC|Fexofenadine|Fexofenadine
C2969975|T201|COMP|60074-2|LNC|Fexofenadine|Fexofenadine
C2969976|T201|COMP|60075-9|LNC|Finasteride|Finasteride
C2969977|T201|COMP|60076-7|LNC|Gallium|Gallium
C2969978|T201|COMP|60077-5|LNC|Ganciclovir|Ganciclovir
C2969979|T201|COMP|60078-3|LNC|Ganciclovir|Ganciclovir
C2969980|T201|COMP|60079-1|LNC|Germanium|Germanium
C2969981|T201|COMP|60090-8|LNC|Indium|Indium
C2969982|T201|COMP|60091-6|LNC|Ketoconazole|Ketoconazole
C2969983|T201|COMP|60092-4|LNC|Ketoconazole|Ketoconazole
C2969984|T201|COMP|60093-2|LNC|Ketoprofen|Ketoprofen
C2969985|T201|COMP|60094-0|LNC|Ketoprofen|Ketoprofen
C2969986|T201|COMP|60095-7|LNC|Loperamide|Loperamide
C2969987|T201|COMP|60096-5|LNC|Loperamide|Loperamide
C2969988|T201|COMP|60097-3|LNC|Loratadine|Loratadine
C2969989|T201|COMP|60098-1|LNC|Loratadine|Loratadine
C2969990|T201|COMP|60099-9|LNC|Loxapine|Loxapine
C2969991|T201|COMP|60100-5|LNC|Loxapine|Loxapine
C2969992|T201|COMP|60101-3|LNC|Molybdenum|Molybdenum
C2969993|T201|COMP|60102-1|LNC|Norvenlafaxine|Norvenlafaxine
C2969994|T201|COMP|60103-9|LNC|Norvenlafaxine|Norvenlafaxine
C2969995|T201|COMP|60104-7|LNC|Norvenlafaxine|Norvenlafaxine
C2969996|T201|COMP|60105-4|LNC|OLANZapine|OLANZapine
C2969997|T201|COMP|60106-2|LNC|OLANZapine|OLANZapine
C2969998|T201|COMP|60107-0|LNC|OLANZapine|OLANZapine
C2969999|T201|COMP|60108-8|LNC|Oxychlordane|Oxychlordane
C2970000|T201|COMP|60109-6|LNC|Oxychlordane|Oxychlordane
C2970001|T201|COMP|60110-4|LNC|Oxyphenbutazone|Oxyphenbutazone
C2970002|T201|COMP|60111-2|LNC|Oxyphenbutazone|Oxyphenbutazone
C2970003|T201|COMP|60112-0|LNC|Oxipurinol|Oxipurinol
C2970004|T201|COMP|60113-8|LNC|Oxypurinol|Oxypurinol
C2970005|T201|COMP|60114-6|LNC|PACLitaxel|PACLitaxel
C2970006|T201|COMP|60115-3|LNC|9-Hydroxyrisperidone|9-Hydroxyrisperidone
C2970007|T201|COMP|60116-1|LNC|9-Hydroxyrisperidone|9-Hydroxyrisperidone
C2970008|T201|COMP|60117-9|LNC|Palladium|Palladium
C2970009|T201|COMP|60118-7|LNC|Palladium|Palladium
C2970010|T201|COMP|60119-5|LNC|Palladium|Palladium
C2970011|T201|COMP|60120-3|LNC|Palladium|Palladium
C2970012|T201|COMP|60121-1|LNC|Pancuronium|Pancuronium
C2970013|T201|COMP|60122-9|LNC|Pancuronium|Pancuronium
C2970014|T201|COMP|60123-7|LNC|Pancuronium|Pancuronium
C2970015|T201|COMP|60124-5|LNC|Pancuronium|Pancuronium
C2970016|T201|COMP|60125-2|LNC|Papaverine|Papaverine
C2970017|T201|COMP|60126-0|LNC|Papaverine|Papaverine
C2970018|T201|COMP|60127-8|LNC|Paramethadione|Paramethadione
C2970019|T201|COMP|60128-6|LNC|Paramethadione|Paramethadione
C2970020|T201|COMP|60129-4|LNC|Paraoxon|Paraoxon
C2970021|T201|COMP|60130-2|LNC|Paraoxon|Paraoxon
C2970022|T201|COMP|60131-0|LNC|Paraoxon|Paraoxon
C2970023|T201|COMP|60132-8|LNC|Parathion|Parathion
C2970024|T201|COMP|60133-6|LNC|Parathion|Parathion
C2970025|T201|COMP|60134-4|LNC|Parathion|Parathion
C2970026|T201|COMP|60135-1|LNC|Pargyline|Pargyline
C2970027|T201|COMP|60136-9|LNC|PARoxetine|PARoxetine
C2970028|T201|COMP|60137-7|LNC|PARoxetine|PARoxetine
C2970029|T201|COMP|60138-5|LNC|PARoxetine|PARoxetine
C2970030|T201|COMP|60139-3|LNC|Pemoline|Pemoline
C2970031|T201|COMP|60140-1|LNC|Penciclovir|Penciclovir
C2970032|T201|COMP|60141-9|LNC|Penciclovir|Penciclovir
C2970033|T201|COMP|60142-7|LNC|Pendimethalin|Pendimethalin
C2970034|T201|COMP|60143-5|LNC|Pendimethalin|Pendimethalin
C2970035|T201|COMP|60144-3|LNC|Pendimethalin|Pendimethalin
C2970036|T201|COMP|60145-0|LNC|Pentane|Pentane
C2970037|T201|COMP|60146-8|LNC|Pentane|Pentane
C2970038|T201|COMP|60147-6|LNC|Pentane|Pentane
C2970039|T201|COMP|60148-4|LNC|Pentane|Pentane
C2970040|T201|COMP|60149-2|LNC|Pentazocine|Pentazocine
C2970041|T201|COMP|60150-0|LNC|Pentazocine|Pentazocine
C2970042|T201|COMP|60151-8|LNC|PENTobarbital|PENTobarbital
C2970043|T201|COMP|60152-6|LNC|PENTobarbital|PENTobarbital
C2970044|T201|COMP|60153-4|LNC|PENTobarbital|PENTobarbital
C2970045|T201|COMP|60154-2|LNC|Pentoxifylline|Pentoxifylline
C2970046|T201|COMP|60155-9|LNC|Pentoxifylline|Pentoxifylline
C2970047|T201|COMP|60156-7|LNC|Perfluorooctanoate|Perfluorooctanoate
C2970048|T201|COMP|60157-5|LNC|Perfluorooctanoate|Perfluorooctanoate
C2970049|T201|COMP|60158-3|LNC|Pergolide|Pergolide
C2970050|T201|COMP|60159-1|LNC|Pergolide|Pergolide
C2970051|T201|COMP|60160-9|LNC|Perphenazine|Perphenazine
C2970052|T201|COMP|60161-7|LNC|Phenacemide|Phenacemide
C2970053|T201|COMP|60162-5|LNC|Phenacemide|Phenacemide
C2970054|T201|COMP|60163-3|LNC|Phenolphthalein|Phenolphthalein
C2970055|T201|COMP|60164-1|LNC|Phensuximide|Phensuximide
C2970056|T201|COMP|60165-8|LNC|Phensuximide|Phensuximide
C2970057|T201|COMP|60166-6|LNC|Platinum|Platinum
C2970058|T201|COMP|60167-4|LNC|Platinum|Platinum
C2970059|T201|COMP|60168-2|LNC|Platinum|Platinum
C2970060|T201|COMP|60169-0|LNC|Rubidium|Rubidium
C2970061|T201|COMP|60170-8|LNC|Silicon|Silicon
C2970062|T201|COMP|60171-6|LNC|Silicon|Silicon
C2970063|T201|COMP|60194-8|LNC|Triamterene|Triamterene
C2970064|T201|COMP|60195-5|LNC|Trichlormethiazide|Trichlormethiazide
C2970065|T201|COMP|60196-3|LNC|Trichlormethiazide|Trichlormethiazide
C2970066|T201|COMP|60197-1|LNC|Triclopyr|Triclopyr
C2970067|T201|COMP|60198-9|LNC|Trifluralin|Trifluralin
C2970068|T201|COMP|60199-7|LNC|Trifluralin|Trifluralin
C2970069|T201|COMP|60200-3|LNC|Trifluralin|Trifluralin
C2970070|T201|COMP|60212-8|LNC|Zolazepam|Zolazepam
C2970071|T201|COMP|60213-6|LNC|Zolazepam|Zolazepam
C2970072|T201|COMP|60235-9|LNC|Hydrogen/Expired gas^1.25H post dose lactose PO|Hydrogen/Expired gas^1.25H post dose lactose PO
C2970075|T201|COMP|60237-5|LNC|Fraxinus excelsior Ab.IgE.RAST class|Fraxinus excelsior Ab.IgE.RAST class
C2970077|T201|COMP|60238-3|LNC|Fraxinus excelsior Ab.IgE|Fraxinus excelsior Ab.IgE
C2970081|T201|COMP|60240-9|LNC|Vespula vulgaris recombinant (rVes v) 5 Ab.IgE|Vespula vulgaris recombinant (rVes v) 5 Ab.IgE
C2970085|T201|COMP|60242-5|LNC|Coagulation ecarin induced|Coagulation ecarin induced
C2970086|T201|COMP|60243-3|LNC|Matrix metallopeptidase 9|Matrix metallopeptidase 9
C2970087|T201|COMP|60244-1|LNC|Androstanolone^8th specimen post XXX challenge|Androstanolone^8th specimen post XXX challenge
C2970088|T201|COMP|60245-8|LNC|Androstanolone^7th specimen post XXX challenge|Androstanolone^7th specimen post XXX challenge
C2970089|T201|COMP|60246-6|LNC|Androstanolone^6th specimen post XXX challenge|Androstanolone^6th specimen post XXX challenge
C2970090|T201|COMP|60247-4|LNC|Androstanolone^5th specimen post XXX challenge|Androstanolone^5th specimen post XXX challenge
C2970091|T201|COMP|60248-2|LNC|Androstanolone^4th specimen post XXX challenge|Androstanolone^4th specimen post XXX challenge
C2970092|T201|COMP|60249-0|LNC|Androstanolone^3rd specimen post XXX challenge|Androstanolone^3rd specimen post XXX challenge
C2970093|T201|COMP|60250-8|LNC|Androstanolone^2nd specimen post XXX challenge|Androstanolone^2nd specimen post XXX challenge
C2970094|T201|COMP|60251-6|LNC|Androstanolone^1st specimen post XXX challenge|Androstanolone^1st specimen post XXX challenge
C2970095|T201|COMP|60252-4|LNC|MGMT gene methylation|MGMT gene methylation
C2970096|T201|COMP|60253-2|LNC|DNA index 4|DNA index 4
C2970097|T201|COMP|60254-0|LNC|Parainfluenza virus 1+2+3 RNA|Parainfluenza virus 1+2+3 RNA
C2970098|T201|COMP|60255-7|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2970099|T201|COMP|60256-5|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2970100|T201|COMP|60257-3|LNC|Bacteria identified|Bacteria identified
C2970101|T201|COMP|60258-1|LNC|Bacteria identified|Bacteria identified
C2970102|T201|COMP|60259-9|LNC|Adenovirus DNA|Adenovirus DNA
C2970103|T201|COMP|60260-7|LNC|Chikungunya virus RNA|Chikungunya virus RNA
C2970104|T201|COMP|60261-5|LNC|Coxiella burnetii DNA|Coxiella burnetii DNA
C2970105|T201|COMP|60262-3|LNC|Dengue virus 1 RNA|Dengue virus 1 RNA
C2970106|T201|COMP|60263-1|LNC|Enterovirus RNA|Enterovirus RNA
C2970107|T201|COMP|60264-9|LNC|Hantavirus Ab|Hantavirus Ab
C2970108|T201|COMP|60265-6|LNC|Human coronavirus RNA|Human coronavirus RNA
C2970109|T201|COMP|60266-4|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C2970110|T201|COMP|60267-2|LNC|Influenza virus C RNA|Influenza virus C RNA
C2970111|T201|COMP|60268-0|LNC|Orientia tsutsugamushi DNA|Orientia tsutsugamushi DNA
C2970112|T201|COMP|60269-8|LNC|Parainfluenza virus 1 RNA|Parainfluenza virus 1 RNA
C2970113|T201|COMP|60270-6|LNC|Rabies virus RNA|Rabies virus RNA
C2970114|T201|COMP|60271-4|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C2970115|T201|COMP|60272-2|LNC|Rickettsia typhus group DNA|Rickettsia typhus group DNA
C2970116|T201|COMP|60273-0|LNC|Rotavirus RNA|Rotavirus RNA
C2970117|T201|COMP|60274-8|LNC|Rubella virus RNA|Rubella virus RNA
C2970118|T201|COMP|60275-5|LNC|SARS coronavirus RNA|SARS coronavirus RNA
C2970119|T201|COMP|60276-3|LNC|oxyCODONE+Oxymorphone cutoff|oxyCODONE+Oxymorphone cutoff
C2970121|T201|COMP|60277-1|LNC|Complement C3 Ag|Complement C3 Ag
C2970122|T201|COMP|60278-9|LNC|Fibrinogen Ag|Fibrinogen Ag
C2970123|T201|COMP|60279-7|LNC|IL28B gene associated variant rs12979860|IL28B gene associated variant rs12979860
C2970127|T201|COMP|60282-1|LNC|ALPRAZolam|ALPRAZolam
C2970128|T201|COMP|60283-9|LNC|Amitriptyline|Amitriptyline
C2970129|T201|COMP|60284-7|LNC|Amobarbital|Amobarbital
C2970130|T201|COMP|60285-4|LNC|Amoxapine|Amoxapine
C2970131|T201|COMP|60286-2|LNC|Ascorbate|Ascorbate
C2970132|T201|COMP|60287-0|LNC|Benztropine|Benztropine
C2970133|T201|COMP|60288-8|LNC|Bromazepam|Bromazepam
C2970134|T201|COMP|60289-6|LNC|Brompheniramine|Brompheniramine
C2970135|T201|COMP|60290-4|LNC|Caffeine|Caffeine
C2970136|T201|COMP|60291-2|LNC|carBAMazepine|carBAMazepine
C2970137|T201|COMP|60292-0|LNC|Chloral hydrate|Chloral hydrate
C2970138|T201|COMP|60293-8|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C2970139|T201|COMP|60294-6|LNC|chlorproMAZINE|chlorproMAZINE
C2970140|T201|COMP|60295-3|LNC|Citalopram|Citalopram
C2970141|T201|COMP|60296-1|LNC|cloBAZam|cloBAZam
C2970142|T201|COMP|60297-9|LNC|clomiPRAMINE|clomiPRAMINE
C2970143|T201|COMP|60298-7|LNC|cloZAPine|cloZAPine
C2970144|T201|COMP|60299-5|LNC|Cotinine|Cotinine
C2970145|T201|COMP|60300-1|LNC|Desipramine|Desipramine
C2970146|T201|COMP|60301-9|LNC|Disopyramide|Disopyramide
C2970147|T201|COMP|60302-7|LNC|Doxepin|Doxepin
C2970148|T201|COMP|60303-5|LNC|Fenoprofen|Fenoprofen
C2970149|T201|COMP|60304-3|LNC|FLUoxetine|FLUoxetine
C2970150|T201|COMP|60305-0|LNC|fluPHENAZine|fluPHENAZine
C2970151|T201|COMP|60306-8|LNC|fluvoxaMINE|fluvoxaMINE
C2970152|T201|COMP|60307-6|LNC|hydrOXYzine|hydrOXYzine
C2970153|T201|COMP|60308-4|LNC|Ibuprofen|Ibuprofen
C2970154|T201|COMP|60319-1|LNC|Naproxen|Naproxen
C2970155|T201|COMP|60320-9|LNC|Nicotine|Nicotine
C2970156|T201|COMP|60321-7|LNC|Norclobazam|Norclobazam
C2970157|T201|COMP|60322-5|LNC|Norclomipramine|Norclomipramine
C2970158|T201|COMP|60323-3|LNC|Nordoxepin|Nordoxepin
C2970159|T201|COMP|60324-1|LNC|Nortriptyline|Nortriptyline
C2970160|T201|COMP|60325-8|LNC|OLANZapine|OLANZapine
C2970161|T201|COMP|60326-6|LNC|OXcarbazepine|OXcarbazepine
C2970162|T201|COMP|60327-4|LNC|PARoxetine|PARoxetine
C2970163|T201|COMP|60328-2|LNC|Pentazocine|Pentazocine
C2970164|T201|COMP|60329-0|LNC|Promazine|Promazine
C2970165|T201|COMP|60330-8|LNC|Propoxyphene|Propoxyphene
C2970166|T201|COMP|60331-6|LNC|Propranolol|Propranolol
C2970167|T201|COMP|60332-4|LNC|QUEtiapine|QUEtiapine
C2970168|T201|COMP|60333-2|LNC|Sulfamethoxazole|Sulfamethoxazole
C2970169|T201|COMP|60334-0|LNC|Thiocyanate|Thiocyanate
C2970170|T201|COMP|60335-7|LNC|traZODone|traZODone
C2970171|T201|COMP|60336-5|LNC|Trimipramine|Trimipramine
C2970172|T201|COMP|60337-3|LNC|Venlafaxine|Venlafaxine
C2970173|T201|COMP|60338-1|LNC|Warfarin|Warfarin
C2970174|T201|COMP|60339-9|LNC|Zopiclone|Zopiclone
C2970175|T201|COMP|60340-7|LNC|Crystals.amorphous|Crystals.amorphous
C2970176|T201|COMP|60348-0|LNC|Prunus dulcis Ab.IgG|Prunus dulcis Ab.IgG
C2970177|T201|COMP|60349-8|LNC|Malus sylvestris Ab.IgG|Malus sylvestris Ab.IgG
C2970178|T201|COMP|60350-6|LNC|Prunus armeniaca Ab.IgG|Prunus armeniaca Ab.IgG
C2970179|T201|COMP|60351-4|LNC|Cynara scolymus Ab.IgG|Cynara scolymus Ab.IgG
C2970180|T201|COMP|60352-2|LNC|Musa spp Ab.IgG|Musa spp Ab.IgG
C2970181|T201|COMP|60353-0|LNC|Bean green Ab.IgG|Bean green Ab.IgG
C2970182|T201|COMP|60354-8|LNC|Bean kidney red Ab.IgG|Bean kidney red Ab.IgG
C2970183|T201|COMP|60355-5|LNC|Bean pinto Ab.IgG|Bean pinto Ab.IgG
C2970184|T201|COMP|60356-3|LNC|Brassica oleracea var italica Ab.IgG|Brassica oleracea var italica Ab.IgG
C2970185|T201|COMP|60357-1|LNC|Brassica oleracea var gemmifera Ab.IgG|Brassica oleracea var gemmifera Ab.IgG
C2970186|T201|COMP|60358-9|LNC|Brassica oleracea var capitata Ab.IgG|Brassica oleracea var capitata Ab.IgG
C2970187|T201|COMP|60359-7|LNC|Cucumis melo cantalupensis Ab.IgG|Cucumis melo cantalupensis Ab.IgG
C2970188|T201|COMP|60360-5|LNC|Daucus carota Ab.IgG|Daucus carota Ab.IgG
C2970189|T201|COMP|60361-3|LNC|Brassica oleracea var botrytis Ab.IgG|Brassica oleracea var botrytis Ab.IgG
C2970190|T201|COMP|60362-1|LNC|Asparagus officinalis Ab.IgG|Asparagus officinalis Ab.IgG
C2970191|T201|COMP|60363-9|LNC|Apium graveolens Ab.IgG|Apium graveolens Ab.IgG
C2970192|T201|COMP|60364-7|LNC|Cheese mold type Ab.IgG|Cheese mold type Ab.IgG
C2970193|T201|COMP|60365-4|LNC|Prunus avium Ab.IgG|Prunus avium Ab.IgG
C2970194|T201|COMP|60366-2|LNC|Capsicum frutescens Ab.IgG|Capsicum frutescens Ab.IgG
C2970195|T201|COMP|60367-0|LNC|Cinnamomum spp Ab.IgG|Cinnamomum spp Ab.IgG
C2970196|T201|COMP|60368-8|LNC|Ruditapes spp Ab.IgG|Ruditapes spp Ab.IgG
C2970197|T201|COMP|60369-6|LNC|Syzygium aromaticum Ab.IgG|Syzygium aromaticum Ab.IgG
C2970198|T201|COMP|60370-4|LNC|Cancer pagurus Ab.IgG|Cancer pagurus Ab.IgG
C2970199|T201|COMP|60371-2|LNC|Cucumis sativus Ab.IgG|Cucumis sativus Ab.IgG
C2970200|T201|COMP|60372-0|LNC|Solanum melongena Ab.IgG|Solanum melongena Ab.IgG
C2970201|T201|COMP|60373-8|LNC|Flounder Ab.IgG|Flounder Ab.IgG
C2970202|T201|COMP|60374-6|LNC|Allium sativum Ab.IgG|Allium sativum Ab.IgG
C2970203|T201|COMP|60375-3|LNC|Zingiber officinale Ab.IgG|Zingiber officinale Ab.IgG
C2970204|T201|COMP|60395-1|LNC|Prunus domestica Ab.IgG|Prunus domestica Ab.IgG
C2970205|T201|COMP|60396-9|LNC|Ipomoea batatas Ab.IgG|Ipomoea batatas Ab.IgG
C2970206|T201|COMP|60397-7|LNC|Raphanus sativus Ab.IgG|Raphanus sativus Ab.IgG
C2970207|T201|COMP|60398-5|LNC|Persea americana Ab.IgG|Persea americana Ab.IgG
C2970208|T201|COMP|60399-3|LNC|Salvia officinalis Ab.IgG|Salvia officinalis Ab.IgG
C2970209|T201|COMP|60400-9|LNC|Salmo salar Ab.IgG|Salmo salar Ab.IgG
C2970210|T201|COMP|60401-7|LNC|Pecten spp Ab.IgG|Pecten spp Ab.IgG
C2970211|T201|COMP|60402-5|LNC|Sesamum indicum Ab.IgG|Sesamum indicum Ab.IgG
C2970212|T201|COMP|60403-3|LNC|Pandalus borealis Ab.IgG|Pandalus borealis Ab.IgG
C2970213|T201|COMP|60404-1|LNC|Snapper red Ab.IgG|Snapper red Ab.IgG
C2970214|T201|COMP|60405-8|LNC|Solea solea Ab.IgG|Solea solea Ab.IgG
C2970215|T201|COMP|60406-6|LNC|Spinacia oleracea Ab.IgG|Spinacia oleracea Ab.IgG
C2970216|T201|COMP|60407-4|LNC|Helianthus annuus seed Ab.IgG|Helianthus annuus seed Ab.IgG
C2970217|T201|COMP|60408-2|LNC|Citrus reticulata Ab.IgG|Citrus reticulata Ab.IgG
C2970218|T201|COMP|60409-0|LNC|Oncorhynchus mykiss Ab.IgG|Oncorhynchus mykiss Ab.IgG
C2970219|T201|COMP|60410-8|LNC|Thunnus albacares Ab.IgG|Thunnus albacares Ab.IgG
C2970220|T201|COMP|60411-6|LNC|Turkey Ab.IgG|Turkey Ab.IgG
C2970221|T201|COMP|60412-4|LNC|Vanilla planifolia Ab.IgG|Vanilla planifolia Ab.IgG
C2970222|T201|COMP|60413-2|LNC|Yeast brewer's Ab.IgG|Yeast brewer's Ab.IgG
C2970223|T201|COMP|60414-0|LNC|Squash zucchini Ab.IgG|Squash zucchini Ab.IgG
C2970224|T201|COMP|60415-7|LNC|Parainfluenza virus 4 RNA|Parainfluenza virus 4 RNA
C2970225|T201|COMP|60416-5|LNC|Parainfluenza virus 3 RNA|Parainfluenza virus 3 RNA
C2970226|T201|COMP|60417-3|LNC|Parainfluenza virus 2 RNA|Parainfluenza virus 2 RNA
C2970227|T201|COMP|60418-1|LNC|Dengue virus 4 RNA|Dengue virus 4 RNA
C2970228|T201|COMP|60419-9|LNC|Dengue virus 3 RNA|Dengue virus 3 RNA
C2970229|T201|COMP|60420-7|LNC|Dengue virus 2 RNA|Dengue virus 2 RNA
C2970232|T201|COMP|60422-3|LNC|Measles virus genotype|Measles virus genotype
C2970233|T201|COMP|60423-1|LNC|Measles virus identified|Measles virus identified
C2970234|T201|COMP|60424-9|LNC|Parainfluenza virus 4 Ag|Parainfluenza virus 4 Ag
C2970235|T201|COMP|60425-6|LNC|Human metapneumovirus Ag|Human metapneumovirus Ag
C2970236|T201|COMP|60426-4|LNC|SARS coronavirus Ab|SARS coronavirus Ab
C2970237|T201|COMP|60427-2|LNC|Norovirus RNA|Norovirus RNA
C2970238|T201|COMP|60428-0|LNC|Toxoplasma gondii Ab.IgA|Toxoplasma gondii Ab.IgA
C2970239|T201|COMP|60429-8|LNC|Enterovirus 71 RNA|Enterovirus 71 RNA
C2970240|T201|COMP|60430-6|LNC|Hepatitis E virus genotype|Hepatitis E virus genotype
C2970244|T201|COMP|60433-0|LNC|Leukocytes|Leukocytes
C2970245|T201|COMP|60434-8|LNC|Cells.CD19+CD103+|Cells.CD19+CD103+
C2970249|T201|COMP|60454-6|LNC|Bixa orellana seed Ab.IgE.RAST class|Bixa orellana seed Ab.IgE.RAST class
C2970251|T201|COMP|60455-3|LNC|Bizarre platelets|Bizarre platelets
C2970252|T201|COMP|60456-1|LNC|Cells.CD3+CD8+CD57+/100 cells|Cells.CD3+CD8+CD57+/100 cells
C2970254|T201|COMP|60457-9|LNC|Cells.CD4+CD26-|Cells.CD4+CD26-
C2970255|T201|COMP|60458-7|LNC|Collection time^6th specimen|Collection time^6th specimen
C2970256|T201|COMP|61139-2|LNC|Toluene diisocyanate (TDI) Ab.IgG|Toluene diisocyanate (TDI) Ab.IgG
C2970257|T201|COMP|61140-0|LNC|Diphenylmethane diisocyanate (MDI) Ab.IgG|Diphenylmethane diisocyanate (MDI) Ab.IgG
C2970258|T201|COMP|60465-2|LNC|Neisseria meningitidis serogroup w135 Ab.IgG|Neisseria meningitidis serogroup w135 Ab.IgG
C2970259|T201|COMP|60466-0|LNC|Neisseria meningitidis serogroup Y Ab.IgG|Neisseria meningitidis serogroup Y Ab.IgG
C2970260|T201|COMP|60467-8|LNC|oxyMORphone|oxyMORphone
C2970261|T201|COMP|60468-6|LNC|PHENobarbital|PHENobarbital
C2970262|T201|COMP|60469-4|LNC|Urate|Urate
C2970263|T201|COMP|60470-2|LNC|Toxocara canis Ab|Toxocara canis Ab
C2970264|T201|COMP|60471-0|LNC|busPIRone|busPIRone
C2970265|T201|COMP|60472-8|LNC|Complement C5.functional|Complement C5.functional
C2970266|T201|COMP|60473-6|LNC|Lymphocytes.vacuolated|Lymphocytes.vacuolated
C2970267|T201|COMP|60474-4|LNC|Reticulocytes|Reticulocytes
C2970269|T201|COMP|60486-8|LNC|MED12 gene targeted mutation analysis|MED12 gene targeted mutation analysis
C2970271|T201|COMP|60487-6|LNC|NPHP1 gene targeted mutation analysis|NPHP1 gene targeted mutation analysis
C2970273|T201|COMP|60488-4|LNC|NPHS2 gene targeted mutation analysis|NPHS2 gene targeted mutation analysis
C2970275|T201|COMP|60489-2|LNC|Streptococcus pyogenes DNA|Streptococcus pyogenes DNA
C2970276|T201|COMP|60490-0|LNC|UMOD gene targeted mutation analysis|UMOD gene targeted mutation analysis
C2970278|T201|COMP|60491-8|LNC|LCA gene targeted mutation analysis|LCA gene targeted mutation analysis
C2970282|T201|COMP|60493-4|LNC|Calcidiol+Calciferol|Calcidiol+Calciferol
C2970284|T201|COMP|60495-9|LNC|MAP2K1 gene targeted mutation analysis|MAP2K1 gene targeted mutation analysis
C2970286|T201|COMP|60496-7|LNC|MAP2K2 gene targeted mutation analysis|MAP2K2 gene targeted mutation analysis
C2970288|T201|COMP|60497-5|LNC|SLC22A5 gene targeted mutation analysis|SLC22A5 gene targeted mutation analysis
C2970306|T201|COMP|60514-7|LNC|6-Acetylcodeine|6-Acetylcodeine
C2970307|T201|COMP|60525-3|LNC|Parechovirus RNA|Parechovirus RNA
C2970308|T201|COMP|60526-1|LNC|Pseudo Pelger Huet cells|Pseudo Pelger Huet cells
C2970310|T201|COMP|60528-7|LNC|Enterovirus subtype|Enterovirus subtype
C2970311|T201|COMP|60529-5|LNC|Influenza virus A H1 2009 pandemic Ab|Influenza virus A H1 2009 pandemic Ab
C2970312|T201|COMP|60530-3|LNC|Influenza virus A H9 RNA|Influenza virus A H9 RNA
C2970313|T201|COMP|60531-1|LNC|Japanese encephalitis virus Ab.IgM|Japanese encephalitis virus Ab.IgM
C2970314|T201|COMP|60532-9|LNC|Japanese encephalitis virus Ab.IgM|Japanese encephalitis virus Ab.IgM
C2970315|T201|COMP|60533-7|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C2970316|T201|COMP|60534-5|LNC|SARS coronavirus RNA|SARS coronavirus RNA
C2970317|T201|COMP|60535-2|LNC|Doripenem|Doripenem
C2970318|T201|COMP|60536-0|LNC|HLA-DQ beta|HLA-DQ beta
C2970319|T201|COMP|60537-8|LNC|CLCN5 gene targeted mutation analysis|CLCN5 gene targeted mutation analysis
C2970321|T201|COMP|60538-6|LNC|Influenza virus A H1+H3+B RNA|Influenza virus A H1+H3+B RNA
C2970322|T201|COMP|60539-4|LNC|Tryptase.beta|Tryptase.beta
C2970323|T201|COMP|60540-2|LNC|HBA2 gene targeted mutation analysis|HBA2 gene targeted mutation analysis
C2970325|T201|COMP|60541-0|LNC|Cytomegalovirus early Ag|Cytomegalovirus early Ag
C2970326|T201|COMP|60542-8|LNC|Mupirocin 5 ug|Mupirocin 5 ug
C2970327|T201|COMP|60543-6|LNC|Mupirocin 200 ug|Mupirocin 200 ug
C2970328|T201|COMP|60544-4|LNC|Giardia lamblia DNA|Giardia lamblia DNA
C2970329|T201|COMP|60545-1|LNC|Cryptosporidium sp DNA|Cryptosporidium sp DNA
C2970330|T201|COMP|60546-9|LNC|Polio virus identified|Polio virus identified
C2970331|T201|COMP|60547-7|LNC|11-Oxo-Androsterone/Creatinine|11-Oxo-Androsterone/Creatinine
C2970332|T201|COMP|60548-5|LNC|11-Oxo-Etiocholanolone/Creatinine|11-Oxo-Etiocholanolone/Creatinine
C2970333|T201|COMP|60549-3|LNC|8-Estriol|8-Estriol
C2970334|T201|COMP|60550-1|LNC|Fascin|Fascin
C2970335|T201|COMP|60551-9|LNC|Interferon.beta 1a Ab|Interferon.beta 1a Ab
C2970336|T201|COMP|60552-7|LNC|Interferon.beta 1b Ab|Interferon.beta 1b Ab
C2970337|T201|COMP|60553-5|LNC|Trypanosoma cruzi Ab|Trypanosoma cruzi Ab
C2970338|T201|COMP|60554-3|LNC|Monocytes.CD59 deficient/100 cells|Monocytes.CD59 deficient/100 cells
C2970349|T201|COMP|60564-2|LNC|Amikacin 1.0 ug/mL|Amikacin 1.0 ug/mL
C2970351|T201|COMP|60565-9|LNC|Amikacin 4.0 ug/mL|Amikacin 4.0 ug/mL
C2970353|T201|COMP|60566-7|LNC|Respiratory pathogens DNA & RNA 12b panel|Respiratory pathogens DNA & RNA 12b panel
C2970355|T201|COMP|60568-3|LNC|Synoptic report|Synoptic report
C2970356|T201|COMP|60569-1|LNC|Report addendum.synoptic|Report addendum.synoptic
C2970357|T201|COMP|60570-9|LNC|Consultation note|Consultation note
C2970358|T201|COMP|60571-7|LNC|Consultation note.synoptic|Consultation note.synoptic
C2970362|T201|COMP|60575-8|LNC|Immunoglobulin heavy chain gene rearrangements|Immunoglobulin heavy chain gene rearrangements
C2970363|T201|COMP|60577-4|LNC|SERPINE1 gene targeted mutation analysis|SERPINE1 gene targeted mutation analysis
C2970364|T201|COMP|60578-2|LNC|TCRG gene rearrangements|TCRG gene rearrangements
C2970365|T201|COMP|60579-0|LNC|TCRG gene rearrangements|TCRG gene rearrangements
C2970366|T201|COMP|60580-8|LNC|TCRG gene rearrangements|TCRG gene rearrangements
C2970367|T201|COMP|60581-6|LNC|TCRB gene rearrangements|TCRB gene rearrangements
C2970368|T201|COMP|60582-4|LNC|TCRB gene rearrangements|TCRB gene rearrangements
C2970369|T201|COMP|60583-2|LNC|TCRB gene rearrangements|TCRB gene rearrangements
C2970370|T201|COMP|60585-7|LNC|Ganglioside GT1b Ab.IgG|Ganglioside GT1b Ab.IgG
C2970371|T201|COMP|60586-5|LNC|Ganglioside GM3 Ab.IgG|Ganglioside GM3 Ab.IgG
C2970372|T201|COMP|60587-3|LNC|Cell count & Differential panel|Cell count & Differential panel
C2970453|T201|COMP|60676-4|LNC|Ethyl sulfate|Ethyl sulfate
C2970454|T201|COMP|60677-2|LNC|Alpha hydroxytriazolam|Alpha hydroxytriazolam
C2970455|T201|COMP|60680-6|LNC|Cortisol.free^30M post dose corticotropin|Cortisol.free^30M post dose corticotropin
C2970456|T201|COMP|60681-4|LNC|Cortisol.free^1H post dose corticotropin|Cortisol.free^1H post dose corticotropin
C2970462|T201|COMP|61298-6|LNC|Picea excelsa Ab.IgE/IgE.total|Picea excelsa Ab.IgE/IgE.total
C2970463|T201|COMP|61299-4|LNC|Pinus strobus Ab.IgE/IgE.total|Pinus strobus Ab.IgE/IgE.total
C2970464|T201|COMP|61300-0|LNC|Pisum sativum Ab.IgE/IgE.total|Pisum sativum Ab.IgE/IgE.total
C2970465|T201|COMP|61301-8|LNC|Plantago lanceolata Ab.IgE/IgE.total|Plantago lanceolata Ab.IgE/IgE.total
C2970466|T201|COMP|61302-6|LNC|Platanus acerifolia Ab.IgE/IgE.total|Platanus acerifolia Ab.IgE/IgE.total
C2970467|T201|COMP|61303-4|LNC|Poa pratensis Ab.IgE/IgE.total|Poa pratensis Ab.IgE/IgE.total
C2970468|T201|COMP|61304-2|LNC|Populus deltoides Ab.IgE/IgE.total|Populus deltoides Ab.IgE/IgE.total
C2970469|T201|COMP|61305-9|LNC|Prosopis juliflora Ab.IgE/IgE.total|Prosopis juliflora Ab.IgE/IgE.total
C2970476|T201|COMP|61029-5|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2970477|T201|COMP|61030-3|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2970478|T201|COMP|61031-1|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2970479|T201|COMP|61032-9|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C2970480|T201|COMP|61033-7|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C2970481|T201|COMP|61034-5|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C2970482|T201|COMP|61035-2|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2970483|T201|COMP|61036-0|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2970484|T201|COMP|61037-8|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2970485|T201|COMP|61038-6|LNC|ALPRAZolam|ALPRAZolam
C2970486|T201|COMP|61039-4|LNC|clonazePAM|clonazePAM
C2970487|T201|COMP|61040-2|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2970488|T201|COMP|61041-0|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2970489|T201|COMP|61042-8|LNC|fentaNYL|fentaNYL
C2970490|T201|COMP|61043-6|LNC|Ketamine|Ketamine
C2970491|T201|COMP|61044-4|LNC|LORazepam|LORazepam
C2970492|T201|COMP|61045-1|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C2970493|T201|COMP|61046-9|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C2970494|T201|COMP|61047-7|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C2970495|T201|COMP|61048-5|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C2970496|T201|COMP|61049-3|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C2970497|T201|COMP|61050-1|LNC|Methylphenidate|Methylphenidate
C2970498|T201|COMP|61051-9|LNC|Nordiazepam|Nordiazepam
C2970499|T201|COMP|61052-7|LNC|Norfentanyl|Norfentanyl
C2970500|T201|COMP|61053-5|LNC|Norfentanyl|Norfentanyl
C2970501|T201|COMP|61054-3|LNC|Normeperidine|Normeperidine
C2970502|T201|COMP|61055-0|LNC|Oxazepam|Oxazepam
C2970503|T201|COMP|61056-8|LNC|Pseudoephedrine|Pseudoephedrine
C2970504|T201|COMP|61057-6|LNC|Pseudoephedrine|Pseudoephedrine
C2970505|T201|COMP|61058-4|LNC|Alpha-Phenyl-2-Piperidine acetate|Alpha-Phenyl-2-Piperidine acetate
C2970506|T201|COMP|61059-2|LNC|Alpha-Phenyl-2-Piperidine acetate|Alpha-Phenyl-2-Piperidine acetate
C2970507|T201|COMP|61060-0|LNC|Temazepam|Temazepam
C2970508|T201|COMP|61061-8|LNC|Temazepam|Temazepam
C2970509|T201|COMP|61062-6|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C2970510|T201|COMP|61063-4|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C2970511|T201|COMP|61064-2|LNC|Triazolam|Triazolam
C2970512|T201|COMP|61065-9|LNC|Lysergate diethylamide|Lysergate diethylamide
C2970513|T201|COMP|61066-7|LNC|Ethanol|Ethanol
C2970514|T201|COMP|61067-5|LNC|Barbiturates|Barbiturates
C2970515|T201|COMP|61070-9|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C2970516|T201|COMP|61071-7|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C2970517|T201|COMP|61072-5|LNC|Alpha hydroxyalprazolam|Alpha hydroxyalprazolam
C2970518|T201|COMP|61073-3|LNC|ALPRAZolam|ALPRAZolam
C2970519|T201|COMP|61074-1|LNC|diazePAM|diazePAM
C2970520|T201|COMP|61075-8|LNC|diphenhydrAMINE|diphenhydrAMINE
C2970521|T201|COMP|61076-6|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C2970522|T201|COMP|61077-4|LNC|fentaNYL|fentaNYL
C2970523|T201|COMP|61078-2|LNC|Flunitrazepam|Flunitrazepam
C2970524|T201|COMP|61079-0|LNC|Flunitrazepam|Flunitrazepam
C2970525|T201|COMP|61080-8|LNC|Flurazepam|Flurazepam
C2970526|T201|COMP|61081-6|LNC|Ketamine|Ketamine
C2970527|T201|COMP|61082-4|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C2970528|T201|COMP|61083-2|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C2970529|T201|COMP|61084-0|LNC|Methylphenidate|Methylphenidate
C2970530|T201|COMP|61085-7|LNC|Nordiazepam|Nordiazepam
C2970531|T201|COMP|61086-5|LNC|Norfentanyl|Norfentanyl
C2970532|T201|COMP|61087-3|LNC|Normeperidine|Normeperidine
C2970533|T201|COMP|61088-1|LNC|Oxazepam|Oxazepam
C2970534|T201|COMP|61089-9|LNC|Pseudoephedrine|Pseudoephedrine
C2970535|T201|COMP|61090-7|LNC|Alpha-Phenyl-2-Piperidine acetate|Alpha-Phenyl-2-Piperidine acetate
C2970536|T201|COMP|61091-5|LNC|Temazepam|Temazepam
C2970537|T201|COMP|61092-3|LNC|Triazolam|Triazolam
C2970538|T201|COMP|61093-1|LNC|Triazolam|Triazolam
C2970539|T201|COMP|61094-9|LNC|Lysergate diethylamide|Lysergate diethylamide
C2970540|T201|COMP|61095-6|LNC|Ethanol|Ethanol
C2970541|T201|COMP|61096-4|LNC|Barbiturates|Barbiturates
C2970542|T201|COMP|61098-0|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C2970545|T201|COMP|61110-3|LNC|ACSL4 gene targeted mutation analysis|ACSL4 gene targeted mutation analysis
C2970547|T201|COMP|61111-1|LNC|Mitochondria tRNA targeted mutation analysis|Mitochondria tRNA targeted mutation analysis
C2970549|T201|COMP|61112-9|LNC|HTLV|HTLV
C2970550|T201|COMP|61113-7|LNC|Immunoglobulin gene rearrangements|Immunoglobulin gene rearrangements
C2970555|T201|COMP|61116-0|LNC|Mitochondria rRNA targeted mutation analysis|Mitochondria rRNA targeted mutation analysis
C2970557|T201|COMP|61117-8|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C2970558|T201|COMP|61252-3|LNC|Cucurbita pepo seed Ab.IgE/IgE.total|Cucurbita pepo seed Ab.IgE/IgE.total
C2970559|T201|COMP|61253-1|LNC|Cupressus arizonica Ab.IgE/IgE.total|Cupressus arizonica Ab.IgE/IgE.total
C2970560|T201|COMP|61254-9|LNC|Cupressus sempervirens Ab.IgE/IgE.total|Cupressus sempervirens Ab.IgE/IgE.total
C2970561|T201|COMP|61255-6|LNC|Cynodon dactylon Ab.IgE/IgE.total|Cynodon dactylon Ab.IgE/IgE.total
C2970562|T201|COMP|61270-5|LNC|Gluten Ab.IgE/IgE.total|Gluten Ab.IgE/IgE.total
C2970563|T201|COMP|61271-3|LNC|Glycine max Ab.IgE/IgE.total|Glycine max Ab.IgE/IgE.total
C2970564|T201|COMP|61272-1|LNC|Helianthus annuus seed Ab.IgE/IgE.total|Helianthus annuus seed Ab.IgE/IgE.total
C2970565|T201|COMP|61273-9|LNC|Hordeum vulgare Ab.IgE/IgE.total|Hordeum vulgare Ab.IgE/IgE.total
C2970566|T201|COMP|61274-7|LNC|House dust Greer Ab.IgE/IgE.total|House dust Greer Ab.IgE/IgE.total
C2970567|T201|COMP|61275-4|LNC|Humulus lupus Ab.IgE/IgE.total|Humulus lupus Ab.IgE/IgE.total
C2970576|T201|COMP|61118-6|LNC|Lymphocytes.cytoplasmic IgG/100 lymphocytes|Lymphocytes.cytoplasmic IgG/100 lymphocytes
C2970578|T201|COMP|61119-4|LNC|Lymphocytes.cytoplasmic IgM/100 lymphocytes|Lymphocytes.cytoplasmic IgM/100 lymphocytes
C2970580|T201|COMP|61120-2|LNC|PM-SCL-100 Ab.IgG|PM-SCL-100 Ab.IgG
C2970581|T201|COMP|61121-0|LNC|Cells.CD8-CD57+/100 cells|Cells.CD8-CD57+/100 cells
C2970582|T201|COMP|61122-8|LNC|Cells.CD8-CD57+|Cells.CD8-CD57+
C2970583|T201|COMP|61123-6|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C2970584|T201|COMP|61124-4|LNC|Granulocytes/100 leukocytes|Granulocytes/100 leukocytes
C2970585|T201|COMP|61125-1|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C2970586|T201|COMP|61126-9|LNC|Blasts/100 cells|Blasts/100 cells
C2970587|T201|COMP|61127-7|LNC|Whitefish Ab.IgG|Whitefish Ab.IgG
C2970588|T201|COMP|61128-5|LNC|Cotinine|Cotinine
C2970591|T201|COMP|61141-8|LNC|Hexamethylene diisocyanate (HDI) Ab.IgG|Hexamethylene diisocyanate (HDI) Ab.IgG
C2970592|T201|COMP|61142-6|LNC|Trimellitic anhydride Ab.IgG|Trimellitic anhydride Ab.IgG
C2970598|T201|COMP|61151-7|LNC|Albumin|Albumin
C2970599|T201|COMP|61152-5|LNC|Albumin|Albumin
C2970600|T201|COMP|61153-3|LNC|Glucose^baseline|Glucose^baseline
C2970601|T201|COMP|61174-9|LNC|17-Hydroxyprogesterone^20M pre XXX challenge|17-Hydroxyprogesterone^20M pre XXX challenge
C2970602|T201|COMP|61175-6|LNC|Polychlorinated biphenyl.Aroclor 1242|Polychlorinated biphenyl.Aroclor 1242
C2970603|T201|COMP|61176-4|LNC|Polychlorinated biphenyl.Aroclor 1248|Polychlorinated biphenyl.Aroclor 1248
C2970604|T201|COMP|61177-2|LNC|Paraneoplastic Ab|Paraneoplastic Ab
C2970605|T201|COMP|61178-0|LNC|Cells.CD79/100 cells|Cells.CD79/100 cells
C2970607|T201|COMP|61179-8|LNC|Leukocyte morphology finding|Leukocyte morphology finding
C2970608|T201|COMP|61180-6|LNC|Hemoglobin|Hemoglobin
C2970609|T201|COMP|61181-4|LNC|Cells counted.total|Cells counted.total
C2970610|T201|COMP|61182-2|LNC|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C2970611|T201|COMP|61183-0|LNC|Cells.myeloperoxidase/100 cells|Cells.myeloperoxidase/100 cells
C2970612|T201|COMP|61184-8|LNC|Spermatozoa.broken tail/100 spermatozoa|Spermatozoa.broken tail/100 spermatozoa
C2970614|T201|COMP|61185-5|LNC|Spermatozoa.thick midpiece/100 spermatozoa|Spermatozoa.thick midpiece/100 spermatozoa
C2970616|T201|COMP|61186-3|LNC|Spermatozoa.thin midpiece/100 spermatozoa|Spermatozoa.thin midpiece/100 spermatozoa
C2970618|T201|COMP|61187-1|LNC|Spermatozoa.bent midpiece/100 spermatozoa|Spermatozoa.bent midpiece/100 spermatozoa
C2970620|T201|COMP|61189-7|LNC|Coagulation tissue factor induced.INR|Coagulation tissue factor induced.INR
C2970621|T201|COMP|61190-5|LNC|Coagulation tissue factor induced|Coagulation tissue factor induced
C2970622|T201|COMP|61191-3|LNC|Coagulation surface induced|Coagulation surface induced
C2970623|T201|COMP|61192-1|LNC|Color|Color
C2970624|T201|COMP|61193-9|LNC|Clarity|Clarity
C2970625|T201|COMP|61194-7|LNC|Cells counted.total|Cells counted.total
C2970626|T201|COMP|61195-4|LNC|Albumin|Albumin
C2970627|T201|COMP|61196-2|LNC|Albumin|Albumin
C2970628|T201|COMP|61197-0|LNC|oxyCODONE+Oxymorphone|oxyCODONE+Oxymorphone
C2970629|T201|COMP|61198-8|LNC|Raltegravir|Raltegravir
C2970630|T201|COMP|61199-6|LNC|HIV 1 integrase gene mutations detected|HIV 1 integrase gene mutations detected
C2970632|T201|COMP|61200-2|LNC|Colorado tick fever virus Ab.IgG|Colorado tick fever virus Ab.IgG
C2970637|T201|COMP|61205-1|LNC|Acer macrophyllum Ab.IgE/IgE.total|Acer macrophyllum Ab.IgE/IgE.total
C2970638|T201|COMP|61206-9|LNC|Acer negundo Ab.IgE/IgE.total|Acer negundo Ab.IgE/IgE.total
C2970639|T201|COMP|61207-7|LNC|Acremonium sp Ab.IgE/IgE.total|Acremonium sp Ab.IgE/IgE.total
C2970640|T201|COMP|61208-5|LNC|Aedes communis Ab.IgE/IgE.total|Aedes communis Ab.IgE/IgE.total
C2970641|T201|COMP|61209-3|LNC|Agaricus hortensis Ab.IgE/IgE.total|Agaricus hortensis Ab.IgE/IgE.total
C2970642|T201|COMP|61210-1|LNC|Allium cepa Ab.IgE/IgE.total|Allium cepa Ab.IgE/IgE.total
C2970643|T201|COMP|61211-9|LNC|Allium sativum Ab.IgE/IgE.total|Allium sativum Ab.IgE/IgE.total
C2970644|T201|COMP|61212-7|LNC|Alnus incana Ab.IgE/IgE.total|Alnus incana Ab.IgE/IgE.total
C2970645|T201|COMP|61213-5|LNC|Lactalbumin alpha Ab.IgE/IgE.total|Lactalbumin alpha Ab.IgE/IgE.total
C2970646|T201|COMP|61214-3|LNC|Ambrosia elatior Ab.IgE/IgE.total|Ambrosia elatior Ab.IgE/IgE.total
C2970647|T201|COMP|61215-0|LNC|Ambrosia trifida Ab.IgE/IgE.total|Ambrosia trifida Ab.IgE/IgE.total
C2970648|T201|COMP|61216-8|LNC|Ananas comosus Ab.IgE/IgE.total|Ananas comosus Ab.IgE/IgE.total
C2970649|T201|COMP|61217-6|LNC|Anthoxanthum odoratum Ab.IgE/IgE.total|Anthoxanthum odoratum Ab.IgE/IgE.total
C2970650|T201|COMP|61218-4|LNC|Apium graveolens Ab.IgE/IgE.total|Apium graveolens Ab.IgE/IgE.total
C2970651|T201|COMP|61219-2|LNC|Arachis hypogaea Ab.IgE/IgE.total|Arachis hypogaea Ab.IgE/IgE.total
C2970652|T201|COMP|61220-0|LNC|Ascaris sp Ab.IgE/IgE.total|Ascaris sp Ab.IgE/IgE.total
C2970653|T201|COMP|61221-8|LNC|Aspergillus niger Ab.IgE/IgE.total|Aspergillus niger Ab.IgE/IgE.total
C2970654|T201|COMP|61222-6|LNC|Aspergillus sp Ab.IgE/IgE.total|Aspergillus sp Ab.IgE/IgE.total
C2970655|T201|COMP|61223-4|LNC|Astacus astacus Ab.IgE/IgE.total|Astacus astacus Ab.IgE/IgE.total
C2970656|T201|COMP|61224-2|LNC|Atriplex lentiformis Ab.IgE/IgE.total|Atriplex lentiformis Ab.IgE/IgE.total
C2970657|T201|COMP|61225-9|LNC|Aureobasidium pullulans Ab.IgE/IgE.total|Aureobasidium pullulans Ab.IgE/IgE.total
C2970658|T201|COMP|61226-7|LNC|Avena sativa Ab.IgE/IgE.total|Avena sativa Ab.IgE/IgE.total
C2970659|T201|COMP|61227-5|LNC|Betula populifolia Ab.IgE/IgE.total|Betula populifolia Ab.IgE/IgE.total
C2970660|T201|COMP|61228-3|LNC|Betula verrucosa Ab.IgE/IgE.total|Betula verrucosa Ab.IgE/IgE.total
C2970662|T201|COMP|61230-9|LNC|Blatella germanica Ab.IgE/IgE.total|Blatella germanica Ab.IgE/IgE.total
C2970663|T201|COMP|61231-7|LNC|Botrytis cinerea Ab.IgE/IgE.total|Botrytis cinerea Ab.IgE/IgE.total
C2970664|T201|COMP|61232-5|LNC|Brassica oleracea var botrytis Ab.IgE/IgE.total|Brassica oleracea var botrytis Ab.IgE/IgE.total
C2970665|T201|COMP|61233-3|LNC|Brassica oleracea var capitata Ab.IgE/IgE.total|Brassica oleracea var capitata Ab.IgE/IgE.total
C2970666|T201|COMP|61234-1|LNC|Brassica oleracea var italica Ab.IgE/IgE.total|Brassica oleracea var italica Ab.IgE/IgE.total
C2970667|T201|COMP|61235-8|LNC|Bromus inermis Ab.IgE/IgE.total|Bromus inermis Ab.IgE/IgE.total
C2970668|T201|COMP|61236-6|LNC|Budgerigar droppings Ab.IgE/IgE.total|Budgerigar droppings Ab.IgE/IgE.total
C2970669|T201|COMP|61237-4|LNC|Budgerigar feather Ab.IgE/IgE.total|Budgerigar feather Ab.IgE/IgE.total
C2970670|T201|COMP|61238-2|LNC|Candida albicans Ab.IgE/IgE.total|Candida albicans Ab.IgE/IgE.total
C2970671|T201|COMP|61239-0|LNC|Capsicum annuum Ab.IgE/IgE.total|Capsicum annuum Ab.IgE/IgE.total
C2970672|T201|COMP|61240-8|LNC|Carya illinoinensis tree Ab.IgE/IgE.total|Carya illinoinensis tree Ab.IgE/IgE.total
C2970673|T201|COMP|61241-6|LNC|Casein Ab.IgE/IgE.total|Casein Ab.IgE/IgE.total
C2970674|T201|COMP|61242-4|LNC|Chaetomium globosum Ab.IgE/IgE.total|Chaetomium globosum Ab.IgE/IgE.total
C2970675|T201|COMP|61243-2|LNC|Chenopodium album Ab.IgE/IgE.total|Chenopodium album Ab.IgE/IgE.total
C2970676|T201|COMP|61244-0|LNC|Cicer arietinus Ab.IgE/IgE.total|Cicer arietinus Ab.IgE/IgE.total
C2970677|T201|COMP|61245-7|LNC|Cinnamomum spp Ab.IgE/IgE.total|Cinnamomum spp Ab.IgE/IgE.total
C2970678|T201|COMP|61246-5|LNC|Citrus limon Ab.IgE/IgE.total|Citrus limon Ab.IgE/IgE.total
C2970679|T201|COMP|61247-3|LNC|Citrus paradisis Ab.IgE/IgE.total|Citrus paradisis Ab.IgE/IgE.total
C2970680|T201|COMP|61248-1|LNC|Citrus sinensis Ab.IgE/IgE.total|Citrus sinensis Ab.IgE/IgE.total
C2970681|T201|COMP|61249-9|LNC|Cladosporium herbarum Ab.IgE/IgE.total|Cladosporium herbarum Ab.IgE/IgE.total
C2970682|T201|COMP|61250-7|LNC|Coffea spp Ab.IgE/IgE.total|Coffea spp Ab.IgE/IgE.total
C2970683|T201|COMP|61251-5|LNC|Cryptomeria japonica Ab.IgE/IgE.total|Cryptomeria japonica Ab.IgE/IgE.total
C2970684|T201|COMP|61276-2|LNC|Insulin porcine Ab.IgE/IgE.total|Insulin porcine Ab.IgE/IgE.total
C2972886|T201|COMP|61277-0|LNC|Hexamethylene diisocyanate (HDI) Ab.IgE/IgE.total|Hexamethylene diisocyanate (HDI) Ab.IgE/IgE.total
C2972887|T201|COMP|61278-8|LNC|Toluene diisocyanate (TDI) Ab.IgE/IgE.total|Toluene diisocyanate (TDI) Ab.IgE/IgE.total
C2972888|T201|COMP|61279-6|LNC|Juglans regia Ab.IgE/IgE.total|Juglans regia Ab.IgE/IgE.total
C2972889|T201|COMP|61280-4|LNC|Lactuca sativa Ab.IgE/IgE.total|Lactuca sativa Ab.IgE/IgE.total
C2972890|T201|COMP|61281-2|LNC|Loligo sp Ab.IgE/IgE.total|Loligo sp Ab.IgE/IgE.total
C2972891|T201|COMP|61282-0|LNC|Lolium perenne Ab.IgE/IgE.total|Lolium perenne Ab.IgE/IgE.total
C2972892|T201|COMP|61283-8|LNC|Macadamia spp Ab.IgE/IgE.total|Macadamia spp Ab.IgE/IgE.total
C2972893|T201|COMP|61284-6|LNC|Melaleuca leucadendron Ab.IgE/IgE.total|Melaleuca leucadendron Ab.IgE/IgE.total
C2972894|T201|COMP|61285-3|LNC|Micropterus salmoides Ab.IgE/IgE.total|Micropterus salmoides Ab.IgE/IgE.total
C2972895|T201|COMP|61286-1|LNC|Morus alba Ab.IgE/IgE.total|Morus alba Ab.IgE/IgE.total
C2972896|T201|COMP|61287-9|LNC|Musa spp Ab.IgE/IgE.total|Musa spp Ab.IgE/IgE.total
C2972897|T201|COMP|61288-7|LNC|Ocimum basilicum Ab.IgE/IgE.total|Ocimum basilicum Ab.IgE/IgE.total
C2972898|T201|COMP|61289-5|LNC|Oncorhynchus mykiss Ab.IgE/IgE.total|Oncorhynchus mykiss Ab.IgE/IgE.total
C2972899|T201|COMP|61290-3|LNC|Origanum vulgare Ab.IgE/IgE.total|Origanum vulgare Ab.IgE/IgE.total
C2972900|T201|COMP|61291-1|LNC|Oryza sativa Ab.IgE/IgE.total|Oryza sativa Ab.IgE/IgE.total
C2972901|T201|COMP|61292-9|LNC|Ostrea edulis Ab.IgE/IgE.total|Ostrea edulis Ab.IgE/IgE.total
C2972902|T201|COMP|61293-7|LNC|Passiflora edulis Ab.IgE/IgE.total|Passiflora edulis Ab.IgE/IgE.total
C2972903|T201|COMP|61294-5|LNC|Persea americana Ab.IgE/IgE.total|Persea americana Ab.IgE/IgE.total
C2972904|T201|COMP|61295-2|LNC|Petroselinum crispum Ab.IgE/IgE.total|Petroselinum crispum Ab.IgE/IgE.total
C2972905|T201|COMP|61296-0|LNC|Phleum pratense Ab.IgE/IgE.total|Phleum pratense Ab.IgE/IgE.total
C2972906|T201|COMP|61297-8|LNC|Phthalic anhydride Ab.IgE/IgE.total|Phthalic anhydride Ab.IgE/IgE.total
C2972907|T201|COMP|61306-7|LNC|Prunus avium Ab.IgE/IgE.total|Prunus avium Ab.IgE/IgE.total
C2972908|T201|COMP|61307-5|LNC|Pyrus communis Ab.IgE/IgE.total|Pyrus communis Ab.IgE/IgE.total
C2972909|T201|COMP|61308-3|LNC|Rhizopus nigricans Ab.IgE/IgE.total|Rhizopus nigricans Ab.IgE/IgE.total
C2972910|T201|COMP|61309-1|LNC|Rumex acetosella Ab.IgE/IgE.total|Rumex acetosella Ab.IgE/IgE.total
C2972911|T201|COMP|61310-9|LNC|Salix caprea Ab.IgE/IgE.total|Salix caprea Ab.IgE/IgE.total
C2972912|T201|COMP|61311-7|LNC|Salsola kali Ab.IgE/IgE.total|Salsola kali Ab.IgE/IgE.total
C2972913|T201|COMP|61312-5|LNC|Secale cereale Ab.IgE/IgE.total|Secale cereale Ab.IgE/IgE.total
C2972914|T201|COMP|61313-3|LNC|Sesamum indicum Ab.IgE/IgE.total|Sesamum indicum Ab.IgE/IgE.total
C2972915|T201|COMP|61314-1|LNC|Sheep wool Ab.IgE/IgE.total|Sheep wool Ab.IgE/IgE.total
C2972916|T201|COMP|61315-8|LNC|Solenopsis invicta Ab.IgE/IgE.total|Solenopsis invicta Ab.IgE/IgE.total
C2972917|T201|COMP|61316-6|LNC|Solidago virgaurea Ab.IgE/IgE.total|Solidago virgaurea Ab.IgE/IgE.total
C2972918|T201|COMP|61317-4|LNC|Spinacia oleracea Ab.IgE/IgE.total|Spinacia oleracea Ab.IgE/IgE.total
C2972919|T201|COMP|61318-2|LNC|Taraxacum vulgare Ab.IgE/IgE.total|Taraxacum vulgare Ab.IgE/IgE.total
C2972920|T201|COMP|61319-0|LNC|Theobroma cacao Ab.IgE/IgE.total|Theobroma cacao Ab.IgE/IgE.total
C2972921|T201|COMP|61320-8|LNC|Trachurus japonicus Ab.IgE/IgE.total|Trachurus japonicus Ab.IgE/IgE.total
C2972922|T201|COMP|61321-6|LNC|Trimellitic anhydride Ab.IgE/IgE.total|Trimellitic anhydride Ab.IgE/IgE.total
C2972923|T201|COMP|61322-4|LNC|Ulmus americana Ab.IgE/IgE.total|Ulmus americana Ab.IgE/IgE.total
C2972924|T201|COMP|61323-2|LNC|Vaccinium oxycoccos Ab.IgE/IgE.total|Vaccinium oxycoccos Ab.IgE/IgE.total
C2972925|T201|COMP|61324-0|LNC|Vanilla planifolia Ab.IgE/IgE.total|Vanilla planifolia Ab.IgE/IgE.total
C2972926|T201|COMP|61325-7|LNC|Vespa crabro Ab.IgE/IgE.total|Vespa crabro Ab.IgE/IgE.total
C2972927|T201|COMP|61326-5|LNC|Xanthium commune Ab.IgE/IgE.total|Xanthium commune Ab.IgE/IgE.total
C2972928|T201|COMP|61327-3|LNC|Zea mays Ab.IgE/IgE.total|Zea mays Ab.IgE/IgE.total
C2972929|T201|COMP|61328-1|LNC|Zingiber officinale Ab.IgE/IgE.total|Zingiber officinale Ab.IgE/IgE.total
C2972930|T201|COMP|61329-9|LNC|Cucumis sativus Ab.IgE/IgE.total|Cucumis sativus Ab.IgE/IgE.total
C2972931|T201|COMP|61330-7|LNC|Pinus edulis Ab.IgE/IgE.total|Pinus edulis Ab.IgE/IgE.total
C2972932|T201|COMP|61331-5|LNC|Beef Ab.IgE/IgE.total|Beef Ab.IgE/IgE.total
C2972933|T201|COMP|61332-3|LNC|Cow milk Ab.IgE/IgE.total|Cow milk Ab.IgE/IgE.total
C2972934|T201|COMP|61333-1|LNC|Dog dander Ab.IgE/IgE.total|Dog dander Ab.IgE/IgE.total
C2972935|T201|COMP|61334-9|LNC|Dog epithelium Ab.IgE/IgE.total|Dog epithelium Ab.IgE/IgE.total
C2972936|T201|COMP|61335-6|LNC|Goat milk Ab.IgE/IgE.total|Goat milk Ab.IgE/IgE.total
C2972937|T201|COMP|61336-4|LNC|Cochineal extract Ab.IgE/IgE.total|Cochineal extract Ab.IgE/IgE.total
C2972938|T201|COMP|61337-2|LNC|Chicken feather Ab.IgE/IgE.total|Chicken feather Ab.IgE/IgE.total
C2972939|T201|COMP|61338-0|LNC|Egg white Ab.IgE/IgE.total|Egg white Ab.IgE/IgE.total
C2972940|T201|COMP|61339-8|LNC|Egg yolk Ab.IgE/IgE.total|Egg yolk Ab.IgE/IgE.total
C2972941|T201|COMP|61340-6|LNC|Cottonseed Ab.IgE/IgE.total|Cottonseed Ab.IgE/IgE.total
C2972942|T201|COMP|61341-4|LNC|Gerbil epithelium Ab.IgE/IgE.total|Gerbil epithelium Ab.IgE/IgE.total
C2972943|T201|COMP|61342-2|LNC|Mouse urine proteins Ab.IgE/IgE.total|Mouse urine proteins Ab.IgE/IgE.total
C2972944|T201|COMP|61343-0|LNC|Ferret epithelium Ab.IgE/IgE.total|Ferret epithelium Ab.IgE/IgE.total
C2972945|T201|COMP|61344-8|LNC|Sheep epithelium Ab.IgE/IgE.total|Sheep epithelium Ab.IgE/IgE.total
C2972946|T201|COMP|61345-5|LNC|Flounder Ab.IgE/IgE.total|Flounder Ab.IgE/IgE.total
C2972947|T201|COMP|61346-3|LNC|Rat urine proteins Ab.IgE/IgE.total|Rat urine proteins Ab.IgE/IgE.total
C2972948|T201|COMP|61347-1|LNC|Pork Ab.IgE/IgE.total|Pork Ab.IgE/IgE.total
C2972949|T201|COMP|61348-9|LNC|Cockatiel droppings Ab.IgE/IgE.total|Cockatiel droppings Ab.IgE/IgE.total
C2972950|T201|COMP|61349-7|LNC|Cockatiel feather Ab.IgE/IgE.total|Cockatiel feather Ab.IgE/IgE.total
C2972956|T201|COMP|61355-4|LNC|Capreomycin 5.0 ug/mL|Capreomycin 5.0 ug/mL
C2972962|T201|COMP|61360-4|LNC|Acinetobacter baumannii DNA|Acinetobacter baumannii DNA
C2972963|T201|COMP|61361-2|LNC|Klebsiella aerogenes DNA|Klebsiella aerogenes DNA
C2972964|T201|COMP|61362-0|LNC|Enterococcus faecalis DNA|Enterococcus faecalis DNA
C2972965|T201|COMP|61363-8|LNC|Adenovirus 3+4+7+21 DNA|Adenovirus 3+4+7+21 DNA
C2972966|T201|COMP|61364-6|LNC|Echovirus+Coxsackievirus RNA|Echovirus+Coxsackievirus RNA
C2972967|T201|COMP|61365-3|LNC|Parainfluenza virus RNA|Parainfluenza virus RNA
C2972968|T201|COMP|61366-1|LNC|Haemophilus influenzae DNA|Haemophilus influenzae DNA
C2972969|T201|COMP|61367-9|LNC|Clostridioides difficile DNA|Clostridioides difficile DNA
C2972970|T201|COMP|61368-7|LNC|Campylobacter jejuni DNA|Campylobacter jejuni DNA
C2972971|T201|COMP|61369-5|LNC|Listeria monocytogenes DNA|Listeria monocytogenes DNA
C2972972|T201|COMP|61370-3|LNC|Salmonella enterica DNA|Salmonella enterica DNA
C2972973|T201|COMP|61371-1|LNC|Vibrio cholerae DNA|Vibrio cholerae DNA
C2972974|T201|COMP|61372-9|LNC|Human papilloma virus 16 DNA|Human papilloma virus 16 DNA
C2972975|T201|COMP|61373-7|LNC|Human papilloma virus 18 DNA|Human papilloma virus 18 DNA
C2972976|T201|COMP|61374-5|LNC|Human papilloma virus 26 DNA|Human papilloma virus 26 DNA
C2972977|T201|COMP|61375-2|LNC|Human papilloma virus 31 DNA|Human papilloma virus 31 DNA
C2972978|T201|COMP|61376-0|LNC|Human papilloma virus 33 DNA|Human papilloma virus 33 DNA
C2972979|T201|COMP|61377-8|LNC|Human papilloma virus 35 DNA|Human papilloma virus 35 DNA
C2972980|T201|COMP|61378-6|LNC|Human papilloma virus 39 DNA|Human papilloma virus 39 DNA
C2972981|T201|COMP|61379-4|LNC|Human papilloma virus 44 DNA|Human papilloma virus 44 DNA
C2972982|T201|COMP|61380-2|LNC|Human papilloma virus 45 DNA|Human papilloma virus 45 DNA
C2972983|T201|COMP|61381-0|LNC|Human papilloma virus 51 DNA|Human papilloma virus 51 DNA
C2972984|T201|COMP|61382-8|LNC|Human papilloma virus 52 DNA|Human papilloma virus 52 DNA
C2972985|T201|COMP|61383-6|LNC|Human papilloma virus 53 DNA|Human papilloma virus 53 DNA
C2972986|T201|COMP|61384-4|LNC|Human papilloma virus 58 DNA|Human papilloma virus 58 DNA
C2972987|T201|COMP|61385-1|LNC|Human papilloma virus 59 DNA|Human papilloma virus 59 DNA
C2972988|T201|COMP|61386-9|LNC|Human papilloma virus 66 DNA|Human papilloma virus 66 DNA
C2972989|T201|COMP|61387-7|LNC|Human papilloma virus 67 DNA|Human papilloma virus 67 DNA
C2972990|T201|COMP|61388-5|LNC|Human papilloma virus 68 DNA|Human papilloma virus 68 DNA
C2972991|T201|COMP|61389-3|LNC|Human papilloma virus 69 DNA|Human papilloma virus 69 DNA
C2972992|T201|COMP|61390-1|LNC|Human papilloma virus 70 DNA|Human papilloma virus 70 DNA
C2972993|T201|COMP|61391-9|LNC|Human papilloma virus 73 DNA|Human papilloma virus 73 DNA
C2972994|T201|COMP|61392-7|LNC|Human papilloma virus 82 DNA|Human papilloma virus 82 DNA
C2972995|T201|COMP|61400-8|LNC|Proteus mirabilis DNA|Proteus mirabilis DNA
C2972996|T201|COMP|61401-6|LNC|Pseudomonas aeruginosa DNA|Pseudomonas aeruginosa DNA
C2972997|T201|COMP|61402-4|LNC|Serratia marcescens DNA|Serratia marcescens DNA
C2972998|T201|COMP|61403-2|LNC|Stenotrophomonas maltophilia DNA|Stenotrophomonas maltophilia DNA
C2972999|T201|COMP|61404-0|LNC|Staphylococcus aureus DNA|Staphylococcus aureus DNA
C2973000|T201|COMP|61405-7|LNC|Staphylococcus epidermidis DNA|Staphylococcus epidermidis DNA
C2973001|T201|COMP|61406-5|LNC|XXX blood group Ab|XXX blood group Ab
C2973002|T201|COMP|61409-9|LNC|Cyclobenzaprine|Cyclobenzaprine
C2973003|T201|COMP|61410-7|LNC|Cyclobenzaprine|Cyclobenzaprine
C2973004|T201|COMP|61412-3|LNC|Desipramine|Desipramine
C2973005|T201|COMP|61413-1|LNC|Desipramine|Desipramine
C2973006|T201|COMP|61415-6|LNC|Doxepin|Doxepin
C2973007|T201|COMP|61416-4|LNC|Doxepin|Doxepin
C2973008|T201|COMP|61418-0|LNC|Imipramine|Imipramine
C2973009|T201|COMP|61419-8|LNC|Imipramine|Imipramine
C2973010|T201|COMP|61421-4|LNC|Norhydrocodone|Norhydrocodone
C2973011|T201|COMP|61422-2|LNC|Norhydrocodone|Norhydrocodone
C2973012|T201|COMP|61424-8|LNC|Noroxycodone|Noroxycodone
C2973013|T201|COMP|61425-5|LNC|Noroxycodone|Noroxycodone
C2973014|T201|COMP|61427-1|LNC|Nortriptyline|Nortriptyline
C2973015|T201|COMP|61428-9|LNC|Nortriptyline|Nortriptyline
C2973016|T201|COMP|61430-5|LNC|Aquaporin 4 water channel Ab|Aquaporin 4 water channel Ab
C2973146|T201|COMP|62321-5|LNC|Severe combined immunodeficiency|Severe combined immunodeficiency
C2973155|T201|COMP|62342-1|LNC|Borrelia burgdorferi Ab.IgG & IgM|Borrelia burgdorferi Ab.IgG & IgM
C2973156|T201|COMP|62234-0|LNC|Albumin|Albumin
C2973157|T201|COMP|62235-7|LNC|Albumin|Albumin
C2973158|T201|COMP|62236-5|LNC|Pyridoxal phosphate|Pyridoxal phosphate
C2973159|T201|COMP|62237-3|LNC|Carbapenem|Carbapenem
C2973160|T201|COMP|62238-1|LNC|Glomerular filtration rate/1.73 sq M.predicted|Glomerular filtration rate/1.73 sq M.predicted
C2973161|T201|COMP|62239-9|LNC|Leukocytes|Leukocytes
C2973162|T201|COMP|62240-7|LNC|Erythrocytes|Erythrocytes
C2973163|T201|COMP|62241-5|LNC|Hematocrit|Hematocrit
C2973164|T201|COMP|62242-3|LNC|Erythrocyte mean corpuscular volume|Erythrocyte mean corpuscular volume
C2973165|T201|COMP|62243-1|LNC|Erythrocyte mean corpuscular hemoglobin|Erythrocyte mean corpuscular hemoglobin
C2973166|T201|COMP|62244-9|LNC|Platelets|Platelets
C2973167|T201|COMP|62245-6|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C2973169|T201|COMP|62247-2|LNC|Erythrocyte distribution width|Erythrocyte distribution width
C2973170|T201|COMP|62248-0|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C2973171|T201|COMP|62249-8|LNC|Reticulocytes|Reticulocytes
C2973172|T201|COMP|62250-6|LNC|Reticulocytes.immature/Reticulocytes.total|Reticulocytes.immature/Reticulocytes.total
C2973173|T201|COMP|62251-4|LNC|Leukocytes|Leukocytes
C2973174|T201|COMP|62252-2|LNC|Cells.CD79/100 cells|Cells.CD79/100 cells
C2973175|T201|COMP|62253-0|LNC|Lipoprotein.alpha|Lipoprotein.alpha
C2973176|T201|COMP|62254-8|LNC|Lipoprotein.pre-beta|Lipoprotein.pre-beta
C2973177|T201|COMP|62255-5|LNC|Lipoprotein insulin resistance score|Lipoprotein insulin resistance score
C2973178|T201|COMP|62256-3|LNC|Bacterial aminoglycoside resistance aacA gene|Bacterial aminoglycoside resistance aacA gene
C2973179|T201|COMP|62257-1|LNC|Cephalosporin resistance gene|Cephalosporin resistance gene
C2973181|T201|COMP|62259-7|LNC|Methicillin resistance gene|Methicillin resistance gene
C2973182|T201|COMP|62260-5|LNC|Bacterial tetracycline resistance tetK+tetM genes|Bacterial tetracycline resistance tetK+tetM genes
C2973183|T201|COMP|62261-3|LNC|Bacterial vancomycin resistance vanA+vanB genes|Bacterial vancomycin resistance vanA+vanB genes
C2973199|T201|COMP|62290-2|LNC|1,25-Dihydroxyvitamin D|1,25-Dihydroxyvitamin D
C2973200|T201|COMP|62291-0|LNC|1,25-Dihydroxyvitamin D2|1,25-Dihydroxyvitamin D2
C2973201|T201|COMP|62292-8|LNC|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3
C2973210|T201|COMP|62301-7|LNC|Lysosomal storage disorders|Lysosomal storage disorders
C2973211|T201|COMP|62302-5|LNC|Lysosomal storage disorders suspected|Lysosomal storage disorders suspected
C2973213|T201|COMP|62304-1|LNC|Fabry disease newborn screening panel|Fabry disease newborn screening panel
C2973214|T201|COMP|62305-8|LNC|Fabry disease|Fabry disease
C2973216|T201|COMP|62307-4|LNC|Krabbe disease newborn screening panel|Krabbe disease newborn screening panel
C2973217|T201|COMP|62308-2|LNC|Krabbe disease|Krabbe disease
C2973219|T201|COMP|62310-8|LNC|Galactosylceramidase|Galactosylceramidase
C2973220|T201|COMP|62311-6|LNC|Gaucher disease newborn screening panel|Gaucher disease newborn screening panel
C2973221|T201|COMP|62312-4|LNC|Gaucher disease|Gaucher disease
C2973223|T201|COMP|62315-7|LNC|Niemann Pick disease A+B newborn screening panel|Niemann Pick disease A+B newborn screening panel
C2973224|T201|COMP|62316-5|LNC|Acid sphingomyelinase|Acid sphingomyelinase
C2973226|T201|COMP|62318-1|LNC|Niemann Pick disease A+B|Niemann Pick disease A+B
C2973228|T201|COMP|62320-7|LNC|T-cell receptor excision circle|T-cell receptor excision circle
C2973229|T201|COMP|62343-9|LNC|Chromosome analysis copy number change panel|Chromosome analysis copy number change panel
C2973230|T201|COMP|62344-7|LNC|Chromosome analysis.metaphase panel|Chromosome analysis.metaphase panel
C2973231|T201|COMP|62345-4|LNC|Chromosome analysis.interphase panel|Chromosome analysis.interphase panel
C2973232|T201|COMP|62346-2|LNC|Chromosome analysis.interphase panel|Chromosome analysis.interphase panel
C2973233|T201|COMP|62347-0|LNC|Chromosome analysis.prenatal panel|Chromosome analysis.prenatal panel
C2973234|T201|COMP|62348-8|LNC|Chromosome analysis panel|Chromosome analysis panel
C2973235|T201|COMP|62349-6|LNC|Chromosome analysis panel|Chromosome analysis panel
C2973236|T201|COMP|62350-4|LNC|Chromosome analysis panel|Chromosome analysis panel
C2973237|T201|COMP|62351-2|LNC|Chromosome analysis panel|Chromosome analysis panel
C2973238|T201|COMP|62352-0|LNC|Chromosome analysis panel|Chromosome analysis panel
C2973239|T201|COMP|62353-8|LNC|Chromosome analysis panel|Chromosome analysis panel
C2973240|T201|COMP|62354-6|LNC|Chromosome analysis.metaphase panel|Chromosome analysis.metaphase panel
C2973241|T201|COMP|62355-3|LNC|Chromosome analysis panel|Chromosome analysis panel
C2973242|T201|COMP|62356-1|LNC|Chromosome analysis result in ISCN expression|Chromosome analysis result in ISCN expression
C2973243|T201|COMP|62357-9|LNC|Chromosome analysis overall interpretation|Chromosome analysis overall interpretation
C2973244|T201|COMP|62358-7|LNC|ISCN band level|ISCN band level
C2973245|T201|COMP|62359-5|LNC|Chromosome banding method|Chromosome banding method
C2973246|T201|COMP|62367-8|LNC|Chromosome analysis panel|Chromosome analysis panel
C2973247|T201|COMP|62368-6|LNC|Cell phase|Cell phase
C2973248|T201|COMP|62369-4|LNC|FISH probe name panel|FISH probe name panel
C2973249|T201|COMP|62370-2|LNC|FISH probe gene name|FISH probe gene name
C2973250|T201|COMP|62371-0|LNC|FISH probe locus|FISH probe locus
C2973251|T201|COMP|62372-8|LNC|FISH probe vendor|FISH probe vendor
C2973252|T201|COMP|62373-6|LNC|Human reference assembly release, UCSC version|Human reference assembly release, UCSC version
C2973253|T201|COMP|62374-4|LNC|Human reference sequence assembly release number|Human reference sequence assembly release number
C2973254|T201|COMP|62375-1|LNC|Microarray platform|Microarray platform
C2973255|T201|COMP|62376-9|LNC|Microarray platform version number|Microarray platform version number
C2973256|T201|COMP|62377-7|LNC|Chromosome copy number change panel|Chromosome copy number change panel
C2973257|T201|COMP|62378-5|LNC|Chromosome copy number change|Chromosome copy number change
C2973258|T201|COMP|62379-3|LNC|Chromosome band involved start|Chromosome band involved start
C2973259|T201|COMP|62380-1|LNC|Chromosome band involved end|Chromosome band involved end
C2973260|T201|COMP|62381-9|LNC|Base pair start coordinate|Base pair start coordinate
C2973261|T201|COMP|62382-7|LNC|Base pair end coordinate|Base pair end coordinate
C2973262|T201|COMP|62383-5|LNC|Flanking normal region before start|Flanking normal region before start
C2973263|T201|COMP|62384-3|LNC|Flanking normal region after end|Flanking normal region after end
C2973264|T201|COMP|62385-0|LNC|Recommendation|Recommendation
C2973265|T201|COMP|62386-8|LNC|Chromosome analysis summary panel|Chromosome analysis summary panel
C2973266|T201|COMP|62388-4|LNC|Hemoglobin A1c/Hemoglobin.total|Hemoglobin A1c/Hemoglobin.total
C2973267|T201|COMP|62389-2|LNC|Chromosome analysis master panel|Chromosome analysis master panel
C2973277|T201|COMP|10330-9|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C2973278|T201|COMP|10329-1|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C2973279|T201|COMP|32503-5|LNC|Cells.CD13+CD33+/100 cells|Cells.CD13+CD33+/100 cells
C2973280|T201|COMP|26572-8|LNC|Cells.CD2+CD7+/100 cells|Cells.CD2+CD7+/100 cells
C2973281|T201|COMP|17097-7|LNC|Cells.CD10+CD20+/100 cells|Cells.CD10+CD20+/100 cells
C2973283|T201|COMP|8104-2|LNC|Cells.CD5+CD20+/100 cells|Cells.CD5+CD20+/100 cells
C3166946|T201|COMP|57645-4|LNC|C peptide^10M pre XXX challenge|C peptide^10M pre XXX challenge
C3167211|T201|COMP|57593-6|LNC|Aldosterone^30M pre XXX challenge|Aldosterone^30M pre XXX challenge
C3167212|T201|COMP|57594-4|LNC|Aldosterone^30M pre XXX challenge|Aldosterone^30M pre XXX challenge
C3167213|T201|COMP|57648-8|LNC|C peptide^5M pre XXX challenge|C peptide^5M pre XXX challenge
C3167214|T201|COMP|57649-6|LNC|C peptide^1H pre XXX challenge|C peptide^1H pre XXX challenge
C3167215|T201|COMP|57650-4|LNC|C peptide^70M pre XXX challenge|C peptide^70M pre XXX challenge
C3167216|T201|COMP|57795-7|LNC|Fecal hydrolysis panel|Fecal hydrolysis panel
C3167217|T201|COMP|57836-9|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C3167218|T201|COMP|57840-1|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C3167219|T201|COMP|57850-0|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C3167221|T201|COMP|58472-2|LNC|Other cells|Other cells
C3167817|T201|COMP|58904-4|LNC|Nucleated cells|Nucleated cells
C3167818|T201|COMP|58905-1|LNC|Nucleated cells|Nucleated cells
C3167819|T201|COMP|58906-9|LNC|Nucleated cells|Nucleated cells
C3167822|T201|COMP|60841-4|LNC|Oxygen content|Oxygen content
C3167827|T201|COMP|59246-9|LNC|Palmitoyl protein thioesterase|Palmitoyl protein thioesterase
C3167828|T201|COMP|59586-8|LNC|HLA Ab.IgG|HLA Ab.IgG
C3168375|T201|COMP|60519-6|LNC|Fatty acids.ethyl esters|Fatty acids.ethyl esters
C3168378|T201|COMP|60678-0|LNC|Protein/Creatinine|Protein/Creatinine
C3168379|T201|COMP|61154-1|LNC|Hepatitis B virus codon L180M|Hepatitis B virus codon L180M
C3168380|T201|COMP|61155-8|LNC|Hepatitis B virus codon L80V|Hepatitis B virus codon L80V
C3168381|T201|COMP|61156-6|LNC|Hepatitis B virus codon V173L|Hepatitis B virus codon V173L
C3168382|T201|COMP|61157-4|LNC|Hepatitis B virus codon M204V|Hepatitis B virus codon M204V
C3168383|T201|COMP|61158-2|LNC|Hepatitis B virus codon M204I|Hepatitis B virus codon M204I
C3168384|T201|COMP|61159-0|LNC|Hepatitis B virus codon M204S|Hepatitis B virus codon M204S
C3168385|T201|COMP|61160-8|LNC|Hepatitis B virus codon A181V|Hepatitis B virus codon A181V
C3168386|T201|COMP|61161-6|LNC|Hepatitis B virus codon A181T|Hepatitis B virus codon A181T
C3168387|T201|COMP|61162-4|LNC|Hepatitis B virus codon N236T|Hepatitis B virus codon N236T
C3168388|T201|COMP|61163-2|LNC|Hepatitis B virus codon A194T|Hepatitis B virus codon A194T
C3168389|T201|COMP|61164-0|LNC|Hepatitis B virus codon T184S|Hepatitis B virus codon T184S
C3168390|T201|COMP|61165-7|LNC|Hepatitis B virus codon T184I|Hepatitis B virus codon T184I
C3168391|T201|COMP|61166-5|LNC|Hepatitis B virus codon S202G|Hepatitis B virus codon S202G
C3168392|T201|COMP|61167-3|LNC|Hepatitis B virus codon S202C|Hepatitis B virus codon S202C
C3168393|T201|COMP|61168-1|LNC|Hepatitis B virus codon S202I|Hepatitis B virus codon S202I
C3168394|T201|COMP|61169-9|LNC|Hepatitis B virus codon I233V|Hepatitis B virus codon I233V
C3168395|T201|COMP|61170-7|LNC|Hepatitis B virus codon M250V|Hepatitis B virus codon M250V
C3168396|T201|COMP|61171-5|LNC|Hepatitis B virus codon M250I|Hepatitis B virus codon M250I
C3168397|T201|COMP|61172-3|LNC|Hepatitis B virus codon M250L|Hepatitis B virus codon M250L
C3168398|T201|COMP|61173-1|LNC|Hepatitis B virus codon L80I|Hepatitis B virus codon L80I
C3168399|T201|COMP|61188-9|LNC|Clindamycin.induced|Clindamycin.induced
C3169258|T201|COMP|61407-3|LNC|Amitriptyline/Creatinine|Amitriptyline/Creatinine
C3169260|T201|COMP|61408-1|LNC|Cyclobenzaprine/Creatinine|Cyclobenzaprine/Creatinine
C3169262|T201|COMP|61411-5|LNC|Desipramine/Creatinine|Desipramine/Creatinine
C3169264|T201|COMP|61414-9|LNC|Doxepin/Creatinine|Doxepin/Creatinine
C3169266|T201|COMP|61417-2|LNC|Imipramine/Creatinine|Imipramine/Creatinine
C3169268|T201|COMP|61420-6|LNC|Norhydrocodone/Creatinine|Norhydrocodone/Creatinine
C3169270|T201|COMP|61423-0|LNC|Noroxycodone/Creatinine|Noroxycodone/Creatinine
C3169272|T201|COMP|61426-3|LNC|Nortriptyline/Creatinine|Nortriptyline/Creatinine
C3169274|T201|COMP|61429-7|LNC|Tapentadol/Creatinine|Tapentadol/Creatinine
C3169284|T201|COMP|63130-9|LNC|Phoenix dactylifera Ab.IgG|Phoenix dactylifera Ab.IgG
C3169285|T201|COMP|63131-7|LNC|Carica papaya Ab.IgG|Carica papaya Ab.IgG
C3169287|T201|COMP|63132-5|LNC|Castanea sativa Ab.IgG|Castanea sativa Ab.IgG
C3169289|T201|COMP|63133-3|LNC|Goat milk Ab.IgG|Goat milk Ab.IgG
C3169290|T201|COMP|63134-1|LNC|Sardina pilchardus Ab.IgG|Sardina pilchardus Ab.IgG
C3169291|T201|COMP|63135-8|LNC|Cicer arietinus Ab.IgG|Cicer arietinus Ab.IgG
C3169293|T201|COMP|63136-6|LNC|Pimenta dioica Ab.IgG|Pimenta dioica Ab.IgG
C3169294|T201|COMP|63137-4|LNC|Astacus astacus Ab.IgG|Astacus astacus Ab.IgG
C3169296|T201|COMP|63138-2|LNC|Humulus lupus Ab.IgG|Humulus lupus Ab.IgG
C3169297|T201|COMP|63139-0|LNC|Wine Vinegar Ab.IgG|Wine Vinegar Ab.IgG
C3169298|T201|COMP|63569-8|LNC|Nuclear Ab pattern|Nuclear Ab pattern
C3169299|T201|COMP|63570-6|LNC|Nuclear Ab pattern|Nuclear Ab pattern
C3169300|T201|COMP|63571-4|LNC|Pancreatic islet cell Ab pattern|Pancreatic islet cell Ab pattern
C3169302|T201|COMP|63572-2|LNC|Time received in laboratory|Time received in laboratory
C3169303|T201|COMP|63574-8|LNC|Staphylococcus sp.coagulase negative DNA|Staphylococcus sp.coagulase negative DNA
C3169359|T201|COMP|62426-2|LNC|Bordetella sp DNA panel|Bordetella sp DNA panel
C3169361|T201|COMP|62427-0|LNC|Bordetella holmesii DNA|Bordetella holmesii DNA
C3169363|T201|COMP|62428-8|LNC|Bordetella sp DNA|Bordetella sp DNA
C3169365|T201|COMP|62429-6|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C3169366|T201|COMP|62430-4|LNC|Eastern equine encephalitis virus Ab.IgM|Eastern equine encephalitis virus Ab.IgM
C3169367|T201|COMP|62431-2|LNC|Eastern equine encephalitis virus Ab.IgG|Eastern equine encephalitis virus Ab.IgG
C3169368|T201|COMP|62432-0|LNC|La Crosse virus Ab.IgM|La Crosse virus Ab.IgM
C3169435|T201|COMP|63458-4|LNC|Artemisia vulgaris native (nArt v) 1 Ab.IgE|Artemisia vulgaris native (nArt v) 1 Ab.IgE
C3169437|T201|COMP|63459-2|LNC|Gliadin peptide Ab.IgG|Gliadin peptide Ab.IgG
C3169438|T201|COMP|63460-0|LNC|HTLV I+II Ab|HTLV I+II Ab
C3169439|T201|COMP|63461-8|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C3169440|T201|COMP|63462-6|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C3169443|T201|COMP|63464-2|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C3169474|T201|COMP|64413-8|LNC|KIR gene allele 2DL1|KIR gene allele 2DL1
C3169476|T201|COMP|64414-6|LNC|KIR gene allele 2DL2|KIR gene allele 2DL2
C3169478|T201|COMP|64415-3|LNC|KIR gene allele 2DL3|KIR gene allele 2DL3
C3169480|T201|COMP|64416-1|LNC|KIR gene allele 2DL4|KIR gene allele 2DL4
C3169482|T201|COMP|64417-9|LNC|Fragile X protein (FMRP)|Fragile X protein (FMRP)
C3169484|T201|COMP|64418-7|LNC|KIR genotyping panel|KIR genotyping panel
C3169486|T201|COMP|64419-5|LNC|KIR gene allele 2DL5|KIR gene allele 2DL5
C3169488|T201|COMP|64420-3|LNC|KIR gene allele 2DS1|KIR gene allele 2DS1
C3169490|T201|COMP|64421-1|LNC|KIR gene allele 2DS2|KIR gene allele 2DS2
C3169492|T201|COMP|64422-9|LNC|KIR gene allele 2DS3|KIR gene allele 2DS3
C3169500|T201|COMP|62418-9|LNC|Glucose/Insulin|Glucose/Insulin
C3169501|T201|COMP|62419-7|LNC|Galectin 3|Galectin 3
C3169502|T201|COMP|62420-5|LNC|Fatty acids.nonesterified^8th specimen post CFst|Fatty acids.nonesterified^8th specimen post CFst
C3169503|T201|COMP|62421-3|LNC|Fatty acids.nonesterified^9th specimen post CFst|Fatty acids.nonesterified^9th specimen post CFst
C3169504|T201|COMP|62422-1|LNC|Fatty acids.nonesterified^10th specimen post CFst|Fatty acids.nonesterified^10th specimen post CFst
C3169505|T201|COMP|62423-9|LNC|Human coronavirus HKU1 RNA|Human coronavirus HKU1 RNA
C3169507|T201|COMP|62424-7|LNC|Human bocavirus DNA|Human bocavirus DNA
C3169509|T201|COMP|62425-4|LNC|Creatinine^post XXX challenge|Creatinine^post XXX challenge
C3169510|T201|COMP|62433-8|LNC|La Crosse virus Ab.IgG|La Crosse virus Ab.IgG
C3169511|T201|COMP|62434-6|LNC|Saint Louis encephalitis virus Ab.IgM|Saint Louis encephalitis virus Ab.IgM
C3169512|T201|COMP|62435-3|LNC|Saint Louis encephalitis virus Ab.IgG|Saint Louis encephalitis virus Ab.IgG
C3169513|T201|COMP|62436-1|LNC|West Nile virus Ab.IgM|West Nile virus Ab.IgM
C3169514|T201|COMP|62437-9|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C3169515|T201|COMP|62438-7|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C3169516|T201|COMP|62439-5|LNC|Erythrocytes.nucleated|Erythrocytes.nucleated
C3169517|T201|COMP|62440-3|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C3169518|T201|COMP|62441-1|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C3169519|T201|COMP|62442-9|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C3169531|T201|COMP|62453-6|LNC|Fatty acids.ethyl esters|Fatty acids.ethyl esters
C3169534|T201|COMP|62455-1|LNC|Coccidioides sp F Ab|Coccidioides sp F Ab
C3169536|T201|COMP|62456-9|LNC|HIV 2 p15 Ab|HIV 2 p15 Ab
C3169538|T201|COMP|62457-7|LNC|Coccidioides sp TP Ab|Coccidioides sp TP Ab
C3169540|T201|COMP|62458-5|LNC|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C3169541|T201|COMP|62459-3|LNC|Coccidioides immitis Ab.IgG|Coccidioides immitis Ab.IgG
C3169542|T201|COMP|62460-1|LNC|Candida sp DNA|Candida sp DNA
C3169543|T201|COMP|62461-9|LNC|Trichomonas vaginalis DNA|Trichomonas vaginalis DNA
C3169544|T201|COMP|62462-7|LNC|Influenza virus A+B RNA|Influenza virus A+B RNA
C3169545|T201|COMP|62463-5|LNC|Enterovirus RNA|Enterovirus RNA
C3169546|T201|COMP|62464-3|LNC|Enterovirus RNA|Enterovirus RNA
C3169547|T201|COMP|62465-0|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C3169548|T201|COMP|62466-8|LNC|BK virus Ab.IgG|BK virus Ab.IgG
C3169550|T201|COMP|62467-6|LNC|Galactomannan Ag|Galactomannan Ag
C3169551|T201|COMP|62468-4|LNC|1,3 beta glucan|1,3 beta glucan
C3169552|T201|COMP|62469-2|LNC|HIV 1 RNA|HIV 1 RNA
C3169553|T201|COMP|62470-0|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C3169554|T201|COMP|62471-8|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C3169555|T201|COMP|62472-6|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C3169556|T201|COMP|62473-4|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C3169557|T201|COMP|62474-2|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C3169558|T201|COMP|62475-9|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C3169559|T201|COMP|62476-7|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C3169560|T201|COMP|62477-5|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C3169561|T201|COMP|62478-3|LNC|Aspergillus fumigatus DNA|Aspergillus fumigatus DNA
C3169563|T201|COMP|62479-1|LNC|Aspergillus terreus DNA|Aspergillus terreus DNA
C3169565|T201|COMP|62480-9|LNC|Adenovirus DNA|Adenovirus DNA
C3169566|T201|COMP|62481-7|LNC|Herpes virus 6A DNA|Herpes virus 6A DNA
C3169568|T201|COMP|62482-5|LNC|Herpes virus 6B DNA|Herpes virus 6B DNA
C3169570|T201|COMP|62483-3|LNC|Herpes virus 6A DNA|Herpes virus 6A DNA
C3169571|T201|COMP|62484-1|LNC|Herpes virus 6B DNA|Herpes virus 6B DNA
C3169572|T201|COMP|62485-8|LNC|Herpes virus 6A DNA|Herpes virus 6A DNA
C3169573|T201|COMP|62486-6|LNC|Herpes virus 6B DNA|Herpes virus 6B DNA
C3169574|T201|COMP|62487-4|LNC|Urobilinogen|Urobilinogen
C3169575|T201|COMP|62488-2|LNC|Ova1 test|Ova1 test
C3169577|T201|COMP|62489-0|LNC|Sulfate.inorganic|Sulfate.inorganic
C3171808|T201|COMP|63193-7|LNC|Artemisia tridentata Ab.IgG|Artemisia tridentata Ab.IgG
C3171809|T201|COMP|63194-5|LNC|Medicago sativa Ab.IgG|Medicago sativa Ab.IgG
C3171810|T201|COMP|63337-0|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C3171811|T201|COMP|63338-8|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C3171812|T201|COMP|63339-6|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C3171813|T201|COMP|63340-4|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C3171814|T201|COMP|63341-2|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C3171853|T201|COMP|62848-7|LNC|Mirtazapine+Normirtazapine|Mirtazapine+Normirtazapine
C3171855|T201|COMP|62849-5|LNC|Venlafaxine+Norvenlafaxine|Venlafaxine+Norvenlafaxine
C3171862|T201|COMP|62857-8|LNC|Micromegakaryocytes|Micromegakaryocytes
C3171863|T201|COMP|62858-6|LNC|Micromegakaryocytes/100 leukocytes|Micromegakaryocytes/100 leukocytes
C3171865|T201|COMP|62859-4|LNC|Rotavirus RNA|Rotavirus RNA
C3171866|T201|COMP|62860-2|LNC|Influenza virus C RNA|Influenza virus C RNA
C3171867|T201|COMP|62861-0|LNC|Enterovirus 71 RNA|Enterovirus 71 RNA
C3171868|T201|COMP|62862-8|LNC|Microsatellite instability|Microsatellite instability
C3171935|T201|COMP|62946-9|LNC|Jamestown canyon virus Ab.IgM|Jamestown canyon virus Ab.IgM
C3171936|T201|COMP|62947-7|LNC|MPL gene.p.Trp515Leu+Trp515Lys+Ser505Asn|MPL gene.p.Trp515Leu+Trp515Lys+Ser505Asn
C3171938|T201|COMP|62948-5|LNC|MPL gene mutations tested for|MPL gene mutations tested for
C3172011|T201|COMP|63042-6|LNC|17-Hydroxyprogesterone/Creatinine|17-Hydroxyprogesterone/Creatinine
C3172012|T201|COMP|63043-4|LNC|Nuclei scored|Nuclei scored
C3172014|T201|COMP|63044-2|LNC|Cotinine|Cotinine
C3172038|T201|COMP|63068-1|LNC|TOP2A gene copy number/Chromosome 17 copy number|TOP2A gene copy number/Chromosome 17 copy number
C3172040|T201|COMP|63069-9|LNC|TOP2A gene|TOP2A gene
C3172041|T201|COMP|63070-7|LNC|TOP2A gene 17q21-22 deletion+duplication|TOP2A gene 17q21-22 deletion+duplication
C3172047|T201|COMP|63075-6|LNC|Dermatophagoides farinae Ab.IgG|Dermatophagoides farinae Ab.IgG
C3172048|T201|COMP|63076-4|LNC|Cat dander Ab.IgG|Cat dander Ab.IgG
C3172049|T201|COMP|63077-2|LNC|Dog dander Ab.IgG|Dog dander Ab.IgG
C3172050|T201|COMP|63078-0|LNC|Fagopyrum esculentum Ab.IgG|Fagopyrum esculentum Ab.IgG
C3172051|T201|COMP|63079-8|LNC|Bean white Ab.IgG|Bean white Ab.IgG
C3172052|T201|COMP|63080-6|LNC|Corylus avellana Ab.IgG|Corylus avellana Ab.IgG
C3172053|T201|COMP|63081-4|LNC|Bertholletia excelsa Ab.IgG|Bertholletia excelsa Ab.IgG
C3172054|T201|COMP|63082-2|LNC|Pepper cayenne Ab.IgG|Pepper cayenne Ab.IgG
C3172055|T201|COMP|63083-0|LNC|Rubus idaeus Ab.IgG|Rubus idaeus Ab.IgG
C3172056|T201|COMP|63084-8|LNC|Cocos nucifera Ab.IgG|Cocos nucifera Ab.IgG
C3172057|T201|COMP|63085-5|LNC|Mytilus edulis Ab.IgG|Mytilus edulis Ab.IgG
C3172058|T201|COMP|63086-3|LNC|Scomber japonicus Ab.IgG|Scomber japonicus Ab.IgG
C3172059|T201|COMP|63087-1|LNC|Panicum milliaceum Ab.IgG|Panicum milliaceum Ab.IgG
C3172060|T201|COMP|63088-9|LNC|Perca spp Ab.IgG|Perca spp Ab.IgG
C3172061|T201|COMP|63089-7|LNC|Cheese parmesan Ab.IgG|Cheese parmesan Ab.IgG
C3172063|T201|COMP|63090-5|LNC|Beta lactoglobulin Ab.IgG|Beta lactoglobulin Ab.IgG
C3172064|T201|COMP|63091-3|LNC|Gluten Ab.IgG|Gluten Ab.IgG
C3172065|T201|COMP|63092-1|LNC|Cheese cheddar type Ab.IgG|Cheese cheddar type Ab.IgG
C3172066|T201|COMP|63093-9|LNC|Actinidia chinensis Ab.IgG|Actinidia chinensis Ab.IgG
C3172067|T201|COMP|63094-7|LNC|Petroselinum crispum Ab.IgG|Petroselinum crispum Ab.IgG
C3172068|T201|COMP|63095-4|LNC|Cucumis melo spp Ab.IgG|Cucumis melo spp Ab.IgG
C3172069|T201|COMP|63096-2|LNC|Mangifera indica Ab.IgG|Mangifera indica Ab.IgG
C3172070|T201|COMP|63097-0|LNC|Cottonseed Ab.IgG|Cottonseed Ab.IgG
C3172071|T201|COMP|63098-8|LNC|Venison Ab.IgG|Venison Ab.IgG
C3172072|T201|COMP|63099-6|LNC|Cheese American Ab.IgG|Cheese American Ab.IgG
C3172073|T201|COMP|63100-2|LNC|Vigna sinensis Ab.IgG|Vigna sinensis Ab.IgG
C3172074|T201|COMP|63101-0|LNC|Duck meat Ab.IgG|Duck meat Ab.IgG
C3172076|T201|COMP|63102-8|LNC|Prunus persica var nucipersica Ab.IgG|Prunus persica var nucipersica Ab.IgG
C3172077|T201|COMP|63103-6|LNC|Cheese swiss Ab.IgG|Cheese swiss Ab.IgG
C3172078|T201|COMP|63104-4|LNC|Vaccinium oxycoccos Ab.IgG|Vaccinium oxycoccos Ab.IgG
C3172079|T201|COMP|63105-1|LNC|Rheum spp Ab.IgG|Rheum spp Ab.IgG
C3172080|T201|COMP|63106-9|LNC|Phaseolus limensis Ab.IgG|Phaseolus limensis Ab.IgG
C3172081|T201|COMP|63107-7|LNC|Linum usitatissimum Ab.IgG|Linum usitatissimum Ab.IgG
C3172083|T201|COMP|63108-5|LNC|Carya illinoinensis nut Ab.IgG|Carya illinoinensis nut Ab.IgG
C3172084|T201|COMP|63109-3|LNC|Anacardium occidentale Ab.IgG|Anacardium occidentale Ab.IgG
C3172085|T201|COMP|63110-1|LNC|Pistacia vera Ab.IgG|Pistacia vera Ab.IgG
C3172086|T201|COMP|63111-9|LNC|Clupea harengus Ab.IgG|Clupea harengus Ab.IgG
C3172087|T201|COMP|63112-7|LNC|Rubus fruticosus Ab.IgG|Rubus fruticosus Ab.IgG
C3172088|T201|COMP|63113-5|LNC|Rabbit Ab.IgG|Rabbit Ab.IgG
C3172089|T201|COMP|63114-3|LNC|Capsicum annuum Ab.IgG|Capsicum annuum Ab.IgG
C3172090|T201|COMP|63115-0|LNC|Papaver somniferum Ab.IgG|Papaver somniferum Ab.IgG
C3172092|T201|COMP|63116-8|LNC|Cucurbita pepo Ab.IgG|Cucurbita pepo Ab.IgG
C3172094|T201|COMP|63117-6|LNC|Carthamus tinctorius Ab.IgG|Carthamus tinctorius Ab.IgG
C3172095|T201|COMP|63118-4|LNC|Lens esculenta Ab.IgG|Lens esculenta Ab.IgG
C3172096|T201|COMP|63119-2|LNC|Honey Ab.IgG|Honey Ab.IgG
C3172097|T201|COMP|63120-0|LNC|Juglans spp Ab.IgG|Juglans spp Ab.IgG
C3172098|T201|COMP|63121-8|LNC|Loligo sp Ab.IgG|Loligo sp Ab.IgG
C3172100|T201|COMP|63122-6|LNC|Anguilla anguilla Ab.IgG|Anguilla anguilla Ab.IgG
C3172102|T201|COMP|63123-4|LNC|Cuminum cyminum Ab.IgG|Cuminum cyminum Ab.IgG
C3172104|T201|COMP|63124-2|LNC|Ocimum basilicum Ab.IgG|Ocimum basilicum Ab.IgG
C3172105|T201|COMP|63125-9|LNC|Thymus vulgaris Ab.IgG|Thymus vulgaris Ab.IgG
C3172106|T201|COMP|63126-7|LNC|Foeniculum vulgare fresh Ab.IgG|Foeniculum vulgare fresh Ab.IgG
C3172108|T201|COMP|63127-5|LNC|Anethum graveolens Ab.IgG|Anethum graveolens Ab.IgG
C3172109|T201|COMP|63128-3|LNC|Laurus nobilis Ab.IgG|Laurus nobilis Ab.IgG
C3172110|T201|COMP|63129-1|LNC|Curry Ab.IgG|Curry Ab.IgG
C3172111|T201|COMP|63140-8|LNC|Gelatin Ab.IgG|Gelatin Ab.IgG
C3172112|T201|COMP|63141-6|LNC|Yogurt Ab.IgG|Yogurt Ab.IgG
C3172113|T201|COMP|63142-4|LNC|Micropterus salmoides Ab.IgG|Micropterus salmoides Ab.IgG
C3172115|T201|COMP|63143-2|LNC|Ictalurus punctatus Ab.IgG|Ictalurus punctatus Ab.IgG
C3172117|T201|COMP|63144-0|LNC|Cichorium intybus Ab.IgG|Cichorium intybus Ab.IgG
C3172119|T201|COMP|63145-7|LNC|Gum arabic Ab.IgG|Gum arabic Ab.IgG
C3172121|T201|COMP|63146-5|LNC|Karaya gum Ab.IgG|Karaya gum Ab.IgG
C3172123|T201|COMP|63147-3|LNC|Armoracia rusticana Ab.IgG|Armoracia rusticana Ab.IgG
C3172124|T201|COMP|63148-1|LNC|Maple syrup Ab.IgG|Maple syrup Ab.IgG
C3172125|T201|COMP|63149-9|LNC|Abelmoschus esculentus Ab.IgG|Abelmoschus esculentus Ab.IgG
C3172127|T201|COMP|63150-7|LNC|Pastinaca sativa Ab.IgG|Pastinaca sativa Ab.IgG
C3172130|T201|COMP|63152-3|LNC|Cynodon dactylon Ab.IgG|Cynodon dactylon Ab.IgG
C3172131|T201|COMP|63153-1|LNC|Sorghum halepense Ab.IgG|Sorghum halepense Ab.IgG
C3172132|T201|COMP|63154-9|LNC|Secale cereale pollen Ab.IgG|Secale cereale pollen Ab.IgG
C3172133|T201|COMP|63155-6|LNC|Triticum aestivum pollen Ab.IgG|Triticum aestivum pollen Ab.IgG
C3172134|T201|COMP|63156-4|LNC|Paspalum notatum Ab.IgG|Paspalum notatum Ab.IgG
C3172135|T201|COMP|63157-2|LNC|House dust Greer Ab.IgG|House dust Greer Ab.IgG
C3172136|T201|COMP|63158-0|LNC|House dust Hollister Stier Ab.IgG|House dust Hollister Stier Ab.IgG
C3172137|T201|COMP|63159-8|LNC|Ctenocephalides sp Ab.IgG|Ctenocephalides sp Ab.IgG
C3172138|T201|COMP|63160-6|LNC|Ricinus communis Ab.IgG|Ricinus communis Ab.IgG
C3172139|T201|COMP|63161-4|LNC|Latex Ab.IgG|Latex Ab.IgG
C3172140|T201|COMP|63162-2|LNC|Curvularia lunata Ab.IgG|Curvularia lunata Ab.IgG
C3172141|T201|COMP|63163-0|LNC|Paecilomyces sp Ab.IgG|Paecilomyces sp Ab.IgG
C3172143|T201|COMP|63164-8|LNC|Penicillium brevicompactum Ab.IgG|Penicillium brevicompactum Ab.IgG
C3172144|T201|COMP|63165-5|LNC|Serpula lacrymans Ab.IgG|Serpula lacrymans Ab.IgG
C3172145|T201|COMP|63166-3|LNC|Aspergillus terreus Ab.IgG|Aspergillus terreus Ab.IgG
C3172147|T201|COMP|63167-1|LNC|Trichophyton mentagrophytes Ab.IgG|Trichophyton mentagrophytes Ab.IgG
C3172148|T201|COMP|63168-9|LNC|Aspergillus amstelodami Ab.IgG|Aspergillus amstelodami Ab.IgG
C3172150|T201|COMP|63169-7|LNC|Aspergillus nidulans Ab.IgG|Aspergillus nidulans Ab.IgG
C3172151|T201|COMP|63170-5|LNC|Helminthosporium interseminatum Ab.IgG|Helminthosporium interseminatum Ab.IgG
C3172153|T201|COMP|63171-3|LNC|Neurospora sitophila Ab.IgG|Neurospora sitophila Ab.IgG
C3172155|T201|COMP|63172-1|LNC|Mucor plumbeus Ab.IgG|Mucor plumbeus Ab.IgG
C3172157|T201|COMP|63173-9|LNC|Mycogone perniciosa Ab.IgG|Mycogone perniciosa Ab.IgG
C3172159|T201|COMP|63174-7|LNC|Spondylocladium sp Ab.IgG|Spondylocladium sp Ab.IgG
C3172160|T201|COMP|63175-4|LNC|Epidermophyton floccosum Ab.IgG|Epidermophyton floccosum Ab.IgG
C3172162|T201|COMP|63176-2|LNC|Algae Ab.IgG|Algae Ab.IgG
C3172164|T201|COMP|63177-0|LNC|Acremonium sp Ab.IgG|Acremonium sp Ab.IgG
C3172165|T201|COMP|63178-8|LNC|Chaetomium globosum Ab.IgG|Chaetomium globosum Ab.IgG
C3172166|T201|COMP|63179-6|LNC|Sphacelotheca cruenta Ab.IgG|Sphacelotheca cruenta Ab.IgG
C3172167|T201|COMP|63180-4|LNC|Nicotiana tabacum Ab.IgG|Nicotiana tabacum Ab.IgG
C3172168|T201|COMP|63181-2|LNC|Juniperus sabinoides Ab.IgG|Juniperus sabinoides Ab.IgG
C3172169|T201|COMP|63182-0|LNC|Quercus alba Ab.IgG|Quercus alba Ab.IgG
C3172170|T201|COMP|63183-8|LNC|Populus deltoides Ab.IgG|Populus deltoides Ab.IgG
C3172171|T201|COMP|63184-6|LNC|Fraxinus americana Ab.IgG|Fraxinus americana Ab.IgG
C3172172|T201|COMP|63185-3|LNC|Prosopis juliflora Ab.IgG|Prosopis juliflora Ab.IgG
C3172173|T201|COMP|63186-1|LNC|Chenopodium album Ab.IgG|Chenopodium album Ab.IgG
C3172174|T201|COMP|63313-1|LNC|Rheumatoid factor|Rheumatoid factor
C3172175|T201|COMP|63314-9|LNC|Rheumatoid factor.IgA|Rheumatoid factor.IgA
C3172176|T201|COMP|63315-6|LNC|Rheumatoid factor.IgM|Rheumatoid factor.IgM
C3172177|T201|COMP|63316-4|LNC|U1 small nuclear ribonucleoprotein 70kD Ab|U1 small nuclear ribonucleoprotein 70kD Ab
C3172178|T201|COMP|63317-2|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C3172179|T201|COMP|63318-0|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C3172180|T201|COMP|63319-8|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C3172181|T201|COMP|63320-6|LNC|Ribosomal Ab|Ribosomal Ab
C3172182|T201|COMP|63321-4|LNC|Ribosomal Ab|Ribosomal Ab
C3172183|T201|COMP|63322-2|LNC|Ribosomal Ab|Ribosomal Ab
C3172184|T201|COMP|63323-0|LNC|Ribosomal Ab|Ribosomal Ab
C3172185|T201|COMP|63324-8|LNC|Ribosomal Ab.IgG|Ribosomal Ab.IgG
C3172186|T201|COMP|63325-5|LNC|Ribosomal Ab.IgG|Ribosomal Ab.IgG
C3172187|T201|COMP|63326-3|LNC|Ribosomal P Ab|Ribosomal P Ab
C3172188|T201|COMP|63327-1|LNC|Ribosomal P Ab|Ribosomal P Ab
C3172189|T201|COMP|63449-3|LNC|Cells.CD3|Cells.CD3
C3172190|T201|COMP|63450-1|LNC|Cells.CD3+CD4+|Cells.CD3+CD4+
C3172191|T201|COMP|63451-9|LNC|Cells.CD3+CD8+|Cells.CD3+CD8+
C3172192|T201|COMP|63452-7|LNC|Cells.CD3-CD7+/100 cells|Cells.CD3-CD7+/100 cells
C3172193|T201|COMP|63453-5|LNC|Gliadin peptide Ab.IgA|Gliadin peptide Ab.IgA
C3172194|T201|COMP|63454-3|LNC|TPMT gene mutations tested for|TPMT gene mutations tested for
C3172196|T201|COMP|63455-0|LNC|Coxiella burnetii phase 1 Ab.IgM|Coxiella burnetii phase 1 Ab.IgM
C3172231|T201|COMP|63187-9|LNC|Salsola kali Ab.IgG|Salsola kali Ab.IgG
C3172232|T201|COMP|63188-7|LNC|Xanthium commune Ab.IgG|Xanthium commune Ab.IgG
C3172233|T201|COMP|63189-5|LNC|Pigweed rough Ab.IgG|Pigweed rough Ab.IgG
C3172234|T201|COMP|63190-3|LNC|Iva ciliata Ab.IgG|Iva ciliata Ab.IgG
C3172235|T201|COMP|63191-1|LNC|Urtica dioica Ab.IgG|Urtica dioica Ab.IgG
C3172236|T201|COMP|63192-9|LNC|Rumex crispus Ab.IgG|Rumex crispus Ab.IgG
C3172237|T201|COMP|63342-0|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C3172238|T201|COMP|63343-8|LNC|Sjogrens syndrome-A extractable nuclear 60kD Ab|Sjogrens syndrome-A extractable nuclear 60kD Ab
C3172239|T201|COMP|63470-9|LNC|Ganglioside GM4 Ab.IgG|Ganglioside GM4 Ab.IgG
C3172240|T201|COMP|63471-7|LNC|Ganglioside GD2 Ab.IgG|Ganglioside GD2 Ab.IgG
C3172241|T201|COMP|63472-5|LNC|Ganglioside GD3 Ab.IgG|Ganglioside GD3 Ab.IgG
C3172242|T201|COMP|63473-3|LNC|Gadus morhua recombinant (rGad c) 1 Ab.IgE|Gadus morhua recombinant (rGad c) 1 Ab.IgE
C3172244|T201|COMP|63474-1|LNC|Albumin|Albumin
C3172245|T201|COMP|63475-8|LNC|BK virus DNA|BK virus DNA
C3172246|T201|COMP|63476-6|LNC|Glycine max recombinant (rGly m) 4 Ab.IgE|Glycine max recombinant (rGly m) 4 Ab.IgE
C3172248|T201|COMP|63477-4|LNC|Arachis hypogaea recombinant (rAra h) 8 Ab.IgE|Arachis hypogaea recombinant (rAra h) 8 Ab.IgE
C3172275|T201|COMP|63195-2|LNC|Helianthus annuus pollen Ab.IgG|Helianthus annuus pollen Ab.IgG
C3172282|T201|COMP|63200-0|LNC|Solidago virgaurea Ab.IgG|Solidago virgaurea Ab.IgG
C3172283|T201|COMP|63201-8|LNC|Beet red Ab.IgG|Beet red Ab.IgG
C3172285|T201|COMP|63202-6|LNC|Morus alba Ab.IgG|Morus alba Ab.IgG
C3172286|T201|COMP|63203-4|LNC|Alnus rugosa Ab.IgG|Alnus rugosa Ab.IgG
C3172287|T201|COMP|63204-2|LNC|Ligustrum vulgare Ab.IgG|Ligustrum vulgare Ab.IgG
C3172288|T201|COMP|63205-9|LNC|Populus tremula Ab.IgG|Populus tremula Ab.IgG
C3172289|T201|COMP|63206-7|LNC|Ambrosia elatior Ab.IgG|Ambrosia elatior Ab.IgG
C3172290|T201|COMP|63207-5|LNC|Franseria acanthicarpa Ab.IgG|Franseria acanthicarpa Ab.IgG
C3172291|T201|COMP|63208-3|LNC|Artemisia vulgaris Ab.IgG|Artemisia vulgaris Ab.IgG
C3172292|T201|COMP|63209-1|LNC|Plantago lanceolata Ab.IgG|Plantago lanceolata Ab.IgG
C3172293|T201|COMP|63210-9|LNC|Actin.smooth muscle Ab|Actin.smooth muscle Ab
C3172294|T201|COMP|63211-7|LNC|Actin.smooth muscle Ab|Actin.smooth muscle Ab
C3172295|T201|COMP|63212-5|LNC|Asialoganglioside GM1 Ab.IgG|Asialoganglioside GM1 Ab.IgG
C3172296|T201|COMP|63213-3|LNC|Bactericidal permeability increasing protein Ab|Bactericidal permeability increasing protein Ab
C3172297|T201|COMP|63214-1|LNC|Bactericidal permeability increasing protein Ab|Bactericidal permeability increasing protein Ab
C3172298|T201|COMP|63215-8|LNC|Cathepsin G Ab|Cathepsin G Ab
C3172299|T201|COMP|63216-6|LNC|CV2 Ab|CV2 Ab
C3172300|T201|COMP|63217-4|LNC|Cyclic citrullinated peptide Ab.IgG|Cyclic citrullinated peptide Ab.IgG
C3172301|T201|COMP|63218-2|LNC|Desmoglein 1 Ab|Desmoglein 1 Ab
C3172302|T201|COMP|63219-0|LNC|Desmoglein 3 Ab|Desmoglein 3 Ab
C3172303|T201|COMP|63220-8|LNC|DNA double strand Ab|DNA double strand Ab
C3172304|T201|COMP|63221-6|LNC|DNA double strand Ab|DNA double strand Ab
C3172305|T201|COMP|63222-4|LNC|DNA double strand Ab|DNA double strand Ab
C3172306|T201|COMP|63223-2|LNC|DNA double strand Ab|DNA double strand Ab
C3172307|T201|COMP|63224-0|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172308|T201|COMP|63225-7|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172309|T201|COMP|63226-5|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172310|T201|COMP|63227-3|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172311|T201|COMP|63228-1|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172312|T201|COMP|63229-9|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172313|T201|COMP|63230-7|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172314|T201|COMP|63231-5|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172315|T201|COMP|63232-3|LNC|DNA double strand Ab.IgM|DNA double strand Ab.IgM
C3172317|T201|COMP|63233-1|LNC|DNA double strand Ab.IgM|DNA double strand Ab.IgM
C3172318|T201|COMP|63234-9|LNC|DNA double strand Ab.IgM|DNA double strand Ab.IgM
C3172319|T201|COMP|63235-6|LNC|DNA double strand Ab.IgM|DNA double strand Ab.IgM
C3172320|T201|COMP|63236-4|LNC|DNA double strand Ab.IgM|DNA double strand Ab.IgM
C3172321|T201|COMP|63237-2|LNC|DNA double strand Ab.IgM|DNA double strand Ab.IgM
C3172322|T201|COMP|63238-0|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C3172323|T201|COMP|63239-8|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C3172324|T201|COMP|63240-6|LNC|Ganglioside GD3 Ab.IgG+IgM|Ganglioside GD3 Ab.IgG+IgM
C3172326|T201|COMP|63241-4|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C3172327|T201|COMP|63242-2|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C3172328|T201|COMP|63243-0|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C3172329|T201|COMP|63244-8|LNC|Ganglioside GM1 Ab.IgG+IgM|Ganglioside GM1 Ab.IgG+IgM
C3172330|T201|COMP|63245-5|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C3172331|T201|COMP|63246-3|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C3172332|T201|COMP|63247-1|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C3172333|T201|COMP|63248-9|LNC|Ganglioside GM2 Ab.IgG|Ganglioside GM2 Ab.IgG
C3172334|T201|COMP|63249-7|LNC|Ganglioside GM2 Ab.IgG+IgM|Ganglioside GM2 Ab.IgG+IgM
C3172336|T201|COMP|63250-5|LNC|Ganglioside GM2 Ab.IgM|Ganglioside GM2 Ab.IgM
C3172337|T201|COMP|63251-3|LNC|Ganglioside GM3 Ab.IgG|Ganglioside GM3 Ab.IgG
C3172338|T201|COMP|63252-1|LNC|Ganglioside GM3 Ab.IgG+IgM|Ganglioside GM3 Ab.IgG+IgM
C3172340|T201|COMP|63253-9|LNC|Ganglioside GM3 Ab.IgM|Ganglioside GM3 Ab.IgM
C3172341|T201|COMP|63254-7|LNC|Ganglioside GQ1b Ab.IgG|Ganglioside GQ1b Ab.IgG
C3172342|T201|COMP|63255-4|LNC|Ganglioside GQ1b Ab.IgM|Ganglioside GQ1b Ab.IgM
C3172343|T201|COMP|63256-2|LNC|Ganglioside GT1a Ab.IgG+IgM|Ganglioside GT1a Ab.IgG+IgM
C3172345|T201|COMP|63257-0|LNC|Ganglioside GT1b Ab.IgG|Ganglioside GT1b Ab.IgG
C3172346|T201|COMP|63258-8|LNC|Ganglioside GT1b Ab.IgG+IgM|Ganglioside GT1b Ab.IgG+IgM
C3172348|T201|COMP|63259-6|LNC|Ganglioside GT1b Ab.IgM|Ganglioside GT1b Ab.IgM
C3172349|T201|COMP|63260-4|LNC|Gliadin Ab.IgA|Gliadin Ab.IgA
C3172350|T201|COMP|63261-2|LNC|Gliadin Ab.IgG|Gliadin Ab.IgG
C3172351|T201|COMP|63262-0|LNC|Glomerular basement membrane Ab|Glomerular basement membrane Ab
C3172352|T201|COMP|63263-8|LNC|Histone Ab|Histone Ab
C3172353|T201|COMP|63264-6|LNC|Histone Ab|Histone Ab
C3172354|T201|COMP|63265-3|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C3172355|T201|COMP|63266-1|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C3172356|T201|COMP|63267-9|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C3172357|T201|COMP|63268-7|LNC|Keratin Ab|Keratin Ab
C3172358|T201|COMP|63269-5|LNC|Ku Ab|Ku Ab
C3172359|T201|COMP|63270-3|LNC|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C3172360|T201|COMP|63271-1|LNC|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C3172361|T201|COMP|63272-9|LNC|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C3172362|T201|COMP|63273-7|LNC|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C3172363|T201|COMP|63274-5|LNC|Liver kidney microsomal 2 Ab|Liver kidney microsomal 2 Ab
C3172365|T201|COMP|63275-2|LNC|Liver kidney microsomal 2 Ab|Liver kidney microsomal 2 Ab
C3172366|T201|COMP|63276-0|LNC|Mi-2 Ab|Mi-2 Ab
C3172367|T201|COMP|63277-8|LNC|Mitochondria Ab|Mitochondria Ab
C3172368|T201|COMP|63278-6|LNC|Mitochondria Ab|Mitochondria Ab
C3172369|T201|COMP|63279-4|LNC|Mitochondria Ab|Mitochondria Ab
C3172370|T201|COMP|63280-2|LNC|Mitochondria Ab|Mitochondria Ab
C3172371|T201|COMP|63281-0|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C3172372|T201|COMP|63282-8|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C3172373|T201|COMP|63283-6|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C3172374|T201|COMP|63284-4|LNC|Mitochondria M5 Ab|Mitochondria M5 Ab
C3172376|T201|COMP|63285-1|LNC|Mitochondria M5 Ab|Mitochondria M5 Ab
C3172377|T201|COMP|63286-9|LNC|Myelin Ab|Myelin Ab
C3172378|T201|COMP|63287-7|LNC|Myelin Ab|Myelin Ab
C3172379|T201|COMP|63288-5|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C3172380|T201|COMP|63289-3|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C3172381|T201|COMP|63290-1|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C3172382|T201|COMP|63291-9|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C3172383|T201|COMP|63292-7|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C3172384|T201|COMP|63293-5|LNC|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C3172385|T201|COMP|63294-3|LNC|Nuclear Ab|Nuclear Ab
C3172386|T201|COMP|63295-0|LNC|Nuclear Ab|Nuclear Ab
C3172387|T201|COMP|63296-8|LNC|Nuclear Ab|Nuclear Ab
C3172388|T201|COMP|63297-6|LNC|Nuclear Ab|Nuclear Ab
C3172389|T201|COMP|63298-4|LNC|Nucleosome Ab|Nucleosome Ab
C3172390|T201|COMP|63299-2|LNC|Nucleosome Ab|Nucleosome Ab
C3172391|T201|COMP|63300-8|LNC|Nucleosome Ab|Nucleosome Ab
C3172392|T201|COMP|63301-6|LNC|Parathyrin Ab|Parathyrin Ab
C3172393|T201|COMP|63302-4|LNC|Parathyrin Ab|Parathyrin Ab
C3172394|T201|COMP|63303-2|LNC|Parietal cell Ab|Parietal cell Ab
C3172395|T201|COMP|63304-0|LNC|Parietal cell Ab|Parietal cell Ab
C3172396|T201|COMP|63305-7|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C3172397|T201|COMP|63306-5|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C3172398|T201|COMP|63307-3|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C3172399|T201|COMP|63308-1|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C3172400|T201|COMP|63309-9|LNC|Proteinase 3 Ab|Proteinase 3 Ab
C3172401|T201|COMP|63310-7|LNC|Proteinase 3 Ab|Proteinase 3 Ab
C3172402|T201|COMP|63311-5|LNC|Proteinase 3 Ab|Proteinase 3 Ab
C3172403|T201|COMP|63312-3|LNC|Purkinje cells Ab|Purkinje cells Ab
C3172404|T201|COMP|63328-9|LNC|RNA polymerase III Ab|RNA polymerase III Ab
C3172405|T201|COMP|63329-7|LNC|RNA polymerase III Ab|RNA polymerase III Ab
C3172406|T201|COMP|63330-5|LNC|Saccharomyces cerevisiae Ab.IgA|Saccharomyces cerevisiae Ab.IgA
C3172407|T201|COMP|63331-3|LNC|Saccharomyces cerevisiae Ab.IgA|Saccharomyces cerevisiae Ab.IgA
C3172408|T201|COMP|63332-1|LNC|Saccharomyces cerevisiae Ab.IgG|Saccharomyces cerevisiae Ab.IgG
C3172409|T201|COMP|63333-9|LNC|Saccharomyces cerevisiae Ab.IgG|Saccharomyces cerevisiae Ab.IgG
C3172410|T201|COMP|63334-7|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C3172411|T201|COMP|63335-4|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C3172412|T201|COMP|63336-2|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C3172413|T201|COMP|63344-6|LNC|Sjogrens syndrome-A extractable nuclear 60kD Ab|Sjogrens syndrome-A extractable nuclear 60kD Ab
C3172414|T201|COMP|63345-3|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C3172415|T201|COMP|63346-1|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C3172416|T201|COMP|63347-9|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C3172417|T201|COMP|63348-7|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C3172418|T201|COMP|63349-5|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C3172419|T201|COMP|63350-3|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C3172420|T201|COMP|63351-1|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C3172421|T201|COMP|63352-9|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C3172422|T201|COMP|63353-7|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C3172423|T201|COMP|63354-5|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C3172424|T201|COMP|63355-2|LNC|Smooth muscle Ab|Smooth muscle Ab
C3172425|T201|COMP|63356-0|LNC|Smooth muscle Ab|Smooth muscle Ab
C3172426|T201|COMP|63357-8|LNC|Smooth muscle Ab|Smooth muscle Ab
C3172427|T201|COMP|63358-6|LNC|Smooth muscle Ab|Smooth muscle Ab
C3172428|T201|COMP|63359-4|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C3172429|T201|COMP|63360-2|LNC|Thyroglobulin Ab|Thyroglobulin Ab
C3172430|T201|COMP|63361-0|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C3172431|T201|COMP|63362-8|LNC|Thyroperoxidase Ab|Thyroperoxidase Ab
C3172432|T201|COMP|63363-6|LNC|Thyrotropin receptor Ab|Thyrotropin receptor Ab
C3172433|T201|COMP|63364-4|LNC|Thyrotropin receptor Ab|Thyrotropin receptor Ab
C3172434|T201|COMP|63365-1|LNC|Thyrotropin receptor Ab|Thyrotropin receptor Ab
C3172435|T201|COMP|63366-9|LNC|Thyrotropin receptor Ab|Thyrotropin receptor Ab
C3172436|T201|COMP|63367-7|LNC|U1 small nuclear ribonucleoprotein Ab|U1 small nuclear ribonucleoprotein Ab
C3172437|T201|COMP|63368-5|LNC|Carbapenem resistance genes|Carbapenem resistance genes
C3172439|T201|COMP|63369-3|LNC|Chronic urticaria index|Chronic urticaria index
C3172441|T201|COMP|63370-1|LNC|Gamma tocopherol|Gamma tocopherol
C3172442|T201|COMP|63371-9|LNC|Ketones^1H post dose glucose|Ketones^1H post dose glucose
C3172443|T201|COMP|63372-7|LNC|Ketones^3H post dose glucose|Ketones^3H post dose glucose
C3172444|T201|COMP|63373-5|LNC|Ketones^4H post dose glucose|Ketones^4H post dose glucose
C3172445|T201|COMP|63374-3|LNC|Fusarium roseum Ab.IgE|Fusarium roseum Ab.IgE
C3172447|T201|COMP|63375-0|LNC|Cyclic citrullinated peptide Ab.IgA+IgG|Cyclic citrullinated peptide Ab.IgA+IgG
C3172448|T201|COMP|63376-8|LNC|Lactoferrin|Lactoferrin
C3172449|T201|COMP|63378-4|LNC|Erythrocyte clumps|Erythrocyte clumps
C3172450|T201|COMP|63379-2|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172451|T201|COMP|63380-0|LNC|Methionine|Methionine
C3172452|T201|COMP|63381-8|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172453|T201|COMP|63382-6|LNC|Glucose^post CFst|Glucose^post CFst
C3172454|T201|COMP|63383-4|LNC|Amphiphysin Ab|Amphiphysin Ab
C3172455|T201|COMP|63384-2|LNC|Asialoganglioside GM1 Ab.IgM|Asialoganglioside GM1 Ab.IgM
C3172456|T201|COMP|63385-9|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172457|T201|COMP|63386-7|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172458|T201|COMP|63387-5|LNC|Elastase Ab|Elastase Ab
C3172459|T201|COMP|63388-3|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C3172460|T201|COMP|63389-1|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C3172461|T201|COMP|63390-9|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C3172462|T201|COMP|63391-7|LNC|Extractable nuclear Ab|Extractable nuclear Ab
C3172463|T201|COMP|63392-5|LNC|Herpes gestationis Ab|Herpes gestationis Ab
C3172464|T201|COMP|63393-3|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C3172465|T201|COMP|63394-1|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C3172466|T201|COMP|63395-8|LNC|Liver cytosol Ab|Liver cytosol Ab
C3172467|T201|COMP|63396-6|LNC|Myelin associated glycoprotein Ab|Myelin associated glycoprotein Ab
C3172468|T201|COMP|63397-4|LNC|Myeloperoxidase Ab|Myeloperoxidase Ab
C3172469|T201|COMP|63398-2|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C3172470|T201|COMP|63399-0|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C3172471|T201|COMP|63400-6|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C3172472|T201|COMP|63401-4|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C3172473|T201|COMP|63402-2|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C3172474|T201|COMP|63403-0|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C3172475|T201|COMP|63404-8|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C3172476|T201|COMP|63405-5|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C3172477|T201|COMP|63406-3|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C3172478|T201|COMP|63407-1|LNC|Thyroid colloidal Ab|Thyroid colloidal Ab
C3172479|T201|COMP|63408-9|LNC|DNA double strand Ab|DNA double strand Ab
C3172480|T201|COMP|63409-7|LNC|DNA double strand Ab|DNA double strand Ab
C3172481|T201|COMP|63410-5|LNC|DNA double strand Ab|DNA double strand Ab
C3172482|T201|COMP|63411-3|LNC|Sjogrens syndrome-A extractable nuclear 60kD Ab|Sjogrens syndrome-A extractable nuclear 60kD Ab
C3172483|T201|COMP|63412-1|LNC|Thyroid colloidal Ab|Thyroid colloidal Ab
C3172484|T201|COMP|63413-9|LNC|Thyroid colloidal Ab|Thyroid colloidal Ab
C3172485|T201|COMP|63414-7|LNC|Pompe disease newborn screening panel|Pompe disease newborn screening panel
C3172486|T201|COMP|63415-4|LNC|Pompe disease|Pompe disease
C3172490|T201|COMP|63418-8|LNC|Lactalbumin alpha Ab.IgG|Lactalbumin alpha Ab.IgG
C3172491|T201|COMP|63419-6|LNC|PIK3CA gene mutations tested for|PIK3CA gene mutations tested for
C3172495|T201|COMP|63421-2|LNC|JAK2 gene exon 12 mutations tested for|JAK2 gene exon 12 mutations tested for
C3172499|T201|COMP|63423-8|LNC|Escherichia coli eaeA gene|Escherichia coli eaeA gene
C3172501|T201|COMP|63424-6|LNC|Bacterial enterohemolysin (ehlyA) gene|Bacterial enterohemolysin (ehlyA) gene
C3172503|T201|COMP|63425-3|LNC|Bacterial heat-labile enterotoxin LT gene|Bacterial heat-labile enterotoxin LT gene
C3172505|T201|COMP|63426-1|LNC|Bacterial heat-stable enterotoxin ST gene|Bacterial heat-stable enterotoxin ST gene
C3172507|T201|COMP|63427-9|LNC|Escherichia coli Stx1 toxin stx1 gene|Escherichia coli Stx1 toxin stx1 gene
C3172509|T201|COMP|63428-7|LNC|Escherichia coli Stx2 toxin stx2 gene|Escherichia coli Stx2 toxin stx2 gene
C3172511|T201|COMP|63429-5|LNC|Bacterial beta-glucuronidase (uidA) gene|Bacterial beta-glucuronidase (uidA) gene
C3172513|T201|COMP|63430-3|LNC|Human coronavirus RNA panel|Human coronavirus RNA panel
C3172515|T201|COMP|63431-1|LNC|Bordetella sp DNA|Bordetella sp DNA
C3172516|T201|COMP|63432-9|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C3172518|T201|COMP|63434-5|LNC|Coxsackievirus A Ab|Coxsackievirus A Ab
C3172519|T201|COMP|63435-2|LNC|Brucella abortus Ab|Brucella abortus Ab
C3172520|T201|COMP|63436-0|LNC|Polistes spp recombinant (rPol d) 5 Ab.IgE|Polistes spp recombinant (rPol d) 5 Ab.IgE
C3172522|T201|COMP|63437-8|LNC|Brucella abortus Ab|Brucella abortus Ab
C3172523|T201|COMP|63438-6|LNC|MAPT gene mutations tested for|MAPT gene mutations tested for
C3172525|T201|COMP|63439-4|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C3172526|T201|COMP|63440-2|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C3172527|T201|COMP|63441-0|LNC|Tissue polypeptide Ag|Tissue polypeptide Ag
C3172528|T201|COMP|63443-6|LNC|Fasciola hepatica Ab|Fasciola hepatica Ab
C3172529|T201|COMP|63444-4|LNC|Somatotropin^7H post XXX challenge|Somatotropin^7H post XXX challenge
C3172530|T201|COMP|63445-1|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C3172531|T201|COMP|63446-9|LNC|Cells.CD3+CD5-/100 cells|Cells.CD3+CD5-/100 cells
C3172533|T201|COMP|63447-7|LNC|Cells.CD3+CD5-|Cells.CD3+CD5-
C3172535|T201|COMP|63448-5|LNC|Cells.CD3+CD5+/100 cells|Cells.CD3+CD5+/100 cells
C3172537|T201|COMP|63465-9|LNC|Brucella sp DNA|Brucella sp DNA
C3172538|T201|COMP|63466-7|LNC|Ganglioside GM3 Ab.IgG|Ganglioside GM3 Ab.IgG
C3172539|T201|COMP|63467-5|LNC|Ganglioside GM3 Ab.IgM|Ganglioside GM3 Ab.IgM
C3172540|T201|COMP|63468-3|LNC|Ganglioside GT1a Ab.IgG|Ganglioside GT1a Ab.IgG
C3172541|T201|COMP|63469-1|LNC|Ganglioside GT1b Ab.IgG|Ganglioside GT1b Ab.IgG
C3172542|T201|COMP|63478-2|LNC|Platelet glycoprotein Ib-Ix Ab|Platelet glycoprotein Ib-Ix Ab
C3172543|T201|COMP|63479-0|LNC|Platelet glycoprotein Ia-IIa Ab|Platelet glycoprotein Ia-IIa Ab
C3172545|T201|COMP|63481-6|LNC|Urea|Urea
C3172546|T201|COMP|63482-4|LNC|Methotrimeprazine|Methotrimeprazine
C3172547|T201|COMP|63483-2|LNC|Penicillium notatum Ab|Penicillium notatum Ab
C3172548|T201|COMP|63484-0|LNC|Actin.filamentous Ab|Actin.filamentous Ab
C3172551|T201|COMP|63486-5|LNC|Nut allergen panel|Nut allergen panel
C3172553|T201|COMP|63487-3|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C3172554|T201|COMP|63488-1|LNC|Epithelial cells.ciliated|Epithelial cells.ciliated
C3172589|T201|COMP|63523-5|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C3172590|T201|COMP|63524-3|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C3172591|T201|COMP|63526-8|LNC|Centromere Ab|Centromere Ab
C3172592|T201|COMP|63527-6|LNC|Centromere Ab|Centromere Ab
C3172593|T201|COMP|63528-4|LNC|Centromere Ab|Centromere Ab
C3172594|T201|COMP|63529-2|LNC|Centromere Ab|Centromere Ab
C3172595|T201|COMP|63530-0|LNC|Centromere Ab|Centromere Ab
C3172596|T201|COMP|63531-8|LNC|Centromere Ab|Centromere Ab
C3172597|T201|COMP|63532-6|LNC|Centromere protein B Ab|Centromere protein B Ab
C3172598|T201|COMP|63533-4|LNC|Centromere protein B Ab|Centromere protein B Ab
C3172599|T201|COMP|63534-2|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172600|T201|COMP|63535-9|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3172601|T201|COMP|63536-7|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C3172602|T201|COMP|63537-5|LNC|Muscle specific receptor tyrosine kinase Ab.IgG|Muscle specific receptor tyrosine kinase Ab.IgG
C3172604|T201|COMP|63538-3|LNC|Myeloperoxidase Ab|Myeloperoxidase Ab
C3172605|T201|COMP|63539-1|LNC|Proteinase 3 Ab|Proteinase 3 Ab
C3172606|T201|COMP|63540-9|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C3172607|T201|COMP|63541-7|LNC|Ribosomal P Ab|Ribosomal P Ab
C3172608|T201|COMP|63542-5|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C3172609|T201|COMP|63543-3|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C3172610|T201|COMP|63544-1|LNC|Sjogrens syndrome-A extractable nuclear 60kD Ab|Sjogrens syndrome-A extractable nuclear 60kD Ab
C3172611|T201|COMP|63545-8|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C3172612|T201|COMP|63546-6|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C3172614|T201|COMP|63548-2|LNC|Smith extractable nuclear B Ab|Smith extractable nuclear B Ab
C3172615|T201|COMP|63549-0|LNC|Albumin.serum-Albumin.periton fld|Albumin.serum-Albumin.periton fld
C3172616|T201|COMP|63551-6|LNC|Pituitary Ab|Pituitary Ab
C3172617|T201|COMP|63552-4|LNC|Macrophages/100 cells|Macrophages/100 cells
C3172619|T201|COMP|63553-2|LNC|Succinylaminoimidazole carboxamide riboside|Succinylaminoimidazole carboxamide riboside
C3172620|T201|COMP|63554-0|LNC|Leukocytes|Leukocytes
C3172621|T201|COMP|63555-7|LNC|Leukocytes|Leukocytes
C3172623|T201|COMP|63557-3|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C3172624|T201|COMP|63558-1|LNC|HLA-DQB1*06:02|HLA-DQB1*06:02
C3172625|T201|COMP|63559-9|LNC|Signal recognition particle Ab|Signal recognition particle Ab
C3172626|T201|COMP|63560-7|LNC|Somatotropin^8.5H post XXX challenge|Somatotropin^8.5H post XXX challenge
C3172627|T201|COMP|63561-5|LNC|Coagulation surface induced actual/Normal|Coagulation surface induced actual/Normal
C3172629|T201|COMP|63562-3|LNC|Japanese encephalitis virus Ab.IgM|Japanese encephalitis virus Ab.IgM
C3172630|T201|COMP|63563-1|LNC|Japanese encephalitis virus Ab.IgM|Japanese encephalitis virus Ab.IgM
C3172633|T201|COMP|63565-6|LNC|Prothionamide|Prothionamide
C3172634|T201|COMP|63566-4|LNC|Basement membrane Ab pattern|Basement membrane Ab pattern
C3172636|T201|COMP|63567-2|LNC|Neutrophil cytoplasmic Ab pattern|Neutrophil cytoplasmic Ab pattern
C3172637|T201|COMP|63568-0|LNC|Neutrophil cytoplasmic Ab pattern|Neutrophil cytoplasmic Ab pattern
C3173208|T201|COMP|64233-0|LNC|Benzylpiperazine|Benzylpiperazine
C3173232|T201|COMP|64966-5|LNC|Triticum aestivum recombinant (rTri a) 14 Ab.IgE|Triticum aestivum recombinant (rTri a) 14 Ab.IgE
C3173234|T201|COMP|64967-3|LNC|Alnus glutinosa recombinant (rAln g) 1 Ab.IgE|Alnus glutinosa recombinant (rAln g) 1 Ab.IgE
C3173238|T201|COMP|64969-9|LNC|Platanus acerifolia recombinant (rPla a) 1 Ab.IgE|Platanus acerifolia recombinant (rPla a) 1 Ab.IgE
C3173240|T201|COMP|64970-7|LNC|Platanus acerifolia recombinant (rPla a) 3 Ab.IgE|Platanus acerifolia recombinant (rPla a) 3 Ab.IgE
C3173242|T201|COMP|64971-5|LNC|Chenopodium album recombinant (rChe a) 1 Ab.IgE|Chenopodium album recombinant (rChe a) 1 Ab.IgE
C3173438|T201|COMP|64012-8|LNC|CEBPA gene targeted mutation analysis|CEBPA gene targeted mutation analysis
C3173440|T201|COMP|64013-6|LNC|Escherichia coli shiga-like toxin 1 & 2|Escherichia coli shiga-like toxin 1 & 2
C3173462|T201|COMP|64038-3|LNC|Adenovirus DNA|Adenovirus DNA
C3173542|T201|COMP|64081-3|LNC|Cells.FMRP/100 lymphocytes|Cells.FMRP/100 lymphocytes
C3173544|T201|COMP|64082-1|LNC|Bilirubin.non-glucuronidated|Bilirubin.non-glucuronidated
C3173545|T201|COMP|64083-9|LNC|MGMT gene methylation score|MGMT gene methylation score
C3173548|T201|COMP|64085-4|LNC|Cells karyotyped.total|Cells karyotyped.total
C3173549|T201|COMP|64086-2|LNC|Cells analyzed|Cells analyzed
C3173550|T201|COMP|64087-0|LNC|ISCN band level|ISCN band level
C3173551|T201|COMP|64088-8|LNC|Karyotype|Karyotype
C3173552|T201|COMP|64089-6|LNC|Cells counted|Cells counted
C3173553|T201|COMP|64090-4|LNC|Chromosome analysis overall interpretation|Chromosome analysis overall interpretation
C3173554|T201|COMP|64091-2|LNC|Cells karyotyped.total|Cells karyotyped.total
C3173555|T201|COMP|64092-0|LNC|Cells analyzed|Cells analyzed
C3173556|T201|COMP|64093-8|LNC|ISCN band level|ISCN band level
C3173557|T201|COMP|64094-6|LNC|Karyotype|Karyotype
C3173558|T201|COMP|64095-3|LNC|Cells counted|Cells counted
C3173559|T201|COMP|64096-1|LNC|Colonies counted|Colonies counted
C3173581|T201|COMP|64116-7|LNC|Hemoglobin observations newborn screening panel|Hemoglobin observations newborn screening panel
C3173583|T201|COMP|64117-5|LNC|Most predominant hemoglobin|Most predominant hemoglobin
C3173585|T201|COMP|64118-3|LNC|Second most predominant hemoglobin|Second most predominant hemoglobin
C3173586|T201|COMP|64119-1|LNC|Third most predominant hemoglobin|Third most predominant hemoglobin
C3173587|T201|COMP|64120-9|LNC|Fourth most predominant hemoglobin|Fourth most predominant hemoglobin
C3173589|T201|COMP|64121-7|LNC|Fifth most predominant hemoglobin|Fifth most predominant hemoglobin
C3173597|T201|COMP|64125-8|LNC|Pregabalin|Pregabalin
C3173598|T201|COMP|64126-6|LNC|Drugs identified|Drugs identified
C3173599|T201|COMP|64127-4|LNC|Methylenedioxyethylamphetamine/Creatinine|Methylenedioxyethylamphetamine/Creatinine
C3173601|T201|COMP|64128-2|LNC|Amobarbital/Creatinine|Amobarbital/Creatinine
C3173603|T201|COMP|64129-0|LNC|N-desalkylflurazepam/Creatinine|N-desalkylflurazepam/Creatinine
C3173605|T201|COMP|64130-8|LNC|diazePAM/Creatinine|diazePAM/Creatinine
C3173607|T201|COMP|64131-6|LNC|Dihydrocodeine/Creatinine|Dihydrocodeine/Creatinine
C3173609|T201|COMP|64132-4|LNC|PENTobarbital/Creatinine|PENTobarbital/Creatinine
C3173611|T201|COMP|64133-2|LNC|PHENobarbital/Creatinine|PHENobarbital/Creatinine
C3173613|T201|COMP|64134-0|LNC|Phentermine/Creatinine|Phentermine/Creatinine
C3173615|T201|COMP|64135-7|LNC|Secobarbital/Creatinine|Secobarbital/Creatinine
C3173617|T201|COMP|64136-5|LNC|Pregabalin/Creatinine|Pregabalin/Creatinine
C3173619|T201|COMP|64137-3|LNC|Pregabalin|Pregabalin
C3173620|T201|COMP|64138-1|LNC|Methylenedioxyamphetamine/Creatinine|Methylenedioxyamphetamine/Creatinine
C3173622|T201|COMP|64139-9|LNC|Butalbital/Creatinine|Butalbital/Creatinine
C3173950|T201|COMP|64412-0|LNC|Mycobacterium sp|Mycobacterium sp
C3173951|T201|COMP|64423-7|LNC|KIR2DS4 gene full variant|KIR2DS4 gene full variant
C3173953|T201|COMP|64424-5|LNC|KIR2DS4 gene deletion variant|KIR2DS4 gene deletion variant
C3173955|T201|COMP|64425-2|LNC|KIR gene allele 2DS5|KIR gene allele 2DS5
C3173957|T201|COMP|64426-0|LNC|KIR gene allele 3DL1|KIR gene allele 3DL1
C3173959|T201|COMP|64427-8|LNC|KIR gene allele 3DL2|KIR gene allele 3DL2
C3173961|T201|COMP|64428-6|LNC|KIR gene allele 3DL3|KIR gene allele 3DL3
C3173963|T201|COMP|64429-4|LNC|KIR gene allele 3DS1|KIR gene allele 3DS1
C3173965|T201|COMP|64430-2|LNC|KIR gene allele 2DP1|KIR gene allele 2DP1
C3173967|T201|COMP|64431-0|LNC|KIR3DP1 gene full variant|KIR3DP1 gene full variant
C3173969|T201|COMP|64432-8|LNC|KIR3DP1 gene deletion variant|KIR3DP1 gene deletion variant
C3173971|T201|COMP|64433-6|LNC|Fragile X protein (FMRP) panel|Fragile X protein (FMRP) panel
C3174140|T201|COMP|64986-3|LNC|Anisakis simplex recombinant (rAni s) 3 Ab.IgE|Anisakis simplex recombinant (rAni s) 3 Ab.IgE
C3174192|T201|COMP|65360-0|LNC|Thyrotropin^pre or post XXX challenge|Thyrotropin^pre or post XXX challenge
C3174193|T201|COMP|65361-8|LNC|Phenytoin^^corrected for albumin|Phenytoin^^corrected for albumin
C3174194|T201|COMP|65362-6|LNC|Magnesium^^corrected for albumin|Magnesium^^corrected for albumin
C3174195|T201|COMP|65363-4|LNC|Glutathione|Glutathione
C3174196|T201|COMP|65364-2|LNC|Cortisol.free/Cortisol.total|Cortisol.free/Cortisol.total
C3174348|T201|COMP|65789-0|LNC|Mouse lipocain native (nMus m) 1 Ab.IgE|Mouse lipocain native (nMus m) 1 Ab.IgE
C3174350|T201|COMP|65790-8|LNC|Dermatophagoides farinae native (nDer f) 1 Ab.IgE|Dermatophagoides farinae native (nDer f) 1 Ab.IgE
C3174352|T201|COMP|65791-6|LNC|Apis mellifera native (nApi m) 4 Ab.IgE|Apis mellifera native (nApi m) 4 Ab.IgE
C3174354|T201|COMP|65792-4|LNC|Armoracia rusticana native (nArm r) HRP Ab.IgE|Armoracia rusticana native (nArm r) HRP Ab.IgE
C3174356|T201|COMP|65793-2|LNC|Blatella germanica native (nBla g) 7 Ab.IgE|Blatella germanica native (nBla g) 7 Ab.IgE
C3174358|T201|COMP|65794-0|LNC|Penaeus monodon native (nPen m) 1 Ab.IgE|Penaeus monodon native (nPen m) 1 Ab.IgE
C3174360|T201|COMP|65795-7|LNC|Actinidia deliciosa native (nAct d) 1 Ab.IgE|Actinidia deliciosa native (nAct d) 1 Ab.IgE
C3174362|T201|COMP|65796-5|LNC|Actinidia deliciosa native (nAct d) 2 Ab.IgE|Actinidia deliciosa native (nAct d) 2 Ab.IgE
C3174658|T201|COMP|65750-2|LNC|Drugs of abuse 5 panel|Drugs of abuse 5 panel
C3174659|T201|COMP|65751-0|LNC|Pathology biopsy report|Pathology biopsy report
C3174660|T201|COMP|65752-8|LNC|Pathology biopsy report|Pathology biopsy report
C3174661|T201|COMP|65753-6|LNC|Pathology biopsy report|Pathology biopsy report
C3174662|T201|COMP|65754-4|LNC|Pathology biopsy report|Pathology biopsy report
C3174663|T201|COMP|65755-1|LNC|Pathology biopsy report|Pathology biopsy report
C3174664|T201|COMP|65757-7|LNC|Pathology biopsy report|Pathology biopsy report
C3174665|T201|COMP|65758-5|LNC|T-cell helper (CD4) subset panel|T-cell helper (CD4) subset panel
C3174853|T201|COMP|64797-4|LNC|Oxygen content|Oxygen content
C3174854|T201|COMP|64798-2|LNC|Oxygen content|Oxygen content
C3174855|T201|COMP|64799-0|LNC|Oxygen content|Oxygen content
C3174856|T201|COMP|64800-6|LNC|Oxygen content|Oxygen content
C3175084|T201|COMP|64959-0|LNC|Actinidia deliciosa recombinant (rAct d) 8 Ab.IgE|Actinidia deliciosa recombinant (rAct d) 8 Ab.IgE
C3175086|T201|COMP|64960-8|LNC|Apium graveolens recombinant (rApi g) 1 Ab.IgE|Apium graveolens recombinant (rApi g) 1 Ab.IgE
C3175088|T201|COMP|64961-6|LNC|Malus domestica recombinant (rMal d) 1 Ab.IgE|Malus domestica recombinant (rMal d) 1 Ab.IgE
C3175151|T201|COMP|64965-7|LNC|Arachis hypogaea recombinant (rAra h) 9 Ab.IgE|Arachis hypogaea recombinant (rAra h) 9 Ab.IgE
C3175153|T201|COMP|64972-3|LNC|Plantago lanceolata recombinant (rPla l) 1 Ab.IgE|Plantago lanceolata recombinant (rPla l) 1 Ab.IgE
C3175155|T201|COMP|64973-1|LNC|Dog recombinant (rCan f) 5 Ab.IgE|Dog recombinant (rCan f) 5 Ab.IgE
C3175157|T201|COMP|64974-9|LNC|Horse recombinant (rEqu c) 1 Ab.IgE|Horse recombinant (rEqu c) 1 Ab.IgE
C3175159|T201|COMP|64975-6|LNC|Cat recombinant (rFel d) 1 Ab.IgE|Cat recombinant (rFel d) 1 Ab.IgE
C3175161|T201|COMP|64976-4|LNC|Cat recombinant (rFel d) 4 Ab.IgE|Cat recombinant (rFel d) 4 Ab.IgE
C3175167|T201|COMP|64979-8|LNC|Blomia tropicalis recombinant (rBlo t) 5 Ab.IgE|Blomia tropicalis recombinant (rBlo t) 5 Ab.IgE
C3175173|T201|COMP|64982-2|LNC|Blatella germanica recombinant (rBla g) 1 Ab.IgE|Blatella germanica recombinant (rBla g) 1 Ab.IgE
C3175175|T201|COMP|64983-0|LNC|Blatella germanica recombinant (rBla g) 2 Ab.IgE|Blatella germanica recombinant (rBla g) 2 Ab.IgE
C3175177|T201|COMP|64984-8|LNC|Blatella germanica recombinant (rBla g) 5 Ab.IgE|Blatella germanica recombinant (rBla g) 5 Ab.IgE
C3175179|T201|COMP|64985-5|LNC|Anisakis simplex recombinant (rAni s) 1 Ab.IgE|Anisakis simplex recombinant (rAni s) 1 Ab.IgE
C3175662|T201|COMP|65318-8|LNC|A little t super little a Ab|A little t super little a Ab
C3175664|T201|COMP|65319-6|LNC|D little u super little a Ab|D little u super little a Ab
C3175666|T201|COMP|65320-4|LNC|F little y3 Ab|F little y3 Ab
C3175668|T201|COMP|65321-2|LNC|G little e Ab|G little e Ab
C3175670|T201|COMP|65322-0|LNC|G little y super little a Ab|G little y super little a Ab
C3175672|T201|COMP|65323-8|LNC|H little e Ab|H little e Ab
C3175674|T201|COMP|65324-6|LNC|J little k3 Ab|J little k3 Ab
C3175676|T201|COMP|65325-3|LNC|K little u Ab|K little u Ab
C3175677|T201|COMP|65326-1|LNC|LAN Ab|LAN Ab
C3175679|T201|COMP|65327-9|LNC|L little u 14 Ab|L little u 14 Ab
C3175681|T201|COMP|65328-7|LNC|LW super little a Ab|LW super little a Ab
C3175683|T201|COMP|65329-5|LNC|M little c C super little c Ab|M little c C super little c Ab
C3175685|T201|COMP|65330-3|LNC|MER Ab|MER Ab
C3175687|T201|COMP|65331-1|LNC|little c E Ab|little c E Ab
C3175689|T201|COMP|65332-9|LNC|Rh32 Ab|Rh32 Ab
C3175690|T201|COMP|65333-7|LNC|S little c super 1 Ab|S little c super 1 Ab
C3175691|T201|COMP|65334-5|LNC|S little c super 2 Ab|S little c super 2 Ab
C3175692|T201|COMP|65335-2|LNC|S little w super little a Ab|S little w super little a Ab
C3175693|T201|COMP|65336-0|LNC|T little m Ab|T little m Ab
C3175694|T201|COMP|65337-8|LNC|T little r super little a Ab|T little r super little a Ab
C3175695|T201|COMP|65338-6|LNC|WES super little b Ab|WES super little b Ab
C3175696|T201|COMP|65339-4|LNC|W little r super little b Ab|W little r super little b Ab
C3175697|T201|COMP|65340-2|LNC|Micafungin|Micafungin
C3175698|T201|COMP|65343-6|LNC|Oxygen^^saturation adjusted to 0.5|Oxygen^^saturation adjusted to 0.5
C3175699|T201|COMP|65344-4|LNC|Glucagon^pre XXX challenge|Glucagon^pre XXX challenge
C3175700|T201|COMP|65345-1|LNC|Glucagon^1st specimen post XXX challenge|Glucagon^1st specimen post XXX challenge
C3175701|T201|COMP|65346-9|LNC|Glucagon^2nd specimen post XXX challenge|Glucagon^2nd specimen post XXX challenge
C3175702|T201|COMP|65347-7|LNC|Glucagon^3rd specimen post XXX challenge|Glucagon^3rd specimen post XXX challenge
C3175703|T201|COMP|65348-5|LNC|Glucagon^4th specimen post XXX challenge|Glucagon^4th specimen post XXX challenge
C3175704|T201|COMP|65349-3|LNC|Glucagon^5th specimen post XXX challenge|Glucagon^5th specimen post XXX challenge
C3175705|T201|COMP|65350-1|LNC|Follitropin^pre or post XXX challenge|Follitropin^pre or post XXX challenge
C3175706|T201|COMP|65351-9|LNC|Triiodothyronine.free^pre or post XXX challenge|Triiodothyronine.free^pre or post XXX challenge
C3175707|T201|COMP|65352-7|LNC|Proinsulin^1st specimen post XXX challenge|Proinsulin^1st specimen post XXX challenge
C3175708|T201|COMP|65353-5|LNC|Proinsulin^2nd specimen post XXX challenge|Proinsulin^2nd specimen post XXX challenge
C3175709|T201|COMP|65354-3|LNC|Proinsulin^3rd specimen post XXX challenge|Proinsulin^3rd specimen post XXX challenge
C3175710|T201|COMP|65355-0|LNC|Proinsulin^4th specimen post XXX challenge|Proinsulin^4th specimen post XXX challenge
C3175711|T201|COMP|65356-8|LNC|Proinsulin^5th specimen post XXX challenge|Proinsulin^5th specimen post XXX challenge
C3175712|T201|COMP|65357-6|LNC|Proinsulin^6th specimen post XXX challenge|Proinsulin^6th specimen post XXX challenge
C3175713|T201|COMP|65358-4|LNC|Proinsulin^7th specimen post XXX challenge|Proinsulin^7th specimen post XXX challenge
C3176084|T201|COMP|65632-2|LNC|Clozapine & Norclozapine panel|Clozapine & Norclozapine panel
C3176086|T201|COMP|65633-0|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C3176087|T201|COMP|65634-8|LNC|Creatinine 24 hour urine panel|Creatinine 24 hour urine panel
C3176244|T201|COMP|65759-3|LNC|T-cell subsets CD4 & CD8 panel|T-cell subsets CD4 & CD8 panel
C3176245|T201|COMP|65761-9|LNC|Lymphocyte subset interpretation|Lymphocyte subset interpretation
C3176247|T201|COMP|65762-7|LNC|Hantavirus Ag|Hantavirus Ag
C3176249|T201|COMP|65763-5|LNC|Neisseria meningitidis Ag|Neisseria meningitidis Ag
C3176250|T201|COMP|65764-3|LNC|Actinidia deliciosa native (nAct d) 5 Ab.IgE|Actinidia deliciosa native (nAct d) 5 Ab.IgE
C3176252|T201|COMP|65765-0|LNC|Corylus avellana native (nCor a) 9 Ab.IgE|Corylus avellana native (nCor a) 9 Ab.IgE
C3176254|T201|COMP|65766-8|LNC|Juglans regia native (nJug r) 1 Ab.IgE|Juglans regia native (nJug r) 1 Ab.IgE
C3176256|T201|COMP|65767-6|LNC|Juglans regia native (nJug r) 2 Ab.IgE|Juglans regia native (nJug r) 2 Ab.IgE
C3176258|T201|COMP|65768-4|LNC|Juglans regia native (nJug r) 3 Ab.IgE|Juglans regia native (nJug r) 3 Ab.IgE
C3176260|T201|COMP|65769-2|LNC|Arachis hypogaea native (nAra h) 1 Ab.IgE|Arachis hypogaea native (nAra h) 1 Ab.IgE
C3176262|T201|COMP|65770-0|LNC|Arachis hypogaea native (nAra h) 2 Ab.IgE|Arachis hypogaea native (nAra h) 2 Ab.IgE
C3176264|T201|COMP|65771-8|LNC|Arachis hypogaea native (nAra h) 3 Ab.IgE|Arachis hypogaea native (nAra h) 3 Ab.IgE
C3176266|T201|COMP|65772-6|LNC|Glycine max native (nGly m) 6 Ab.IgE|Glycine max native (nGly m) 6 Ab.IgE
C3176268|T201|COMP|65773-4|LNC|Fagopyrum esculentum native (nFag e) 2 Ab.IgE|Fagopyrum esculentum native (nFag e) 2 Ab.IgE
C3176270|T201|COMP|65774-2|LNC|Triticum aestivum native (nTri a) aA_TI Ab.IgE|Triticum aestivum native (nTri a) aA_TI Ab.IgE
C3176272|T201|COMP|65775-9|LNC|Cynodon dactylon native (nCyn d) 1 Ab.IgE|Cynodon dactylon native (nCyn d) 1 Ab.IgE
C3176274|T201|COMP|65776-7|LNC|Betula verrucosa native (nBet v) 1 Ab.IgE|Betula verrucosa native (nBet v) 1 Ab.IgE
C3176276|T201|COMP|65777-5|LNC|Cryptomeria japonica native (nCry j) 1 Ab.IgE|Cryptomeria japonica native (nCry j) 1 Ab.IgE
C3176278|T201|COMP|65778-3|LNC|Cupressus arizonica native (nCup a) 1 Ab.IgE|Cupressus arizonica native (nCup a) 1 Ab.IgE
C3176280|T201|COMP|65779-1|LNC|Olea europaea native (nOle e) 7 Ab.IgE|Olea europaea native (nOle e) 7 Ab.IgE
C3176282|T201|COMP|65780-9|LNC|Olea europaea recombinant (rOle e) 9 Ab.IgE|Olea europaea recombinant (rOle e) 9 Ab.IgE
C3176284|T201|COMP|65781-7|LNC|Platanus acerifolia native (nPla a) 2 Ab.IgE|Platanus acerifolia native (nPla a) 2 Ab.IgE
C3176286|T201|COMP|65782-5|LNC|Ambrosia artemisiifolia native (nAmb a) 1 Ab.IgE|Ambrosia artemisiifolia native (nAmb a) 1 Ab.IgE
C3176288|T201|COMP|65783-3|LNC|Artemisia vulgaris native (nArt v) 3 Ab.IgE|Artemisia vulgaris native (nArt v) 3 Ab.IgE
C3176290|T201|COMP|65784-1|LNC|Salsola kali native (nSal k) 1 Ab.IgE|Salsola kali native (nSal k) 1 Ab.IgE
C3176294|T201|COMP|65786-6|LNC|Penaeus monodon native (nPen m) 2 Ab.IgE|Penaeus monodon native (nPen m) 2 Ab.IgE
C3176296|T201|COMP|65787-4|LNC|Penaeus monodon native (nPen m) 4 Ab.IgE|Penaeus monodon native (nPen m) 4 Ab.IgE
C3176298|T201|COMP|65788-2|LNC|Horse serum albumin native (nEqu c) 3 Ab.IgE|Horse serum albumin native (nEqu c) 3 Ab.IgE
C3176300|T201|COMP|65807-0|LNC|Tapentadol|Tapentadol
C3176301|T201|COMP|65808-8|LNC|Nortapentadol|Nortapentadol
C3176303|T201|COMP|65809-6|LNC|Kingella kingae DNA|Kingella kingae DNA
C3176305|T201|COMP|65810-4|LNC|SEPT9 gene methylation|SEPT9 gene methylation
C3176316|T201|COMP|65818-7|LNC|Medication XXX|Medication XXX
C3176355|T201|COMP|65844-3|LNC|Date of observation|Date of observation
C3176378|T201|COMP|65866-6|LNC|Methacholine|Methacholine
C3202994|T201|COMP|7518-4|LNC|Cucumis melo spp Ab.IgE|Cucumis melo spp Ab.IgE
C3202995|T201|COMP|7176-1|LNC|Cucumis melo spp Ab.IgG|Cucumis melo spp Ab.IgG
C3202996|T201|COMP|15600-0|LNC|Cucumis melo spp Ab.IgE.RAST class|Cucumis melo spp Ab.IgE.RAST class
C3202997|T201|COMP|6172-1|LNC|Cucumis melo spp Ab.IgE|Cucumis melo spp Ab.IgE
C3202998|T201|COMP|7175-3|LNC|Cucumis melo spp Ab.IgE|Cucumis melo spp Ab.IgE
C3258478|T201|COMP|62201-9|LNC|XXX microorganism DNA|XXX microorganism DNA
C3258479|T201|COMP|62202-7|LNC|XXX microorganism DNA|XXX microorganism DNA
C3258483|T201|COMP|61099-8|LNC|Collection date^3rd specimen|Collection date^3rd specimen
C3258484|T201|COMP|61100-4|LNC|Collection date^2nd specimen|Collection date^2nd specimen
C3258818|T201|COMP|63550-8|LNC|Calcium magnesium phosphate/Total|Calcium magnesium phosphate/Total
C3258825|T201|COMP|66143-9|LNC|Monocytes|Monocytes
C3258826|T201|COMP|66144-7|LNC|Lymphocytes.variant|Lymphocytes.variant
C3258827|T201|COMP|66145-4|LNC|Leukocytes other|Leukocytes other
C3258828|T201|COMP|66146-2|LNC|Reticulocytes|Reticulocytes
C3258829|T201|COMP|66147-0|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C3258830|T201|COMP|66148-8|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C3258848|T201|COMP|66130-6|LNC|Fentanyl+Norfentanyl|Fentanyl+Norfentanyl
C3258849|T201|COMP|66131-4|LNC|Norbuprenorphine|Norbuprenorphine
C3258850|T201|COMP|66132-2|LNC|Mononuclear+Mesothelial cells/100 leukocytes|Mononuclear+Mesothelial cells/100 leukocytes
C3258852|T201|COMP|66133-0|LNC|Mononuclear cells.atypical/100 leukocytes|Mononuclear cells.atypical/100 leukocytes
C3258854|T201|COMP|66134-8|LNC|Blasts|Blasts
C3258855|T201|COMP|66135-5|LNC|Promyelocytes|Promyelocytes
C3258856|T201|COMP|66136-3|LNC|Myelocytes|Myelocytes
C3258879|T201|COMP|65756-9|LNC|Salmonella sp serovar|Salmonella sp serovar
C3258882|T201|COMP|66107-4|LNC|Pathology biopsy report|Pathology biopsy report
C3258883|T201|COMP|66108-2|LNC|Pathology biopsy report|Pathology biopsy report
C3258884|T201|COMP|66109-0|LNC|Pathology biopsy report|Pathology biopsy report
C3258885|T201|COMP|66110-8|LNC|Pathology biopsy report|Pathology biopsy report
C3258886|T201|COMP|66111-6|LNC|Pathology biopsy report|Pathology biopsy report
C3258887|T201|COMP|66112-4|LNC|Pathology biopsy report|Pathology biopsy report
C3258888|T201|COMP|66113-2|LNC|Pathology biopsy report|Pathology biopsy report
C3258889|T201|COMP|66114-0|LNC|Pathology biopsy report|Pathology biopsy report
C3258890|T201|COMP|66115-7|LNC|Pathology biopsy report|Pathology biopsy report
C3258891|T201|COMP|66116-5|LNC|Pathology biopsy report|Pathology biopsy report
C3258892|T201|COMP|66117-3|LNC|Pathology biopsy report|Pathology biopsy report
C3258893|T201|COMP|66118-1|LNC|Pathology biopsy report|Pathology biopsy report
C3258894|T201|COMP|66119-9|LNC|Pathology biopsy report|Pathology biopsy report
C3258895|T201|COMP|66120-7|LNC|Pathology biopsy report|Pathology biopsy report
C3258896|T201|COMP|66121-5|LNC|Pathology biopsy report|Pathology biopsy report
C3258897|T201|COMP|66122-3|LNC|Pathology biopsy report|Pathology biopsy report
C3258898|T201|COMP|66123-1|LNC|Pathology biopsy report|Pathology biopsy report
C3258899|T201|COMP|66124-9|LNC|Pathology biopsy report|Pathology biopsy report
C3258900|T201|COMP|66125-6|LNC|Pathology biopsy report|Pathology biopsy report
C3258901|T201|COMP|66126-4|LNC|Cholesterol.in VLDL|Cholesterol.in VLDL
C3258902|T201|COMP|66127-2|LNC|Amphetamine|Amphetamine
C3258903|T201|COMP|66128-0|LNC|chlordiazePOXIDE/Creatinine|chlordiazePOXIDE/Creatinine
C3258905|T201|COMP|66129-8|LNC|Fentanyl+Norfentanyl|Fentanyl+Norfentanyl
C3258969|T201|COMP|66137-1|LNC|Metamyelocytes|Metamyelocytes
C3258970|T201|COMP|66138-9|LNC|Neutrophils.band form|Neutrophils.band form
C3258971|T201|COMP|66139-7|LNC|Neutrophils|Neutrophils
C3258972|T201|COMP|66140-5|LNC|Lymphocytes|Lymphocytes
C3258973|T201|COMP|66141-3|LNC|Eosinophils|Eosinophils
C3258974|T201|COMP|66142-1|LNC|Basophils|Basophils
C3258979|T201|COMP|66481-3|LNC|Protein.monoclonal band 2|Protein.monoclonal band 2
C3258980|T201|COMP|66482-1|LNC|OmpC Ab.IgA|OmpC Ab.IgA
C3258981|T201|COMP|66483-9|LNC|Heparin.unfractionated|Heparin.unfractionated
C3258982|T201|COMP|66484-7|LNC|DNA single strand Ab|DNA single strand Ab
C3258983|T201|COMP|66485-4|LNC|Brucella sp Ab.IgG & IgM|Brucella sp Ab.IgG & IgM
C3258985|T201|COMP|66884-8|LNC|Skin Ab.IgG pattern|Skin Ab.IgG pattern
C3258986|T201|COMP|66885-5|LNC|Bacterial 16S rRNA sequencing|Bacterial 16S rRNA sequencing
C3259279|T201|COMP|66441-7|LNC|Beta hydroxybutyrate|Beta hydroxybutyrate
C3259280|T201|COMP|66444-1|LNC|Blatella germanica recombinant (rBla g) 4 Ab.IgE|Blatella germanica recombinant (rBla g) 4 Ab.IgE
C3259282|T201|COMP|66445-8|LNC|Cyprinus carpio recombinant (rCyp c) 1 Ab.IgE|Cyprinus carpio recombinant (rCyp c) 1 Ab.IgE
C3259284|T201|COMP|66446-6|LNC|Daucus carota recombinant (rDau c) 1 Ab.IgE|Daucus carota recombinant (rDau c) 1 Ab.IgE
C3259286|T201|COMP|66447-4|LNC|Euroglyphus maynei recombinant (rEur m) 2 Ab.IgE|Euroglyphus maynei recombinant (rEur m) 2 Ab.IgE
C3259288|T201|COMP|66448-2|LNC|Latex recombinant (rHev b) 6 Ab.IgE|Latex recombinant (rHev b) 6 Ab.IgE
C3259331|T201|COMP|66753-5|LNC|Clot formation^after addition of heparinase|Clot formation^after addition of heparinase
C3259335|T201|COMP|66756-8|LNC|Clotting time^after addition of heparinase|Clotting time^after addition of heparinase
C3259336|T201|COMP|66757-6|LNC|Clot lysis estimate|Clot lysis estimate
C3259342|T201|COMP|67151-1|LNC|Troponin T.cardiac|Troponin T.cardiac
C3259389|T201|COMP|66449-0|LNC|Mercurialis annua recombinant (rMer a) 1 Ab.IgE|Mercurialis annua recombinant (rMer a) 1 Ab.IgE
C3259391|T201|COMP|66450-8|LNC|Olea europaea native (nOle e) 2 Ab.IgE|Olea europaea native (nOle e) 2 Ab.IgE
C3259393|T201|COMP|66451-6|LNC|Penaeus indicus native (nPen i) 11 Ab.IgE|Penaeus indicus native (nPen i) 11 Ab.IgE
C3259395|T201|COMP|66452-4|LNC|Triticum aestivum native (nTri a) 18 Ab.IgE|Triticum aestivum native (nTri a) 18 Ab.IgE
C3259397|T201|COMP|66453-2|LNC|M little c D super little d Ab|M little c D super little d Ab
C3259418|T201|COMP|66489-6|LNC|CYP2C19 gene targeted mutation analysis|CYP2C19 gene targeted mutation analysis
C3259419|T201|COMP|66491-2|LNC|Urease^2nd specimen|Urease^2nd specimen
C3259420|T201|COMP|66492-0|LNC|Urease^3rd specimen|Urease^3rd specimen
C3259421|T201|COMP|66493-8|LNC|Epstein Barr virus nuclear 1 Ab.IgG|Epstein Barr virus nuclear 1 Ab.IgG
C3259422|T201|COMP|66494-6|LNC|Spermatozoa.acrosome defects/100 spermatozoa|Spermatozoa.acrosome defects/100 spermatozoa
C3259424|T201|COMP|66495-3|LNC|Spermatozoa.abnormal head shape/100 spermatozoa|Spermatozoa.abnormal head shape/100 spermatozoa
C3259426|T201|COMP|66496-1|LNC|Spermatozoa.abnormal head size/100 spermatozoa|Spermatozoa.abnormal head size/100 spermatozoa
C3259428|T201|COMP|66497-9|LNC|Spermatozoa.double forms/100 spermatozoa|Spermatozoa.double forms/100 spermatozoa
C3259430|T201|COMP|66498-7|LNC|Spermatozoa.multiple defects/100 spermatozoa|Spermatozoa.multiple defects/100 spermatozoa
C3259432|T201|COMP|66499-5|LNC|Cholesterol.in VLDL.beta|Cholesterol.in VLDL.beta
C3259435|T201|COMP|66502-6|LNC|HBA1 gene targeted mutation analysis|HBA1 gene targeted mutation analysis
C3259660|T201|COMP|66853-3|LNC|Myeloperoxidase|Myeloperoxidase
C3259727|T201|COMP|66714-7|LNC|Vespula vulgaris recombinant (rVes v) 1 Ab.IgE|Vespula vulgaris recombinant (rVes v) 1 Ab.IgE
C3259731|T201|COMP|66716-2|LNC|Chlorhexidine Ab.IgE.RAST class|Chlorhexidine Ab.IgE.RAST class
C3259733|T201|COMP|66717-0|LNC|Chlorhexidine Ab.IgE|Chlorhexidine Ab.IgE
C3259736|T201|COMP|66719-6|LNC|Adenovirus DNA|Adenovirus DNA
C3259737|T201|COMP|66720-4|LNC|Adenovirus DNA|Adenovirus DNA
C3259738|T201|COMP|66721-2|LNC|Adenovirus DNA|Adenovirus DNA
C3259739|T201|COMP|66722-0|LNC|Adenovirus DNA|Adenovirus DNA
C3259740|T201|COMP|66723-8|LNC|Adenovirus DNA|Adenovirus DNA
C3259741|T201|COMP|66724-6|LNC|Adenovirus DNA|Adenovirus DNA
C3259742|T201|COMP|66725-3|LNC|Adenovirus DNA|Adenovirus DNA
C3259743|T201|COMP|66726-1|LNC|Adenovirus DNA|Adenovirus DNA
C3259744|T201|COMP|66727-9|LNC|Adenovirus DNA|Adenovirus DNA
C3259745|T201|COMP|66728-7|LNC|Adenovirus DNA|Adenovirus DNA
C3259746|T201|COMP|66729-5|LNC|Adenovirus DNA|Adenovirus DNA
C3259747|T201|COMP|66730-3|LNC|Adenovirus DNA|Adenovirus DNA
C3259748|T201|COMP|66731-1|LNC|Adenovirus DNA|Adenovirus DNA
C3259749|T201|COMP|66732-9|LNC|Corticotropin|Corticotropin
C3259750|T201|COMP|66733-7|LNC|Cortisol^afternoon specimen|Cortisol^afternoon specimen
C3259752|T201|COMP|66736-0|LNC|Normalized silica clotting time|Normalized silica clotting time
C3259753|T201|COMP|66737-8|LNC|CYP2C19 gene.c.1A>G(*4)|CYP2C19 gene.c.1A>G(*4)
C3259755|T201|COMP|66738-6|LNC|CYP2C19 gene.c.358T>C(*8)|CYP2C19 gene.c.358T>C(*8)
C3259757|T201|COMP|66739-4|LNC|CYP2C19 gene.c.395G>A(*6)|CYP2C19 gene.c.395G>A(*6)
C3259759|T201|COMP|66740-2|LNC|CYP2C19 gene.c.636G>A(*3)|CYP2C19 gene.c.636G>A(*3)
C3259761|T201|COMP|66741-0|LNC|CYP2C19 gene.c.681G>A(*2)|CYP2C19 gene.c.681G>A(*2)
C3259763|T201|COMP|66742-8|LNC|CYP2C19 gene.c.806C>T(*17)|CYP2C19 gene.c.806C>T(*17)
C3259765|T201|COMP|66743-6|LNC|CYP2C19 gene.c.IVS5+2T>A(*7)|CYP2C19 gene.c.IVS5+2T>A(*7)
C3259767|T201|COMP|66744-4|LNC|Heparin/body weight|Heparin/body weight
C3259769|T201|COMP|66745-1|LNC|Coagulum lysis^30M post maximum clot amplitude|Coagulum lysis^30M post maximum clot amplitude
C3259770|T201|COMP|66747-7|LNC|Clotting time|Clotting time
C3259771|T201|COMP|66748-5|LNC|Clot angle|Clot angle
C3259773|T201|COMP|66749-3|LNC|Circulatory assist status|Circulatory assist status
C3259775|T201|COMP|66750-1|LNC|Clot angle^after addition of heparinase|Clot angle^after addition of heparinase
C3259776|T201|COMP|66751-9|LNC|Clot strength|Clot strength
C3259778|T201|COMP|66752-7|LNC|Clot strength^after addition of heparinase|Clot strength^after addition of heparinase
C3259779|T201|COMP|66759-2|LNC|Heparin neutralization|Heparin neutralization
C3259780|T201|COMP|66760-0|LNC|Coagulation index|Coagulation index
C3259782|T201|COMP|66761-8|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C3259783|T201|COMP|66764-2|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C3259784|T201|COMP|66765-9|LNC|Albumin.pericard fld/Albumin.SerPl|Albumin.pericard fld/Albumin.SerPl
C3259786|T201|COMP|66766-7|LNC|Albumin.periton fld/Albumin.SerPl|Albumin.periton fld/Albumin.SerPl
C3259788|T201|COMP|66767-5|LNC|Vanillylmandelate/body weight|Vanillylmandelate/body weight
C3259790|T201|COMP|66768-3|LNC|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C3259791|T201|COMP|66769-1|LNC|Triglyceride|Triglyceride
C3259950|T201|COMP|66874-9|LNC|FMR1 gene activation|FMR1 gene activation
C3259952|T201|COMP|66875-6|LNC|FMR1 gene methylation/methylated+unmethylated|FMR1 gene methylation/methylated+unmethylated
C3259954|T201|COMP|66876-4|LNC|FMR1 gene premutation/premutation+full mutation|FMR1 gene premutation/premutation+full mutation
C3259956|T201|COMP|66877-2|LNC|Skin Ab pattern|Skin Ab pattern
C3259957|T201|COMP|66878-0|LNC|Skin Ab|Skin Ab
C3259958|T201|COMP|66879-8|LNC|Skin Ab.IgG|Skin Ab.IgG
C3259959|T201|COMP|66880-6|LNC|Skin Ab.IgG pattern|Skin Ab.IgG pattern
C3259960|T201|COMP|66881-4|LNC|Skin Ab.IgG|Skin Ab.IgG
C3259961|T201|COMP|66882-2|LNC|Skin Ab.IgG|Skin Ab.IgG
C3259962|T201|COMP|66883-0|LNC|Skin Ab.IgG|Skin Ab.IgG
C3260037|T201|COMP|66950-7|LNC|MALT1 18q21 gene rearrangements|MALT1 18q21 gene rearrangements
C3260251|T201|COMP|67126-3|LNC|Cannabinoids.synthetic|Cannabinoids.synthetic
C3260253|T201|COMP|67127-1|LNC|Cellularity assessment|Cellularity assessment
C3260255|T201|COMP|67128-9|LNC|Leukocytes.abnormal/100 leukocytes|Leukocytes.abnormal/100 leukocytes
C3260547|T201|COMP|67561-1|LNC|Corynebacterium diphtheriae DNA|Corynebacterium diphtheriae DNA
C3260549|T201|COMP|67562-9|LNC|Achromobacter sp DNA|Achromobacter sp DNA
C3260551|T201|COMP|67563-7|LNC|Legionella micdadei DNA|Legionella micdadei DNA
C3260554|T201|COMP|67568-6|LNC|Circulating tumor cells.breast|Circulating tumor cells.breast
C3260556|T201|COMP|67569-4|LNC|Streptococcus pyogenes M protein (emm) gene|Streptococcus pyogenes M protein (emm) gene
C3260622|T201|COMP|68380-5|LNC|Chromatin Ab|Chromatin Ab
C3260626|T201|COMP|68384-7|LNC|Specific gravity|Specific gravity
C3260627|T201|COMP|68385-4|LNC|Glomerular basement membrane Ab|Glomerular basement membrane Ab
C3260628|T201|COMP|68386-2|LNC|Glomerular basement membrane Ab.IgG|Glomerular basement membrane Ab.IgG
C3261131|T201|COMP|67866-4|LNC|Babesia identification panel|Babesia identification panel
C3261133|T201|COMP|68389-6|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3261134|T201|COMP|68391-2|LNC|Specimen volume|Specimen volume
C3261135|T201|COMP|68392-0|LNC|Basophils|Basophils
C3261136|T201|COMP|68393-8|LNC|Basophils|Basophils
C3261137|T201|COMP|68394-6|LNC|Basophils|Basophils
C3261138|T201|COMP|68395-3|LNC|Basophils|Basophils
C3261139|T201|COMP|68396-1|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C3261140|T201|COMP|68397-9|LNC|Basophils|Basophils
C3261141|T201|COMP|68398-7|LNC|Eosinophils|Eosinophils
C3261142|T201|COMP|68399-5|LNC|Eosinophils|Eosinophils
C3261143|T201|COMP|68400-1|LNC|Eosinophils|Eosinophils
C3261165|T201|COMP|68541-2|LNC|HYDROmorphone|HYDROmorphone
C3261166|T201|COMP|68542-0|LNC|Codeine|Codeine
C3261167|T201|COMP|68543-8|LNC|oxyCODONE|oxyCODONE
C3261168|T201|COMP|68544-6|LNC|HYDROcodone|HYDROcodone
C3261169|T201|COMP|68545-3|LNC|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C3261170|T201|COMP|68548-7|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C3261171|T201|COMP|68549-5|LNC|U2 small nuclear ribonucleoprotein Ab|U2 small nuclear ribonucleoprotein Ab
C3261229|T201|COMP|67725-2|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C3261230|T201|COMP|67726-0|LNC|Rickettsia sp DNA|Rickettsia sp DNA
C3261273|T201|COMP|67767-4|LNC|HEDIS 2012 panel|HEDIS 2012 panel
C3261301|T201|COMP|67790-6|LNC|Thromboelastography panel|Thromboelastography panel
C3261328|T201|COMP|67805-2|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C3261329|T201|COMP|67806-0|LNC|Measles virus Ag|Measles virus Ag
C3261330|T201|COMP|67807-8|LNC|Mumps virus Ag|Mumps virus Ag
C3261331|T201|COMP|67808-6|LNC|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C3261332|T201|COMP|67809-4|LNC|Parainfluenza virus 2 Ag|Parainfluenza virus 2 Ag
C3261333|T201|COMP|67810-2|LNC|Parainfluenza virus 3 Ag|Parainfluenza virus 3 Ag
C3261334|T201|COMP|67811-0|LNC|Parainfluenza virus 4 Ag|Parainfluenza virus 4 Ag
C3261335|T201|COMP|67812-8|LNC|Varicella zoster virus Ag|Varicella zoster virus Ag
C3261336|T201|COMP|67813-6|LNC|Fatty casts|Fatty casts
C3261337|T201|COMP|67814-4|LNC|Granulocytic cells/100 cells|Granulocytic cells/100 cells
C3261339|T201|COMP|67815-1|LNC|HTLV I Ab|HTLV I Ab
C3261340|T201|COMP|67816-9|LNC|Trisomy 18+Trisomy 13 risk|Trisomy 18+Trisomy 13 risk
C3261341|T201|COMP|67818-5|LNC|Parainfluenza virus 4a RNA|Parainfluenza virus 4a RNA
C3261342|T201|COMP|67819-3|LNC|Parainfluenza virus 4b RNA|Parainfluenza virus 4b RNA
C3261343|T201|COMP|67820-1|LNC|Human metapneumovirus A RNA|Human metapneumovirus A RNA
C3261345|T201|COMP|67821-9|LNC|Human metapneumovirus B RNA|Human metapneumovirus B RNA
C3261347|T201|COMP|67822-7|LNC|Fentanyl & Norfentanyl panel|Fentanyl & Norfentanyl panel
C3261349|T201|COMP|67826-8|LNC|Neutrophils|Neutrophils
C3261350|T201|COMP|67827-6|LNC|Lymphocytes|Lymphocytes
C3261351|T201|COMP|67828-4|LNC|Macrophages|Macrophages
C3261352|T201|COMP|67829-2|LNC|Eosinophils|Eosinophils
C3261353|T201|COMP|67830-0|LNC|Leukocytes other|Leukocytes other
C3261354|T201|COMP|67831-8|LNC|Erythrocytes|Erythrocytes
C3261355|T201|COMP|67832-6|LNC|Neutrophils|Neutrophils
C3261356|T201|COMP|67833-4|LNC|Lymphocytes|Lymphocytes
C3261357|T201|COMP|67834-2|LNC|Macrophages|Macrophages
C3261358|T201|COMP|67835-9|LNC|Eosinophils|Eosinophils
C3261359|T201|COMP|67836-7|LNC|Leukocytes other|Leukocytes other
C3261360|T201|COMP|67837-5|LNC|Cells counted.total|Cells counted.total
C3261361|T201|COMP|67838-3|LNC|Mephedrone|Mephedrone
C3261378|T201|COMP|67848-2|LNC|Leukocyte clumps|Leukocyte clumps
C3261385|T201|COMP|67867-2|LNC|Babesia sp identified|Babesia sp identified
C3261446|T201|COMP|68434-0|LNC|Leukocytes|Leukocytes
C3261447|T201|COMP|68435-7|LNC|Erythrocytes|Erythrocytes
C3261448|T201|COMP|68436-5|LNC|Appearance|Appearance
C3261449|T201|COMP|68437-3|LNC|Smudge cells|Smudge cells
C3261450|T201|COMP|68438-1|LNC|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3
C3261451|T201|COMP|68439-9|LNC|Gabapentin|Gabapentin
C3261452|T201|COMP|68440-7|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C3261453|T201|COMP|69031-3|LNC|Enterocyte Ab.IgA|Enterocyte Ab.IgA
C3261461|T201|COMP|68961-2|LNC|HIV 1 Ab|HIV 1 Ab
C3261462|T201|COMP|68962-0|LNC|Phenylbutazone|Phenylbutazone
C3261463|T201|COMP|68963-8|LNC|Collection date & time|Collection date & time
C3261464|T201|COMP|68964-6|LNC|Lan Ag|Lan Ag
C3261465|T201|COMP|68965-3|LNC|R little g Ag|R little g Ag
C3261466|T201|COMP|68966-1|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C3261467|T201|COMP|68967-9|LNC|Dantu Ab|Dantu Ab
C3261870|T201|COMP|68123-9|LNC|Circulating tumor cells.prostate|Circulating tumor cells.prostate
C3261872|T201|COMP|68124-7|LNC|Circulating tumor cells.colon|Circulating tumor cells.colon
C3262196|T201|COMP|68314-4|LNC|Meperidine & Normeperidine panel|Meperidine & Normeperidine panel
C3262197|T201|COMP|68315-1|LNC|Transcortin & Cortisol.free panel|Transcortin & Cortisol.free panel
C3262198|T201|COMP|68317-7|LNC|Metanephrine, Normetanephrine & Creatinine panel|Metanephrine, Normetanephrine & Creatinine panel
C3262199|T201|COMP|68318-5|LNC|Hypoglycemics panel|Hypoglycemics panel
C3262201|T201|COMP|68320-1|LNC|Polio virus Ab panel|Polio virus Ab panel
C3262207|T201|COMP|68324-3|LNC|von Willebrand factor.activity actual/Normal|von Willebrand factor.activity actual/Normal
C3262209|T201|COMP|68327-6|LNC|Age|Age
C3262210|T201|COMP|68328-4|LNC|Previous fetus defect|Previous fetus defect
C3262263|T201|COMP|68363-1|LNC|Oxygen saturation|Oxygen saturation
C3262264|T201|COMP|68364-9|LNC|Pincer cells|Pincer cells
C3262265|T201|COMP|68366-4|LNC|Bacteria identified|Bacteria identified
C3262266|T201|COMP|68367-2|LNC|Bilirubin|Bilirubin
C3262267|T201|COMP|68368-0|LNC|Leukocytes|Leukocytes
C3262268|T201|COMP|68369-8|LNC|Nuclear Ab|Nuclear Ab
C3262269|T201|COMP|68370-6|LNC|Nuclear Ab|Nuclear Ab
C3262270|T201|COMP|68371-4|LNC|Nuclear Ab|Nuclear Ab
C3262271|T201|COMP|68372-2|LNC|Nuclear Ab|Nuclear Ab
C3262272|T201|COMP|68373-0|LNC|Nuclear Ab|Nuclear Ab
C3262273|T201|COMP|68374-8|LNC|Nuclear Ab|Nuclear Ab
C3262274|T201|COMP|68375-5|LNC|Nuclear Ab|Nuclear Ab
C3262275|T201|COMP|68376-3|LNC|Nuclear Ab|Nuclear Ab
C3262276|T201|COMP|68378-9|LNC|Leukocytes.disintegrated/100 leukocytes|Leukocytes.disintegrated/100 leukocytes
C3262277|T201|COMP|68379-7|LNC|Phenylbutazone|Phenylbutazone
C3262278|T201|COMP|68387-0|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C3262279|T201|COMP|68388-8|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3262280|T201|COMP|68401-9|LNC|Eosinophils|Eosinophils
C3262281|T201|COMP|68402-7|LNC|Eosinophils|Eosinophils
C3262282|T201|COMP|68403-5|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C3262283|T201|COMP|68404-3|LNC|Lymphocytes|Lymphocytes
C3262284|T201|COMP|68405-0|LNC|Lymphocytes|Lymphocytes
C3262285|T201|COMP|68406-8|LNC|Lymphocytes.abnormal/100 leukocytes|Lymphocytes.abnormal/100 leukocytes
C3262286|T201|COMP|68407-6|LNC|Lymphocytes|Lymphocytes
C3262287|T201|COMP|68408-4|LNC|Macrophages|Macrophages
C3262288|T201|COMP|68409-2|LNC|Macrophages|Macrophages
C3262289|T201|COMP|68410-0|LNC|Macrophages|Macrophages
C3262290|T201|COMP|68411-8|LNC|Macrophages|Macrophages
C3262291|T201|COMP|68412-6|LNC|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C3262292|T201|COMP|68413-4|LNC|Macrophages|Macrophages
C3262293|T201|COMP|68414-2|LNC|Mesothelial cells|Mesothelial cells
C3262294|T201|COMP|68415-9|LNC|Mesothelial cells|Mesothelial cells
C3262295|T201|COMP|68416-7|LNC|Mesothelial cells|Mesothelial cells
C3262296|T201|COMP|68417-5|LNC|Mesothelial cells|Mesothelial cells
C3262297|T201|COMP|68418-3|LNC|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C3262298|T201|COMP|68419-1|LNC|Mesothelial cells|Mesothelial cells
C3262299|T201|COMP|68420-9|LNC|Monocytes|Monocytes
C3262300|T201|COMP|68421-7|LNC|Monocytes|Monocytes
C3262301|T201|COMP|68422-5|LNC|Monocytes|Monocytes
C3262302|T201|COMP|68423-3|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C3262303|T201|COMP|68424-1|LNC|Monocytes|Monocytes
C3262304|T201|COMP|68425-8|LNC|Neutrophils|Neutrophils
C3262305|T201|COMP|68426-6|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C3262306|T201|COMP|68427-4|LNC|Neutrophils|Neutrophils
C3262307|T201|COMP|68428-2|LNC|Leukocytes other|Leukocytes other
C3262308|T201|COMP|68429-0|LNC|Leukocytes other|Leukocytes other
C3262309|T201|COMP|68430-8|LNC|Leukocytes other|Leukocytes other
C3262310|T201|COMP|68431-6|LNC|Leukocytes other|Leukocytes other
C3262311|T201|COMP|68432-4|LNC|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C3262312|T201|COMP|68433-2|LNC|Leukocytes other|Leukocytes other
C3262313|T201|COMP|68441-5|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C3262332|T201|COMP|68452-2|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C3262333|T201|COMP|68453-0|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C3262334|T201|COMP|68454-8|LNC|Phenylbutazone|Phenylbutazone
C3262335|T201|COMP|68455-5|LNC|Appearance|Appearance
C3262338|T201|COMP|68457-1|LNC|Enterovirus & Parechovirus A RNA|Enterovirus & Parechovirus A RNA
C3262340|T201|COMP|68458-9|LNC|Trichomonas sp identified|Trichomonas sp identified
C3262342|T201|COMP|68460-5|LNC|Picornavirus Ag|Picornavirus Ag
C3262344|T201|COMP|68463-9|LNC|Rilpivirine|Rilpivirine
C3262345|T201|COMP|68464-7|LNC|Insulin^1.25H post XXX challenge|Insulin^1.25H post XXX challenge
C3262346|T201|COMP|68465-4|LNC|Insulin^1.75H post XXX challenge|Insulin^1.75H post XXX challenge
C3262347|T201|COMP|68466-2|LNC|Epstein-Barr virus-encoded RNA 1|Epstein-Barr virus-encoded RNA 1
C3262348|T201|COMP|68467-0|LNC|APOB+LDLR+PCSK9 gene targeted mutation analysis|APOB+LDLR+PCSK9 gene targeted mutation analysis
C3262388|T201|COMP|68502-4|LNC|Treponema pallidum Ab.IgG & IgM panel|Treponema pallidum Ab.IgG & IgM panel
C3262456|T201|COMP|69032-1|LNC|Enterocyte Ab.IgM|Enterocyte Ab.IgM
C3262458|T201|COMP|69033-9|LNC|Buprenorphine & Norbuprenorphine panel|Buprenorphine & Norbuprenorphine panel
C3262474|T201|COMP|69021-4|LNC|Amphetamines panel|Amphetamines panel
C3262476|T201|COMP|69022-2|LNC|Methamphetamine|Methamphetamine
C3262477|T201|COMP|69023-0|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C3262478|T201|COMP|69024-8|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C3262479|T201|COMP|69025-5|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C3262480|T201|COMP|69026-3|LNC|Opiates panel|Opiates panel
C3262481|T201|COMP|69027-1|LNC|Morphine|Morphine
C3262482|T201|COMP|69028-9|LNC|oxyMORphone|oxyMORphone
C3262485|T201|COMP|69030-5|LNC|Enterocyte Ab.IgG|Enterocyte Ab.IgG
C3262755|T201|COMP|68901-8|LNC|Erythrocytes|Erythrocytes
C3262756|T201|COMP|68902-6|LNC|Erythrocytes|Erythrocytes
C3262757|T201|COMP|68903-4|LNC|Erythrocytes|Erythrocytes
C3262758|T201|COMP|68910-9|LNC|Teratozoospermia index|Teratozoospermia index
C3262759|T201|COMP|68911-7|LNC|Lactate^post exercise|Lactate^post exercise
C3262760|T201|COMP|68912-5|LNC|Erythrocytes|Erythrocytes
C3262761|T201|COMP|68913-3|LNC|Voltage-gated potassium channel Ab|Voltage-gated potassium channel Ab
C3262765|T201|COMP|68917-4|LNC|Parathyrin.intact^20M post excision|Parathyrin.intact^20M post excision
C3262766|T201|COMP|68919-0|LNC|Somatotropin^15M post exercise|Somatotropin^15M post exercise
C3262767|T201|COMP|68923-2|LNC|Cancer Ag 125|Cancer Ag 125
C3262768|T201|COMP|68924-0|LNC|Cancer Ag 72-4|Cancer Ag 72-4
C3262769|T201|COMP|68925-7|LNC|Cancer Ag 72-4|Cancer Ag 72-4
C3262770|T201|COMP|68926-5|LNC|Cancer Ag 72-4|Cancer Ag 72-4
C3262771|T201|COMP|68927-3|LNC|Cytokeratin 19|Cytokeratin 19
C3262772|T201|COMP|68928-1|LNC|Cytokeratin 19|Cytokeratin 19
C3262773|T201|COMP|68929-9|LNC|Cytokeratin 19|Cytokeratin 19
C3262774|T201|COMP|68930-7|LNC|Albumin/Globulin|Albumin/Globulin
C3262775|T201|COMP|68931-5|LNC|Catecholamines.free|Catecholamines.free
C3262776|T201|COMP|68932-3|LNC|IgA.secretory|IgA.secretory
C3262777|T201|COMP|68933-1|LNC|IgA.secretory|IgA.secretory
C3262778|T201|COMP|68934-9|LNC|Heat shock protein 60 Ab|Heat shock protein 60 Ab
C3262780|T201|COMP|68935-6|LNC|LDL.oxidized Ab|LDL.oxidized Ab
C3262781|T201|COMP|68936-4|LNC|Saccharomyces cerevisiae Ab|Saccharomyces cerevisiae Ab
C3262782|T201|COMP|68937-2|LNC|Acetylcholine receptor Ab|Acetylcholine receptor Ab
C3262783|T201|COMP|68938-0|LNC|Cytokeratin 19|Cytokeratin 19
C3262784|T201|COMP|68939-8|LNC|Enolase.neuron specific|Enolase.neuron specific
C3262785|T201|COMP|68940-6|LNC|Somatotropin^90M post exercise|Somatotropin^90M post exercise
C3262786|T201|COMP|68941-4|LNC|Somatotropin^110M post exercise|Somatotropin^110M post exercise
C3262787|T201|COMP|68942-2|LNC|Somatotropin^130M post exercise|Somatotropin^130M post exercise
C3262788|T201|COMP|68944-8|LNC|Listeria monocytogenes Ab.IgG|Listeria monocytogenes Ab.IgG
C3262789|T201|COMP|68945-5|LNC|Cells.CD3+CD5+|Cells.CD3+CD5+
C3262790|T201|COMP|68946-3|LNC|SERPINA10 gene mutations tested for|SERPINA10 gene mutations tested for
C3262792|T201|COMP|68947-1|LNC|ATP1A2 gene mutations tested for|ATP1A2 gene mutations tested for
C3262794|T201|COMP|68952-1|LNC|Enolase.neuron specific|Enolase.neuron specific
C3262795|T201|COMP|68954-7|LNC|Streptococcus pyogenes rRNA|Streptococcus pyogenes rRNA
C3262796|T201|COMP|68955-4|LNC|Ketones|Ketones
C3262797|T201|COMP|68956-2|LNC|DNA double strand Ab.IgG|DNA double strand Ab.IgG
C3262799|T201|COMP|68959-6|LNC|Specimen condition|Specimen condition
C3262800|T201|COMP|68960-4|LNC|Myoglobin|Myoglobin
C3262801|T201|COMP|68968-7|LNC|H little y super little a Ab|H little y super little a Ab
C3262803|T201|COMP|68970-3|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C3262804|T201|COMP|68971-1|LNC|Color|Color
C3262805|T201|COMP|68972-9|LNC|Lupinus albus seed Ab.IgE.RAST Class|Lupinus albus seed Ab.IgE.RAST Class
C3262807|T201|COMP|68973-7|LNC|IgA.intrathecally synthesized/IgA.total|IgA.intrathecally synthesized/IgA.total
C3262809|T201|COMP|68974-5|LNC|IgG.intrathecally synthesized/IgG.total|IgG.intrathecally synthesized/IgG.total
C3262811|T201|COMP|68975-2|LNC|IgM.intrathecally synthesized/IgM.total|IgM.intrathecally synthesized/IgM.total
C3262813|T201|COMP|68976-0|LNC|Pseudomonas aeruginosa alkaline protease Ab|Pseudomonas aeruginosa alkaline protease Ab
C3262814|T201|COMP|68977-8|LNC|Pseudomonas aeruginosa elastase Ab|Pseudomonas aeruginosa elastase Ab
C3262815|T201|COMP|68978-6|LNC|Pseudomonas aeruginosa exotoxin A Ab|Pseudomonas aeruginosa exotoxin A Ab
C3262816|T201|COMP|68986-9|LNC|Influenza virus A H5a RNA|Influenza virus A H5a RNA
C3262818|T201|COMP|68987-7|LNC|Influenza virus A H5b RNA|Influenza virus A H5b RNA
C3262820|T201|COMP|68989-3|LNC|Performing laboratory|Performing laboratory
C3262821|T201|COMP|68990-1|LNC|Performing laboratory medical director|Performing laboratory medical director
C3262824|T201|COMP|68992-7|LNC|Specimen-related information panel|Specimen-related information panel
C3262825|T201|COMP|68993-5|LNC|Human RNase P RNA|Human RNase P RNA
C3262827|T201|COMP|68994-3|LNC|Performing laboratory name|Performing laboratory name
C3262838|T201|COMP|69003-2|LNC|Mononuclear cells.atypical/100 leukocytes|Mononuclear cells.atypical/100 leukocytes
C3262839|T201|COMP|69004-0|LNC|Granulocytes.immature/100 leukocytes|Granulocytes.immature/100 leukocytes
C3262840|T201|COMP|69005-7|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C3262841|T201|COMP|69006-5|LNC|Granulocytes.immature/100 leukocytes|Granulocytes.immature/100 leukocytes
C3262842|T201|COMP|69007-3|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C3262843|T201|COMP|69008-1|LNC|Cocaine panel|Cocaine panel
C3262844|T201|COMP|69009-9|LNC|Cocaine|Cocaine
C3262845|T201|COMP|69010-7|LNC|Benzoylecgonine|Benzoylecgonine
C3262846|T201|COMP|69011-5|LNC|Cocaethylene|Cocaethylene
C3262847|T201|COMP|69012-3|LNC|3-Hydroxybenzoylecgonine|3-Hydroxybenzoylecgonine
C3262856|T201|COMP|69017-2|LNC|Granulocytes.immature/100 leukocytes|Granulocytes.immature/100 leukocytes
C3262858|T201|COMP|69040-4|LNC|Chronic urticaria index panel|Chronic urticaria index panel
C3262867|T201|COMP|69047-9|LNC|Geneticist review|Geneticist review
C3262869|T201|COMP|69048-7|LNC|Immunologist review|Immunologist review
C3262871|T201|COMP|69049-5|LNC|Coagulation specialist review|Coagulation specialist review
C3262873|T201|COMP|69050-3|LNC|Toxicologist review|Toxicologist review
C3262874|T201|COMP|69051-1|LNC|Urinalysis specialist review|Urinalysis specialist review
C3262875|T201|COMP|69052-9|LNC|Flow cytometry specialist review|Flow cytometry specialist review
C3262877|T201|COMP|69053-7|LNC|Endocrinologist review|Endocrinologist review
C3263111|T201|COMP|69322-6|LNC|Health insurance plan benefits comment|Health insurance plan benefits comment
C3263156|T201|COMP|69353-1|LNC|HIV 2 RNA|HIV 2 RNA
C3263158|T201|COMP|69354-9|LNC|HIV 2 RNA|HIV 2 RNA
C3263159|T201|COMP|69355-6|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C3263160|T201|COMP|69356-4|LNC|oxyCODONE|oxyCODONE
C3263161|T201|COMP|69357-2|LNC|Amylase^post CFst|Amylase^post CFst
C3263162|T201|COMP|69358-0|LNC|Cells.HPV E6+E7 mRNA/cells|Cells.HPV E6+E7 mRNA/cells
C3263164|T201|COMP|69359-8|LNC|Amylase^2nd specimen post XXX challenge|Amylase^2nd specimen post XXX challenge
C3263165|T201|COMP|69360-6|LNC|Amylase^1st specimen post XXX challenge|Amylase^1st specimen post XXX challenge
C3263166|T201|COMP|69361-4|LNC|PCA3 score|PCA3 score
C3263167|T201|COMP|69362-2|LNC|PCA3 score|PCA3 score
C3263168|T201|COMP|69363-0|LNC|SERPINA10 gene targeted mutation analysis|SERPINA10 gene targeted mutation analysis
C3263170|T201|COMP|69364-8|LNC|ATP1A2 gene targeted mutation analysis|ATP1A2 gene targeted mutation analysis
C3263174|T201|COMP|69366-3|LNC|Bordetella pertussis Ab.IgA|Bordetella pertussis Ab.IgA
C3263175|T201|COMP|69367-1|LNC|Bordetella pertussis Ab.IgG|Bordetella pertussis Ab.IgG
C3263176|T201|COMP|69368-9|LNC|Bordetella pertussis Ab.IgM|Bordetella pertussis Ab.IgM
C3263177|T201|COMP|69369-7|LNC|Blood group antibody screen|Blood group antibody screen
C3263178|T201|COMP|69370-5|LNC|A1 Ab|A1 Ab
C3263179|T201|COMP|69371-3|LNC|B Ab|B Ab
C3263181|T201|COMP|69373-9|LNC|Passive D Ab|Passive D Ab
C3263200|T201|COMP|69383-8|LNC|AGXT gene targeted mutation analysis|AGXT gene targeted mutation analysis
C3263223|T201|COMP|69405-9|LNC|Glomerular filtration rate/1.73 sq M.predicted|Glomerular filtration rate/1.73 sq M.predicted
C3263245|T201|COMP|69429-9|LNC|Metabolic rate^resting|Metabolic rate^resting
C3263348|T201|COMP|69545-2|LNC|DNA region of interest start|DNA region of interest start
C3263350|T201|COMP|69546-0|LNC|DNA region of interest stop|DNA region of interest stop
C3263352|T201|COMP|69547-8|LNC|Reference nucleotide|Reference nucleotide
C3263353|T201|COMP|69548-6|LNC|Genetic variant assessment|Genetic variant assessment
C3263355|T201|COMP|69549-4|LNC|Genetic knowledge reference|Genetic knowledge reference
C3263357|T201|COMP|69550-2|LNC|Genetic knowledge reference|Genetic knowledge reference
C3263358|T201|COMP|69551-0|LNC|Variable nucleotide|Variable nucleotide
C3263693|T201|COMP|69039-6|LNC|Enterocyte Ab panel|Enterocyte Ab panel
C3263694|T201|COMP|66746-9|LNC|Specimen type|Specimen type
C3263708|T201|COMP|66735-2|LNC|Cortisol^AM peak specimen|Cortisol^AM peak specimen
C3481469|T201|COMP|48577-1|LNC|HFE gene.c.845G>A|HFE gene.c.845G>A
C3481470|T201|COMP|48579-7|LNC|HFE gene.c.187C>G|HFE gene.c.187C>G
C3481473|T201|COMP|66762-6|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C3481474|T201|COMP|66763-4|LNC|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C3481499|T201|COMP|68546-1|LNC|Mycoplasma hominis DNA|Mycoplasma hominis DNA
C3481500|T201|COMP|68547-9|LNC|Ureaplasma sp DNA|Ureaplasma sp DNA
C3481501|T201|COMP|68969-5|LNC|Activated clotting time|Activated clotting time
C3481505|T201|COMP|68325-0|LNC|Coagulation thrombin induced actual/Normal|Coagulation thrombin induced actual/Normal
C3481507|T201|COMP|68326-8|LNC|Coagulation reptilase induced actual/Normal|Coagulation reptilase induced actual/Normal
C3481524|T201|COMP|68377-1|LNC|Ribonucleoprotein extractable nuclear 63kD Ab|Ribonucleoprotein extractable nuclear 63kD Ab
C3481525|T201|COMP|69773-0|LNC|Dicarboxyoleylcarnitine (C18:1-DC)|Dicarboxyoleylcarnitine (C18:1-DC)
C3481526|T201|COMP|69774-8|LNC|Propionylcarnitine (C3)|Propionylcarnitine (C3)
C3481527|T201|COMP|69775-5|LNC|Stearoylcarnitine (C18)|Stearoylcarnitine (C18)
C3481528|T201|COMP|69776-3|LNC|Suberylcarnitine (C8-DC)/Creatinine|Suberylcarnitine (C8-DC)/Creatinine
C3481530|T201|COMP|69777-1|LNC|Suberylcarnitine (C8-DC)|Suberylcarnitine (C8-DC)
C3481531|T201|COMP|69778-9|LNC|Suberylcarnitine (C8-DC)|Suberylcarnitine (C8-DC)
C3481532|T201|COMP|69779-7|LNC|Suberylcarnitine (C8-DC)|Suberylcarnitine (C8-DC)
C3481533|T201|COMP|69780-5|LNC|2-Hydroxyisovalerate|2-Hydroxyisovalerate
C3481534|T201|COMP|69781-3|LNC|2-Hydroxyisovalerate|2-Hydroxyisovalerate
C3481535|T201|COMP|69782-1|LNC|2-Hydroxyphenylacetate|2-Hydroxyphenylacetate
C3481536|T201|COMP|69783-9|LNC|2-Hydroxyphenylacetate|2-Hydroxyphenylacetate
C3481537|T201|COMP|69784-7|LNC|2-Hydroxysebacate|2-Hydroxysebacate
C3481538|T201|COMP|69785-4|LNC|2-Hydroxysebacate|2-Hydroxysebacate
C3481539|T201|COMP|69786-2|LNC|2-Methylacetoacetate|2-Methylacetoacetate
C3481540|T201|COMP|69787-0|LNC|2-Methylacetoacetate|2-Methylacetoacetate
C3481541|T201|COMP|69788-8|LNC|2-Methyl-3-Hydroxybutyrate|2-Methyl-3-Hydroxybutyrate
C3481542|T201|COMP|69789-6|LNC|2-Methyl-3-Hydroxybutyrate|2-Methyl-3-Hydroxybutyrate
C3481543|T201|COMP|69790-4|LNC|2-Methylbutyrylglycine|2-Methylbutyrylglycine
C3481544|T201|COMP|69791-2|LNC|Tetradecadienoylcarnitine (C14:2)/Creatinine|Tetradecadienoylcarnitine (C14:2)/Creatinine
C3481546|T201|COMP|69792-0|LNC|Tetradecadienoylcarnitine (C14:2)|Tetradecadienoylcarnitine (C14:2)
C3481547|T201|COMP|70132-6|LNC|Rickettsia typhus group Ab.IgG^2nd specimen|Rickettsia typhus group Ab.IgG^2nd specimen
C3481548|T201|COMP|70133-4|LNC|Rickettsia typhus group Ab.IgM^1st specimen|Rickettsia typhus group Ab.IgM^1st specimen
C3481549|T201|COMP|70134-2|LNC|Rickettsia typhus group Ab.IgM^2nd specimen|Rickettsia typhus group Ab.IgM^2nd specimen
C3481552|T201|COMP|70138-3|LNC|Amphetamines|Amphetamines
C3481553|T201|COMP|70139-1|LNC|Barbiturates|Barbiturates
C3481554|T201|COMP|70140-9|LNC|Benzodiazepines|Benzodiazepines
C3481555|T201|COMP|70141-7|LNC|Benzodiazepines|Benzodiazepines
C3481556|T201|COMP|68948-9|LNC|Candida albicans Ab|Candida albicans Ab
C3481557|T201|COMP|68949-7|LNC|Ehrlichia chaffeensis Ab|Ehrlichia chaffeensis Ab
C3481558|T201|COMP|68950-5|LNC|Herpes virus 8 Ab.IgG|Herpes virus 8 Ab.IgG
C3481559|T201|COMP|68951-3|LNC|Pyruvate^20M post XXX challenge|Pyruvate^20M post XXX challenge
C3481561|T201|COMP|70008-8|LNC|Enterovirus Ab.IgM|Enterovirus Ab.IgM
C3481562|T201|COMP|70009-6|LNC|Enterovirus Ab.IgM|Enterovirus Ab.IgM
C3481563|T201|COMP|70010-4|LNC|Enterovirus Ab.IgG|Enterovirus Ab.IgG
C3481565|T201|COMP|70011-2|LNC|Enterovirus Ab.IgG|Enterovirus Ab.IgG
C3481566|T201|COMP|70012-0|LNC|Coxsackievirus Ab.IgM|Coxsackievirus Ab.IgM
C3481568|T201|COMP|70013-8|LNC|Coxsackievirus Ab.IgG|Coxsackievirus Ab.IgG
C3481606|T201|COMP|68943-0|LNC|Voltage-gated potassium channel Ab|Voltage-gated potassium channel Ab
C3481607|T201|COMP|68979-4|LNC|Rivaroxaban|Rivaroxaban
C3481608|T201|COMP|68980-2|LNC|Dabigatran|Dabigatran
C3481609|T201|COMP|68981-0|LNC|Argatroban|Argatroban
C3481610|T201|COMP|68982-8|LNC|PFGE panel|PFGE panel
C3481611|T201|COMP|68983-6|LNC|National (USA) PFGE pattern|National (USA) PFGE pattern
C3481612|T201|COMP|68985-1|LNC|Bacteria antigenic formula|Bacteria antigenic formula
C3481613|T201|COMP|68988-5|LNC|Local PFGE pattern|Local PFGE pattern
C3481614|T201|COMP|69018-0|LNC|Lymphocyte proliferation mitogen panel|Lymphocyte proliferation mitogen panel
C3481619|T201|COMP|69042-0|LNC|Lymphocyte proliferation antigen panel|Lymphocyte proliferation antigen panel
C3481647|T201|COMP|70197-9|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C3481648|T201|COMP|70198-7|LNC|Acetaminophen|Acetaminophen
C3481649|T201|COMP|70199-5|LNC|Bilirubin|Bilirubin
C3481650|T201|COMP|70200-1|LNC|Cholesterol.in HDL/Cholesterol.total|Cholesterol.in HDL/Cholesterol.total
C3481651|T201|COMP|70201-9|LNC|Cholesterol.in IDL|Cholesterol.in IDL
C3481652|T201|COMP|70202-7|LNC|Cholesterol.in IDL+Cholesterol.in VLDL 3|Cholesterol.in IDL+Cholesterol.in VLDL 3
C3481653|T201|COMP|70203-5|LNC|Cholesterol.in VLDL 3|Cholesterol.in VLDL 3
C3481662|T201|COMP|69478-6|LNC|AGXT gene deletion+duplication|AGXT gene deletion+duplication
C3481666|T201|COMP|69480-2|LNC|CFTR gene deletion+duplication|CFTR gene deletion+duplication
C3481668|T201|COMP|69481-0|LNC|ACVRL1 gene+ENG gene deletion+duplication|ACVRL1 gene+ENG gene deletion+duplication
C3481674|T201|COMP|69571-8|LNC|Bacterial vaginosis DNA & score panel|Bacterial vaginosis DNA & score panel
C3481675|T201|COMP|69572-6|LNC|ERCC1 Ag|ERCC1 Ag
C3481676|T201|COMP|69573-4|LNC|Tiglylcarnitine+methylcrotonylcarnitine (C5:1)|Tiglylcarnitine+methylcrotonylcarnitine (C5:1)
C3481677|T201|COMP|69574-2|LNC|Furazolidone|Furazolidone
C3481678|T201|COMP|69575-9|LNC|Campylobacter jejuni Ab|Campylobacter jejuni Ab
C3481679|T201|COMP|69576-7|LNC|Campylobacter fetus Ab|Campylobacter fetus Ab
C3481680|T201|COMP|69577-5|LNC|Hepatitis E virus RNA|Hepatitis E virus RNA
C3481683|T201|COMP|69579-1|LNC|Local PFGE event description|Local PFGE event description
C3481684|T201|COMP|69580-9|LNC|Local assigning authority|Local assigning authority
C3481685|T201|COMP|69581-7|LNC|National (USA) PFGE cluster code or CDC cluster|National (USA) PFGE cluster code or CDC cluster
C3481686|T201|COMP|69582-5|LNC|PFGE restriction enzyme|PFGE restriction enzyme
C3481687|T201|COMP|69895-1|LNC|Service comment 68|Service comment 68
C3481688|T201|COMP|69896-9|LNC|Service comment 69|Service comment 69
C3481689|T201|COMP|69897-7|LNC|Service comment 70|Service comment 70
C3481690|T201|COMP|69898-5|LNC|Service comment 71|Service comment 71
C3481691|T201|COMP|69899-3|LNC|Service comment 72|Service comment 72
C3481692|T201|COMP|69900-9|LNC|Service comment 73|Service comment 73
C3481693|T201|COMP|69901-7|LNC|Service comment 74|Service comment 74
C3481694|T201|COMP|69902-5|LNC|Service comment 75|Service comment 75
C3481695|T201|COMP|69903-3|LNC|Service comment 76|Service comment 76
C3481703|T201|COMP|69410-9|LNC|Haemophilus influenzae|Haemophilus influenzae
C3481704|T201|COMP|69419-0|LNC|Cholesterol.in LDL|Cholesterol.in LDL
C3481705|T201|COMP|69420-8|LNC|Heterophile Ab|Heterophile Ab
C3481706|T201|COMP|69421-6|LNC|Corylus avellana recombinant (rCor a) 1 Ab.IgE|Corylus avellana recombinant (rCor a) 1 Ab.IgE
C3481708|T201|COMP|69422-4|LNC|Carnitine.free (C0)|Carnitine.free (C0)
C3481709|T201|COMP|69423-2|LNC|Rosner index|Rosner index
C3481710|T201|COMP|69424-0|LNC|Nitrogen|Nitrogen
C3481711|T201|COMP|69425-7|LNC|Calcium|Calcium
C3481712|T201|COMP|69426-5|LNC|Medical director review|Medical director review
C3481713|T201|COMP|69427-3|LNC|Supervisor review|Supervisor review
C3481723|T201|COMP|69486-9|LNC|LDLR gene deletion+duplication|LDLR gene deletion+duplication
C3481725|T201|COMP|69487-7|LNC|TNFRSF13B gene full mutation analysis|TNFRSF13B gene full mutation analysis
C3481731|T201|COMP|69922-3|LNC|(Beef+Chicken+Pork) Ab.IgE|(Beef+Chicken+Pork) Ab.IgE
C3481732|T201|COMP|69923-1|LNC|European tick borne encephalitis virus Ab.IgM|European tick borne encephalitis virus Ab.IgM
C3481733|T201|COMP|69924-9|LNC|European tick borne encephalitis virus Ab.IgM|European tick borne encephalitis virus Ab.IgM
C3481736|T201|COMP|69926-4|LNC|European tick borne encephalitis virus Ab.IgG|European tick borne encephalitis virus Ab.IgG
C3481737|T201|COMP|69927-2|LNC|European tick borne encephalitis virus Ab.IgG|European tick borne encephalitis virus Ab.IgG
C3481740|T201|COMP|69929-8|LNC|Respiratory syncytial virus Ab.IgA|Respiratory syncytial virus Ab.IgA
C3481799|T201|COMP|69553-6|LNC|Lactose tolerance|Lactose tolerance
C3481800|T201|COMP|69554-4|LNC|Lactose tolerance panel^dosage unspecified|Lactose tolerance panel^dosage unspecified
C3481801|T201|COMP|69555-1|LNC|Lactose tolerance panel^dosage unspecified|Lactose tolerance panel^dosage unspecified
C3481802|T201|COMP|69556-9|LNC|Ku Ab|Ku Ab
C3481803|T201|COMP|69557-7|LNC|OJ Ab|OJ Ab
C3481804|T201|COMP|69558-5|LNC|Ma1 Ab|Ma1 Ab
C3481805|T201|COMP|69559-3|LNC|Ma1 Ab|Ma1 Ab
C3481806|T201|COMP|69560-1|LNC|Enolase.neuron specific|Enolase.neuron specific
C3481807|T201|COMP|69561-9|LNC|Thyrotropin|Thyrotropin
C3481808|T201|COMP|69562-7|LNC|Candida albicans DNA|Candida albicans DNA
C3481809|T201|COMP|69563-5|LNC|Candida glabrata DNA|Candida glabrata DNA
C3481810|T201|COMP|69564-3|LNC|Bacterial vaginosis score|Bacterial vaginosis score
C3481811|T201|COMP|69565-0|LNC|Atopobium vaginae DNA|Atopobium vaginae DNA
C3481812|T201|COMP|69566-8|LNC|Bacterial vaginosis associated bacterium 2 DNA|Bacterial vaginosis associated bacterium 2 DNA
C3481813|T201|COMP|69567-6|LNC|Megasphaera sp type 1 DNA|Megasphaera sp type 1 DNA
C3481814|T201|COMP|69568-4|LNC|Bacterial vaginosis|Bacterial vaginosis
C3481818|T201|COMP|69668-2|LNC|HIV 1 & 2 Ab|HIV 1 & 2 Ab
C3481823|T201|COMP|69738-3|LNC|Differential panel, method unspecified|Differential panel, method unspecified
C3481824|T201|COMP|69739-1|LNC|Drugs of abuse panel|Drugs of abuse panel
C3481825|T201|COMP|69740-9|LNC|Cell count panel|Cell count panel
C3481826|T201|COMP|69741-7|LNC|Differential panel|Differential panel
C3481827|T201|COMP|69742-5|LNC|CBC W Differential panel, method unspecified|CBC W Differential panel, method unspecified
C3481837|T201|COMP|69765-6|LNC|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C3481838|T201|COMP|69766-4|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C3481839|T201|COMP|69767-2|LNC|La Crosse virus RNA|La Crosse virus RNA
C3481840|T201|COMP|69768-0|LNC|2-Oxoadipate|2-Oxoadipate
C3481841|T201|COMP|69769-8|LNC|Dicarboxyoleylcarnitine (C18:1-DC)/Creatinine|Dicarboxyoleylcarnitine (C18:1-DC)/Creatinine
C3481843|T201|COMP|69770-6|LNC|Dicarboxyoleylcarnitine (C18:1-DC)|Dicarboxyoleylcarnitine (C18:1-DC)
C3481844|T201|COMP|69771-4|LNC|Dicarboxyoleylcarnitine (C18:1-DC)|Dicarboxyoleylcarnitine (C18:1-DC)
C3481845|T201|COMP|69772-2|LNC|Orotate|Orotate
C3481846|T201|COMP|69793-8|LNC|Tetradecadienoylcarnitine (C14:2)|Tetradecadienoylcarnitine (C14:2)
C3481847|T201|COMP|69794-6|LNC|Tetradecadienoylcarnitine (C14:2)|Tetradecadienoylcarnitine (C14:2)
C3481850|T201|COMP|69796-1|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C3481851|T201|COMP|69797-9|LNC|1-Hydroxymidazolam|1-Hydroxymidazolam
C3481852|T201|COMP|69798-7|LNC|2,5-dimethoxy-4-bromoamphetamine|2,5-dimethoxy-4-bromoamphetamine
C3481853|T201|COMP|69799-5|LNC|21-Deoxycorticosterone|21-Deoxycorticosterone
C3481854|T201|COMP|69800-1|LNC|Methyl ethyl ketone|Methyl ethyl ketone
C3481855|T201|COMP|69801-9|LNC|2-Oxoadipate|2-Oxoadipate
C3481856|T201|COMP|69802-7|LNC|Alpha ketoglutarate|Alpha ketoglutarate
C3481857|T201|COMP|69803-5|LNC|Alpha ketoglutarate|Alpha ketoglutarate
C3481858|T201|COMP|69804-3|LNC|2-Oxoisocaproate|2-Oxoisocaproate
C3481860|T201|COMP|69806-8|LNC|2-Dechloroethylifosfamide^post dose ifosfamide|2-Dechloroethylifosfamide^post dose ifosfamide
C3481861|T201|COMP|69807-6|LNC|2-Dechloroethylifosfamide^pre dose ifosfamide|2-Dechloroethylifosfamide^pre dose ifosfamide
C3481862|T201|COMP|69808-4|LNC|2-Dechloroethylifosfamide^pre dose ifosfamide|2-Dechloroethylifosfamide^pre dose ifosfamide
C3481863|T201|COMP|69809-2|LNC|2-Dechloroethylifosfamide^1D post dose ifosfamide|2-Dechloroethylifosfamide^1D post dose ifosfamide
C3481864|T201|COMP|69810-0|LNC|2-Dechloroethylifosfamide^1D post dose ifosfamide|2-Dechloroethylifosfamide^1D post dose ifosfamide
C3481865|T201|COMP|69811-8|LNC|2-Dechloroethylifosfamide^2D post dose ifosfamide|2-Dechloroethylifosfamide^2D post dose ifosfamide
C3481866|T201|COMP|69812-6|LNC|2-Dechloroethylifosfamide^2D post dose ifosfamide|2-Dechloroethylifosfamide^2D post dose ifosfamide
C3481867|T201|COMP|69813-4|LNC|2-Dechloroethylifosfamide^3D post dose ifosfamide|2-Dechloroethylifosfamide^3D post dose ifosfamide
C3481868|T201|COMP|69814-2|LNC|2-Dechloroethylifosfamide^3D post dose ifosfamide|2-Dechloroethylifosfamide^3D post dose ifosfamide
C3481869|T201|COMP|69815-9|LNC|2-Dechloroethylifosfamide^4D post dose ifosfamide|2-Dechloroethylifosfamide^4D post dose ifosfamide
C3481870|T201|COMP|69816-7|LNC|2-Dechloroethylifosfamide^4D post dose ifosfamide|2-Dechloroethylifosfamide^4D post dose ifosfamide
C3481871|T201|COMP|69817-5|LNC|2-Dechloroethylifosfamide^5D post dose ifosfamide|2-Dechloroethylifosfamide^5D post dose ifosfamide
C3481872|T201|COMP|69818-3|LNC|2-Dechloroethylifosfamide^5D post dose ifosfamide|2-Dechloroethylifosfamide^5D post dose ifosfamide
C3481873|T201|COMP|69819-1|LNC|2-Dechloroethylifosfamide^6D post dose ifosfamide|2-Dechloroethylifosfamide^6D post dose ifosfamide
C3481874|T201|COMP|69820-9|LNC|2-Dechloroethylifosfamide^6D post dose ifosfamide|2-Dechloroethylifosfamide^6D post dose ifosfamide
C3481875|T201|COMP|69821-7|LNC|2-Dechloroethylifosfamide^6D post dose ifosfamide|2-Dechloroethylifosfamide^6D post dose ifosfamide
C3481876|T201|COMP|69822-5|LNC|2-Dechloroethylifosfamide^7D post dose ifosfamide|2-Dechloroethylifosfamide^7D post dose ifosfamide
C3481877|T201|COMP|69823-3|LNC|2-Dechloroethylifosfamide^7D post dose ifosfamide|2-Dechloroethylifosfamide^7D post dose ifosfamide
C3481878|T201|COMP|69824-1|LNC|2-Dechloroethylifosfamide^7D post dose ifosfamide|2-Dechloroethylifosfamide^7D post dose ifosfamide
C3481879|T201|COMP|69825-8|LNC|2-Ethylhydracrylate|2-Ethylhydracrylate
C3481880|T201|COMP|69826-6|LNC|2-Ethylhydracrylate|2-Ethylhydracrylate
C3481881|T201|COMP|69827-4|LNC|2-Methylglutarate|2-Methylglutarate
C3481882|T201|COMP|69828-2|LNC|Methylsuccinate|Methylsuccinate
C3481883|T201|COMP|69829-0|LNC|Methylsuccinate|Methylsuccinate
C3481884|T201|COMP|69830-8|LNC|3,4-Dihydroxyphenylacetate|3,4-Dihydroxyphenylacetate
C3481885|T201|COMP|69831-6|LNC|3,4-Dihydroxyphenylacetate/Creatinine|3,4-Dihydroxyphenylacetate/Creatinine
C3481886|T201|COMP|69832-4|LNC|3-Hydroxy,3-Methylglutarate|3-Hydroxy,3-Methylglutarate
C3481887|T201|COMP|69833-2|LNC|3-Hydroxy,3-Methylglutarate|3-Hydroxy,3-Methylglutarate
C3481888|T201|COMP|69834-0|LNC|3-Hydroxy,3-Methylglutarate|3-Hydroxy,3-Methylglutarate
C3481889|T201|COMP|69835-7|LNC|3-Hydroxyadipate|3-Hydroxyadipate
C3481890|T201|COMP|69836-5|LNC|3-Hydroxyadipate|3-Hydroxyadipate
C3481891|T201|COMP|69837-3|LNC|3-Hydroxyglutarate|3-Hydroxyglutarate
C3481892|T201|COMP|69838-1|LNC|2-Hydroxy-3-Methylvalerate|2-Hydroxy-3-Methylvalerate
C3481893|T201|COMP|69839-9|LNC|2-Hydroxy-3-Methylvalerate|2-Hydroxy-3-Methylvalerate
C3481894|T201|COMP|69840-7|LNC|2-Hydroxyadipate|2-Hydroxyadipate
C3481895|T201|COMP|69841-5|LNC|2-Hydroxyadipate|2-Hydroxyadipate
C3481896|T201|COMP|69842-3|LNC|Alpha hydroxybutyrate|Alpha hydroxybutyrate
C3481897|T201|COMP|69843-1|LNC|Alpha hydroxybutyrate|Alpha hydroxybutyrate
C3481898|T201|COMP|69844-9|LNC|2-Hydroxyglutarate|2-Hydroxyglutarate
C3481899|T201|COMP|69845-6|LNC|2-Hydroxyglutarate|2-Hydroxyglutarate
C3481900|T201|COMP|69846-4|LNC|2-Hydroxyisobutyrate|2-Hydroxyisobutyrate
C3481901|T201|COMP|69847-2|LNC|2-Hydroxyisobutyrate|2-Hydroxyisobutyrate
C3481902|T201|COMP|69848-0|LNC|2-Hydroxyisocaproate|2-Hydroxyisocaproate
C3481903|T201|COMP|69849-8|LNC|2-Hydroxyisocaproate|2-Hydroxyisocaproate
C3481904|T201|COMP|69850-6|LNC|3-Hydroxyglutarate|3-Hydroxyglutarate
C3481905|T201|COMP|69851-4|LNC|3-Hydroxyglutarate|3-Hydroxyglutarate
C3481906|T201|COMP|69852-2|LNC|3-Hydroxyisobutyrate|3-Hydroxyisobutyrate
C3481907|T201|COMP|69853-0|LNC|3-Hydroxyisobutyrate|3-Hydroxyisobutyrate
C3481930|T201|COMP|69868-8|LNC|Service comment 41|Service comment 41
C3481931|T201|COMP|69869-6|LNC|Service comment 42|Service comment 42
C3481932|T201|COMP|69870-4|LNC|Service comment 43|Service comment 43
C3481933|T201|COMP|69871-2|LNC|Service comment 44|Service comment 44
C3481934|T201|COMP|69872-0|LNC|Service comment 45|Service comment 45
C3481935|T201|COMP|69873-8|LNC|Service comment 46|Service comment 46
C3481936|T201|COMP|69874-6|LNC|Service comment 47|Service comment 47
C3481937|T201|COMP|69875-3|LNC|Service comment 48|Service comment 48
C3481938|T201|COMP|69876-1|LNC|Service comment 49|Service comment 49
C3481939|T201|COMP|69877-9|LNC|Service comment 50|Service comment 50
C3481940|T201|COMP|69878-7|LNC|Service comment 51|Service comment 51
C3481941|T201|COMP|69879-5|LNC|Service comment 52|Service comment 52
C3481942|T201|COMP|69880-3|LNC|Service comment 53|Service comment 53
C3481943|T201|COMP|69881-1|LNC|Service comment 54|Service comment 54
C3481944|T201|COMP|69882-9|LNC|Service comment 55|Service comment 55
C3481945|T201|COMP|69883-7|LNC|Service comment 56|Service comment 56
C3481946|T201|COMP|69884-5|LNC|Service comment 57|Service comment 57
C3481947|T201|COMP|69885-2|LNC|Service comment 58|Service comment 58
C3481948|T201|COMP|69886-0|LNC|Service comment 59|Service comment 59
C3481949|T201|COMP|69887-8|LNC|Service comment 60|Service comment 60
C3481950|T201|COMP|69888-6|LNC|Service comment 61|Service comment 61
C3481951|T201|COMP|69889-4|LNC|Service comment 62|Service comment 62
C3481952|T201|COMP|69890-2|LNC|Service comment 63|Service comment 63
C3481953|T201|COMP|69891-0|LNC|Service comment 64|Service comment 64
C3481954|T201|COMP|69892-8|LNC|Service comment 65|Service comment 65
C3481955|T201|COMP|69893-6|LNC|Service comment 66|Service comment 66
C3481956|T201|COMP|69894-4|LNC|Service comment 67|Service comment 67
C3481957|T201|COMP|69904-1|LNC|Service comment 77|Service comment 77
C3481958|T201|COMP|69905-8|LNC|Service comment 78|Service comment 78
C3481959|T201|COMP|69906-6|LNC|Service comment 79|Service comment 79
C3481960|T201|COMP|69907-4|LNC|Service comment 80|Service comment 80
C3481963|T201|COMP|69910-8|LNC|Basophils+Mast cells/100 leukocytes|Basophils+Mast cells/100 leukocytes
C3481965|T201|COMP|69913-2|LNC|Basophils+Mast cells/100 leukocytes|Basophils+Mast cells/100 leukocytes
C3481966|T201|COMP|69916-5|LNC|Basophils+Mast cells/100 leukocytes|Basophils+Mast cells/100 leukocytes
C3481967|T201|COMP|69918-1|LNC|Coagulation thrombin induced.high dose|Coagulation thrombin induced.high dose
C3481970|T201|COMP|69920-7|LNC|Adenovirus Ab.IgA|Adenovirus Ab.IgA
C3481972|T201|COMP|69921-5|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C3481973|T201|COMP|69930-6|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C3481975|T201|COMP|69933-0|LNC|Ureaplasma parvum DNA|Ureaplasma parvum DNA
C3481976|T201|COMP|69934-8|LNC|Ureaplasma urealyticum+Ureaplasma parvum DNA|Ureaplasma urealyticum+Ureaplasma parvum DNA
C3481977|T201|COMP|69935-5|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C3481978|T201|COMP|69936-3|LNC|Gardnerella vaginalis DNA|Gardnerella vaginalis DNA
C3481979|T201|COMP|69937-1|LNC|Trichomonas vaginalis DNA|Trichomonas vaginalis DNA
C3481980|T201|COMP|69938-9|LNC|Astrovirus RNA|Astrovirus RNA
C3481981|T201|COMP|69939-7|LNC|Trichophyton rubrum DNA|Trichophyton rubrum DNA
C3481982|T201|COMP|69941-3|LNC|Glucose^20M post dose lactose PO|Glucose^20M post dose lactose PO
C3481983|T201|COMP|69942-1|LNC|Glucose^40M post dose lactose PO|Glucose^40M post dose lactose PO
C3481984|T201|COMP|69943-9|LNC|Glucose^20M post 50 g lactose PO|Glucose^20M post 50 g lactose PO
C3481985|T201|COMP|69944-7|LNC|Glucose^40M post 50 g lactose PO|Glucose^40M post 50 g lactose PO
C3481986|T201|COMP|69945-4|LNC|Insulin-like growth factor binding protein 1|Insulin-like growth factor binding protein 1
C3481987|T201|COMP|69946-2|LNC|Treponema pallidum Ab.IgM|Treponema pallidum Ab.IgM
C3481988|T201|COMP|69947-0|LNC|Triglyceride|Triglyceride
C3481989|T201|COMP|69948-8|LNC|Bordetella parapertussis Ab.IgG|Bordetella parapertussis Ab.IgG
C3481990|T201|COMP|69949-6|LNC|Epstein Barr virus capsid Ab.IgG avidity|Epstein Barr virus capsid Ab.IgG avidity
C3481992|T201|COMP|69950-4|LNC|Hemoglobin|Hemoglobin
C3481993|T201|COMP|69951-2|LNC|Amylase.pancreatic/Creatinine|Amylase.pancreatic/Creatinine
C3481995|T201|COMP|69952-0|LNC|Liver kidney microsomal 1 Ab.IgG|Liver kidney microsomal 1 Ab.IgG
C3481996|T201|COMP|69953-8|LNC|Purkinje cell cytoplasmic type 1 Ab.IgG|Purkinje cell cytoplasmic type 1 Ab.IgG
C3481997|T201|COMP|69954-6|LNC|Neuronal nuclear type 2 Ab.IgG|Neuronal nuclear type 2 Ab.IgG
C3481998|T201|COMP|69955-3|LNC|Intestinal goblet cell Ab|Intestinal goblet cell Ab
C3481999|T201|COMP|69956-1|LNC|Human upstream binding factor Ab.IgG|Human upstream binding factor Ab.IgG
C3482000|T201|COMP|69957-9|LNC|Proteinase 3 Ab.IgG|Proteinase 3 Ab.IgG
C3482004|T201|COMP|69961-1|LNC|Hepatitis E virus RNA|Hepatitis E virus RNA
C3482005|T201|COMP|69962-9|LNC|Respiratory syncytial virus Ab.IgM|Respiratory syncytial virus Ab.IgM
C3482007|T201|COMP|69964-5|LNC|Bicarbonate^^standard|Bicarbonate^^standard
C3482008|T201|COMP|69965-2|LNC|Clinical cytogeneticist review|Clinical cytogeneticist review
C3482032|T201|COMP|70014-6|LNC|Parainfluenza virus 1+2+3+4 Ab.IgA|Parainfluenza virus 1+2+3+4 Ab.IgA
C3482033|T201|COMP|70015-3|LNC|Streptococcus sp DNA|Streptococcus sp DNA
C3482034|T201|COMP|70016-1|LNC|Staphylococcus sp.coagulase negative DNA|Staphylococcus sp.coagulase negative DNA
C3482035|T201|COMP|70017-9|LNC|Parainfluenza virus 1+2+3+4 Ab.IgM|Parainfluenza virus 1+2+3+4 Ab.IgM
C3482036|T201|COMP|70018-7|LNC|Staphylococcus haemolyticus DNA|Staphylococcus haemolyticus DNA
C3482037|T201|COMP|70019-5|LNC|Klebsiella oxytoca DNA|Klebsiella oxytoca DNA
C3482038|T201|COMP|70020-3|LNC|Bacteroides fragilis DNA|Bacteroides fragilis DNA
C3482040|T201|COMP|70106-0|LNC|Methotrexate^9th specimen|Methotrexate^9th specimen
C3482041|T201|COMP|70107-8|LNC|SERPINC1 gene mutations tested for|SERPINC1 gene mutations tested for
C3482043|T201|COMP|70108-6|LNC|Glutathione S-transferase T1 Ab|Glutathione S-transferase T1 Ab
C3482044|T201|COMP|70109-4|LNC|Number of chromosome 13 present|Number of chromosome 13 present
C3482045|T201|COMP|70110-2|LNC|Number of chromosome 18 present|Number of chromosome 18 present
C3482046|T201|COMP|70111-0|LNC|Number of chromosome 21 present|Number of chromosome 21 present
C3482079|T201|COMP|70664-8|LNC|Parathyrin.intact intraoperative percent change|Parathyrin.intact intraoperative percent change
C3482080|T201|COMP|70665-5|LNC|Cold agglutinin|Cold agglutinin
C3482099|T201|COMP|70021-1|LNC|Salmonella typhi DNA|Salmonella typhi DNA
C3482100|T201|COMP|70022-9|LNC|Candida albicans DNA|Candida albicans DNA
C3482101|T201|COMP|70023-7|LNC|Candida tropicalis DNA|Candida tropicalis DNA
C3482103|T201|COMP|70024-5|LNC|Candida parapsilosis DNA|Candida parapsilosis DNA
C3482105|T201|COMP|70025-2|LNC|Candida krusei DNA|Candida krusei DNA
C3482107|T201|COMP|70026-0|LNC|Candida glabrata DNA|Candida glabrata DNA
C3482108|T201|COMP|70027-8|LNC|Dermatophytes chitin synthase 1 (chs1) gene|Dermatophytes chitin synthase 1 (chs1) gene
C3482110|T201|COMP|70028-6|LNC|Megakaryocytic nuclei/100 leukocytes|Megakaryocytic nuclei/100 leukocytes
C3482112|T201|COMP|70032-8|LNC|Platelets.reticulated/platelets.total|Platelets.reticulated/platelets.total
C3482114|T201|COMP|70033-6|LNC|Ragocytes/100 leukocytes|Ragocytes/100 leukocytes
C3482116|T201|COMP|70034-4|LNC|Lipophages/100 leukocytes|Lipophages/100 leukocytes
C3482118|T201|COMP|70035-1|LNC|Siderophages/100 leukocytes|Siderophages/100 leukocytes
C3482120|T201|COMP|70036-9|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C3482121|T201|COMP|70037-7|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C3482122|T201|COMP|70038-5|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C3482123|T201|COMP|70039-3|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C3482124|T201|COMP|70040-1|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C3482125|T201|COMP|70041-9|LNC|FSHB gene.c.-211G>T|FSHB gene.c.-211G>T
C3482127|T201|COMP|70042-7|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C3482128|T201|COMP|70043-5|LNC|Mononuclear cells|Mononuclear cells
C3482129|T201|COMP|70044-3|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C3482130|T201|COMP|70045-0|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C3482131|T201|COMP|70046-8|LNC|Mononuclear cells|Mononuclear cells
C3482132|T201|COMP|70047-6|LNC|Mononuclear cells|Mononuclear cells
C3482133|T201|COMP|70048-4|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C3482134|T201|COMP|70049-2|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C3482135|T201|COMP|70050-0|LNC|Mononuclear cells|Mononuclear cells
C3482136|T201|COMP|70051-8|LNC|Multiple inhalant allergen Ab.IgE|Multiple inhalant allergen Ab.IgE
C3482137|T201|COMP|70052-6|LNC|Hantavirus hantaan Ab.IgG|Hantavirus hantaan Ab.IgG
C3482138|T201|COMP|70053-4|LNC|Hantavirus hantaan Ab.IgM|Hantavirus hantaan Ab.IgM
C3482139|T201|COMP|70054-2|LNC|Hantavirus dobrova Ab.IgM|Hantavirus dobrova Ab.IgM
C3482140|T201|COMP|70055-9|LNC|Hantavirus dobrova Ab.IgG|Hantavirus dobrova Ab.IgG
C3482141|T201|COMP|70056-7|LNC|Hantavirus saaremaa Ab.IgG|Hantavirus saaremaa Ab.IgG
C3482142|T201|COMP|70057-5|LNC|Hantavirus saaremaa Ab.IgM|Hantavirus saaremaa Ab.IgM
C3482143|T201|COMP|70058-3|LNC|Hantavirus puumala Ab.IgM|Hantavirus puumala Ab.IgM
C3482144|T201|COMP|70059-1|LNC|Hantavirus puumala Ab.IgG|Hantavirus puumala Ab.IgG
C3482145|T201|COMP|70060-9|LNC|Hantavirus seoul Ab.IgG|Hantavirus seoul Ab.IgG
C3482146|T201|COMP|70061-7|LNC|Human papilloma virus 16 & 18 DNA|Human papilloma virus 16 & 18 DNA
C3482147|T201|COMP|70065-8|LNC|Enterovirus Ag|Enterovirus Ag
C3482148|T201|COMP|70066-6|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C3482149|T201|COMP|70067-4|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C3482151|T201|COMP|70069-0|LNC|Streptococcus intermedius DNA|Streptococcus intermedius DNA
C3482152|T201|COMP|70070-8|LNC|Streptococcus anginosus DNA|Streptococcus anginosus DNA
C3482153|T201|COMP|70071-6|LNC|Streptococcus constellatus DNA|Streptococcus constellatus DNA
C3482154|T201|COMP|70072-4|LNC|Amyloid beta 40 peptide|Amyloid beta 40 peptide
C3482156|T201|COMP|70073-2|LNC|Amyloid beta 40 peptide|Amyloid beta 40 peptide
C3482157|T201|COMP|70074-0|LNC|Angiotensin II^supine|Angiotensin II^supine
C3482158|T201|COMP|70075-7|LNC|Interleukin 1 alpha|Interleukin 1 alpha
C3482159|T201|COMP|70076-5|LNC|Interleukin 1 alpha|Interleukin 1 alpha
C3482160|T201|COMP|70077-3|LNC|Interleukin 2|Interleukin 2
C3482161|T201|COMP|70078-1|LNC|Interleukin 2|Interleukin 2
C3482162|T201|COMP|70079-9|LNC|Interleukin 3|Interleukin 3
C3482163|T201|COMP|70080-7|LNC|Interleukin 3|Interleukin 3
C3482164|T201|COMP|70081-5|LNC|Interleukin 3|Interleukin 3
C3482165|T201|COMP|70082-3|LNC|Interleukin 4|Interleukin 4
C3482166|T201|COMP|70083-1|LNC|Interleukin 4|Interleukin 4
C3482167|T201|COMP|70084-9|LNC|Interleukin 5|Interleukin 5
C3482168|T201|COMP|70085-6|LNC|Interleukin 5|Interleukin 5
C3482169|T201|COMP|70086-4|LNC|Interleukin 7|Interleukin 7
C3482170|T201|COMP|70087-2|LNC|Interleukin 7|Interleukin 7
C3482171|T201|COMP|70088-0|LNC|Interleukin 7|Interleukin 7
C3482172|T201|COMP|70089-8|LNC|Interleukin 13|Interleukin 13
C3482173|T201|COMP|70090-6|LNC|Interleukin 13|Interleukin 13
C3482174|T201|COMP|70091-4|LNC|Prostaglandin E2|Prostaglandin E2
C3482175|T201|COMP|70092-2|LNC|Prostaglandin E1|Prostaglandin E1
C3482176|T201|COMP|70093-0|LNC|Prostaglandin E1|Prostaglandin E1
C3482177|T201|COMP|70094-8|LNC|Prostaglandin F2 alpha|Prostaglandin F2 alpha
C3482178|T201|COMP|70095-5|LNC|Prostaglandin F2 alpha|Prostaglandin F2 alpha
C3482179|T201|COMP|70096-3|LNC|Thyrotropin releasing hormone|Thyrotropin releasing hormone
C3482182|T201|COMP|70098-9|LNC|Methotrexate^10th specimen|Methotrexate^10th specimen
C3482183|T201|COMP|70099-7|LNC|Methotrexate^2nd specimen|Methotrexate^2nd specimen
C3482184|T201|COMP|70100-3|LNC|Methotrexate^3rd specimen|Methotrexate^3rd specimen
C3482185|T201|COMP|70101-1|LNC|Methotrexate^4th specimen|Methotrexate^4th specimen
C3482186|T201|COMP|70102-9|LNC|Methotrexate^5th specimen|Methotrexate^5th specimen
C3482187|T201|COMP|70103-7|LNC|Methotrexate^6th specimen|Methotrexate^6th specimen
C3482188|T201|COMP|70104-5|LNC|Methotrexate^7th specimen|Methotrexate^7th specimen
C3482189|T201|COMP|70105-2|LNC|Methotrexate^8th specimen|Methotrexate^8th specimen
C3482203|T201|COMP|70121-9|LNC|Francisella tularensis Ab.IgG|Francisella tularensis Ab.IgG
C3482204|T201|COMP|70122-7|LNC|Epithelial cells.squamous|Epithelial cells.squamous
C3482205|T201|COMP|70123-5|LNC|Epithelial cells.ciliated|Epithelial cells.ciliated
C3482206|T201|COMP|70124-3|LNC|Erythrocytes|Erythrocytes
C3482207|T201|COMP|70125-0|LNC|Yeast.hyphae|Yeast.hyphae
C3482208|T201|COMP|70126-8|LNC|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C3482214|T201|COMP|70131-8|LNC|Rickettsia typhus group Ab.IgG^1st specimen|Rickettsia typhus group Ab.IgG^1st specimen
C3482215|T201|COMP|70142-5|LNC|Benzodiazepines|Benzodiazepines
C3482216|T201|COMP|70143-3|LNC|Cannabinoids|Cannabinoids
C3482217|T201|COMP|70144-1|LNC|Cannabinoids|Cannabinoids
C3482218|T201|COMP|70149-0|LNC|Methadone|Methadone
C3482219|T201|COMP|70154-0|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C3482220|T201|COMP|70155-7|LNC|Barbiturates|Barbiturates
C3482234|T201|COMP|70165-6|LNC|Trichomonas vaginalis rRNA|Trichomonas vaginalis rRNA
C3482235|T201|COMP|70166-4|LNC|Trichomonas vaginalis rRNA|Trichomonas vaginalis rRNA
C3482236|T201|COMP|70167-2|LNC|Trichomonas vaginalis rRNA|Trichomonas vaginalis rRNA
C3482237|T201|COMP|70168-0|LNC|Hematocrit|Hematocrit
C3482238|T201|COMP|70169-8|LNC|Hematocrit|Hematocrit
C3482239|T201|COMP|70170-6|LNC|Erythrocytes.nucleated/100 cells|Erythrocytes.nucleated/100 cells
C3482240|T201|COMP|70171-4|LNC|Erythrocytes.nucleated/100 cells|Erythrocytes.nucleated/100 cells
C3482241|T201|COMP|70172-2|LNC|Neisseria meningitidis serogroup|Neisseria meningitidis serogroup
C3482242|T201|COMP|70173-0|LNC|JC virus Ab|JC virus Ab
C3482243|T201|COMP|70174-8|LNC|Dicarboxytetradecenoylcarnitine (C14:1-DC)|Dicarboxytetradecenoylcarnitine (C14:1-DC)
C3482244|T201|COMP|70175-5|LNC|Dicarboxytetradecenoylcarnitine (C14:1-DC)|Dicarboxytetradecenoylcarnitine (C14:1-DC)
C3482245|T201|COMP|70176-3|LNC|Dicarboxytetradecenoylcarnitine (C14:1-DC)|Dicarboxytetradecenoylcarnitine (C14:1-DC)
C3482246|T201|COMP|70177-1|LNC|Dicarboxytetradecenoylcarnitine (C14:1-DC)|Dicarboxytetradecenoylcarnitine (C14:1-DC)
C3482247|T201|COMP|70178-9|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C3482248|T201|COMP|70179-7|LNC|1-Methylhistidine|1-Methylhistidine
C3482249|T201|COMP|70180-5|LNC|Alpha aminoadipate|Alpha aminoadipate
C3482250|T201|COMP|70181-3|LNC|Alpha aminobutyrate|Alpha aminobutyrate
C3482266|T201|COMP|70204-3|LNC|Cholesterol.non HDL|Cholesterol.non HDL
C3482267|T201|COMP|70205-0|LNC|clonazePAM|clonazePAM
C3482268|T201|COMP|70206-8|LNC|Codeine|Codeine
C3482269|T201|COMP|70207-6|LNC|Estrogen|Estrogen
C3482270|T201|COMP|70208-4|LNC|Glucose^pre 100 g glucose PO|Glucose^pre 100 g glucose PO
C3482271|T201|COMP|70209-2|LNC|Haptoglobin|Haptoglobin
C3482272|T201|COMP|70210-0|LNC|Morphine|Morphine
C3482273|T201|COMP|70211-8|LNC|Mycophenolate|Mycophenolate
C3482274|T201|COMP|70212-6|LNC|Nordiazepam|Nordiazepam
C3482275|T201|COMP|70213-4|LNC|Nordiazepam|Nordiazepam
C3482276|T201|COMP|70214-2|LNC|Oxazepam|Oxazepam
C3482277|T201|COMP|70215-9|LNC|oxyCODONE|oxyCODONE
C3482278|T201|COMP|70216-7|LNC|Salicylates|Salicylates
C3482279|T201|COMP|70217-5|LNC|Thyroxine.free|Thyroxine.free
C3482280|T201|COMP|70218-3|LNC|Triglyceride|Triglyceride
C3482281|T201|COMP|70219-1|LNC|Basic metabolic 2008 panel with ionized calcium|Basic metabolic 2008 panel with ionized calcium
C3482290|T201|COMP|70239-9|LNC|Testosterone|Testosterone
C3482291|T201|COMP|70240-7|LNC|Testosterone.free|Testosterone.free
C3482292|T201|COMP|70241-5|LNC|HIV 1 RNA|HIV 1 RNA
C3482295|T201|COMP|70243-1|LNC|CLN3 gene exon 7+8 deletion|CLN3 gene exon 7+8 deletion
C3482297|T201|COMP|70244-9|LNC|CFTR gene.c.394delTT|CFTR gene.c.394delTT
C3482299|T201|COMP|70245-6|LNC|PAH gene.p.Arg408Trp|PAH gene.p.Arg408Trp
C3482300|T201|COMP|70246-4|LNC|CCR2 gene.p.Val64Ile|CCR2 gene.p.Val64Ile
C3482302|T201|COMP|70247-2|LNC|CCR5 gene.c.794_825del|CCR5 gene.c.794_825del
C3482304|T201|COMP|70248-0|LNC|GALT gene.p.Gln188Arg|GALT gene.p.Gln188Arg
C3482306|T201|COMP|70251-4|LNC|Pyruvate dehydrogenase Ab.IgG|Pyruvate dehydrogenase Ab.IgG
C3482307|T201|COMP|70252-2|LNC|Islet cell 512 Ab.IgG|Islet cell 512 Ab.IgG
C3482308|T201|COMP|70253-0|LNC|Islet cell 512 Ab.IgG|Islet cell 512 Ab.IgG
C3482309|T201|COMP|70254-8|LNC|Follitropin Ab.IgG|Follitropin Ab.IgG
C3482311|T201|COMP|70255-5|LNC|Follitropin Ab.IgA|Follitropin Ab.IgA
C3482313|T201|COMP|70256-3|LNC|Nuclear Ab.IgG|Nuclear Ab.IgG
C3482315|T201|COMP|70258-9|LNC|Amylase.pancreatic|Amylase.pancreatic
C3482316|T201|COMP|70259-7|LNC|Triglyceride.pericard fld/Triglyceride.serum|Triglyceride.pericard fld/Triglyceride.serum
C3482318|T201|COMP|70260-5|LNC|Triglyceride.periton fld/Triglyceride.serum|Triglyceride.periton fld/Triglyceride.serum
C3482320|T201|COMP|70261-3|LNC|Cholesterol.periton fld/Cholesterol.serum|Cholesterol.periton fld/Cholesterol.serum
C3482322|T201|COMP|70262-1|LNC|Amylase.periton fld/Amylase.serum|Amylase.periton fld/Amylase.serum
C3482324|T201|COMP|70263-9|LNC|Cholesterol.pericard fld/Cholesterol.serum|Cholesterol.pericard fld/Cholesterol.serum
C3482326|T201|COMP|70264-7|LNC|Creatinine.plr fld/Creatinine.serum|Creatinine.plr fld/Creatinine.serum
C3482328|T201|COMP|70265-4|LNC|Protein.pericard fld/Protein.serum|Protein.pericard fld/Protein.serum
C3482330|T201|COMP|70266-2|LNC|Creatinine.periton fld/Creatinine.serum|Creatinine.periton fld/Creatinine.serum
C3482332|T201|COMP|70267-0|LNC|Protein.periton fld/Protein.serum|Protein.periton fld/Protein.serum
C3482334|T201|COMP|70268-8|LNC|Cholesterol.plr fld/Cholesterol.serum|Cholesterol.plr fld/Cholesterol.serum
C3482336|T201|COMP|70269-6|LNC|Triglyceride.plr fld/Triglyceride.serum|Triglyceride.plr fld/Triglyceride.serum
C3482338|T201|COMP|70270-4|LNC|Amylase.pancreatic|Amylase.pancreatic
C3482344|T201|COMP|70275-3|LNC|t(X;11)(q13.1;q23)(FOXO4,MLL) fusion transcript|t(X;11)(q13.1;q23)(FOXO4,MLL) fusion transcript
C3482346|T201|COMP|70276-1|LNC|t(1;11)(p32;q23)(EPS15,MLL) fusion transcript|t(1;11)(p32;q23)(EPS15,MLL) fusion transcript
C3482348|T201|COMP|70277-9|LNC|t(3;5)(q25.1;q35.1)(MLF1,NPM1) fusion transcript|t(3;5)(q25.1;q35.1)(MLF1,NPM1) fusion transcript
C3482350|T201|COMP|70278-7|LNC|t(3;21)(q26;q22.3)(MECOM,RUNX1) fusion transcript|t(3;21)(q26;q22.3)(MECOM,RUNX1) fusion transcript
C3482352|T201|COMP|70279-5|LNC|t(5;17)(q25.1;q21.1)(NPM1,RARA) fusion transcript|t(5;17)(q25.1;q21.1)(NPM1,RARA) fusion transcript
C3482354|T201|COMP|70280-3|LNC|t(6;11)(q27;q23)(MLLT4,MLL) fusion transcript|t(6;11)(q27;q23)(MLLT4,MLL) fusion transcript
C3482356|T201|COMP|70281-1|LNC|t(9;9)(q34;q34)(NUP214,SET) fusion transcript|t(9;9)(q34;q34)(NUP214,SET) fusion transcript
C3482358|T201|COMP|70282-9|LNC|t(9;12)(q34.1;p13)(ABL1,ETV6) fusion transcript|t(9;12)(q34.1;p13)(ABL1,ETV6) fusion transcript
C3482360|T201|COMP|70283-7|LNC|t(11;17)(q23;q21)(MLL,MLLT6) fusion transcript|t(11;17)(q23;q21)(MLL,MLLT6) fusion transcript
C3482364|T201|COMP|70285-2|LNC|t(11;19)(q23;p13.1)(MLL,ELL) fusion transcript|t(11;19)(q23;p13.1)(MLL,ELL) fusion transcript
C3482366|T201|COMP|70286-0|LNC|t(12;22)(p13;q12.1)(ETV6,MN1) fusion transcript|t(12;22)(p13;q12.1)(ETV6,MN1) fusion transcript
C3482368|T201|COMP|70287-8|LNC|t(16;21)(p11.2;q22.3)(FUS,ERG) fusion transcript|t(16;21)(p11.2;q22.3)(FUS,ERG) fusion transcript
C3482370|T201|COMP|70288-6|LNC|t(17;19)(q22;p13.3)(HLF,TCF3) fusion transcript|t(17;19)(q22;p13.3)(HLF,TCF3) fusion transcript
C3482372|T201|COMP|70289-4|LNC|Del(1)(p32p32)(STIL,TAL1) fusion transcript|Del(1)(p32p32)(STIL,TAL1) fusion transcript
C3482376|T201|COMP|70292-8|LNC|Blastocystis hominis DNA|Blastocystis hominis DNA
C3482380|T201|COMP|70294-4|LNC|Entamoeba sp DNA|Entamoeba sp DNA
C3482382|T201|COMP|70295-1|LNC|Dientamoeba fragilis DNA|Dientamoeba fragilis DNA
C3482384|T201|COMP|70296-9|LNC|Plesiomonas shigelloides DNA|Plesiomonas shigelloides DNA
C3482410|T201|COMP|70666-3|LNC|Cold agglutinin|Cold agglutinin
C3482411|T201|COMP|70667-1|LNC|Cold agglutinin|Cold agglutinin
C3482453|T201|COMP|71425-3|LNC|Natriuretic peptide.B prohormone N-Terminal|Natriuretic peptide.B prohormone N-Terminal
C3482454|T201|COMP|71426-1|LNC|C reactive protein|C reactive protein
C3482455|T201|COMP|71427-9|LNC|Fibrin D-dimer FEU|Fibrin D-dimer FEU
C3482458|T201|COMP|71429-5|LNC|Campylobacter sp DNA.diarrheagenic|Campylobacter sp DNA.diarrheagenic
C3482460|T201|COMP|71430-3|LNC|oxyCODONE+Oxymorphone|oxyCODONE+Oxymorphone
C3482769|T201|COMP|70568-1|LNC|Plasmodium knowlesi DNA|Plasmodium knowlesi DNA
C3482770|T201|COMP|70569-9|LNC|Plasmodium sp Ag|Plasmodium sp Ag
C3483025|T201|COMP|70850-3|LNC|Burkholderia mallei|Burkholderia mallei
C3483026|T201|COMP|70851-1|LNC|Burkholderia pseudomallei|Burkholderia pseudomallei
C3483027|T201|COMP|70852-9|LNC|Burkholderia pseudomallei DNA|Burkholderia pseudomallei DNA
C3483029|T201|COMP|70853-7|LNC|Burkholderia mallei DNA|Burkholderia mallei DNA
C3483031|T201|COMP|70854-5|LNC|Burkholderia mallei Ag|Burkholderia mallei Ag
C3483032|T201|COMP|70855-2|LNC|Burkholderia pseudomallei Ag|Burkholderia pseudomallei Ag
C3483033|T201|COMP|70856-0|LNC|Rabies virus Ab|Rabies virus Ab
C3483034|T201|COMP|70857-8|LNC|Rabies virus Ab|Rabies virus Ab
C3483035|T201|COMP|70858-6|LNC|Rabies virus Ab|Rabies virus Ab
C3483036|T201|COMP|70859-4|LNC|Rabies virus Ab|Rabies virus Ab
C3483037|T201|COMP|70860-2|LNC|Rabies virus Ab.IgG|Rabies virus Ab.IgG
C3483038|T201|COMP|70861-0|LNC|Rabies virus Ab.IgG|Rabies virus Ab.IgG
C3483039|T201|COMP|70862-8|LNC|Rabies virus Ab.IgM|Rabies virus Ab.IgM
C3483040|T201|COMP|70863-6|LNC|Rabies virus Ab.IgM|Rabies virus Ab.IgM
C3483041|T201|COMP|70864-4|LNC|Rabies virus Ab.IgM|Rabies virus Ab.IgM
C3483042|T201|COMP|70865-1|LNC|Rabies virus Ab.IgM|Rabies virus Ab.IgM
C3483043|T201|COMP|70866-9|LNC|Rabies virus strain identified|Rabies virus strain identified
C3483044|T201|COMP|70867-7|LNC|Rabies virus strain identified|Rabies virus strain identified
C3483122|T201|COMP|70907-1|LNC|Cryptococcus sp rRNA gene|Cryptococcus sp rRNA gene
C3483124|T201|COMP|70908-9|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C3483125|T201|COMP|70909-7|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C3483126|T201|COMP|70910-5|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C3483127|T201|COMP|70911-3|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C3483181|T201|COMP|70970-9|LNC|Cryoglobulin|Cryoglobulin
C3483285|T201|COMP|71358-6|LNC|GJB3 gene targeted mutation analysis|GJB3 gene targeted mutation analysis
C3483287|T201|COMP|71359-4|LNC|Y chromosome AZFa region deletion|Y chromosome AZFa region deletion
C3483289|T201|COMP|71360-2|LNC|Y chromosome AZFb region deletion|Y chromosome AZFb region deletion
C3483291|T201|COMP|71361-0|LNC|Y chromosome AZFc region deletion|Y chromosome AZFc region deletion
C3483295|T201|COMP|71365-1|LNC|Alkaline phosphatase.intestinal 2|Alkaline phosphatase.intestinal 2
C3483296|T201|COMP|71366-9|LNC|Alkaline phosphatase.intestinal 3|Alkaline phosphatase.intestinal 3
C3483297|T201|COMP|71367-7|LNC|Alkaline phosphatase.placental 2|Alkaline phosphatase.placental 2
C3483299|T201|COMP|71368-5|LNC|Desmosome Ab.IgG|Desmosome Ab.IgG
C3483301|T201|COMP|71883-3|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C3483302|T201|COMP|71884-1|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C3483303|T201|COMP|71885-8|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C3483304|T201|COMP|71886-6|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C3483305|T201|COMP|71887-4|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C3483306|T201|COMP|71888-2|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C3483307|T201|COMP|71889-0|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C3483308|T201|COMP|71890-8|LNC|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C3483310|T201|COMP|71892-4|LNC|Cortisone^AM peak specimen|Cortisone^AM peak specimen
C3483457|T201|COMP|71592-0|LNC|Hemoglobinopathies conditions suspected|Hemoglobinopathies conditions suspected
C3483458|T201|COMP|71593-8|LNC|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C3483632|T201|COMP|71355-2|LNC|SLC26A5 gene.c.-53-2A>G|SLC26A5 gene.c.-53-2A>G
C3483633|T201|COMP|71356-0|LNC|TPMT gene.c.238G>C+460G>A+719A>G|TPMT gene.c.238G>C+460G>A+719A>G
C3483634|T201|COMP|71357-8|LNC|PDGFRA gene exon 18 targeted mutation analysis|PDGFRA gene exon 18 targeted mutation analysis
C3483636|T201|COMP|71369-3|LNC|Neutrophils.dysplastic|Neutrophils.dysplastic
C3483646|T201|COMP|71377-6|LNC|Legionella sp|Legionella sp
C3483647|T201|COMP|71378-4|LNC|Leptospira sp|Leptospira sp
C3483655|T201|COMP|71386-7|LNC|Hepcidin 25 peptide|Hepcidin 25 peptide
C3483656|T201|COMP|71387-5|LNC|Spermatozoa.motile^post ejaculate|Spermatozoa.motile^post ejaculate
C3483754|T201|COMP|71456-8|LNC|Nitrofural|Nitrofural
C3483867|T201|COMP|71689-4|LNC|Mononuclear cells|Mononuclear cells
C3483868|T201|COMP|71690-2|LNC|Nucleated cells|Nucleated cells
C3483869|T201|COMP|71691-0|LNC|Hematopoietic progenitor cells|Hematopoietic progenitor cells
C3483870|T201|COMP|71692-8|LNC|Platelets.reticulated|Platelets.reticulated
C3483871|T201|COMP|71693-6|LNC|Platelets.reticulated/100 platelets|Platelets.reticulated/100 platelets
C3483872|T201|COMP|71694-4|LNC|Hemoglobin|Hemoglobin
C3483873|T201|COMP|71695-1|LNC|Granulocytes.immature/100 leukocytes|Granulocytes.immature/100 leukocytes
C3483874|T201|COMP|71696-9|LNC|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C3483875|T201|COMP|71697-7|LNC|Mononuclear cells/100 leukocytes|Mononuclear cells/100 leukocytes
C3483876|T201|COMP|71698-5|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C3483877|T201|COMP|71699-3|LNC|Flavivirus Ag|Flavivirus Ag
C3483879|T201|COMP|71700-9|LNC|Rotavirus RNA|Rotavirus RNA
C3483880|T201|COMP|71701-7|LNC|Rotavirus dsRNA|Rotavirus dsRNA
C3483881|T201|COMP|71702-5|LNC|Rotavirus dsRNA|Rotavirus dsRNA
C3483882|T201|COMP|71843-7|LNC|Oxygen saturation|Oxygen saturation
C3483883|T201|COMP|71844-5|LNC|Oxygen saturation|Oxygen saturation
C3483884|T201|COMP|71845-2|LNC|Oxygen saturation|Oxygen saturation
C3483885|T201|COMP|71846-0|LNC|Oxygen saturation|Oxygen saturation
C3483886|T201|COMP|71847-8|LNC|Oxygen saturation|Oxygen saturation
C3483887|T201|COMP|71848-6|LNC|Oxygen saturation|Oxygen saturation
C3483888|T201|COMP|71849-4|LNC|Oxygen saturation|Oxygen saturation
C3483889|T201|COMP|71850-2|LNC|Oxygen saturation|Oxygen saturation
C3483890|T201|COMP|71851-0|LNC|Oxygen saturation|Oxygen saturation
C3483891|T201|COMP|71852-8|LNC|Oxygen saturation|Oxygen saturation
C3483896|T201|COMP|71853-6|LNC|Oxygen saturation|Oxygen saturation
C3483897|T201|COMP|71854-4|LNC|Deoxyhemoglobin/Hemoglobin.total|Deoxyhemoglobin/Hemoglobin.total
C3483898|T201|COMP|71855-1|LNC|Hemoglobin.other/Hemoglobin.total|Hemoglobin.other/Hemoglobin.total
C3483899|T201|COMP|71856-9|LNC|Hemoglobin.other/Hemoglobin.total|Hemoglobin.other/Hemoglobin.total
C3483900|T201|COMP|71857-7|LNC|Hemoglobin S/Hemoglobin.total|Hemoglobin S/Hemoglobin.total
C3483901|T201|COMP|71858-5|LNC|Hemoglobin S/Hemoglobin.total|Hemoglobin S/Hemoglobin.total
C3483904|T201|COMP|72111-8|LNC|Sapovirus RNA|Sapovirus RNA
C3483920|T201|COMP|71703-3|LNC|Rotavirus Ab.IgG|Rotavirus Ab.IgG
C3483921|T201|COMP|71704-1|LNC|Rotavirus Ab.IgA|Rotavirus Ab.IgA
C3483922|T201|COMP|71705-8|LNC|Rotavirus Ab|Rotavirus Ab
C3483923|T201|COMP|71706-6|LNC|Marburg virus Ab.IgM|Marburg virus Ab.IgM
C3483924|T201|COMP|71707-4|LNC|Marburg virus Ab.IgG|Marburg virus Ab.IgG
C3483925|T201|COMP|71708-2|LNC|Marburg virus Ag|Marburg virus Ag
C3483926|T201|COMP|71709-0|LNC|Lassa virus Ab.IgM|Lassa virus Ab.IgM
C3483927|T201|COMP|71710-8|LNC|Lassa virus Ab.IgG|Lassa virus Ab.IgG
C3483928|T201|COMP|71711-6|LNC|Ebola virus Ab.IgM|Ebola virus Ab.IgM
C3483930|T201|COMP|71712-4|LNC|Ebola virus Ab.IgM|Ebola virus Ab.IgM
C3483931|T201|COMP|71713-2|LNC|Pyruvate kinase|Pyruvate kinase
C3483932|T201|COMP|71714-0|LNC|Brucella abortus Ab|Brucella abortus Ab
C3483933|T201|COMP|71715-7|LNC|Brucella abortus Ab.IgG1+IgG2|Brucella abortus Ab.IgG1+IgG2
C3483935|T201|COMP|71716-5|LNC|Brucella suis Ab|Brucella suis Ab
C3483936|T201|COMP|71717-3|LNC|Brucella suis Ab|Brucella suis Ab
C3483937|T201|COMP|71718-1|LNC|Enterococcus sp DNA|Enterococcus sp DNA
C3483938|T201|COMP|71719-9|LNC|Mycobacterium avium complex DNA|Mycobacterium avium complex DNA
C3483984|T201|COMP|71759-5|LNC|Rotavirus RNA|Rotavirus RNA
C3483985|T201|COMP|71760-3|LNC|Rotavirus identified|Rotavirus identified
C3483986|T201|COMP|71761-1|LNC|Rotavirus identified|Rotavirus identified
C3483987|T201|COMP|71762-9|LNC|Rotavirus Ab.IgA|Rotavirus Ab.IgA
C3483988|T201|COMP|71763-7|LNC|Rotavirus Ab.IgA|Rotavirus Ab.IgA
C3483989|T201|COMP|71764-5|LNC|Rotavirus Ab|Rotavirus Ab
C3483990|T201|COMP|71765-2|LNC|Rotavirus Ab|Rotavirus Ab
C3483992|T201|COMP|71767-8|LNC|Ebola virus Ab.IgG|Ebola virus Ab.IgG
C3483994|T201|COMP|71768-6|LNC|Ebola virus Ag|Ebola virus Ag
C3483995|T201|COMP|71769-4|LNC|Marburg virus Ab.IgG|Marburg virus Ab.IgG
C3483996|T201|COMP|71770-2|LNC|Ebola virus Ab.IgG|Ebola virus Ab.IgG
C3483997|T201|COMP|71771-0|LNC|Marburg virus Ab.IgM|Marburg virus Ab.IgM
C3483998|T201|COMP|71772-8|LNC|Mitogen stimulated gamma interferon|Mitogen stimulated gamma interferon
C3484002|T201|COMP|71776-9|LNC|Gamma interferon background|Gamma interferon background
C3484005|T201|COMP|71778-5|LNC|Rift valley fever virus Ag|Rift valley fever virus Ag
C3484006|T201|COMP|71779-3|LNC|Rift valley fever virus Ab.IgM|Rift valley fever virus Ab.IgM
C3484007|T201|COMP|71780-1|LNC|Rift valley fever virus Ab.IgG|Rift valley fever virus Ab.IgG
C3484008|T201|COMP|71781-9|LNC|Rift valley fever virus Ab.IgM|Rift valley fever virus Ab.IgM
C3484009|T201|COMP|71782-7|LNC|Yellow fever virus Ab.IgM|Yellow fever virus Ab.IgM
C3484010|T201|COMP|71783-5|LNC|Yellow fever virus Ab|Yellow fever virus Ab
C3484011|T201|COMP|71784-3|LNC|Rift valley fever virus Ab.IgG|Rift valley fever virus Ab.IgG
C3484016|T201|COMP|71788-4|LNC|Neisseria meningitidis DNA|Neisseria meningitidis DNA
C3484019|T201|COMP|71790-0|LNC|Calcium|Calcium
C3484020|T201|COMP|71792-6|LNC|Procollagen type III.N-terminal propeptide|Procollagen type III.N-terminal propeptide
C3484021|T201|COMP|71793-4|LNC|Treponema pallidum Ab|Treponema pallidum Ab
C3484025|T201|COMP|71797-5|LNC|Protoporphyrin.zinc|Protoporphyrin.zinc
C3484034|T201|COMP|71804-9|LNC|Serotonin|Serotonin
C3484035|T201|COMP|71805-6|LNC|Cortisol.free/Cortisone.free|Cortisol.free/Cortisone.free
C3484058|T201|COMP|71828-8|LNC|Hematocrit|Hematocrit
C3484059|T201|COMP|71829-6|LNC|Hematocrit|Hematocrit
C3484060|T201|COMP|71830-4|LNC|Hematocrit|Hematocrit
C3484061|T201|COMP|71831-2|LNC|Hematocrit|Hematocrit
C3484062|T201|COMP|71832-0|LNC|Hematocrit|Hematocrit
C3484063|T201|COMP|71833-8|LNC|Hematocrit|Hematocrit
C3484064|T201|COMP|71834-6|LNC|Cryoglobulin/Serum.total|Cryoglobulin/Serum.total
C3484066|T201|COMP|71836-1|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C3484067|T201|COMP|71837-9|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C3484068|T201|COMP|71838-7|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C3484069|T201|COMP|71839-5|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C3484070|T201|COMP|71840-3|LNC|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C3484071|T201|COMP|71841-1|LNC|Oxygen saturation|Oxygen saturation
C3484072|T201|COMP|71842-9|LNC|Oxygen saturation|Oxygen saturation
C3484073|T201|COMP|71859-3|LNC|Hemoglobin S/Hemoglobin.total|Hemoglobin S/Hemoglobin.total
C3484074|T201|COMP|71860-1|LNC|Hemoglobin M/Hemoglobin.total|Hemoglobin M/Hemoglobin.total
C3484075|T201|COMP|71861-9|LNC|Hemoglobin Lepore/Hemoglobin.total|Hemoglobin Lepore/Hemoglobin.total
C3484076|T201|COMP|71862-7|LNC|Hemoglobin H/Hemoglobin.total|Hemoglobin H/Hemoglobin.total
C3484077|T201|COMP|71863-5|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C3484078|T201|COMP|71864-3|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C3484079|T201|COMP|71865-0|LNC|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C3484080|T201|COMP|71866-8|LNC|Hemoglobin E/Hemoglobin.total|Hemoglobin E/Hemoglobin.total
C3484081|T201|COMP|71867-6|LNC|Hemoglobin D/Hemoglobin.total|Hemoglobin D/Hemoglobin.total
C3484082|T201|COMP|71868-4|LNC|Hemoglobin D/Hemoglobin.total|Hemoglobin D/Hemoglobin.total
C3484083|T201|COMP|71869-2|LNC|Hemoglobin C/Hemoglobin.total|Hemoglobin C/Hemoglobin.total
C3484084|T201|COMP|71870-0|LNC|Hemoglobin C/Hemoglobin.total|Hemoglobin C/Hemoglobin.total
C3484085|T201|COMP|71871-8|LNC|Hemoglobin Barts/Hemoglobin.total|Hemoglobin Barts/Hemoglobin.total
C3484086|T201|COMP|71872-6|LNC|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C3484087|T201|COMP|71873-4|LNC|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C3484088|T201|COMP|71874-2|LNC|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C3484089|T201|COMP|71875-9|LNC|Hemoglobin A1c/Hemoglobin.total|Hemoglobin A1c/Hemoglobin.total
C3484090|T201|COMP|71876-7|LNC|Hemoglobin A/Hemoglobin.total|Hemoglobin A/Hemoglobin.total
C3484091|T201|COMP|71877-5|LNC|Hemoglobin A/Hemoglobin.total|Hemoglobin A/Hemoglobin.total
C3484092|T201|COMP|71878-3|LNC|Hemoglobin A/Hemoglobin.total|Hemoglobin A/Hemoglobin.total
C3484093|T201|COMP|71879-1|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C3484094|T201|COMP|71880-9|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C3484095|T201|COMP|71881-7|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C3484096|T201|COMP|71882-5|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C3484097|T201|COMP|71893-2|LNC|Cortisone^PM trough specimen|Cortisone^PM trough specimen
C3484098|T201|COMP|71894-0|LNC|Cortisone.free|Cortisone.free
C3484229|T201|COMP|72103-5|LNC|Acute & chronic leukemia fusion transcript panel|Acute & chronic leukemia fusion transcript panel
C3484387|T201|COMP|20993-2|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C3484388|T201|COMP|23908-7|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C3484389|T201|COMP|17297-3|LNC|Mycobacterium tuberculosis rRNA|Mycobacterium tuberculosis rRNA
C3494486|T201|COMP|71791-8|LNC|Metanephrines|Metanephrines
C3496299|T201|COMP|72512-7|LNC|VKORC1 gene targeted mutation analysis|VKORC1 gene targeted mutation analysis
C3496495|T201|COMP|72199-3|LNC|HEDIS 2013 panel|HEDIS 2013 panel
C3533356|T201|COMP|72627-3|LNC|Barbiturates|Barbiturates
C3533357|T201|COMP|72457-5|LNC|Desmin Ab|Desmin Ab
C3533358|T201|COMP|72433-6|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C3533361|T201|COMP|72824-6|LNC|Del(17)(p13)|Del(17)(p13)
C3533362|T201|COMP|72823-8|LNC|Staphylococcus aureus enterotoxin C sec gene|Staphylococcus aureus enterotoxin C sec gene
C3533363|T201|COMP|72822-0|LNC|Staphylococcus aureus enterotoxin D sed gene|Staphylococcus aureus enterotoxin D sed gene
C3533364|T201|COMP|72821-2|LNC|Creatinine|Creatinine
C3533365|T201|COMP|72820-4|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C3533366|T201|COMP|72819-6|LNC|Acetaminophen/Creatinine|Acetaminophen/Creatinine
C3533367|T201|COMP|72818-8|LNC|AM-2201 4-hydroxypentyl/Creatinine|AM-2201 4-hydroxypentyl/Creatinine
C3533368|T201|COMP|72817-0|LNC|AM-2201 4-hydroxypentyl|AM-2201 4-hydroxypentyl
C3533369|T201|COMP|72816-2|LNC|DOPamine|DOPamine
C3533370|T201|COMP|72815-4|LNC|DULoxetine/Creatinine|DULoxetine/Creatinine
C3533371|T201|COMP|72814-7|LNC|DULoxetine|DULoxetine
C3533372|T201|COMP|72813-9|LNC|FLUoxetine/Creatinine|FLUoxetine/Creatinine
C3533373|T201|COMP|72812-1|LNC|Norfluoxetine/Creatinine|Norfluoxetine/Creatinine
C3533374|T201|COMP|72811-3|LNC|Gabapentin/Creatinine|Gabapentin/Creatinine
C3533375|T201|COMP|72810-5|LNC|Gabapentin|Gabapentin
C3533376|T201|COMP|72809-7|LNC|JWH-018 carboxylated/Creatinine|JWH-018 carboxylated/Creatinine
C3533377|T201|COMP|72808-9|LNC|JWH-018 carboxylated|JWH-018 carboxylated
C3533378|T201|COMP|72807-1|LNC|JWH-073 carboxylated/Creatinine|JWH-073 carboxylated/Creatinine
C3533379|T201|COMP|72806-3|LNC|JWH-073 carboxylated|JWH-073 carboxylated
C3533380|T201|COMP|72805-5|LNC|JWH-210 5-carboxypentyl/Creatinine|JWH-210 5-carboxypentyl/Creatinine
C3533381|T201|COMP|72804-8|LNC|JWH-210 5-carboxypentyl|JWH-210 5-carboxypentyl
C3533382|T201|COMP|72803-0|LNC|JWH-250 5-carboxypentyl/Creatinine|JWH-250 5-carboxypentyl/Creatinine
C3533383|T201|COMP|72802-2|LNC|JWH-250 5-carboxypentyl|JWH-250 5-carboxypentyl
C3533384|T201|COMP|72801-4|LNC|Ketamine/Creatinine|Ketamine/Creatinine
C3533385|T201|COMP|72800-6|LNC|Norketamine/Creatinine|Norketamine/Creatinine
C3533386|T201|COMP|72799-0|LNC|Norketamine|Norketamine
C3533387|T201|COMP|72798-2|LNC|Methylenedioxypyrovalerone/Creatinine|Methylenedioxypyrovalerone/Creatinine
C3533388|T201|COMP|72797-4|LNC|Methylenedioxypyrovalerone|Methylenedioxypyrovalerone
C3533389|T201|COMP|72796-6|LNC|Mephedrone/Creatinine|Mephedrone/Creatinine
C3533390|T201|COMP|72795-8|LNC|Mephedrone|Mephedrone
C3533391|T201|COMP|72794-1|LNC|Methylone/Creatinine|Methylone/Creatinine
C3533392|T201|COMP|72793-3|LNC|Methylone|Methylone
C3533393|T201|COMP|72792-5|LNC|Methylphenidate/Creatinine|Methylphenidate/Creatinine
C3533394|T201|COMP|72791-7|LNC|Alpha-Phenyl-2-Piperidine acetate/Creatinine|Alpha-Phenyl-2-Piperidine acetate/Creatinine
C3533395|T201|COMP|72790-9|LNC|Alpha-Phenyl-2-Piperidine acetate|Alpha-Phenyl-2-Piperidine acetate
C3533396|T201|COMP|72789-1|LNC|Naltrexone/Creatinine|Naltrexone/Creatinine
C3533397|T201|COMP|72788-3|LNC|6-Beta naltrexone/Creatinine|6-Beta naltrexone/Creatinine
C3533398|T201|COMP|72787-5|LNC|6-Beta naltrexone|6-Beta naltrexone
C3533399|T201|COMP|72786-7|LNC|Cotinine|Cotinine
C3533400|T201|COMP|72785-9|LNC|PARoxetine/Creatinine|PARoxetine/Creatinine
C3533401|T201|COMP|72784-2|LNC|PARoxetine|PARoxetine
C3533402|T201|COMP|72783-4|LNC|JWH-018 pentanoate/Creatinine|JWH-018 pentanoate/Creatinine
C3533403|T201|COMP|72782-6|LNC|JWH-018 pentanoate|JWH-018 pentanoate
C3533404|T201|COMP|72781-8|LNC|JWH-018 pentanol/Creatinine|JWH-018 pentanol/Creatinine
C3533405|T201|COMP|72780-0|LNC|JWH-018 pentanol|JWH-018 pentanol
C3533406|T201|COMP|72779-2|LNC|JWH-073 butanoate/Creatinine|JWH-073 butanoate/Creatinine
C3533407|T201|COMP|72778-4|LNC|JWH-073 butanoate|JWH-073 butanoate
C3533408|T201|COMP|72757-8|LNC|Benzodiazepines|Benzodiazepines
C3533409|T201|COMP|72756-0|LNC|ALPRAZolam|ALPRAZolam
C3533410|T201|COMP|72755-2|LNC|clonazePAM|clonazePAM
C3533411|T201|COMP|72754-5|LNC|LORazepam|LORazepam
C3533412|T201|COMP|72753-7|LNC|HYDROcodone|HYDROcodone
C3533413|T201|COMP|72752-9|LNC|Morphine|Morphine
C3533414|T201|COMP|72751-1|LNC|oxyCODONE|oxyCODONE
C3533415|T201|COMP|72750-3|LNC|oxyCODONE|oxyCODONE
C3533416|T201|COMP|72749-5|LNC|Meperidine|Meperidine
C3533417|T201|COMP|72748-7|LNC|Meprobamate|Meprobamate
C3533418|T201|COMP|72747-9|LNC|N-Nortramadol|N-Nortramadol
C3533419|T201|COMP|72746-1|LNC|Norbuprenorphine|Norbuprenorphine
C3533420|T201|COMP|72745-3|LNC|Norfentanyl|Norfentanyl
C3533421|T201|COMP|72744-6|LNC|Norhydrocodone|Norhydrocodone
C3533422|T201|COMP|72743-8|LNC|Normeperidine|Normeperidine
C3533423|T201|COMP|72742-0|LNC|Noroxycodone|Noroxycodone
C3533424|T201|COMP|72741-2|LNC|Nortramadol|Nortramadol
C3533425|T201|COMP|72740-4|LNC|traMADol|traMADol
C3533426|T201|COMP|72739-6|LNC|Nordiazepam|Nordiazepam
C3533427|T201|COMP|72738-8|LNC|Temazepam|Temazepam
C3533428|T201|COMP|72737-0|LNC|Cocaine|Cocaine
C3533429|T201|COMP|72736-2|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C3533430|T201|COMP|72735-4|LNC|Methamphetamine|Methamphetamine
C3533431|T201|COMP|72734-7|LNC|Methadone|Methadone
C3533432|T201|COMP|72733-9|LNC|HYDROmorphone|HYDROmorphone
C3533433|T201|COMP|72732-1|LNC|Mitragynine|Mitragynine
C3533434|T201|COMP|72731-3|LNC|7-Hydroxymitragynine|7-Hydroxymitragynine
C3533435|T201|COMP|72730-5|LNC|Mitragynine/Creatinine|Mitragynine/Creatinine
C3533436|T201|COMP|72729-7|LNC|7-Hydroxymitragynine/Creatinine|7-Hydroxymitragynine/Creatinine
C3533437|T201|COMP|72728-9|LNC|Del(13)(q14)|Del(13)(q14)
C3533438|T201|COMP|72727-1|LNC|Del(13)(q14) & del(17)(p13)|Del(13)(q14) & del(17)(p13)
C3533439|T201|COMP|72726-3|LNC|t(4;14)(p16;q32)(FGFR3,IGH) fusion transcript|t(4;14)(p16;q32)(FGFR3,IGH) fusion transcript
C3533440|T201|COMP|72725-5|LNC|t(11;14)(q13.2;q32)(MYEOV,IGH) fusion transcript|t(11;14)(q13.2;q32)(MYEOV,IGH) fusion transcript
C3533441|T201|COMP|72724-8|LNC|PM-SCL-75 Ab.IgG|PM-SCL-75 Ab.IgG
C3533442|T201|COMP|72723-0|LNC|Base excess.100% oxygenated^^standard|Base excess.100% oxygenated^^standard
C3533443|T201|COMP|72722-2|LNC|Base excess.100% oxygenated^^standard|Base excess.100% oxygenated^^standard
C3533444|T201|COMP|72721-4|LNC|Base excess.100% oxygenated^^standard|Base excess.100% oxygenated^^standard
C3533445|T201|COMP|72720-6|LNC|Base excess.100% oxygenated^^standard|Base excess.100% oxygenated^^standard
C3533446|T201|COMP|72697-6|LNC|CYP3A5 gene.c.6986A>G(*3)|CYP3A5 gene.c.6986A>G(*3)
C3533447|T201|COMP|72696-8|LNC|SLC40A1 gene targeted mutation analysis|SLC40A1 gene targeted mutation analysis
C3533448|T201|COMP|72695-0|LNC|Erythrocyte enzyme panel|Erythrocyte enzyme panel
C3533449|T201|COMP|72694-3|LNC|Cholinesterase activity panel|Cholinesterase activity panel
C3533450|T201|COMP|72679-4|LNC|Bile acid|Bile acid
C3533451|T201|COMP|72678-6|LNC|Venlafaxine+Norvenlafaxine^trough|Venlafaxine+Norvenlafaxine^trough
C3533452|T201|COMP|72677-8|LNC|Salicylates^trough|Salicylates^trough
C3533453|T201|COMP|72676-0|LNC|Sirolimus^trough|Sirolimus^trough
C3533454|T201|COMP|72675-2|LNC|Sotalol^trough|Sotalol^trough
C3533455|T201|COMP|72674-5|LNC|Sulfamethoxazole^trough|Sulfamethoxazole^trough
C3533456|T201|COMP|72673-7|LNC|Theophylline^trough|Theophylline^trough
C3533457|T201|COMP|72672-9|LNC|traZODone^trough|traZODone^trough
C3533458|T201|COMP|72671-1|LNC|Everolimus^trough|Everolimus^trough
C3533460|T201|COMP|72669-5|LNC|Mianserin^trough|Mianserin^trough
C3533461|T201|COMP|72668-7|LNC|Mirtazapine^trough|Mirtazapine^trough
C3533462|T201|COMP|72667-9|LNC|Mycophenolate^trough|Mycophenolate^trough
C3533463|T201|COMP|72666-1|LNC|Nitrazepam^trough|Nitrazepam^trough
C3533464|T201|COMP|72665-3|LNC|Trans,trans-muconate|Trans,trans-muconate
C3533465|T201|COMP|72664-6|LNC|Phosphofructokinase|Phosphofructokinase
C3533466|T201|COMP|72663-8|LNC|Bisphosphoglycerate mutase|Bisphosphoglycerate mutase
C3533467|T201|COMP|72662-0|LNC|Extrinsic coagulation factor activity 4 panel|Extrinsic coagulation factor activity 4 panel
C3533468|T201|COMP|72661-2|LNC|Intrinsic coagulation factor activity 4 panel|Intrinsic coagulation factor activity 4 panel
C3533469|T201|COMP|72660-4|LNC|Beta-trace protein|Beta-trace protein
C3533470|T201|COMP|72659-6|LNC|OXcarbazepine^trough|OXcarbazepine^trough
C3533471|T201|COMP|72658-8|LNC|PARoxetine^trough|PARoxetine^trough
C3533472|T201|COMP|72657-0|LNC|Procainamide^trough|Procainamide^trough
C3533473|T201|COMP|72656-2|LNC|risperiDONE^trough|risperiDONE^trough
C3533474|T201|COMP|72649-7|LNC|Glucose.serum-glucose.perition fld|Glucose.serum-glucose.perition fld
C3533475|T201|COMP|72648-9|LNC|Glucose.serum-glucose.synv fld|Glucose.serum-glucose.synv fld
C3533476|T201|COMP|72647-1|LNC|Albumin.serum-albumin.plr fld|Albumin.serum-albumin.plr fld
C3533477|T201|COMP|72646-3|LNC|Albumin.serum-albumin.pericard fld|Albumin.serum-albumin.pericard fld
C3533482|T201|COMP|72635-6|LNC|PENTobarbital|PENTobarbital
C3533483|T201|COMP|72634-9|LNC|Temazepam|Temazepam
C3533484|T201|COMP|72633-1|LNC|Benzodiazepines|Benzodiazepines
C3533485|T201|COMP|72632-3|LNC|Butalbital|Butalbital
C3533486|T201|COMP|72631-5|LNC|Amobarbital|Amobarbital
C3533487|T201|COMP|72630-7|LNC|PENTobarbital|PENTobarbital
C3533488|T201|COMP|72629-9|LNC|Secobarbital|Secobarbital
C3533489|T201|COMP|72628-1|LNC|PHENobarbital|PHENobarbital
C3533490|T201|COMP|72626-5|LNC|Methadone|Methadone
C3533491|T201|COMP|72625-7|LNC|Dabigatran|Dabigatran
C3533492|T201|COMP|72624-0|LNC|Rivaroxaban|Rivaroxaban
C3533493|T201|COMP|72623-2|LNC|inFLIXimab Ab|inFLIXimab Ab
C3533494|T201|COMP|72622-4|LNC|Propoxyphene|Propoxyphene
C3533495|T201|COMP|72621-6|LNC|Propoxyphene|Propoxyphene
C3533496|T201|COMP|72620-8|LNC|Norpropoxyphene|Norpropoxyphene
C3533497|T201|COMP|72619-0|LNC|Norpropoxyphene|Norpropoxyphene
C3533498|T201|COMP|72618-2|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C3533499|T201|COMP|72617-4|LNC|Propoxyphene|Propoxyphene
C3533500|T201|COMP|72616-6|LNC|Benzodiazepines|Benzodiazepines
C3533501|T201|COMP|72615-8|LNC|Nordiazepam|Nordiazepam
C3533502|T201|COMP|72614-1|LNC|Oxazepam|Oxazepam
C3533503|T201|COMP|72613-3|LNC|Oxazepam|Oxazepam
C3533504|T201|COMP|72612-5|LNC|ALPRAZolam|ALPRAZolam
C3533505|T201|COMP|72611-7|LNC|diazePAM|diazePAM
C3533506|T201|COMP|72610-9|LNC|diazePAM|diazePAM
C3533507|T201|COMP|72609-1|LNC|Nonsteroidal antiinflammatory drugs|Nonsteroidal antiinflammatory drugs
C3533508|T201|COMP|72608-3|LNC|Apixaban|Apixaban
C3533509|T201|COMP|72607-5|LNC|Streptococcus agalactiae|Streptococcus agalactiae
C3533510|T201|COMP|72606-7|LNC|Hepatitis D virus genotype|Hepatitis D virus genotype
C3533511|T201|COMP|72605-9|LNC|Cytomegalovirus glycoprotein genotype|Cytomegalovirus glycoprotein genotype
C3533512|T201|COMP|72604-2|LNC|Insulin^4.5H post 75 g glucose PO|Insulin^4.5H post 75 g glucose PO
C3533513|T201|COMP|72603-4|LNC|Beta hydroxybutyrate+Acetoacetate|Beta hydroxybutyrate+Acetoacetate
C3533514|T201|COMP|72602-6|LNC|Beta hydroxybutyrate+Acetoacetate^post meal|Beta hydroxybutyrate+Acetoacetate^post meal
C3533515|T201|COMP|72601-8|LNC|Beta hydroxybutyrate+Acetoacetate^pre-meal|Beta hydroxybutyrate+Acetoacetate^pre-meal
C3533516|T201|COMP|72600-0|LNC|Albumin/Protein.total|Albumin/Protein.total
C3533517|T201|COMP|72599-4|LNC|Albumin/Protein.total|Albumin/Protein.total
C3533518|T201|COMP|72598-6|LNC|Albumin/Protein.total|Albumin/Protein.total
C3533519|T201|COMP|72597-8|LNC|Albumin/Protein.total|Albumin/Protein.total
C3533520|T201|COMP|72596-0|LNC|Albumin/Protein.total|Albumin/Protein.total
C3533521|T201|COMP|72595-2|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C3533522|T201|COMP|72594-5|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C3533523|T201|COMP|72593-7|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C3533524|T201|COMP|72592-9|LNC|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C3533525|T201|COMP|72591-1|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C3533526|T201|COMP|72590-3|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C3533527|T201|COMP|72589-5|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C3533528|T201|COMP|72574-7|LNC|Coproporphyrin/Porphyrins.total|Coproporphyrin/Porphyrins.total
C3533529|T201|COMP|72573-9|LNC|Uroporphyrin/Porphyrins.total|Uroporphyrin/Porphyrins.total
C3533530|T201|COMP|72572-1|LNC|Amylase.salivary/Amylase.total|Amylase.salivary/Amylase.total
C3533531|T201|COMP|72571-3|LNC|Amylase.pancreatic/Amylase.total|Amylase.pancreatic/Amylase.total
C3533532|T201|COMP|72570-5|LNC|Cholinesterase.chloride inhibited/Cholinesterase|Cholinesterase.chloride inhibited/Cholinesterase
C3533533|T201|COMP|72569-7|LNC|Cholinesterase^dibucaine/Cholinesterase|Cholinesterase^dibucaine/Cholinesterase
C3533534|T201|COMP|72568-9|LNC|Cholinesterase.fluoride inhibited/Cholinesterase|Cholinesterase.fluoride inhibited/Cholinesterase
C3533535|T201|COMP|72567-1|LNC|Cholinesterase.RO 020683 inhibited/Cholinesterase|Cholinesterase.RO 020683 inhibited/Cholinesterase
C3533536|T201|COMP|72566-3|LNC|Cholinesterase.scoline inhibited/Cholinesterase|Cholinesterase.scoline inhibited/Cholinesterase
C3533537|T201|COMP|72565-5|LNC|Creatine kinase.BB/Creatine kinase.total|Creatine kinase.BB/Creatine kinase.total
C3533538|T201|COMP|72564-8|LNC|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C3533539|T201|COMP|72563-0|LNC|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C3533540|T201|COMP|72562-2|LNC|Creatine kinase.MM/Creatine kinase.total|Creatine kinase.MM/Creatine kinase.total
C3533542|T201|COMP|72560-6|LNC|HIV integrase inhibitor susceptibility panel|HIV integrase inhibitor susceptibility panel
C3533543|T201|COMP|72559-8|LNC|HIV integrase inhibitor susceptibility panel|HIV integrase inhibitor susceptibility panel
C3533544|T201|COMP|72558-0|LNC|Etravirine|Etravirine
C3533545|T201|COMP|72557-2|LNC|Rilpivirine|Rilpivirine
C3533575|T201|COMP|72526-7|LNC|Elvitegravir|Elvitegravir
C3533576|T201|COMP|72525-9|LNC|Raltegravir|Raltegravir
C3533577|T201|COMP|72524-2|LNC|Myelin Ab|Myelin Ab
C3533578|T201|COMP|72523-4|LNC|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C3533579|T201|COMP|72522-6|LNC|p-ANCA formalin resistant Ab.IgG|p-ANCA formalin resistant Ab.IgG
C3533580|T201|COMP|72521-8|LNC|p-ANCA formalin sensitive Ab.IgG|p-ANCA formalin sensitive Ab.IgG
C3533581|T201|COMP|72520-0|LNC|FLT3 gene.p.Asp835+Ile836|FLT3 gene.p.Asp835+Ile836
C3533583|T201|COMP|72518-4|LNC|CHEK2 gene.c.470C>T & 1100delC|CHEK2 gene.c.470C>T & 1100delC
C3533584|T201|COMP|72517-6|LNC|Spermatozoa^post ejaculate|Spermatozoa^post ejaculate
C3533585|T201|COMP|72516-8|LNC|Glucose|Glucose
C3533586|T201|COMP|72515-0|LNC|Myeloperoxidase Ab.IgG|Myeloperoxidase Ab.IgG
C3533588|T201|COMP|72511-9|LNC|CYP2B6 gene targeted mutation analysis|CYP2B6 gene targeted mutation analysis
C3533591|T201|COMP|72508-5|LNC|UGT1A1 gene.c.A(TA)7TAA(*28)|UGT1A1 gene.c.A(TA)7TAA(*28)
C3533592|T201|COMP|72507-7|LNC|VKORC1 gene.c.1173C>T|VKORC1 gene.c.1173C>T
C3533593|T201|COMP|72506-9|LNC|ABCB1 gene.c.3435C>T|ABCB1 gene.c.3435C>T
C3533594|T201|COMP|72505-1|LNC|Exserohilum rostratum DNA|Exserohilum rostratum DNA
C3533595|T201|COMP|72504-4|LNC|CV2 Ab|CV2 Ab
C3533596|T201|COMP|72503-6|LNC|WT1 gene exon 1+2 transcript/control transcript|WT1 gene exon 1+2 transcript/control transcript
C3533598|T201|COMP|72501-0|LNC|Homocyst(e)ine^6H post dose methionine|Homocyst(e)ine^6H post dose methionine
C3533599|T201|COMP|72500-2|LNC|Homocyst(e)ine^post CFst|Homocyst(e)ine^post CFst
C3533600|T201|COMP|72499-7|LNC|Oval fat bodies (globules)|Oval fat bodies (globules)
C3533601|T201|COMP|72498-9|LNC|Tripeptidyl peptidase I|Tripeptidyl peptidase I
C3533602|T201|COMP|72497-1|LNC|Dihydropteridine reductase|Dihydropteridine reductase
C3533603|T201|COMP|72496-3|LNC|DNA double strand|DNA double strand
C3533604|T201|COMP|72495-5|LNC|Candida parapsilosis DNA|Candida parapsilosis DNA
C3533605|T201|COMP|72494-8|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C3533606|T201|COMP|72493-0|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C3533607|T201|COMP|72492-2|LNC|Paraoxonase-arylesterase 1|Paraoxonase-arylesterase 1
C3533608|T201|COMP|72491-4|LNC|Bile acid|Bile acid
C3533609|T201|COMP|72490-6|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C3533610|T201|COMP|72489-8|LNC|Androstenedione|Androstenedione
C3533611|T201|COMP|72488-0|LNC|Beta 2 glycoprotein 1 Ab.IgG & IgM panel|Beta 2 glycoprotein 1 Ab.IgG & IgM panel
C3533612|T201|COMP|72487-2|LNC|TF gene full mutation analysis|TF gene full mutation analysis
C3533613|T201|COMP|72486-4|LNC|Laboratory director name|Laboratory director name
C3533614|T201|COMP|72485-6|LNC|Tapentadol|Tapentadol
C3533615|T201|COMP|72484-9|LNC|BK virus subtype|BK virus subtype
C3533616|T201|COMP|72483-1|LNC|BK virus subtype|BK virus subtype
C3533617|T201|COMP|72482-3|LNC|BK virus subtype|BK virus subtype
C3533618|T201|COMP|72481-5|LNC|Candida sp 6 panel|Candida sp 6 panel
C3533619|T201|COMP|72478-1|LNC|Synthetic cannabinoids panel|Synthetic cannabinoids panel
C3533620|T201|COMP|72475-7|LNC|Methadone+Metabolite|Methadone+Metabolite
C3533621|T201|COMP|72474-0|LNC|JWH-122 5-hydroxypentyl|JWH-122 5-hydroxypentyl
C3533622|T201|COMP|72473-2|LNC|JWH-398 5-hydroxypentyl|JWH-398 5-hydroxypentyl
C3533623|T201|COMP|72460-9|LNC|JWH-073 3-hydroxybutyl|JWH-073 3-hydroxybutyl
C3533624|T201|COMP|72459-1|LNC|JWH-018 4+5-hydroxypentyl|JWH-018 4+5-hydroxypentyl
C3533625|T201|COMP|72458-3|LNC|Myosin Ab|Myosin Ab
C3533626|T201|COMP|72456-7|LNC|Benzodiazepines|Benzodiazepines
C3533627|T201|COMP|72455-9|LNC|Amobarbital|Amobarbital
C3533628|T201|COMP|72454-2|LNC|Butalbital|Butalbital
C3533629|T201|COMP|72453-4|LNC|PHENobarbital|PHENobarbital
C3533630|T201|COMP|72452-6|LNC|Secobarbital|Secobarbital
C3533631|T201|COMP|72451-8|LNC|Barbiturates|Barbiturates
C3533632|T201|COMP|72450-0|LNC|3-Hydroxyisovalerate|3-Hydroxyisovalerate
C3533633|T201|COMP|72449-2|LNC|3-Hydroxyisovalerate|3-Hydroxyisovalerate
C3533634|T201|COMP|72448-4|LNC|3-Hydroxysebacate|3-Hydroxysebacate
C3533635|T201|COMP|72447-6|LNC|3-Hydroxysebacate|3-Hydroxysebacate
C3533636|T201|COMP|72446-8|LNC|3-Hydroxysuberate|3-Hydroxysuberate
C3533637|T201|COMP|72445-0|LNC|3-Hydroxysuberate|3-Hydroxysuberate
C3533638|T201|COMP|72444-3|LNC|3-Hydroxytetradecanedioate|3-Hydroxytetradecanedioate
C3533639|T201|COMP|72443-5|LNC|3-Methyladipate|3-Methyladipate
C3533640|T201|COMP|72442-7|LNC|3-Methylcrotonylglycine|3-Methylcrotonylglycine
C3533641|T201|COMP|72441-9|LNC|3-Methylcrotonylglycine|3-Methylcrotonylglycine
C3533642|T201|COMP|72440-1|LNC|3-Methylglutaconate|3-Methylglutaconate
C3533643|T201|COMP|72439-3|LNC|3-Methylglutarate|3-Methylglutarate
C3533644|T201|COMP|72438-5|LNC|3-Methylglutarate|3-Methylglutarate
C3533645|T201|COMP|72437-7|LNC|Phenyllactate|Phenyllactate
C3533646|T201|COMP|72436-9|LNC|Phenylpyruvate|Phenylpyruvate
C3533647|T201|COMP|72435-1|LNC|4,5-Dihydroxyhexanoate|4,5-Dihydroxyhexanoate
C3533648|T201|COMP|72434-4|LNC|4,5-Dihydroxyhexanolactone|4,5-Dihydroxyhexanolactone
C3533649|T201|COMP|72432-8|LNC|4-Hydroxyphenylacetate|4-Hydroxyphenylacetate
C3533650|T201|COMP|72431-0|LNC|4-Hydroxyphenylacetate|4-Hydroxyphenylacetate
C3533651|T201|COMP|72430-2|LNC|4-Hydroxyphenyllactate|4-Hydroxyphenyllactate
C3533652|T201|COMP|72429-4|LNC|4-Hydroxyphenyllactate|4-Hydroxyphenyllactate
C3533653|T201|COMP|72428-6|LNC|4-Hydroxyphenylpyruvate|4-Hydroxyphenylpyruvate
C3533654|T201|COMP|72427-8|LNC|4-Hydroxyphenylpyruvate|4-Hydroxyphenylpyruvate
C3533655|T201|COMP|72426-0|LNC|5-Hydroxyhexanoate|5-Hydroxyhexanoate
C3533656|T201|COMP|72425-2|LNC|7-Hydroxyoctanoate|7-Hydroxyoctanoate
C3533657|T201|COMP|72424-5|LNC|3-Methylhistidine/Amino acids.total|3-Methylhistidine/Amino acids.total
C3533658|T201|COMP|72423-7|LNC|3-Methylhistidine|3-Methylhistidine
C3533659|T201|COMP|72422-9|LNC|Gamma aminobutyrate|Gamma aminobutyrate
C3533660|T201|COMP|72421-1|LNC|Bacterial vancomycin resistance vanB gene|Bacterial vancomycin resistance vanB gene
C3533661|T201|COMP|72420-3|LNC|Gamma aminobutyrate.free|Gamma aminobutyrate.free
C3533662|T201|COMP|72419-5|LNC|Beta hydroxybutyrate/Acetoacetate^post meal|Beta hydroxybutyrate/Acetoacetate^post meal
C3533663|T201|COMP|72418-7|LNC|Beta hydroxybutyrate/Acetoacetate^pre-meal|Beta hydroxybutyrate/Acetoacetate^pre-meal
C3533664|T201|COMP|72417-9|LNC|Beta hydroxybutyrate^pre-meal|Beta hydroxybutyrate^pre-meal
C3533665|T201|COMP|72416-1|LNC|Beta hydroxybutyrate^post meal|Beta hydroxybutyrate^post meal
C3533666|T201|COMP|72415-3|LNC|Acetoacetate^post meal|Acetoacetate^post meal
C3533667|T201|COMP|72414-6|LNC|Acetoacetate^pre-meal|Acetoacetate^pre-meal
C3533668|T201|COMP|72413-8|LNC|BK virus subtype|BK virus subtype
C3533669|T201|COMP|72412-0|LNC|BK virus subtype|BK virus subtype
C3533670|T201|COMP|72411-2|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C3533671|T201|COMP|72410-4|LNC|Testosterone^pre dose HCG|Testosterone^pre dose HCG
C3533672|T201|COMP|72409-6|LNC|Testosterone^post dose HCG|Testosterone^post dose HCG
C3533674|T201|COMP|72407-0|LNC|Benzoylecgonine|Benzoylecgonine
C3533675|T201|COMP|72406-2|LNC|Norchlordiazepoxide|Norchlordiazepoxide
C3533676|T201|COMP|72405-4|LNC|Cocaine|Cocaine
C3533677|T201|COMP|72404-7|LNC|3-epi-25-Hydroxyvitamin D2|3-epi-25-Hydroxyvitamin D2
C3533678|T201|COMP|72403-9|LNC|3-epi-25-Hydroxyvitamin D3|3-epi-25-Hydroxyvitamin D3
C3533679|T201|COMP|72402-1|LNC|oxyCODONE|oxyCODONE
C3533680|T201|COMP|72401-3|LNC|Propoxyphene|Propoxyphene
C3533681|T201|COMP|72400-5|LNC|Methadone|Methadone
C3533682|T201|COMP|72399-9|LNC|Amobarbital|Amobarbital
C3533683|T201|COMP|72398-1|LNC|Butalbital|Butalbital
C3533684|T201|COMP|72397-3|LNC|Secobarbital|Secobarbital
C3533685|T201|COMP|72396-5|LNC|PHENobarbital|PHENobarbital
C3533686|T201|COMP|72395-7|LNC|Differential panel|Differential panel
C3533687|T201|COMP|72394-0|LNC|Cell count panel|Cell count panel
C3533688|T201|COMP|72393-2|LNC|Cell count & Differential panel|Cell count & Differential panel
C3533689|T201|COMP|72392-4|LNC|Cortisol/Cortisone|Cortisol/Cortisone
C3533690|T201|COMP|72391-6|LNC|Candida tropicalis DNA|Candida tropicalis DNA
C3533691|T201|COMP|72390-8|LNC|Candida lusitaniae DNA|Candida lusitaniae DNA
C3533692|T201|COMP|72389-0|LNC|Candida krusei DNA|Candida krusei DNA
C3533693|T201|COMP|72376-7|LNC|Hepatitis C virus Ab|Hepatitis C virus Ab
C3533694|T201|COMP|72375-9|LNC|Microscopic method|Microscopic method
C3533695|T201|COMP|72374-2|LNC|Virus identified|Virus identified
C3533696|T201|COMP|72373-4|LNC|Virus identified|Virus identified
C3533700|T201|COMP|72368-4|LNC|t(11;14)(q13;q32)(CCND1,IGH) fusion transcript|t(11;14)(q13;q32)(CCND1,IGH) fusion transcript
C3533701|T201|COMP|72367-6|LNC|Influenza virus A+B Ag|Influenza virus A+B Ag
C3533702|T201|COMP|72366-8|LNC|Influenza virus A & B Ag|Influenza virus A & B Ag
C3533703|T201|COMP|72365-0|LNC|Influenza virus A & B Ag|Influenza virus A & B Ag
C3533704|T201|COMP|72364-3|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C3533705|T201|COMP|72362-7|LNC|Starch granules|Starch granules
C3533706|T201|COMP|72361-9|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C3533707|T201|COMP|72360-1|LNC|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C3533709|T201|COMP|72356-9|LNC|Influenza virus A & B Ag|Influenza virus A & B Ag
C3533715|T201|COMP|72348-6|LNC|Leukocytes|Leukocytes
C3533716|T201|COMP|72347-8|LNC|Neutrophils|Neutrophils
C3533717|T201|COMP|72346-0|LNC|Round cells|Round cells
C3533718|T201|COMP|72345-2|LNC|Neutrophils/100 round cells|Neutrophils/100 round cells
C3533719|T201|COMP|72344-5|LNC|Monocytes/100 round cells|Monocytes/100 round cells
C3533720|T201|COMP|72343-7|LNC|Monocytes/100 round cells|Monocytes/100 round cells
C3533721|T201|COMP|72342-9|LNC|Neutrophils/100 round cells|Neutrophils/100 round cells
C3533722|T201|COMP|72341-1|LNC|Amyloid bodies|Amyloid bodies
C3533723|T201|COMP|72340-3|LNC|Bacteria|Bacteria
C3533724|T201|COMP|72339-5|LNC|Lecithin|Lecithin
C3533725|T201|COMP|72338-7|LNC|Erythrocytes|Erythrocytes
C3533726|T201|COMP|72337-9|LNC|Protein S Ag|Protein S Ag
C3533730|T201|COMP|72333-8|LNC|JAK2 gene.p.Val617Phe|JAK2 gene.p.Val617Phe
C3533731|T201|COMP|72332-0|LNC|Nucleated cells/100 round cells|Nucleated cells/100 round cells
C3533732|T201|COMP|72331-2|LNC|Anucleated bodies/100 round cells|Anucleated bodies/100 round cells
C3533733|T201|COMP|72330-4|LNC|Nucleated cells/100 round cells|Nucleated cells/100 round cells
C3533734|T201|COMP|72329-6|LNC|Anucleated bodies/100 round cells|Anucleated bodies/100 round cells
C3533735|T201|COMP|72328-8|LNC|HLA-A+B+C Ab.IgG|HLA-A+B+C Ab.IgG
C3533736|T201|COMP|72327-0|LNC|Amphiphysin Ab.IgG|Amphiphysin Ab.IgG
C3533740|T201|COMP|72323-9|LNC|HLA-DP+DQ+DR Ab.IgG|HLA-DP+DQ+DR Ab.IgG
C3533741|T201|COMP|72322-1|LNC|HLA-A+B+C Ab.IgG|HLA-A+B+C Ab.IgG
C3533742|T201|COMP|72321-3|LNC|HLA-DP+DQ+DR Ab.IgG|HLA-DP+DQ+DR Ab.IgG
C3533743|T201|COMP|72320-5|LNC|Mitochondria M2-3E Ab.IgG|Mitochondria M2-3E Ab.IgG
C3533744|T201|COMP|72318-9|LNC|Centromere protein A Ab.IgG|Centromere protein A Ab.IgG
C3533745|T201|COMP|72317-1|LNC|RNA polymerase III RP11 Ab.IgG|RNA polymerase III RP11 Ab.IgG
C3533746|T201|COMP|72316-3|LNC|RNA polymerase III RP155 Ab.IgG|RNA polymerase III RP155 Ab.IgG
C3533747|T201|COMP|72315-5|LNC|Platelet-derived growth factor receptor Ab.IgG|Platelet-derived growth factor receptor Ab.IgG
C3533748|T201|COMP|72314-8|LNC|Th-To Ab.IgG|Th-To Ab.IgG
C3533754|T201|COMP|72308-0|LNC|Brucella sp Ab.IgG^1st specimen|Brucella sp Ab.IgG^1st specimen
C3533755|T201|COMP|72307-2|LNC|Brucella sp Ab.IgG^2nd specimen|Brucella sp Ab.IgG^2nd specimen
C3533756|T201|COMP|72306-4|LNC|Nicotinurate|Nicotinurate
C3533773|T201|COMP|72280-1|LNC|Rh immune globulin expiration|Rh immune globulin expiration
C3533775|T201|COMP|72278-5|LNC|Specimen volume|Specimen volume
C3533776|T201|COMP|72277-7|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C3533780|T201|COMP|72273-6|LNC|Blood product ordered|Blood product ordered
C3533781|T201|COMP|72272-8|LNC|Amylase & triacylglycerol lipase panel|Amylase & triacylglycerol lipase panel
C3533782|T201|COMP|72271-0|LNC|Creatinine^pre contrast|Creatinine^pre contrast
C3533783|T201|COMP|72270-2|LNC|Urea nitrogen^pre contrast|Urea nitrogen^pre contrast
C3533784|T201|COMP|72262-9|LNC|Methemoglobin|Methemoglobin
C3533785|T201|COMP|72261-1|LNC|Bilirubin excess|Bilirubin excess
C3533786|T201|COMP|72260-3|LNC|Tau protein.phosphorylated 181|Tau protein.phosphorylated 181
C3533787|T201|COMP|72259-5|LNC|Adefovir|Adefovir
C3533788|T201|COMP|72258-7|LNC|Malondialdehyde|Malondialdehyde
C3533809|T201|COMP|72224-9|LNC|Pathologic casts|Pathologic casts
C3533810|T201|COMP|72223-1|LNC|Yeast|Yeast
C3533819|T201|COMP|72206-6|LNC|Epstein Barr virus nuclear 1 Ab.IgG & IgM|Epstein Barr virus nuclear 1 Ab.IgG & IgM
C3533822|T201|COMP|72203-3|LNC|Parathyrin.intact intraoperative panel|Parathyrin.intact intraoperative panel
C3533848|T201|COMP|72174-6|LNC|Rotavirus Ag|Rotavirus Ag
C3533851|T201|COMP|72171-2|LNC|Glucose tolerance 2H panel|Glucose tolerance 2H panel
C3533853|T201|COMP|72168-8|LNC|Ofloxacin 1.5 ug/mL|Ofloxacin 1.5 ug/mL
C3533856|T201|COMP|72163-9|LNC|Leukocytes|Leukocytes
C3533857|T201|COMP|72162-1|LNC|Erythrocytes|Erythrocytes
C3533858|T201|COMP|72161-3|LNC|Epithelial cells|Epithelial cells
C3533859|T201|COMP|72160-5|LNC|Holo-transcobalamin II|Holo-transcobalamin II
C3533860|T201|COMP|72159-7|LNC|Inulin renal clearance/1.73 sq M|Inulin renal clearance/1.73 sq M
C3533861|T201|COMP|72158-9|LNC|Apo-transcobalamin I|Apo-transcobalamin I
C3533862|T201|COMP|72157-1|LNC|Apo-transcobalamin II|Apo-transcobalamin II
C3533874|T201|COMP|72827-9|LNC|dic(9;20)(p11-13;q11)(wcp9+,wcp20+)|dic(9;20)(p11-13;q11)(wcp9+,wcp20+)
C3533876|T201|COMP|72825-3|LNC|Phencyclidine|Phencyclidine
C3533877|T201|COMP|72588-7|LNC|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C3533878|T201|COMP|72587-9|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C3533879|T201|COMP|72586-1|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C3533880|T201|COMP|72585-3|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C3533881|T201|COMP|72584-6|LNC|Beta globulin/Protein.total|Beta globulin/Protein.total
C3533882|T201|COMP|72583-8|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C3533883|T201|COMP|72582-0|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C3533884|T201|COMP|72581-2|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C3533885|T201|COMP|72580-4|LNC|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C3533886|T201|COMP|72579-6|LNC|Prealbumin/Protein.total|Prealbumin/Protein.total
C3533887|T201|COMP|72578-8|LNC|Prealbumin/Protein.total|Prealbumin/Protein.total
C3533888|T201|COMP|72577-0|LNC|Protein.monoclonal/Protein.total|Protein.monoclonal/Protein.total
C3533890|T201|COMP|72575-4|LNC|Macroprolactin/Prolactin|Macroprolactin/Prolactin
C3533892|T201|COMP|72268-6|LNC|Streptococcus pyogenes exotoxin B speB gene|Streptococcus pyogenes exotoxin B speB gene
C3533894|T201|COMP|72266-0|LNC|Influenza virus A Ab.IgA|Influenza virus A Ab.IgA
C3533895|T201|COMP|72265-2|LNC|Influenza virus B Ab.IgA|Influenza virus B Ab.IgA
C3533897|T201|COMP|72263-7|LNC|Oxyhemoglobin|Oxyhemoglobin
C3533911|T201|COMP|72777-6|LNC|JWH-018 butanol/Creatinine|JWH-018 butanol/Creatinine
C3533912|T201|COMP|72776-8|LNC|JWH-018 butanol|JWH-018 butanol
C3533913|T201|COMP|72775-0|LNC|Venlafaxine/Creatinine|Venlafaxine/Creatinine
C3533914|T201|COMP|72774-3|LNC|Venlafaxine|Venlafaxine
C3533915|T201|COMP|72773-5|LNC|Norvenlafaxine/Creatinine|Norvenlafaxine/Creatinine
C3533916|T201|COMP|72772-7|LNC|Norvenlafaxine|Norvenlafaxine
C3533917|T201|COMP|72771-9|LNC|Zolpidem/Creatinine|Zolpidem/Creatinine
C3533918|T201|COMP|72770-1|LNC|Zolpidem|Zolpidem
C3533919|T201|COMP|72769-3|LNC|Zolpidem phenyl-4-carboxylate/Creatinine|Zolpidem phenyl-4-carboxylate/Creatinine
C3533920|T201|COMP|72768-5|LNC|Zolpidem phenyl-4-carboxylate|Zolpidem phenyl-4-carboxylate
C3533921|T201|COMP|72766-9|LNC|oxyMORphone|oxyMORphone
C3533922|T201|COMP|72765-1|LNC|Phencyclidine|Phencyclidine
C3533923|T201|COMP|72764-4|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C3533924|T201|COMP|72763-6|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C3533925|T201|COMP|72762-8|LNC|Buprenorphine|Buprenorphine
C3533926|T201|COMP|72761-0|LNC|Carisoprodol|Carisoprodol
C3533927|T201|COMP|72760-2|LNC|fentaNYL|fentaNYL
C3533928|T201|COMP|72759-4|LNC|Codeine|Codeine
C3533929|T201|COMP|72758-6|LNC|Amphetamine|Amphetamine
C3533930|T201|COMP|72388-2|LNC|Methadone|Methadone
C3533931|T201|COMP|72387-4|LNC|Methadone|Methadone
C3533932|T201|COMP|72386-6|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C3533933|T201|COMP|72385-8|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C3533934|T201|COMP|72384-1|LNC|Meperidine+Normeperidine|Meperidine+Normeperidine
C3533935|T201|COMP|72383-3|LNC|HER2|HER2
C3533936|T201|COMP|72382-5|LNC|HER2|HER2
C3533937|T201|COMP|72381-7|LNC|ALPRAZolam|ALPRAZolam
C3533938|T201|COMP|72380-9|LNC|LORazepam|LORazepam
C3533939|T201|COMP|72379-1|LNC|Cannabinoids.synthetic|Cannabinoids.synthetic
C3533940|T201|COMP|72378-3|LNC|Oxazepam|Oxazepam
C3533941|T201|COMP|72377-5|LNC|Nordiazepam|Nordiazepam
C3533943|T201|COMP|72466-6|LNC|JWH-250 5-hydroxypentyl|JWH-250 5-hydroxypentyl
C3533944|T201|COMP|72465-8|LNC|JWH-073 butanoate|JWH-073 butanoate
C3533945|T201|COMP|72464-1|LNC|JWH-073 4-hydroxybutyl|JWH-073 4-hydroxybutyl
C3533946|T201|COMP|72463-3|LNC|AM-2201 4-hydroxypentyl|AM-2201 4-hydroxypentyl
C3533947|T201|COMP|72462-5|LNC|JWH-200 4-Hydroxyindole|JWH-200 4-Hydroxyindole
C3533948|T201|COMP|72461-7|LNC|JWH-018 pentanoate|JWH-018 pentanoate
C3533949|T201|COMP|72220-7|LNC|Macrophages|Macrophages
C3533950|T201|COMP|72219-9|LNC|Lymphocytes|Lymphocytes
C3533955|T201|COMP|71680-3|LNC|Basophils/leukocytes|Basophils/leukocytes
C3533956|T201|COMP|71679-5|LNC|Eosinophils/leukocytes|Eosinophils/leukocytes
C3533957|T201|COMP|71678-7|LNC|Lymphocytes/leukocytes|Lymphocytes/leukocytes
C3533958|T201|COMP|71677-9|LNC|Monocytes/leukocytes|Monocytes/leukocytes
C3533959|T201|COMP|71676-1|LNC|Neutrophils/leukocytes|Neutrophils/leukocytes
C3533960|T201|COMP|71675-3|LNC|Basophils/leukocytes|Basophils/leukocytes
C3533961|T201|COMP|71674-6|LNC|Eosinophils/leukocytes|Eosinophils/leukocytes
C3533962|T201|COMP|71673-8|LNC|Lymphocytes/leukocytes|Lymphocytes/leukocytes
C3533963|T201|COMP|71672-0|LNC|Monocytes/leukocytes|Monocytes/leukocytes
C3533964|T201|COMP|71671-2|LNC|Neutrophils/leukocytes|Neutrophils/leukocytes
C3533965|T201|COMP|71670-4|LNC|Neutrophils.band form/leukocytes|Neutrophils.band form/leukocytes
C3533966|T201|COMP|71669-6|LNC|Blasts/leukocytes|Blasts/leukocytes
C3533967|T201|COMP|71668-8|LNC|Metamyelocytes/leukocytes|Metamyelocytes/leukocytes
C3533968|T201|COMP|71667-0|LNC|Myelocytes/leukocytes|Myelocytes/leukocytes
C3533969|T201|COMP|71666-2|LNC|Promyelocytes/leukocytes|Promyelocytes/leukocytes
C3533970|T201|COMP|71665-4|LNC|Lymphocytes.variant/leukocytes|Lymphocytes.variant/leukocytes
C3533971|T201|COMP|71664-7|LNC|Smudge cells/leukocytes|Smudge cells/leukocytes
C3533972|T201|COMP|71663-9|LNC|Plasma cells/leukocytes|Plasma cells/leukocytes
C3533973|T201|COMP|71662-1|LNC|Basophils/leukocytes|Basophils/leukocytes
C3533974|T201|COMP|71661-3|LNC|Eosinophils/leukocytes|Eosinophils/leukocytes
C3533975|T201|COMP|71660-5|LNC|Lymphocytes/leukocytes|Lymphocytes/leukocytes
C3533976|T201|COMP|71659-7|LNC|Monocytes/leukocytes|Monocytes/leukocytes
C3533977|T201|COMP|71658-9|LNC|Neutrophils/leukocytes|Neutrophils/leukocytes
C3533978|T201|COMP|71657-1|LNC|Neutrophils.band form/leukocytes|Neutrophils.band form/leukocytes
C3533979|T201|COMP|71656-3|LNC|Blasts/leukocytes|Blasts/leukocytes
C3533980|T201|COMP|71655-5|LNC|Metamyelocytes/leukocytes|Metamyelocytes/leukocytes
C3533981|T201|COMP|71654-8|LNC|Myelocytes/leukocytes|Myelocytes/leukocytes
C3533982|T201|COMP|71653-0|LNC|Promyelocytes/leukocytes|Promyelocytes/leukocytes
C3533983|T201|COMP|71652-2|LNC|Plasma cells/leukocytes|Plasma cells/leukocytes
C3533984|T201|COMP|71651-4|LNC|Macrophages/leukocytes|Macrophages/leukocytes
C3533985|T201|COMP|71650-6|LNC|Neutrophils.segmented/leukocytes|Neutrophils.segmented/leukocytes
C3533986|T201|COMP|71649-8|LNC|Lymphocytes/leukocytes|Lymphocytes/leukocytes
C3533987|T201|COMP|71648-0|LNC|Monocytes/leukocytes|Monocytes/leukocytes
C3533988|T201|COMP|71647-2|LNC|Basophils/leukocytes|Basophils/leukocytes
C3533989|T201|COMP|71646-4|LNC|Eosinophils/leukocytes|Eosinophils/leukocytes
C3533990|T201|COMP|71645-6|LNC|Neutrophils.band form/leukocytes|Neutrophils.band form/leukocytes
C3533991|T201|COMP|71644-9|LNC|Blasts/leukocytes|Blasts/leukocytes
C3533992|T201|COMP|71643-1|LNC|Metamyelocytes/leukocytes|Metamyelocytes/leukocytes
C3533993|T201|COMP|71642-3|LNC|Promyelocytes/leukocytes|Promyelocytes/leukocytes
C3533994|T201|COMP|71641-5|LNC|Macrophages/leukocytes|Macrophages/leukocytes
C3533995|T201|COMP|71640-7|LNC|Mesothelial cells/leukocytes|Mesothelial cells/leukocytes
C3533996|T201|COMP|71639-9|LNC|Monocytes+Macrophages/leukocytes|Monocytes+Macrophages/leukocytes
C3533997|T201|COMP|71638-1|LNC|Unidentified cells/leukocytes|Unidentified cells/leukocytes
C3533998|T201|COMP|71637-3|LNC|Unspecified cells/leukocytes|Unspecified cells/leukocytes
C3533999|T201|COMP|71636-5|LNC|Plasma cells/leukocytes|Plasma cells/leukocytes
C3534000|T201|COMP|71635-7|LNC|Neutrophils/leukocytes|Neutrophils/leukocytes
C3534001|T201|COMP|71634-0|LNC|Lymphocytes/leukocytes|Lymphocytes/leukocytes
C3534002|T201|COMP|71633-2|LNC|Monocytes/leukocytes|Monocytes/leukocytes
C3534003|T201|COMP|71632-4|LNC|Eosinophils/leukocytes|Eosinophils/leukocytes
C3534004|T201|COMP|71631-6|LNC|Basophils/leukocytes|Basophils/leukocytes
C3534005|T201|COMP|71630-8|LNC|Leukocytes other/leukocytes|Leukocytes other/leukocytes
C3534006|T201|COMP|71629-0|LNC|Mononuclear cells/leukocytes|Mononuclear cells/leukocytes
C3534007|T201|COMP|71628-2|LNC|Macrophages/leukocytes|Macrophages/leukocytes
C3534008|T201|COMP|71627-4|LNC|Polymorphonuclear cells/leukocytes|Polymorphonuclear cells/leukocytes
C3534009|T201|COMP|71626-6|LNC|Mesothelial cells/leukocytes|Mesothelial cells/leukocytes
C3534010|T201|COMP|71625-8|LNC|Neutrophils/leukocytes|Neutrophils/leukocytes
C3534011|T201|COMP|71624-1|LNC|Lymphocytes/leukocytes|Lymphocytes/leukocytes
C3534012|T201|COMP|71623-3|LNC|Monocytes/leukocytes|Monocytes/leukocytes
C3534013|T201|COMP|71622-5|LNC|Eosinophils/leukocytes|Eosinophils/leukocytes
C3534014|T201|COMP|71621-7|LNC|Basophils/leukocytes|Basophils/leukocytes
C3534015|T201|COMP|71613-4|LNC|Eosinophils/leukocytes|Eosinophils/leukocytes
C3534016|T201|COMP|71612-6|LNC|Basophils/leukocytes|Basophils/leukocytes
C3534017|T201|COMP|71611-8|LNC|Leukocytes other/leukocytes|Leukocytes other/leukocytes
C3534018|T201|COMP|71610-0|LNC|Mononuclear cells/leukocytes|Mononuclear cells/leukocytes
C3534019|T201|COMP|71609-2|LNC|Macrophages/leukocytes|Macrophages/leukocytes
C3534020|T201|COMP|71608-4|LNC|Polymorphonuclear cells/leukocytes|Polymorphonuclear cells/leukocytes
C3534021|T201|COMP|71607-6|LNC|Mesothelial cells/leukocytes|Mesothelial cells/leukocytes
C3534022|T201|COMP|71606-8|LNC|Neutrophils/leukocytes|Neutrophils/leukocytes
C3534023|T201|COMP|71605-0|LNC|Lymphocytes/leukocytes|Lymphocytes/leukocytes
C3534024|T201|COMP|71604-3|LNC|Monocytes/leukocytes|Monocytes/leukocytes
C3534025|T201|COMP|71603-5|LNC|Eosinophils/leukocytes|Eosinophils/leukocytes
C3534026|T201|COMP|71602-7|LNC|Basophils/leukocytes|Basophils/leukocytes
C3534027|T201|COMP|71601-9|LNC|Leukocytes other/leukocytes|Leukocytes other/leukocytes
C3534028|T201|COMP|71600-1|LNC|Macrophages/leukocytes|Macrophages/leukocytes
C3534029|T201|COMP|71599-5|LNC|Mesothelial cells/leukocytes|Mesothelial cells/leukocytes
C3534030|T201|COMP|71598-7|LNC|Neutrophils/leukocytes|Neutrophils/leukocytes
C3534031|T201|COMP|71597-9|LNC|Lymphocytes/leukocytes|Lymphocytes/leukocytes
C3534032|T201|COMP|71596-1|LNC|Eosinophils/leukocytes|Eosinophils/leukocytes
C3534033|T201|COMP|71595-3|LNC|Basophils/leukocytes|Basophils/leukocytes
C3534034|T201|COMP|71594-6|LNC|Macrophages/leukocytes|Macrophages/leukocytes
C3534036|T201|COMP|72680-2|LNC|Macroprolactin|Macroprolactin
C3534037|T201|COMP|72655-4|LNC|Aldolase|Aldolase
C3534038|T201|COMP|72654-7|LNC|SNRPN gene 15q11 deletion+duplication|SNRPN gene 15q11 deletion+duplication
C3534039|T201|COMP|72653-9|LNC|Subtelomere analysis.short arm|Subtelomere analysis.short arm
C3534040|T201|COMP|72652-1|LNC|Subtelomere analysis.long arm|Subtelomere analysis.long arm
C3534041|T201|COMP|72651-3|LNC|Glucose.serum-glucose.plr fld|Glucose.serum-glucose.plr fld
C3534042|T201|COMP|72650-5|LNC|Glucose.serum-glucose.pericard fld|Glucose.serum-glucose.pericard fld
C3534043|T201|COMP|72472-4|LNC|UR-144 pentanoate|UR-144 pentanoate
C3534044|T201|COMP|72471-6|LNC|UR-144 4+5-hydroxypentyl|UR-144 4+5-hydroxypentyl
C3534045|T201|COMP|72470-8|LNC|MAM-2201 pentanoate|MAM-2201 pentanoate
C3534046|T201|COMP|72469-0|LNC|RCS-4 5-carboxypentyl|RCS-4 5-carboxypentyl
C3534047|T201|COMP|72468-2|LNC|RCS-4 5-hydroxypentyl|RCS-4 5-hydroxypentyl
C3534048|T201|COMP|72467-4|LNC|JWH-250 5-carboxypentyl|JWH-250 5-carboxypentyl
C3534049|T201|COMP|71620-9|LNC|Leukocytes other/leukocytes|Leukocytes other/leukocytes
C3534050|T201|COMP|71619-1|LNC|Mononuclear cells/leukocytes|Mononuclear cells/leukocytes
C3534051|T201|COMP|71618-3|LNC|Macrophages/leukocytes|Macrophages/leukocytes
C3534052|T201|COMP|71617-5|LNC|Polymorphonuclear cells/leukocytes|Polymorphonuclear cells/leukocytes
C3534053|T201|COMP|71616-7|LNC|Neutrophils/leukocytes|Neutrophils/leukocytes
C3534054|T201|COMP|71615-9|LNC|Lymphocytes/leukocytes|Lymphocytes/leukocytes
C3534055|T201|COMP|71614-2|LNC|Monocytes/leukocytes|Monocytes/leukocytes
C3534057|T201|COMP|58469-8|LNC|Cells|Cells
C3534060|T201|COMP|51752-4|LNC|Heptaporphyrin/Creatinine|Heptaporphyrin/Creatinine
C3539901|T201|COMP|73913-6|LNC|Glycine CSF/Glycine plas|Glycine CSF/Glycine plas
C3539903|T201|COMP|73901-1|LNC|Cells.CD3-CD8-CD57+/100 lymphocytes|Cells.CD3-CD8-CD57+/100 lymphocytes
C3539904|T201|COMP|73900-3|LNC|Cells.CD3-CD8-CD57+/100 leukocytes|Cells.CD3-CD8-CD57+/100 leukocytes
C3541304|T201|COMP|73904-5|LNC|Cells.CD3-CD57+/100 lymphocytes|Cells.CD3-CD57+/100 lymphocytes
C3541305|T201|COMP|73903-7|LNC|Cells.CD3-CD57+/100 leukocytes|Cells.CD3-CD57+/100 leukocytes
C3541866|T201|COMP|72922-8|LNC|HNA 1a-1a Ab|HNA 1a-1a Ab
C3654067|T201|COMP|73610-8|LNC|Sarafloxacin|Sarafloxacin
C3654068|T201|COMP|73586-0|LNC|Tedizolid|Tedizolid
C3654069|T201|COMP|73582-9|LNC|Anion gap 4|Anion gap 4
C3654070|T201|COMP|72907-9|LNC|HNA genotype panel|HNA genotype panel
C3654071|T201|COMP|72899-8|LNC|Isoleucine+Leucine|Isoleucine+Leucine
C3654072|T201|COMP|73914-4|LNC|JWH-018|JWH-018
C3654073|T201|COMP|73887-2|LNC|Tetrahydrocorticosterone|Tetrahydrocorticosterone
C3654074|T201|COMP|73880-7|LNC|Cortisone.free|Cortisone.free
C3654075|T201|COMP|73862-5|LNC|Allo-tetrahydrocortisol|Allo-tetrahydrocortisol
C3654076|T201|COMP|72480-7|LNC|Barbiturates panel|Barbiturates panel
C3654077|T201|COMP|73687-6|LNC|Methylenedioxypyrovalerone|Methylenedioxypyrovalerone
C3654078|T201|COMP|73979-7|LNC|Keyhole limpet hemocyanin Ab panel|Keyhole limpet hemocyanin Ab panel
C3654079|T201|COMP|73978-9|LNC|von Willebrand factor.activity|von Willebrand factor.activity
C3654080|T201|COMP|73972-2|LNC|Morphine.free|Morphine.free
C3654082|T201|COMP|73970-6|LNC|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3654083|T201|COMP|73969-8|LNC|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3654084|T201|COMP|73968-0|LNC|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3654086|T201|COMP|73962-3|LNC|Candida sp rRNA|Candida sp rRNA
C3654088|T201|COMP|73960-7|LNC|Bacteria identified|Bacteria identified
C3654090|T201|COMP|73954-0|LNC|JWH-398 5-hydroxypentyl|JWH-398 5-hydroxypentyl
C3654091|T201|COMP|73953-2|LNC|JWH-073|JWH-073
C3654092|T201|COMP|73952-4|LNC|AM-2201|AM-2201
C3654093|T201|COMP|73951-6|LNC|RCS-4|RCS-4
C3654094|T201|COMP|73950-8|LNC|JWH-250|JWH-250
C3654095|T201|COMP|73949-0|LNC|JWH-018|JWH-018
C3654096|T201|COMP|73948-2|LNC|JWH-122|JWH-122
C3654097|T201|COMP|73947-4|LNC|JWH-398|JWH-398
C3654098|T201|COMP|73946-6|LNC|JWH-200|JWH-200
C3654099|T201|COMP|73945-8|LNC|UR-144|UR-144
C3654100|T201|COMP|73944-1|LNC|MAM-2201|MAM-2201
C3654101|T201|COMP|73943-3|LNC|Cannabinoids.synthetic|Cannabinoids.synthetic
C3654102|T201|COMP|73942-5|LNC|Buprenorphine|Buprenorphine
C3654103|T201|COMP|73941-7|LNC|6-Monoacetylmorphine.free|6-Monoacetylmorphine.free
C3654104|T201|COMP|73940-9|LNC|HYDROmorphone.free|HYDROmorphone.free
C3654105|T201|COMP|73939-1|LNC|HYDROcodone.free|HYDROcodone.free
C3654106|T201|COMP|73938-3|LNC|fentaNYL|fentaNYL
C3654107|T201|COMP|73937-5|LNC|Norfentanyl|Norfentanyl
C3654108|T201|COMP|73936-7|LNC|fentaNYL|fentaNYL
C3654109|T201|COMP|73935-9|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C3654110|T201|COMP|73934-2|LNC|Meperidine|Meperidine
C3654111|T201|COMP|73933-4|LNC|Normeperidine|Normeperidine
C3654112|T201|COMP|73932-6|LNC|traMADol|traMADol
C3654113|T201|COMP|73931-8|LNC|Propanol|Propanol
C3654114|T201|COMP|73930-0|LNC|RCS-4 5-carboxypentyl|RCS-4 5-carboxypentyl
C3654115|T201|COMP|73929-2|LNC|JWH-250 5-carboxypentyl|JWH-250 5-carboxypentyl
C3654116|T201|COMP|73928-4|LNC|JWH-250 5-hydroxypentyl|JWH-250 5-hydroxypentyl
C3654117|T201|COMP|73927-6|LNC|JWH-073 butanoate|JWH-073 butanoate
C3654118|T201|COMP|73926-8|LNC|JWH-073 4-hydroxybutyl|JWH-073 4-hydroxybutyl
C3654119|T201|COMP|73925-0|LNC|AM-2201 4-hydroxypentyl|AM-2201 4-hydroxypentyl
C3654120|T201|COMP|73924-3|LNC|JWH-200 4-Hydroxyindole|JWH-200 4-Hydroxyindole
C3654121|T201|COMP|73923-5|LNC|JWH-018 pentanoate|JWH-018 pentanoate
C3654122|T201|COMP|73922-7|LNC|RCS-4 5-hydroxypentyl|RCS-4 5-hydroxypentyl
C3654123|T201|COMP|73921-9|LNC|JWH-073 3-hydroxybutyl|JWH-073 3-hydroxybutyl
C3654124|T201|COMP|73920-1|LNC|JWH-018 4+5-hydroxypentyl|JWH-018 4+5-hydroxypentyl
C3654125|T201|COMP|73919-3|LNC|MAM-2201 pentanoate|MAM-2201 pentanoate
C3654126|T201|COMP|73918-5|LNC|JWH-073|JWH-073
C3654127|T201|COMP|73917-7|LNC|JWH-250 4+5-hydroxypentyl|JWH-250 4+5-hydroxypentyl
C3654128|T201|COMP|73916-9|LNC|1,3-Dimethylamylamine|1,3-Dimethylamylamine
C3654129|T201|COMP|73915-1|LNC|1,3-Dimethylamylamine|1,3-Dimethylamylamine
C3654130|T201|COMP|73912-8|LNC|DOG1 Ag|DOG1 Ag
C3654131|T201|COMP|73911-0|LNC|SOX10 Ag|SOX10 Ag
C3654132|T201|COMP|73910-2|LNC|PAX8 Ag|PAX8 Ag
C3654133|T201|COMP|73909-4|LNC|D2-40 Ag|D2-40 Ag
C3654134|T201|COMP|73908-6|LNC|Alloisoleucine/Creatinine|Alloisoleucine/Creatinine
C3654135|T201|COMP|73907-8|LNC|Polio virus identified|Polio virus identified
C3654136|T201|COMP|73906-0|LNC|HIV 1+2 Ab.IgG|HIV 1+2 Ab.IgG
C3654137|T201|COMP|73905-2|LNC|HIV 1+2 Ab.IgG|HIV 1+2 Ab.IgG
C3654138|T201|COMP|73902-9|LNC|Cells.CD3-CD57+|Cells.CD3-CD57+
C3654139|T201|COMP|73899-7|LNC|Cells.CD3-CD8-CD57+|Cells.CD3-CD8-CD57+
C3654140|T201|COMP|73898-9|LNC|Cells.CD8-CD57+/100 lymphocytes|Cells.CD8-CD57+/100 lymphocytes
C3654141|T201|COMP|73897-1|LNC|Chronic lyme disease panel|Chronic lyme disease panel
C3654142|T201|COMP|73895-5|LNC|Hemoglobin|Hemoglobin
C3654143|T201|COMP|73894-8|LNC|Tetrahydrocortisone|Tetrahydrocortisone
C3654144|T201|COMP|73893-0|LNC|Tetrahydrocortisone|Tetrahydrocortisone
C3654145|T201|COMP|73892-2|LNC|Tetrahydrocortisol|Tetrahydrocortisol
C3654146|T201|COMP|73891-4|LNC|Tetrahydrocortisol|Tetrahydrocortisol
C3654147|T201|COMP|73890-6|LNC|Tetrahydrocortisol|Tetrahydrocortisol
C3654148|T201|COMP|73889-8|LNC|Tetrahydrocorticosterone|Tetrahydrocorticosterone
C3654149|T201|COMP|73888-0|LNC|Tetrahydrocorticosterone|Tetrahydrocorticosterone
C3654150|T201|COMP|73886-4|LNC|Steroid fractions panel|Steroid fractions panel
C3654151|T201|COMP|73885-6|LNC|Steroid fractions panel|Steroid fractions panel
C3654152|T201|COMP|73884-9|LNC|Steroid fractions interpretation|Steroid fractions interpretation
C3654153|T201|COMP|73883-1|LNC|Glycolate|Glycolate
C3654154|T201|COMP|73882-3|LNC|Glycolate|Glycolate
C3654155|T201|COMP|73881-5|LNC|Cortisone.free|Cortisone.free
C3654156|T201|COMP|73879-9|LNC|Catecholamine metabolites & creatinine panel|Catecholamine metabolites & creatinine panel
C3654157|T201|COMP|73878-1|LNC|Beta cortolone|Beta cortolone
C3654158|T201|COMP|73877-3|LNC|Beta cortolone|Beta cortolone
C3654159|T201|COMP|73876-5|LNC|Beta cortolone|Beta cortolone
C3654160|T201|COMP|73875-7|LNC|Androstenetriol|Androstenetriol
C3654161|T201|COMP|73874-0|LNC|Androstenetriol|Androstenetriol
C3654162|T201|COMP|73873-2|LNC|Androstenetriol|Androstenetriol
C3654163|T201|COMP|73872-4|LNC|Alpha cortolone|Alpha cortolone
C3654164|T201|COMP|73871-6|LNC|Alpha cortolone|Alpha cortolone
C3654165|T201|COMP|73870-8|LNC|Alpha cortolone|Alpha cortolone
C3654166|T201|COMP|73869-0|LNC|Alpha cortol|Alpha cortol
C3654167|T201|COMP|73868-2|LNC|Alpha cortol|Alpha cortol
C3654168|T201|COMP|73867-4|LNC|Alpha cortol|Alpha cortol
C3654169|T201|COMP|73866-6|LNC|Catecholamines 3 & creatinine panel|Catecholamines 3 & creatinine panel
C3654170|T201|COMP|73865-8|LNC|Catecholamines 3 panel|Catecholamines 3 panel
C3654171|T201|COMP|73864-1|LNC|Allo-tetrahydrocortisol|Allo-tetrahydrocortisol
C3654172|T201|COMP|73863-3|LNC|Allo-tetrahydrocortisol|Allo-tetrahydrocortisol
C3654173|T201|COMP|73861-7|LNC|Allo-tetrahydrocorticosterone|Allo-tetrahydrocorticosterone
C3654174|T201|COMP|73860-9|LNC|Allo-tetrahydrocorticosterone|Allo-tetrahydrocorticosterone
C3654175|T201|COMP|73859-1|LNC|Allo-tetrahydrocorticosterone|Allo-tetrahydrocorticosterone
C3654176|T201|COMP|73858-3|LNC|Allo-pregnanediol|Allo-pregnanediol
C3654177|T201|COMP|73857-5|LNC|Allo-pregnanediol|Allo-pregnanediol
C3654178|T201|COMP|73856-7|LNC|Allo-pregnanediol|Allo-pregnanediol
C3654179|T201|COMP|73855-9|LNC|Aldosterone-18-glucuronide|Aldosterone-18-glucuronide
C3654180|T201|COMP|73854-2|LNC|Aldosterone-18-glucuronide|Aldosterone-18-glucuronide
C3654181|T201|COMP|73853-4|LNC|Aldosterone-18-glucuronide|Aldosterone-18-glucuronide
C3654182|T201|COMP|73852-6|LNC|7-Dehydrocholesterol & 8-Dehydrocholesterol panel|7-Dehydrocholesterol & 8-Dehydrocholesterol panel
C3654183|T201|COMP|73851-8|LNC|18-Beta glycyrrhetinate|18-Beta glycyrrhetinate
C3654184|T201|COMP|73850-0|LNC|18-Beta glycyrrhetinate|18-Beta glycyrrhetinate
C3654185|T201|COMP|73849-2|LNC|16-Ketoandrostenediol|16-Ketoandrostenediol
C3654186|T201|COMP|73848-4|LNC|16-Ketoandrostenediol|16-Ketoandrostenediol
C3654187|T201|COMP|73847-6|LNC|16-Ketoandrostenediol|16-Ketoandrostenediol
C3654188|T201|COMP|73846-8|LNC|16-Alpha hydroxydehydroepiandrosterone|16-Alpha hydroxydehydroepiandrosterone
C3654189|T201|COMP|73845-0|LNC|16-Alpha hydroxydehydroepiandrosterone|16-Alpha hydroxydehydroepiandrosterone
C3654190|T201|COMP|73844-3|LNC|16-Alpha hydroxydehydroepiandrosterone|16-Alpha hydroxydehydroepiandrosterone
C3654191|T201|COMP|73843-5|LNC|Tetrahydrodeoxycortisol|Tetrahydrodeoxycortisol
C3654192|T201|COMP|73842-7|LNC|Tetrahydrodeoxycortisol|Tetrahydrodeoxycortisol
C3654193|T201|COMP|73841-9|LNC|Tetrahydrodeoxycortisol|Tetrahydrodeoxycortisol
C3654194|T201|COMP|73840-1|LNC|11-Dehydrotetrahydrocorticosterone|11-Dehydrotetrahydrocorticosterone
C3654195|T201|COMP|73839-3|LNC|11-Dehydrotetrahydrocorticosterone|11-Dehydrotetrahydrocorticosterone
C3654196|T201|COMP|73838-5|LNC|11-Dehydrotetrahydrocorticosterone|11-Dehydrotetrahydrocorticosterone
C3654197|T201|COMP|73837-7|LNC|Galactose-alpha-1,3-galactose Ab.IgE|Galactose-alpha-1,3-galactose Ab.IgE
C3654198|T201|COMP|73836-9|LNC|Bacteria.fluoroquinolone resistant identified|Bacteria.fluoroquinolone resistant identified
C3654200|T201|COMP|73829-4|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C3654201|T201|COMP|73828-6|LNC|Flunitrazepam|Flunitrazepam
C3654202|T201|COMP|73827-8|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C3654203|T201|COMP|73826-0|LNC|Flurazepam+N-desalkylflurazepam|Flurazepam+N-desalkylflurazepam
C3654204|T201|COMP|73825-2|LNC|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3654205|T201|COMP|73824-5|LNC|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3654206|T201|COMP|73823-7|LNC|Cocaine+Benzoylecgonine|Cocaine+Benzoylecgonine
C3654207|T201|COMP|73822-9|LNC|Fetal chromosome X & Y aneuploidy|Fetal chromosome X & Y aneuploidy
C3654208|T201|COMP|73821-1|LNC|Fetal chromosome X & Y aneuploidy risk|Fetal chromosome X & Y aneuploidy risk
C3654209|T201|COMP|73819-5|LNC|Platelet factor 4 heparin complex induced Ab.IgG|Platelet factor 4 heparin complex induced Ab.IgG
C3654210|T201|COMP|73818-7|LNC|Platelet factor 4 heparin complex induced Ab.IgG|Platelet factor 4 heparin complex induced Ab.IgG
C3654211|T201|COMP|73817-9|LNC|Percent heparin inhibition|Percent heparin inhibition
C3654212|T201|COMP|73816-1|LNC|Platelet factor 4 heparin complex induced Ab.IgG|Platelet factor 4 heparin complex induced Ab.IgG
C3654219|T201|COMP|73809-6|LNC|B cell+T cell crossmatch|B cell+T cell crossmatch
C3654220|T201|COMP|73808-8|LNC|B cell+T cell crossmatch|B cell+T cell crossmatch
C3654221|T201|COMP|73807-0|LNC|B cell+T cell crossmatch.autologous|B cell+T cell crossmatch.autologous
C3654241|T201|COMP|73755-1|LNC|Adenovirus B+E DNA|Adenovirus B+E DNA
C3654242|T201|COMP|73754-4|LNC|Adenovirus C DNA|Adenovirus C DNA
C3654243|T201|COMP|73753-6|LNC|oxyCODONE|oxyCODONE
C3654244|T201|COMP|73752-8|LNC|Reagin Ab & Treponema pallidum Ab.IgG & IgM|Reagin Ab & Treponema pallidum Ab.IgG & IgM
C3654245|T201|COMP|73751-0|LNC|5p15.2 chromosome deletion|5p15.2 chromosome deletion
C3654246|T201|COMP|73750-2|LNC|RAI1 gene 17p11.2 deletion+duplication|RAI1 gene 17p11.2 deletion+duplication
C3654247|T201|COMP|73749-4|LNC|4p16.3 chromosome deletion|4p16.3 chromosome deletion
C3654248|T201|COMP|73748-6|LNC|APOB gene.p.Arg3500Gln & Arg3500Trp|APOB gene.p.Arg3500Gln & Arg3500Trp
C3654249|T201|COMP|73747-8|LNC|Keyhole limpet hemocyanin Ab.IgM|Keyhole limpet hemocyanin Ab.IgM
C3654250|T201|COMP|73746-0|LNC|Keyhole limpet hemocyanin Ab.IgG|Keyhole limpet hemocyanin Ab.IgG
C3654251|T201|COMP|73745-2|LNC|Keyhole limpet hemocyanin Ab.IgA|Keyhole limpet hemocyanin Ab.IgA
C3654258|T201|COMP|73733-8|LNC|Bacteria biotype|Bacteria biotype
C3654260|T201|COMP|73731-2|LNC|Transaldolase|Transaldolase
C3654261|T201|COMP|73730-4|LNC|Lysergate diethylamide|Lysergate diethylamide
C3654262|T201|COMP|73729-6|LNC|Meperidine|Meperidine
C3654263|T201|COMP|73728-8|LNC|Norcocaine|Norcocaine
C3654264|T201|COMP|73727-0|LNC|Methadone|Methadone
C3654265|T201|COMP|73726-2|LNC|Lysergate diethylamide|Lysergate diethylamide
C3654266|T201|COMP|73725-4|LNC|Bile acid panel|Bile acid panel
C3654267|T201|COMP|73724-7|LNC|Bile acid dihydroxy & trihydroxy panel|Bile acid dihydroxy & trihydroxy panel
C3654268|T201|COMP|73723-9|LNC|Riboflavin|Riboflavin
C3654269|T201|COMP|73722-1|LNC|Bile acid|Bile acid
C3654270|T201|COMP|73721-3|LNC|Rocuronium Ab.IgE|Rocuronium Ab.IgE
C3654271|T201|COMP|73720-5|LNC|Pholcodine Ab.IgE|Pholcodine Ab.IgE
C3654272|T201|COMP|73719-7|LNC|Glycine max native (nGly m) 5 Ab.IgE|Glycine max native (nGly m) 5 Ab.IgE
C3654282|T201|COMP|73703-1|LNC|Path report.preliminary diagnosis|Path report.preliminary diagnosis
C3654283|T201|COMP|73702-3|LNC|Neisseria meningitidis serosubtype|Neisseria meningitidis serosubtype
C3654284|T201|COMP|73701-5|LNC|Multiple carboxylase deficiency|Multiple carboxylase deficiency
C3654285|T201|COMP|73699-1|LNC|Number of prior CCHD screens|Number of prior CCHD screens
C3654286|T201|COMP|73697-5|LNC|CCHD newborn screening protocol used|CCHD newborn screening protocol used
C3654290|T201|COMP|73693-4|LNC|African swine fever virus DNA|African swine fever virus DNA
C3654291|T201|COMP|73692-6|LNC|Escitalopram|Escitalopram
C3654292|T201|COMP|73691-8|LNC|Glimepiride|Glimepiride
C3654293|T201|COMP|73690-0|LNC|Nateglinide|Nateglinide
C3654294|T201|COMP|73689-2|LNC|Repaglinide|Repaglinide
C3654295|T201|COMP|73688-4|LNC|Danazol|Danazol
C3654296|T201|COMP|73686-8|LNC|Methylone|Methylone
C3654297|T201|COMP|73685-0|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C3654298|T201|COMP|73684-3|LNC|Atovaquone|Atovaquone
C3654299|T201|COMP|73683-5|LNC|Busulfan^trough|Busulfan^trough
C3654300|T201|COMP|73682-7|LNC|CYP2D6 gene allele 1|CYP2D6 gene allele 1
C3654301|T201|COMP|73681-9|LNC|CYP2D6 gene allele 2|CYP2D6 gene allele 2
C3654302|T201|COMP|73680-1|LNC|Mycophenolate^peak|Mycophenolate^peak
C3654303|T201|COMP|73679-3|LNC|SORAfenib|SORAfenib
C3654304|T201|COMP|73678-5|LNC|Topotecan^trough|Topotecan^trough
C3654305|T201|COMP|73677-7|LNC|Valproate^peak|Valproate^peak
C3654306|T201|COMP|73676-9|LNC|Voriconazole^trough|Voriconazole^trough
C3654307|T201|COMP|73675-1|LNC|Adenosine triphosphate/Adenosine diphosphate|Adenosine triphosphate/Adenosine diphosphate
C3654308|T201|COMP|73967-2|LNC|Noninvasive prenatal fetal aneuploidy test panel|Noninvasive prenatal fetal aneuploidy test panel
C3654309|T201|COMP|73966-4|LNC|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3654313|T201|COMP|73737-9|LNC|Phospholipase A2 receptor Ab.IgG|Phospholipase A2 receptor Ab.IgG
C3654315|T201|COMP|73735-3|LNC|ACADVL gene full mutation analysis|ACADVL gene full mutation analysis
C3654316|T201|COMP|73674-4|LNC|Streptococcus pneumoniae serotype|Streptococcus pneumoniae serotype
C3654317|T201|COMP|73673-6|LNC|Yersinia enterocolitica serotype|Yersinia enterocolitica serotype
C3654318|T201|COMP|73672-8|LNC|Salmonella sp phage type|Salmonella sp phage type
C3654319|T201|COMP|73671-0|LNC|Legionella pneumophila serogroup|Legionella pneumophila serogroup
C3654320|T201|COMP|73670-2|LNC|Bacteria producing coagulase+protein A|Bacteria producing coagulase+protein A
C3654321|T201|COMP|73664-5|LNC|Yersinia adhesion protein YadA|Yersinia adhesion protein YadA
C3654322|T201|COMP|73663-7|LNC|Barbiturates panel|Barbiturates panel
C3654323|T201|COMP|73662-9|LNC|Benzodiazepines panel|Benzodiazepines panel
C3654324|T201|COMP|73661-1|LNC|Methadone panel|Methadone panel
C3654325|T201|COMP|73660-3|LNC|Propoxyphene panel|Propoxyphene panel
C3654326|T201|COMP|73659-5|LNC|HIV 2 subtype|HIV 2 subtype
C3654327|T201|COMP|73658-7|LNC|HIV 1 subtype|HIV 1 subtype
C3654328|T201|COMP|73657-9|LNC|Varicella zoster virus ORF36 genotype|Varicella zoster virus ORF36 genotype
C3654329|T201|COMP|73656-1|LNC|Varicella zoster virus ORF28 genotype|Varicella zoster virus ORF28 genotype
C3654330|T201|COMP|73655-3|LNC|Hepatitis C virus NS5 gene mutations detected|Hepatitis C virus NS5 gene mutations detected
C3654331|T201|COMP|73654-6|LNC|Hepatitis C virus NS3 gene mutations detected|Hepatitis C virus NS3 gene mutations detected
C3654332|T201|COMP|73653-8|LNC|Apramycin|Apramycin
C3654333|T201|COMP|73652-0|LNC|Apramycin|Apramycin
C3654334|T201|COMP|73651-2|LNC|Besifloxacin|Besifloxacin
C3654335|T201|COMP|73650-4|LNC|Ceftaroline|Ceftaroline
C3654336|T201|COMP|73649-6|LNC|Ceftaroline+Avibactam|Ceftaroline+Avibactam
C3654337|T201|COMP|73648-8|LNC|cefTAZidime+Avibactam|cefTAZidime+Avibactam
C3654338|T201|COMP|73647-0|LNC|Ceftolozane+Tazobactam|Ceftolozane+Tazobactam
C3654339|T201|COMP|73646-2|LNC|Danofloxacin|Danofloxacin
C3654340|T201|COMP|73645-4|LNC|Faropenem|Faropenem
C3654341|T201|COMP|73644-7|LNC|Fidaxomicin|Fidaxomicin
C3654342|T201|COMP|73643-9|LNC|Finafloxacin|Finafloxacin
C3654343|T201|COMP|73642-1|LNC|Iclaprim|Iclaprim
C3654344|T201|COMP|73641-3|LNC|Marbofloxacin|Marbofloxacin
C3654345|T201|COMP|73640-5|LNC|Nitazoxanide|Nitazoxanide
C3654346|T201|COMP|73639-7|LNC|Omadacycline|Omadacycline
C3654347|T201|COMP|73638-9|LNC|Ormetroprim+Sulfamethoxazole|Ormetroprim+Sulfamethoxazole
C3654348|T201|COMP|73637-1|LNC|Plazomicin|Plazomicin
C3654349|T201|COMP|73636-3|LNC|Premafloxacin|Premafloxacin
C3654350|T201|COMP|73635-5|LNC|Razupenem|Razupenem
C3654351|T201|COMP|73634-8|LNC|rifAXIMin|rifAXIMin
C3654352|T201|COMP|73633-0|LNC|Sarafloxacin|Sarafloxacin
C3654353|T201|COMP|73632-2|LNC|Solithromycin|Solithromycin
C3654354|T201|COMP|73631-4|LNC|Tedizolid|Tedizolid
C3654355|T201|COMP|73630-6|LNC|Telavancin|Telavancin
C3654356|T201|COMP|73629-8|LNC|Tizoxanide|Tizoxanide
C3654357|T201|COMP|73628-0|LNC|Besifloxacin|Besifloxacin
C3654358|T201|COMP|73627-2|LNC|Ceftaroline|Ceftaroline
C3654359|T201|COMP|73626-4|LNC|Ceftaroline+Avibactam|Ceftaroline+Avibactam
C3654360|T201|COMP|73625-6|LNC|cefTAZidime+Avibactam|cefTAZidime+Avibactam
C3654361|T201|COMP|73624-9|LNC|Ceftolozane+Tazobactam|Ceftolozane+Tazobactam
C3654362|T201|COMP|73623-1|LNC|Danofloxacin|Danofloxacin
C3654363|T201|COMP|73622-3|LNC|Faropenem|Faropenem
C3654364|T201|COMP|73621-5|LNC|Fidaxomicin|Fidaxomicin
C3654365|T201|COMP|73620-7|LNC|Finafloxacin|Finafloxacin
C3654366|T201|COMP|73619-9|LNC|Iclaprim|Iclaprim
C3654367|T201|COMP|73618-1|LNC|Marbofloxacin|Marbofloxacin
C3654368|T201|COMP|73617-3|LNC|Nitazoxanide|Nitazoxanide
C3654369|T201|COMP|73616-5|LNC|Omadacycline|Omadacycline
C3654370|T201|COMP|73615-7|LNC|Ormetroprim+Sulfamethoxazole|Ormetroprim+Sulfamethoxazole
C3654371|T201|COMP|73614-0|LNC|Plazomicin|Plazomicin
C3654372|T201|COMP|73613-2|LNC|Premafloxacin|Premafloxacin
C3654373|T201|COMP|73612-4|LNC|Razupenem|Razupenem
C3654374|T201|COMP|73611-6|LNC|rifAXIMin|rifAXIMin
C3654375|T201|COMP|73609-0|LNC|Solithromycin|Solithromycin
C3654376|T201|COMP|73608-2|LNC|Tedizolid|Tedizolid
C3654377|T201|COMP|73607-4|LNC|Tizoxanide|Tizoxanide
C3654378|T201|COMP|73606-6|LNC|Besifloxacin|Besifloxacin
C3654379|T201|COMP|73605-8|LNC|Ceftaroline|Ceftaroline
C3654380|T201|COMP|73604-1|LNC|Ceftaroline+Avibactam|Ceftaroline+Avibactam
C3654381|T201|COMP|73603-3|LNC|cefTAZidime+Avibactam|cefTAZidime+Avibactam
C3654382|T201|COMP|73602-5|LNC|Ceftolozane+Tazobactam|Ceftolozane+Tazobactam
C3654383|T201|COMP|73601-7|LNC|Danofloxacin|Danofloxacin
C3654384|T201|COMP|73600-9|LNC|Faropenem|Faropenem
C3654385|T201|COMP|73599-3|LNC|Fidaxomicin|Fidaxomicin
C3654386|T201|COMP|73598-5|LNC|Finafloxacin|Finafloxacin
C3654387|T201|COMP|73597-7|LNC|Iclaprim|Iclaprim
C3654388|T201|COMP|73596-9|LNC|Marbofloxacin|Marbofloxacin
C3654389|T201|COMP|73595-1|LNC|Nitazoxanide|Nitazoxanide
C3654390|T201|COMP|73594-4|LNC|Omadacycline|Omadacycline
C3654391|T201|COMP|73593-6|LNC|Ormetroprim+Sulfamethoxazole|Ormetroprim+Sulfamethoxazole
C3654392|T201|COMP|73592-8|LNC|Plazomicin|Plazomicin
C3654393|T201|COMP|73591-0|LNC|Premafloxacin|Premafloxacin
C3654394|T201|COMP|73590-2|LNC|Razupenem|Razupenem
C3654395|T201|COMP|73589-4|LNC|rifAXIMin|rifAXIMin
C3654396|T201|COMP|73588-6|LNC|Sarafloxacin|Sarafloxacin
C3654397|T201|COMP|73587-8|LNC|Solithromycin|Solithromycin
C3654398|T201|COMP|73585-2|LNC|Tizoxanide|Tizoxanide
C3654399|T201|COMP|73584-5|LNC|Norcitalopram|Norcitalopram
C3654400|T201|COMP|73583-7|LNC|Molybdenum/Creatinine|Molybdenum/Creatinine
C3654401|T201|COMP|73581-1|LNC|Anion gap 4|Anion gap 4
C3654402|T201|COMP|73580-3|LNC|Anion gap 4|Anion gap 4
C3654403|T201|COMP|73579-5|LNC|Anion gap 4|Anion gap 4
C3654404|T201|COMP|73573-8|LNC|Magnesium.ionized^^adjusted to pH 7.4|Magnesium.ionized^^adjusted to pH 7.4
C3654405|T201|COMP|73572-0|LNC|Magnesium.ionized|Magnesium.ionized
C3654406|T201|COMP|73571-2|LNC|Osmol gap|Osmol gap
C3654407|T201|COMP|73570-4|LNC|Testosterone/Epitestosterone|Testosterone/Epitestosterone
C3654410|T201|COMP|73567-0|LNC|Propoxyphene|Propoxyphene
C3654411|T201|COMP|73566-2|LNC|Dextrorphan|Dextrorphan
C3654412|T201|COMP|73565-4|LNC|Trenbolone|Trenbolone
C3654413|T201|COMP|73564-7|LNC|Alpha hydroxytriazolam|Alpha hydroxytriazolam
C3654414|T201|COMP|73563-9|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C3654415|T201|COMP|73562-1|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C3654416|T201|COMP|73561-3|LNC|Insulin-like growth factor-I|Insulin-like growth factor-I
C3654417|T201|COMP|73560-5|LNC|Mumps virus Ab.IgG & IgM|Mumps virus Ab.IgG & IgM
C3654418|T201|COMP|73559-7|LNC|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C3654420|T201|COMP|73557-1|LNC|Thyroxine.free|Thyroxine.free
C3654421|T201|COMP|73556-3|LNC|Platelet Ab.IgM|Platelet Ab.IgM
C3654422|T201|COMP|73555-5|LNC|Abciximab induced platelet Ab.IgG|Abciximab induced platelet Ab.IgG
C3654423|T201|COMP|73554-8|LNC|Abciximab induced platelet Ab.IgM|Abciximab induced platelet Ab.IgM
C3654424|T201|COMP|73553-0|LNC|Abciximab induced platelet Ab|Abciximab induced platelet Ab
C3654425|T201|COMP|73552-2|LNC|Drug induced platelet Ab|Drug induced platelet Ab
C3654426|T201|COMP|73551-4|LNC|Acarbose induced platelet Ab.IgG|Acarbose induced platelet Ab.IgG
C3654427|T201|COMP|73550-6|LNC|Acarbose induced platelet Ab.IgM|Acarbose induced platelet Ab.IgM
C3654428|T201|COMP|73549-8|LNC|Acebutolol induced platelet Ab.IgG|Acebutolol induced platelet Ab.IgG
C3654429|T201|COMP|73548-0|LNC|Acebutolol induced platelet Ab.IgM|Acebutolol induced platelet Ab.IgM
C3654430|T201|COMP|73547-2|LNC|Acetaminophen induced platelet Ab.IgM|Acetaminophen induced platelet Ab.IgM
C3654431|T201|COMP|73546-4|LNC|Acetaminophen induced platelet Ab.IgG|Acetaminophen induced platelet Ab.IgG
C3654432|T201|COMP|73545-6|LNC|Acyclovir induced platelet Ab.IgM|Acyclovir induced platelet Ab.IgM
C3654433|T201|COMP|73544-9|LNC|Acyclovir induced platelet Ab.IgG|Acyclovir induced platelet Ab.IgG
C3654434|T201|COMP|73543-1|LNC|Albuterol induced platelet Ab.IgG|Albuterol induced platelet Ab.IgG
C3654435|T201|COMP|73542-3|LNC|Albuterol induced platelet Ab.IgM|Albuterol induced platelet Ab.IgM
C3654436|T201|COMP|73541-5|LNC|Alendronate induced platelet Ab.IgG|Alendronate induced platelet Ab.IgG
C3654437|T201|COMP|73540-7|LNC|Alendronate induced platelet Ab.IgM|Alendronate induced platelet Ab.IgM
C3654438|T201|COMP|73539-9|LNC|Allopurinol induced platelet Ab.IgM|Allopurinol induced platelet Ab.IgM
C3654439|T201|COMP|73538-1|LNC|Allopurinol induced platelet Ab.IgG|Allopurinol induced platelet Ab.IgG
C3654440|T201|COMP|73537-3|LNC|ALPRAZolam induced platelet Ab.IgG|ALPRAZolam induced platelet Ab.IgG
C3654441|T201|COMP|73536-5|LNC|ALPRAZolam induced platelet Ab.IgM|ALPRAZolam induced platelet Ab.IgM
C3654442|T201|COMP|73535-7|LNC|Amiodarone induced platelet Ab.IgM|Amiodarone induced platelet Ab.IgM
C3654443|T201|COMP|73958-1|LNC|Cholesterol esterase|Cholesterol esterase
C3654444|T201|COMP|73957-3|LNC|UR-144 pentanoate|UR-144 pentanoate
C3654445|T201|COMP|73956-5|LNC|JWH-122 5-hydroxypentyl|JWH-122 5-hydroxypentyl
C3654446|T201|COMP|73955-7|LNC|UR-144 4+5-hydroxypentyl|UR-144 4+5-hydroxypentyl
C3654448|T201|COMP|73976-3|LNC|Cells.CD158b/100 cells|Cells.CD158b/100 cells
C3654449|T201|COMP|73975-5|LNC|Cells.CD158a/100 cells|Cells.CD158a/100 cells
C3654450|T201|COMP|73974-8|LNC|Cells.CD158e/100 cells|Cells.CD158e/100 cells
C3654451|T201|COMP|73973-0|LNC|O-nortramadol|O-nortramadol
C3654452|T201|COMP|73834-4|LNC|Bacteria.carbapenem resistant identified|Bacteria.carbapenem resistant identified
C3654453|T201|COMP|73833-6|LNC|Legionella sp Ab|Legionella sp Ab
C3654468|T201|COMP|73578-7|LNC|Anion gap 4|Anion gap 4
C3654469|T201|COMP|73577-9|LNC|Anion gap 4|Anion gap 4
C3654470|T201|COMP|73576-1|LNC|Anion gap 4|Anion gap 4
C3654472|T201|COMP|73574-6|LNC|Acyclovir|Acyclovir
C3654473|T201|COMP|73534-0|LNC|Amiodarone induced platelet Ab.IgG|Amiodarone induced platelet Ab.IgG
C3654474|T201|COMP|73533-2|LNC|Amitriptyline induced platelet Ab.IgM|Amitriptyline induced platelet Ab.IgM
C3654475|T201|COMP|73532-4|LNC|Amitriptyline induced platelet Ab.IgG|Amitriptyline induced platelet Ab.IgG
C3654476|T201|COMP|73531-6|LNC|amLODIPine induced platelet Ab.IgG|amLODIPine induced platelet Ab.IgG
C3654477|T201|COMP|73530-8|LNC|amLODIPine induced platelet Ab.IgM|amLODIPine induced platelet Ab.IgM
C3654478|T201|COMP|73529-0|LNC|amLODIPine+Benazepril induced platelet Ab.IgM|amLODIPine+Benazepril induced platelet Ab.IgM
C3654479|T201|COMP|73528-2|LNC|amLODIPine+Benazepril induced platelet Ab.IgG|amLODIPine+Benazepril induced platelet Ab.IgG
C3654480|T201|COMP|73527-4|LNC|Amoxicillin induced platelet Ab.IgG|Amoxicillin induced platelet Ab.IgG
C3654481|T201|COMP|73526-6|LNC|Amoxicillin induced platelet Ab.IgM|Amoxicillin induced platelet Ab.IgM
C3654482|T201|COMP|73525-8|LNC|Amoxicillin+Clavulanate induced platelet Ab.IgG|Amoxicillin+Clavulanate induced platelet Ab.IgG
C3654483|T201|COMP|73524-1|LNC|Amoxicillin+Clavulanate induced platelet Ab.IgM|Amoxicillin+Clavulanate induced platelet Ab.IgM
C3654484|T201|COMP|73523-3|LNC|Ampicillin induced platelet Ab.IgG|Ampicillin induced platelet Ab.IgG
C3654485|T201|COMP|73522-5|LNC|Ampicillin induced platelet Ab.IgM|Ampicillin induced platelet Ab.IgM
C3654486|T201|COMP|73521-7|LNC|Argatroban induced platelet Ab.IgM|Argatroban induced platelet Ab.IgM
C3654487|T201|COMP|73520-9|LNC|Argatroban induced platelet Ab.IgG|Argatroban induced platelet Ab.IgG
C3654488|T201|COMP|73519-1|LNC|Acetylsalicylate induced platelet Ab.IgM|Acetylsalicylate induced platelet Ab.IgM
C3654489|T201|COMP|73518-3|LNC|Acetylsalicylate induced platelet Ab.IgG|Acetylsalicylate induced platelet Ab.IgG
C3654490|T201|COMP|73517-5|LNC|Atenolol induced platelet Ab.IgM|Atenolol induced platelet Ab.IgM
C3654491|T201|COMP|73516-7|LNC|Atenolol induced platelet Ab.IgG|Atenolol induced platelet Ab.IgG
C3654492|T201|COMP|73515-9|LNC|Atomoxetine induced platelet Ab.IgG|Atomoxetine induced platelet Ab.IgG
C3654493|T201|COMP|73514-2|LNC|Atomoxetine induced platelet Ab.IgM|Atomoxetine induced platelet Ab.IgM
C3654494|T201|COMP|73513-4|LNC|Atorvastatin induced platelet Ab.IgG|Atorvastatin induced platelet Ab.IgG
C3654495|T201|COMP|73512-6|LNC|Atorvastatin induced platelet Ab.IgM|Atorvastatin induced platelet Ab.IgM
C3654496|T201|COMP|73511-8|LNC|Azithromycin induced platelet Ab.IgG|Azithromycin induced platelet Ab.IgG
C3654497|T201|COMP|73506-8|LNC|Benazepril induced platelet Ab.IgG|Benazepril induced platelet Ab.IgG
C3654498|T201|COMP|73505-0|LNC|Benztropine induced platelet Ab.IgM|Benztropine induced platelet Ab.IgM
C3654499|T201|COMP|73504-3|LNC|Benztropine induced platelet Ab.IgG|Benztropine induced platelet Ab.IgG
C3654500|T201|COMP|73503-5|LNC|Bivalirudin induced platelet Ab.IgG|Bivalirudin induced platelet Ab.IgG
C3654501|T201|COMP|73502-7|LNC|Bivalirudin induced platelet Ab.IgM|Bivalirudin induced platelet Ab.IgM
C3654502|T201|COMP|73501-9|LNC|Budesonide induced platelet Ab.IgG|Budesonide induced platelet Ab.IgG
C3654503|T201|COMP|73500-1|LNC|Budesonide induced platelet Ab.IgM|Budesonide induced platelet Ab.IgM
C3654504|T201|COMP|73499-6|LNC|Bumetanide induced platelet Ab.IgG|Bumetanide induced platelet Ab.IgG
C3654505|T201|COMP|73498-8|LNC|Bumetanide induced platelet Ab.IgM|Bumetanide induced platelet Ab.IgM
C3654506|T201|COMP|73497-0|LNC|buPROPion induced platelet Ab.IgM|buPROPion induced platelet Ab.IgM
C3654507|T201|COMP|73496-2|LNC|buPROPion induced platelet Ab.IgG|buPROPion induced platelet Ab.IgG
C3654508|T201|COMP|73495-4|LNC|busPIRone induced platelet Ab.IgG|busPIRone induced platelet Ab.IgG
C3654509|T201|COMP|73494-7|LNC|busPIRone induced platelet Ab.IgM|busPIRone induced platelet Ab.IgM
C3654512|T201|COMP|73491-3|LNC|Candesartan induced platelet Ab.IgG|Candesartan induced platelet Ab.IgG
C3654513|T201|COMP|73490-5|LNC|Candesartan induced platelet Ab.IgM|Candesartan induced platelet Ab.IgM
C3654514|T201|COMP|73489-7|LNC|Captopril induced platelet Ab.IgG|Captopril induced platelet Ab.IgG
C3654515|T201|COMP|73488-9|LNC|Captopril induced platelet Ab.IgM|Captopril induced platelet Ab.IgM
C3654516|T201|COMP|73487-1|LNC|carBAMazepine induced platelet Ab.IgM|carBAMazepine induced platelet Ab.IgM
C3654517|T201|COMP|73486-3|LNC|carBAMazepine induced platelet Ab.IgG|carBAMazepine induced platelet Ab.IgG
C3654518|T201|COMP|73485-5|LNC|Carbidopa induced platelet Ab.IgG|Carbidopa induced platelet Ab.IgG
C3654519|T201|COMP|73484-8|LNC|Carbidopa induced platelet Ab.IgM|Carbidopa induced platelet Ab.IgM
C3654520|T201|COMP|73483-0|LNC|Carisoprodol induced platelet Ab.IgG|Carisoprodol induced platelet Ab.IgG
C3654521|T201|COMP|73482-2|LNC|Carisoprodol induced platelet Ab.IgM|Carisoprodol induced platelet Ab.IgM
C3654522|T201|COMP|73481-4|LNC|Carvedilol induced platelet Ab.IgG|Carvedilol induced platelet Ab.IgG
C3654523|T201|COMP|73480-6|LNC|Carvedilol induced platelet Ab.IgM|Carvedilol induced platelet Ab.IgM
C3654524|T201|COMP|73479-8|LNC|Casanthranol induced platelet Ab.IgG|Casanthranol induced platelet Ab.IgG
C3654525|T201|COMP|73478-0|LNC|Casanthranol induced platelet Ab.IgM|Casanthranol induced platelet Ab.IgM
C3654526|T201|COMP|73477-2|LNC|Caspofungin induced platelet Ab.IgG|Caspofungin induced platelet Ab.IgG
C3654527|T201|COMP|73476-4|LNC|Caspofungin induced platelet Ab.IgM|Caspofungin induced platelet Ab.IgM
C3654528|T201|COMP|73475-6|LNC|Cefadroxil induced platelet Ab.IgG|Cefadroxil induced platelet Ab.IgG
C3654529|T201|COMP|73474-9|LNC|Cefadroxil induced platelet Ab.IgM|Cefadroxil induced platelet Ab.IgM
C3654530|T201|COMP|73473-1|LNC|ceFAZolin induced platelet Ab.IgM|ceFAZolin induced platelet Ab.IgM
C3654531|T201|COMP|73472-3|LNC|ceFAZolin induced platelet Ab.IgG|ceFAZolin induced platelet Ab.IgG
C3654532|T201|COMP|73471-5|LNC|Cefepime induced platelet Ab.IgG|Cefepime induced platelet Ab.IgG
C3654533|T201|COMP|73470-7|LNC|Cefepime induced platelet Ab.IgM|Cefepime induced platelet Ab.IgM
C3654534|T201|COMP|73469-9|LNC|cefTAZidime induced platelet Ab.IgM|cefTAZidime induced platelet Ab.IgM
C3654535|T201|COMP|73468-1|LNC|cefTAZidime induced platelet Ab.IgG|cefTAZidime induced platelet Ab.IgG
C3654536|T201|COMP|73467-3|LNC|Ceftizoxime induced platelet Ab.IgM|Ceftizoxime induced platelet Ab.IgM
C3654537|T201|COMP|73466-5|LNC|Ceftizoxime induced platelet Ab.IgG|Ceftizoxime induced platelet Ab.IgG
C3654538|T201|COMP|73465-7|LNC|cefTRIAXone induced platelet Ab.IgM|cefTRIAXone induced platelet Ab.IgM
C3654539|T201|COMP|73464-0|LNC|cefTRIAXone induced platelet Ab.IgG|cefTRIAXone induced platelet Ab.IgG
C3654540|T201|COMP|73463-2|LNC|Cefuroxime induced platelet Ab.IgM|Cefuroxime induced platelet Ab.IgM
C3654541|T201|COMP|73462-4|LNC|Cefuroxime induced platelet Ab.IgG|Cefuroxime induced platelet Ab.IgG
C3654542|T201|COMP|73461-6|LNC|Celecoxib induced platelet Ab.IgG|Celecoxib induced platelet Ab.IgG
C3654543|T201|COMP|73460-8|LNC|Celecoxib induced platelet Ab.IgM|Celecoxib induced platelet Ab.IgM
C3654544|T201|COMP|73459-0|LNC|Cephalexin induced platelet Ab.IgM|Cephalexin induced platelet Ab.IgM
C3654545|T201|COMP|73453-3|LNC|chlorproPAMIDE induced platelet Ab.IgG|chlorproPAMIDE induced platelet Ab.IgG
C3654546|T201|COMP|73452-5|LNC|chlorproPAMIDE induced platelet Ab.IgM|chlorproPAMIDE induced platelet Ab.IgM
C3654547|T201|COMP|73451-7|LNC|Chlorthalidone induced platelet Ab.IgG|Chlorthalidone induced platelet Ab.IgG
C3654548|T201|COMP|73450-9|LNC|Chlorthalidone induced platelet Ab.IgM|Chlorthalidone induced platelet Ab.IgM
C3654549|T201|COMP|73449-1|LNC|Cilastatin induced platelet Ab.IgM|Cilastatin induced platelet Ab.IgM
C3654550|T201|COMP|73448-3|LNC|Cilastatin induced platelet Ab.IgG|Cilastatin induced platelet Ab.IgG
C3654551|T201|COMP|73447-5|LNC|Cimetidine induced platelet Ab.IgG|Cimetidine induced platelet Ab.IgG
C3654552|T201|COMP|73446-7|LNC|Cimetidine induced platelet Ab.IgM|Cimetidine induced platelet Ab.IgM
C3654553|T201|COMP|73445-9|LNC|Ciprofloxacin induced platelet Ab.IgG|Ciprofloxacin induced platelet Ab.IgG
C3654554|T201|COMP|73444-2|LNC|Ciprofloxacin induced platelet Ab.IgM|Ciprofloxacin induced platelet Ab.IgM
C3654555|T201|COMP|73443-4|LNC|Citalopram induced platelet Ab.IgG|Citalopram induced platelet Ab.IgG
C3654556|T201|COMP|73442-6|LNC|Citalopram induced platelet Ab.IgM|Citalopram induced platelet Ab.IgM
C3654557|T201|COMP|73441-8|LNC|Clarithromycin induced platelet Ab.IgG|Clarithromycin induced platelet Ab.IgG
C3654558|T201|COMP|73440-0|LNC|Clarithromycin induced platelet Ab.IgM|Clarithromycin induced platelet Ab.IgM
C3654559|T201|COMP|73439-2|LNC|Clavulanate induced platelet Ab.IgG|Clavulanate induced platelet Ab.IgG
C3654560|T201|COMP|73438-4|LNC|Clavulanate induced platelet Ab.IgM|Clavulanate induced platelet Ab.IgM
C3654561|T201|COMP|73437-6|LNC|Clindamycin induced platelet Ab.IgG|Clindamycin induced platelet Ab.IgG
C3654562|T201|COMP|73436-8|LNC|Clindamycin induced platelet Ab.IgM|Clindamycin induced platelet Ab.IgM
C3654563|T201|COMP|73435-0|LNC|clonazePAM induced platelet Ab.IgM|clonazePAM induced platelet Ab.IgM
C3654564|T201|COMP|73434-3|LNC|clonazePAM induced platelet Ab.IgG|clonazePAM induced platelet Ab.IgG
C3654565|T201|COMP|73433-5|LNC|cloNIDine induced platelet Ab.IgG|cloNIDine induced platelet Ab.IgG
C3654566|T201|COMP|73432-7|LNC|cloNIDine induced platelet Ab.IgM|cloNIDine induced platelet Ab.IgM
C3654567|T201|COMP|73431-9|LNC|Clopidogrel induced platelet Ab.IgM|Clopidogrel induced platelet Ab.IgM
C3654568|T201|COMP|73430-1|LNC|Clopidogrel induced platelet Ab.IgG|Clopidogrel induced platelet Ab.IgG
C3654569|T201|COMP|73429-3|LNC|Colchicine induced platelet Ab.IgM|Colchicine induced platelet Ab.IgM
C3654570|T201|COMP|73428-5|LNC|Colchicine induced platelet Ab.IgG|Colchicine induced platelet Ab.IgG
C3654571|T201|COMP|73427-7|LNC|cycloSPORINE induced platelet Ab.IgG|cycloSPORINE induced platelet Ab.IgG
C3654572|T201|COMP|73426-9|LNC|cycloSPORINE induced platelet Ab.IgM|cycloSPORINE induced platelet Ab.IgM
C3654573|T201|COMP|73425-1|LNC|Amphetamine induced platelet Ab.IgG|Amphetamine induced platelet Ab.IgG
C3654574|T201|COMP|73424-4|LNC|Amphetamine induced platelet Ab.IgM|Amphetamine induced platelet Ab.IgM
C3654575|T201|COMP|73416-0|LNC|dilTIAZem induced platelet Ab.IgG|dilTIAZem induced platelet Ab.IgG
C3654576|T201|COMP|73415-2|LNC|diphenhydrAMINE induced platelet Ab.IgG|diphenhydrAMINE induced platelet Ab.IgG
C3654577|T201|COMP|73414-5|LNC|diphenhydrAMINE induced platelet Ab.IgM|diphenhydrAMINE induced platelet Ab.IgM
C3654578|T201|COMP|73413-7|LNC|Diphenoxylate+Atropine induced platelet Ab.IgG|Diphenoxylate+Atropine induced platelet Ab.IgG
C3654579|T201|COMP|73412-9|LNC|Diphenoxylate+Atropine induced platelet Ab.IgM|Diphenoxylate+Atropine induced platelet Ab.IgM
C3654580|T201|COMP|73411-1|LNC|Dipyridamole induced platelet Ab.IgG|Dipyridamole induced platelet Ab.IgG
C3654581|T201|COMP|73410-3|LNC|Dipyridamole induced platelet Ab.IgM|Dipyridamole induced platelet Ab.IgM
C3654582|T201|COMP|73409-5|LNC|Docusate induced platelet Ab.IgG|Docusate induced platelet Ab.IgG
C3654583|T201|COMP|73408-7|LNC|Docusate induced platelet Ab.IgM|Docusate induced platelet Ab.IgM
C3654584|T201|COMP|73407-9|LNC|Donepezil induced platelet Ab.IgM|Donepezil induced platelet Ab.IgM
C3654585|T201|COMP|73406-1|LNC|Donepezil induced platelet Ab.IgG|Donepezil induced platelet Ab.IgG
C3654586|T201|COMP|73405-3|LNC|Doxazosin induced platelet Ab.IgM|Doxazosin induced platelet Ab.IgM
C3654587|T201|COMP|73404-6|LNC|Doxazosin induced platelet Ab.IgG|Doxazosin induced platelet Ab.IgG
C3654588|T201|COMP|73403-8|LNC|Doxycycline induced platelet Ab.IgM|Doxycycline induced platelet Ab.IgM
C3654589|T201|COMP|73402-0|LNC|Doxycycline induced platelet Ab.IgG|Doxycycline induced platelet Ab.IgG
C3654590|T201|COMP|73401-2|LNC|Enalapril induced platelet Ab.IgG|Enalapril induced platelet Ab.IgG
C3654591|T201|COMP|73400-4|LNC|Enalapril induced platelet Ab.IgM|Enalapril induced platelet Ab.IgM
C3654592|T201|COMP|73399-8|LNC|Erythropoietin induced platelet Ab.IgG|Erythropoietin induced platelet Ab.IgG
C3654593|T201|COMP|73398-0|LNC|Erythropoietin induced platelet Ab.IgM|Erythropoietin induced platelet Ab.IgM
C3654594|T201|COMP|73397-2|LNC|Eptifibatide induced platelet Ab.IgG|Eptifibatide induced platelet Ab.IgG
C3654595|T201|COMP|73396-4|LNC|Eptifibatide induced platelet Ab.IgM|Eptifibatide induced platelet Ab.IgM
C3654596|T201|COMP|73395-6|LNC|Erythromycin induced platelet Ab.IgG|Erythromycin induced platelet Ab.IgG
C3654597|T201|COMP|73394-9|LNC|Erythromycin induced platelet Ab.IgM|Erythromycin induced platelet Ab.IgM
C3654598|T201|COMP|73393-1|LNC|Escitalopram induced platelet Ab.IgG|Escitalopram induced platelet Ab.IgG
C3654599|T201|COMP|73392-3|LNC|Escitalopram induced platelet Ab.IgM|Escitalopram induced platelet Ab.IgM
C3654600|T201|COMP|73391-5|LNC|Esomeprazole induced platelet Ab.IgG|Esomeprazole induced platelet Ab.IgG
C3654601|T201|COMP|73390-7|LNC|Esomeprazole induced platelet Ab.IgM|Esomeprazole induced platelet Ab.IgM
C3654602|T201|COMP|73384-0|LNC|Fenofibrate induced platelet Ab.IgM|Fenofibrate induced platelet Ab.IgM
C3654603|T201|COMP|73383-2|LNC|fentaNYL induced platelet Ab.IgM|fentaNYL induced platelet Ab.IgM
C3654604|T201|COMP|73382-4|LNC|fentaNYL induced platelet Ab.IgG|fentaNYL induced platelet Ab.IgG
C3654605|T201|COMP|73381-6|LNC|Fexofenadine induced platelet Ab.IgG|Fexofenadine induced platelet Ab.IgG
C3654606|T201|COMP|73380-8|LNC|Fexofenadine induced platelet Ab.IgM|Fexofenadine induced platelet Ab.IgM
C3654607|T201|COMP|73379-0|LNC|Finasteride induced platelet Ab.IgG|Finasteride induced platelet Ab.IgG
C3654608|T201|COMP|73378-2|LNC|Finasteride induced platelet Ab.IgM|Finasteride induced platelet Ab.IgM
C3654609|T201|COMP|73377-4|LNC|Fluconazole induced platelet Ab.IgM|Fluconazole induced platelet Ab.IgM
C3654610|T201|COMP|73376-6|LNC|Fluconazole induced platelet Ab.IgG|Fluconazole induced platelet Ab.IgG
C3654611|T201|COMP|73375-8|LNC|FLUoxetine induced platelet Ab.IgG|FLUoxetine induced platelet Ab.IgG
C3654612|T201|COMP|73374-1|LNC|FLUoxetine induced platelet Ab.IgM|FLUoxetine induced platelet Ab.IgM
C3654613|T201|COMP|73373-3|LNC|Fluvastatin induced platelet Ab.IgM|Fluvastatin induced platelet Ab.IgM
C3654614|T201|COMP|73372-5|LNC|Fluvastatin induced platelet Ab.IgG|Fluvastatin induced platelet Ab.IgG
C3654615|T201|COMP|73371-7|LNC|Fosinopril induced platelet Ab.IgG|Fosinopril induced platelet Ab.IgG
C3654616|T201|COMP|73365-9|LNC|Gentamicin induced platelet Ab.IgG|Gentamicin induced platelet Ab.IgG
C3654617|T201|COMP|73364-2|LNC|Gentamicin induced platelet Ab.IgM|Gentamicin induced platelet Ab.IgM
C3654618|T201|COMP|73363-4|LNC|Glimepiride induced platelet Ab.IgG|Glimepiride induced platelet Ab.IgG
C3654619|T201|COMP|73362-6|LNC|Glimepiride induced platelet Ab.IgM|Glimepiride induced platelet Ab.IgM
C3654620|T201|COMP|73361-8|LNC|glipiZIDE induced platelet Ab.IgM|glipiZIDE induced platelet Ab.IgM
C3654621|T201|COMP|73360-0|LNC|glipiZIDE induced platelet Ab.IgG|glipiZIDE induced platelet Ab.IgG
C3654622|T201|COMP|73359-2|LNC|glyBURIDE induced platelet Ab.IgG|glyBURIDE induced platelet Ab.IgG
C3654623|T201|COMP|73358-4|LNC|glyBURIDE induced platelet Ab.IgM|glyBURIDE induced platelet Ab.IgM
C3654624|T201|COMP|73357-6|LNC|Haloperidol induced platelet Ab.IgM|Haloperidol induced platelet Ab.IgM
C3654625|T201|COMP|73356-8|LNC|Haloperidol induced platelet Ab.IgG|Haloperidol induced platelet Ab.IgG
C3654626|T201|COMP|73355-0|LNC|hydrALAZINE induced platelet Ab.IgG|hydrALAZINE induced platelet Ab.IgG
C3654627|T201|COMP|73354-3|LNC|hydrALAZINE induced platelet Ab.IgM|hydrALAZINE induced platelet Ab.IgM
C3654628|T201|COMP|73353-5|LNC|hydroCHLOROthiazide induced platelet Ab.IgG|hydroCHLOROthiazide induced platelet Ab.IgG
C3654629|T201|COMP|73352-7|LNC|hydroCHLOROthiazide induced platelet Ab.IgM|hydroCHLOROthiazide induced platelet Ab.IgM
C3654632|T201|COMP|73349-3|LNC|HYDROcodone induced platelet Ab.IgG|HYDROcodone induced platelet Ab.IgG
C3654633|T201|COMP|73348-5|LNC|HYDROcodone induced platelet Ab.IgM|HYDROcodone induced platelet Ab.IgM
C3654634|T201|COMP|73347-7|LNC|HYDROcodone+Acetaminophen induced platelet Ab.IgG|HYDROcodone+Acetaminophen induced platelet Ab.IgG
C3654635|T201|COMP|73346-9|LNC|HYDROcodone+Acetaminophen induced platelet Ab.IgM|HYDROcodone+Acetaminophen induced platelet Ab.IgM
C3654638|T201|COMP|73343-6|LNC|Hydrocortisone induced platelet Ab.IgM|Hydrocortisone induced platelet Ab.IgM
C3654639|T201|COMP|73342-8|LNC|Hydrocortisone induced platelet Ab.IgG|Hydrocortisone induced platelet Ab.IgG
C3654640|T201|COMP|73341-0|LNC|HYDROmorphone induced platelet Ab.IgG|HYDROmorphone induced platelet Ab.IgG
C3654641|T201|COMP|73340-2|LNC|HYDROmorphone induced platelet Ab.IgM|HYDROmorphone induced platelet Ab.IgM
C3654642|T201|COMP|73339-4|LNC|hydrOXYzine induced platelet Ab.IgG|hydrOXYzine induced platelet Ab.IgG
C3654643|T201|COMP|73338-6|LNC|hydrOXYzine induced platelet Ab.IgM|hydrOXYzine induced platelet Ab.IgM
C3654644|T201|COMP|73337-8|LNC|Ibuprofen induced platelet Ab.IgM|Ibuprofen induced platelet Ab.IgM
C3654645|T201|COMP|73336-0|LNC|Ibuprofen induced platelet Ab.IgG|Ibuprofen induced platelet Ab.IgG
C3654646|T201|COMP|73335-2|LNC|Imipenem induced platelet Ab.IgM|Imipenem induced platelet Ab.IgM
C3654647|T201|COMP|73334-5|LNC|Imipenem induced platelet Ab.IgG|Imipenem induced platelet Ab.IgG
C3654648|T201|COMP|73333-7|LNC|Imipenem+Cilastatin induced platelet Ab.IgG|Imipenem+Cilastatin induced platelet Ab.IgG
C3654649|T201|COMP|73332-9|LNC|Imipenem+Cilastatin induced platelet Ab.IgM|Imipenem+Cilastatin induced platelet Ab.IgM
C3654650|T201|COMP|73331-1|LNC|Ipratropium induced platelet Ab.IgG|Ipratropium induced platelet Ab.IgG
C3654651|T201|COMP|73330-3|LNC|Ipratropium induced platelet Ab.IgM|Ipratropium induced platelet Ab.IgM
C3654652|T201|COMP|73329-5|LNC|Irbesartan induced platelet Ab.IgG|Irbesartan induced platelet Ab.IgG
C3654653|T201|COMP|73328-7|LNC|Irbesartan induced platelet Ab.IgM|Irbesartan induced platelet Ab.IgM
C3654656|T201|COMP|73325-3|LNC|Isosorbide induced platelet Ab.IgG|Isosorbide induced platelet Ab.IgG
C3654657|T201|COMP|73324-6|LNC|Isosorbide induced platelet Ab.IgM|Isosorbide induced platelet Ab.IgM
C3654658|T201|COMP|73319-6|LNC|Lansoprazole induced platelet Ab.IgG|Lansoprazole induced platelet Ab.IgG
C3654659|T201|COMP|73318-8|LNC|Lansoprazole induced platelet Ab.IgM|Lansoprazole induced platelet Ab.IgM
C3654660|T201|COMP|73317-0|LNC|Lepirudin induced platelet Ab.IgG|Lepirudin induced platelet Ab.IgG
C3654661|T201|COMP|73316-2|LNC|Lepirudin induced platelet Ab.IgM|Lepirudin induced platelet Ab.IgM
C3654662|T201|COMP|73315-4|LNC|Leuprolide induced platelet Ab.IgG|Leuprolide induced platelet Ab.IgG
C3654663|T201|COMP|73314-7|LNC|Leuprolide induced platelet Ab.IgM|Leuprolide induced platelet Ab.IgM
C3654664|T201|COMP|73313-9|LNC|Levalbuterol induced platelet Ab.IgG|Levalbuterol induced platelet Ab.IgG
C3654665|T201|COMP|73312-1|LNC|Levalbuterol induced platelet Ab.IgM|Levalbuterol induced platelet Ab.IgM
C3654666|T201|COMP|73311-3|LNC|levETIRAcetam induced platelet Ab.IgG|levETIRAcetam induced platelet Ab.IgG
C3654667|T201|COMP|73310-5|LNC|levETIRAcetam induced platelet Ab.IgM|levETIRAcetam induced platelet Ab.IgM
C3654668|T201|COMP|73309-7|LNC|Levodopa induced platelet Ab.IgG|Levodopa induced platelet Ab.IgG
C3654669|T201|COMP|73308-9|LNC|Levodopa induced platelet Ab.IgM|Levodopa induced platelet Ab.IgM
C3654670|T201|COMP|73307-1|LNC|levoFLOXacin induced platelet Ab.IgG|levoFLOXacin induced platelet Ab.IgG
C3654671|T201|COMP|73306-3|LNC|levoFLOXacin induced platelet Ab.IgM|levoFLOXacin induced platelet Ab.IgM
C3654672|T201|COMP|73305-5|LNC|Lidocaine induced platelet Ab.IgG|Lidocaine induced platelet Ab.IgG
C3654673|T201|COMP|73304-8|LNC|Lidocaine induced platelet Ab.IgM|Lidocaine induced platelet Ab.IgM
C3654674|T201|COMP|73303-0|LNC|Linezolid induced platelet Ab.IgM|Linezolid induced platelet Ab.IgM
C3654675|T201|COMP|73302-2|LNC|Linezolid induced platelet Ab.IgG|Linezolid induced platelet Ab.IgG
C3654676|T201|COMP|73301-4|LNC|Lisinopril induced platelet Ab.IgG|Lisinopril induced platelet Ab.IgG
C3654677|T201|COMP|73295-8|LNC|LORazepam induced platelet Ab.IgG|LORazepam induced platelet Ab.IgG
C3654678|T201|COMP|73294-1|LNC|LORazepam induced platelet Ab.IgM|LORazepam induced platelet Ab.IgM
C3654679|T201|COMP|73293-3|LNC|Losartan induced platelet Ab.IgM|Losartan induced platelet Ab.IgM
C3654680|T201|COMP|73292-5|LNC|Losartan induced platelet Ab.IgG|Losartan induced platelet Ab.IgG
C3654681|T201|COMP|73291-7|LNC|Lovastatin induced platelet Ab.IgG|Lovastatin induced platelet Ab.IgG
C3654682|T201|COMP|73290-9|LNC|Lovastatin induced platelet Ab.IgM|Lovastatin induced platelet Ab.IgM
C3654683|T201|COMP|73289-1|LNC|Meropenem induced platelet Ab.IgG|Meropenem induced platelet Ab.IgG
C3654684|T201|COMP|73288-3|LNC|Meropenem induced platelet Ab.IgM|Meropenem induced platelet Ab.IgM
C3654685|T201|COMP|73287-5|LNC|metFORMIN induced platelet Ab.IgG|metFORMIN induced platelet Ab.IgG
C3654686|T201|COMP|73286-7|LNC|metFORMIN induced platelet Ab.IgM|metFORMIN induced platelet Ab.IgM
C3654687|T201|COMP|73285-9|LNC|Methocarbamol induced platelet Ab.IgG|Methocarbamol induced platelet Ab.IgG
C3654688|T201|COMP|73284-2|LNC|Methocarbamol induced platelet Ab.IgM|Methocarbamol induced platelet Ab.IgM
C3654689|T201|COMP|73283-4|LNC|Methotrexate induced platelet Ab.IgG|Methotrexate induced platelet Ab.IgG
C3654690|T201|COMP|73282-6|LNC|Methotrexate induced platelet Ab.IgM|Methotrexate induced platelet Ab.IgM
C3654691|T201|COMP|73281-8|LNC|Methyldopa induced platelet Ab.IgG|Methyldopa induced platelet Ab.IgG
C3654692|T201|COMP|73280-0|LNC|Methyldopa induced platelet Ab.IgM|Methyldopa induced platelet Ab.IgM
C3654693|T201|COMP|73279-2|LNC|Methylphenidate induced platelet Ab.IgM|Methylphenidate induced platelet Ab.IgM
C3654694|T201|COMP|73278-4|LNC|Methylphenidate induced platelet Ab.IgG|Methylphenidate induced platelet Ab.IgG
C3654695|T201|COMP|73277-6|LNC|Methylprednisolone induced platelet Ab.IgG|Methylprednisolone induced platelet Ab.IgG
C3654696|T201|COMP|73276-8|LNC|Methylprednisolone induced platelet Ab.IgM|Methylprednisolone induced platelet Ab.IgM
C3654697|T201|COMP|73275-0|LNC|Metoclopramide induced platelet Ab.IgG|Metoclopramide induced platelet Ab.IgG
C3654698|T201|COMP|73274-3|LNC|Metoclopramide induced platelet Ab.IgM|Metoclopramide induced platelet Ab.IgM
C3654699|T201|COMP|73273-5|LNC|Metoprolol induced platelet Ab.IgG|Metoprolol induced platelet Ab.IgG
C3654700|T201|COMP|73272-7|LNC|Metoprolol induced platelet Ab.IgM|Metoprolol induced platelet Ab.IgM
C3654701|T201|COMP|73271-9|LNC|metroNIDAZOLE induced platelet Ab.IgG|metroNIDAZOLE induced platelet Ab.IgG
C3654702|T201|COMP|73270-1|LNC|metroNIDAZOLE induced platelet Ab.IgM|metroNIDAZOLE induced platelet Ab.IgM
C3654703|T201|COMP|73269-3|LNC|Midazolam induced platelet Ab.IgG|Midazolam induced platelet Ab.IgG
C3654704|T201|COMP|73268-5|LNC|Midazolam induced platelet Ab.IgM|Midazolam induced platelet Ab.IgM
C3654705|T201|COMP|73267-7|LNC|Milrinone induced platelet Ab.IgM|Milrinone induced platelet Ab.IgM
C3654706|T201|COMP|73266-9|LNC|Milrinone induced platelet Ab.IgG|Milrinone induced platelet Ab.IgG
C3654707|T201|COMP|73265-1|LNC|Minocycline induced platelet Ab.IgG|Minocycline induced platelet Ab.IgG
C3654708|T201|COMP|73264-4|LNC|Minocycline induced platelet Ab.IgM|Minocycline induced platelet Ab.IgM
C3654709|T201|COMP|73263-6|LNC|Minoxidil induced platelet Ab.IgG|Minoxidil induced platelet Ab.IgG
C3654710|T201|COMP|73262-8|LNC|Minoxidil induced platelet Ab.IgM|Minoxidil induced platelet Ab.IgM
C3654711|T201|COMP|73261-0|LNC|Mirtazapine induced platelet Ab.IgG|Mirtazapine induced platelet Ab.IgG
C3654712|T201|COMP|73260-2|LNC|Mirtazapine induced platelet Ab.IgM|Mirtazapine induced platelet Ab.IgM
C3654713|T201|COMP|73259-4|LNC|Montelukast induced platelet Ab.IgG|Montelukast induced platelet Ab.IgG
C3654714|T201|COMP|73258-6|LNC|Montelukast induced platelet Ab.IgM|Montelukast induced platelet Ab.IgM
C3654715|T201|COMP|73257-8|LNC|Morphine induced platelet Ab.IgG|Morphine induced platelet Ab.IgG
C3654716|T201|COMP|73256-0|LNC|Morphine induced platelet Ab.IgM|Morphine induced platelet Ab.IgM
C3654717|T201|COMP|73255-2|LNC|Moxifloxacin induced platelet Ab.IgM|Moxifloxacin induced platelet Ab.IgM
C3654718|T201|COMP|73254-5|LNC|Moxifloxacin induced platelet Ab.IgG|Moxifloxacin induced platelet Ab.IgG
C3654719|T201|COMP|73253-7|LNC|Mycophenolate induced platelet Ab.IgG|Mycophenolate induced platelet Ab.IgG
C3654720|T201|COMP|73252-9|LNC|Mycophenolate induced platelet Ab.IgM|Mycophenolate induced platelet Ab.IgM
C3654721|T201|COMP|73251-1|LNC|Nafcillin induced platelet Ab.IgG|Nafcillin induced platelet Ab.IgG
C3654722|T201|COMP|73250-3|LNC|Nafcillin induced platelet Ab.IgM|Nafcillin induced platelet Ab.IgM
C3654723|T201|COMP|73249-5|LNC|Naproxen induced platelet Ab.IgG|Naproxen induced platelet Ab.IgG
C3654724|T201|COMP|73248-7|LNC|Naproxen induced platelet Ab.IgM|Naproxen induced platelet Ab.IgM
C3654725|T201|COMP|73247-9|LNC|Niacin+Lovastatin induced platelet Ab.IgG|Niacin+Lovastatin induced platelet Ab.IgG
C3654726|T201|COMP|73246-1|LNC|Niacin+Lovastatin induced platelet Ab.IgM|Niacin+Lovastatin induced platelet Ab.IgM
C3654727|T201|COMP|73245-3|LNC|NIFEdipine induced platelet Ab.IgG|NIFEdipine induced platelet Ab.IgG
C3654728|T201|COMP|73244-6|LNC|NIFEdipine induced platelet Ab.IgM|NIFEdipine induced platelet Ab.IgM
C3654729|T201|COMP|73243-8|LNC|Nitrofurantoin induced platelet Ab.IgG|Nitrofurantoin induced platelet Ab.IgG
C3654730|T201|COMP|73242-0|LNC|Nitrofurantoin induced platelet Ab.IgM|Nitrofurantoin induced platelet Ab.IgM
C3654731|T201|COMP|73235-4|LNC|OLANZapine induced platelet Ab.IgG|OLANZapine induced platelet Ab.IgG
C3654732|T201|COMP|73234-7|LNC|OLANZapine induced platelet Ab.IgM|OLANZapine induced platelet Ab.IgM
C3654733|T201|COMP|73233-9|LNC|Omeprazole induced platelet Ab.IgG|Omeprazole induced platelet Ab.IgG
C3654734|T201|COMP|73232-1|LNC|Omeprazole induced platelet Ab.IgM|Omeprazole induced platelet Ab.IgM
C3654735|T201|COMP|73231-3|LNC|Ondansetron induced platelet Ab.IgG|Ondansetron induced platelet Ab.IgG
C3654736|T201|COMP|73230-5|LNC|Ondansetron induced platelet Ab.IgM|Ondansetron induced platelet Ab.IgM
C3654737|T201|COMP|73229-7|LNC|Oxacillin induced platelet Ab.IgG|Oxacillin induced platelet Ab.IgG
C3654738|T201|COMP|73228-9|LNC|Oxacillin induced platelet Ab.IgM|Oxacillin induced platelet Ab.IgM
C3654739|T201|COMP|73227-1|LNC|Oxaliplatin induced platelet Ab.IgG|Oxaliplatin induced platelet Ab.IgG
C3654740|T201|COMP|73226-3|LNC|Oxaliplatin induced platelet Ab.IgM|Oxaliplatin induced platelet Ab.IgM
C3654741|T201|COMP|73225-5|LNC|OXcarbazepine induced platelet Ab.IgM|OXcarbazepine induced platelet Ab.IgM
C3654742|T201|COMP|73224-8|LNC|OXcarbazepine induced platelet Ab.IgG|OXcarbazepine induced platelet Ab.IgG
C3654743|T201|COMP|73223-0|LNC|oxyCODONE induced platelet Ab.IgM|oxyCODONE induced platelet Ab.IgM
C3654744|T201|COMP|73222-2|LNC|oxyCODONE induced platelet Ab.IgG|oxyCODONE induced platelet Ab.IgG
C3654747|T201|COMP|73219-8|LNC|Pantoprazole induced platelet Ab.IgG|Pantoprazole induced platelet Ab.IgG
C3654748|T201|COMP|73218-0|LNC|Pantoprazole induced platelet Ab.IgM|Pantoprazole induced platelet Ab.IgM
C3654749|T201|COMP|73217-2|LNC|Papaverine induced platelet Ab.IgM|Papaverine induced platelet Ab.IgM
C3654750|T201|COMP|73216-4|LNC|Papaverine induced platelet Ab.IgG|Papaverine induced platelet Ab.IgG
C3654751|T201|COMP|73215-6|LNC|PARoxetine induced platelet Ab.IgG|PARoxetine induced platelet Ab.IgG
C3654752|T201|COMP|73214-9|LNC|PARoxetine induced platelet Ab.IgM|PARoxetine induced platelet Ab.IgM
C3654753|T201|COMP|73213-1|LNC|Penicillin induced platelet Ab.IgG|Penicillin induced platelet Ab.IgG
C3654754|T201|COMP|73212-3|LNC|Penicillin induced platelet Ab.IgM|Penicillin induced platelet Ab.IgM
C3654755|T201|COMP|73211-5|LNC|Perphenazine induced platelet Ab.IgG|Perphenazine induced platelet Ab.IgG
C3654756|T201|COMP|73210-7|LNC|Perphenazine induced platelet Ab.IgM|Perphenazine induced platelet Ab.IgM
C3654757|T201|COMP|73209-9|LNC|PHENobarbital induced platelet Ab.IgG|PHENobarbital induced platelet Ab.IgG
C3654758|T201|COMP|73208-1|LNC|PHENobarbital induced platelet Ab.IgM|PHENobarbital induced platelet Ab.IgM
C3654759|T201|COMP|73207-3|LNC|Phenytoin induced platelet Ab.IgM|Phenytoin induced platelet Ab.IgM
C3654760|T201|COMP|73206-5|LNC|Phenytoin induced platelet Ab.IgG|Phenytoin induced platelet Ab.IgG
C3654761|T201|COMP|73205-7|LNC|Pioglitazone induced platelet Ab.IgG|Pioglitazone induced platelet Ab.IgG
C3654762|T201|COMP|73204-0|LNC|Pioglitazone induced platelet Ab.IgM|Pioglitazone induced platelet Ab.IgM
C3654763|T201|COMP|73203-2|LNC|Piperacillin induced platelet Ab.IgM|Piperacillin induced platelet Ab.IgM
C3654764|T201|COMP|73202-4|LNC|Piperacillin induced platelet Ab.IgG|Piperacillin induced platelet Ab.IgG
C3654765|T201|COMP|73201-6|LNC|Piperacillin+Tazobactam induced platelet Ab.IgG|Piperacillin+Tazobactam induced platelet Ab.IgG
C3654766|T201|COMP|73200-8|LNC|Piperacillin+Tazobactam induced platelet Ab.IgM|Piperacillin+Tazobactam induced platelet Ab.IgM
C3654767|T201|COMP|73199-2|LNC|Pravastatin induced platelet Ab.IgG|Pravastatin induced platelet Ab.IgG
C3654768|T201|COMP|73198-4|LNC|Pravastatin induced platelet Ab.IgM|Pravastatin induced platelet Ab.IgM
C3654769|T201|COMP|73197-6|LNC|predniSONE induced platelet Ab.IgG|predniSONE induced platelet Ab.IgG
C3654770|T201|COMP|73196-8|LNC|predniSONE induced platelet Ab.IgM|predniSONE induced platelet Ab.IgM
C3654771|T201|COMP|73195-0|LNC|Primidone induced platelet Ab.IgG|Primidone induced platelet Ab.IgG
C3654772|T201|COMP|73194-3|LNC|Primidone induced platelet Ab.IgM|Primidone induced platelet Ab.IgM
C3654773|T201|COMP|73193-5|LNC|Procainamide induced platelet Ab.IgG|Procainamide induced platelet Ab.IgG
C3654774|T201|COMP|73192-7|LNC|Procainamide induced platelet Ab.IgM|Procainamide induced platelet Ab.IgM
C3654775|T201|COMP|73191-9|LNC|Propoxyphene induced platelet Ab.IgM|Propoxyphene induced platelet Ab.IgM
C3654776|T201|COMP|73190-1|LNC|Propoxyphene induced platelet Ab.IgG|Propoxyphene induced platelet Ab.IgG
C3654779|T201|COMP|73187-7|LNC|Propranolol induced platelet Ab.IgG|Propranolol induced platelet Ab.IgG
C3654780|T201|COMP|73186-9|LNC|Propranolol induced platelet Ab.IgM|Propranolol induced platelet Ab.IgM
C3654781|T201|COMP|73185-1|LNC|Pseudoephedrine induced platelet Ab.IgG|Pseudoephedrine induced platelet Ab.IgG
C3654782|T201|COMP|73184-4|LNC|Pseudoephedrine induced platelet Ab.IgM|Pseudoephedrine induced platelet Ab.IgM
C3654783|T201|COMP|73183-6|LNC|QUEtiapine induced platelet Ab.IgG|QUEtiapine induced platelet Ab.IgG
C3654784|T201|COMP|73182-8|LNC|QUEtiapine induced platelet Ab.IgM|QUEtiapine induced platelet Ab.IgM
C3654785|T201|COMP|73181-0|LNC|Quinapril induced platelet Ab.IgG|Quinapril induced platelet Ab.IgG
C3654786|T201|COMP|73180-2|LNC|Quinapril induced platelet Ab.IgM|Quinapril induced platelet Ab.IgM
C3654787|T201|COMP|73179-4|LNC|quiNIDine induced platelet Ab.IgM|quiNIDine induced platelet Ab.IgM
C3654788|T201|COMP|73178-6|LNC|quiNIDine induced platelet Ab.IgG|quiNIDine induced platelet Ab.IgG
C3654789|T201|COMP|73177-8|LNC|quiNINE induced platelet Ab.IgG|quiNINE induced platelet Ab.IgG
C3654790|T201|COMP|73176-0|LNC|quiNINE induced platelet Ab.IgM|quiNINE induced platelet Ab.IgM
C3654791|T201|COMP|73175-2|LNC|RABEprazole induced platelet Ab.IgM|RABEprazole induced platelet Ab.IgM
C3654792|T201|COMP|73174-5|LNC|RABEprazole induced platelet Ab.IgG|RABEprazole induced platelet Ab.IgG
C3654793|T201|COMP|73173-7|LNC|Raloxifene induced platelet Ab.IgG|Raloxifene induced platelet Ab.IgG
C3654794|T201|COMP|73172-9|LNC|Raloxifene induced platelet Ab.IgM|Raloxifene induced platelet Ab.IgM
C3654795|T201|COMP|73171-1|LNC|Ramipril induced platelet Ab.IgG|Ramipril induced platelet Ab.IgG
C3654796|T201|COMP|73170-3|LNC|Ramipril induced platelet Ab.IgM|Ramipril induced platelet Ab.IgM
C3654797|T201|COMP|73169-5|LNC|raNITIdine induced platelet Ab.IgM|raNITIdine induced platelet Ab.IgM
C3654798|T201|COMP|73168-7|LNC|raNITIdine induced platelet Ab.IgG|raNITIdine induced platelet Ab.IgG
C3654799|T201|COMP|73167-9|LNC|rifAMPin induced platelet Ab.IgM|rifAMPin induced platelet Ab.IgM
C3654800|T201|COMP|73166-1|LNC|rifAMPin induced platelet Ab.IgG|rifAMPin induced platelet Ab.IgG
C3654801|T201|COMP|73165-3|LNC|Risedronate induced platelet Ab.IgG|Risedronate induced platelet Ab.IgG
C3654802|T201|COMP|73164-6|LNC|Risedronate induced platelet Ab.IgM|Risedronate induced platelet Ab.IgM
C3654803|T201|COMP|73163-8|LNC|risperiDONE induced platelet Ab.IgG|risperiDONE induced platelet Ab.IgG
C3654804|T201|COMP|73162-0|LNC|risperiDONE induced platelet Ab.IgM|risperiDONE induced platelet Ab.IgM
C3654805|T201|COMP|73161-2|LNC|Rofecoxib induced platelet Ab.IgM|Rofecoxib induced platelet Ab.IgM
C3654806|T201|COMP|73160-4|LNC|Rofecoxib induced platelet Ab.IgG|Rofecoxib induced platelet Ab.IgG
C3654807|T201|COMP|73159-6|LNC|Rosiglitazone induced platelet Ab.IgG|Rosiglitazone induced platelet Ab.IgG
C3654808|T201|COMP|73158-8|LNC|Rosiglitazone induced platelet Ab.IgM|Rosiglitazone induced platelet Ab.IgM
C3654809|T201|COMP|73157-0|LNC|Rosuvastatin induced platelet Ab.IgG|Rosuvastatin induced platelet Ab.IgG
C3654810|T201|COMP|73156-2|LNC|Rosuvastatin induced platelet Ab.IgM|Rosuvastatin induced platelet Ab.IgM
C3654811|T201|COMP|73155-4|LNC|Sertraline induced platelet Ab.IgG|Sertraline induced platelet Ab.IgG
C3654812|T201|COMP|73154-7|LNC|Sertraline induced platelet Ab.IgM|Sertraline induced platelet Ab.IgM
C3654813|T201|COMP|73153-9|LNC|Sildenafil citrate induced platelet Ab.IgG|Sildenafil citrate induced platelet Ab.IgG
C3654814|T201|COMP|73152-1|LNC|Sildenafil citrate induced platelet Ab.IgM|Sildenafil citrate induced platelet Ab.IgM
C3654815|T201|COMP|73151-3|LNC|Simethicone induced platelet Ab.IgG|Simethicone induced platelet Ab.IgG
C3654816|T201|COMP|73150-5|LNC|Simethicone induced platelet Ab.IgM|Simethicone induced platelet Ab.IgM
C3654817|T201|COMP|73149-7|LNC|Simvastatin induced platelet Ab.IgG|Simvastatin induced platelet Ab.IgG
C3654818|T201|COMP|73148-9|LNC|Simvastatin induced platelet Ab.IgM|Simvastatin induced platelet Ab.IgM
C3654819|T201|COMP|73147-1|LNC|Sotalol induced platelet Ab.IgM|Sotalol induced platelet Ab.IgM
C3654820|T201|COMP|73146-3|LNC|Sotalol induced platelet Ab.IgG|Sotalol induced platelet Ab.IgG
C3654821|T201|COMP|73145-5|LNC|Spironolactone induced platelet Ab.IgM|Spironolactone induced platelet Ab.IgM
C3654822|T201|COMP|73144-8|LNC|Spironolactone induced platelet Ab.IgG|Spironolactone induced platelet Ab.IgG
C3654823|T201|COMP|73143-0|LNC|Sucralfate induced platelet Ab.IgG|Sucralfate induced platelet Ab.IgG
C3654824|T201|COMP|73142-2|LNC|Sucralfate induced platelet Ab.IgM|Sucralfate induced platelet Ab.IgM
C3654825|T201|COMP|73141-4|LNC|Sulfamethoxazole induced platelet Ab.IgM|Sulfamethoxazole induced platelet Ab.IgM
C3654826|T201|COMP|73140-6|LNC|Sulfamethoxazole induced platelet Ab.IgG|Sulfamethoxazole induced platelet Ab.IgG
C3654827|T201|COMP|73139-8|LNC|sulfaSALAzine induced platelet Ab.IgG|sulfaSALAzine induced platelet Ab.IgG
C3654828|T201|COMP|73138-0|LNC|sulfaSALAzine induced platelet Ab.IgM|sulfaSALAzine induced platelet Ab.IgM
C3654829|T201|COMP|73137-2|LNC|sulfiSOXAZOLE induced platelet Ab.IgG|sulfiSOXAZOLE induced platelet Ab.IgG
C3654830|T201|COMP|73136-4|LNC|sulfiSOXAZOLE induced platelet Ab.IgM|sulfiSOXAZOLE induced platelet Ab.IgM
C3654831|T201|COMP|73135-6|LNC|Sulindac induced platelet Ab.IgG|Sulindac induced platelet Ab.IgG
C3654832|T201|COMP|73134-9|LNC|Sulindac induced platelet Ab.IgM|Sulindac induced platelet Ab.IgM
C3654833|T201|COMP|73133-1|LNC|Tacrolimus induced platelet Ab.IgG|Tacrolimus induced platelet Ab.IgG
C3654834|T201|COMP|73132-3|LNC|Tacrolimus induced platelet Ab.IgM|Tacrolimus induced platelet Ab.IgM
C3654835|T201|COMP|73131-5|LNC|Tamoxifen induced platelet Ab.IgG|Tamoxifen induced platelet Ab.IgG
C3654836|T201|COMP|73130-7|LNC|Tamoxifen induced platelet Ab.IgM|Tamoxifen induced platelet Ab.IgM
C3654837|T201|COMP|73129-9|LNC|Tamsulosin induced platelet Ab.IgG|Tamsulosin induced platelet Ab.IgG
C3654838|T201|COMP|73128-1|LNC|Tamsulosin induced platelet Ab.IgM|Tamsulosin induced platelet Ab.IgM
C3654839|T201|COMP|73127-3|LNC|Tazobactam induced platelet Ab.IgG|Tazobactam induced platelet Ab.IgG
C3654840|T201|COMP|73126-5|LNC|Tazobactam induced platelet Ab.IgM|Tazobactam induced platelet Ab.IgM
C3654841|T201|COMP|73125-7|LNC|Telmisartan induced platelet Ab.IgG|Telmisartan induced platelet Ab.IgG
C3654842|T201|COMP|73124-0|LNC|Telmisartan induced platelet Ab.IgM|Telmisartan induced platelet Ab.IgM
C3654843|T201|COMP|73123-2|LNC|Terazosin induced platelet Ab.IgG|Terazosin induced platelet Ab.IgG
C3654844|T201|COMP|73122-4|LNC|Terazosin induced platelet Ab.IgM|Terazosin induced platelet Ab.IgM
C3654845|T201|COMP|73121-6|LNC|Tetracycline induced platelet Ab.IgG|Tetracycline induced platelet Ab.IgG
C3654846|T201|COMP|73120-8|LNC|Tetracycline induced platelet Ab.IgM|Tetracycline induced platelet Ab.IgM
C3654847|T201|COMP|73119-0|LNC|Timolol induced platelet Ab.IgG|Timolol induced platelet Ab.IgG
C3654848|T201|COMP|73118-2|LNC|Timolol induced platelet Ab.IgM|Timolol induced platelet Ab.IgM
C3654849|T201|COMP|73117-4|LNC|Tirofiban induced platelet Ab.IgG|Tirofiban induced platelet Ab.IgG
C3654850|T201|COMP|73116-6|LNC|Tirofiban induced platelet Ab.IgM|Tirofiban induced platelet Ab.IgM
C3654851|T201|COMP|73115-8|LNC|Tobramycin induced platelet Ab.IgG|Tobramycin induced platelet Ab.IgG
C3654852|T201|COMP|73114-1|LNC|Tobramycin induced platelet Ab.IgM|Tobramycin induced platelet Ab.IgM
C3654853|T201|COMP|73113-3|LNC|Tolterodine induced platelet Ab.IgM|Tolterodine induced platelet Ab.IgM
C3654854|T201|COMP|73112-5|LNC|Tolterodine induced platelet Ab.IgG|Tolterodine induced platelet Ab.IgG
C3654855|T201|COMP|73111-7|LNC|Topiramate induced platelet Ab.IgG|Topiramate induced platelet Ab.IgG
C3654856|T201|COMP|73110-9|LNC|Topiramate induced platelet Ab.IgM|Topiramate induced platelet Ab.IgM
C3654857|T201|COMP|73109-1|LNC|traMADol induced platelet Ab.IgG|traMADol induced platelet Ab.IgG
C3654858|T201|COMP|73108-3|LNC|traMADol induced platelet Ab.IgM|traMADol induced platelet Ab.IgM
C3654859|T201|COMP|73107-5|LNC|Triamcinolone induced platelet Ab.IgG|Triamcinolone induced platelet Ab.IgG
C3654860|T201|COMP|73106-7|LNC|Triamcinolone induced platelet Ab.IgM|Triamcinolone induced platelet Ab.IgM
C3654861|T201|COMP|73105-9|LNC|Triamterene induced platelet Ab.IgM|Triamterene induced platelet Ab.IgM
C3654862|T201|COMP|73104-2|LNC|Triamterene induced platelet Ab.IgG|Triamterene induced platelet Ab.IgG
C3654863|T201|COMP|73103-4|LNC|Triazolam induced platelet Ab.IgM|Triazolam induced platelet Ab.IgM
C3654864|T201|COMP|73102-6|LNC|Triazolam induced platelet Ab.IgG|Triazolam induced platelet Ab.IgG
C3654865|T201|COMP|73101-8|LNC|Trimethoprim induced platelet Ab.IgM|Trimethoprim induced platelet Ab.IgM
C3654866|T201|COMP|73100-0|LNC|Trimethoprim induced platelet Ab.IgG|Trimethoprim induced platelet Ab.IgG
C3654867|T201|COMP|73099-4|LNC|Ursodeoxycholate induced platelet Ab.IgM|Ursodeoxycholate induced platelet Ab.IgM
C3654868|T201|COMP|73098-6|LNC|Ursodeoxycholate induced platelet Ab.IgG|Ursodeoxycholate induced platelet Ab.IgG
C3654869|T201|COMP|73097-8|LNC|valACYclovir induced platelet Ab.IgM|valACYclovir induced platelet Ab.IgM
C3654870|T201|COMP|73091-1|LNC|Valproate induced platelet Ab.IgG|Valproate induced platelet Ab.IgG
C3654871|T201|COMP|73090-3|LNC|Valproate induced platelet Ab.IgM|Valproate induced platelet Ab.IgM
C3654872|T201|COMP|73089-5|LNC|Valsartan induced platelet Ab.IgM|Valsartan induced platelet Ab.IgM
C3654873|T201|COMP|73088-7|LNC|Valsartan induced platelet Ab.IgG|Valsartan induced platelet Ab.IgG
C3654874|T201|COMP|73087-9|LNC|Vancomycin induced platelet Ab.IgM|Vancomycin induced platelet Ab.IgM
C3654875|T201|COMP|73086-1|LNC|Vancomycin induced platelet Ab.IgG|Vancomycin induced platelet Ab.IgG
C3654876|T201|COMP|73085-3|LNC|Venlafaxine induced platelet Ab.IgG|Venlafaxine induced platelet Ab.IgG
C3654877|T201|COMP|73084-6|LNC|Venlafaxine induced platelet Ab.IgM|Venlafaxine induced platelet Ab.IgM
C3654878|T201|COMP|73083-8|LNC|Verapamil induced platelet Ab.IgG|Verapamil induced platelet Ab.IgG
C3654879|T201|COMP|73082-0|LNC|Verapamil induced platelet Ab.IgM|Verapamil induced platelet Ab.IgM
C3654880|T201|COMP|73081-2|LNC|Voriconazole induced platelet Ab.IgG|Voriconazole induced platelet Ab.IgG
C3654881|T201|COMP|73080-4|LNC|Voriconazole induced platelet Ab.IgM|Voriconazole induced platelet Ab.IgM
C3654882|T201|COMP|73079-6|LNC|Warfarin induced platelet Ab.IgM|Warfarin induced platelet Ab.IgM
C3654883|T201|COMP|73078-8|LNC|Warfarin induced platelet Ab.IgG|Warfarin induced platelet Ab.IgG
C3654884|T201|COMP|73077-0|LNC|Neutrophil Ab.IgG|Neutrophil Ab.IgG
C3654885|T201|COMP|73076-2|LNC|Neutrophil Ab.IgM|Neutrophil Ab.IgM
C3654886|T201|COMP|73075-4|LNC|Drug induced neutrophil Ab|Drug induced neutrophil Ab
C3654887|T201|COMP|73074-7|LNC|Acetaminophen induced neutrophil Ab.IgM|Acetaminophen induced neutrophil Ab.IgM
C3654888|T201|COMP|73073-9|LNC|Acetaminophen induced neutrophil Ab.IgG|Acetaminophen induced neutrophil Ab.IgG
C3654889|T201|COMP|73072-1|LNC|Alendronate induced neutrophil Ab.IgG|Alendronate induced neutrophil Ab.IgG
C3654890|T201|COMP|73071-3|LNC|Alendronate induced neutrophil Ab.IgM|Alendronate induced neutrophil Ab.IgM
C3654891|T201|COMP|73070-5|LNC|Allopurinol induced neutrophil Ab.IgG|Allopurinol induced neutrophil Ab.IgG
C3654892|T201|COMP|73069-7|LNC|Allopurinol induced neutrophil Ab.IgM|Allopurinol induced neutrophil Ab.IgM
C3654893|T201|COMP|73068-9|LNC|Amiodarone induced neutrophil Ab.IgG|Amiodarone induced neutrophil Ab.IgG
C3654894|T201|COMP|73067-1|LNC|Amiodarone induced neutrophil Ab.IgM|Amiodarone induced neutrophil Ab.IgM
C3654895|T201|COMP|73066-3|LNC|Amitriptyline induced neutrophil Ab.IgG|Amitriptyline induced neutrophil Ab.IgG
C3654896|T201|COMP|73065-5|LNC|Amitriptyline induced neutrophil Ab.IgM|Amitriptyline induced neutrophil Ab.IgM
C3654897|T201|COMP|73064-8|LNC|amLODIPine induced neutrophil Ab.IgG|amLODIPine induced neutrophil Ab.IgG
C3654898|T201|COMP|73063-0|LNC|amLODIPine induced neutrophil Ab.IgM|amLODIPine induced neutrophil Ab.IgM
C3654899|T201|COMP|73062-2|LNC|Amoxicillin induced neutrophil Ab.IgG|Amoxicillin induced neutrophil Ab.IgG
C3654900|T201|COMP|73061-4|LNC|Amoxicillin induced neutrophil Ab.IgM|Amoxicillin induced neutrophil Ab.IgM
C3654901|T201|COMP|73060-6|LNC|Ampicillin induced neutrophil Ab.IgG|Ampicillin induced neutrophil Ab.IgG
C3654902|T201|COMP|73059-8|LNC|Ampicillin induced neutrophil Ab.IgM|Ampicillin induced neutrophil Ab.IgM
C3654903|T201|COMP|73058-0|LNC|Acetylsalicylate induced neutrophil Ab.IgG|Acetylsalicylate induced neutrophil Ab.IgG
C3654904|T201|COMP|73057-2|LNC|Acetylsalicylate induced neutrophil Ab.IgM|Acetylsalicylate induced neutrophil Ab.IgM
C3654905|T201|COMP|73056-4|LNC|Atenolol induced neutrophil Ab.IgG|Atenolol induced neutrophil Ab.IgG
C3654906|T201|COMP|73055-6|LNC|Atenolol induced neutrophil Ab.IgM|Atenolol induced neutrophil Ab.IgM
C3654907|T201|COMP|73054-9|LNC|Atorvastatin induced neutrophil Ab.IgG|Atorvastatin induced neutrophil Ab.IgG
C3654908|T201|COMP|73053-1|LNC|Atorvastatin induced neutrophil Ab.IgM|Atorvastatin induced neutrophil Ab.IgM
C3654909|T201|COMP|73052-3|LNC|buPROPion induced neutrophil Ab.IgG|buPROPion induced neutrophil Ab.IgG
C3654910|T201|COMP|73051-5|LNC|buPROPion induced neutrophil Ab.IgM|buPROPion induced neutrophil Ab.IgM
C3654911|T201|COMP|73050-7|LNC|carBAMazepine induced neutrophil Ab.IgG|carBAMazepine induced neutrophil Ab.IgG
C3654912|T201|COMP|73049-9|LNC|carBAMazepine induced neutrophil Ab.IgM|carBAMazepine induced neutrophil Ab.IgM
C3654913|T201|COMP|73048-1|LNC|ceFAZolin induced neutrophil Ab.IgG|ceFAZolin induced neutrophil Ab.IgG
C3654914|T201|COMP|73047-3|LNC|ceFAZolin induced neutrophil Ab.IgM|ceFAZolin induced neutrophil Ab.IgM
C3654915|T201|COMP|73046-5|LNC|Cefepime induced neutrophil Ab.IgG|Cefepime induced neutrophil Ab.IgG
C3654916|T201|COMP|73045-7|LNC|Cefepime induced neutrophil Ab.IgM|Cefepime induced neutrophil Ab.IgM
C3654917|T201|COMP|73044-0|LNC|cefTAZidime induced neutrophil Ab.IgG|cefTAZidime induced neutrophil Ab.IgG
C3654918|T201|COMP|73043-2|LNC|cefTAZidime induced neutrophil Ab.IgM|cefTAZidime induced neutrophil Ab.IgM
C3654919|T201|COMP|73042-4|LNC|cefTRIAXone induced neutrophil Ab.IgG|cefTRIAXone induced neutrophil Ab.IgG
C3654920|T201|COMP|73041-6|LNC|cefTRIAXone induced neutrophil Ab.IgM|cefTRIAXone induced neutrophil Ab.IgM
C3654921|T201|COMP|73040-8|LNC|Celecoxib induced neutrophil Ab.IgG|Celecoxib induced neutrophil Ab.IgG
C3654922|T201|COMP|73039-0|LNC|Celecoxib induced neutrophil Ab.IgM|Celecoxib induced neutrophil Ab.IgM
C3654923|T201|COMP|73038-2|LNC|Ciprofloxacin induced neutrophil Ab.IgG|Ciprofloxacin induced neutrophil Ab.IgG
C3654924|T201|COMP|73037-4|LNC|Ciprofloxacin induced neutrophil Ab.IgM|Ciprofloxacin induced neutrophil Ab.IgM
C3654925|T201|COMP|73036-6|LNC|Citalopram induced neutrophil Ab.IgG|Citalopram induced neutrophil Ab.IgG
C3654926|T201|COMP|73035-8|LNC|Citalopram induced neutrophil Ab.IgM|Citalopram induced neutrophil Ab.IgM
C3654927|T201|COMP|73034-1|LNC|Clindamycin induced neutrophil Ab.IgG|Clindamycin induced neutrophil Ab.IgG
C3654928|T201|COMP|73033-3|LNC|Clindamycin induced neutrophil Ab.IgM|Clindamycin induced neutrophil Ab.IgM
C3654929|T201|COMP|73032-5|LNC|cloNIDine induced neutrophil Ab.IgG|cloNIDine induced neutrophil Ab.IgG
C3654930|T201|COMP|73031-7|LNC|cloNIDine induced neutrophil Ab.IgM|cloNIDine induced neutrophil Ab.IgM
C3654931|T201|COMP|73030-9|LNC|Clopidogrel induced neutrophil Ab.IgG|Clopidogrel induced neutrophil Ab.IgG
C3654932|T201|COMP|73029-1|LNC|Clopidogrel induced neutrophil Ab.IgM|Clopidogrel induced neutrophil Ab.IgM
C3654933|T201|COMP|73028-3|LNC|Enalapril induced neutrophil Ab.IgG|Enalapril induced neutrophil Ab.IgG
C3654934|T201|COMP|73027-5|LNC|Enalapril induced neutrophil Ab.IgM|Enalapril induced neutrophil Ab.IgM
C3654935|T201|COMP|73026-7|LNC|Escitalopram induced neutrophil Ab.IgG|Escitalopram induced neutrophil Ab.IgG
C3654936|T201|COMP|73025-9|LNC|Escitalopram induced neutrophil Ab.IgM|Escitalopram induced neutrophil Ab.IgM
C3654937|T201|COMP|73024-2|LNC|Fenofibrate induced neutrophil Ab.IgG|Fenofibrate induced neutrophil Ab.IgG
C3654938|T201|COMP|73015-0|LNC|Gabapentin induced neutrophil Ab.IgM|Gabapentin induced neutrophil Ab.IgM
C3654939|T201|COMP|73014-3|LNC|Gentamicin induced neutrophil Ab.IgG|Gentamicin induced neutrophil Ab.IgG
C3654940|T201|COMP|73013-5|LNC|Gentamicin induced neutrophil Ab.IgM|Gentamicin induced neutrophil Ab.IgM
C3654941|T201|COMP|73012-7|LNC|hydroCHLOROthiazide induced neutrophil Ab.IgG|hydroCHLOROthiazide induced neutrophil Ab.IgG
C3654942|T201|COMP|73006-9|LNC|levETIRAcetam induced neutrophil Ab.IgG|levETIRAcetam induced neutrophil Ab.IgG
C3654943|T201|COMP|73005-1|LNC|levETIRAcetam induced neutrophil Ab.IgM|levETIRAcetam induced neutrophil Ab.IgM
C3654944|T201|COMP|73004-4|LNC|levoFLOXacin induced neutrophil Ab.IgG|levoFLOXacin induced neutrophil Ab.IgG
C3654945|T201|COMP|73003-6|LNC|levoFLOXacin induced neutrophil Ab.IgM|levoFLOXacin induced neutrophil Ab.IgM
C3654946|T201|COMP|73002-8|LNC|Lisinopril induced neutrophil Ab.IgG|Lisinopril induced neutrophil Ab.IgG
C3654947|T201|COMP|73001-0|LNC|Lisinopril induced neutrophil Ab.IgM|Lisinopril induced neutrophil Ab.IgM
C3654948|T201|COMP|73000-2|LNC|Loratadine induced neutrophil Ab.IgG|Loratadine induced neutrophil Ab.IgG
C3654949|T201|COMP|72999-6|LNC|Loratadine induced neutrophil Ab.IgM|Loratadine induced neutrophil Ab.IgM
C3654950|T201|COMP|72998-8|LNC|Losartan induced neutrophil Ab.IgG|Losartan induced neutrophil Ab.IgG
C3654951|T201|COMP|72997-0|LNC|Losartan induced neutrophil Ab.IgM|Losartan induced neutrophil Ab.IgM
C3654952|T201|COMP|72996-2|LNC|metFORMIN induced neutrophil Ab.IgG|metFORMIN induced neutrophil Ab.IgG
C3654953|T201|COMP|72995-4|LNC|metFORMIN induced neutrophil Ab.IgM|metFORMIN induced neutrophil Ab.IgM
C3654954|T201|COMP|72994-7|LNC|Methylphenidate induced neutrophil Ab.IgG|Methylphenidate induced neutrophil Ab.IgG
C3654955|T201|COMP|72993-9|LNC|Methylphenidate induced neutrophil Ab.IgM|Methylphenidate induced neutrophil Ab.IgM
C3654956|T201|COMP|72992-1|LNC|Metoclopramide induced neutrophil Ab.IgG|Metoclopramide induced neutrophil Ab.IgG
C3654957|T201|COMP|72991-3|LNC|Metoclopramide induced neutrophil Ab.IgM|Metoclopramide induced neutrophil Ab.IgM
C3654958|T201|COMP|72990-5|LNC|Metoprolol induced neutrophil Ab.IgG|Metoprolol induced neutrophil Ab.IgG
C3654959|T201|COMP|72989-7|LNC|Metoprolol induced neutrophil Ab.IgM|Metoprolol induced neutrophil Ab.IgM
C3654960|T201|COMP|72988-9|LNC|Montelukast induced neutrophil Ab.IgG|Montelukast induced neutrophil Ab.IgG
C3654961|T201|COMP|72987-1|LNC|Montelukast induced neutrophil Ab.IgM|Montelukast induced neutrophil Ab.IgM
C3654962|T201|COMP|72986-3|LNC|Mycophenolate induced neutrophil Ab.IgG|Mycophenolate induced neutrophil Ab.IgG
C3654963|T201|COMP|72985-5|LNC|Mycophenolate induced neutrophil Ab.IgM|Mycophenolate induced neutrophil Ab.IgM
C3654964|T201|COMP|72984-8|LNC|OLANZapine induced neutrophil Ab.IgG|OLANZapine induced neutrophil Ab.IgG
C3654965|T201|COMP|72983-0|LNC|OLANZapine induced neutrophil Ab.IgM|OLANZapine induced neutrophil Ab.IgM
C3654966|T201|COMP|72982-2|LNC|Omeprazole induced neutrophil Ab.IgG|Omeprazole induced neutrophil Ab.IgG
C3654967|T201|COMP|72981-4|LNC|Omeprazole induced neutrophil Ab.IgM|Omeprazole induced neutrophil Ab.IgM
C3654968|T201|COMP|72980-6|LNC|Pantoprazole induced neutrophil Ab.IgG|Pantoprazole induced neutrophil Ab.IgG
C3654969|T201|COMP|72979-8|LNC|Pantoprazole induced neutrophil Ab.IgM|Pantoprazole induced neutrophil Ab.IgM
C3654970|T201|COMP|72978-0|LNC|PARoxetine induced neutrophil Ab.IgG|PARoxetine induced neutrophil Ab.IgG
C3654971|T201|COMP|72977-2|LNC|PARoxetine induced neutrophil Ab.IgM|PARoxetine induced neutrophil Ab.IgM
C3654972|T201|COMP|72976-4|LNC|Penicillin induced neutrophil Ab.IgG|Penicillin induced neutrophil Ab.IgG
C3654973|T201|COMP|72975-6|LNC|Penicillin induced neutrophil Ab.IgM|Penicillin induced neutrophil Ab.IgM
C3654974|T201|COMP|72974-9|LNC|PHENobarbital induced neutrophil Ab.IgG|PHENobarbital induced neutrophil Ab.IgG
C3654975|T201|COMP|72973-1|LNC|PHENobarbital induced neutrophil Ab.IgM|PHENobarbital induced neutrophil Ab.IgM
C3654976|T201|COMP|72972-3|LNC|Phenytoin induced neutrophil Ab.IgG|Phenytoin induced neutrophil Ab.IgG
C3654977|T201|COMP|72971-5|LNC|Phenytoin induced neutrophil Ab.IgM|Phenytoin induced neutrophil Ab.IgM
C3654978|T201|COMP|72964-0|LNC|quiNINE induced neutrophil Ab.IgG|quiNINE induced neutrophil Ab.IgG
C3654979|T201|COMP|72963-2|LNC|quiNINE induced neutrophil Ab.IgM|quiNINE induced neutrophil Ab.IgM
C3654980|T201|COMP|72962-4|LNC|Ramipril induced neutrophil Ab.IgG|Ramipril induced neutrophil Ab.IgG
C3654981|T201|COMP|72961-6|LNC|Ramipril induced neutrophil Ab.IgM|Ramipril induced neutrophil Ab.IgM
C3654982|T201|COMP|72960-8|LNC|raNITIdine induced neutrophil Ab.IgG|raNITIdine induced neutrophil Ab.IgG
C3654983|T201|COMP|72959-0|LNC|raNITIdine induced neutrophil Ab.IgM|raNITIdine induced neutrophil Ab.IgM
C3654984|T201|COMP|72958-2|LNC|risperiDONE induced neutrophil Ab.IgG|risperiDONE induced neutrophil Ab.IgG
C3654985|T201|COMP|72957-4|LNC|risperiDONE induced neutrophil Ab.IgM|risperiDONE induced neutrophil Ab.IgM
C3654986|T201|COMP|72956-6|LNC|Sertraline induced neutrophil Ab.IgG|Sertraline induced neutrophil Ab.IgG
C3654987|T201|COMP|72955-8|LNC|Sertraline induced neutrophil Ab.IgM|Sertraline induced neutrophil Ab.IgM
C3654988|T201|COMP|72954-1|LNC|Sildenafil citrate induced neutrophil Ab.IgG|Sildenafil citrate induced neutrophil Ab.IgG
C3654989|T201|COMP|72953-3|LNC|Sildenafil citrate induced neutrophil Ab.IgM|Sildenafil citrate induced neutrophil Ab.IgM
C3654990|T201|COMP|72952-5|LNC|Simvastatin induced neutrophil Ab.IgG|Simvastatin induced neutrophil Ab.IgG
C3654991|T201|COMP|72951-7|LNC|Simvastatin induced neutrophil Ab.IgM|Simvastatin induced neutrophil Ab.IgM
C3654992|T201|COMP|72950-9|LNC|Spironolactone induced neutrophil Ab.IgG|Spironolactone induced neutrophil Ab.IgG
C3654993|T201|COMP|72949-1|LNC|Spironolactone induced neutrophil Ab.IgM|Spironolactone induced neutrophil Ab.IgM
C3654994|T201|COMP|72948-3|LNC|Sulfamethoxazole induced neutrophil Ab.IgG|Sulfamethoxazole induced neutrophil Ab.IgG
C3654995|T201|COMP|72947-5|LNC|Sulfamethoxazole induced neutrophil Ab.IgM|Sulfamethoxazole induced neutrophil Ab.IgM
C3654996|T201|COMP|72946-7|LNC|Tacrolimus induced neutrophil Ab.IgG|Tacrolimus induced neutrophil Ab.IgG
C3654997|T201|COMP|72945-9|LNC|Tacrolimus induced neutrophil Ab.IgM|Tacrolimus induced neutrophil Ab.IgM
C3654998|T201|COMP|72944-2|LNC|Tazobactam induced neutrophil Ab.IgG|Tazobactam induced neutrophil Ab.IgG
C3654999|T201|COMP|72943-4|LNC|Tazobactam induced neutrophil Ab.IgM|Tazobactam induced neutrophil Ab.IgM
C3655000|T201|COMP|72942-6|LNC|Terazosin induced neutrophil Ab.IgG|Terazosin induced neutrophil Ab.IgG
C3655001|T201|COMP|72941-8|LNC|Terazosin induced neutrophil Ab.IgM|Terazosin induced neutrophil Ab.IgM
C3655002|T201|COMP|72940-0|LNC|Topiramate induced neutrophil Ab.IgG|Topiramate induced neutrophil Ab.IgG
C3655003|T201|COMP|72939-2|LNC|Topiramate induced neutrophil Ab.IgM|Topiramate induced neutrophil Ab.IgM
C3655004|T201|COMP|72938-4|LNC|Trimethoprim induced neutrophil Ab.IgG|Trimethoprim induced neutrophil Ab.IgG
C3655005|T201|COMP|72937-6|LNC|Trimethoprim induced neutrophil Ab.IgM|Trimethoprim induced neutrophil Ab.IgM
C3655006|T201|COMP|72936-8|LNC|Valproate induced neutrophil Ab.IgG|Valproate induced neutrophil Ab.IgG
C3655007|T201|COMP|72935-0|LNC|Valproate induced neutrophil Ab.IgM|Valproate induced neutrophil Ab.IgM
C3655008|T201|COMP|72917-8|LNC|HNA 5 genotype|HNA 5 genotype
C3655009|T201|COMP|72916-0|LNC|HNA 1b-1b Ab|HNA 1b-1b Ab
C3655010|T201|COMP|72915-2|LNC|HNA 1a-1b Ab|HNA 1a-1b Ab
C3655011|T201|COMP|72914-5|LNC|HNA 1c Ab|HNA 1c Ab
C3655012|T201|COMP|72913-7|LNC|HNA 2 Ab|HNA 2 Ab
C3655013|T201|COMP|72912-9|LNC|HNA 4a-4a Ab|HNA 4a-4a Ab
C3655014|T201|COMP|72911-1|LNC|HNA 4b-4b Ab|HNA 4b-4b Ab
C3655015|T201|COMP|72910-3|LNC|HNA 4a-4b Ab|HNA 4a-4b Ab
C3655016|T201|COMP|72909-5|LNC|Drug induced neutrophil Ab panel|Drug induced neutrophil Ab panel
C3655017|T201|COMP|72908-7|LNC|Drug induced platelet Ab panel|Drug induced platelet Ab panel
C3655018|T201|COMP|72906-1|LNC|HNA Ab panel|HNA Ab panel
C3655019|T201|COMP|72905-3|LNC|Neutrophil Ab & HLA Ab screen panel|Neutrophil Ab & HLA Ab screen panel
C3655020|T201|COMP|72904-6|LNC|Formate|Formate
C3655021|T201|COMP|72903-8|LNC|Urea|Urea
C3655022|T201|COMP|72902-0|LNC|Insulin^1H post 75 g glucose PO|Insulin^1H post 75 g glucose PO
C3655023|T201|COMP|72901-2|LNC|Insulin^2H post 75 g glucose PO|Insulin^2H post 75 g glucose PO
C3655024|T201|COMP|72900-4|LNC|Insulin^3H post 75 g glucose PO|Insulin^3H post 75 g glucose PO
C3655025|T201|COMP|72898-0|LNC|Bilirubin|Bilirubin
C3655026|T201|COMP|72897-2|LNC|Xanthine|Xanthine
C3655027|T201|COMP|72896-4|LNC|Glucose^15M post dose lactose PO|Glucose^15M post dose lactose PO
C3655028|T201|COMP|72895-6|LNC|Glucose^2.5H post dose lactose PO|Glucose^2.5H post dose lactose PO
C3655029|T201|COMP|72894-9|LNC|Telavancin|Telavancin
C3655030|T201|COMP|72893-1|LNC|Doripenem|Doripenem
C3655032|T201|COMP|72891-5|LNC|Staphylococcus protein A spa gene|Staphylococcus protein A spa gene
C3655033|T201|COMP|72890-7|LNC|Progesterone.free/Progesterone.total|Progesterone.free/Progesterone.total
C3655034|T201|COMP|72889-9|LNC|Progesterone.free|Progesterone.free
C3655038|T201|COMP|72885-7|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C3655039|T201|COMP|72884-0|LNC|CYP1A2 gene targeted mutation analysis|CYP1A2 gene targeted mutation analysis
C3655040|T201|COMP|72883-2|LNC|CYP2E1 gene targeted mutation analysis|CYP2E1 gene targeted mutation analysis
C3655041|T201|COMP|72882-4|LNC|CYP2B6 gene targeted mutation analysis|CYP2B6 gene targeted mutation analysis
C3655042|T201|COMP|72881-6|LNC|UGT2B15 gene targeted mutation analysis|UGT2B15 gene targeted mutation analysis
C3655048|T201|COMP|72875-8|LNC|JWH-073 butanol|JWH-073 butanol
C3655049|T201|COMP|72874-1|LNC|JWH-073 butanol/Creatinine|JWH-073 butanol/Creatinine
C3655050|T201|COMP|72873-3|LNC|Estradiol|Estradiol
C3655051|T201|COMP|72872-5|LNC|MCM6 gene.c.-13910C>T & -13915T>G|MCM6 gene.c.-13910C>T & -13915T>G
C3655061|T201|COMP|72862-6|LNC|Hepatitis C virus resistance panel|Hepatitis C virus resistance panel
C3655062|T201|COMP|72861-8|LNC|Ganciclovir|Ganciclovir
C3655063|T201|COMP|72860-0|LNC|Telaprevir|Telaprevir
C3655064|T201|COMP|72859-2|LNC|Boceprevir|Boceprevir
C3655065|T201|COMP|72858-4|LNC|Enfuvirtide|Enfuvirtide
C3655066|T201|COMP|72857-6|LNC|Dolutegravir|Dolutegravir
C3655067|T201|COMP|72856-8|LNC|Cidofovir|Cidofovir
C3655068|T201|COMP|72855-0|LNC|Cidofovir|Cidofovir
C3655069|T201|COMP|72854-3|LNC|Ganciclovir|Ganciclovir
C3655070|T201|COMP|72853-5|LNC|Maribavir|Maribavir
C3655071|T201|COMP|72852-7|LNC|Cytomegalovirus resistance panel|Cytomegalovirus resistance panel
C3655072|T201|COMP|72851-9|LNC|Hepatitis B virus codon 84|Hepatitis B virus codon 84
C3655073|T201|COMP|72850-1|LNC|Hepatitis B virus codon 85|Hepatitis B virus codon 85
C3655074|T201|COMP|72849-3|LNC|Hepatitis B virus codon 169|Hepatitis B virus codon 169
C3655075|T201|COMP|72848-5|LNC|Hepatitis B virus codon 184|Hepatitis B virus codon 184
C3655076|T201|COMP|72847-7|LNC|Hepatitis B virus codon 191|Hepatitis B virus codon 191
C3655077|T201|COMP|72846-9|LNC|Hepatitis B virus codon 194|Hepatitis B virus codon 194
C3655078|T201|COMP|72845-1|LNC|Hepatitis B virus codon 202|Hepatitis B virus codon 202
C3655079|T201|COMP|72844-4|LNC|Hepatitis B virus codon 214|Hepatitis B virus codon 214
C3655080|T201|COMP|72833-7|LNC|Cytomegalovirus UL97 gene mutations detected|Cytomegalovirus UL97 gene mutations detected
C3655084|T201|COMP|73669-4|LNC|Bacteria producing DNAse|Bacteria producing DNAse
C3655085|T201|COMP|73668-6|LNC|Bacteria soluble by bile|Bacteria soluble by bile
C3655086|T201|COMP|73667-8|LNC|Bacteria producing hippuricase|Bacteria producing hippuricase
C3655087|T201|COMP|73666-0|LNC|Streptococcus.beta-hemolytic|Streptococcus.beta-hemolytic
C3655088|T201|COMP|73665-2|LNC|Optochin|Optochin
C3655089|T201|COMP|73370-9|LNC|Fosinopril induced platelet Ab.IgM|Fosinopril induced platelet Ab.IgM
C3655090|T201|COMP|73369-1|LNC|Furosemide induced platelet Ab.IgG|Furosemide induced platelet Ab.IgG
C3655091|T201|COMP|73368-3|LNC|Furosemide induced platelet Ab.IgM|Furosemide induced platelet Ab.IgM
C3655092|T201|COMP|73367-5|LNC|Gabapentin induced platelet Ab.IgG|Gabapentin induced platelet Ab.IgG
C3655093|T201|COMP|73366-7|LNC|Gabapentin induced platelet Ab.IgM|Gabapentin induced platelet Ab.IgM
C3655094|T201|COMP|73300-6|LNC|Lisinopril induced platelet Ab.IgM|Lisinopril induced platelet Ab.IgM
C3655095|T201|COMP|73299-0|LNC|Loperamide induced platelet Ab.IgG|Loperamide induced platelet Ab.IgG
C3655096|T201|COMP|73298-2|LNC|Loperamide induced platelet Ab.IgM|Loperamide induced platelet Ab.IgM
C3655097|T201|COMP|72930-1|LNC|Warfarin induced neutrophil Ab.IgG|Warfarin induced neutrophil Ab.IgG
C3655098|T201|COMP|72929-3|LNC|Warfarin induced neutrophil Ab.IgM|Warfarin induced neutrophil Ab.IgM
C3655099|T201|COMP|72928-5|LNC|Secobarbital|Secobarbital
C3655100|T201|COMP|72927-7|LNC|Urea|Urea
C3655101|T201|COMP|72926-9|LNC|Urea|Urea
C3655102|T201|COMP|72925-1|LNC|Bilirubin|Bilirubin
C3655103|T201|COMP|72924-4|LNC|Barium|Barium
C3655104|T201|COMP|72923-6|LNC|Specimen source|Specimen source
C3655105|T201|COMP|72921-0|LNC|HNA 1 genotype|HNA 1 genotype
C3655106|T201|COMP|72920-2|LNC|HNA 1c genotype|HNA 1c genotype
C3655107|T201|COMP|72919-4|LNC|HNA 3 genotype|HNA 3 genotype
C3655108|T201|COMP|72918-6|LNC|HNA 4 genotype|HNA 4 genotype
C3655109|T201|COMP|72479-9|LNC|Drugs of abuse panel|Drugs of abuse panel
C3655110|T201|COMP|72476-5|LNC|Methadone panel|Methadone panel
C3655111|T201|COMP|73323-8|LNC|ISOtretinoin induced platelet Ab.IgG|ISOtretinoin induced platelet Ab.IgG
C3655112|T201|COMP|73322-0|LNC|ISOtretinoin induced platelet Ab.IgM|ISOtretinoin induced platelet Ab.IgM
C3655113|T201|COMP|73321-2|LNC|Ketorolac induced platelet Ab.IgG|Ketorolac induced platelet Ab.IgG
C3655114|T201|COMP|73320-4|LNC|Ketorolac induced platelet Ab.IgM|Ketorolac induced platelet Ab.IgM
C3655115|T201|COMP|73023-4|LNC|Fenofibrate induced neutrophil Ab.IgM|Fenofibrate induced neutrophil Ab.IgM
C3655116|T201|COMP|73022-6|LNC|Fexofenadine induced neutrophil Ab.IgG|Fexofenadine induced neutrophil Ab.IgG
C3655117|T201|COMP|73021-8|LNC|Fexofenadine induced neutrophil Ab.IgM|Fexofenadine induced neutrophil Ab.IgM
C3655118|T201|COMP|73020-0|LNC|Fluconazole induced neutrophil Ab.IgG|Fluconazole induced neutrophil Ab.IgG
C3655119|T201|COMP|72934-3|LNC|Vancomycin induced neutrophil Ab.IgG|Vancomycin induced neutrophil Ab.IgG
C3655120|T201|COMP|72933-5|LNC|Vancomycin induced neutrophil Ab.IgM|Vancomycin induced neutrophil Ab.IgM
C3655121|T201|COMP|72932-7|LNC|Venlafaxine induced neutrophil Ab.IgG|Venlafaxine induced neutrophil Ab.IgG
C3655122|T201|COMP|72931-9|LNC|Venlafaxine induced neutrophil Ab.IgM|Venlafaxine induced neutrophil Ab.IgM
C3655123|T201|COMP|72838-6|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C3655124|T201|COMP|72837-8|LNC|Bacterial vancomycin resistance vanC1 gene|Bacterial vancomycin resistance vanC1 gene
C3655125|T201|COMP|72836-0|LNC|Bacterial vancomycin resistance vanC2+vanC3 genes|Bacterial vancomycin resistance vanC2+vanC3 genes
C3655126|T201|COMP|72835-2|LNC|Raltegravir|Raltegravir
C3655127|T201|COMP|72834-5|LNC|Foscarnet|Foscarnet
C3655128|T201|COMP|73510-0|LNC|Azithromycin induced platelet Ab.IgM|Azithromycin induced platelet Ab.IgM
C3655129|T201|COMP|73509-2|LNC|Aztreonam induced platelet Ab.IgG|Aztreonam induced platelet Ab.IgG
C3655130|T201|COMP|73508-4|LNC|Aztreonam induced platelet Ab.IgM|Aztreonam induced platelet Ab.IgM
C3655131|T201|COMP|73507-6|LNC|Benazepril induced platelet Ab.IgM|Benazepril induced platelet Ab.IgM
C3655132|T201|COMP|73458-2|LNC|Cephalexin induced platelet Ab.IgG|Cephalexin induced platelet Ab.IgG
C3655133|T201|COMP|73457-4|LNC|chlordiazePOXIDE induced platelet Ab.IgG|chlordiazePOXIDE induced platelet Ab.IgG
C3655134|T201|COMP|73456-6|LNC|chlordiazePOXIDE induced platelet Ab.IgM|chlordiazePOXIDE induced platelet Ab.IgM
C3655135|T201|COMP|73455-8|LNC|chlorproMAZINE induced platelet Ab.IgM|chlorproMAZINE induced platelet Ab.IgM
C3655136|T201|COMP|73454-1|LNC|chlorproMAZINE induced platelet Ab.IgG|chlorproMAZINE induced platelet Ab.IgG
C3655137|T201|COMP|73389-9|LNC|Ezetimibe induced platelet Ab.IgG|Ezetimibe induced platelet Ab.IgG
C3655138|T201|COMP|73388-1|LNC|Ezetimibe induced platelet Ab.IgM|Ezetimibe induced platelet Ab.IgM
C3655139|T201|COMP|73387-3|LNC|Famotidine induced platelet Ab.IgG|Famotidine induced platelet Ab.IgG
C3655140|T201|COMP|73386-5|LNC|Famotidine induced platelet Ab.IgM|Famotidine induced platelet Ab.IgM
C3655141|T201|COMP|73385-7|LNC|Fenofibrate induced platelet Ab.IgG|Fenofibrate induced platelet Ab.IgG
C3655142|T201|COMP|73096-0|LNC|valACYclovir induced platelet Ab.IgG|valACYclovir induced platelet Ab.IgG
C3655143|T201|COMP|73095-2|LNC|Valdecoxib induced platelet Ab.IgM|Valdecoxib induced platelet Ab.IgM
C3655144|T201|COMP|73094-5|LNC|Valdecoxib induced platelet Ab.IgG|Valdecoxib induced platelet Ab.IgG
C3655145|T201|COMP|73093-7|LNC|valGANciclovir induced platelet Ab.IgG|valGANciclovir induced platelet Ab.IgG
C3655146|T201|COMP|73092-9|LNC|valGANciclovir induced platelet Ab.IgM|valGANciclovir induced platelet Ab.IgM
C3655147|T201|COMP|73019-2|LNC|Fluconazole induced neutrophil Ab.IgM|Fluconazole induced neutrophil Ab.IgM
C3655148|T201|COMP|73018-4|LNC|Furosemide induced neutrophil Ab.IgG|Furosemide induced neutrophil Ab.IgG
C3655149|T201|COMP|73017-6|LNC|Furosemide induced neutrophil Ab.IgM|Furosemide induced neutrophil Ab.IgM
C3655150|T201|COMP|73016-8|LNC|Gabapentin induced neutrophil Ab.IgG|Gabapentin induced neutrophil Ab.IgG
C3655151|T201|COMP|72843-6|LNC|Hepatitis B virus codon 215|Hepatitis B virus codon 215
C3655152|T201|COMP|72842-8|LNC|Hepatitis B virus codon 233|Hepatitis B virus codon 233
C3655153|T201|COMP|72841-0|LNC|Hepatitis B virus codon 237|Hepatitis B virus codon 237
C3655154|T201|COMP|72840-2|LNC|Hepatitis B virus codon 250|Hepatitis B virus codon 250
C3655155|T201|COMP|72839-4|LNC|Famciclovir|Famciclovir
C3655156|T201|COMP|73423-6|LNC|diazePAM induced platelet Ab.IgG|diazePAM induced platelet Ab.IgG
C3655157|T201|COMP|73422-8|LNC|diazePAM induced platelet Ab.IgM|diazePAM induced platelet Ab.IgM
C3655158|T201|COMP|73421-0|LNC|Dicyclomine induced platelet Ab.IgG|Dicyclomine induced platelet Ab.IgG
C3655159|T201|COMP|73420-2|LNC|Dicyclomine induced platelet Ab.IgM|Dicyclomine induced platelet Ab.IgM
C3655160|T201|COMP|73419-4|LNC|Digoxin induced platelet Ab.IgM|Digoxin induced platelet Ab.IgM
C3655161|T201|COMP|73418-6|LNC|Digoxin induced platelet Ab.IgG|Digoxin induced platelet Ab.IgG
C3655162|T201|COMP|73417-8|LNC|dilTIAZem induced platelet Ab.IgM|dilTIAZem induced platelet Ab.IgM
C3655163|T201|COMP|73241-2|LNC|Nitroglycerin induced platelet Ab.IgG|Nitroglycerin induced platelet Ab.IgG
C3655164|T201|COMP|73240-4|LNC|Nitroglycerin induced platelet Ab.IgM|Nitroglycerin induced platelet Ab.IgM
C3655165|T201|COMP|73239-6|LNC|Nizatidine induced platelet Ab.IgG|Nizatidine induced platelet Ab.IgG
C3655166|T201|COMP|73238-8|LNC|Nizatidine induced platelet Ab.IgM|Nizatidine induced platelet Ab.IgM
C3655167|T201|COMP|73237-0|LNC|Nystatin induced platelet Ab.IgG|Nystatin induced platelet Ab.IgG
C3655168|T201|COMP|73236-2|LNC|Nystatin induced platelet Ab.IgM|Nystatin induced platelet Ab.IgM
C3655169|T201|COMP|72970-7|LNC|Piperacillin induced neutrophil Ab.IgG|Piperacillin induced neutrophil Ab.IgG
C3655170|T201|COMP|72969-9|LNC|Piperacillin induced neutrophil Ab.IgM|Piperacillin induced neutrophil Ab.IgM
C3655171|T201|COMP|72968-1|LNC|QUEtiapine induced neutrophil Ab.IgG|QUEtiapine induced neutrophil Ab.IgG
C3655172|T201|COMP|72967-3|LNC|QUEtiapine induced neutrophil Ab.IgM|QUEtiapine induced neutrophil Ab.IgM
C3655173|T201|COMP|72966-5|LNC|quiNIDine induced neutrophil Ab.IgG|quiNIDine induced neutrophil Ab.IgG
C3655174|T201|COMP|72965-7|LNC|quiNIDine induced neutrophil Ab.IgM|quiNIDine induced neutrophil Ab.IgM
C3655175|T201|COMP|73297-4|LNC|Loratadine induced platelet Ab.IgG|Loratadine induced platelet Ab.IgG
C3655176|T201|COMP|73296-6|LNC|Loratadine induced platelet Ab.IgM|Loratadine induced platelet Ab.IgM
C3655177|T201|COMP|73011-9|LNC|hydroCHLOROthiazide induced neutrophil Ab.IgM|hydroCHLOROthiazide induced neutrophil Ab.IgM
C3655178|T201|COMP|73010-1|LNC|Ibuprofen induced neutrophil Ab.IgG|Ibuprofen induced neutrophil Ab.IgG
C3655179|T201|COMP|73009-3|LNC|Ibuprofen induced neutrophil Ab.IgM|Ibuprofen induced neutrophil Ab.IgM
C3655180|T201|COMP|73008-5|LNC|Lansoprazole induced neutrophil Ab.IgG|Lansoprazole induced neutrophil Ab.IgG
C3655181|T201|COMP|73007-7|LNC|Lansoprazole induced neutrophil Ab.IgM|Lansoprazole induced neutrophil Ab.IgM
C3655182|T201|COMP|70148-2|LNC|Methadone|Methadone
C3655183|T201|COMP|70147-4|LNC|Methadone|Methadone
C3655184|T201|COMP|70146-6|LNC|Benzoylecgonine|Benzoylecgonine
C3655185|T201|COMP|70145-8|LNC|Cannabinoids|Cannabinoids
C3655186|T201|COMP|70151-6|LNC|Opiates|Opiates
C3655187|T201|COMP|70150-8|LNC|Opiates|Opiates
C3655188|T201|COMP|70137-5|LNC|Sample icteric|Sample icteric
C3655189|T201|COMP|70153-2|LNC|Sample hemolyzed|Sample hemolyzed
C3655190|T201|COMP|70152-4|LNC|Triiodothyronine/Thyroxine|Triiodothyronine/Thyroxine
C3655191|T201|COMP|66951-5|LNC|Complement C1.functional|Complement C1.functional
C3665475|T201|COMP|74239-5|LNC|HEDIS 2014 Value Set - carBAMazepine Level|HEDIS 2014 Value Set - carBAMazepine Level
C3665673|T201|COMP|74245-2|LNC|HEDIS 2014-2016 Value Set - Group A Strep Tests|HEDIS 2014-2016 Value Set - Group A Strep Tests
C3668843|T201|COMP|74243-7|LNC|HEDIS 2014-2016 Value Set - FOBT|HEDIS 2014-2016 Value Set - FOBT
C3668845|T201|COMP|74250-2|LNC|HEDIS 2014, 2015 Value Set - Lead Tests|HEDIS 2014, 2015 Value Set - Lead Tests
C3668847|T201|COMP|74258-5|LNC|HEDIS 2014 Value Set - Sexual Activity|HEDIS 2014 Value Set - Sexual Activity
C3668994|T201|COMP|74261-9|LNC|HEDIS 2014 Value Set - Phenytoin Level|HEDIS 2014 Value Set - Phenytoin Level
C3668995|T201|COMP|74253-6|LNC|HEDIS 2014 Value Set - Pregnancy Tests|HEDIS 2014 Value Set - Pregnancy Tests
C3668997|T201|COMP|74254-4|LNC|HEDIS 2014-2018 Value Set - Rh|HEDIS 2014-2018 Value Set - Rh
C3669003|T201|COMP|74255-1|LNC|HEDIS 2014-2018 Value Set - Rubella Antibody|HEDIS 2014-2018 Value Set - Rubella Antibody
C3669004|T201|COMP|74256-9|LNC|HEDIS 2014-2019 Value Set - Serum Creatinine|HEDIS 2014-2019 Value Set - Serum Creatinine
C3669006|T201|COMP|74252-8|LNC|HEDIS 2014 Value Set - PHENobarbital Level|HEDIS 2014 Value Set - PHENobarbital Level
C3669007|T201|COMP|74257-7|LNC|HEDIS 2014-2016 Value Set - Serum Potassium|HEDIS 2014-2016 Value Set - Serum Potassium
C3669142|T201|COMP|74240-3|LNC|HEDIS 2014-2020 Value Set - Cervical Cytology|HEDIS 2014-2020 Value Set - Cervical Cytology
C3669146|T201|COMP|74262-7|LNC|HEDIS 2014-2018 Value Set - Toxoplasma Antibody|HEDIS 2014-2018 Value Set - Toxoplasma Antibody
C3669187|T201|COMP|74235-3|LNC|HEDIS 2014-2019 Value Set - ABO|HEDIS 2014-2019 Value Set - ABO
C3669192|T201|COMP|74260-1|LNC|HEDIS 2014 Value Set - Valproic Acid Level|HEDIS 2014 Value Set - Valproic Acid Level
C3669194|T201|COMP|74234-6|LNC|HEDIS 2014 Value Sets|HEDIS 2014 Value Sets
C3669302|T201|COMP|74397-1|LNC|Reticulocytes/100 erythrocytes|Reticulocytes/100 erythrocytes
C3669323|T201|COMP|74237-9|LNC|HEDIS 2014, 2015 Value Set - ABO and Rh|HEDIS 2014, 2015 Value Set - ABO and Rh
C3669325|T201|COMP|74238-7|LNC|HEDIS 2014 Value Set - Blood Urea Nitrogen|HEDIS 2014 Value Set - Blood Urea Nitrogen
C3669326|T201|COMP|74241-1|LNC|HEDIS 2014-2016 Value Set - Chlamydia Tests|HEDIS 2014-2016 Value Set - Chlamydia Tests
C3669331|T201|COMP|74244-5|LNC|HEDIS 2014 Value Set - Glucose Tests|HEDIS 2014 Value Set - Glucose Tests
C3669334|T201|COMP|74246-0|LNC|HEDIS 2014 Value Set - HbA1c Tests|HEDIS 2014 Value Set - HbA1c Tests
C3669338|T201|COMP|74249-4|LNC|HEDIS 2014 Value Set - LDL-C Tests|HEDIS 2014 Value Set - LDL-C Tests
C3671182|T201|COMP|74411-0|LNC|Consistency|Consistency
C3699321|T201|COMP|74138-9|LNC|Monocytes.immature|Monocytes.immature
C3699322|T201|COMP|74139-7|LNC|Mononuclear cells|Mononuclear cells
C3699323|T201|COMP|74140-5|LNC|Granulocytes|Granulocytes
C3699324|T201|COMP|74141-3|LNC|Granulocytes/100 leukocytes|Granulocytes/100 leukocytes
C3699325|T201|COMP|74142-1|LNC|Granulocytes|Granulocytes
C3699326|T201|COMP|74143-9|LNC|Granulocytes/100 leukocytes|Granulocytes/100 leukocytes
C3699327|T201|COMP|74032-4|LNC|Arbovirus Ab.IgM panel|Arbovirus Ab.IgM panel
C3699329|T201|COMP|74033-2|LNC|Arbovirus Ab.IgM|Arbovirus Ab.IgM
C3699330|T201|COMP|74034-0|LNC|MAML2 11q21 gene rearrangements|MAML2 11q21 gene rearrangements
C3699332|T201|COMP|74035-7|LNC|Prion protein.abnormal|Prion protein.abnormal
C3699333|T201|COMP|74036-5|LNC|Prion protein.abnormal|Prion protein.abnormal
C3699334|T201|COMP|74112-4|LNC|Bromadiolone|Bromadiolone
C3699335|T201|COMP|74113-2|LNC|Coumafuryl|Coumafuryl
C3699336|T201|COMP|74114-0|LNC|Coumatetralyl|Coumatetralyl
C3699337|T201|COMP|74115-7|LNC|Difenacoum|Difenacoum
C3699338|T201|COMP|74116-5|LNC|Adalimumab Ab|Adalimumab Ab
C3699342|T201|COMP|73982-1|LNC|Bacterial carbapenem resistance blaNDM gene|Bacterial carbapenem resistance blaNDM gene
C3699346|T201|COMP|73984-7|LNC|Hemoglobin.other|Hemoglobin.other
C3699347|T201|COMP|73987-0|LNC|2,2',3,4,4',5-Hexachlorobiphenyl|2,2',3,4,4',5-Hexachlorobiphenyl
C3699349|T201|COMP|73988-8|LNC|2,2',4,5,5'-Pentachlorobiphenyl|2,2',4,5,5'-Pentachlorobiphenyl
C3699350|T201|COMP|73989-6|LNC|2,3',4,4',5-Pentachlorobiphenyl|2,3',4,4',5-Pentachlorobiphenyl
C3699351|T201|COMP|73990-4|LNC|2,3',4',5-Tetrachlorobiphenyl|2,3',4',5-Tetrachlorobiphenyl
C3699353|T201|COMP|73991-2|LNC|2,2',5,5'-Tetrachlorobiphenyl|2,2',5,5'-Tetrachlorobiphenyl
C3699354|T201|COMP|73992-0|LNC|2,2',5-Trichlorobiphenyl|2,2',5-Trichlorobiphenyl
C3699355|T201|COMP|73993-8|LNC|Polychlorinated biphenyl|Polychlorinated biphenyl
C3699356|T201|COMP|73994-6|LNC|Polychlorinated biphenyl|Polychlorinated biphenyl
C3699357|T201|COMP|73995-3|LNC|Mitragynine|Mitragynine
C3699358|T201|COMP|73996-1|LNC|oxyCODONE|oxyCODONE
C3699359|T201|COMP|73997-9|LNC|Ibuprofen|Ibuprofen
C3699360|T201|COMP|73998-7|LNC|25H-NBOMe|25H-NBOMe
C3699362|T201|COMP|73999-5|LNC|2C-C-NBOMe|2C-C-NBOMe
C3699364|T201|COMP|74000-1|LNC|25I-NBOMe|25I-NBOMe
C3699366|T201|COMP|74001-9|LNC|NBOMe|NBOMe
C3699368|T201|COMP|74002-7|LNC|Tungsten/Creatinine|Tungsten/Creatinine
C3699370|T201|COMP|74003-5|LNC|CYP3A4 gene.c.-392A>G (*1B)|CYP3A4 gene.c.-392A>G (*1B)
C3699372|T201|COMP|74004-3|LNC|ABCB1 gene targeted mutation analysis|ABCB1 gene targeted mutation analysis
C3699378|T201|COMP|74007-6|LNC|CYP3A4 gene targeted mutation analysis|CYP3A4 gene targeted mutation analysis
C3699391|T201|COMP|74031-6|LNC|Arbovirus identified|Arbovirus identified
C3699392|T201|COMP|74037-3|LNC|Transmissible spongiform encephalopathy|Transmissible spongiform encephalopathy
C3699393|T201|COMP|74038-1|LNC|Influenza virus A H1 RNA|Influenza virus A H1 RNA
C3699394|T201|COMP|74039-9|LNC|Influenza virus A H3 RNA|Influenza virus A H3 RNA
C3699395|T201|COMP|74040-7|LNC|Influenza virus A N2 RNA|Influenza virus A N2 RNA
C3699461|T201|COMP|74082-9|LNC|Urea|Urea
C3699462|T201|COMP|74083-7|LNC|Norolanzapine|Norolanzapine
C3699463|T201|COMP|74084-5|LNC|Glucose^15M post 50 g lactose PO|Glucose^15M post 50 g lactose PO
C3699464|T201|COMP|74085-2|LNC|Isocoproporphyrin|Isocoproporphyrin
C3699465|T201|COMP|74086-0|LNC|Pentacarboxylporphyrin III|Pentacarboxylporphyrin III
C3699466|T201|COMP|74087-8|LNC|Hexacarboxylporphyrin III|Hexacarboxylporphyrin III
C3699467|T201|COMP|74088-6|LNC|Heptacarboxylporphyrin III|Heptacarboxylporphyrin III
C3699468|T201|COMP|74089-4|LNC|Pentacarboxylporphyrin III/Creatinine|Pentacarboxylporphyrin III/Creatinine
C3699470|T201|COMP|74090-2|LNC|Hexacarboxylporphyrin III/Creatinine|Hexacarboxylporphyrin III/Creatinine
C3699472|T201|COMP|74091-0|LNC|Heptacarboxylporphyrin III/Creatinine|Heptacarboxylporphyrin III/Creatinine
C3699474|T201|COMP|74092-8|LNC|Acidity.titratable|Acidity.titratable
C3699475|T201|COMP|74093-6|LNC|Gliquidone|Gliquidone
C3699476|T201|COMP|74094-4|LNC|Gliclazide|Gliclazide
C3699477|T201|COMP|74095-1|LNC|Didesmethylcitalopram|Didesmethylcitalopram
C3699478|T201|COMP|74096-9|LNC|Tacrolimus|Tacrolimus
C3699479|T201|COMP|74097-7|LNC|Tacrolimus|Tacrolimus
C3699480|T201|COMP|74098-5|LNC|Endothelin|Endothelin
C3699481|T201|COMP|74099-3|LNC|Neutrophil gelatinase-associated lipocalin|Neutrophil gelatinase-associated lipocalin
C3699482|T201|COMP|74100-9|LNC|Nitrate+Nitrite|Nitrate+Nitrite
C3699483|T201|COMP|74101-7|LNC|Tissue inhibitor of metalloproteinases 1|Tissue inhibitor of metalloproteinases 1
C3699484|T201|COMP|74102-5|LNC|Matrix metallopeptidase 2|Matrix metallopeptidase 2
C3699486|T201|COMP|74103-3|LNC|Neutrophil gelatinase-associated lipocalin|Neutrophil gelatinase-associated lipocalin
C3699487|T201|COMP|74104-1|LNC|Alpha-amanitin+gamma-amanitin|Alpha-amanitin+gamma-amanitin
C3699489|T201|COMP|74105-8|LNC|Oxygen saturation|Oxygen saturation
C3699490|T201|COMP|74106-6|LNC|Proteinase 3 Ab.IgG|Proteinase 3 Ab.IgG
C3699491|T201|COMP|74107-4|LNC|Warfarin|Warfarin
C3699492|T201|COMP|74108-2|LNC|Meperidine|Meperidine
C3699493|T201|COMP|74109-0|LNC|4-hydroxycoumarins|4-hydroxycoumarins
C3699494|T201|COMP|74110-8|LNC|traMADol|traMADol
C3699495|T201|COMP|74111-6|LNC|Brodifacoum|Brodifacoum
C3699496|T201|COMP|74117-3|LNC|Adalimumab|Adalimumab
C3699497|T201|COMP|74118-1|LNC|P27 Ag|P27 Ag
C3699498|T201|COMP|74119-9|LNC|P504S Ag|P504S Ag
C3699500|T201|COMP|74120-7|LNC|PDGFR-alpha Ag|PDGFR-alpha Ag
C3699502|T201|COMP|74121-5|LNC|Perforin Ag|Perforin Ag
C3699504|T201|COMP|74122-3|LNC|Ubiquitin Ag|Ubiquitin Ag
C3699506|T201|COMP|74123-1|LNC|Phospho-S6 ribosomal protein Ag|Phospho-S6 ribosomal protein Ag
C3699508|T201|COMP|74124-9|LNC|Blood group 8 Ag|Blood group 8 Ag
C3699510|T201|COMP|74125-6|LNC|Mesothelin Ag|Mesothelin Ag
C3699512|T201|COMP|74126-4|LNC|Mucin-4 Ag|Mucin-4 Ag
C3699514|T201|COMP|74127-2|LNC|Akt1 phosphate Ag|Akt1 phosphate Ag
C3699516|T201|COMP|74128-0|LNC|Neuroblastoma 84 Ag|Neuroblastoma 84 Ag
C3699518|T201|COMP|74129-8|LNC|Transforming growth factor alpha Ag|Transforming growth factor alpha Ag
C3699520|T201|COMP|74130-6|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C3699521|T201|COMP|74131-4|LNC|Morphine|Morphine
C3699522|T201|COMP|74132-2|LNC|Aromatic solvents|Aromatic solvents
C3699523|T201|COMP|74133-0|LNC|Volatiles|Volatiles
C3699524|T201|COMP|74134-8|LNC|Ezogabine|Ezogabine
C3699525|T201|COMP|74135-5|LNC|N-acetyl ezogabine|N-acetyl ezogabine
C3699527|T201|COMP|74136-3|LNC|fentaNYL|fentaNYL
C3699528|T201|COMP|74137-1|LNC|Norfentanyl|Norfentanyl
C3699529|T201|COMP|74337-7|LNC|MICA*012 Ab.IgG|MICA*012 Ab.IgG
C3699531|T201|COMP|74338-5|LNC|MICA*011 Ab.IgG|MICA*011 Ab.IgG
C3699533|T201|COMP|74339-3|LNC|MICA*009 Ab.IgG|MICA*009 Ab.IgG
C3699535|T201|COMP|74340-1|LNC|MICA*008 Ab.IgG|MICA*008 Ab.IgG
C3699537|T201|COMP|74341-9|LNC|MICA*007 Ab.IgG|MICA*007 Ab.IgG
C3699539|T201|COMP|74418-5|LNC|Measles virus Ab.IgG|Measles virus Ab.IgG
C3699540|T201|COMP|74419-3|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C3699541|T201|COMP|74420-1|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C3699542|T201|COMP|74421-9|LNC|Mumps virus Ab.IgM|Mumps virus Ab.IgM
C3699545|T201|COMP|74157-9|LNC|Cannabinoids|Cannabinoids
C3699555|T201|COMP|74167-8|LNC|Opiates|Opiates
C3699556|T201|COMP|74168-6|LNC|Barbiturates|Barbiturates
C3699557|T201|COMP|74169-4|LNC|Cocaine|Cocaine
C3699558|T201|COMP|74170-2|LNC|Ceftaroline|Ceftaroline
C3699585|T201|COMP|74184-3|LNC|Lymphocytes.clefted|Lymphocytes.clefted
C3699629|T201|COMP|74469-8|LNC|Glucose-6-Phosphate dehydrogenase/Pyruvate kinase|Glucose-6-Phosphate dehydrogenase/Pyruvate kinase
C3699643|T201|COMP|74214-8|LNC|Apixaban|Apixaban
C3699644|T201|COMP|74215-5|LNC|Rivaroxaban|Rivaroxaban
C3699645|T201|COMP|74216-3|LNC|Fondaparinux|Fondaparinux
C3699646|T201|COMP|74217-1|LNC|Fondaparinux|Fondaparinux
C3699647|T201|COMP|74218-9|LNC|Apixaban|Apixaban
C3699650|T201|COMP|74220-5|LNC|Dabigatran|Dabigatran
C3699651|T201|COMP|74222-1|LNC|Reviewed material & summary of stains|Reviewed material & summary of stains
C3699653|T201|COMP|74223-9|LNC|Immunohistochemical stains|Immunohistochemical stains
C3699654|T201|COMP|74224-7|LNC|Disease category|Disease category
C3699656|T201|COMP|74225-4|LNC|Cytochemical stains|Cytochemical stains
C3699658|T201|COMP|74226-2|LNC|Plasma cells assessment|Plasma cells assessment
C3699660|T201|COMP|74227-0|LNC|Other observations|Other observations
C3699662|T201|COMP|74228-8|LNC|Myelopoiesis assessment|Myelopoiesis assessment
C3699664|T201|COMP|74229-6|LNC|Megakaryopoiesis assessment|Megakaryopoiesis assessment
C3699666|T201|COMP|74230-4|LNC|Lymphocytes assessment|Lymphocytes assessment
C3699668|T201|COMP|74231-2|LNC|Erythropoiesis assessment|Erythropoiesis assessment
C3699670|T201|COMP|74232-0|LNC|Cellularity assessment|Cellularity assessment
C3699671|T201|COMP|74233-8|LNC|Blasts assessment|Blasts assessment
C3699673|T201|COMP|74236-1|LNC|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C3699674|T201|COMP|74263-5|LNC|Dabigatran|Dabigatran
C3699681|T201|COMP|74279-1|LNC|Gamma interferon.negative control spot count|Gamma interferon.negative control spot count
C3699704|T201|COMP|74294-0|LNC|Isovaleric acidemia|Isovaleric acidemia
C3699705|T201|COMP|74295-7|LNC|Hydroxymethylglutaryl CoA lyase deficiency|Hydroxymethylglutaryl CoA lyase deficiency
C3699706|T201|COMP|74296-5|LNC|3-Methylcrotonyl-CoA carboxylase deficiency|3-Methylcrotonyl-CoA carboxylase deficiency
C3699707|T201|COMP|74297-3|LNC|Isobutyryl-CoA dehydrogenase deficiency|Isobutyryl-CoA dehydrogenase deficiency
C3699708|T201|COMP|74298-1|LNC|Short-chain acyl-CoA dehydrogenase deficiency|Short-chain acyl-CoA dehydrogenase deficiency
C3699709|T201|COMP|74299-9|LNC|Tyrosine/Phenylalanine^post therapeutic diet|Tyrosine/Phenylalanine^post therapeutic diet
C3699711|T201|COMP|74300-5|LNC|Phenylalanine/Tyrosine^post therapeutic diet|Phenylalanine/Tyrosine^post therapeutic diet
C3699712|T201|COMP|74301-3|LNC|Succinylacetone^post therapeutic diet|Succinylacetone^post therapeutic diet
C3699713|T201|COMP|74302-1|LNC|Tyrosine^post therapeutic diet|Tyrosine^post therapeutic diet
C3699714|T201|COMP|74303-9|LNC|Phenylalanine^post therapeutic diet|Phenylalanine^post therapeutic diet
C3699740|T201|COMP|74319-5|LNC|MICA*051 Ab.IgG|MICA*051 Ab.IgG
C3699742|T201|COMP|74320-3|LNC|MICA*050 Ab.IgG|MICA*050 Ab.IgG
C3699744|T201|COMP|74321-1|LNC|MICA*046 Ab.IgG|MICA*046 Ab.IgG
C3699746|T201|COMP|74322-9|LNC|MICA*043 Ab.IgG|MICA*043 Ab.IgG
C3699748|T201|COMP|74323-7|LNC|MICA*042 Ab.IgG|MICA*042 Ab.IgG
C3699750|T201|COMP|74324-5|LNC|MICA*041 Ab.IgG|MICA*041 Ab.IgG
C3699752|T201|COMP|74325-2|LNC|MICA*037 Ab.IgG|MICA*037 Ab.IgG
C3699754|T201|COMP|74326-0|LNC|MICA*036 Ab.IgG|MICA*036 Ab.IgG
C3699756|T201|COMP|74327-8|LNC|MICA*033 Ab.IgG|MICA*033 Ab.IgG
C3699758|T201|COMP|74328-6|LNC|MICA*030 Ab.IgG|MICA*030 Ab.IgG
C3699760|T201|COMP|74329-4|LNC|MICA*029 Ab.IgG|MICA*029 Ab.IgG
C3699762|T201|COMP|74330-2|LNC|MICA*028 Ab.IgG|MICA*028 Ab.IgG
C3699764|T201|COMP|74331-0|LNC|MICA*024 Ab.IgG|MICA*024 Ab.IgG
C3699766|T201|COMP|74332-8|LNC|MICA*019 Ab.IgG|MICA*019 Ab.IgG
C3699768|T201|COMP|74333-6|LNC|MICA*018 Ab.IgG|MICA*018 Ab.IgG
C3699770|T201|COMP|74334-4|LNC|MICA*017 Ab.IgG|MICA*017 Ab.IgG
C3699772|T201|COMP|74335-1|LNC|MICA*016 Ab.IgG|MICA*016 Ab.IgG
C3699774|T201|COMP|74336-9|LNC|MICA*015 Ab.IgG|MICA*015 Ab.IgG
C3699776|T201|COMP|74342-7|LNC|MICA*006 Ab.IgG|MICA*006 Ab.IgG
C3699778|T201|COMP|74343-5|LNC|MICA*005 Ab.IgG|MICA*005 Ab.IgG
C3699780|T201|COMP|74344-3|LNC|MICA*004 Ab.IgG|MICA*004 Ab.IgG
C3699782|T201|COMP|74345-0|LNC|MICA*002 Ab.IgG|MICA*002 Ab.IgG
C3699784|T201|COMP|74346-8|LNC|MICA*001 Ab.IgG|MICA*001 Ab.IgG
C3699786|T201|COMP|74347-6|LNC|Leukocyte aggregates|Leukocyte aggregates
C3699788|T201|COMP|74348-4|LNC|Bacteria identified|Bacteria identified
C3699789|T201|COMP|74349-2|LNC|Lactose^post CFst|Lactose^post CFst
C3699791|T201|COMP|74351-8|LNC|Glucose|Glucose
C3699792|T201|COMP|74352-6|LNC|Cryoglobulin & cryofibrinogen panel|Cryoglobulin & cryofibrinogen panel
C3699794|T201|COMP|74353-4|LNC|Sodium & Potassium panel|Sodium & Potassium panel
C3699795|T201|COMP|74354-2|LNC|Epithelial cells/100 leukocytes|Epithelial cells/100 leukocytes
C3699797|T201|COMP|74355-9|LNC|Bacteria identified|Bacteria identified
C3699798|T201|COMP|74356-7|LNC|Bacteria identified|Bacteria identified
C3699799|T201|COMP|74357-5|LNC|Lymphocytes.immunoblastic|Lymphocytes.immunoblastic
C3699800|T201|COMP|74358-3|LNC|Adenine phosphoribosyltransferase|Adenine phosphoribosyltransferase
C3699801|T201|COMP|74359-1|LNC|Cholesterol ester transfer protein actual/normal|Cholesterol ester transfer protein actual/normal
C3699803|T201|COMP|74360-9|LNC|Cortisone|Cortisone
C3699804|T201|COMP|74361-7|LNC|Dehydroepiandrosterone|Dehydroepiandrosterone
C3699807|T201|COMP|74363-3|LNC|N,N-dimethylarginine|N,N-dimethylarginine
C3699808|T201|COMP|74364-1|LNC|Oxytocin|Oxytocin
C3699809|T201|COMP|74365-8|LNC|Palmitoyl protein thioesterase|Palmitoyl protein thioesterase
C3699810|T201|COMP|74366-6|LNC|Clorazepate^trough|Clorazepate^trough
C3699811|T201|COMP|74367-4|LNC|Norfluoxetine^trough|Norfluoxetine^trough
C3699812|T201|COMP|74368-2|LNC|Apelin|Apelin
C3699813|T201|COMP|74369-0|LNC|Nitric oxide|Nitric oxide
C3699814|T201|COMP|74370-8|LNC|Cotinine|Cotinine
C3699815|T201|COMP|74371-6|LNC|Cotinine|Cotinine
C3699816|T201|COMP|74372-4|LNC|Acetyl fentaNYL|Acetyl fentaNYL
C3699818|T201|COMP|74373-2|LNC|cloNIDine|cloNIDine
C3699819|T201|COMP|74374-0|LNC|2,4,4'-Trichlorobiphenyl|2,4,4'-Trichlorobiphenyl
C3699820|T201|COMP|74375-7|LNC|2,2',3,5'-Tetrachlorobiphenyl|2,2',3,5'-Tetrachlorobiphenyl
C3699822|T201|COMP|74376-5|LNC|2,2',4,4',5,5'-Hexachlorobiphenyl|2,2',4,4',5,5'-Hexachlorobiphenyl
C3699823|T201|COMP|74377-3|LNC|Baclofen|Baclofen
C3699824|T201|COMP|74378-1|LNC|Meperidine|Meperidine
C3699825|T201|COMP|74379-9|LNC|Morphine|Morphine
C3699826|T201|COMP|74380-7|LNC|HYDROmorphone|HYDROmorphone
C3699827|T201|COMP|74381-5|LNC|Midazolam|Midazolam
C3699828|T201|COMP|74382-3|LNC|Bupivacaine|Bupivacaine
C3699829|T201|COMP|74383-1|LNC|fentaNYL|fentaNYL
C3699830|T201|COMP|74384-9|LNC|Specimen container|Specimen container
C3699831|T201|COMP|74385-6|LNC|Normirtazapine|Normirtazapine
C3699832|T201|COMP|74386-4|LNC|Normirtazapine|Normirtazapine
C3699833|T201|COMP|74387-2|LNC|Normirtazapine|Normirtazapine
C3699834|T201|COMP|74388-0|LNC|Normirtazapine|Normirtazapine
C3699835|T201|COMP|74389-8|LNC|Normirtazapine|Normirtazapine
C3699836|T201|COMP|74390-6|LNC|Baclofen|Baclofen
C3699837|T201|COMP|74391-4|LNC|Baclofen|Baclofen
C3699838|T201|COMP|74392-2|LNC|Zopiclone|Zopiclone
C3699839|T201|COMP|74393-0|LNC|Reticulocytes.immature/100 erythrocytes|Reticulocytes.immature/100 erythrocytes
C3699841|T201|COMP|74394-8|LNC|Normoblasts|Normoblasts
C3699842|T201|COMP|74395-5|LNC|Blasts|Blasts
C3699843|T201|COMP|74396-3|LNC|Large unstained cells/100 leukocytes|Large unstained cells/100 leukocytes
C3699844|T201|COMP|74398-9|LNC|Neutrophils|Neutrophils
C3699845|T201|COMP|74399-7|LNC|Monocytes|Monocytes
C3699846|T201|COMP|74400-3|LNC|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C3699847|T201|COMP|74401-1|LNC|Lymphocytes|Lymphocytes
C3699848|T201|COMP|74402-9|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C3699849|T201|COMP|74403-7|LNC|Normoblasts/100 leukocytes|Normoblasts/100 leukocytes
C3699850|T201|COMP|74404-5|LNC|Eosinophils|Eosinophils
C3699851|T201|COMP|74405-2|LNC|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C3699852|T201|COMP|74406-0|LNC|Basophils|Basophils
C3699853|T201|COMP|74407-8|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C3699856|T201|COMP|74409-4|LNC|MICA Ab.IgG panel|MICA Ab.IgG panel
C3699858|T201|COMP|74410-2|LNC|Polychlorinated biphenyl panel|Polychlorinated biphenyl panel
C3699860|T201|COMP|74412-8|LNC|CBC W Differential panel|CBC W Differential panel
C3699862|T201|COMP|74413-6|LNC|Differential panel|Differential panel
C3699863|T201|COMP|74414-4|LNC|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C3699864|T201|COMP|74415-1|LNC|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C3699865|T201|COMP|74416-9|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C3699866|T201|COMP|74417-7|LNC|Measles virus Ab.IgM|Measles virus Ab.IgM
C3699867|T201|COMP|74422-7|LNC|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C3699868|T201|COMP|74423-5|LNC|Enterovirus RNA|Enterovirus RNA
C3699869|T201|COMP|74424-3|LNC|Enterovirus RNA|Enterovirus RNA
C3699870|T201|COMP|74425-0|LNC|Myelocytes.neutrophilic/100 leukocytes|Myelocytes.neutrophilic/100 leukocytes
C3699872|T201|COMP|74426-8|LNC|Myelocytes.neutrophilic/100 cells|Myelocytes.neutrophilic/100 cells
C3699874|T201|COMP|74427-6|LNC|Myelocytes.eosinophilic/100 leukocytes|Myelocytes.eosinophilic/100 leukocytes
C3699876|T201|COMP|74428-4|LNC|Metamyelocytes.neutrophilic/100 leukocytes|Metamyelocytes.neutrophilic/100 leukocytes
C3699878|T201|COMP|74429-2|LNC|Metamyelocytes.eosinophilic/100 cells|Metamyelocytes.eosinophilic/100 cells
C3699880|T201|COMP|74430-0|LNC|3-Hydroxykynurenin|3-Hydroxykynurenin
C3699881|T201|COMP|74431-8|LNC|Acetoacetate|Acetoacetate
C3699882|T201|COMP|74432-6|LNC|Cholestanol|Cholestanol
C3699883|T201|COMP|74433-4|LNC|Cholestanol/Cholesterol|Cholestanol/Cholesterol
C3699885|T201|COMP|74434-2|LNC|Bilirubin/Total|Bilirubin/Total
C3699886|T201|COMP|74435-9|LNC|Cholesterol.non-esterified/Cholesterol.total|Cholesterol.non-esterified/Cholesterol.total
C3699888|T201|COMP|74436-7|LNC|D-lactate|D-lactate
C3699889|T201|COMP|74437-5|LNC|Galactokinase|Galactokinase
C3699890|T201|COMP|74438-3|LNC|Lactose/Creatinine|Lactose/Creatinine
C3699892|T201|COMP|74439-1|LNC|Gamma aminobutyrate free and total panel|Gamma aminobutyrate free and total panel
C3699894|T201|COMP|74440-9|LNC|Pemptoporphyrin|Pemptoporphyrin
C3699896|T201|COMP|74441-7|LNC|Porphobilinogen/Creatinine|Porphobilinogen/Creatinine
C3699897|T201|COMP|74442-5|LNC|Pyridoxal phosphate|Pyridoxal phosphate
C3699898|T201|COMP|74443-3|LNC|Sucrose/Creatinine^post XXX g sugar solution PO|Sucrose/Creatinine^post XXX g sugar solution PO
C3699900|T201|COMP|74444-1|LNC|Thiamine pyrophosphate|Thiamine pyrophosphate
C3699901|T201|COMP|74445-8|LNC|Porphyrin fractions panel|Porphyrin fractions panel
C3699902|T201|COMP|74446-6|LNC|Calculus analysis panel|Calculus analysis panel
C3699904|T201|COMP|74447-4|LNC|Sugars and polyols panel|Sugars and polyols panel
C3699906|T201|COMP|74448-2|LNC|Sugars and polyols pattern|Sugars and polyols pattern
C3699908|T201|COMP|74450-8|LNC|Other cells|Other cells
C3699909|T201|COMP|74451-6|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C3699910|T201|COMP|74452-4|LNC|Platelet distribution width|Platelet distribution width
C3699911|T201|COMP|74453-2|LNC|Histiocytes/100 cells|Histiocytes/100 cells
C3699912|T201|COMP|74454-0|LNC|Normoblasts|Normoblasts
C3699913|T201|COMP|74455-7|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C3699914|T201|COMP|74456-5|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C3699915|T201|COMP|74457-3|LNC|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C3699916|T201|COMP|74458-1|LNC|Large unstained cells/100 leukocytes|Large unstained cells/100 leukocytes
C3699917|T201|COMP|74459-9|LNC|Granulocytes.immature/100 leukocytes|Granulocytes.immature/100 leukocytes
C3699918|T201|COMP|74460-7|LNC|Blasts/100 leukocytes|Blasts/100 leukocytes
C3699919|T201|COMP|74461-5|LNC|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C3699920|T201|COMP|74462-3|LNC|Basophils/100 leukocytes|Basophils/100 leukocytes
C3699921|T201|COMP|74463-1|LNC|Normoblasts/100 leukocytes|Normoblasts/100 leukocytes
C3699922|T201|COMP|74464-9|LNC|Platelets|Platelets
C3699932|T201|COMP|74475-5|LNC|Middle east respiratory syndrome coronavirus RNA|Middle east respiratory syndrome coronavirus RNA
C3699942|T201|COMP|74481-3|LNC|Tyrosine/Phenylalanine|Tyrosine/Phenylalanine
C3699943|T201|COMP|74483-9|LNC|Homocitrulline|Homocitrulline
C3699944|T201|COMP|74484-7|LNC|Argininosuccinate|Argininosuccinate
C3715002|T201|COMP|75091-9|LNC|Catechol/Creatinine|Catechol/Creatinine
C3831801|T201|COMP|74952-3|LNC|Lymphocyte proliferation|Lymphocyte proliferation
C3833389|T201|COMP|74859-0|LNC|Ethanol|Ethanol
C3833418|T201|COMP|74820-2|LNC|Plasma cells.centrocytes/100 leukocytes|Plasma cells.centrocytes/100 leukocytes
C3833429|T201|COMP|74814-5|LNC|Plasma cells.centroblasts/100 leukocytes|Plasma cells.centroblasts/100 leukocytes
C3846734|T201|COMP|74652-9|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C3846736|T201|COMP|75150-3|LNC|Inosine|Inosine
C3846737|T201|COMP|74532-3|LNC|Energy content|Energy content
C3846738|T201|COMP|75095-0|LNC|Docosahexaenoate|Docosahexaenoate
C3846739|T201|COMP|75080-2|LNC|N-acetyl-L-aspartate|N-acetyl-L-aspartate
C3846740|T201|COMP|74492-0|LNC|PAX5 & CD43 Ag|PAX5 & CD43 Ag
C3846741|T201|COMP|74850-9|LNC|Lymphoblasts/100 cells|Lymphoblasts/100 cells
C3846742|T201|COMP|74914-3|LNC|Acylglycines panel|Acylglycines panel
C3846743|T201|COMP|74993-7|LNC|Chloride & sodium panel|Chloride & sodium panel
C3846744|T201|COMP|74970-5|LNC|Acetylsalicylate^trough|Acetylsalicylate^trough
C3846745|T201|COMP|74865-7|LNC|IgA.lambda|IgA.lambda
C3846746|T201|COMP|75269-1|LNC|Bacteria identified|Bacteria identified
C3846747|T201|COMP|75268-3|LNC|Leucine/Phenylalanine|Leucine/Phenylalanine
C3846750|T201|COMP|75265-9|LNC|Blood group antibody screen|Blood group antibody screen
C3846751|T201|COMP|75264-2|LNC|Blood group antibody screen|Blood group antibody screen
C3846752|T201|COMP|75263-4|LNC|Blood group antibody screen|Blood group antibody screen
C3846769|T201|COMP|75242-8|LNC|Antipsychotics|Antipsychotics
C3846770|T201|COMP|75241-0|LNC|Procalcitonin|Procalcitonin
C3846771|T201|COMP|75240-2|LNC|Meat fibers|Meat fibers
C3846772|T201|COMP|75239-4|LNC|Albumin.ischemia modified|Albumin.ischemia modified
C3846774|T201|COMP|75237-8|LNC|Erythrocytes|Erythrocytes
C3846775|T201|COMP|75236-0|LNC|Crystals|Crystals
C3846776|T201|COMP|75235-2|LNC|Vilazodone|Vilazodone
C3846777|T201|COMP|75234-5|LNC|Norvenlafaxine|Norvenlafaxine
C3846778|T201|COMP|75233-7|LNC|Norsertraline|Norsertraline
C3846779|T201|COMP|75232-9|LNC|Norcitalopram|Norcitalopram
C3846780|T201|COMP|75231-1|LNC|Nefazodone|Nefazodone
C3846781|T201|COMP|75230-3|LNC|m-Chlorophenylpiperazine|m-Chlorophenylpiperazine
C3846782|T201|COMP|75229-5|LNC|DULoxetine|DULoxetine
C3846783|T201|COMP|75228-7|LNC|Carisoprodol+Meprobamate|Carisoprodol+Meprobamate
C3846784|T201|COMP|75227-9|LNC|Baclofen|Baclofen
C3846785|T201|COMP|75226-1|LNC|8-Hydroxyamoxapine|8-Hydroxyamoxapine
C3846786|T201|COMP|75225-3|LNC|Glutarylcarnitine (C5-DC)/Carnitine (C0)|Glutarylcarnitine (C5-DC)/Carnitine (C0)
C3846787|T201|COMP|75224-6|LNC|Chediak-Higashi cells|Chediak-Higashi cells
C3846788|T201|COMP|75223-8|LNC|Dengue virus Ab.IgG & IgM|Dengue virus Ab.IgG & IgM
C3846791|T201|COMP|75217-0|LNC|Biotinidase|Biotinidase
C3846793|T201|COMP|75215-4|LNC|Ornithine/Citrulline|Ornithine/Citrulline
C3846794|T201|COMP|75214-7|LNC|Arginine/Ornithine|Arginine/Ornithine
C3846796|T201|COMP|75212-1|LNC|Malonylcarnitine (C3-DC)/Decanoylcarnitine (C10)|Malonylcarnitine (C3-DC)/Decanoylcarnitine (C10)
C3846797|T201|COMP|75211-3|LNC|Propionylcarnitine (C3)+Palmitoylcarnitine (C16)|Propionylcarnitine (C3)+Palmitoylcarnitine (C16)
C3846841|T201|COMP|75160-2|LNC|Adenosine/Creatinine|Adenosine/Creatinine
C3846842|T201|COMP|75159-4|LNC|Uridine|Uridine
C3846843|T201|COMP|75158-6|LNC|Allantoine|Allantoine
C3846844|T201|COMP|75157-8|LNC|Deoxyinosine|Deoxyinosine
C3846845|T201|COMP|75156-0|LNC|Thymidine|Thymidine
C3846846|T201|COMP|75155-2|LNC|Allantoine/Creatinine|Allantoine/Creatinine
C3846847|T201|COMP|75154-5|LNC|Inosine|Inosine
C3846848|T201|COMP|75153-7|LNC|Thymine|Thymine
C3846849|T201|COMP|75152-9|LNC|Uracil|Uracil
C3846850|T201|COMP|75151-1|LNC|Acadesine/Creatinine|Acadesine/Creatinine
C3846851|T201|COMP|75149-5|LNC|Deoxyguanosine|Deoxyguanosine
C3846852|T201|COMP|75148-7|LNC|Orotidine|Orotidine
C3846853|T201|COMP|75147-9|LNC|Succinylaminoimidazole carboxamide riboside|Succinylaminoimidazole carboxamide riboside
C3846854|T201|COMP|75146-1|LNC|Succinylaminoimidazole carboxamide riboside|Succinylaminoimidazole carboxamide riboside
C3846855|T201|COMP|75145-3|LNC|Succinyladenosine|Succinyladenosine
C3846856|T201|COMP|75144-6|LNC|Xanthine|Xanthine
C3846858|T201|COMP|75137-0|LNC|Acadesine|Acadesine
C3846859|T201|COMP|75136-2|LNC|Adenosine|Adenosine
C3846860|T201|COMP|75135-4|LNC|Hypoxanthine|Hypoxanthine
C3846861|T201|COMP|75134-7|LNC|Deoxyguanosine|Deoxyguanosine
C3846862|T201|COMP|75133-9|LNC|Adenine|Adenine
C3846863|T201|COMP|75132-1|LNC|Oxipurinol/Creatinine|Oxipurinol/Creatinine
C3846864|T201|COMP|75131-3|LNC|Adenine|Adenine
C3846865|T201|COMP|75130-5|LNC|Uridine|Uridine
C3846866|T201|COMP|75129-7|LNC|Xanthine|Xanthine
C3846867|T201|COMP|75128-9|LNC|Uracil|Uracil
C3846868|T201|COMP|75127-1|LNC|Deoxyinosine|Deoxyinosine
C3846869|T201|COMP|75126-3|LNC|Orotate|Orotate
C3846870|T201|COMP|75125-5|LNC|Orotidine|Orotidine
C3846871|T201|COMP|75124-8|LNC|Deoxyadenosine|Deoxyadenosine
C3846872|T201|COMP|75123-0|LNC|Hypoxanthine|Hypoxanthine
C3846873|T201|COMP|75122-2|LNC|Deoxyadenosine|Deoxyadenosine
C3846874|T201|COMP|75121-4|LNC|Thymine|Thymine
C3846875|T201|COMP|75120-6|LNC|Octanoate|Octanoate
C3846876|T201|COMP|75119-8|LNC|Gamma linolenate|Gamma linolenate
C3846877|T201|COMP|75118-0|LNC|Octadecanoate|Octadecanoate
C3846878|T201|COMP|75117-2|LNC|Linoleate|Linoleate
C3846879|T201|COMP|75116-4|LNC|Decanoate|Decanoate
C3846880|T201|COMP|75115-6|LNC|Palmitate|Palmitate
C3846881|T201|COMP|75114-9|LNC|Fatty acids pattern|Fatty acids pattern
C3846882|T201|COMP|75113-1|LNC|Alpha linolenate|Alpha linolenate
C3846883|T201|COMP|75112-3|LNC|Docosatetraenoate|Docosatetraenoate
C3846884|T201|COMP|75111-5|LNC|Palmitoleate|Palmitoleate
C3846885|T201|COMP|75110-7|LNC|Arachidonate|Arachidonate
C3846886|T201|COMP|75109-9|LNC|Fatty acids.very long chain.C22:1n9|Fatty acids.very long chain.C22:1n9
C3846887|T201|COMP|75108-1|LNC|Arachidate|Arachidate
C3846888|T201|COMP|75107-3|LNC|Pentadecanoate|Pentadecanoate
C3846889|T201|COMP|75106-5|LNC|Mead acid|Mead acid
C3846890|T201|COMP|75105-7|LNC|Fatty acids.very long chain.C26:1|Fatty acids.very long chain.C26:1
C3846891|T201|COMP|75104-0|LNC|Fatty acids.very long chain.C24:0|Fatty acids.very long chain.C24:0
C3846892|T201|COMP|75103-2|LNC|Myristate|Myristate
C3846893|T201|COMP|75102-4|LNC|Oleate|Oleate
C3846894|T201|COMP|75101-6|LNC|Fatty acids.very long chain.C22:0|Fatty acids.very long chain.C22:0
C3846895|T201|COMP|75100-8|LNC|Fatty acids|Fatty acids
C3846896|T201|COMP|75099-2|LNC|Laurate|Laurate
C3846897|T201|COMP|75098-4|LNC|Nervonate|Nervonate
C3846898|T201|COMP|75097-6|LNC|Eicosapentaenoate|Eicosapentaenoate
C3846899|T201|COMP|75096-8|LNC|Fatty acids.very long chain.C26:0|Fatty acids.very long chain.C26:0
C3846901|T201|COMP|75093-5|LNC|Galactose^post therapeutic diet|Galactose^post therapeutic diet
C3846902|T201|COMP|75092-7|LNC|Birth date|Birth date
C3846903|T201|COMP|75090-1|LNC|Isocitrate|Isocitrate
C3846904|T201|COMP|75089-3|LNC|5-Oxoproline|5-Oxoproline
C3846905|T201|COMP|75088-5|LNC|3-Indolelactate|3-Indolelactate
C3846906|T201|COMP|75087-7|LNC|Adipate|Adipate
C3846907|T201|COMP|75086-9|LNC|Catecholamine metabolites pattern|Catecholamine metabolites pattern
C3846908|T201|COMP|75085-1|LNC|Homogentisate/Creatinine|Homogentisate/Creatinine
C3846909|T201|COMP|75084-4|LNC|Sebacate|Sebacate
C3846910|T201|COMP|75083-6|LNC|Aconitate|Aconitate
C3846911|T201|COMP|75081-0|LNC|Fumarate|Fumarate
C3846912|T201|COMP|75079-4|LNC|Succinylacetone|Succinylacetone
C3846913|T201|COMP|75078-6|LNC|3-Hydroxydodecanoate/Creatinine|3-Hydroxydodecanoate/Creatinine
C3846914|T201|COMP|75077-8|LNC|Quinolinate|Quinolinate
C3846915|T201|COMP|75076-0|LNC|Vanillate|Vanillate
C3846916|T201|COMP|75075-2|LNC|4-Hydroxybenzoate|4-Hydroxybenzoate
C3846917|T201|COMP|75073-7|LNC|Suberate|Suberate
C3846918|T201|COMP|75072-9|LNC|Mandelate|Mandelate
C3846919|T201|COMP|75071-1|LNC|Acetaminophen/Creatinine|Acetaminophen/Creatinine
C3846920|T201|COMP|75070-3|LNC|Catechol|Catechol
C3846921|T201|COMP|75069-5|LNC|Hippurate|Hippurate
C3846922|T201|COMP|75068-7|LNC|Malate|Malate
C3846923|T201|COMP|75067-9|LNC|Indole-3-Acetate|Indole-3-Acetate
C3846924|T201|COMP|75066-1|LNC|Pantothenate|Pantothenate
C3846925|T201|COMP|75065-3|LNC|Benzoate|Benzoate
C3846926|T201|COMP|75064-6|LNC|Vanillylmandelate|Vanillylmandelate
C3846927|T201|COMP|75063-8|LNC|Glycerate|Glycerate
C3846928|T201|COMP|75062-0|LNC|Phenylacetate|Phenylacetate
C3846929|T201|COMP|75061-2|LNC|Malonate|Malonate
C3846930|T201|COMP|75060-4|LNC|Pantothenate/Creatinine|Pantothenate/Creatinine
C3846931|T201|COMP|75059-6|LNC|Transaldolase|Transaldolase
C3846932|T201|COMP|75058-8|LNC|Thymidine phosphorylase|Thymidine phosphorylase
C3846933|T201|COMP|75057-0|LNC|Sialidase|Sialidase
C3846934|T201|COMP|75056-2|LNC|Pyridoxal phosphate|Pyridoxal phosphate
C3846935|T201|COMP|75055-4|LNC|Glutaryl CoA dehydrogenase|Glutaryl CoA dehydrogenase
C3846936|T201|COMP|75049-7|LNC|Thiosulfate|Thiosulfate
C3846937|T201|COMP|75048-9|LNC|Tetrahydrofolate|Tetrahydrofolate
C3846938|T201|COMP|75047-1|LNC|Sialate|Sialate
C3846939|T201|COMP|75046-3|LNC|Sialate|Sialate
C3846940|T201|COMP|75045-5|LNC|Sialate|Sialate
C3846941|T201|COMP|75044-8|LNC|Sepiapterin/Creatinine|Sepiapterin/Creatinine
C3846942|T201|COMP|75043-0|LNC|Pyridoxine|Pyridoxine
C3846943|T201|COMP|75042-2|LNC|Pyridoxal|Pyridoxal
C3846944|T201|COMP|75041-4|LNC|Pyridoxal|Pyridoxal
C3846945|T201|COMP|75040-6|LNC|D-lactate|D-lactate
C3846946|T201|COMP|75023-2|LNC|Basophils.CD63/100 basophils|Basophils.CD63/100 basophils
C3846947|T201|COMP|75022-4|LNC|Fat.Microscopic Observation|Fat.Microscopic Observation
C3846948|T201|COMP|75021-6|LNC|OLANZapine panel|OLANZapine panel
C3846949|T201|COMP|75020-8|LNC|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript
C3846955|T201|COMP|75014-1|LNC|t(9;12)(q34.1;p13)(ABL1,ETV6) fusion transcript|t(9;12)(q34.1;p13)(ABL1,ETV6) fusion transcript
C3846957|T201|COMP|75012-5|LNC|t(4;11)(q21.3;q23)(AFF1,MLL) fusion transcript|t(4;11)(q21.3;q23)(AFF1,MLL) fusion transcript
C3846958|T201|COMP|75011-7|LNC|t(15;17)(q24.1;q21.1)(PML,RARA) fusion transcript|t(15;17)(q24.1;q21.1)(PML,RARA) fusion transcript
C3846960|T201|COMP|75009-1|LNC|CEBPA gene full mutation analysis|CEBPA gene full mutation analysis
C3846961|T201|COMP|75008-3|LNC|Canis familiaris native (nCan f) 1 Ab.IgE|Canis familiaris native (nCan f) 1 Ab.IgE
C3846962|T201|COMP|75007-5|LNC|Aspergillus restrictus native (nAsp r) 1 Ab.IgE|Aspergillus restrictus native (nAsp r) 1 Ab.IgE
C3846965|T201|COMP|75004-2|LNC|(Beef+Chicken+Pork+Lamb) Ab.IgE|(Beef+Chicken+Pork+Lamb) Ab.IgE
C3846968|T201|COMP|75001-8|LNC|Coproporphyrin 3/Coproporphyrin.total|Coproporphyrin 3/Coproporphyrin.total
C3846969|T201|COMP|75000-0|LNC|Coproporphyrin 3/Coproporphyrin.total|Coproporphyrin 3/Coproporphyrin.total
C3846970|T201|COMP|74999-4|LNC|5,10-Methylenetetrahydrofolate reductase|5,10-Methylenetetrahydrofolate reductase
C3846971|T201|COMP|74998-6|LNC|5,10-Methylenetetrahydrofolate reductase|5,10-Methylenetetrahydrofolate reductase
C3846972|T201|COMP|74997-8|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C3846973|T201|COMP|74996-0|LNC|Alkaline phosphatase.bone|Alkaline phosphatase.bone
C3846974|T201|COMP|74995-2|LNC|Osteocalcin|Osteocalcin
C3846975|T201|COMP|74994-5|LNC|Collagen crosslinked C-telopeptide|Collagen crosslinked C-telopeptide
C3846976|T201|COMP|74992-9|LNC|Amylase|Amylase
C3846977|T201|COMP|74991-1|LNC|Amino acids panel|Amino acids panel
C3846978|T201|COMP|74990-3|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C3846979|T201|COMP|74989-5|LNC|Pentacarboxylporphyrins|Pentacarboxylporphyrins
C3846980|T201|COMP|74988-7|LNC|Hexacarboxylporphyrin|Hexacarboxylporphyrin
C3846981|T201|COMP|74987-9|LNC|Pericyazine^trough|Pericyazine^trough
C3846982|T201|COMP|74986-1|LNC|Hydroxychloroquine^trough|Hydroxychloroquine^trough
C3846983|T201|COMP|74985-3|LNC|ALPRAZolam^trough|ALPRAZolam^trough
C3846984|T201|COMP|74984-6|LNC|5,10-Methylenetetrahydrofolate reductase|5,10-Methylenetetrahydrofolate reductase
C3846985|T201|COMP|74983-8|LNC|Phenytoin.free^trough|Phenytoin.free^trough
C3846986|T201|COMP|74982-0|LNC|FLUoxetine^trough|FLUoxetine^trough
C3846987|T201|COMP|74981-2|LNC|Pimozide^trough|Pimozide^trough
C3846988|T201|COMP|74974-7|LNC|carBAMazepine.free^trough|carBAMazepine.free^trough
C3846989|T201|COMP|74973-9|LNC|carBAMazepine^trough|carBAMazepine^trough
C3846990|T201|COMP|74972-1|LNC|9-Hydroxyrisperidone^trough|9-Hydroxyrisperidone^trough
C3846991|T201|COMP|74971-3|LNC|Clopenthixol^trough|Clopenthixol^trough
C3846992|T201|COMP|74969-7|LNC|Methotrimeprazine^trough|Methotrimeprazine^trough
C3846993|T201|COMP|74968-9|LNC|Norsertraline^trough|Norsertraline^trough
C3846994|T201|COMP|74967-1|LNC|Adrenal cortex Ab.IgG|Adrenal cortex Ab.IgG
C3846995|T201|COMP|74966-3|LNC|Acetaminophen^trough|Acetaminophen^trough
C3846996|T201|COMP|74965-5|LNC|Haloperidol^trough|Haloperidol^trough
C3846997|T201|COMP|74964-8|LNC|Gabapentin^trough|Gabapentin^trough
C3846998|T201|COMP|74963-0|LNC|Promethazine^trough|Promethazine^trough
C3846999|T201|COMP|74962-2|LNC|Maprotiline^trough|Maprotiline^trough
C3847000|T201|COMP|74961-4|LNC|10-Hydroxycarbazepine^trough|10-Hydroxycarbazepine^trough
C3847001|T201|COMP|74960-6|LNC|valGANciclovir^trough|valGANciclovir^trough
C3847002|T201|COMP|74959-8|LNC|fluvoxaMINE^trough|fluvoxaMINE^trough
C3847003|T201|COMP|74958-0|LNC|clomiPRAMINE^trough|clomiPRAMINE^trough
C3847004|T201|COMP|74957-2|LNC|Succinylacetone|Succinylacetone
C3847005|T201|COMP|74956-4|LNC|chlordiazePOXIDE^trough|chlordiazePOXIDE^trough
C3847006|T201|COMP|74955-6|LNC|Cyproheptadine^trough|Cyproheptadine^trough
C3847007|T201|COMP|74954-9|LNC|Isomaltase|Isomaltase
C3847008|T201|COMP|74953-1|LNC|Macroprolactin|Macroprolactin
C3847009|T201|COMP|74951-5|LNC|E-10-Hydroxynortriptyline^trough|E-10-Hydroxynortriptyline^trough
C3847010|T201|COMP|74950-7|LNC|Galactocerebrosidase|Galactocerebrosidase
C3847011|T201|COMP|74949-9|LNC|Perphenazine^trough|Perphenazine^trough
C3847012|T201|COMP|74948-1|LNC|Fluoxetine+Norfluoxetine^trough|Fluoxetine+Norfluoxetine^trough
C3847013|T201|COMP|74947-3|LNC|Norclomipramine^trough|Norclomipramine^trough
C3847014|T201|COMP|74946-5|LNC|Normirtazapine^trough|Normirtazapine^trough
C3847015|T201|COMP|74945-7|LNC|Clomipramine+Norclomipramine^trough|Clomipramine+Norclomipramine^trough
C3847016|T201|COMP|74944-0|LNC|lamoTRIgine^trough|lamoTRIgine^trough
C3847017|T201|COMP|74943-2|LNC|busPIRone^trough|busPIRone^trough
C3847018|T201|COMP|74942-4|LNC|Kynurenin|Kynurenin
C3847019|T201|COMP|74941-6|LNC|Moclobemide|Moclobemide
C3847020|T201|COMP|74940-8|LNC|Moclobemide^trough|Moclobemide^trough
C3847021|T201|COMP|74939-0|LNC|Vigabatrin^trough|Vigabatrin^trough
C3847022|T201|COMP|74938-2|LNC|Lidocaine^trough|Lidocaine^trough
C3847023|T201|COMP|74937-4|LNC|Chlorprothixene^trough|Chlorprothixene^trough
C3847024|T201|COMP|74936-6|LNC|QUEtiapine^trough|QUEtiapine^trough
C3847025|T201|COMP|74935-8|LNC|Palmitoyl protein thioesterase|Palmitoyl protein thioesterase
C3847026|T201|COMP|74934-1|LNC|fluPHENAZine^trough|fluPHENAZine^trough
C3847027|T201|COMP|74933-3|LNC|N-desalkylflurazepam^trough|N-desalkylflurazepam^trough
C3847028|T201|COMP|74932-5|LNC|Citalopram^trough|Citalopram^trough
C3847029|T201|COMP|74931-7|LNC|ARIPiprazole^trough|ARIPiprazole^trough
C3847030|T201|COMP|74930-9|LNC|3-Hydroxykynurenin|3-Hydroxykynurenin
C3847031|T201|COMP|74929-1|LNC|Fluspirilene^trough|Fluspirilene^trough
C3847032|T201|COMP|74928-3|LNC|Allopurinol^trough|Allopurinol^trough
C3847033|T201|COMP|74927-5|LNC|Pipamperone^trough|Pipamperone^trough
C3847034|T201|COMP|74926-7|LNC|PHENobarbital^trough|PHENobarbital^trough
C3847035|T201|COMP|74925-9|LNC|Flupenthixol^trough|Flupenthixol^trough
C3847036|T201|COMP|74924-2|LNC|Nortriptyline^trough|Nortriptyline^trough
C3847037|T201|COMP|74923-4|LNC|Temazepam^trough|Temazepam^trough
C3847038|T201|COMP|74922-6|LNC|N-acetyl-L-aspartate|N-acetyl-L-aspartate
C3847039|T201|COMP|74921-8|LNC|Norclobazam^trough|Norclobazam^trough
C3847040|T201|COMP|74920-0|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C3847041|T201|COMP|74919-2|LNC|Caffeine^trough|Caffeine^trough
C3847042|T201|COMP|74918-4|LNC|Fatty acids|Fatty acids
C3847043|T201|COMP|74917-6|LNC|CXCL13 Ag|CXCL13 Ag
C3847044|T201|COMP|74916-8|LNC|Metoprolol^trough|Metoprolol^trough
C3847045|T201|COMP|74915-0|LNC|Sulpiride^trough|Sulpiride^trough
C3847046|T201|COMP|74913-5|LNC|Escitalopram^trough|Escitalopram^trough
C3847047|T201|COMP|74912-7|LNC|Primidone^trough|Primidone^trough
C3847048|T201|COMP|74911-9|LNC|Sertraline^trough|Sertraline^trough
C3847049|T201|COMP|74909-3|LNC|Calcium oxalate dihydrate/Total|Calcium oxalate dihydrate/Total
C3847050|T201|COMP|74908-5|LNC|3-ketoacyl-CoA thiolase|3-ketoacyl-CoA thiolase
C3847051|T201|COMP|74907-7|LNC|Beta sitosterol|Beta sitosterol
C3847052|T201|COMP|74906-9|LNC|Bilirubin|Bilirubin
C3847053|T201|COMP|74905-1|LNC|Desmosterol|Desmosterol
C3847054|T201|COMP|74904-4|LNC|DOPamine|DOPamine
C3847055|T201|COMP|74903-6|LNC|Fatty acids|Fatty acids
C3847056|T201|COMP|74902-8|LNC|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C3847057|T201|COMP|74901-0|LNC|Gamma tocopherol|Gamma tocopherol
C3847058|T201|COMP|74900-2|LNC|Lactulose/Creatinine^post XXX g sugar solution PO|Lactulose/Creatinine^post XXX g sugar solution PO
C3847059|T201|COMP|74899-6|LNC|Lactulose/mannitol^post XXX g sugar solution PO|Lactulose/mannitol^post XXX g sugar solution PO
C3847060|T201|COMP|74898-8|LNC|Lanosterol|Lanosterol
C3847061|T201|COMP|74897-0|LNC|Lithocholate|Lithocholate
C3847062|T201|COMP|74896-2|LNC|Lactate|Lactate
C3847063|T201|COMP|74895-4|LNC|Maltose/Creatinine|Maltose/Creatinine
C3847064|T201|COMP|74894-7|LNC|Mannitol^post XXX g sugar solution PO|Mannitol^post XXX g sugar solution PO
C3847065|T201|COMP|74893-9|LNC|Mannose/Creatinine|Mannose/Creatinine
C3847066|T201|COMP|74892-1|LNC|Medium-chain Acyl CoA dehydrogenase|Medium-chain Acyl CoA dehydrogenase
C3847067|T201|COMP|74891-3|LNC|Medium-chain Acyl CoA dehydrogenase|Medium-chain Acyl CoA dehydrogenase
C3847068|T201|COMP|74890-5|LNC|Inositol.free/Creatinine|Inositol.free/Creatinine
C3847069|T201|COMP|74889-7|LNC|Phosphate|Phosphate
C3847070|T201|COMP|74888-9|LNC|Sterols panel|Sterols panel
C3847071|T201|COMP|74887-1|LNC|Stigmastanol|Stigmastanol
C3847072|T201|COMP|74886-3|LNC|Stigmasterol|Stigmasterol
C3847073|T201|COMP|74885-5|LNC|HER2 panel|HER2 panel
C3847074|T201|COMP|74884-8|LNC|Valine^post therapeutic diet|Valine^post therapeutic diet
C3847075|T201|COMP|74883-0|LNC|Ornithine^post therapeutic diet|Ornithine^post therapeutic diet
C3847076|T201|COMP|74882-2|LNC|Leucine^post therapeutic diet|Leucine^post therapeutic diet
C3847077|T201|COMP|74881-4|LNC|Isoleucine^post therapeutic diet|Isoleucine^post therapeutic diet
C3847078|T201|COMP|74880-6|LNC|Hydroxyproline^post therapeutic diet|Hydroxyproline^post therapeutic diet
C3847079|T201|COMP|74879-8|LNC|Galactose 1 phosphate^post therapeutic diet|Galactose 1 phosphate^post therapeutic diet
C3847080|T201|COMP|74878-0|LNC|Carnitine.free (C0)^post therapeutic diet|Carnitine.free (C0)^post therapeutic diet
C3847081|T201|COMP|74877-2|LNC|Argininosuccinate^post therapeutic diet|Argininosuccinate^post therapeutic diet
C3847082|T201|COMP|74876-4|LNC|Arginine^post therapeutic diet|Arginine^post therapeutic diet
C3847083|T201|COMP|74875-6|LNC|Alloisoleucine^post therapeutic diet|Alloisoleucine^post therapeutic diet
C3847084|T201|COMP|74874-9|LNC|Metabolic disorder therapy monitoring panel|Metabolic disorder therapy monitoring panel
C3847085|T201|COMP|74873-1|LNC|Metabolic disorder being monitored|Metabolic disorder being monitored
C3847086|T201|COMP|74872-3|LNC|21-Deoxycortisol|21-Deoxycortisol
C3847087|T201|COMP|74871-5|LNC|Rivaroxaban|Rivaroxaban
C3847088|T201|COMP|74870-7|LNC|IgM.kappa/IgM.lambda|IgM.kappa/IgM.lambda
C3847089|T201|COMP|74864-0|LNC|IgA.kappa|IgA.kappa
C3847090|T201|COMP|74863-2|LNC|IgG.lambda|IgG.lambda
C3847091|T201|COMP|74862-4|LNC|IgG.kappa|IgG.kappa
C3847092|T201|COMP|74861-6|LNC|Chromosome 17 copy number/nucleus|Chromosome 17 copy number/nucleus
C3847093|T201|COMP|74860-8|LNC|HER2 gene copy number/nucleus|HER2 gene copy number/nucleus
C3847094|T201|COMP|74858-2|LNC|Hepatitis E virus genotypes 1+2+3+4 RNA|Hepatitis E virus genotypes 1+2+3+4 RNA
C3847095|T201|COMP|74857-4|LNC|West Nile Virus RNA|West Nile Virus RNA
C3847097|T201|COMP|74855-8|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C3847098|T201|COMP|74854-1|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C3847099|T201|COMP|74846-7|LNC|Snowshoe hare virus Ab.IgM|Snowshoe hare virus Ab.IgM
C3847100|T201|COMP|74845-9|LNC|Sindbis virus Ab|Sindbis virus Ab
C3847101|T201|COMP|74844-2|LNC|Baylisascaris sp Ab.IgG|Baylisascaris sp Ab.IgG
C3847102|T201|COMP|74843-4|LNC|Baylisascaris sp Ab.IgG|Baylisascaris sp Ab.IgG
C3847103|T201|COMP|74842-6|LNC|Cells.CD25|Cells.CD25
C3847104|T201|COMP|74841-8|LNC|Cells.CD8+CD57+/100 cells|Cells.CD8+CD57+/100 cells
C3847105|T201|COMP|74840-0|LNC|Cells.CD56|Cells.CD56
C3847106|T201|COMP|74839-2|LNC|Cells.CD3-CD4+/100 cells|Cells.CD3-CD4+/100 cells
C3847107|T201|COMP|74838-4|LNC|Cells.CD34|Cells.CD34
C3847108|T201|COMP|74837-6|LNC|Cells.CD20|Cells.CD20
C3847109|T201|COMP|74830-1|LNC|Toxoplasma gondii Ab.IgA|Toxoplasma gondii Ab.IgA
C3847110|T201|COMP|74829-3|LNC|Snowshoe hare virus Ab.IgG|Snowshoe hare virus Ab.IgG
C3847111|T201|COMP|74828-5|LNC|Snowshoe hare virus Ab|Snowshoe hare virus Ab
C3847112|T201|COMP|74827-7|LNC|Snowshoe hare virus Ab|Snowshoe hare virus Ab
C3847113|T201|COMP|74826-9|LNC|Semliki forest virus Ab|Semliki forest virus Ab
C3847114|T201|COMP|74825-1|LNC|Saint Louis encephalitis virus Ab|Saint Louis encephalitis virus Ab
C3847115|T201|COMP|74824-4|LNC|Powassan virus Ab|Powassan virus Ab
C3847116|T201|COMP|74823-6|LNC|Jamestown canyon virus Ab|Jamestown canyon virus Ab
C3847117|T201|COMP|74822-8|LNC|Clostridioides difficile toxin B tcdB gene|Clostridioides difficile toxin B tcdB gene
C3847118|T201|COMP|74821-0|LNC|Chikungunya virus Ab|Chikungunya virus Ab
C3847119|T201|COMP|74819-4|LNC|Promazine|Promazine
C3847120|T201|COMP|74818-6|LNC|Desomorphine|Desomorphine
C3847121|T201|COMP|74817-8|LNC|Desomorphine|Desomorphine
C3847122|T201|COMP|74816-0|LNC|Bacteria identified|Bacteria identified
C3847123|T201|COMP|74815-2|LNC|Ascaris sp Ab.IgG|Ascaris sp Ab.IgG
C3847124|T201|COMP|74813-7|LNC|Nucleated cells|Nucleated cells
C3847125|T201|COMP|74812-9|LNC|Mirtazapine|Mirtazapine
C3847126|T201|COMP|74811-1|LNC|Dihydrocodeine|Dihydrocodeine
C3847127|T201|COMP|74810-3|LNC|Acetyl fentaNYL|Acetyl fentaNYL
C3847128|T201|COMP|74805-3|LNC|Penicillium sp Ab.IgG|Penicillium sp Ab.IgG
C3847129|T201|COMP|74804-6|LNC|Fructose challenge|Fructose challenge
C3847130|T201|COMP|74803-8|LNC|Lactose challenge|Lactose challenge
C3847131|T201|COMP|74802-0|LNC|Glucose challenge|Glucose challenge
C3847132|T201|COMP|74795-6|LNC|Total thyroxine binding capacity|Total thyroxine binding capacity
C3847133|T201|COMP|74794-9|LNC|Thyroid hormone binding ratio|Thyroid hormone binding ratio
C3847134|T201|COMP|74793-1|LNC|Thyroid hormone uptake|Thyroid hormone uptake
C3847135|T201|COMP|74792-3|LNC|Fructose.PO|Fructose.PO
C3847136|T201|COMP|74791-5|LNC|Lactulose challenge|Lactulose challenge
C3847137|T201|COMP|74785-7|LNC|Influenza virus B Victoria lineage RNA|Influenza virus B Victoria lineage RNA
C3847138|T201|COMP|74784-0|LNC|Influenza virus B lineage RNA|Influenza virus B lineage RNA
C3847139|T201|COMP|74783-2|LNC|Malignant cells|Malignant cells
C3847142|T201|COMP|74780-8|LNC|CPT1A gene.c.1436C>T|CPT1A gene.c.1436C>T
C3847143|T201|COMP|74779-0|LNC|Human papilloma virus 11 DNA|Human papilloma virus 11 DNA
C3847144|T201|COMP|74778-2|LNC|Human papilloma virus 11 DNA|Human papilloma virus 11 DNA
C3847145|T201|COMP|74777-4|LNC|Human papilloma virus 6 DNA|Human papilloma virus 6 DNA
C3847146|T201|COMP|74776-6|LNC|Human papilloma virus 6 DNA|Human papilloma virus 6 DNA
C3847147|T201|COMP|74775-8|LNC|Platelets|Platelets
C3847148|T201|COMP|74774-1|LNC|Glucose|Glucose
C3847149|T201|COMP|74773-3|LNC|Immunoglobulin light chains & heavy chains panel|Immunoglobulin light chains & heavy chains panel
C3847153|T201|COMP|74769-1|LNC|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C3847154|T201|COMP|74768-3|LNC|5-hydroxytryptophan|5-hydroxytryptophan
C3847155|T201|COMP|74767-5|LNC|Tryptophan|Tryptophan
C3847156|T201|COMP|74766-7|LNC|Bordetella pertussis.pertussis toxin 100 Ab.IgG|Bordetella pertussis.pertussis toxin 100 Ab.IgG
C3847157|T201|COMP|74765-9|LNC|Bordetella pertussis.pertussis toxin Ab.IgA|Bordetella pertussis.pertussis toxin Ab.IgA
C3847160|T201|COMP|74762-6|LNC|Megasphaera sp DNA|Megasphaera sp DNA
C3847161|T201|COMP|74761-8|LNC|Microcytes/100 erythrocytes|Microcytes/100 erythrocytes
C3847162|T201|COMP|74760-0|LNC|HYDROcodone & metabolites panel|HYDROcodone & metabolites panel
C3847163|T201|COMP|74759-2|LNC|Yeast|Yeast
C3847164|T201|COMP|74758-4|LNC|Ethyl sulfate+Ethyl glucuronide|Ethyl sulfate+Ethyl glucuronide
C3847166|T201|COMP|74756-8|LNC|Soluble fms-like tyrosine kinase-1|Soluble fms-like tyrosine kinase-1
C3847167|T201|COMP|74755-0|LNC|Placental growth factor|Placental growth factor
C3847168|T201|COMP|74754-3|LNC|Blood group antigens present|Blood group antigens present
C3847169|T201|COMP|74753-5|LNC|Blood group antigens present|Blood group antigens present
C3847170|T201|COMP|74752-7|LNC|Porcine epidemic diarrhea virus RNA|Porcine epidemic diarrhea virus RNA
C3847171|T201|COMP|74751-9|LNC|Collection time|Collection time
C3847172|T201|COMP|74750-1|LNC|Lymphocytes.clefted|Lymphocytes.clefted
C3847173|T201|COMP|74749-3|LNC|Gram positive blood culture panel|Gram positive blood culture panel
C3847174|T201|COMP|74748-5|LNC|Staphylococcus sp tuf gene|Staphylococcus sp tuf gene
C3847175|T201|COMP|74747-7|LNC|Staphylococcus aureus gyrB gene|Staphylococcus aureus gyrB gene
C3847176|T201|COMP|74746-9|LNC|Staphylococcus epidermidis hsp60 gene|Staphylococcus epidermidis hsp60 gene
C3847177|T201|COMP|74745-1|LNC|Bacterial methicillin resistance (mecA) gene|Bacterial methicillin resistance (mecA) gene
C3847178|T201|COMP|74744-4|LNC|Staphylococcus lugdunensis sodA gene|Staphylococcus lugdunensis sodA gene
C3847179|T201|COMP|74743-6|LNC|Enterococcus faecalis hsp60 gene|Enterococcus faecalis hsp60 gene
C3847180|T201|COMP|74742-8|LNC|Bacterial vancomycin resistance vanA gene|Bacterial vancomycin resistance vanA gene
C3847181|T201|COMP|74741-0|LNC|Bacterial vancomycin resistance vanB gene|Bacterial vancomycin resistance vanB gene
C3847182|T201|COMP|75054-7|LNC|Glutaryl CoA dehydrogenase|Glutaryl CoA dehydrogenase
C3847183|T201|COMP|75053-9|LNC|Alpha-L-iduronidase|Alpha-L-iduronidase
C3847184|T201|COMP|75052-1|LNC|Adenosine deaminase|Adenosine deaminase
C3847185|T201|COMP|75051-3|LNC|Xylose/Creatinine|Xylose/Creatinine
C3847186|T201|COMP|75050-5|LNC|Ubiquinone 10|Ubiquinone 10
C3847187|T201|COMP|74980-4|LNC|LORazepam^trough|LORazepam^trough
C3847188|T201|COMP|74979-6|LNC|Urate|Urate
C3847190|T201|COMP|74977-0|LNC|Transferrin|Transferrin
C3847191|T201|COMP|74976-2|LNC|Phenytoin^trough|Phenytoin^trough
C3847192|T201|COMP|74975-4|LNC|Nordiazepam^trough|Nordiazepam^trough
C3847194|T201|COMP|74835-0|LNC|Porphyrin fractions panel|Porphyrin fractions panel
C3847195|T201|COMP|74834-3|LNC|MARS2 gene full mutation analysis|MARS2 gene full mutation analysis
C3847196|T201|COMP|74833-5|LNC|ACAT1 gene full mutation analysis|ACAT1 gene full mutation analysis
C3847197|T201|COMP|74832-7|LNC|OLANZapine|OLANZapine
C3847198|T201|COMP|74831-9|LNC|Metanephrine & Normetanephrine panel|Metanephrine & Normetanephrine panel
C3847199|T201|COMP|74740-2|LNC|Streptococcus sp tuf gene|Streptococcus sp tuf gene
C3847200|T201|COMP|74739-4|LNC|Streptococcus agalactiae hsp60 gene|Streptococcus agalactiae hsp60 gene
C3847201|T201|COMP|74738-6|LNC|Streptococcus anginosus group gyrB gene|Streptococcus anginosus group gyrB gene
C3847202|T201|COMP|74737-8|LNC|Streptococcus pneumoniae gryB gene|Streptococcus pneumoniae gryB gene
C3847203|T201|COMP|74736-0|LNC|Streptococcus pyogenes hsp60 gene|Streptococcus pyogenes hsp60 gene
C3847204|T201|COMP|74735-2|LNC|Health data repository|Health data repository
C3847205|T201|COMP|74729-5|LNC|Adrenoleukodystrophy protein|Adrenoleukodystrophy protein
C3847226|T201|COMP|74699-0|LNC|Cefuroxime|Cefuroxime
C3847228|T201|COMP|74697-4|LNC|Acamprosate|Acamprosate
C3847229|T201|COMP|74696-6|LNC|Magnesium|Magnesium
C3847232|T201|COMP|74692-5|LNC|MT-ND6 gene.m.14459G>A|MT-ND6 gene.m.14459G>A
C3847233|T201|COMP|74691-7|LNC|Round Cells|Round Cells
C3847234|T201|COMP|74690-9|LNC|D little u Ag|D little u Ag
C3847235|T201|COMP|74689-1|LNC|Nucleated cells|Nucleated cells
C3847236|T201|COMP|74688-3|LNC|Sodium^post dialysis|Sodium^post dialysis
C3847237|T201|COMP|74687-5|LNC|Glucose|Glucose
C3847238|T201|COMP|74686-7|LNC|Glucose|Glucose
C3847239|T201|COMP|74685-9|LNC|Sodium|Sodium
C3847240|T201|COMP|74684-2|LNC|Carbon dioxide^post dialysis|Carbon dioxide^post dialysis
C3847241|T201|COMP|74683-4|LNC|Ethyl sulfate|Ethyl sulfate
C3847242|T201|COMP|74682-6|LNC|Trichloroethanol.free|Trichloroethanol.free
C3847243|T201|COMP|74680-0|LNC|Amphetamine|Amphetamine
C3847243|T201|COMP|74681-8|LNC|Amphetamines|Amphetamines
C3847244|T201|COMP|74679-2|LNC|Benzoylecgonine|Benzoylecgonine
C3847245|T201|COMP|74678-4|LNC|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C3847246|T201|COMP|74677-6|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C3847247|T201|COMP|74676-8|LNC|Carbapenemase|Carbapenemase
C3847248|T201|COMP|74675-0|LNC|Codeine|Codeine
C3847249|T201|COMP|74674-3|LNC|Chlorinated solvents|Chlorinated solvents
C3847250|T201|COMP|74673-5|LNC|Ethanol|Ethanol
C3847251|T201|COMP|74672-7|LNC|Carisoprodol+Meprobamate|Carisoprodol+Meprobamate
C3847252|T201|COMP|74671-9|LNC|Cocaine|Cocaine
C3847253|T201|COMP|74670-1|LNC|Cocaine+Metabolites|Cocaine+Metabolites
C3847254|T201|COMP|74669-3|LNC|Lactobacillus sp DNA|Lactobacillus sp DNA
C3847255|T201|COMP|74668-5|LNC|Gardnerella vaginalis DNA|Gardnerella vaginalis DNA
C3847256|T201|COMP|74667-7|LNC|Atopobium vaginae DNA|Atopobium vaginae DNA
C3847257|T201|COMP|74666-9|LNC|Monoclonal band observed|Monoclonal band observed
C3847258|T201|COMP|74665-1|LNC|Monoclonal band observed|Monoclonal band observed
C3847259|T201|COMP|74664-4|LNC|Zolpidem|Zolpidem
C3847260|T201|COMP|74663-6|LNC|Zaleplon|Zaleplon
C3847261|T201|COMP|74662-8|LNC|Sertraline|Sertraline
C3847262|T201|COMP|74661-0|LNC|Phosphatidylethanol|Phosphatidylethanol
C3847263|T201|COMP|74660-2|LNC|Phencyclidine|Phencyclidine
C3847264|T201|COMP|74659-4|LNC|oxyMORphone|oxyMORphone
C3847265|T201|COMP|74658-6|LNC|oxyCODONE+Oxymorphone|oxyCODONE+Oxymorphone
C3847266|T201|COMP|74657-8|LNC|oxyCODONE|oxyCODONE
C3847267|T201|COMP|74656-0|LNC|Opiates|Opiates
C3847268|T201|COMP|74655-2|LNC|Norsertraline|Norsertraline
C3847269|T201|COMP|74654-5|LNC|Morphine|Morphine
C3847270|T201|COMP|74653-7|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C3847271|T201|COMP|74651-1|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C3847272|T201|COMP|74650-3|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C3847273|T201|COMP|74649-5|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C3847274|T201|COMP|74648-7|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C3847275|T201|COMP|74647-9|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C3847276|T201|COMP|74646-1|LNC|Methamphetamine|Methamphetamine
C3847277|T201|COMP|74645-3|LNC|HYDROmorphone|HYDROmorphone
C3847278|T201|COMP|75039-8|LNC|Biopterin|Biopterin
C3847279|T201|COMP|75038-0|LNC|Bile acid pattern|Bile acid pattern
C3847280|T201|COMP|75027-3|LNC|Mesoporphyrin/Porphyrins.total|Mesoporphyrin/Porphyrins.total
C3847281|T201|COMP|75026-5|LNC|Deuteroporphyrin/Porphyrins.total|Deuteroporphyrin/Porphyrins.total
C3847282|T201|COMP|75025-7|LNC|Coproporphyrin 3/Porphyrins.total|Coproporphyrin 3/Porphyrins.total
C3847283|T201|COMP|75024-0|LNC|Coproporphyrin 1/Porphyrins.total|Coproporphyrin 1/Porphyrins.total
C3847284|T201|COMP|74869-9|LNC|IgA.kappa/IgA.lambda|IgA.kappa/IgA.lambda
C3847285|T201|COMP|74868-1|LNC|IgG.kappa/IgG.lambda|IgG.kappa/IgG.lambda
C3847286|T201|COMP|74867-3|LNC|IgM.lambda|IgM.lambda
C3847287|T201|COMP|74866-5|LNC|IgM.kappa|IgM.kappa
C3847288|T201|COMP|74790-7|LNC|Glucose challenge panel|Glucose challenge panel
C3847289|T201|COMP|74789-9|LNC|Fructose challenge panel|Fructose challenge panel
C3847290|T201|COMP|74788-1|LNC|Lactulose challenge panel|Lactulose challenge panel
C3847292|T201|COMP|74786-5|LNC|Influenza virus B Yamagata lineage RNA|Influenza virus B Yamagata lineage RNA
C3847293|T201|COMP|74733-7|LNC|Mycobacterium sp rRNA|Mycobacterium sp rRNA
C3847294|T201|COMP|74732-9|LNC|Listeria sp (tuf) gene|Listeria sp (tuf) gene
C3847295|T201|COMP|74731-1|LNC|Gram positive bacteria identified|Gram positive bacteria identified
C3847296|T201|COMP|74730-3|LNC|Oligosaccharides pattern|Oligosaccharides pattern
C3847297|T201|COMP|74640-4|LNC|Monoclonal band 3 observed|Monoclonal band 3 observed
C3847298|T201|COMP|74639-6|LNC|Monoclonal band 2 observed|Monoclonal band 2 observed
C3847299|T201|COMP|74638-8|LNC|Monoclonal band 3 observed|Monoclonal band 3 observed
C3847300|T201|COMP|74637-0|LNC|Protein.monoclonal band 2|Protein.monoclonal band 2
C3847301|T201|COMP|74636-2|LNC|Protein.monoclonal band 3|Protein.monoclonal band 3
C3847302|T201|COMP|74635-4|LNC|Bacterial vaginosis DNA panel|Bacterial vaginosis DNA panel
C3847303|T201|COMP|74634-7|LNC|Dimethylacetal panel|Dimethylacetal panel
C3847304|T201|COMP|74633-9|LNC|Dimethylacetal panel|Dimethylacetal panel
C3847305|T201|COMP|74632-1|LNC|Glycosaminoglycans|Glycosaminoglycans
C3847306|T201|COMP|74631-3|LNC|Glycosaminoglycans/Creatinine|Glycosaminoglycans/Creatinine
C3847309|T201|COMP|74628-9|LNC|Adipoylcarnitine (C6-DC)|Adipoylcarnitine (C6-DC)
C3847310|T201|COMP|74627-1|LNC|1,1-Dimethoxyhexadecane|1,1-Dimethoxyhexadecane
C3847311|T201|COMP|74626-3|LNC|1,1-Dimethoxyhexadecane|1,1-Dimethoxyhexadecane
C3847312|T201|COMP|74625-5|LNC|1,1-Dimethoxyhexadecane/palmitate|1,1-Dimethoxyhexadecane/palmitate
C3847313|T201|COMP|74624-8|LNC|1,1-Dimethoxyhexadecane/palmitate|1,1-Dimethoxyhexadecane/palmitate
C3847314|T201|COMP|74623-0|LNC|1,1-Dimethoxy-(9Z)octadecene|1,1-Dimethoxy-(9Z)octadecene
C3847315|T201|COMP|74622-2|LNC|1,1-Dimethoxy-(9Z)octadecene|1,1-Dimethoxy-(9Z)octadecene
C3847316|T201|COMP|74621-4|LNC|1,1-Dimethoxy-(9Z)octadecene/oleate|1,1-Dimethoxy-(9Z)octadecene/oleate
C3847317|T201|COMP|74620-6|LNC|1,1-Dimethoxy-(9Z)octadecene/oleate|1,1-Dimethoxy-(9Z)octadecene/oleate
C3847318|T201|COMP|74619-8|LNC|1,1-Dimethoxyoctadecane|1,1-Dimethoxyoctadecane
C3847319|T201|COMP|74618-0|LNC|1,1-Dimethoxyoctadecane|1,1-Dimethoxyoctadecane
C3847320|T201|COMP|74617-2|LNC|1,1-Dimethoxyoctadecane/octadecanoate|1,1-Dimethoxyoctadecane/octadecanoate
C3847321|T201|COMP|74616-4|LNC|1,1-Dimethoxyoctadecane/octadecanoate|1,1-Dimethoxyoctadecane/octadecanoate
C3847322|T201|COMP|74615-6|LNC|Fatty acids.very long chain.C22:0|Fatty acids.very long chain.C22:0
C3847323|T201|COMP|74614-9|LNC|Fatty acids.very long chain.C26:0|Fatty acids.very long chain.C26:0
C3847324|T201|COMP|74613-1|LNC|Fatty acids.very long chain.C24:0|Fatty acids.very long chain.C24:0
C3847325|T201|COMP|74612-3|LNC|Decanoylcarnitine (C10)|Decanoylcarnitine (C10)
C3847326|T201|COMP|74611-5|LNC|Decenoylcarnitine (C10:1)|Decenoylcarnitine (C10:1)
C3847327|T201|COMP|74610-7|LNC|Decadienoylcarnitine (C10:2)|Decadienoylcarnitine (C10:2)
C3847328|T201|COMP|74609-9|LNC|Sebacylcarnitine (C10-DC)|Sebacylcarnitine (C10-DC)
C3847329|T201|COMP|74608-1|LNC|Dodecanoylcarnitine (C12)|Dodecanoylcarnitine (C12)
C3847330|T201|COMP|74607-3|LNC|Dodecenoylcarnitine (C12:1)|Dodecenoylcarnitine (C12:1)
C3847331|T201|COMP|74606-5|LNC|Tetradecanoylcarnitine (C14)|Tetradecanoylcarnitine (C14)
C3847332|T201|COMP|74605-7|LNC|Tetradecenoylcarnitine (C14:1)|Tetradecenoylcarnitine (C14:1)
C3847333|T201|COMP|74604-0|LNC|3-Hydroxymyristoleylcarnitine (C14:1-OH)|3-Hydroxymyristoleylcarnitine (C14:1-OH)
C3847334|T201|COMP|74603-2|LNC|Tetradecadienoylcarnitine (C14:2)|Tetradecadienoylcarnitine (C14:2)
C3847335|T201|COMP|74602-4|LNC|3-Hydroxytetradecanoylcarnitine (C14-OH)|3-Hydroxytetradecanoylcarnitine (C14-OH)
C3847336|T201|COMP|74601-6|LNC|Palmitoylcarnitine (C16)|Palmitoylcarnitine (C16)
C3847337|T201|COMP|74600-8|LNC|Palmitoleylcarnitine (C16:1)|Palmitoleylcarnitine (C16:1)
C3847338|T201|COMP|74599-2|LNC|3-Hydroxypalmitoleylcarnitine (C16:1-OH)|3-Hydroxypalmitoleylcarnitine (C16:1-OH)
C3847339|T201|COMP|74598-4|LNC|Dicarboxypalmitoylcarnitine (C16-DC)|Dicarboxypalmitoylcarnitine (C16-DC)
C3847340|T201|COMP|74597-6|LNC|3-Hydroxypalmitoylcarnitine (C16-OH)|3-Hydroxypalmitoylcarnitine (C16-OH)
C3847341|T201|COMP|74596-8|LNC|Butyrylcarnitine (C4)|Butyrylcarnitine (C4)
C3847342|T201|COMP|74595-0|LNC|3-Hydroxybutyrylcarnitine (C4-OH)|3-Hydroxybutyrylcarnitine (C4-OH)
C3847343|T201|COMP|74594-3|LNC|Hexanoylcarnitine (C6)|Hexanoylcarnitine (C6)
C3847344|T201|COMP|74593-5|LNC|Adipoylcarnitine (C6-DC)|Adipoylcarnitine (C6-DC)
C3847345|T201|COMP|74592-7|LNC|Octanoylcarnitine (C8)|Octanoylcarnitine (C8)
C3847346|T201|COMP|74591-9|LNC|Suberylcarnitine (C8-DC)|Suberylcarnitine (C8-DC)
C3847347|T201|COMP|74590-1|LNC|NADH cytochrome C reductase/Citrate synthase|NADH cytochrome C reductase/Citrate synthase
C3847348|T201|COMP|74589-3|LNC|Succinate dehydrogenase/Citrate synthase|Succinate dehydrogenase/Citrate synthase
C3847349|T201|COMP|74588-5|LNC|Succinate cytochrome C reductase|Succinate cytochrome C reductase
C3847350|T201|COMP|74587-7|LNC|Succinate cytochrome C reductase/Citrate synthase|Succinate cytochrome C reductase/Citrate synthase
C3847351|T201|COMP|74586-9|LNC|Coenzyme Q cytochrome C reductase|Coenzyme Q cytochrome C reductase
C3847353|T201|COMP|74584-4|LNC|Cytochrome C oxidase/Citrate synthase|Cytochrome C oxidase/Citrate synthase
C3847354|T201|COMP|74583-6|LNC|Fatty acids.very long chain.C24:0/C22:0|Fatty acids.very long chain.C24:0/C22:0
C3847355|T201|COMP|74582-8|LNC|Fatty acids.very long chain.C26:0/C22:0|Fatty acids.very long chain.C26:0/C22:0
C3847356|T201|COMP|74581-0|LNC|Fumarase|Fumarase
C3847357|T201|COMP|74580-2|LNC|Fumarase|Fumarase
C3847358|T201|COMP|74579-4|LNC|Pyruvate dehydrogenase E1|Pyruvate dehydrogenase E1
C3847359|T201|COMP|74578-6|LNC|Pyruvate dehydrogenase complex|Pyruvate dehydrogenase complex
C3847360|T201|COMP|74577-8|LNC|Pyruvate dehydrogenase complex|Pyruvate dehydrogenase complex
C3847361|T201|COMP|74545-5|LNC|Tryptophan-related indole profiling panel|Tryptophan-related indole profiling panel
C3847362|T201|COMP|74544-8|LNC|Tocopherols|Tocopherols
C3847363|T201|COMP|74542-2|LNC|Pyruvate kinase/Glucose-6-Phosphate dehydrogenase|Pyruvate kinase/Glucose-6-Phosphate dehydrogenase
C3847364|T201|COMP|74541-4|LNC|Surfactant pulmonary-associated protein D|Surfactant pulmonary-associated protein D
C3847365|T201|COMP|74540-6|LNC|Hexenoylcarnitine (C6:1)|Hexenoylcarnitine (C6:1)
C3847366|T201|COMP|74539-8|LNC|Neisseria meningitidis serogroup A DNA|Neisseria meningitidis serogroup A DNA
C3847367|T201|COMP|74538-0|LNC|Neisseria meningitidis serogroup B DNA|Neisseria meningitidis serogroup B DNA
C3847368|T201|COMP|74537-2|LNC|Neisseria meningitidis serogroup C DNA|Neisseria meningitidis serogroup C DNA
C3847369|T201|COMP|74536-4|LNC|Neisseria meningitidis serogroup w135 DNA|Neisseria meningitidis serogroup w135 DNA
C3847370|T201|COMP|74535-6|LNC|Neisseria meningitidis serogroup X DNA|Neisseria meningitidis serogroup X DNA
C3847371|T201|COMP|74534-9|LNC|Neisseria meningitidis serogroup Y DNA|Neisseria meningitidis serogroup Y DNA
C3847372|T201|COMP|74531-5|LNC|Dicarboxytetradecanoylcarnitine (C14-DC)|Dicarboxytetradecanoylcarnitine (C14-DC)
C3847373|T201|COMP|74530-7|LNC|Dicarboxypalmitoleylcarnitine (C16:1-DC)|Dicarboxypalmitoleylcarnitine (C16:1-DC)
C3847374|T201|COMP|74529-9|LNC|Dicarboxyhexenoylcarnitine (C6:1-DC)|Dicarboxyhexenoylcarnitine (C6:1-DC)
C3847375|T201|COMP|74528-1|LNC|Dicarboxyeicosanoylcarnitine (C20-DC)|Dicarboxyeicosanoylcarnitine (C20-DC)
C3847378|T201|COMP|74525-7|LNC|Dehydrosebacylcarnitine (C10:1-DC)|Dehydrosebacylcarnitine (C10:1-DC)
C3847379|T201|COMP|74524-0|LNC|Decatrienoylcarnitine (C10:3)|Decatrienoylcarnitine (C10:3)
C3847380|T201|COMP|74523-2|LNC|Nonanoylcarnitine (C9)|Nonanoylcarnitine (C9)
C3847381|T201|COMP|74522-4|LNC|Complement lectin pathway actual/normal|Complement lectin pathway actual/normal
C3847382|T201|COMP|74521-6|LNC|Complement total hemolytic CH50 actual/normal|Complement total hemolytic CH50 actual/normal
C3847383|T201|COMP|74520-8|LNC|Complement alternate pathway AH50 actual/normal|Complement alternate pathway AH50 actual/normal
C3847384|T201|COMP|74519-0|LNC|Complement activity panel|Complement activity panel
C3847385|T201|COMP|74518-2|LNC|Clara cell protein 16|Clara cell protein 16
C3847386|T201|COMP|74517-4|LNC|Cholesterol sulfate|Cholesterol sulfate
C3847387|T201|COMP|74516-6|LNC|Calcium|Calcium
C3847388|T201|COMP|74515-8|LNC|Bile acid|Bile acid
C3847389|T201|COMP|74514-1|LNC|Amino acids panel|Amino acids panel
C3847390|T201|COMP|74513-3|LNC|Alpha tocopherol|Alpha tocopherol
C3847391|T201|COMP|74512-5|LNC|Chemokine (C-C motif) ligand 18|Chemokine (C-C motif) ligand 18
C3847392|T201|COMP|74511-7|LNC|COMT gene.c.1947G>A|COMT gene.c.1947G>A
C3847393|T201|COMP|74510-9|LNC|3-Hydroxyeicosanoylcarnitine (C20-OH)|3-Hydroxyeicosanoylcarnitine (C20-OH)
C3847394|T201|COMP|74509-1|LNC|3-Hydroxydecanoylcarnitine (C10-OH)|3-Hydroxydecanoylcarnitine (C10-OH)
C3847395|T201|COMP|74508-3|LNC|16-Alpha hydroxypregnenolone|16-Alpha hydroxypregnenolone
C3847396|T201|COMP|74507-5|LNC|16-Alpha hydroxypregnenolone|16-Alpha hydroxypregnenolone
C3847397|T201|COMP|74506-7|LNC|16-Alpha hydroxypregnenolone|16-Alpha hydroxypregnenolone
C3847398|T201|COMP|74505-9|LNC|16-Beta,18-dihydroxydehydroepiandrosterone|16-Beta,18-dihydroxydehydroepiandrosterone
C3847399|T201|COMP|74504-2|LNC|16-Beta,18-dihydroxydehydroepiandrosterone|16-Beta,18-dihydroxydehydroepiandrosterone
C3847400|T201|COMP|74503-4|LNC|16-Beta,18-dihydroxydehydroepiandrosterone|16-Beta,18-dihydroxydehydroepiandrosterone
C3847406|T201|COMP|74494-6|LNC|CD34 & Coagulation factor XIII Ag|CD34 & Coagulation factor XIII Ag
C3847408|T201|COMP|74487-0|LNC|P504S & p63 & Cytokeratin 903 Ag|P504S & p63 & Cytokeratin 903 Ag
C3847409|T201|COMP|74486-2|LNC|Cytokeratin 5 & p63 & Cytokeratin AE1 Ag|Cytokeratin 5 & p63 & Cytokeratin AE1 Ag
C3847410|T201|COMP|74485-4|LNC|CD3 & CD20 Ag|CD3 & CD20 Ag
C3847411|T201|COMP|75143-8|LNC|Deoxyuridine|Deoxyuridine
C3847412|T201|COMP|75142-0|LNC|Adenosine|Adenosine
C3847413|T201|COMP|75141-2|LNC|Acadesine|Acadesine
C3847414|T201|COMP|75140-4|LNC|Allantoine|Allantoine
C3847415|T201|COMP|75139-6|LNC|Urate|Urate
C3847417|T201|COMP|75029-9|LNC|Zanamivir|Zanamivir
C3847418|T201|COMP|75028-1|LNC|Protoporphyrin/Porphyrins.total|Protoporphyrin/Porphyrins.total
C3847419|T201|COMP|74809-5|LNC|von Willebrand factor.activity actual/Normal|von Willebrand factor.activity actual/Normal
C3847421|T201|COMP|74807-9|LNC|Transferrin receptor.soluble/log Ferritin index|Transferrin receptor.soluble/log Ferritin index
C3847422|T201|COMP|74806-1|LNC|Lithium^trough|Lithium^trough
C3847430|T201|COMP|74493-8|LNC|PAX5 & CD5 Ag|PAX5 & CD5 Ag
C3847431|T201|COMP|74491-2|LNC|Cytokeratin 7 & Thyroid transcription factor 1 Ag|Cytokeratin 7 & Thyroid transcription factor 1 Ag
C3847432|T201|COMP|74490-4|LNC|PAX5 & BCL2 Ag|PAX5 & BCL2 Ag
C3847433|T201|COMP|74489-6|LNC|Melan-A & Ki67 Ag|Melan-A & Ki67 Ag
C3847434|T201|COMP|74853-3|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C3847435|T201|COMP|74852-5|LNC|Mesothelial cells/100 cells|Mesothelial cells/100 cells
C3847436|T201|COMP|74851-7|LNC|Blasts/100 cells|Blasts/100 cells
C3847437|T201|COMP|74849-1|LNC|Plasma cells/100 cells|Plasma cells/100 cells
C3847438|T201|COMP|74848-3|LNC|Lymphocytes/100 cells|Lymphocytes/100 cells
C3847439|T201|COMP|74847-5|LNC|Toxoplasma gondii Ab.IgE|Toxoplasma gondii Ab.IgE
C3847440|T201|COMP|74644-6|LNC|HYDROcodone|HYDROcodone
C3847441|T201|COMP|74643-8|LNC|Aromatic solvents|Aromatic solvents
C3847442|T201|COMP|74642-0|LNC|1,3-Dichlorobenzene|1,3-Dichlorobenzene
C3847443|T201|COMP|74641-2|LNC|Monoclonal band 2 observed|Monoclonal band 2 observed
C3847444|T201|COMP|74576-0|LNC|Tripeptidyl peptidase I|Tripeptidyl peptidase I
C3847445|T201|COMP|74575-2|LNC|Pyruvate dehydrogenase E1|Pyruvate dehydrogenase E1
C3847446|T201|COMP|74574-5|LNC|Macroscopic observation|Macroscopic observation
C3847466|T201|COMP|75037-2|LNC|2-Hydroxyglutarate|2-Hydroxyglutarate
C3847467|T201|COMP|75036-4|LNC|2-Hydroxyglutarate|2-Hydroxyglutarate
C3847468|T201|COMP|75035-6|LNC|Oxytocin|Oxytocin
C3847469|T201|COMP|75034-9|LNC|NPM1 gene targeted mutation analysis|NPM1 gene targeted mutation analysis
C3847470|T201|COMP|75033-1|LNC|MPL gene mutations tested for|MPL gene mutations tested for
C3847471|T201|COMP|75032-3|LNC|CEBPA gene full mutation analysis|CEBPA gene full mutation analysis
C3853549|T201|COMP|3508-9|LNC|Codeine|Codeine
C3853700|T201|COMP|40570-4|LNC|Blasts|Blasts
C3853701|T201|COMP|19233-6|LNC|Bicarbonate^^standard|Bicarbonate^^standard
C3853749|T201|COMP|34722-9|LNC|EGR2 gene targeted mutation analysis|EGR2 gene targeted mutation analysis
C3853765|T201|COMP|41110-8|LNC|CSTB gene targeted mutation analysis|CSTB gene targeted mutation analysis
C3853766|T201|COMP|39018-7|LNC|Coliform bacteria|Coliform bacteria
C3853768|T201|COMP|12286-1|LNC|Drugs identified|Drugs identified
C3853769|T201|COMP|59022-4|LNC|HLA-DRB3|HLA-DRB3
C3853782|T201|COMP|41112-4|LNC|CMT axonal gene targeted mutation analysis|CMT axonal gene targeted mutation analysis
C3853783|T201|COMP|41117-3|LNC|AS+PWS gene targeted mutation analysis|AS+PWS gene targeted mutation analysis
C3853785|T201|COMP|41120-7|LNC|ALDOB gene targeted mutation analysis|ALDOB gene targeted mutation analysis
C3853853|T201|COMP|56656-2|LNC|Fluoride/Creatinine|Fluoride/Creatinine
C3853963|T201|COMP|75574-4|LNC|22q11.2 deletion prior risk|22q11.2 deletion prior risk
C3853964|T201|COMP|75568-6|LNC|Monosomy X prior risk|Monosomy X prior risk
C3853965|T201|COMP|75566-0|LNC|Monosomy X prior risk|Monosomy X prior risk
C3853966|T201|COMP|75546-2|LNC|Trisomy 13 prior risk|Trisomy 13 prior risk
C3853967|T201|COMP|75550-4|LNC|Trisomy 13 prior risk|Trisomy 13 prior risk
C3853968|T201|COMP|75556-1|LNC|Trisomy 18 prior risk|Trisomy 18 prior risk
C3853969|T201|COMP|75554-6|LNC|Trisomy 18 prior risk|Trisomy 18 prior risk
C3853970|T201|COMP|75562-9|LNC|Trisomy 21 prior risk|Trisomy 21 prior risk
C3853971|T201|COMP|75560-3|LNC|Trisomy 21 prior risk|Trisomy 21 prior risk
C3853983|T201|COMP|75888-8|LNC|HCV RNA screening tests - Meaningful Use set|HCV RNA screening tests - Meaningful Use set
C3854191|T201|COMP|75863-1|LNC|HEDIS 2015-2018 Value Set - Digoxin Level|HEDIS 2015-2018 Value Set - Digoxin Level
C3854194|T201|COMP|75864-9|LNC|HEDIS 2015-2018 Value Set - Glucose Tests|HEDIS 2015-2018 Value Set - Glucose Tests
C3854195|T201|COMP|75862-3|LNC|HEDIS 2015-2020 Value Set - HbA1c Tests|HEDIS 2015-2020 Value Set - HbA1c Tests
C3854197|T201|COMP|75861-5|LNC|HEDIS 2015-2020 Value Set - LDL-C Tests|HEDIS 2015-2020 Value Set - LDL-C Tests
C3854201|T201|COMP|75865-6|LNC|HEDIS 2015-2018 Value Set - PSA Test Exclusion|HEDIS 2015-2018 Value Set - PSA Test Exclusion
C3854203|T201|COMP|75866-4|LNC|HEDIS 2015-2018 Value Set - PSA Tests|HEDIS 2015-2018 Value Set - PSA Tests
C3854205|T201|COMP|75868-0|LNC|HEDIS 2015 Value Sets|HEDIS 2015 Value Sets
C3854207|T201|COMP|75974-6|LNC|KRAS gene targeted mutation analysis|KRAS gene targeted mutation analysis
C3861011|T201|COMP|75599-1|LNC|1p36 deletion prior risk|1p36 deletion prior risk
C3864290|T201|COMP|75575-1|LNC|22q11.2 deletion prior risk|22q11.2 deletion prior risk
C3864940|T201|COMP|75598-3|LNC|1p36 deletion prior risk|1p36 deletion prior risk
C3864941|T201|COMP|75711-2|LNC|Date of autopsy|Date of autopsy
C3869944|T201|COMP|76090-0|LNC|Erythrocytes.hyperchromic/100 erythrocytes|Erythrocytes.hyperchromic/100 erythrocytes
C3869945|T201|COMP|76089-2|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C3869946|T201|COMP|76088-4|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C3869947|T201|COMP|76087-6|LNC|Parainfluenza virus 4 RNA|Parainfluenza virus 4 RNA
C3869948|T201|COMP|76086-8|LNC|Parainfluenza virus 3 RNA|Parainfluenza virus 3 RNA
C3869949|T201|COMP|76085-0|LNC|Parainfluenza virus 2 RNA|Parainfluenza virus 2 RNA
C3869950|T201|COMP|76084-3|LNC|Parainfluenza virus 1 RNA|Parainfluenza virus 1 RNA
C3869954|T201|COMP|76080-1|LNC|Influenza virus B RNA|Influenza virus B RNA
C3869955|T201|COMP|76079-3|LNC|Influenza virus B RNA|Influenza virus B RNA
C3869956|T201|COMP|76078-5|LNC|Influenza virus A RNA|Influenza virus A RNA
C3869957|T201|COMP|76077-7|LNC|Influenza virus A RNA|Influenza virus A RNA
C3869958|T201|COMP|76076-9|LNC|Haemophilus ducreyi DNA|Haemophilus ducreyi DNA
C3869959|T201|COMP|76075-1|LNC|Galactomannan Ag|Galactomannan Ag
C3869960|T201|COMP|76074-4|LNC|Enterovirus RNA|Enterovirus RNA
C3869961|T201|COMP|76073-6|LNC|Fungus identified|Fungus identified
C3869962|T201|COMP|76072-8|LNC|Enterovirus D68 RNA|Enterovirus D68 RNA
C3869963|T201|COMP|76071-0|LNC|Aspergillus sp DNA|Aspergillus sp DNA
C3869964|T201|COMP|76070-2|LNC|Adenovirus DNA|Adenovirus DNA
C3869965|T201|COMP|76069-4|LNC|Erythrocytes.hypochromic/100 erythrocytes|Erythrocytes.hypochromic/100 erythrocytes
C3869966|T201|COMP|76068-6|LNC|MBL2 gene targeted mutation analysis|MBL2 gene targeted mutation analysis
C3869972|T201|COMP|76062-9|LNC|Schistocytes/100 cells|Schistocytes/100 cells
C3869975|T201|COMP|76045-4|LNC|Moxifloxacin 2.0 ug/mL|Moxifloxacin 2.0 ug/mL
C3869976|T201|COMP|76044-7|LNC|Moxifloxacin 1.0 ug/mL|Moxifloxacin 1.0 ug/mL
C3869977|T201|COMP|76043-9|LNC|Moxifloxacin 0.5 ug/mL|Moxifloxacin 0.5 ug/mL
C3869978|T201|COMP|76042-1|LNC|levoFLOXacin 4.0 ug/mL|levoFLOXacin 4.0 ug/mL
C3869979|T201|COMP|76041-3|LNC|levoFLOXacin 2.0 ug/mL|levoFLOXacin 2.0 ug/mL
C3869980|T201|COMP|76040-5|LNC|levoFLOXacin 1.0 ug/mL|levoFLOXacin 1.0 ug/mL
C3869981|T201|COMP|76039-7|LNC|Interleukin 2 receptor.soluble|Interleukin 2 receptor.soluble
C3869982|T201|COMP|76038-9|LNC|Tripeptidyl peptidase I|Tripeptidyl peptidase I
C3869983|T201|COMP|76037-1|LNC|GALT gene full mutation analysis|GALT gene full mutation analysis
C3869984|T201|COMP|76036-3|LNC|GLA gene full mutation analysis|GLA gene full mutation analysis
C3869985|T201|COMP|76035-5|LNC|ARSA gene full mutation analysis|ARSA gene full mutation analysis
C3869986|T201|COMP|76034-8|LNC|GAA gene full mutation analysis|GAA gene full mutation analysis
C3869987|T201|COMP|76033-0|LNC|HEXA gene full mutation analysis|HEXA gene full mutation analysis
C3869988|T201|COMP|76032-2|LNC|SGSH gene full mutation analysis|SGSH gene full mutation analysis
C3869989|T201|COMP|76031-4|LNC|NPC1 gene full mutation analysis|NPC1 gene full mutation analysis
C3869990|T201|COMP|76030-6|LNC|IDS gene full mutation analysis|IDS gene full mutation analysis
C3869991|T201|COMP|76029-8|LNC|HEXB gene full mutation analysis|HEXB gene full mutation analysis
C3869992|T201|COMP|76028-0|LNC|IDUA gene full mutation analysis|IDUA gene full mutation analysis
C3869993|T201|COMP|76027-2|LNC|Mannose-6-phosphate isomerase|Mannose-6-phosphate isomerase
C3869994|T201|COMP|76026-4|LNC|Phosphomannomutase 2|Phosphomannomutase 2
C3869995|T201|COMP|76025-6|LNC|Arylsulfatase C|Arylsulfatase C
C3869996|T201|COMP|76024-9|LNC|Sialate/Creatinine|Sialate/Creatinine
C3869997|T201|COMP|76023-1|LNC|N-acetyl-L-aspartate/Creatinine|N-acetyl-L-aspartate/Creatinine
C3869998|T201|COMP|76022-3|LNC|8(9)-Cholestenol|8(9)-Cholestenol
C3869999|T201|COMP|76021-5|LNC|Delta aPTT|Delta aPTT
C3870000|T201|COMP|76020-7|LNC|Delta dRVVT|Delta dRVVT
C3870001|T201|COMP|75983-7|LNC|Fetal chromosome 21 trisomy|Fetal chromosome 21 trisomy
C3870002|T201|COMP|75982-9|LNC|Fetal chromosome 18 trisomy|Fetal chromosome 18 trisomy
C3870003|T201|COMP|75981-1|LNC|Fetal chromosome 13 trisomy|Fetal chromosome 13 trisomy
C3870004|T201|COMP|75980-3|LNC|Fetal chromosome 13+18+21+X+Y aneuploidy|Fetal chromosome 13+18+21+X+Y aneuploidy
C3870005|T201|COMP|75979-5|LNC|Fetal chromosome 13 trisomy|Fetal chromosome 13 trisomy
C3870006|T201|COMP|75978-7|LNC|Fetal chromosome 18 trisomy|Fetal chromosome 18 trisomy
C3870007|T201|COMP|75977-9|LNC|Fetal chromosome X & Y aneuploidy|Fetal chromosome X & Y aneuploidy
C3870008|T201|COMP|75976-1|LNC|Fetal chromosome 21 trisomy|Fetal chromosome 21 trisomy
C3870009|T201|COMP|75975-3|LNC|Fetal chromosome 13+18+21 trisomy|Fetal chromosome 13+18+21 trisomy
C3870010|T201|COMP|75913-4|LNC|dRVVT.hexagonal phase phospholipid actual/Normal|dRVVT.hexagonal phase phospholipid actual/Normal
C3870034|T201|COMP|75887-0|LNC|HCV antibody RIBA tests - Meaningful Use set|HCV antibody RIBA tests - Meaningful Use set
C3870035|T201|COMP|75886-2|LNC|HCV antibody screening tests - Meaningful Use set|HCV antibody screening tests - Meaningful Use set
C3870037|T201|COMP|75883-9|LNC|dRVVT.hexagonal phase phospholipid|dRVVT.hexagonal phase phospholipid
C3870040|T201|COMP|75880-5|LNC|14-3-3 eta Ag|14-3-3 eta Ag
C3870050|T201|COMP|75860-7|LNC|Hepatitis A virus RNA & Parvovirus B19 DNA panel|Hepatitis A virus RNA & Parvovirus B19 DNA panel
C3870051|T201|COMP|75858-1|LNC|Sterols panel|Sterols panel
C3870089|T201|COMP|75819-3|LNC|Erythrocyte chromasia|Erythrocyte chromasia
C3870094|T201|COMP|75811-0|LNC|Antipsychotics|Antipsychotics
C3870128|T201|COMP|75771-6|LNC|Trifluoperazine|Trifluoperazine
C3870129|T201|COMP|75770-8|LNC|Thioridazine|Thioridazine
C3870130|T201|COMP|75769-0|LNC|Promazine|Promazine
C3870131|T201|COMP|75768-2|LNC|Prochlorperazine|Prochlorperazine
C3870132|T201|COMP|75767-4|LNC|Mesoridazine|Mesoridazine
C3870133|T201|COMP|75766-6|LNC|fluPHENAZine|fluPHENAZine
C3870134|T201|COMP|75765-8|LNC|Triprolidine|Triprolidine
C3870135|T201|COMP|75764-1|LNC|Tripelennamine|Tripelennamine
C3870136|T201|COMP|75763-3|LNC|Orphenadrine|Orphenadrine
C3870137|T201|COMP|75762-5|LNC|Methapyrilene|Methapyrilene
C3870138|T201|COMP|75761-7|LNC|Doxylamine|Doxylamine
C3870139|T201|COMP|75760-9|LNC|Haloperidol|Haloperidol
C3870140|T201|COMP|75759-1|LNC|Chlorpheniramine|Chlorpheniramine
C3870141|T201|COMP|75758-3|LNC|Brompheniramine|Brompheniramine
C3870142|T201|COMP|75757-5|LNC|Chlamydia sp Ab|Chlamydia sp Ab
C3870143|T201|COMP|75756-7|LNC|Bacteria identified|Bacteria identified
C3870144|T201|COMP|75755-9|LNC|Staphylococcus aureus.methicillin susceptible DNA|Staphylococcus aureus.methicillin susceptible DNA
C3870145|T201|COMP|75754-2|LNC|Streptobacillus moniliformis DNA|Streptobacillus moniliformis DNA
C3870146|T201|COMP|75753-4|LNC|Bacterial vancomycin resistance vanD gene|Bacterial vancomycin resistance vanD gene
C3870156|T201|COMP|75741-9|LNC|Beta sitosterol|Beta sitosterol
C3870157|T201|COMP|75740-1|LNC|Lathosterol|Lathosterol
C3870158|T201|COMP|75739-3|LNC|Desmosterol|Desmosterol
C3870159|T201|COMP|75738-5|LNC|Campesterol|Campesterol
C3870160|T201|COMP|75737-7|LNC|Lysophosphatidylcholine(18:0)|Lysophosphatidylcholine(18:0)
C3870161|T201|COMP|75736-9|LNC|Lysophosphatidylcholine(16:0)|Lysophosphatidylcholine(16:0)
C3870165|T201|COMP|75732-8|LNC|HTR2C gene.c.-759C>T|HTR2C gene.c.-759C>T
C3870166|T201|COMP|75731-0|LNC|HTR2A gene.c.102T>C|HTR2A gene.c.102T>C
C3870167|T201|COMP|75725-2|LNC|CYP1A2 gene.c.-729C>T|CYP1A2 gene.c.-729C>T
C3870168|T201|COMP|75724-5|LNC|CYP1A2 gene.c.558C>A|CYP1A2 gene.c.558C>A
C3870169|T201|COMP|75723-7|LNC|CYP1A2 gene.c.2385G>A|CYP1A2 gene.c.2385G>A
C3870170|T201|COMP|75722-9|LNC|CYP1A2 gene.c.-163C>A|CYP1A2 gene.c.-163C>A
C3870171|T201|COMP|75721-1|LNC|CYP1A2 gene.c.5166G>A|CYP1A2 gene.c.5166G>A
C3870172|T201|COMP|75720-3|LNC|CYP1A2 gene.c.5090C>T|CYP1A2 gene.c.5090C>T
C3870173|T201|COMP|75719-5|LNC|CYP1A2 gene.c.-3860G>A|CYP1A2 gene.c.-3860G>A
C3870174|T201|COMP|75718-7|LNC|CYP1A2 gene.c.3533G>A|CYP1A2 gene.c.3533G>A
C3870175|T201|COMP|75717-9|LNC|CYP1A2 gene.c.3497G>A|CYP1A2 gene.c.3497G>A
C3870176|T201|COMP|75716-1|LNC|CYP1A2 gene.c.2499A>T|CYP1A2 gene.c.2499A>T
C3870177|T201|COMP|75715-3|LNC|CYP1A2 gene.c.2473G>A|CYP1A2 gene.c.2473G>A
C3870178|T201|COMP|75714-6|LNC|CYP1A2 gene.c.-2467delT|CYP1A2 gene.c.-2467delT
C3870179|T201|COMP|75713-8|LNC|CYP1A2 gene.c.125C>G|CYP1A2 gene.c.125C>G
C3870180|T201|COMP|75712-0|LNC|Microscopic description|Microscopic description
C3870181|T201|COMP|75710-4|LNC|Coccidioides immitis+posadasii Ab.IgM|Coccidioides immitis+posadasii Ab.IgM
C3870182|T201|COMP|75709-6|LNC|Calcitonin|Calcitonin
C3870183|T201|COMP|75708-8|LNC|Bruton tyrosine kinase|Bruton tyrosine kinase
C3870194|T201|COMP|75697-3|LNC|Bilirubin fractions panel|Bilirubin fractions panel
C3870196|T201|COMP|75695-7|LNC|Human papilloma virus 18 DNA|Human papilloma virus 18 DNA
C3870197|T201|COMP|75694-0|LNC|Human papilloma virus 18+45 E6+E7 mRNA|Human papilloma virus 18+45 E6+E7 mRNA
C3870198|T201|COMP|75693-2|LNC|Fetal sex|Fetal sex
C3870200|T201|COMP|75690-8|LNC|Enterococcus faecium hsp60 gene|Enterococcus faecium hsp60 gene
C3870201|T201|COMP|75689-0|LNC|Iron panel|Iron panel
C3870202|T201|COMP|75688-2|LNC|Gram negative bacteria identified|Gram negative bacteria identified
C3870203|T201|COMP|75684-1|LNC|Bacterial carbapenem resistance blaNDM gene|Bacterial carbapenem resistance blaNDM gene
C3870204|T201|COMP|75683-3|LNC|Bacterial carbapenem resistance blaKPC gene|Bacterial carbapenem resistance blaKPC gene
C3870206|T201|COMP|75681-7|LNC|Pseudomonas aeruginosa (sodA) gene|Pseudomonas aeruginosa (sodA) gene
C3870207|T201|COMP|75680-9|LNC|Klebsiella oxytoca (ompA) gene|Klebsiella oxytoca (ompA) gene
C3870208|T201|COMP|75679-1|LNC|Klebsiella pneumoniae yggE gene|Klebsiella pneumoniae yggE gene
C3870209|T201|COMP|75678-3|LNC|Escherichia coli (oppA) gene|Escherichia coli (oppA) gene
C3870210|T201|COMP|75677-5|LNC|Proteus sp (atpD) gene|Proteus sp (atpD) gene
C3870211|T201|COMP|75676-7|LNC|Enterobacter sp (gyrB+metB) genes|Enterobacter sp (gyrB+metB) genes
C3870212|T201|COMP|75675-9|LNC|Citrobacter sp (ompA+mrkC) genes|Citrobacter sp (ompA+mrkC) genes
C3870213|T201|COMP|75674-2|LNC|Acinetobacter sp (rpsA) gene|Acinetobacter sp (rpsA) gene
C3870214|T201|COMP|75673-4|LNC|Gram negative blood culture panel|Gram negative blood culture panel
C3870219|T201|COMP|75668-4|LNC|Fetal sex|Fetal sex
C3870220|T201|COMP|75667-6|LNC|Electrolytes 3 panel|Electrolytes 3 panel
C3870221|T201|COMP|75666-8|LNC|HIV 1+2 Ab & HIV1 p24 Ag|HIV 1+2 Ab & HIV1 p24 Ag
C3870222|T201|COMP|75665-0|LNC|Ova & parasites identified|Ova & parasites identified
C3870223|T201|COMP|75664-3|LNC|Human papilloma virus 16 DNA|Human papilloma virus 16 DNA
C3870224|T201|COMP|75663-5|LNC|Prolymphocytes|Prolymphocytes
C3870225|T201|COMP|75662-7|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C3870226|T201|COMP|75661-9|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C3870227|T201|COMP|75660-1|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C3870228|T201|COMP|75659-3|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C3870229|T201|COMP|75658-5|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C3870230|T201|COMP|75657-7|LNC|Mononuclear cells|Mononuclear cells
C3870231|T201|COMP|75656-9|LNC|Mononuclear cells|Mononuclear cells
C3870232|T201|COMP|75650-2|LNC|Sulfonamide|Sulfonamide
C3870233|T201|COMP|75649-4|LNC|Mitragynine+7-Hydroxymitragynine|Mitragynine+7-Hydroxymitragynine
C3870234|T201|COMP|75643-7|LNC|7-Hydroxymitragynine|7-Hydroxymitragynine
C3870235|T201|COMP|75642-9|LNC|Urate/Creatinine|Urate/Creatinine
C3870236|T201|COMP|75641-1|LNC|Electrolytes 3 panel|Electrolytes 3 panel
C3870237|T201|COMP|75640-3|LNC|Lysozyme|Lysozyme
C3870239|T201|COMP|75638-7|LNC|Homocarnosine|Homocarnosine
C3870240|T201|COMP|75637-9|LNC|Glucose^45M post 50 g lactose PO|Glucose^45M post 50 g lactose PO
C3870242|T201|COMP|75635-3|LNC|Rheumatoid arthritis disease activity panel|Rheumatoid arthritis disease activity panel
C3870243|T201|COMP|75634-6|LNC|Rheumatoid arthritis disease activity score level|Rheumatoid arthritis disease activity score level
C3870244|T201|COMP|75633-8|LNC|Rheumatoid arthritis disease activity score|Rheumatoid arthritis disease activity score
C3870245|T201|COMP|75632-0|LNC|Resistin|Resistin
C3870246|T201|COMP|75631-2|LNC|Stromelysin-1|Stromelysin-1
C3870247|T201|COMP|75630-4|LNC|Interstitial collagenase|Interstitial collagenase
C3870249|T201|COMP|75628-8|LNC|Vascular endothelial growth factor A|Vascular endothelial growth factor A
C3870250|T201|COMP|75627-0|LNC|Vascular cell adhesion molecule 1|Vascular cell adhesion molecule 1
C3870253|T201|COMP|75622-1|LNC|HIV 1 & 2 tests - Meaningful Use set|HIV 1 & 2 tests - Meaningful Use set
C3870263|T201|COMP|75608-0|LNC|Citation|Citation
C3870264|T201|COMP|75607-2|LNC|Paternal sample received|Paternal sample received
C3870265|T201|COMP|75606-4|LNC|Cell-free DNA.fetal/Cell-free DNA.total|Cell-free DNA.fetal/Cell-free DNA.total
C3870266|T201|COMP|75605-6|LNC|Cell-free DNA.fetal/Cell-free DNA.total|Cell-free DNA.fetal/Cell-free DNA.total
C3870267|T201|COMP|75604-9|LNC|Fetal sex|Fetal sex
C3870269|T201|COMP|75602-3|LNC|Fetal 1p36 deletion risk|Fetal 1p36 deletion risk
C3870270|T201|COMP|75601-5|LNC|Fetal 1p36 deletion risk|Fetal 1p36 deletion risk
C3870271|T201|COMP|75600-7|LNC|Fetal 1p36 deletion risk|Fetal 1p36 deletion risk
C3870273|T201|COMP|75596-7|LNC|Fetal 5p deletion risk|Fetal 5p deletion risk
C3870274|T201|COMP|75595-9|LNC|Fetal 5p deletion risk|Fetal 5p deletion risk
C3870275|T201|COMP|75594-2|LNC|Fetal 5p deletion risk|Fetal 5p deletion risk
C3870276|T201|COMP|75593-4|LNC|5p deletion prior risk|5p deletion prior risk
C3870277|T201|COMP|75592-6|LNC|5p deletion prior risk|5p deletion prior risk
C3870279|T201|COMP|75590-0|LNC|Fetal Angelman syndrome risk|Fetal Angelman syndrome risk
C3870280|T201|COMP|75589-2|LNC|Fetal Angelman syndrome risk|Fetal Angelman syndrome risk
C3870281|T201|COMP|75588-4|LNC|Fetal Angelman syndrome risk|Fetal Angelman syndrome risk
C3870282|T201|COMP|75587-6|LNC|Angelman syndrome prior risk|Angelman syndrome prior risk
C3870283|T201|COMP|75586-8|LNC|Angelman syndrome prior risk|Angelman syndrome prior risk
C3870285|T201|COMP|75584-3|LNC|Fetal Prader-Willi syndrome risk|Fetal Prader-Willi syndrome risk
C3870287|T201|COMP|75647-8|LNC|Meperidine|Meperidine
C3870288|T201|COMP|75646-0|LNC|Ethylene glycol|Ethylene glycol
C3870289|T201|COMP|75645-2|LNC|Butabarbital|Butabarbital
C3870290|T201|COMP|75644-5|LNC|Amphetamine+Methamphetamine|Amphetamine+Methamphetamine
C3870291|T201|COMP|75583-5|LNC|Fetal Prader-Willi syndrome risk|Fetal Prader-Willi syndrome risk
C3870292|T201|COMP|75582-7|LNC|Fetal Prader-Willi syndrome risk|Fetal Prader-Willi syndrome risk
C3870293|T201|COMP|75581-9|LNC|Prader-Willi syndrome prior risk|Prader-Willi syndrome prior risk
C3870294|T201|COMP|75580-1|LNC|Prader-Willi syndrome prior risk|Prader-Willi syndrome prior risk
C3870296|T201|COMP|75578-5|LNC|Fetal 22q11.2 deletion risk|Fetal 22q11.2 deletion risk
C3870297|T201|COMP|75577-7|LNC|Fetal 22q11.2 deletion risk|Fetal 22q11.2 deletion risk
C3870298|T201|COMP|75576-9|LNC|Fetal 22q11.2 deletion risk|Fetal 22q11.2 deletion risk
C3870299|T201|COMP|75573-6|LNC|Genetic counselor comment on fetal Triploidy risk|Genetic counselor comment on fetal Triploidy risk
C3870300|T201|COMP|75572-8|LNC|Fetal triploidy risk|Fetal triploidy risk
C3870302|T201|COMP|75570-2|LNC|Fetal monosomy X risk|Fetal monosomy X risk
C3870303|T201|COMP|75569-4|LNC|Fetal monosomy X risk|Fetal monosomy X risk
C3870304|T201|COMP|75567-8|LNC|Fetal monosomy X risk|Fetal monosomy X risk
C3870306|T201|COMP|75564-5|LNC|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3870307|T201|COMP|75563-7|LNC|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3870308|T201|COMP|75561-1|LNC|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3870310|T201|COMP|75558-7|LNC|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3870311|T201|COMP|75557-9|LNC|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3870312|T201|COMP|75555-3|LNC|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3870314|T201|COMP|75552-0|LNC|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3870315|T201|COMP|75551-2|LNC|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3870317|T201|COMP|75548-8|LNC|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3870320|T201|COMP|75540-5|LNC|Hepatitis A virus RNA+Parvovirus B19 DNA|Hepatitis A virus RNA+Parvovirus B19 DNA
C3870335|T201|COMP|75518-1|LNC|Bacteria identified|Bacteria identified
C3870336|T201|COMP|75517-3|LNC|Protein.monoclonal band 4|Protein.monoclonal band 4
C3870337|T201|COMP|75516-5|LNC|Cortisol.free|Cortisol.free
C3870339|T201|COMP|75514-0|LNC|Lupus anticoagulant two screening tests W Reflex|Lupus anticoagulant two screening tests W Reflex
C3870340|T201|COMP|75513-2|LNC|DRVVT with 1:1 Pooled Normal Plasma|DRVVT with 1:1 Pooled Normal Plasma
C3870341|T201|COMP|75512-4|LNC|DRVVT with 1:1 Pooled Normal Plasma actual/Normal|DRVVT with 1:1 Pooled Normal Plasma actual/Normal
C3870342|T201|COMP|75511-6|LNC|DRVVT percent correction|DRVVT percent correction
C3870418|T201|COMP|75411-9|LNC|Ebola Zaire virus RNA|Ebola Zaire virus RNA
C3870419|T201|COMP|75410-1|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C3870420|T201|COMP|75409-3|LNC|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C3870421|T201|COMP|75408-5|LNC|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C3870422|T201|COMP|75402-8|LNC|GCDH gene targeted mutation analysis|GCDH gene targeted mutation analysis
C3870423|T201|COMP|75401-0|LNC|GCDH gene full mutation analysis|GCDH gene full mutation analysis
C3870424|T201|COMP|75400-2|LNC|KCNJ11 gene full mutation analysis|KCNJ11 gene full mutation analysis
C3870425|T201|COMP|75399-6|LNC|HNF4A gene full mutation analysis|HNF4A gene full mutation analysis
C3870426|T201|COMP|75398-8|LNC|HNF1B gene full mutation analysis|HNF1B gene full mutation analysis
C3870427|T201|COMP|75397-0|LNC|HNF1A gene full mutation analysis|HNF1A gene full mutation analysis
C3870429|T201|COMP|75395-4|LNC|AIP gene full mutation analysis|AIP gene full mutation analysis
C3870430|T201|COMP|75394-7|LNC|Chromosome uniparental disomy|Chromosome uniparental disomy
C3870431|T201|COMP|75393-9|LNC|HTT gene.CAG repeats|HTT gene.CAG repeats
C3870432|T201|COMP|75392-1|LNC|FXN gene.GAA repeats|FXN gene.GAA repeats
C3870433|T201|COMP|75391-3|LNC|FGFR3 gene targeted mutation analysis|FGFR3 gene targeted mutation analysis
C3870434|T201|COMP|75390-5|LNC|APP gene targeted mutation analysis|APP gene targeted mutation analysis
C3870435|T201|COMP|75389-7|LNC|CDKN1B gene full mutation analysis|CDKN1B gene full mutation analysis
C3870436|T201|COMP|75383-0|LNC|DMD gene deletion+duplication|DMD gene deletion+duplication
C3870439|T201|COMP|75380-6|LNC|SERPING1 gene targeted mutation analysis|SERPING1 gene targeted mutation analysis
C3870440|T201|COMP|75379-8|LNC|Norbuprenorphine|Norbuprenorphine
C3870441|T201|COMP|75378-0|LNC|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C3870442|T201|COMP|75377-2|LNC|Dengue virus NS1 Ag|Dengue virus NS1 Ag
C3870443|T201|COMP|75376-4|LNC|Siderocytes.HPF|Siderocytes.HPF
C3870444|T201|COMP|75375-6|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C3870445|T201|COMP|75370-7|LNC|Norbuprenorphine|Norbuprenorphine
C3870446|T201|COMP|75369-9|LNC|Diuretics|Diuretics
C3870447|T201|COMP|75368-1|LNC|Buprenorphine|Buprenorphine
C3870448|T201|COMP|75367-3|LNC|Buprenorphine|Buprenorphine
C3870449|T201|COMP|75366-5|LNC|Lactate|Lactate
C3870451|T201|COMP|75364-0|LNC|Urea|Urea
C3870452|T201|COMP|75363-2|LNC|Creatinine|Creatinine
C3870453|T201|COMP|75362-4|LNC|Tapentadol glucuronide|Tapentadol glucuronide
C3870454|T201|COMP|75359-0|LNC|Bacteria identified|Bacteria identified
C3870455|T201|COMP|75358-2|LNC|Bacteria identified|Bacteria identified
C3870456|T201|COMP|75357-4|LNC|Bacteria identified|Bacteria identified
C3870457|T201|COMP|75356-6|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C3870458|T201|COMP|75355-8|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C3870459|T201|COMP|75354-1|LNC|Other cells|Other cells
C3870460|T201|COMP|75353-3|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C3870461|T201|COMP|75352-5|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C3870462|T201|COMP|75351-7|LNC|Other cells|Other cells
C3870463|T201|COMP|75350-9|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C3870464|T201|COMP|75349-1|LNC|Other cells|Other cells
C3870465|T201|COMP|75347-5|LNC|Tapentadol|Tapentadol
C3870466|T201|COMP|75346-7|LNC|Promethazine|Promethazine
C3870490|T201|COMP|75308-7|LNC|Fetal blood|Fetal blood
C3870510|T201|COMP|75271-7|LNC|Other cells/100 cells|Other cells/100 cells
C3870511|T201|COMP|75270-9|LNC|Promethazine|Promethazine
C3870520|T201|COMP|75815-1|LNC|Antipsychotics drug panel|Antipsychotics drug panel
C3870521|T201|COMP|75814-4|LNC|Antihistamines panel|Antihistamines panel
C3870522|T201|COMP|75813-6|LNC|Promethazine|Promethazine
C3870523|T201|COMP|75812-8|LNC|Antihistamines|Antihistamines
C3870525|T201|COMP|75543-9|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C3870526|T201|COMP|75542-1|LNC|Hepatitis A virus RNA|Hepatitis A virus RNA
C3870527|T201|COMP|75541-3|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C3870528|T201|COMP|75374-9|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C3870529|T201|COMP|75373-1|LNC|Erythrocytes.fetal/2000 erythrocytes|Erythrocytes.fetal/2000 erythrocytes
C3870530|T201|COMP|75372-3|LNC|Hexane|Hexane
C3870531|T201|COMP|75371-5|LNC|Bartlett score|Bartlett score
C3870532|T201|COMP|75730-2|LNC|HTR2C gene.c.796G>C|HTR2C gene.c.796G>C
C3870533|T201|COMP|75729-4|LNC|HTR2A gene.c.1354C>T|HTR2A gene.c.1354C>T
C3870534|T201|COMP|75728-6|LNC|HTR2A gene.c.74C>A|HTR2A gene.c.74C>A
C3870535|T201|COMP|75727-8|LNC|HTR2A gene.c.IVS2+54538A>G|HTR2A gene.c.IVS2+54538A>G
C3870536|T201|COMP|75726-0|LNC|HTR2A gene.c.-1438G>A|HTR2A gene.c.-1438G>A
C3870537|T201|COMP|75687-4|LNC|Bacterial carbapenem resistance blaOXA gene|Bacterial carbapenem resistance blaOXA gene
C3870538|T201|COMP|75686-6|LNC|Bacterial carbapenem resistance blaIMP gene|Bacterial carbapenem resistance blaIMP gene
C3870539|T201|COMP|75685-8|LNC|Bacterial carbapenem resistance blaVIM gene|Bacterial carbapenem resistance blaVIM gene
C3870540|T201|COMP|75655-1|LNC|Mononuclear cells|Mononuclear cells
C3870541|T201|COMP|75654-4|LNC|Manual differential comment|Manual differential comment
C3870542|T201|COMP|75653-6|LNC|Manual differential comment|Manual differential comment
C3870543|T201|COMP|75652-8|LNC|Lymphocytes.immature|Lymphocytes.immature
C3870544|T201|COMP|75651-0|LNC|Tetrahydrocannabivarin|Tetrahydrocannabivarin
C3870545|T201|COMP|75407-7|LNC|Hepatitis B virus little e Ab|Hepatitis B virus little e Ab
C3870546|T201|COMP|75406-9|LNC|Human papilloma virus 16 & 18+45 E6+E7 mRNA|Human papilloma virus 16 & 18+45 E6+E7 mRNA
C3870547|T201|COMP|75405-1|LNC|Glucose^1.5H post dose triple bolus|Glucose^1.5H post dose triple bolus
C3870548|T201|COMP|75404-4|LNC|West Nile virus Ab|West Nile virus Ab
C3870549|T201|COMP|75403-6|LNC|PDHA1 gene full mutation analysis|PDHA1 gene full mutation analysis
C3870562|T201|COMP|75387-1|LNC|INS gene full mutation analysis|INS gene full mutation analysis
C3870564|T201|COMP|75385-5|LNC|DMD gene deletion+duplication|DMD gene deletion+duplication
C3870565|T201|COMP|75384-8|LNC|PMP22 gene deletion+duplication|PMP22 gene deletion+duplication
C3888327|T201|COMP|77309-3|LNC|Acylcarnitine pattern|Acylcarnitine pattern
C4018866|T201|COMP|77012-3|LNC|Fetal chromosome 18 trisomy|Fetal chromosome 18 trisomy
C4018867|T201|COMP|77011-5|LNC|Fetal chromosome 21 trisomy|Fetal chromosome 21 trisomy
C4018884|T201|COMP|77381-2|LNC|Protein fractions panel|Protein fractions panel
C4019049|T201|COMP|76397-9|LNC|Lymph node involvement|Lymph node involvement
C4019186|T201|COMP|77013-1|LNC|Fetal chromosome 13 trisomy|Fetal chromosome 13 trisomy
C4036469|T201|COMP|77764-9|LNC|Buprenorphine cutoff|Buprenorphine cutoff
C4036471|T201|COMP|76681-6|LNC|Color^3rd tube|Color^3rd tube
C4036476|T201|COMP|76483-7|LNC|Apolipoprotein A-I|Apolipoprotein A-I
C4036477|T201|COMP|76149-4|LNC|Tulathromycin|Tulathromycin
C4036481|T201|COMP|78036-1|LNC|Fibers|Fibers
C4036482|T201|COMP|78035-3|LNC|Fibers|Fibers
C4036493|T201|COMP|78015-5|LNC|HLA-B|HLA-B
C4036494|T201|COMP|78014-8|LNC|HLA-A|HLA-A
C4036495|T201|COMP|78013-0|LNC|HLA-A & B & DRB & DQB1 panel|HLA-A & B & DRB & DQB1 panel
C4036496|T201|COMP|78011-4|LNC|Schistocytes/100 cells|Schistocytes/100 cells
C4036497|T201|COMP|78010-6|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C4036498|T201|COMP|78009-8|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C4036499|T201|COMP|78008-0|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C4036500|T201|COMP|78007-2|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C4036501|T201|COMP|78006-4|LNC|Glomerular filtration rate/1.73 sq M|Glomerular filtration rate/1.73 sq M
C4036503|T201|COMP|78004-9|LNC|Staphylococcus aureus.vancomycin resistance|Staphylococcus aureus.vancomycin resistance
C4036506|T201|COMP|78001-5|LNC|Cytomegalovirus pp65 Ag/100000 PMN cells|Cytomegalovirus pp65 Ag/100000 PMN cells
C4036516|T201|COMP|77964-5|LNC|Cholesterol crystals|Cholesterol crystals
C4036518|T201|COMP|77948-8|LNC|Cells.FLAER/100 cells|Cells.FLAER/100 cells
C4036519|T201|COMP|77947-0|LNC|Cells.CD9/100 cells|Cells.CD9/100 cells
C4036520|T201|COMP|77946-2|LNC|Cells.CD42b/100 cells|Cells.CD42b/100 cells
C4036521|T201|COMP|77945-4|LNC|Cells.CD4+CD3-/100 cells|Cells.CD4+CD3-/100 cells
C4036522|T201|COMP|77944-7|LNC|Cells.CD11a/100 cells|Cells.CD11a/100 cells
C4036523|T201|COMP|77943-9|LNC|Schistosoma mansoni+haematobium+intercalatum|Schistosoma mansoni+haematobium+intercalatum
C4036524|T201|COMP|77942-1|LNC|Cells.CD8+CD3-/100 cells|Cells.CD8+CD3-/100 cells
C4036526|T201|COMP|77940-5|LNC|Albumin|Albumin
C4036527|T201|COMP|77939-7|LNC|Corticotropin^45M post XXX challenge|Corticotropin^45M post XXX challenge
C4036528|T201|COMP|77938-9|LNC|Cortisol^124H post XXX challenge|Cortisol^124H post XXX challenge
C4036529|T201|COMP|77937-1|LNC|Cortisol^12H post XXX challenge|Cortisol^12H post XXX challenge
C4036530|T201|COMP|77936-3|LNC|Cortisol^10.5H post XXX challenge|Cortisol^10.5H post XXX challenge
C4036531|T201|COMP|77935-5|LNC|Cortisol^10H post XXX challenge|Cortisol^10H post XXX challenge
C4036532|T201|COMP|77934-8|LNC|Cortisol^9.5H post XXX challenge|Cortisol^9.5H post XXX challenge
C4036533|T201|COMP|77933-0|LNC|Cortisol^9H post XXX challenge|Cortisol^9H post XXX challenge
C4036534|T201|COMP|77932-2|LNC|Cortisol^8H post XXX challenge|Cortisol^8H post XXX challenge
C4036535|T201|COMP|77931-4|LNC|Cortisol^6H post XXX challenge|Cortisol^6H post XXX challenge
C4036536|T201|COMP|77930-6|LNC|Cortisol^4H post XXX challenge|Cortisol^4H post XXX challenge
C4036537|T201|COMP|77929-8|LNC|Cortisol^3.5H post XXX challenge|Cortisol^3.5H post XXX challenge
C4036538|T201|COMP|77928-0|LNC|Cortisol^75M post XXX challenge|Cortisol^75M post XXX challenge
C4036539|T201|COMP|77927-2|LNC|Cortisol^5M post XXX challenge|Cortisol^5M post XXX challenge
C4036540|T201|COMP|77926-4|LNC|Cortisol^3M post XXX challenge|Cortisol^3M post XXX challenge
C4036541|T201|COMP|77925-6|LNC|Cortisol^10M post XXX challenge|Cortisol^10M post XXX challenge
C4036570|T201|COMP|77888-6|LNC|OLANZapine|OLANZapine
C4036571|T201|COMP|77887-8|LNC|OLANZapine cutoff|OLANZapine cutoff
C4036572|T201|COMP|77886-0|LNC|Nortriptyline cutoff|Nortriptyline cutoff
C4036573|T201|COMP|77885-2|LNC|Ethyl sulfate cutoff|Ethyl sulfate cutoff
C4036574|T201|COMP|77884-5|LNC|Dehydroaripiprazole|Dehydroaripiprazole
C4036575|T201|COMP|77883-7|LNC|QUEtiapine cutoff|QUEtiapine cutoff
C4036576|T201|COMP|77882-9|LNC|Dehydroaripiprazole cutoff|Dehydroaripiprazole cutoff
C4036577|T201|COMP|77881-1|LNC|risperiDONE cutoff|risperiDONE cutoff
C4036578|T201|COMP|77880-3|LNC|risperiDONE|risperiDONE
C4036579|T201|COMP|77879-5|LNC|Tapentadol cutoff|Tapentadol cutoff
C4036580|T201|COMP|77878-7|LNC|Ziprasidone cutoff|Ziprasidone cutoff
C4036581|T201|COMP|77877-9|LNC|Ziprasidone|Ziprasidone
C4036582|T201|COMP|77876-1|LNC|Phencyclidine cutoff|Phencyclidine cutoff
C4036607|T201|COMP|78019-7|LNC|Toscana virus Ab.IgM|Toscana virus Ab.IgM
C4036608|T201|COMP|78018-9|LNC|Toscana virus Ab.IgG|Toscana virus Ab.IgG
C4036609|T201|COMP|78017-1|LNC|HLA-DQB1|HLA-DQB1
C4036610|T201|COMP|78016-3|LNC|HLA-DRB|HLA-DRB
C4036615|T201|COMP|77791-2|LNC|Benzoylecgonine cutoff|Benzoylecgonine cutoff
C4036616|T201|COMP|77790-4|LNC|Cocaine cutoff|Cocaine cutoff
C4036618|T201|COMP|77788-8|LNC|cloZAPine cutoff|cloZAPine cutoff
C4036619|T201|COMP|77787-0|LNC|Buprenorphine cutoff|Buprenorphine cutoff
C4036623|T201|COMP|77781-3|LNC|Pregabalin cutoff|Pregabalin cutoff
C4036624|T201|COMP|77780-5|LNC|oxyMORphone cutoff|oxyMORphone cutoff
C4036625|T201|COMP|77779-7|LNC|Noroxycodone cutoff|Noroxycodone cutoff
C4036626|T201|COMP|77778-9|LNC|Noroxycodone cutoff|Noroxycodone cutoff
C4036627|T201|COMP|77777-1|LNC|Normeperidine cutoff|Normeperidine cutoff
C4036628|T201|COMP|77776-3|LNC|Norhydrocodone cutoff|Norhydrocodone cutoff
C4036629|T201|COMP|77775-5|LNC|Norfentanyl cutoff|Norfentanyl cutoff
C4036630|T201|COMP|77774-8|LNC|Norbuprenorphine cutoff|Norbuprenorphine cutoff
C4036631|T201|COMP|77773-0|LNC|Morphine cutoff|Morphine cutoff
C4036632|T201|COMP|77772-2|LNC|Methylenedioxyethylamphetamine cutoff|Methylenedioxyethylamphetamine cutoff
C4036633|T201|COMP|77771-4|LNC|JWH-081 5-hydroxypentyl|JWH-081 5-hydroxypentyl
C4036634|T201|COMP|77770-6|LNC|HYDROmorphone cutoff|HYDROmorphone cutoff
C4036635|T201|COMP|77769-8|LNC|Ethyl glucuronide cutoff|Ethyl glucuronide cutoff
C4036636|T201|COMP|77768-0|LNC|Ethanol cutoff|Ethanol cutoff
C4036637|T201|COMP|77767-2|LNC|Codeine cutoff|Codeine cutoff
C4036638|T201|COMP|77766-4|LNC|clonazePAM cutoff|clonazePAM cutoff
C4036639|T201|COMP|77765-6|LNC|Citalopram+Escitalopram|Citalopram+Escitalopram
C4036640|T201|COMP|77763-1|LNC|ALPRAZolam cutoff|ALPRAZolam cutoff
C4036641|T201|COMP|77762-3|LNC|Alpha hydroxyalprazolam cutoff|Alpha hydroxyalprazolam cutoff
C4036642|T201|COMP|77761-5|LNC|ARIPiprazole|ARIPiprazole
C4036643|T201|COMP|77760-7|LNC|ARIPiprazole cutoff|ARIPiprazole cutoff
C4036644|T201|COMP|77759-9|LNC|9-Hydroxyrisperidone cutoff|9-Hydroxyrisperidone cutoff
C4036645|T201|COMP|77758-1|LNC|7-Hydroxyquetiapine cutoff|7-Hydroxyquetiapine cutoff
C4036646|T201|COMP|77757-3|LNC|7-Hydroxyquetiapine|7-Hydroxyquetiapine
C4036647|T201|COMP|77756-5|LNC|7-Aminoclonazepam cutoff|7-Aminoclonazepam cutoff
C4036648|T201|COMP|77755-7|LNC|6-Monoacetylmorphine cutoff|6-Monoacetylmorphine cutoff
C4036652|T201|COMP|77751-6|LNC|TMEM216 gene.c.218G>T|TMEM216 gene.c.218G>T
C4036653|T201|COMP|77750-8|LNC|DLD gene targeted mutation analysis|DLD gene targeted mutation analysis
C4036654|T201|COMP|77749-0|LNC|CLRN1 gene.c.144T>G|CLRN1 gene.c.144T>G
C4036655|T201|COMP|77748-2|LNC|PCDH15 gene.c.733C>T|PCDH15 gene.c.733C>T
C4036656|T201|COMP|77747-4|LNC|HTLV II gp46-II Ab|HTLV II gp46-II Ab
C4036657|T201|COMP|77746-6|LNC|HTLV I gp46-I Ab|HTLV I gp46-I Ab
C4036658|T201|COMP|77740-9|LNC|Norcotinine|Norcotinine
C4036659|T201|COMP|77739-1|LNC|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C4036665|T201|COMP|77733-4|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C4036666|T201|COMP|77732-6|LNC|oxyCODONE+oxymorphone|oxyCODONE+oxymorphone
C4036667|T201|COMP|77731-8|LNC|oxyCODONE+oxymorphone|oxyCODONE+oxymorphone
C4036668|T201|COMP|77730-0|LNC|oxyCODONE|oxyCODONE
C4036669|T201|COMP|77729-2|LNC|oxyMORphone|oxyMORphone
C4036671|T201|COMP|77727-6|LNC|XXX allergen basophil bound Ab|XXX allergen basophil bound Ab
C4036710|T201|COMP|77685-6|LNC|HIV 1 & 2 Ab.IgG|HIV 1 & 2 Ab.IgG
C4036711|T201|COMP|77684-9|LNC|Legionella pneumophila 1 Ag|Legionella pneumophila 1 Ag
C4036712|T201|COMP|77683-1|LNC|Thrombin activatable fibrinolysis inhibitor|Thrombin activatable fibrinolysis inhibitor
C4036714|T201|COMP|77681-5|LNC|Glucose^11H post XXX challenge|Glucose^11H post XXX challenge
C4036715|T201|COMP|77680-7|LNC|Renin^4H post XXX challenge|Renin^4H post XXX challenge
C4036718|T201|COMP|77677-3|LNC|Glucose^2H post meal|Glucose^2H post meal
C4036719|T201|COMP|77671-6|LNC|Gastrin^1M post XXX challenge|Gastrin^1M post XXX challenge
C4036720|T201|COMP|77669-0|LNC|Calcitonin^30M post XXX challenge|Calcitonin^30M post XXX challenge
C4036721|T201|COMP|77668-2|LNC|Calcitonin^5M post XXX challenge|Calcitonin^5M post XXX challenge
C4036722|T201|COMP|77667-4|LNC|Calcitonin^2M post XXX challenge|Calcitonin^2M post XXX challenge
C4036723|T201|COMP|77666-6|LNC|Bacterial methicillin resistance mecA mRNA|Bacterial methicillin resistance mecA mRNA
C4036724|T201|COMP|77665-8|LNC|Dexamethasone|Dexamethasone
C4036725|T201|COMP|77664-1|LNC|Aneuploid G1 phase cell population 2 peak channel|Aneuploid G1 phase cell population 2 peak channel
C4036726|T201|COMP|77663-3|LNC|Aneuploid G1 phase cell population peak channel|Aneuploid G1 phase cell population peak channel
C4036727|T201|COMP|77662-5|LNC|Diploid G1 phase cell population peak channel|Diploid G1 phase cell population peak channel
C4036728|T201|COMP|77656-7|LNC|Cells.diploid.S phase/100 cells|Cells.diploid.S phase/100 cells
C4036729|T201|COMP|77649-2|LNC|17-Hydroxyprogesterone^10M post XXX challenge|17-Hydroxyprogesterone^10M post XXX challenge
C4036732|T201|COMP|77646-8|LNC|HLA-DR Ab.IgG|HLA-DR Ab.IgG
C4036733|T201|COMP|77645-0|LNC|HLA-DQ Ab.IgG|HLA-DQ Ab.IgG
C4036734|T201|COMP|77644-3|LNC|HLA-DP Ab.IgG|HLA-DP Ab.IgG
C4036735|T201|COMP|77643-5|LNC|HLA-C Ab.IgG|HLA-C Ab.IgG
C4036736|T201|COMP|77642-7|LNC|HLA-B Ab.IgG|HLA-B Ab.IgG
C4036737|T201|COMP|77641-9|LNC|HLA-A Ab.IgG|HLA-A Ab.IgG
C4036738|T201|COMP|77640-1|LNC|HLA class I & II Ab.IgG|HLA class I & II Ab.IgG
C4036739|T201|COMP|77639-3|LNC|HLA class I & II Ab.IgG panel|HLA class I & II Ab.IgG panel
C4036740|T201|COMP|77638-5|LNC|HLA-DP & DQ & DR (class II) Ab.IgG panel|HLA-DP & DQ & DR (class II) Ab.IgG panel
C4036741|T201|COMP|77637-7|LNC|HLA-A & B & C (class I) Ab.IgG panel|HLA-A & B & C (class I) Ab.IgG panel
C4036742|T201|COMP|77636-9|LNC|HLA-C|HLA-C
C4036743|T201|COMP|77635-1|LNC|C9orf72 gene.GGGGCC repeats|C9orf72 gene.GGGGCC repeats
C4036744|T201|COMP|77634-4|LNC|FUS gene targeted mutation analysis|FUS gene targeted mutation analysis
C4036745|T201|COMP|77633-6|LNC|TARDBP gene targeted mutation analysis|TARDBP gene targeted mutation analysis
C4036746|T201|COMP|77632-8|LNC|ANG gene targeted mutation analysis|ANG gene targeted mutation analysis
C4036747|T201|COMP|77631-0|LNC|VAPB gene targeted mutation analysis|VAPB gene targeted mutation analysis
C4036748|T201|COMP|77630-2|LNC|ALS2 gene targeted mutation analysis|ALS2 gene targeted mutation analysis
C4036749|T201|COMP|77629-4|LNC|PARK7 gene targeted mutation analysis|PARK7 gene targeted mutation analysis
C4036750|T201|COMP|77628-6|LNC|PSEN2 gene targeted mutation analysis|PSEN2 gene targeted mutation analysis
C4036751|T201|COMP|77627-8|LNC|HBB gene full mutation analysis|HBB gene full mutation analysis
C4036752|T201|COMP|77626-0|LNC|Pyruvate kinase|Pyruvate kinase
C4036753|T201|COMP|77625-2|LNC|ENG gene full mutation analysis|ENG gene full mutation analysis
C4036754|T201|COMP|77624-5|LNC|SMAD4 gene full mutation analysis|SMAD4 gene full mutation analysis
C4036755|T201|COMP|77623-7|LNC|Thyrotropin^2.5H post XXX challenge|Thyrotropin^2.5H post XXX challenge
C4036756|T201|COMP|77622-9|LNC|Natriuretic peptide.B prohormone N-Terminal|Natriuretic peptide.B prohormone N-Terminal
C4036757|T201|COMP|77621-1|LNC|Natriuretic peptide.B prohormone N-Terminal|Natriuretic peptide.B prohormone N-Terminal
C4036758|T201|COMP|77620-3|LNC|Arginase-1|Arginase-1
C4036759|T201|COMP|77924-9|LNC|Enterobacteriaceae.carbapenem resistant|Enterobacteriaceae.carbapenem resistant
C4036762|T201|COMP|77619-5|LNC|Fetal chromosome 13+18+21+Y aneuploidy|Fetal chromosome 13+18+21+Y aneuploidy
C4036765|T201|COMP|77616-1|LNC|Liver fibrosis score|Liver fibrosis score
C4036767|T201|COMP|77614-6|LNC|Calcitonin^10M post XXX challenge|Calcitonin^10M post XXX challenge
C4036768|T201|COMP|77613-8|LNC|Calcitonin^1M post XXX challenge|Calcitonin^1M post XXX challenge
C4036769|T201|COMP|77612-0|LNC|C peptide^45M post XXX challenge|C peptide^45M post XXX challenge
C4036770|T201|COMP|77611-2|LNC|C peptide^4H post XXX challenge|C peptide^4H post XXX challenge
C4036771|T201|COMP|77610-4|LNC|C peptide^15M post XXX challenge|C peptide^15M post XXX challenge
C4036772|T201|COMP|77609-6|LNC|Aldosterone^4H post XXX challenge|Aldosterone^4H post XXX challenge
C4036788|T201|COMP|77563-5|LNC|Leukocyte esterase|Leukocyte esterase
C4036853|T201|COMP|77496-8|LNC|Clostridium perfringens|Clostridium perfringens
C4036854|T201|COMP|77495-0|LNC|Bacillus cereus|Bacillus cereus
C4036885|T201|COMP|77452-1|LNC|Bilirubin|Bilirubin
C4036889|T201|COMP|77447-1|LNC|Nordiazepam|Nordiazepam
C4036934|T201|COMP|77400-0|LNC|Human papilloma virus 18 DNA|Human papilloma virus 18 DNA
C4036935|T201|COMP|77399-4|LNC|Human papilloma virus 16 DNA|Human papilloma virus 16 DNA
C4036937|T201|COMP|77397-8|LNC|ABO & Rh group|ABO & Rh group
C4036938|T201|COMP|77396-0|LNC|Human papilloma virus 16 DNA|Human papilloma virus 16 DNA
C4036939|T201|COMP|77395-2|LNC|Human papilloma virus 18 DNA|Human papilloma virus 18 DNA
C4036942|T201|COMP|77392-9|LNC|Parainfluenza virus 3 Ag|Parainfluenza virus 3 Ag
C4036943|T201|COMP|77391-1|LNC|Parainfluenza virus 2 Ag|Parainfluenza virus 2 Ag
C4036944|T201|COMP|77390-3|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C4036945|T201|COMP|77389-5|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C4036946|T201|COMP|77388-7|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C4036947|T201|COMP|77387-9|LNC|Parainfluenza virus 3 Ag|Parainfluenza virus 3 Ag
C4036948|T201|COMP|77386-1|LNC|Parainfluenza virus 2 Ag|Parainfluenza virus 2 Ag
C4036949|T201|COMP|77385-3|LNC|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C4036950|T201|COMP|77384-6|LNC|Influenza virus B Ag|Influenza virus B Ag
C4036957|T201|COMP|77373-9|LNC|Lathosterol|Lathosterol
C4036958|T201|COMP|77372-1|LNC|3-Methoxytyramine.free|3-Methoxytyramine.free
C4036959|T201|COMP|77371-3|LNC|Brassicasterol|Brassicasterol
C4036960|T201|COMP|77370-5|LNC|Procollagen type I.N-terminal propeptide|Procollagen type I.N-terminal propeptide
C4036961|T201|COMP|77369-7|LNC|HIV 1 RNA|HIV 1 RNA
C4036962|T201|COMP|77368-9|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C4036963|T201|COMP|77367-1|LNC|Cholinesterase^dibucaine|Cholinesterase^dibucaine
C4036965|T201|COMP|77365-5|LNC|Nitrogen panel|Nitrogen panel
C4036966|T201|COMP|77364-8|LNC|Tryptophan, kynurenin & 3-hydroxykynurenin panel|Tryptophan, kynurenin & 3-hydroxykynurenin panel
C4036967|T201|COMP|77363-0|LNC|N-tau methylimidazoleacetate/Creatinine|N-tau methylimidazoleacetate/Creatinine
C4036968|T201|COMP|77362-2|LNC|N-tau methylimidazoleacetate/Creatinine|N-tau methylimidazoleacetate/Creatinine
C4036969|T201|COMP|77361-4|LNC|Triglyceride|Triglyceride
C4036970|T201|COMP|77360-6|LNC|Triglyceride|Triglyceride
C4036971|T201|COMP|77359-8|LNC|Protein|Protein
C4036972|T201|COMP|77358-0|LNC|Nitrogen|Nitrogen
C4036973|T201|COMP|77357-2|LNC|Nitrogen|Nitrogen
C4036974|T201|COMP|77356-4|LNC|Non-hematopoietic stem cells/100 leukocytes|Non-hematopoietic stem cells/100 leukocytes
C4036975|T201|COMP|77355-6|LNC|Non-hematopoietic stem cells/100 leukocytes|Non-hematopoietic stem cells/100 leukocytes
C4036979|T201|COMP|77350-7|LNC|Erythropoietin Ab|Erythropoietin Ab
C4036980|T201|COMP|77349-9|LNC|Everolimus^trough|Everolimus^trough
C4036981|T201|COMP|77348-1|LNC|Tacrolimus^trough|Tacrolimus^trough
C4036982|T201|COMP|77347-3|LNC|Beta-2 transferrin panel|Beta-2 transferrin panel
C4036983|T201|COMP|77346-5|LNC|Enterobius vermicularis^3rd specimen|Enterobius vermicularis^3rd specimen
C4036984|T201|COMP|77345-7|LNC|Enterobius vermicularis^2nd specimen|Enterobius vermicularis^2nd specimen
C4036985|T201|COMP|77344-0|LNC|Colony count|Colony count
C4036986|T201|COMP|77343-2|LNC|Gamma globulin|Gamma globulin
C4036987|T201|COMP|77342-4|LNC|Beta 1 globulin|Beta 1 globulin
C4036988|T201|COMP|77341-6|LNC|Anion gap 4|Anion gap 4
C4036989|T201|COMP|77340-8|LNC|Alpha 1 globulin|Alpha 1 globulin
C4036990|T201|COMP|77334-1|LNC|Norpropoxyphene|Norpropoxyphene
C4036991|T201|COMP|77333-3|LNC|Imipramine+Desipramine|Imipramine+Desipramine
C4036992|T201|COMP|77332-5|LNC|Morphine|Morphine
C4036993|T201|COMP|77331-7|LNC|Nortrimipramine|Nortrimipramine
C4036994|T201|COMP|77330-9|LNC|Protriptyline|Protriptyline
C4036995|T201|COMP|77329-1|LNC|Temazepam|Temazepam
C4036996|T201|COMP|77328-3|LNC|Methadone|Methadone
C4036997|T201|COMP|77327-5|LNC|Triazolam|Triazolam
C4036998|T201|COMP|77326-7|LNC|LORazepam|LORazepam
C4036999|T201|COMP|77325-9|LNC|N-desalkylflurazepam|N-desalkylflurazepam
C4037000|T201|COMP|77324-2|LNC|Flurazepam|Flurazepam
C4037001|T201|COMP|77323-4|LNC|diazePAM|diazePAM
C4037002|T201|COMP|77322-6|LNC|Amitriptyline+Nortriptyline|Amitriptyline+Nortriptyline
C4037003|T201|COMP|77321-8|LNC|Cyanide|Cyanide
C4037004|T201|COMP|77320-0|LNC|Benzoylecgonine|Benzoylecgonine
C4037005|T201|COMP|77319-2|LNC|Allergen.miscellaneous Ab.IgE.RAST class|Allergen.miscellaneous Ab.IgE.RAST class
C4037014|T201|COMP|77307-7|LNC|Lead|Lead
C4037062|T201|COMP|77955-3|LNC|Yellow fever virus Ab.IgM|Yellow fever virus Ab.IgM
C4037063|T201|COMP|77954-6|LNC|Yellow fever virus Ab.IgG|Yellow fever virus Ab.IgG
C4037064|T201|COMP|77953-8|LNC|West Nile virus Ab.IgG|West Nile virus Ab.IgG
C4037065|T201|COMP|77952-0|LNC|Trypanosoma cruzi Ab|Trypanosoma cruzi Ab
C4037066|T201|COMP|77951-2|LNC|Toscana virus Ab.IgG|Toscana virus Ab.IgG
C4037067|T201|COMP|77745-8|LNC|HTLV I p19-I Ab|HTLV I p19-I Ab
C4037068|T201|COMP|77744-1|LNC|HTLV I & II Ab band pattern|HTLV I & II Ab band pattern
C4037069|T201|COMP|77743-3|LNC|Toxocara sp Ab|Toxocara sp Ab
C4037070|T201|COMP|77742-5|LNC|HTLV I & II panel|HTLV I & II panel
C4037071|T201|COMP|77741-7|LNC|Streptavidin|Streptavidin
C4037072|T201|COMP|77676-5|LNC|Gastrin^30M post XXX challenge|Gastrin^30M post XXX challenge
C4037073|T201|COMP|77675-7|LNC|Gastrin^15M post XXX challenge|Gastrin^15M post XXX challenge
C4037074|T201|COMP|77674-0|LNC|Gastrin^10M post XXX challenge|Gastrin^10M post XXX challenge
C4037075|T201|COMP|77673-2|LNC|Gastrin^5M post XXX challenge|Gastrin^5M post XXX challenge
C4037076|T201|COMP|77672-4|LNC|Gastrin^3M post XXX challenge|Gastrin^3M post XXX challenge
C4037077|T201|COMP|77581-7|LNC|Alpha 2 globulin|Alpha 2 globulin
C4037080|T201|COMP|77250-9|LNC|Mumps virus IgG & IgM panel|Mumps virus IgG & IgM panel
C4037105|T201|COMP|77220-2|LNC|Niobium|Niobium
C4037107|T201|COMP|77216-0|LNC|Parotid secretory protein Ab.IgM|Parotid secretory protein Ab.IgM
C4037108|T201|COMP|77215-2|LNC|Parotid secretory protein Ab.IgG|Parotid secretory protein Ab.IgG
C4037109|T201|COMP|77214-5|LNC|Parotid secretory protein Ab.IgA|Parotid secretory protein Ab.IgA
C4037110|T201|COMP|77213-7|LNC|Carbonic anhydrase 6 Ab.IgM|Carbonic anhydrase 6 Ab.IgM
C4037111|T201|COMP|77212-9|LNC|Carbonic anhydrase 6 Ab.IgG|Carbonic anhydrase 6 Ab.IgG
C4037112|T201|COMP|77211-1|LNC|Carbonic anhydrase 6 Ab.IgA|Carbonic anhydrase 6 Ab.IgA
C4037113|T201|COMP|77210-3|LNC|Salivary gland protein 1 Ab.IgG|Salivary gland protein 1 Ab.IgG
C4037114|T201|COMP|77209-5|LNC|Salivary gland protein 1 Ab.IgM|Salivary gland protein 1 Ab.IgM
C4037115|T201|COMP|77208-7|LNC|Salivary gland protein 1 Ab.IgA|Salivary gland protein 1 Ab.IgA
C4037116|T201|COMP|77207-9|LNC|Naloxone|Naloxone
C4037117|T201|COMP|77206-1|LNC|Norbuprenorphine|Norbuprenorphine
C4037119|T201|COMP|77193-1|LNC|Bacteria identified|Bacteria identified
C4037120|T201|COMP|77192-3|LNC|Prealbumin|Prealbumin
C4037122|T201|COMP|77189-9|LNC|Zirconium/Creatinine|Zirconium/Creatinine
C4037123|T201|COMP|77188-1|LNC|Zirconium|Zirconium
C4037124|T201|COMP|77187-3|LNC|Zirconium|Zirconium
C4037125|T201|COMP|77186-5|LNC|Uranium|Uranium
C4037126|T201|COMP|77185-7|LNC|Uranium|Uranium
C4037127|T201|COMP|77175-8|LNC|Coxiella burnetii phase 1 & 2 Ab.IgG & IgM panel|Coxiella burnetii phase 1 & 2 Ab.IgG & IgM panel
C4037128|T201|COMP|77174-1|LNC|CALR gene exon 9 targeted mutation analysis|CALR gene exon 9 targeted mutation analysis
C4037129|T201|COMP|77173-3|LNC|Hepatocyte growth factor receptor Ag|Hepatocyte growth factor receptor Ag
C4037130|T201|COMP|77172-5|LNC|KIT gene exon 9 targeted mutation analysis|KIT gene exon 9 targeted mutation analysis
C4037131|T201|COMP|77171-7|LNC|KIT gene exon 11 targeted mutation analysis|KIT gene exon 11 targeted mutation analysis
C4037132|T201|COMP|77170-9|LNC|PDGFRA gene.p.Asp842Val|PDGFRA gene.p.Asp842Val
C4037133|T201|COMP|77169-1|LNC|cycloSPORINE^1H post dose|cycloSPORINE^1H post dose
C4037134|T201|COMP|77168-3|LNC|cycloSPORINE^4H post dose|cycloSPORINE^4H post dose
C4037135|T201|COMP|77167-5|LNC|cycloSPORINE^3H post dose|cycloSPORINE^3H post dose
C4037136|T201|COMP|77166-7|LNC|Chlamydia sp Ab.IgG & IgM panel|Chlamydia sp Ab.IgG & IgM panel
C4037138|T201|COMP|77164-2|LNC|Karyotype|Karyotype
C4037139|T201|COMP|77163-4|LNC|Alpha-1-Microglobulin|Alpha-1-Microglobulin
C4037140|T201|COMP|77162-6|LNC|Anidulafungin|Anidulafungin
C4037142|T201|COMP|77159-2|LNC|Erythrocytes.ghost cells|Erythrocytes.ghost cells
C4037143|T201|COMP|77158-4|LNC|Albumin|Albumin
C4037150|T201|COMP|77151-9|LNC|Energy content panel|Energy content panel
C4037151|T201|COMP|77150-1|LNC|Energy content|Energy content
C4037152|T201|COMP|77149-3|LNC|Specimen.dry weight/total|Specimen.dry weight/total
C4037153|T201|COMP|77148-5|LNC|Albumin|Albumin
C4037154|T201|COMP|77147-7|LNC|Glomerular filtration rate/1.73 sq M.predicted|Glomerular filtration rate/1.73 sq M.predicted
C4037155|T201|COMP|77146-9|LNC|Amylase|Amylase
C4037156|T201|COMP|77145-1|LNC|Glucose^post CFst|Glucose^post CFst
C4037157|T201|COMP|77144-4|LNC|Alanine aminotransferase|Alanine aminotransferase
C4037158|T201|COMP|77135-2|LNC|Glucose|Glucose
C4037160|T201|COMP|77133-7|LNC|LCA5 gene full mutation analysis|LCA5 gene full mutation analysis
C4037162|T201|COMP|77131-1|LNC|CDHR1 gene full mutation analysis|CDHR1 gene full mutation analysis
C4037164|T201|COMP|77129-5|LNC|CERKL gene full mutation analysis|CERKL gene full mutation analysis
C4037166|T201|COMP|77127-9|LNC|USH1C gene full mutation analysis|USH1C gene full mutation analysis
C4037168|T201|COMP|77125-3|LNC|PCDH15 gene full mutation analysis|PCDH15 gene full mutation analysis
C4037170|T201|COMP|77123-8|LNC|GPR98 gene full mutation analysis|GPR98 gene full mutation analysis
C4037172|T201|COMP|77121-2|LNC|DFNB31 gene full mutation analysis|DFNB31 gene full mutation analysis
C4037174|T201|COMP|77119-6|LNC|RPGR gene full mutation analysis|RPGR gene full mutation analysis
C4037176|T201|COMP|77117-0|LNC|RPGRIP1 gene full mutation analysis|RPGRIP1 gene full mutation analysis
C4037178|T201|COMP|77115-4|LNC|FKBP10 gene full mutation analysis|FKBP10 gene full mutation analysis
C4037179|T201|COMP|77114-7|LNC|FBN1 gene full mutation analysis|FBN1 gene full mutation analysis
C4037181|T201|COMP|77112-1|LNC|PLOD3 gene full mutation analysis|PLOD3 gene full mutation analysis
C4037183|T201|COMP|77110-5|LNC|KARS gene full mutation analysis|KARS gene full mutation analysis
C4037185|T201|COMP|77108-9|LNC|AARS2 gene full mutation analysis|AARS2 gene full mutation analysis
C4037187|T201|COMP|77106-3|LNC|SARS2 gene full mutation analysis|SARS2 gene full mutation analysis
C4037189|T201|COMP|77104-8|LNC|HARS2 gene full mutation analysis|HARS2 gene full mutation analysis
C4037191|T201|COMP|77102-2|LNC|NARS2 gene full mutation analysis|NARS2 gene full mutation analysis
C4037193|T201|COMP|77100-6|LNC|MRPS18A gene full mutation analysis|MRPS18A gene full mutation analysis
C4037195|T201|COMP|77098-2|LNC|MRPL44 gene full mutation analysis|MRPL44 gene full mutation analysis
C4037197|T201|COMP|77096-6|LNC|MRPS22 gene full mutation analysis|MRPS22 gene full mutation analysis
C4037199|T201|COMP|77094-1|LNC|MRPS2 gene full mutation analysis|MRPS2 gene full mutation analysis
C4037201|T201|COMP|77092-5|LNC|MRRF gene full mutation analysis|MRRF gene full mutation analysis
C4037203|T201|COMP|77090-9|LNC|TFB1M gene full mutation analysis|TFB1M gene full mutation analysis
C4037205|T201|COMP|77088-3|LNC|GFM1 gene full mutation analysis|GFM1 gene full mutation analysis
C4037208|T201|COMP|77080-0|LNC|SERPINF1 gene full mutation analysis|SERPINF1 gene full mutation analysis
C4037210|T201|COMP|77078-4|LNC|MTFMT gene full mutation analysis|MTFMT gene full mutation analysis
C4037212|T201|COMP|77076-8|LNC|MRPL40 gene full mutation analysis|MRPL40 gene full mutation analysis
C4037214|T201|COMP|77074-3|LNC|C12orf65 gene full mutation analysis|C12orf65 gene full mutation analysis
C4037216|T201|COMP|77072-7|LNC|ATP5A1 gene full mutation analysis|ATP5A1 gene full mutation analysis
C4037218|T201|COMP|77070-1|LNC|PLOD2 gene full mutation analysis|PLOD2 gene full mutation analysis
C4037220|T201|COMP|77068-5|LNC|AGA gene full mutation analysis|AGA gene full mutation analysis
C4037221|T201|COMP|77067-7|LNC|SEPT9 gene targeted mutation analysis|SEPT9 gene targeted mutation analysis
C4037223|T201|COMP|77065-1|LNC|AHCY gene full mutation analysis|AHCY gene full mutation analysis
C4037225|T201|COMP|77063-6|LNC|TAT gene full mutation analysis|TAT gene full mutation analysis
C4037227|T201|COMP|77061-0|LNC|HPD gene full mutation analysis|HPD gene full mutation analysis
C4037229|T201|COMP|77059-4|LNC|GNMT gene full mutation analysis|GNMT gene full mutation analysis
C4037231|T201|COMP|77057-8|LNC|CYP17A1 gene full mutation analysis|CYP17A1 gene full mutation analysis
C4037233|T201|COMP|77055-2|LNC|CYP11B1 gene full mutation analysis|CYP11B1 gene full mutation analysis
C4037235|T201|COMP|77053-7|LNC|MTR gene full mutation analysis|MTR gene full mutation analysis
C4037237|T201|COMP|77051-1|LNC|IFITM5 gene full mutation analysis|IFITM5 gene full mutation analysis
C4037239|T201|COMP|77049-5|LNC|SUGCT gene full mutation analysis|SUGCT gene full mutation analysis
C4037241|T201|COMP|77047-9|LNC|ACSF3 gene full mutation analysis|ACSF3 gene full mutation analysis
C4037243|T201|COMP|77045-3|LNC|ACADSB gene full mutation analysis|ACADSB gene full mutation analysis
C4037245|T201|COMP|77043-8|LNC|ACAD8 gene full mutation analysis|ACAD8 gene full mutation analysis
C4037246|T201|COMP|77042-0|LNC|t(6;9)(p22;q34)(DEK,NUP214) fusion transcript|t(6;9)(p22;q34)(DEK,NUP214) fusion transcript
C4037249|T201|COMP|77039-6|LNC|t(12;21)(p13;q22.3)(ETV6,RUNX1) fusion transcript|t(12;21)(p13;q22.3)(ETV6,RUNX1) fusion transcript
C4037250|T201|COMP|77038-8|LNC|t(14;18)(q32;q21.3)(IGH,BCL2) fusion transcript|t(14;18)(q32;q21.3)(IGH,BCL2) fusion transcript
C4037251|T201|COMP|77037-0|LNC|t(11;14)(q13;q32)(CCND1,IGH) fusion transcript|t(11;14)(q13;q32)(CCND1,IGH) fusion transcript
C4037252|T201|COMP|77036-2|LNC|t(11;18)(q21;q21)(BIRC3,MALT1) fusion transcript|t(11;18)(q21;q21)(BIRC3,MALT1) fusion transcript
C4037253|T201|COMP|77035-4|LNC|t(14;18)(q32;q21)(IGH,MALT1) fusion transcript|t(14;18)(q32;q21)(IGH,MALT1) fusion transcript
C4037255|T201|COMP|77033-9|LNC|t(14;16)(q32;q23)(IGH,MAF) fusion transcript|t(14;16)(q32;q23)(IGH,MAF) fusion transcript
C4037256|T201|COMP|77032-1|LNC|t(8;14)(q24;q32)(MYC,IGH) fusion transcript|t(8;14)(q24;q32)(MYC,IGH) fusion transcript
C4037257|T201|COMP|77031-3|LNC|t(15;17)(q24.1;q21.1)(PML,RARA) fusion transcript|t(15;17)(q24.1;q21.1)(PML,RARA) fusion transcript
C4037258|T201|COMP|77030-5|LNC|t(1;19)(q23.3;p13.3)(PBX1,TCF3) fusion transcript|t(1;19)(q23.3;p13.3)(PBX1,TCF3) fusion transcript
C4037259|T201|COMP|77029-7|LNC|Respiratory pathogens DNA & RNA 14 panel|Respiratory pathogens DNA & RNA 14 panel
C4037260|T201|COMP|77028-9|LNC|Influenza virus A H1 2009 pandemic RNA|Influenza virus A H1 2009 pandemic RNA
C4037261|T201|COMP|77027-1|LNC|Influenza virus A H3 RNA|Influenza virus A H3 RNA
C4037262|T201|COMP|77026-3|LNC|Influenza virus A H1 RNA|Influenza virus A H1 RNA
C4037263|T201|COMP|77025-5|LNC|Rhinovirus RNA|Rhinovirus RNA
C4037264|T201|COMP|77024-8|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C4037267|T201|COMP|77017-2|LNC|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C4037268|T201|COMP|77016-4|LNC|Fetal RhD antigen|Fetal RhD antigen
C4037269|T201|COMP|77015-6|LNC|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C4037270|T201|COMP|77014-9|LNC|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C4037271|T201|COMP|77010-7|LNC|Urea^post dialysis/pre dialysis|Urea^post dialysis/pre dialysis
C4037272|T201|COMP|77009-9|LNC|Porphyrin fractions panel|Porphyrin fractions panel
C4037273|T201|COMP|77008-1|LNC|Human coronavirus 229E+OC43 RNA|Human coronavirus 229E+OC43 RNA
C4037450|T201|COMP|77961-1|LNC|cloZAPine|cloZAPine
C4037451|T201|COMP|77960-3|LNC|Penicillin.parenteral|Penicillin.parenteral
C4037452|T201|COMP|77958-7|LNC|Dengue virus 1 & 2 & 3 & 4 RNA|Dengue virus 1 & 2 & 3 & 4 RNA
C4037453|T201|COMP|77957-9|LNC|Yersinia enterocolitica O:9 Ab.IgG|Yersinia enterocolitica O:9 Ab.IgG
C4037454|T201|COMP|77956-1|LNC|Yersinia enterocolitica O:3 Ab.IgG|Yersinia enterocolitica O:3 Ab.IgG
C4037455|T201|COMP|77950-4|LNC|Toscana virus Ab.IgM|Toscana virus Ab.IgM
C4037456|T201|COMP|77949-6|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C4037462|T201|COMP|77655-9|LNC|Cells.diploid/100 cells|Cells.diploid/100 cells
C4037463|T201|COMP|77654-2|LNC|Cells.diploid.G2 phase/100 cells|Cells.diploid.G2 phase/100 cells
C4037465|T201|COMP|77652-6|LNC|C peptide^5H post XXX challenge|C peptide^5H post XXX challenge
C4037466|T201|COMP|77651-8|LNC|C peptide^75M post XXX challenge|C peptide^75M post XXX challenge
C4037467|T201|COMP|77650-0|LNC|17-Hydroxyprogesterone^15M post XXX challenge|17-Hydroxyprogesterone^15M post XXX challenge
C4037468|T201|COMP|77608-8|LNC|Androstenedione^30M post XXX challenge|Androstenedione^30M post XXX challenge
C4037469|T201|COMP|77607-0|LNC|Cortisol^1M post XXX challenge|Cortisol^1M post XXX challenge
C4037471|T201|COMP|77605-4|LNC|Influenza virus A H5 icA RNA|Influenza virus A H5 icA RNA
C4037475|T201|COMP|77254-1|LNC|Albumin/Creatinine|Albumin/Creatinine
C4037476|T201|COMP|77253-3|LNC|Albumin/Creatinine|Albumin/Creatinine
C4037477|T201|COMP|77184-0|LNC|Niobium/Creatinine|Niobium/Creatinine
C4037478|T201|COMP|77183-2|LNC|Niobium|Niobium
C4037479|T201|COMP|77182-4|LNC|Niobium|Niobium
C4037480|T201|COMP|77181-6|LNC|Niobium|Niobium
C4037481|T201|COMP|77180-8|LNC|Niobium|Niobium
C4037482|T201|COMP|77179-0|LNC|Niobium|Niobium
C4037483|T201|COMP|77178-2|LNC|Boron|Boron
C4037484|T201|COMP|77177-4|LNC|IgG|IgG
C4037485|T201|COMP|77176-6|LNC|Hepatitis B virus little e Ag & Ab panel|Hepatitis B virus little e Ag & Ab panel
C4037499|T201|COMP|76773-1|LNC|Heptacarboxylporphyrin|Heptacarboxylporphyrin
C4037500|T201|COMP|76772-3|LNC|Plasmodium falciparum Ag|Plasmodium falciparum Ag
C4037501|T201|COMP|76771-5|LNC|Respiratory pathogens RNA 8 panel|Respiratory pathogens RNA 8 panel
C4037502|T201|COMP|76770-7|LNC|Trace elements panel|Trace elements panel
C4037503|T201|COMP|76769-9|LNC|Hemoglobin|Hemoglobin
C4037504|T201|COMP|76768-1|LNC|Hemoglobin|Hemoglobin
C4037505|T201|COMP|76767-3|LNC|Schistosoma sp identified|Schistosoma sp identified
C4037506|T201|COMP|76766-5|LNC|Treponema pallidum PolA gene|Treponema pallidum PolA gene
C4037507|T201|COMP|76765-7|LNC|Phosphatidylcholine.saturated|Phosphatidylcholine.saturated
C4037555|T201|COMP|76705-3|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C4037556|T201|COMP|76699-8|LNC|Filaria identified|Filaria identified
C4037559|T201|COMP|76693-1|LNC|Bacteria identified|Bacteria identified
C4037560|T201|COMP|76692-3|LNC|Fungus identified|Fungus identified
C4037561|T201|COMP|76688-1|LNC|Alpha-1-acid glycoprotein/Creatinine|Alpha-1-acid glycoprotein/Creatinine
C4037562|T201|COMP|76683-2|LNC|Mean platelet component|Mean platelet component
C4037563|T201|COMP|76682-4|LNC|Color^4th tube|Color^4th tube
C4037564|T201|COMP|76680-8|LNC|Color^2nd tube|Color^2nd tube
C4037565|T201|COMP|76679-0|LNC|Color^1st tube|Color^1st tube
C4037566|T201|COMP|76672-5|LNC|Glucose^4th tube|Glucose^4th tube
C4037567|T201|COMP|76671-7|LNC|Glucose^3rd tube|Glucose^3rd tube
C4037568|T201|COMP|76670-9|LNC|Glucose^2nd tube|Glucose^2nd tube
C4037569|T201|COMP|76669-1|LNC|Glucose^1st tube|Glucose^1st tube
C4037570|T201|COMP|76668-3|LNC|Protein^4th tube|Protein^4th tube
C4037573|T201|COMP|76660-0|LNC|Phosphatidylethanol|Phosphatidylethanol
C4037574|T201|COMP|76659-2|LNC|Antipsychotics drug panel|Antipsychotics drug panel
C4037575|T201|COMP|76658-4|LNC|Zirconium|Zirconium
C4037576|T201|COMP|76657-6|LNC|Iodine|Iodine
C4037577|T201|COMP|76656-8|LNC|Phosphate|Phosphate
C4037578|T201|COMP|76655-0|LNC|Tungsten|Tungsten
C4037579|T201|COMP|76654-3|LNC|Beryllium|Beryllium
C4037580|T201|COMP|76653-5|LNC|Barium|Barium
C4037581|T201|COMP|76652-7|LNC|Thorium|Thorium
C4037582|T201|COMP|76651-9|LNC|Zinc transporter 8 Ab|Zinc transporter 8 Ab
C4037583|T201|COMP|76650-1|LNC|Gadolinium|Gadolinium
C4037584|T201|COMP|76649-3|LNC|Germanium|Germanium
C4037585|T201|COMP|76648-5|LNC|Palladium|Palladium
C4037586|T201|COMP|76647-7|LNC|Strontium|Strontium
C4037595|T201|COMP|76633-7|LNC|Glomerular filtration rate/1.73 sq M.predicted|Glomerular filtration rate/1.73 sq M.predicted
C4037596|T201|COMP|76632-9|LNC|Enterovirus sp|Enterovirus sp
C4037597|T201|COMP|76631-1|LNC|Albumin|Albumin
C4037598|T201|COMP|76630-3|LNC|Amylase|Amylase
C4037599|T201|COMP|76629-5|LNC|Glucose^post CFst|Glucose^post CFst
C4037600|T201|COMP|76628-7|LNC|Norovirus genogroup I & II RNA|Norovirus genogroup I & II RNA
C4037601|T201|COMP|76627-9|LNC|Rifapentine|Rifapentine
C4037602|T201|COMP|76626-1|LNC|Measles virus|Measles virus
C4037603|T201|COMP|76625-3|LNC|Alanine aminotransferase|Alanine aminotransferase
C4037604|T201|COMP|76624-6|LNC|Mitochondrial respiratory chain enzyme analysis|Mitochondrial respiratory chain enzyme analysis
C4037606|T201|COMP|76622-0|LNC|Lysosomal acid lipase|Lysosomal acid lipase
C4037607|T201|COMP|76621-2|LNC|Lysosomal acid lipase panel|Lysosomal acid lipase panel
C4037608|T201|COMP|76620-4|LNC|Mitochondrial respiratory chain enzymes|Mitochondrial respiratory chain enzymes
C4037609|T201|COMP|76619-6|LNC|Mitochondrial respiratory chain enzymes|Mitochondrial respiratory chain enzymes
C4037610|T201|COMP|76618-8|LNC|Mitochondrial respiratory chain enzymes|Mitochondrial respiratory chain enzymes
C4037611|T201|COMP|76617-0|LNC|Mitochondrial respiratory chain enzymes|Mitochondrial respiratory chain enzymes
C4037612|T201|COMP|76616-2|LNC|Mitochondrial respiratory chain enzymes|Mitochondrial respiratory chain enzymes
C4037613|T201|COMP|76615-4|LNC|Lysosomal acid lipase|Lysosomal acid lipase
C4037614|T201|COMP|76614-7|LNC|Lysosomal acid lipase|Lysosomal acid lipase
C4037616|T201|COMP|76612-1|LNC|Enterococcus faecalis cpn60 gene|Enterococcus faecalis cpn60 gene
C4037617|T201|COMP|76611-3|LNC|Klebsiella pneumoniae phoE gene|Klebsiella pneumoniae phoE gene
C4037618|T201|COMP|76610-5|LNC|Streptococcus agalactiae cfb gene|Streptococcus agalactiae cfb gene
C4037619|T201|COMP|76609-7|LNC|Streptococcus pyogenes csrS gene|Streptococcus pyogenes csrS gene
C4037620|T201|COMP|76608-9|LNC|Candida albicans its gene|Candida albicans its gene
C4037621|T201|COMP|77205-3|LNC|Buprenorphine|Buprenorphine
C4037622|T201|COMP|77204-6|LNC|Buprenorphine|Buprenorphine
C4037624|T201|COMP|77202-0|LNC|Laboratory comment|Laboratory comment
C4037625|T201|COMP|77201-2|LNC|Buprenorphine+Norbuprenorphine|Buprenorphine+Norbuprenorphine
C4037626|T201|COMP|77200-4|LNC|SI gene targeted mutation analysis|SI gene targeted mutation analysis
C4037628|T201|COMP|77143-6|LNC|Carbon dioxide|Carbon dioxide
C4037629|T201|COMP|77142-8|LNC|Potassium|Potassium
C4037630|T201|COMP|77141-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C4037631|T201|COMP|77140-2|LNC|Creatinine|Creatinine
C4037632|T201|COMP|77086-7|LNC|TYROBP gene full mutation analysis|TYROBP gene full mutation analysis
C4037634|T201|COMP|77084-2|LNC|ALPL gene full mutation analysis|ALPL gene full mutation analysis
C4037636|T201|COMP|77082-6|LNC|FARS2 gene full mutation analysis|FARS2 gene full mutation analysis
C4037642|T201|COMP|77661-7|LNC|Cells.aneuploid.S phase population 2/100 cells|Cells.aneuploid.S phase population 2/100 cells
C4037643|T201|COMP|77660-9|LNC|Cells.aneuploid.G2 phase population 2/100 cells|Cells.aneuploid.G2 phase population 2/100 cells
C4037644|T201|COMP|77659-1|LNC|Cells.aneuploid.S phase population/100 cells|Cells.aneuploid.S phase population/100 cells
C4037645|T201|COMP|77658-3|LNC|Cells.aneuploid.G2 phase population/100 cells|Cells.aneuploid.G2 phase population/100 cells
C4037646|T201|COMP|77657-5|LNC|Cells.diploid.G1 phase/100 cells|Cells.diploid.G1 phase/100 cells
C4037659|T201|COMP|77023-0|LNC|Respiratory syncytial virus B RNA|Respiratory syncytial virus B RNA
C4037660|T201|COMP|77022-2|LNC|Respiratory syncytial virus A RNA|Respiratory syncytial virus A RNA
C4037661|T201|COMP|77021-4|LNC|Fetal Y chromosome|Fetal Y chromosome
C4037662|T201|COMP|77020-6|LNC|Fetal Y chromosome|Fetal Y chromosome
C4037667|T201|COMP|76687-3|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C4037669|T201|COMP|76685-7|LNC|Platelet dry mass distribution width|Platelet dry mass distribution width
C4037670|T201|COMP|76684-0|LNC|Mean platelet dry mass|Mean platelet dry mass
C4037676|T201|COMP|76667-5|LNC|Protein^3rd tube|Protein^3rd tube
C4037677|T201|COMP|76666-7|LNC|Protein^2nd tube|Protein^2nd tube
C4037678|T201|COMP|76665-9|LNC|Protein^1st tube|Protein^1st tube
C4037679|T201|COMP|76664-2|LNC|Fetal chromosome X & Y aneuploidy|Fetal chromosome X & Y aneuploidy
C4037681|T201|COMP|76607-1|LNC|Enterococcus faecium sodA gene|Enterococcus faecium sodA gene
C4037682|T201|COMP|76606-3|LNC|Pseudomonas aeruginosa regA gene|Pseudomonas aeruginosa regA gene
C4037683|T201|COMP|76605-5|LNC|Staphylococcus aureus sau3AI gene|Staphylococcus aureus sau3AI gene
C4037684|T201|COMP|76604-8|LNC|Serratia marcescens gyrB gene|Serratia marcescens gyrB gene
C4037685|T201|COMP|76603-0|LNC|Bacterial 16S rRNA|Bacterial 16S rRNA
C4037686|T201|COMP|76602-2|LNC|Haemophilus influenzae lex2 gene|Haemophilus influenzae lex2 gene
C4037687|T201|COMP|76601-4|LNC|Moraxella catarrhalis g1b gene|Moraxella catarrhalis g1b gene
C4037688|T201|COMP|76600-6|LNC|Streptococcus pneumoniae nanA gene|Streptococcus pneumoniae nanA gene
C4037689|T201|COMP|76599-0|LNC|Enterococcus faecalis cpn60 gene|Enterococcus faecalis cpn60 gene
C4037690|T201|COMP|76598-2|LNC|Klebsiella pneumoniae phoE gene|Klebsiella pneumoniae phoE gene
C4037691|T201|COMP|76597-4|LNC|Streptococcus agalactiae cfb gene|Streptococcus agalactiae cfb gene
C4037692|T201|COMP|76596-6|LNC|Streptococcus pyogenes csrS gene|Streptococcus pyogenes csrS gene
C4037693|T201|COMP|76595-8|LNC|Candida albicans its gene|Candida albicans its gene
C4037694|T201|COMP|76594-1|LNC|Enterococcus faecium sodA gene|Enterococcus faecium sodA gene
C4037695|T201|COMP|76593-3|LNC|Pseudomonas aeruginosa regA gene|Pseudomonas aeruginosa regA gene
C4037696|T201|COMP|76592-5|LNC|Staphylococcus aureus sau3AI gene|Staphylococcus aureus sau3AI gene
C4037697|T201|COMP|76591-7|LNC|Serratia marcescens gyrB gene|Serratia marcescens gyrB gene
C4037698|T201|COMP|76590-9|LNC|Bacterial 16S rRNA|Bacterial 16S rRNA
C4037699|T201|COMP|76589-1|LNC|Haemophilus influenzae lex2 gene|Haemophilus influenzae lex2 gene
C4037700|T201|COMP|76588-3|LNC|Moraxella catarrhalis g1b gene|Moraxella catarrhalis g1b gene
C4037701|T201|COMP|76587-5|LNC|Streptococcus pneumoniae nanA gene|Streptococcus pneumoniae nanA gene
C4037702|T201|COMP|76586-7|LNC|ENT microorganism gene identification panel|ENT microorganism gene identification panel
C4037703|T201|COMP|76585-9|LNC|Wound microorganism gene identification panel|Wound microorganism gene identification panel
C4037704|T201|COMP|76579-2|LNC|Enterococcus faecium sodA gene|Enterococcus faecium sodA gene
C4037705|T201|COMP|76578-4|LNC|Pseudomonas aeruginosa regA gene|Pseudomonas aeruginosa regA gene
C4037706|T201|COMP|76577-6|LNC|Staphylococcus aureus sau3AI gene|Staphylococcus aureus sau3AI gene
C4037707|T201|COMP|76576-8|LNC|Serratia marcescens gyrB gene|Serratia marcescens gyrB gene
C4037708|T201|COMP|76575-0|LNC|Bacterial 16S rRNA|Bacterial 16S rRNA
C4037709|T201|COMP|76574-3|LNC|Haemophilus influenzae lex2 gene|Haemophilus influenzae lex2 gene
C4037710|T201|COMP|76573-5|LNC|Moraxella catarrhalis g1b gene|Moraxella catarrhalis g1b gene
C4037711|T201|COMP|76572-7|LNC|Streptococcus pneumoniae nanA gene|Streptococcus pneumoniae nanA gene
C4037737|T201|COMP|76540-4|LNC|Pathology diagnosis ICD code|Pathology diagnosis ICD code
C4037738|T201|COMP|76524-8|LNC|Acetone|Acetone
C4037746|T201|COMP|76497-7|LNC|Polymorphonuclear cells|Polymorphonuclear cells
C4037747|T201|COMP|76496-9|LNC|Complement C4|Complement C4
C4037748|T201|COMP|76495-1|LNC|Titanium|Titanium
C4037749|T201|COMP|76494-4|LNC|Tacrolimus|Tacrolimus
C4037750|T201|COMP|76493-6|LNC|Nitrazepam|Nitrazepam
C4037751|T201|COMP|76492-8|LNC|Amphetamine+Methamphetamine|Amphetamine+Methamphetamine
C4037752|T201|COMP|76491-0|LNC|IgM|IgM
C4037753|T201|COMP|76490-2|LNC|IgG|IgG
C4037754|T201|COMP|76489-4|LNC|IgG|IgG
C4037755|T201|COMP|76488-6|LNC|IgE|IgE
C4037756|T201|COMP|76487-8|LNC|IgA|IgA
C4037757|T201|COMP|76486-0|LNC|C reactive protein|C reactive protein
C4037758|T201|COMP|76485-2|LNC|C reactive protein|C reactive protein
C4037759|T201|COMP|76484-5|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C4037760|T201|COMP|76482-9|LNC|Apolipoprotein B|Apolipoprotein B
C4037761|T201|COMP|76481-1|LNC|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C4037762|T201|COMP|76480-3|LNC|Albumin|Albumin
C4037763|T201|COMP|76479-5|LNC|Acetylcholinesterase|Acetylcholinesterase
C4037764|T201|COMP|76478-7|LNC|Acetylcholinesterase panel|Acetylcholinesterase panel
C4037765|T201|COMP|76475-3|LNC|Cortisone.free|Cortisone.free
C4037766|T201|COMP|76474-6|LNC|Ghrelin|Ghrelin
C4037778|T201|COMP|76413-4|LNC|Sheep prion protein codon 112|Sheep prion protein codon 112
C4037779|T201|COMP|76412-6|LNC|Sheep prion protein codon 141|Sheep prion protein codon 141
C4037780|T201|COMP|76411-8|LNC|Neutrophils|Neutrophils
C4037781|T201|COMP|76410-0|LNC|Neutrophils.band form|Neutrophils.band form
C4037782|T201|COMP|76409-2|LNC|Lymphocytes|Lymphocytes
C4037783|T201|COMP|76408-4|LNC|Monocytes+Macrophages|Monocytes+Macrophages
C4037784|T201|COMP|76407-6|LNC|Eosinophils|Eosinophils
C4037785|T201|COMP|76406-8|LNC|Basophils|Basophils
C4037786|T201|COMP|76405-0|LNC|Metamyelocytes|Metamyelocytes
C4037787|T201|COMP|76404-3|LNC|Promyelocytes|Promyelocytes
C4037788|T201|COMP|76403-5|LNC|Blasts|Blasts
C4037789|T201|COMP|76402-7|LNC|Myelocytes|Myelocytes
C4037790|T201|COMP|76401-9|LNC|Albumin/Creatinine|Albumin/Creatinine
C4037792|T201|COMP|76399-5|LNC|Troponin I.cardiac|Troponin I.cardiac
C4037829|T201|COMP|76352-4|LNC|Testosterone/Cortisol|Testosterone/Cortisol
C4037830|T201|COMP|76351-6|LNC|Methotrexate polyglutamates|Methotrexate polyglutamates
C4037831|T201|COMP|76350-8|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C4037832|T201|COMP|76349-0|LNC|clonazePAM|clonazePAM
C4037833|T201|COMP|76348-2|LNC|Pregnancy associated plasma protein A^^adjusted|Pregnancy associated plasma protein A^^adjusted
C4037834|T201|COMP|76347-4|LNC|Dehydroepiandrosterone sulfate/cortisol|Dehydroepiandrosterone sulfate/cortisol
C4037835|T201|COMP|76346-6|LNC|Microorganism identified|Microorganism identified
C4037837|T201|COMP|76341-7|LNC|Protoporphyrin|Protoporphyrin
C4037838|T201|COMP|76340-9|LNC|Porcine deltacoronavirus RNA|Porcine deltacoronavirus RNA
C4037839|T201|COMP|76339-1|LNC|Porcine deltacoronavirus RNA|Porcine deltacoronavirus RNA
C4037840|T201|COMP|76338-3|LNC|Porcine epidemic diarrhea virus RNA|Porcine epidemic diarrhea virus RNA
C4037841|T201|COMP|76150-2|LNC|Cefquinome|Cefquinome
C4037842|T201|COMP|76148-6|LNC|Pradofloxacin|Pradofloxacin
C4037843|T201|COMP|76147-8|LNC|Cefovecin|Cefovecin
C4037844|T201|COMP|76146-0|LNC|Tosufloxacin|Tosufloxacin
C4037845|T201|COMP|76145-2|LNC|Prulifloxacin|Prulifloxacin
C4037846|T201|COMP|76144-5|LNC|Cefteram|Cefteram
C4037847|T201|COMP|76143-7|LNC|Cefcapene|Cefcapene
C4037848|T201|COMP|76142-9|LNC|Lymphocytes.immature|Lymphocytes.immature
C4037850|T201|COMP|76140-3|LNC|Reticulocytes.hypochromic/100 erythrocytes|Reticulocytes.hypochromic/100 erythrocytes
C4037851|T201|COMP|76139-5|LNC|Reticulocyte hemoglobin distribution width|Reticulocyte hemoglobin distribution width
C4037852|T201|COMP|76138-7|LNC|Reticulocyte distribution width|Reticulocyte distribution width
C4037853|T201|COMP|76137-9|LNC|Platelet component distribution width|Platelet component distribution width
C4037854|T201|COMP|76132-0|LNC|Sucrose/Creatinine|Sucrose/Creatinine
C4037855|T201|COMP|76091-8|LNC|Respiratory pathogens DNA & RNA 4 panel|Respiratory pathogens DNA & RNA 4 panel
C4037856|T201|COMP|77383-8|LNC|Influenza virus A Ag|Influenza virus A Ag
C4037857|T201|COMP|77382-0|LNC|Adenovirus Ag|Adenovirus Ag
C4037859|T201|COMP|77339-0|LNC|Indocyanine green^15M post dose indocyanine green|Indocyanine green^15M post dose indocyanine green
C4037860|T201|COMP|77338-2|LNC|Indocyanine green^1M post dose indocyanine green|Indocyanine green^1M post dose indocyanine green
C4037861|T201|COMP|77337-4|LNC|Trimipramine+Nortrimipramine|Trimipramine+Nortrimipramine
C4037862|T201|COMP|77336-6|LNC|Oxazepam|Oxazepam
C4037863|T201|COMP|77335-8|LNC|Propoxyphene+Norpropoxyphene|Propoxyphene+Norpropoxyphene
C4037864|T201|COMP|77139-4|LNC|Sodium|Sodium
C4037865|T201|COMP|77138-6|LNC|Chloride|Chloride
C4037866|T201|COMP|77137-8|LNC|Bilirubin|Bilirubin
C4037867|T201|COMP|77136-0|LNC|Urea|Urea
C4037868|T201|COMP|76678-2|LNC|Appearance^4th tube|Appearance^4th tube
C4037869|T201|COMP|76677-4|LNC|Appearance^3rd tube|Appearance^3rd tube
C4037870|T201|COMP|76676-6|LNC|Appearance^2nd tube|Appearance^2nd tube
C4037871|T201|COMP|76675-8|LNC|Appearance^1st tube|Appearance^1st tube
C4037872|T201|COMP|76674-1|LNC|Leukocytes^1st tube|Leukocytes^1st tube
C4037873|T201|COMP|76673-3|LNC|Erythrocytes^1st tube|Erythrocytes^1st tube
C4037874|T201|COMP|76584-2|LNC|Enterococcus faecalis cpn60 gene|Enterococcus faecalis cpn60 gene
C4037875|T201|COMP|76583-4|LNC|Klebsiella pneumoniae phoE gene|Klebsiella pneumoniae phoE gene
C4037876|T201|COMP|76582-6|LNC|Streptococcus agalactiae cfb gene|Streptococcus agalactiae cfb gene
C4037877|T201|COMP|76581-8|LNC|Streptococcus pyogenes csrS gene|Streptococcus pyogenes csrS gene
C4037878|T201|COMP|76580-0|LNC|Candida albicans its gene|Candida albicans its gene
C4037880|T201|COMP|76414-2|LNC|Sheep prion protein codon 136|Sheep prion protein codon 136
C4037911|T201|COMP|76416-7|LNC|Sheep prion protein codon 171|Sheep prion protein codon 171
C4037912|T201|COMP|76415-9|LNC|Sheep prion protein codon 154|Sheep prion protein codon 154
C4037913|T201|COMP|74910-1|LNC|Porphyrin fractions & creatinine panel|Porphyrin fractions & creatinine panel
C4049659|T201|COMP|80402-1|LNC|Egg source|Egg source
C4049754|T201|COMP|80352-8|LNC|Environment temperature during transport|Environment temperature during transport
C4049778|T201|COMP|79265-5|LNC|Urea nitrogen^overnight dwell|Urea nitrogen^overnight dwell
C4050442|T201|COMP|79264-8|LNC|Glucose^overnight dwell|Glucose^overnight dwell
C4050490|T201|COMP|79568-2|LNC|ABCD1 gene targeted mutation analysis|ABCD1 gene targeted mutation analysis
C4050491|T201|COMP|79401-6|LNC|HBB gene full mutation analysis|HBB gene full mutation analysis
C4050496|T201|COMP|79544-3|LNC|HEDIS 2016 Value Sets|HEDIS 2016 Value Sets
C4050497|T201|COMP|79543-5|LNC|HEDIS 2016-2019 Value Set - ABO and Rh|HEDIS 2016-2019 Value Set - ABO and Rh
C4050528|T201|COMP|79263-0|LNC|Creatinine^overnight dwell|Creatinine^overnight dwell
C4050529|T201|COMP|79542-7|LNC|HEDIS 2016 Value Set - HPV Vaccine Administered|HEDIS 2016 Value Set - HPV Vaccine Administered
C4050530|T201|COMP|79541-9|LNC|HEDIS 2016-2020 Value Set - Lead Tests|HEDIS 2016-2020 Value Set - Lead Tests
C4050531|T201|COMP|79540-1|LNC|HEDIS 2016-2018 Value Set - PHQ-9 Total Score|HEDIS 2016-2018 Value Set - PHQ-9 Total Score
C4050532|T201|COMP|79539-3|LNC|HEDIS 2016-2018 Value Set - Urine Protein Tests|HEDIS 2016-2018 Value Set - Urine Protein Tests
C4050534|T201|COMP|79155-8|LNC|HIV 1 tropism|HIV 1 tropism
C4069288|T201|COMP|79768-8|LNC|Platelet dense bodies|Platelet dense bodies
C4069290|T201|COMP|79623-5|LNC|Alpha aminoisobutyrate/Creatinine|Alpha aminoisobutyrate/Creatinine
C4069292|T201|COMP|79512-0|LNC|Vanilloylglycine|Vanilloylglycine
C4069293|T201|COMP|79476-8|LNC|Ethylmalonate|Ethylmalonate
C4069294|T201|COMP|79495-8|LNC|Azelate|Azelate
C4069295|T201|COMP|78991-7|LNC|Flavin adenine dinucleotide|Flavin adenine dinucleotide
C4069296|T201|COMP|79299-4|LNC|D- & L-2-hydroxyglutarate pattern|D- & L-2-hydroxyglutarate pattern
C4069297|T201|COMP|79284-6|LNC|Carnitine biosynthesis intermediates panel|Carnitine biosynthesis intermediates panel
C4069298|T201|COMP|78963-6|LNC|Mannose-6-phosphate isomerase|Mannose-6-phosphate isomerase
C4069299|T201|COMP|78887-7|LNC|Trans-3-Hydroxycotinine|Trans-3-Hydroxycotinine
C4069300|T201|COMP|79162-4|LNC|Chlordiazepoxide & Norchlordiazepoxide panel|Chlordiazepoxide & Norchlordiazepoxide panel
C4069301|T201|COMP|79648-2|LNC|D-serine|D-serine
C4069303|T201|COMP|78780-4|LNC|Alminoprofen|Alminoprofen
C4069304|T201|COMP|78747-3|LNC|Peritoneal equilibration test panel|Peritoneal equilibration test panel
C4069316|T201|COMP|80123-3|LNC|Alizapride|Alizapride
C4069366|T201|COMP|80426-0|LNC|Hepatitis D virus RNA|Hepatitis D virus RNA
C4069367|T201|COMP|80425-2|LNC|Beta-N-acetylhexosaminidase.A|Beta-N-acetylhexosaminidase.A
C4069368|T201|COMP|80424-5|LNC|Inosine triphosphate pyrophosphatase|Inosine triphosphate pyrophosphatase
C4069384|T201|COMP|80398-1|LNC|Unique identifier|Unique identifier
C4069391|T201|COMP|80382-5|LNC|Influenza virus A Ag|Influenza virus A Ag
C4069392|T201|COMP|80381-7|LNC|Influenza virus A & B Ag panel|Influenza virus A & B Ag panel
C4069393|T201|COMP|80373-4|LNC|Helicobacter pylori Ag|Helicobacter pylori Ag
C4069394|T201|COMP|80372-6|LNC|Hemoglobin.gastrointestinal|Hemoglobin.gastrointestinal
C4069395|T201|COMP|80371-8|LNC|Chitotriosidase|Chitotriosidase
C4069396|T201|COMP|80370-0|LNC|Biotinidase|Biotinidase
C4069397|T201|COMP|80369-2|LNC|Neisseria sp identified|Neisseria sp identified
C4069398|T201|COMP|80368-4|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C4069399|T201|COMP|80367-6|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C4069400|T201|COMP|80366-8|LNC|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C4069401|T201|COMP|80365-0|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C4069402|T201|COMP|80364-3|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C4069403|T201|COMP|80363-5|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C4069404|T201|COMP|80362-7|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C4069405|T201|COMP|80361-9|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C4069406|T201|COMP|80360-1|LNC|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C4069412|T201|COMP|80354-4|LNC|Herpes simplex virus 1 & 2 DNA panel|Herpes simplex virus 1 & 2 DNA panel
C4069417|T201|COMP|80348-6|LNC|Escherichia coli enteropathogenic eae gene|Escherichia coli enteropathogenic eae gene
C4069447|T201|COMP|80244-7|LNC|Mycoplasma hyopneumoniae DNA|Mycoplasma hyopneumoniae DNA
C4069464|T201|COMP|80223-1|LNC|Cells.CD4/100 lymphocytes|Cells.CD4/100 lymphocytes
C4069465|T201|COMP|80222-3|LNC|Cells.CD8/100 lymphocytes|Cells.CD8/100 lymphocytes
C4069466|T201|COMP|80221-5|LNC|N-methyl-D-aspartate receptor Ab.IgG|N-methyl-D-aspartate receptor Ab.IgG
C4069467|T201|COMP|80220-7|LNC|N-methyl-D-aspartate receptor Ab.IgG|N-methyl-D-aspartate receptor Ab.IgG
C4069469|T201|COMP|80218-1|LNC|Mycoplasma hyopneumoniae Ab sample/Buffer control|Mycoplasma hyopneumoniae Ab sample/Buffer control
C4069470|T201|COMP|80217-3|LNC|Mycoplasma hyopneumoniae Ag|Mycoplasma hyopneumoniae Ag
C4069472|T201|COMP|80215-7|LNC|Beta blockers|Beta blockers
C4069473|T201|COMP|80214-0|LNC|Beta blockers|Beta blockers
C4069474|T201|COMP|80213-2|LNC|Beta blockers|Beta blockers
C4069475|T201|COMP|80212-4|LNC|Beta blockers|Beta blockers
C4069476|T201|COMP|80211-6|LNC|Beryllium|Beryllium
C4069477|T201|COMP|80210-8|LNC|Beryllium|Beryllium
C4069478|T201|COMP|80209-0|LNC|Barium|Barium
C4069479|T201|COMP|80208-2|LNC|Leishmania infantum+donovani Ab.IgG|Leishmania infantum+donovani Ab.IgG
C4069480|T201|COMP|80207-4|LNC|Leishmania infantum+donovani Ab.IgM|Leishmania infantum+donovani Ab.IgM
C4069483|T201|COMP|80204-1|LNC|Influenza virus A & B identified|Influenza virus A & B identified
C4069484|T201|COMP|80203-3|LNC|HIV 1 & 2 Ab|HIV 1 & 2 Ab
C4069485|T201|COMP|80201-7|LNC|Alizapride|Alizapride
C4069486|T201|COMP|80200-9|LNC|Nonsteroidal antiinflammatory drugs|Nonsteroidal antiinflammatory drugs
C4069487|T201|COMP|80199-3|LNC|Nonsteroidal antiinflammatory drugs|Nonsteroidal antiinflammatory drugs
C4069488|T201|COMP|80198-5|LNC|Nonsteroidal antiinflammatory drugs|Nonsteroidal antiinflammatory drugs
C4069489|T201|COMP|80197-7|LNC|Antihistamines|Antihistamines
C4069490|T201|COMP|80196-9|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C4069491|T201|COMP|80195-1|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C4069492|T201|COMP|80194-4|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C4069493|T201|COMP|80193-6|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C4069495|T201|COMP|80189-4|LNC|Galactosamine|Galactosamine
C4069496|T201|COMP|80188-6|LNC|JAK2 gene exon 14 targeted mutation analysis|JAK2 gene exon 14 targeted mutation analysis
C4069497|T201|COMP|80187-8|LNC|JAK2 gene exon 14 targeted mutation analysis|JAK2 gene exon 14 targeted mutation analysis
C4069498|T201|COMP|80186-0|LNC|JAK2 gene exon 12 targeted mutation analysis|JAK2 gene exon 12 targeted mutation analysis
C4069499|T201|COMP|80185-2|LNC|Xanthopterin/Creatinine|Xanthopterin/Creatinine
C4069500|T201|COMP|80184-5|LNC|Xanthopterin|Xanthopterin
C4069501|T201|COMP|80183-7|LNC|Xanthopterin|Xanthopterin
C4069502|T201|COMP|80182-9|LNC|S-adenosylmethionine/Creatinine|S-adenosylmethionine/Creatinine
C4069507|T201|COMP|80177-9|LNC|S-adenosylmethionine|S-adenosylmethionine
C4069508|T201|COMP|80176-1|LNC|S-adenosylhomocysteine/Creatinine|S-adenosylhomocysteine/Creatinine
C4069509|T201|COMP|80175-3|LNC|S-adenosylhomocysteine|S-adenosylhomocysteine
C4069510|T201|COMP|80174-6|LNC|S-adenosylhomocysteine|S-adenosylhomocysteine
C4069511|T201|COMP|80173-8|LNC|Pterins pattern|Pterins pattern
C4069512|T201|COMP|80172-0|LNC|Pterins pattern|Pterins pattern
C4069513|T201|COMP|80171-2|LNC|Pterins pattern|Pterins pattern
C4069514|T201|COMP|80170-4|LNC|Pterins panel|Pterins panel
C4069515|T201|COMP|80169-6|LNC|Pterins panel|Pterins panel
C4069516|T201|COMP|80168-8|LNC|Pterins panel|Pterins panel
C4069517|T201|COMP|80167-0|LNC|2-Amino-4-hydroxypteridine/Creatinine|2-Amino-4-hydroxypteridine/Creatinine
C4069518|T201|COMP|80166-2|LNC|2-Amino-4-hydroxypteridine|2-Amino-4-hydroxypteridine
C4069519|T201|COMP|80165-4|LNC|2-Amino-4-hydroxypteridine|2-Amino-4-hydroxypteridine
C4069520|T201|COMP|80164-7|LNC|Bile alcohols pattern|Bile alcohols pattern
C4069521|T201|COMP|80163-9|LNC|Bile alcohols panel|Bile alcohols panel
C4069522|T201|COMP|80162-1|LNC|Bile alcohols|Bile alcohols
C4069525|T201|COMP|80159-7|LNC|27-Norcholestanehexol/Creatinine|27-Norcholestanehexol/Creatinine
C4069526|T201|COMP|80158-9|LNC|Galactosylhydroxylysine/Creatinine|Galactosylhydroxylysine/Creatinine
C4069527|T201|COMP|80157-1|LNC|Etiocholanolone|Etiocholanolone
C4069528|T201|COMP|80156-3|LNC|3-Methoxytyramine/Creatinine|3-Methoxytyramine/Creatinine
C4069529|T201|COMP|80155-5|LNC|Soluble CD27|Soluble CD27
C4069535|T201|COMP|80387-4|LNC|HIV 1+2 Ab|HIV 1+2 Ab
C4069536|T201|COMP|80386-6|LNC|Bladder tumor Ag|Bladder tumor Ag
C4069537|T201|COMP|80385-8|LNC|Choriogonadotropin (pregnancy test)|Choriogonadotropin (pregnancy test)
C4069538|T201|COMP|80384-1|LNC|Choriogonadotropin (pregnancy test)|Choriogonadotropin (pregnancy test)
C4069539|T201|COMP|80383-3|LNC|Influenza virus B Ag|Influenza virus B Ag
C4069545|T201|COMP|80154-8|LNC|Monolysocardiolipin/cardiolipin|Monolysocardiolipin/cardiolipin
C4069546|T201|COMP|80153-0|LNC|Soluble CD27|Soluble CD27
C4069547|T201|COMP|80152-2|LNC|N-methylhistamine/Creatinine|N-methylhistamine/Creatinine
C4069548|T201|COMP|80151-4|LNC|Brucella abortus Ab.IgG|Brucella abortus Ab.IgG
C4069549|T201|COMP|80150-6|LNC|Trimeprazine|Trimeprazine
C4069550|T201|COMP|80149-8|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C4069551|T201|COMP|80148-0|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C4069552|T201|COMP|80147-2|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C4069553|T201|COMP|80146-4|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C4069554|T201|COMP|80145-6|LNC|Silver|Silver
C4069555|T201|COMP|80144-9|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C4069556|T201|COMP|80143-1|LNC|Atazanavir|Atazanavir
C4069557|T201|COMP|80142-3|LNC|Atazanavir|Atazanavir
C4069558|T201|COMP|80141-5|LNC|Arsenic|Arsenic
C4069559|T201|COMP|80140-7|LNC|Antimony|Antimony
C4069560|T201|COMP|80139-9|LNC|Antimony|Antimony
C4069561|T201|COMP|80138-1|LNC|Antimony|Antimony
C4069562|T201|COMP|80137-3|LNC|Antihistamines|Antihistamines
C4069563|T201|COMP|80136-5|LNC|Antihistamines|Antihistamines
C4069564|T201|COMP|80135-7|LNC|Amphetamine|Amphetamine
C4069565|T201|COMP|80134-0|LNC|Amphetamine|Amphetamine
C4069566|T201|COMP|80133-2|LNC|Amoxicillin|Amoxicillin
C4069567|T201|COMP|80132-4|LNC|amLODIPine|amLODIPine
C4069568|T201|COMP|80131-6|LNC|Amisulpride|Amisulpride
C4069569|T201|COMP|80130-8|LNC|Amisulpride|Amisulpride
C4069570|T201|COMP|80129-0|LNC|Amisulpride|Amisulpride
C4069571|T201|COMP|80128-2|LNC|Amisulpride|Amisulpride
C4069572|T201|COMP|80127-4|LNC|Aluminum|Aluminum
C4069573|T201|COMP|80126-6|LNC|Aluminum|Aluminum
C4069574|T201|COMP|80125-8|LNC|Aluminum|Aluminum
C4069575|T201|COMP|80124-1|LNC|Alminoprofen|Alminoprofen
C4069576|T201|COMP|80122-5|LNC|Alfentanil|Alfentanil
C4069577|T201|COMP|80121-7|LNC|Acyclovir|Acyclovir
C4069578|T201|COMP|80120-9|LNC|Acenocoumarol|Acenocoumarol
C4069579|T201|COMP|80119-1|LNC|Acebutolol|Acebutolol
C4069580|T201|COMP|80118-3|LNC|Abacavir|Abacavir
C4069581|T201|COMP|80117-5|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C4069582|T201|COMP|80116-7|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C4069583|T201|COMP|80115-9|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C4069584|T201|COMP|80114-2|LNC|2-Oxo-3-Hydroxy-Lysergate diethylamide|2-Oxo-3-Hydroxy-Lysergate diethylamide
C4069585|T201|COMP|80113-4|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C4069586|T201|COMP|80112-6|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C4069587|T201|COMP|80111-8|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C4069598|T201|COMP|80100-1|LNC|D-2-hydroxyglutarate/Creatinine|D-2-hydroxyglutarate/Creatinine
C4069599|T201|COMP|80099-5|LNC|L-2-hydroxyglutarate/Creatinine|L-2-hydroxyglutarate/Creatinine
C4069600|T201|COMP|80098-7|LNC|Glucosamine/Creatinine|Glucosamine/Creatinine
C4069601|T201|COMP|80097-9|LNC|Glycyl-4-hydroxyproline|Glycyl-4-hydroxyproline
C4069602|T201|COMP|80096-1|LNC|Glutamylphenylalanine|Glutamylphenylalanine
C4069603|T201|COMP|80095-3|LNC|Galactosamine/Creatinine|Galactosamine/Creatinine
C4069604|T201|COMP|80094-6|LNC|Glutamylphenylalanine/Creatinine|Glutamylphenylalanine/Creatinine
C4069605|T201|COMP|80093-8|LNC|Glucosamine|Glucosamine
C4069606|T201|COMP|80092-0|LNC|Glycyl-4-hydroxyproline/Creatinine|Glycyl-4-hydroxyproline/Creatinine
C4069927|T201|COMP|79722-5|LNC|SLCO1B1 gene product functional interpretation|SLCO1B1 gene product functional interpretation
C4069934|T201|COMP|79712-6|LNC|HLA-A*31:01|HLA-A*31:01
C4069935|T201|COMP|79711-8|LNC|HLA-B*58:01|HLA-B*58:01
C4069936|T201|COMP|79710-0|LNC|Potassium|Potassium
C4069937|T201|COMP|79709-2|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C4069938|T201|COMP|79708-4|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C4069939|T201|COMP|79707-6|LNC|Fatty acids.very long chain.C26:1/C22:0|Fatty acids.very long chain.C26:1/C22:0
C4069940|T201|COMP|79706-8|LNC|Octadecatetraenoate|Octadecatetraenoate
C4069941|T201|COMP|79705-0|LNC|Eicosadienoate|Eicosadienoate
C4069942|T201|COMP|79704-3|LNC|Homo-gamma linolenate|Homo-gamma linolenate
C4069943|T201|COMP|79703-5|LNC|cis-13-Eicosenoate|cis-13-Eicosenoate
C4069944|T201|COMP|79702-7|LNC|cis-13-Eicosenoate|cis-13-Eicosenoate
C4069945|T201|COMP|79701-9|LNC|Fatty acids.very long chain.C22:1n9|Fatty acids.very long chain.C22:1n9
C4069946|T201|COMP|79700-1|LNC|cis-11,14-Eicosadienoate|cis-11,14-Eicosadienoate
C4069947|T201|COMP|79699-5|LNC|cis-11-Eicosenoate|cis-11-Eicosenoate
C4069948|T201|COMP|79698-7|LNC|Docosadienoate|Docosadienoate
C4069949|T201|COMP|79697-9|LNC|Docosadienoate|Docosadienoate
C4069950|T201|COMP|79696-1|LNC|cis-11-Eicosenoate|cis-11-Eicosenoate
C4069951|T201|COMP|79695-3|LNC|Octadecatetraenoate|Octadecatetraenoate
C4069952|T201|COMP|79694-6|LNC|Eicosadienoate|Eicosadienoate
C4069953|T201|COMP|79693-8|LNC|5,6-Dihydrouracil|5,6-Dihydrouracil
C4069954|T201|COMP|79692-0|LNC|2,8-Dihydroxyadenine|2,8-Dihydroxyadenine
C4069955|T201|COMP|79691-2|LNC|Oxipurinol|Oxipurinol
C4069956|T201|COMP|79690-4|LNC|Guanine|Guanine
C4069957|T201|COMP|79689-6|LNC|Allopurinol|Allopurinol
C4069958|T201|COMP|79688-8|LNC|5-hydroxymethyluracil|5-hydroxymethyluracil
C4069959|T201|COMP|79687-0|LNC|2,8-Dihydroxyadenine/Creatinine|2,8-Dihydroxyadenine/Creatinine
C4069960|T201|COMP|79686-2|LNC|5-hydroxymethyluracil|5-hydroxymethyluracil
C4069961|T201|COMP|79685-4|LNC|5,6-Dihydrouracil/Creatinine|5,6-Dihydrouracil/Creatinine
C4069962|T201|COMP|79684-7|LNC|Cytidine/Creatinine|Cytidine/Creatinine
C4069963|T201|COMP|79683-9|LNC|Cytosine|Cytosine
C4069964|T201|COMP|79682-1|LNC|5,6-Dihydrouracil|5,6-Dihydrouracil
C4069965|T201|COMP|79681-3|LNC|Allopurinol/Creatinine|Allopurinol/Creatinine
C4069966|T201|COMP|79680-5|LNC|2,8-Dihydroxyadenine|2,8-Dihydroxyadenine
C4069967|T201|COMP|79679-7|LNC|5-Aminoimidazole-4-carboxamide|5-Aminoimidazole-4-carboxamide
C4069968|T201|COMP|79678-9|LNC|5,6-Dihydrouridine/Creatinine|5,6-Dihydrouridine/Creatinine
C4069969|T201|COMP|79677-1|LNC|Purine & Pyrimidine pattern|Purine & Pyrimidine pattern
C4069970|T201|COMP|79676-3|LNC|5,6-Dihydrouridine|5,6-Dihydrouridine
C4069971|T201|COMP|79675-5|LNC|Cytidine|Cytidine
C4069972|T201|COMP|79674-8|LNC|Pseudouridine|Pseudouridine
C4069973|T201|COMP|79673-0|LNC|Purine & Pyrimidine panel|Purine & Pyrimidine panel
C4069974|T201|COMP|79672-2|LNC|5-Aminoimidazole-4-carboxamide/Creatinine|5-Aminoimidazole-4-carboxamide/Creatinine
C4069975|T201|COMP|79671-4|LNC|Cytidine|Cytidine
C4069976|T201|COMP|79670-6|LNC|Guanosine|Guanosine
C4069977|T201|COMP|79669-8|LNC|Dihydrothymine|Dihydrothymine
C4069978|T201|COMP|79668-0|LNC|Purine & Pyrimidine panel|Purine & Pyrimidine panel
C4069979|T201|COMP|79667-2|LNC|5,6-Dihydrouridine|5,6-Dihydrouridine
C4069980|T201|COMP|79666-4|LNC|Purine & Pyrimidine pattern|Purine & Pyrimidine pattern
C4069981|T201|COMP|79665-6|LNC|Purine & Pyrimidine panel|Purine & Pyrimidine panel
C4069982|T201|COMP|79664-9|LNC|N-carbamoyl beta alanine|N-carbamoyl beta alanine
C4069983|T201|COMP|79663-1|LNC|Guanine|Guanine
C4069984|T201|COMP|79662-3|LNC|Allopurinol|Allopurinol
C4069985|T201|COMP|79661-5|LNC|Dihydroorotate|Dihydroorotate
C4069986|T201|COMP|79660-7|LNC|Guanosine|Guanosine
C4069987|T201|COMP|79659-9|LNC|Purine & Pyrimidine pattern|Purine & Pyrimidine pattern
C4069988|T201|COMP|79658-1|LNC|Cytosine/Creatinine|Cytosine/Creatinine
C4069989|T201|COMP|79657-3|LNC|Pseudouridine|Pseudouridine
C4069990|T201|COMP|79656-5|LNC|N-carbamoyl beta alanine|N-carbamoyl beta alanine
C4069991|T201|COMP|79655-7|LNC|Cytosine|Cytosine
C4069992|T201|COMP|79654-0|LNC|Dihydroorotate|Dihydroorotate
C4069993|T201|COMP|79653-2|LNC|Dihydroorotate|Dihydroorotate
C4069994|T201|COMP|79652-4|LNC|5-Aminoimidazole-4-carboxamide|5-Aminoimidazole-4-carboxamide
C4069995|T201|COMP|79651-6|LNC|Dihydrothymine|Dihydrothymine
C4069997|T201|COMP|79639-1|LNC|N,N'-dimethylarginine/Creatinine|N,N'-dimethylarginine/Creatinine
C4069999|T201|COMP|79637-5|LNC|Glutathione.oxidized/Creatinine|Glutathione.oxidized/Creatinine
C4070000|T201|COMP|79636-7|LNC|Aspartylglycosamine/Creatinine|Aspartylglycosamine/Creatinine
C4070001|T201|COMP|79635-9|LNC|N,N-dimethylarginine/Creatinine|N,N-dimethylarginine/Creatinine
C4070002|T201|COMP|79634-2|LNC|N6-Acetyl-L-lysine/Creatinine|N6-Acetyl-L-lysine/Creatinine
C4070003|T201|COMP|79633-4|LNC|L-leucyl-L-proline|L-leucyl-L-proline
C4070004|T201|COMP|79632-6|LNC|Homocarnosine/Creatinine|Homocarnosine/Creatinine
C4070005|T201|COMP|79631-8|LNC|L-homoserine|L-homoserine
C4070007|T201|COMP|79629-2|LNC|R-beta aminoisobutyrate|R-beta aminoisobutyrate
C4070008|T201|COMP|79628-4|LNC|Formiminoglutamate|Formiminoglutamate
C4070009|T201|COMP|79627-6|LNC|N-alpha acetyllysine/Creatinine|N-alpha acetyllysine/Creatinine
C4070010|T201|COMP|79626-8|LNC|L-leucyl-L-proline/Creatinine|L-leucyl-L-proline/Creatinine
C4070011|T201|COMP|79625-0|LNC|Aspartylglycine/Creatinine|Aspartylglycine/Creatinine
C4070012|T201|COMP|79624-3|LNC|5-S-cysteinyldopa|5-S-cysteinyldopa
C4070013|T201|COMP|79622-7|LNC|R-beta aminoisobutyrate/Creatinine|R-beta aminoisobutyrate/Creatinine
C4070014|T201|COMP|79621-9|LNC|Phenylalanine & Tyrosine panel|Phenylalanine & Tyrosine panel
C4070015|T201|COMP|79620-1|LNC|Formiminoglutamate/Creatinine|Formiminoglutamate/Creatinine
C4070016|T201|COMP|79619-3|LNC|S-beta aminoisobutyrate/Creatinine|S-beta aminoisobutyrate/Creatinine
C4070017|T201|COMP|79611-0|LNC|Prolylhydroxyproline/Creatinine|Prolylhydroxyproline/Creatinine
C4070018|T201|COMP|79610-2|LNC|D-serine|D-serine
C4070019|T201|COMP|79609-4|LNC|Glutathione.oxidized|Glutathione.oxidized
C4070020|T201|COMP|79608-6|LNC|2-Methyltyrosine|2-Methyltyrosine
C4070021|T201|COMP|79607-8|LNC|Saccharopine|Saccharopine
C4070022|T201|COMP|79606-0|LNC|Cysteate|Cysteate
C4070024|T201|COMP|79604-5|LNC|S-beta aminoisobutyrate|S-beta aminoisobutyrate
C4070026|T201|COMP|79602-9|LNC|Homocarnosine|Homocarnosine
C4070027|T201|COMP|79601-1|LNC|L-serine|L-serine
C4070028|T201|COMP|79600-3|LNC|Glutathione.reduced|Glutathione.reduced
C4070029|T201|COMP|79599-7|LNC|Cysteate/Creatinine|Cysteate/Creatinine
C4070031|T201|COMP|79597-1|LNC|N-monomethylarginine/Creatinine|N-monomethylarginine/Creatinine
C4070032|T201|COMP|79596-3|LNC|D-serine/Creatinine|D-serine/Creatinine
C4070033|T201|COMP|79595-5|LNC|N,N'-dimethylarginine|N,N'-dimethylarginine
C4070034|T201|COMP|79594-8|LNC|Glycylproline/Creatinine|Glycylproline/Creatinine
C4070035|T201|COMP|79593-0|LNC|Allocystathionine/Creatinine|Allocystathionine/Creatinine
C4070036|T201|COMP|79592-2|LNC|Homocitrulline/Creatinine|Homocitrulline/Creatinine
C4070037|T201|COMP|79591-4|LNC|N-alpha acetyllysine|N-alpha acetyllysine
C4070038|T201|COMP|79590-6|LNC|Alpha aminoisobutyrate|Alpha aminoisobutyrate
C4070039|T201|COMP|79589-8|LNC|Aspartylglycosamine|Aspartylglycosamine
C4070040|T201|COMP|79588-0|LNC|Prolylhydroxyproline|Prolylhydroxyproline
C4070041|T201|COMP|79587-2|LNC|L-homoarginine/Creatinine|L-homoarginine/Creatinine
C4070043|T201|COMP|79585-6|LNC|Aspartylglycine|Aspartylglycine
C4070046|T201|COMP|79582-3|LNC|Beta-ureidoisobutyrate|Beta-ureidoisobutyrate
C4070047|T201|COMP|79581-5|LNC|Alanylproline|Alanylproline
C4070049|T201|COMP|79579-9|LNC|Alanylproline/Creatinine|Alanylproline/Creatinine
C4070050|T201|COMP|79578-1|LNC|N6-Acetyl-L-lysine|N6-Acetyl-L-lysine
C4070051|T201|COMP|79577-3|LNC|Levodopa/Creatinine|Levodopa/Creatinine
C4070052|T201|COMP|79576-5|LNC|Allocystathionine|Allocystathionine
C4070054|T201|COMP|79574-0|LNC|Folate & tryptophan & metabolites pattern|Folate & tryptophan & metabolites pattern
C4070056|T201|COMP|79572-4|LNC|Folate & tryptophan & metabolites panel|Folate & tryptophan & metabolites panel
C4070057|T201|COMP|79571-6|LNC|BCHE gene full mutation analysis|BCHE gene full mutation analysis
C4070060|T201|COMP|79567-4|LNC|Lysophosphatidylcholine(26:0)|Lysophosphatidylcholine(26:0)
C4070061|T201|COMP|79566-6|LNC|Collection method|Collection method
C4070062|T201|COMP|79564-1|LNC|Mucopolysaccharidosis type I|Mucopolysaccharidosis type I
C4070078|T201|COMP|79538-5|LNC|Formate|Formate
C4070088|T201|COMP|79528-6|LNC|5-Hydroxymethyl-2-Furoate|5-Hydroxymethyl-2-Furoate
C4070089|T201|COMP|79527-8|LNC|4-Deoxythreonate/Creatinine|4-Deoxythreonate/Creatinine
C4070090|T201|COMP|79526-0|LNC|3,5-Dihydroxybenzoate|3,5-Dihydroxybenzoate
C4070091|T201|COMP|79525-2|LNC|3-Hydroxysebacate.unsaturated|3-Hydroxysebacate.unsaturated
C4070092|T201|COMP|79524-5|LNC|P-cresol|P-cresol
C4070093|T201|COMP|79523-7|LNC|3-(3-Hydroxyphenyl)propanoate|3-(3-Hydroxyphenyl)propanoate
C4070094|T201|COMP|79522-9|LNC|2,5-Furandicarboxylate/Creatinine|2,5-Furandicarboxylate/Creatinine
C4070095|T201|COMP|79521-1|LNC|Lactyl lactate|Lactyl lactate
C4070096|T201|COMP|79520-3|LNC|4-Deoxythreonate|4-Deoxythreonate
C4070097|T201|COMP|79519-5|LNC|Pimelate|Pimelate
C4070098|T201|COMP|79518-7|LNC|3-Hydroxybenzoate/Creatinine|3-Hydroxybenzoate/Creatinine
C4070099|T201|COMP|79517-9|LNC|Desaminotyrosine/Creatinine|Desaminotyrosine/Creatinine
C4070100|T201|COMP|79516-1|LNC|Octenedioate|Octenedioate
C4070101|T201|COMP|79515-3|LNC|Gentisate|Gentisate
C4070102|T201|COMP|79514-6|LNC|N-acetyltyrosine|N-acetyltyrosine
C4070103|T201|COMP|79513-8|LNC|1,4-Cyclohexanediol|1,4-Cyclohexanediol
C4070104|T201|COMP|79511-2|LNC|Suberylglycine|Suberylglycine
C4070105|T201|COMP|79510-4|LNC|3-Hydroxyhippurate|3-Hydroxyhippurate
C4070106|T201|COMP|79509-6|LNC|Decenedioate|Decenedioate
C4070107|T201|COMP|79508-8|LNC|4-Hydroxymandelate|4-Hydroxymandelate
C4070108|T201|COMP|79507-0|LNC|P-cresol/Creatinine|P-cresol/Creatinine
C4070109|T201|COMP|79506-2|LNC|Desaminotyrosine|Desaminotyrosine
C4070110|T201|COMP|79505-4|LNC|4-Hydroxy-3-Methoxyphenyllactate|4-Hydroxy-3-Methoxyphenyllactate
C4070111|T201|COMP|79504-7|LNC|Levulinate/Creatinine|Levulinate/Creatinine
C4070112|T201|COMP|79503-9|LNC|4-Hydroxyhippurate|4-Hydroxyhippurate
C4070113|T201|COMP|79502-1|LNC|4-Hydroxyvalerate|4-Hydroxyvalerate
C4070114|T201|COMP|79501-3|LNC|3-Hydroxyhippurate/Creatinine|3-Hydroxyhippurate/Creatinine
C4070115|T201|COMP|79500-5|LNC|Furoylglycine/Creatinine|Furoylglycine/Creatinine
C4070116|T201|COMP|79499-0|LNC|Catecholamine metabolites panel|Catecholamine metabolites panel
C4070117|T201|COMP|79498-2|LNC|4-Hydroxyhippurate/Creatinine|4-Hydroxyhippurate/Creatinine
C4070118|T201|COMP|79497-4|LNC|3-Hydroxybenzoate|3-Hydroxybenzoate
C4070119|T201|COMP|79496-6|LNC|Hydantoin-5-propionate|Hydantoin-5-propionate
C4070120|T201|COMP|79484-2|LNC|Levulinate|Levulinate
C4070121|T201|COMP|79483-4|LNC|Vanilloylglycine/Creatinine|Vanilloylglycine/Creatinine
C4070122|T201|COMP|79482-6|LNC|3-(3-Hydroxyphenyl)propanoate/Creatinine|3-(3-Hydroxyphenyl)propanoate/Creatinine
C4070123|T201|COMP|79481-8|LNC|Hydantoin-5-propionate/Creatinine|Hydantoin-5-propionate/Creatinine
C4070124|T201|COMP|79480-0|LNC|3,4-Dihydroxyhydrocinnamate|3,4-Dihydroxyhydrocinnamate
C4070125|T201|COMP|79479-2|LNC|3-Hydroxyadipate 3,6-lactone|3-Hydroxyadipate 3,6-lactone
C4070126|T201|COMP|79478-4|LNC|Salicylurate/Creatinine|Salicylurate/Creatinine
C4070127|T201|COMP|79477-6|LNC|5-Hydroxymethyl-2-Furoate/Creatinine|5-Hydroxymethyl-2-Furoate/Creatinine
C4070128|T201|COMP|79475-0|LNC|2,5-Furandicarboxylate|2,5-Furandicarboxylate
C4070129|T201|COMP|79474-3|LNC|3,4-Dihydroxybutyrate/Creatinine|3,4-Dihydroxybutyrate/Creatinine
C4070130|T201|COMP|79473-5|LNC|Hexanoylglycine|Hexanoylglycine
C4070131|T201|COMP|79472-7|LNC|Phenylpropionylglycine|Phenylpropionylglycine
C4070132|T201|COMP|79471-9|LNC|1,4-Cyclohexanediol/Creatinine|1,4-Cyclohexanediol/Creatinine
C4070133|T201|COMP|79470-1|LNC|Uridine monophosphate synthetase|Uridine monophosphate synthetase
C4070134|T201|COMP|79469-3|LNC|Uridine diphosphate glucose-4-Epimerase|Uridine diphosphate glucose-4-Epimerase
C4070135|T201|COMP|79468-5|LNC|Thiopurine methyltransferase|Thiopurine methyltransferase
C4070136|T201|COMP|79467-7|LNC|Purine nucleoside phosphorylase|Purine nucleoside phosphorylase
C4070137|T201|COMP|79466-9|LNC|Purine nucleoside phosphorylase|Purine nucleoside phosphorylase
C4070138|T201|COMP|79465-1|LNC|Porphobilinogen synthase|Porphobilinogen synthase
C4070139|T201|COMP|79464-4|LNC|Phosphorylase|Phosphorylase
C4070140|T201|COMP|79463-6|LNC|N-Acetylgalactosamine-4-Sulfatase|N-Acetylgalactosamine-4-Sulfatase
C4070141|T201|COMP|79462-8|LNC|Iduronate-2-Sulfatase|Iduronate-2-Sulfatase
C4070142|T201|COMP|79461-0|LNC|Hypoxanthine phosphoribosyltransferase|Hypoxanthine phosphoribosyltransferase
C4070143|T201|COMP|79460-2|LNC|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C4070144|T201|COMP|79459-4|LNC|Dihydropteridine reductase|Dihydropteridine reductase
C4070145|T201|COMP|79458-6|LNC|Beta-N-acetylhexosaminidase|Beta-N-acetylhexosaminidase
C4070146|T201|COMP|79457-8|LNC|Beta glucuronidase|Beta glucuronidase
C4070147|T201|COMP|79456-0|LNC|Arginase|Arginase
C4070148|T201|COMP|79455-2|LNC|Alpha-N-acetylgalactosaminidase|Alpha-N-acetylgalactosaminidase
C4070149|T201|COMP|79454-5|LNC|Alpha fucosidase|Alpha fucosidase
C4070150|T201|COMP|79453-7|LNC|Alcohol dehydrogenase|Alcohol dehydrogenase
C4070151|T201|COMP|79452-9|LNC|Adenylosuccinate lyase|Adenylosuccinate lyase
C4070152|T201|COMP|79451-1|LNC|Adenosine deaminase|Adenosine deaminase
C4070153|T201|COMP|79450-3|LNC|Adenine phosphoribosyltransferase|Adenine phosphoribosyltransferase
C4070154|T201|COMP|79449-5|LNC|Formate|Formate
C4070157|T201|COMP|79446-1|LNC|Pericyazine|Pericyazine
C4070158|T201|COMP|79445-3|LNC|Fluspirilene|Fluspirilene
C4070193|T201|COMP|79644-1|LNC|L-homoserine/Creatinine|L-homoserine/Creatinine
C4070194|T201|COMP|79643-3|LNC|5-S-cysteinyldopa/Creatinine|5-S-cysteinyldopa/Creatinine
C4070196|T201|COMP|79641-7|LNC|Glutathione.reduced/Creatinine|Glutathione.reduced/Creatinine
C4070197|T201|COMP|79640-9|LNC|Saccharopine/Creatinine|Saccharopine/Creatinine
C4070198|T201|COMP|79494-1|LNC|Pimelate/Creatinine|Pimelate/Creatinine
C4070199|T201|COMP|79493-3|LNC|3-Hydroxysuberate.unsaturated|3-Hydroxysuberate.unsaturated
C4070200|T201|COMP|79492-5|LNC|Furoylglycine|Furoylglycine
C4070201|T201|COMP|79491-7|LNC|3-Hydroxyphenylacetate|3-Hydroxyphenylacetate
C4070202|T201|COMP|79427-1|LNC|Platelets|Platelets
C4070203|T201|COMP|79426-3|LNC|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C4070204|T201|COMP|79425-5|LNC|Bacteria identified|Bacteria identified
C4070209|T201|COMP|79420-6|LNC|Allergen.miscellaneous Ab.IgE|Allergen.miscellaneous Ab.IgE
C4070211|T201|COMP|79418-0|LNC|EPCAM gene exons 8 & 9 deletion+duplication|EPCAM gene exons 8 & 9 deletion+duplication
C4070212|T201|COMP|79417-2|LNC|PMS2 gene deletion+duplication|PMS2 gene deletion+duplication
C4070213|T201|COMP|79416-4|LNC|MLH1 gene deletion+duplication|MLH1 gene deletion+duplication
C4070214|T201|COMP|79415-6|LNC|MSH2 gene deletion+duplication|MSH2 gene deletion+duplication
C4070215|T201|COMP|79414-9|LNC|MSH6 gene deletion+duplication|MSH6 gene deletion+duplication
C4070216|T201|COMP|79413-1|LNC|Dothiepin+Nordothiepin^trough|Dothiepin+Nordothiepin^trough
C4070217|T201|COMP|79412-3|LNC|Mianserin trough & Normianserin panel|Mianserin trough & Normianserin panel
C4070218|T201|COMP|79411-5|LNC|Creatine transport protein|Creatine transport protein
C4070219|T201|COMP|79410-7|LNC|Penfluridol^trough|Penfluridol^trough
C4070221|T201|COMP|79408-1|LNC|Clobazam & norclobazam panel|Clobazam & norclobazam panel
C4070222|T201|COMP|79407-3|LNC|Catecholamine metabolites pattern|Catecholamine metabolites pattern
C4070223|T201|COMP|79406-5|LNC|IgM clearance/Albumin clearance|IgM clearance/Albumin clearance
C4070224|T201|COMP|79405-7|LNC|1,4-Alpha glucan branching enzyme|1,4-Alpha glucan branching enzyme
C4070225|T201|COMP|79404-0|LNC|Adenosine deaminase|Adenosine deaminase
C4070226|T201|COMP|79403-2|LNC|Nitrogen|Nitrogen
C4070227|T201|COMP|79402-4|LNC|Niacin|Niacin
C4070228|T201|COMP|79400-8|LNC|Vanillylmandelate|Vanillylmandelate
C4070229|T201|COMP|79399-2|LNC|Synovial fluid analysis panel|Synovial fluid analysis panel
C4070230|T201|COMP|79398-4|LNC|Prolactin isoforms pattern|Prolactin isoforms pattern
C4070231|T201|COMP|79397-6|LNC|Pistacia lentiscus Ab.IgE|Pistacia lentiscus Ab.IgE
C4070232|T201|COMP|79396-8|LNC|NADH:ubiquinone reductase|NADH:ubiquinone reductase
C4070233|T201|COMP|79395-0|LNC|NADH:ubiquinone reductase|NADH:ubiquinone reductase
C4070234|T201|COMP|79394-3|LNC|Hepatocyte growth factor|Hepatocyte growth factor
C4070235|T201|COMP|79393-5|LNC|Flavin mononucleotide|Flavin mononucleotide
C4070236|T201|COMP|79392-7|LNC|Catecholamine metabolites pattern|Catecholamine metabolites pattern
C4070237|T201|COMP|79391-9|LNC|Catecholamine metabolites panel|Catecholamine metabolites panel
C4070238|T201|COMP|79390-1|LNC|Gastrointestinal pathogens identified|Gastrointestinal pathogens identified
C4070239|T201|COMP|79389-3|LNC|Rotavirus A nsp5 gene|Rotavirus A nsp5 gene
C4070241|T201|COMP|79387-7|LNC|Escherichia coli Stx2 toxin stx2 gene|Escherichia coli Stx2 toxin stx2 gene
C4070242|T201|COMP|79386-9|LNC|Escherichia coli Stx1 toxin stx1 gene|Escherichia coli Stx1 toxin stx1 gene
C4070243|T201|COMP|79385-1|LNC|Yersinia enterocolitica recN gene|Yersinia enterocolitica recN gene
C4070245|T201|COMP|79379-4|LNC|HIV 1 RNA+proviral DNA|HIV 1 RNA+proviral DNA
C4070246|T201|COMP|79377-8|LNC|Naltrexol|Naltrexol
C4070247|T201|COMP|79376-0|LNC|Microscopic observation^3rd specimen|Microscopic observation^3rd specimen
C4070248|T201|COMP|79375-2|LNC|Microscopic observation^2nd specimen|Microscopic observation^2nd specimen
C4070262|T201|COMP|79342-2|LNC|Carnitine biosynthesis intermediates pattern|Carnitine biosynthesis intermediates pattern
C4070263|T201|COMP|79341-4|LNC|Carnitine biosynthesis intermediates pattern|Carnitine biosynthesis intermediates pattern
C4070264|T201|COMP|79340-6|LNC|Carnitine biosynthesis intermediates pattern|Carnitine biosynthesis intermediates pattern
C4070265|T201|COMP|79339-8|LNC|Carnitine biosynthesis intermediates pattern|Carnitine biosynthesis intermediates pattern
C4070266|T201|COMP|79338-0|LNC|Hypoglycemics.oral|Hypoglycemics.oral
C4070267|T201|COMP|79337-2|LNC|Hypoglycemics.oral|Hypoglycemics.oral
C4070268|T201|COMP|79336-4|LNC|Hypoglycemics.oral|Hypoglycemics.oral
C4070269|T201|COMP|79335-6|LNC|Hypoglycemics.oral|Hypoglycemics.oral
C4070270|T201|COMP|79334-9|LNC|Hypoglycemics.oral|Hypoglycemics.oral
C4070271|T201|COMP|79333-1|LNC|Viscosity|Viscosity
C4070272|T201|COMP|79332-3|LNC|L-2-hydroxyglutarate|L-2-hydroxyglutarate
C4070273|T201|COMP|79331-5|LNC|Trimethyllysine/Creatinine|Trimethyllysine/Creatinine
C4070274|T201|COMP|79330-7|LNC|Trimethyllysine|Trimethyllysine
C4070275|T201|COMP|79329-9|LNC|Trimethyllysine|Trimethyllysine
C4070276|T201|COMP|79328-1|LNC|Trimethyllysine|Trimethyllysine
C4070277|T201|COMP|79327-3|LNC|Sterols pattern|Sterols pattern
C4070278|T201|COMP|79326-5|LNC|Squalene|Squalene
C4070281|T201|COMP|79323-2|LNC|7-Isobiopterin/Creatinine|7-Isobiopterin/Creatinine
C4070282|T201|COMP|79322-4|LNC|Lysophosphatidylcholine(26:0)|Lysophosphatidylcholine(26:0)
C4070283|T201|COMP|79321-6|LNC|Lysophosphatidylcholine(26:0)|Lysophosphatidylcholine(26:0)
C4070284|T201|COMP|79320-8|LNC|Lysophosphatidylcholine(26:0)|Lysophosphatidylcholine(26:0)
C4070285|T201|COMP|79319-0|LNC|L-2-hydroxyglutarate|L-2-hydroxyglutarate
C4070286|T201|COMP|79318-2|LNC|L-2-hydroxyglutarate|L-2-hydroxyglutarate
C4070287|T201|COMP|79317-4|LNC|L-2-hydroxyglutarate|L-2-hydroxyglutarate
C4070288|T201|COMP|79316-6|LNC|Isoxanthopterin|Isoxanthopterin
C4070289|T201|COMP|79315-8|LNC|Gamma butyrobetaine/Trimethyllysine|Gamma butyrobetaine/Trimethyllysine
C4070290|T201|COMP|79314-1|LNC|Gamma butyrobetaine/Trimethyllysine|Gamma butyrobetaine/Trimethyllysine
C4070291|T201|COMP|79313-3|LNC|Gamma butyrobetaine/Trimethyllysine|Gamma butyrobetaine/Trimethyllysine
C4070292|T201|COMP|79312-5|LNC|Gamma butyrobetaine/Trimethyllysine|Gamma butyrobetaine/Trimethyllysine
C4070293|T201|COMP|79311-7|LNC|Gamma butyrobetaine/Creatinine|Gamma butyrobetaine/Creatinine
C4070294|T201|COMP|79310-9|LNC|Gamma butyrobetaine|Gamma butyrobetaine
C4070295|T201|COMP|79309-1|LNC|Gamma butyrobetaine|Gamma butyrobetaine
C4070296|T201|COMP|79308-3|LNC|Gamma butyrobetaine|Gamma butyrobetaine
C4070297|T201|COMP|79307-5|LNC|D-2-hydroxyglutarate|D-2-hydroxyglutarate
C4070298|T201|COMP|79306-7|LNC|D-2-hydroxyglutarate|D-2-hydroxyglutarate
C4070299|T201|COMP|79305-9|LNC|D-2-hydroxyglutarate|D-2-hydroxyglutarate
C4070300|T201|COMP|79304-2|LNC|D-2-hydroxyglutarate|D-2-hydroxyglutarate
C4070301|T201|COMP|79303-4|LNC|D- & L-2-hydroxyglutarate pattern|D- & L-2-hydroxyglutarate pattern
C4070302|T201|COMP|79302-6|LNC|D- & L-2-hydroxyglutarate pattern|D- & L-2-hydroxyglutarate pattern
C4070303|T201|COMP|79301-8|LNC|D- & L-2-hydroxyglutarate pattern|D- & L-2-hydroxyglutarate pattern
C4070304|T201|COMP|79300-0|LNC|D- & L-2-hydroxyglutarate pattern|D- & L-2-hydroxyglutarate pattern
C4070305|T201|COMP|79298-6|LNC|D- & L-2-hydroxyglutarate panel|D- & L-2-hydroxyglutarate panel
C4070306|T201|COMP|79297-8|LNC|D- & L-2-hydroxyglutarate panel|D- & L-2-hydroxyglutarate panel
C4070307|T201|COMP|79296-0|LNC|D- & L-2-hydroxyglutarate panel|D- & L-2-hydroxyglutarate panel
C4070308|T201|COMP|79295-2|LNC|D- & L-2-hydroxyglutarate panel|D- & L-2-hydroxyglutarate panel
C4070309|T201|COMP|79294-5|LNC|D- & L-2-hydroxyglutarate panel|D- & L-2-hydroxyglutarate panel
C4070310|T201|COMP|79293-7|LNC|Creatine & guanidinoacetate pattern|Creatine & guanidinoacetate pattern
C4070311|T201|COMP|79292-9|LNC|Creatine, guanidinoacetate & creatinine pattern|Creatine, guanidinoacetate & creatinine pattern
C4070312|T201|COMP|79291-1|LNC|Creatine & guanidinoacetate pattern|Creatine & guanidinoacetate pattern
C4070313|T201|COMP|79290-3|LNC|Creatine, guanidinoacetate & creatinine panel|Creatine, guanidinoacetate & creatinine panel
C4070314|T201|COMP|79289-5|LNC|Creatine & guanidinoacetate panel|Creatine & guanidinoacetate panel
C4070315|T201|COMP|79288-7|LNC|Creatine & guanidinoacetate panel|Creatine & guanidinoacetate panel
C4070316|T201|COMP|79287-9|LNC|Carnitine biosynthesis intermediates panel|Carnitine biosynthesis intermediates panel
C4070317|T201|COMP|79286-1|LNC|Carnitine biosynthesis intermediates panel|Carnitine biosynthesis intermediates panel
C4070318|T201|COMP|79285-3|LNC|Carnitine biosynthesis intermediates panel|Carnitine biosynthesis intermediates panel
C4070319|T201|COMP|79283-8|LNC|C29 dicarboxylate|C29 dicarboxylate
C4070320|T201|COMP|79282-0|LNC|Biopterin/Biopterin+Neopterin|Biopterin/Biopterin+Neopterin
C4070321|T201|COMP|79281-2|LNC|Arabinose/Creatinine|Arabinose/Creatinine
C4070322|T201|COMP|79280-4|LNC|Alpha-aminoadipic semialdehyde|Alpha-aminoadipic semialdehyde
C4070323|T201|COMP|79279-6|LNC|Alpha-aminoadipic semialdehyde|Alpha-aminoadipic semialdehyde
C4070324|T201|COMP|79278-8|LNC|8-lathosterol|8-lathosterol
C4070325|T201|COMP|79277-0|LNC|7-lathosterol|7-lathosterol
C4070326|T201|COMP|79276-2|LNC|7,8-Dihydrobiopterin|7,8-Dihydrobiopterin
C4070327|T201|COMP|79275-4|LNC|3-Hydroxytrimethyl-L-lysine/Trimethyllysine|3-Hydroxytrimethyl-L-lysine/Trimethyllysine
C4070328|T201|COMP|79274-7|LNC|3-Hydroxytrimethyl-L-lysine/Trimethyllysine|3-Hydroxytrimethyl-L-lysine/Trimethyllysine
C4070329|T201|COMP|79273-9|LNC|3-Hydroxytrimethyl-L-lysine/Trimethyllysine|3-Hydroxytrimethyl-L-lysine/Trimethyllysine
C4070330|T201|COMP|79272-1|LNC|3-Hydroxytrimethyl-L-lysine/Trimethyllysine|3-Hydroxytrimethyl-L-lysine/Trimethyllysine
C4070331|T201|COMP|79271-3|LNC|3-Hydroxytrimethyl-L-lysine/Creatinine|3-Hydroxytrimethyl-L-lysine/Creatinine
C4070332|T201|COMP|79270-5|LNC|3-Hydroxytrimethyl-L-lysine|3-Hydroxytrimethyl-L-lysine
C4070333|T201|COMP|79269-7|LNC|3-Hydroxytrimethyl-L-lysine|3-Hydroxytrimethyl-L-lysine
C4070334|T201|COMP|79268-9|LNC|3-Hydroxytrimethyl-L-lysine|3-Hydroxytrimethyl-L-lysine
C4070335|T201|COMP|79266-3|LNC|Lead|Lead
C4070336|T201|COMP|79262-2|LNC|Methamphetamine cutoff|Methamphetamine cutoff
C4070337|T201|COMP|79261-4|LNC|HYDROcodone cutoff|HYDROcodone cutoff
C4070338|T201|COMP|79260-6|LNC|fentaNYL cutoff|fentaNYL cutoff
C4070339|T201|COMP|79259-8|LNC|fentaNYL cutoff|fentaNYL cutoff
C4070340|T201|COMP|79258-0|LNC|Meprobamate cutoff|Meprobamate cutoff
C4070341|T201|COMP|79252-3|LNC|Nordiazepam cutoff|Nordiazepam cutoff
C4070342|T201|COMP|79251-5|LNC|diazePAM cutoff|diazePAM cutoff
C4070344|T201|COMP|79249-9|LNC|Methadone cutoff|Methadone cutoff
C4070345|T201|COMP|79248-1|LNC|Methylenedioxyethylamphetamine cutoff|Methylenedioxyethylamphetamine cutoff
C4070346|T201|COMP|79247-3|LNC|Methylenedioxymethamphetamine cutoff|Methylenedioxymethamphetamine cutoff
C4070347|T201|COMP|79246-5|LNC|Methedrone|Methedrone
C4070348|T201|COMP|79245-7|LNC|Triazolam cutoff|Triazolam cutoff
C4070349|T201|COMP|79244-0|LNC|Ethylone cutoff|Ethylone cutoff
C4070350|T201|COMP|79243-2|LNC|Ethylone|Ethylone
C4070351|T201|COMP|79242-4|LNC|Methylone cutoff|Methylone cutoff
C4070352|T201|COMP|79241-6|LNC|Methedrone cutoff|Methedrone cutoff
C4070353|T201|COMP|79240-8|LNC|Tapentadol cutoff|Tapentadol cutoff
C4070354|T201|COMP|79239-0|LNC|Ethyl glucuronide cutoff|Ethyl glucuronide cutoff
C4070355|T201|COMP|79238-2|LNC|Methylenedioxypyrovalerone cutoff|Methylenedioxypyrovalerone cutoff
C4070356|T201|COMP|79237-4|LNC|Mephedrone cutoff|Mephedrone cutoff
C4070357|T201|COMP|79236-6|LNC|Methcathinone cutoff|Methcathinone cutoff
C4070358|T201|COMP|79235-8|LNC|Butylone cutoff|Butylone cutoff
C4070359|T201|COMP|79234-1|LNC|Butylone|Butylone
C4070360|T201|COMP|79233-3|LNC|Naphyrone cutoff|Naphyrone cutoff
C4070361|T201|COMP|79232-5|LNC|Naphyrone|Naphyrone
C4070362|T201|COMP|79231-7|LNC|Amoxapine|Amoxapine
C4070363|T201|COMP|79230-9|LNC|Amiodarone|Amiodarone
C4070364|T201|COMP|79229-1|LNC|Amitriptyline|Amitriptyline
C4070365|T201|COMP|79223-4|LNC|Atenolol|Atenolol
C4070366|T201|COMP|79222-6|LNC|Benzodiazepines|Benzodiazepines
C4070367|T201|COMP|79221-8|LNC|Steroid fractions panel|Steroid fractions panel
C4070368|T201|COMP|79220-0|LNC|Steroid fractions interpretation|Steroid fractions interpretation
C4070375|T201|COMP|79212-7|LNC|Fetal microdeletions risk|Fetal microdeletions risk
C4070376|T201|COMP|79211-9|LNC|Fetal chromosome X & Y aneuploidy risk|Fetal chromosome X & Y aneuploidy risk
C4070377|T201|COMP|79210-1|LNC|FLT3 gene internal tandem duplication|FLT3 gene internal tandem duplication
C4070378|T201|COMP|79209-3|LNC|t(2;3)(q13;p25)(PAX8,PPARG) fusion transcript|t(2;3)(q13;p25)(PAX8,PPARG) fusion transcript
C4070381|T201|COMP|79206-9|LNC|inv(2)(p21;p23)(EML4,ALK) fusion transcript|inv(2)(p21;p23)(EML4,ALK) fusion transcript
C4070382|T201|COMP|79205-1|LNC|Somatotropin^1.5H post dose arginine+insulin|Somatotropin^1.5H post dose arginine+insulin
C4070383|T201|COMP|79204-4|LNC|Somatotropin^1.25H post dose arginine+insulin|Somatotropin^1.25H post dose arginine+insulin
C4070384|T201|COMP|79203-6|LNC|Somatotropin^1H post dose arginine+insulin|Somatotropin^1H post dose arginine+insulin
C4070385|T201|COMP|79202-8|LNC|Somatotropin^45M post dose arginine+insulin|Somatotropin^45M post dose arginine+insulin
C4070386|T201|COMP|79201-0|LNC|Somatotropin^30M post dose arginine+insulin|Somatotropin^30M post dose arginine+insulin
C4070387|T201|COMP|79200-2|LNC|Somatotropin^2.5H post dose arginine+insulin|Somatotropin^2.5H post dose arginine+insulin
C4070388|T201|COMP|79199-6|LNC|Somatotropin^15M post dose arginine+insulin|Somatotropin^15M post dose arginine+insulin
C4070389|T201|COMP|79198-8|LNC|Somatotropin^2.25H post dose arginine+insulin|Somatotropin^2.25H post dose arginine+insulin
C4070390|T201|COMP|79197-0|LNC|Somatotropin^2H post dose arginine+insulin|Somatotropin^2H post dose arginine+insulin
C4070391|T201|COMP|79196-2|LNC|Glucose^1H post dose arginine+insulin|Glucose^1H post dose arginine+insulin
C4070392|T201|COMP|79195-4|LNC|Glucose^45M post dose arginine+insulin|Glucose^45M post dose arginine+insulin
C4070393|T201|COMP|79194-7|LNC|Glucose^30M post dose arginine+insulin|Glucose^30M post dose arginine+insulin
C4070394|T201|COMP|79193-9|LNC|Glucose^15M post dose arginine+insulin|Glucose^15M post dose arginine+insulin
C4070396|T201|COMP|79190-5|LNC|Zika virus RNA|Zika virus RNA
C4070397|T201|COMP|79189-7|LNC|Hepatitis C virus core Ag|Hepatitis C virus core Ag
C4070399|T201|COMP|79187-1|LNC|Cells.CD3+CD4+CD8+|Cells.CD3+CD4+CD8+
C4070400|T201|COMP|79186-3|LNC|Cells.CD3+CD4+CD8+/100 cells|Cells.CD3+CD4+CD8+/100 cells
C4070401|T201|COMP|79184-8|LNC|Last name|Last name
C4070402|T201|COMP|79178-0|LNC|4-Hydroxycyclohexylacetate/creatinine|4-Hydroxycyclohexylacetate/creatinine
C4070404|T201|COMP|79176-4|LNC|Somatotropin^30M post XXX challenge|Somatotropin^30M post XXX challenge
C4070405|T201|COMP|79175-6|LNC|Somatotropin^1H post XXX challenge|Somatotropin^1H post XXX challenge
C4070406|T201|COMP|79174-9|LNC|Somatotropin^1.5H post XXX challenge|Somatotropin^1.5H post XXX challenge
C4070407|T201|COMP|79173-1|LNC|Somatotropin^2H post XXX challenge|Somatotropin^2H post XXX challenge
C4070408|T201|COMP|79172-3|LNC|Somatotropin^2.5H post XXX challenge|Somatotropin^2.5H post XXX challenge
C4070409|T201|COMP|79171-5|LNC|Malus domestica recombinant (rMal d) 4 Ab.IgE|Malus domestica recombinant (rMal d) 4 Ab.IgE
C4070410|T201|COMP|79170-7|LNC|Prunus avium recombinant (rPru av) 1 Ab.IgE|Prunus avium recombinant (rPru av) 1 Ab.IgE
C4070411|T201|COMP|79169-9|LNC|Prunus avium recombinant (rPru av) 3 Ab.IgE|Prunus avium recombinant (rPru av) 3 Ab.IgE
C4070412|T201|COMP|79168-1|LNC|Prunus avium recombinant (rPru av) 4 Ab.IgE|Prunus avium recombinant (rPru av) 4 Ab.IgE
C4070413|T201|COMP|79167-3|LNC|Apis mellifera recombinant (rApi m) 2 Ab.IgE|Apis mellifera recombinant (rApi m) 2 Ab.IgE
C4070414|T201|COMP|79166-5|LNC|Prunus persica native (nPru p) 3 Ab.IgE|Prunus persica native (nPru p) 3 Ab.IgE
C4070416|T201|COMP|79164-0|LNC|CES1 gene.c.428G>A|CES1 gene.c.428G>A
C4070417|T201|COMP|79163-2|LNC|Z-10-Hydroxynortriptyline|Z-10-Hydroxynortriptyline
C4070418|T201|COMP|79154-1|LNC|Alizapride|Alizapride
C4070419|T201|COMP|79153-3|LNC|Alfentanil|Alfentanil
C4070420|T201|COMP|79152-5|LNC|Acenocoumarol|Acenocoumarol
C4070422|T201|COMP|79149-1|LNC|Trimeprazine|Trimeprazine
C4070423|T201|COMP|79148-3|LNC|traMADol|traMADol
C4070424|T201|COMP|79147-5|LNC|traMADol|traMADol
C4070425|T201|COMP|79146-7|LNC|Tapentadol|Tapentadol
C4070426|T201|COMP|79145-9|LNC|Tapentadol|Tapentadol
C4070427|T201|COMP|79135-0|LNC|Acebutolol|Acebutolol
C4070428|T201|COMP|79134-3|LNC|Abacavir|Abacavir
C4070429|T201|COMP|79133-5|LNC|9-Hydroxyrisperidone|9-Hydroxyrisperidone
C4070430|T201|COMP|79132-7|LNC|4-Hydroxymidazolam|4-Hydroxymidazolam
C4070431|T201|COMP|79131-9|LNC|1-Hydroxymidazolam|1-Hydroxymidazolam
C4070432|T201|COMP|79130-1|LNC|Platelet aggregation.ristocetin induced^500 ug/mL|Platelet aggregation.ristocetin induced^500 ug/mL
C4070433|T201|COMP|79129-3|LNC|Uroporphyrin 3 isomer/Creatinine|Uroporphyrin 3 isomer/Creatinine
C4070434|T201|COMP|79128-5|LNC|Uroporphyrin 3 isomer|Uroporphyrin 3 isomer
C4070435|T201|COMP|79127-7|LNC|Uroporphyrin 1 isomer/Creatinine|Uroporphyrin 1 isomer/Creatinine
C4070436|T201|COMP|79126-9|LNC|Uroporphyrin 1 isomer|Uroporphyrin 1 isomer
C4070437|T201|COMP|79125-1|LNC|Hawkinsin|Hawkinsin
C4070454|T201|COMP|79102-0|LNC|Heart transplant acute cellular rejection risk|Heart transplant acute cellular rejection risk
C4070555|T201|COMP|78995-8|LNC|Prolactin.monomeric/Prolactin|Prolactin.monomeric/Prolactin
C4070556|T201|COMP|78994-1|LNC|Prolactin.monomeric|Prolactin.monomeric
C4070557|T201|COMP|78993-3|LNC|Prolactin isoforms panel|Prolactin isoforms panel
C4070558|T201|COMP|78992-5|LNC|Melatonin|Melatonin
C4070559|T201|COMP|78990-9|LNC|Flavin adenine dinucleotide|Flavin adenine dinucleotide
C4070560|T201|COMP|78989-1|LNC|Cryoglobulin|Cryoglobulin
C4070561|T201|COMP|78988-3|LNC|Cortisol|Cortisol
C4070562|T201|COMP|78987-5|LNC|Provasopressin.C-terminal|Provasopressin.C-terminal
C4070563|T201|COMP|78986-7|LNC|Prolactin.dimeric/Prolactin|Prolactin.dimeric/Prolactin
C4070564|T201|COMP|78985-9|LNC|Prolactin.dimeric|Prolactin.dimeric
C4070565|T201|COMP|78984-2|LNC|Macroprolactin/Prolactin|Macroprolactin/Prolactin
C4070566|T201|COMP|78983-4|LNC|4-Hydroxy-3-Methoxyphenyllactate|4-Hydroxy-3-Methoxyphenyllactate
C4070573|T201|COMP|78972-7|LNC|CYP2C8 gene targeted mutation analysis|CYP2C8 gene targeted mutation analysis
C4070574|T201|COMP|78971-9|LNC|Phosphomannomutase 1|Phosphomannomutase 1
C4070575|T201|COMP|78970-1|LNC|Phosphomannomutase 1|Phosphomannomutase 1
C4070576|T201|COMP|78969-3|LNC|Neurofilament heavy chain Ab|Neurofilament heavy chain Ab
C4070577|T201|COMP|78968-5|LNC|Benperidol|Benperidol
C4070578|T201|COMP|78967-7|LNC|Sedoheptulose/Creatinine|Sedoheptulose/Creatinine
C4070579|T201|COMP|78966-9|LNC|S-adenosylmethionine|S-adenosylmethionine
C4070580|T201|COMP|78965-1|LNC|Neurofilament medium chain Ab|Neurofilament medium chain Ab
C4070581|T201|COMP|78964-4|LNC|N-acetylaspartylglutamate|N-acetylaspartylglutamate
C4070582|T201|COMP|78962-8|LNC|IgG clearance/Transferrin clearance|IgG clearance/Transferrin clearance
C4070583|T201|COMP|78961-0|LNC|IgG clearance/Albumin clearance|IgG clearance/Albumin clearance
C4070584|T201|COMP|78960-2|LNC|Aldosterone & renin concentration panel|Aldosterone & renin concentration panel
C4070585|T201|COMP|78959-4|LNC|Hyocholate|Hyocholate
C4070586|T201|COMP|78958-6|LNC|Cathepsin A|Cathepsin A
C4070603|T201|COMP|78922-2|LNC|Respiratory pathogens DNA & RNA panel|Respiratory pathogens DNA & RNA panel
C4070605|T201|COMP|78920-6|LNC|cycloSPORINE|cycloSPORINE
C4070622|T201|COMP|78894-3|LNC|Liver fibrosis score|Liver fibrosis score
C4070623|T201|COMP|78893-5|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C4070624|T201|COMP|78892-7|LNC|Silver|Silver
C4070625|T201|COMP|78891-9|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C4070626|T201|COMP|78890-1|LNC|Barium|Barium
C4070627|T201|COMP|78889-3|LNC|Tricyclic antidepressants|Tricyclic antidepressants
C4070628|T201|COMP|78888-5|LNC|Trimeprazine|Trimeprazine
C4070629|T201|COMP|78886-9|LNC|Venlafaxine cutoff|Venlafaxine cutoff
C4070630|T201|COMP|78885-1|LNC|traZODone cutoff|traZODone cutoff
C4070631|T201|COMP|78884-4|LNC|Lurasidone|Lurasidone
C4070632|T201|COMP|78883-6|LNC|Triazolam|Triazolam
C4070633|T201|COMP|78882-8|LNC|Sertraline cutoff|Sertraline cutoff
C4070634|T201|COMP|78881-0|LNC|RCS-4 5-hydroxypentyl cutoff|RCS-4 5-hydroxypentyl cutoff
C4070635|T201|COMP|78880-2|LNC|RCS-4 5-hydroxypentyl|RCS-4 5-hydroxypentyl
C4070636|T201|COMP|78879-4|LNC|RCS-4 5-carboxypentyl cutoff|RCS-4 5-carboxypentyl cutoff
C4070637|T201|COMP|78878-6|LNC|RCS-4 5-carboxypentyl|RCS-4 5-carboxypentyl
C4070638|T201|COMP|78877-8|LNC|QUEtiapine|QUEtiapine
C4070639|T201|COMP|78876-0|LNC|Pheniramine|Pheniramine
C4070640|T201|COMP|78875-2|LNC|PARoxetine cutoff|PARoxetine cutoff
C4070641|T201|COMP|78874-5|LNC|oxyMORphone|oxyMORphone
C4070642|T201|COMP|78873-7|LNC|oxyCODONE|oxyCODONE
C4070643|T201|COMP|78872-9|LNC|OPC3373|OPC3373
C4070644|T201|COMP|78871-1|LNC|OPC3373 cutoff|OPC3373 cutoff
C4070645|T201|COMP|78870-3|LNC|OPC3373|OPC3373
C4070646|T201|COMP|78869-5|LNC|Norvenlafaxine cutoff|Norvenlafaxine cutoff
C4070647|T201|COMP|78868-7|LNC|Norhydrocodone cutoff|Norhydrocodone cutoff
C4070648|T201|COMP|78867-9|LNC|Norfentanyl cutoff|Norfentanyl cutoff
C4070649|T201|COMP|78866-1|LNC|Norbuprenorphine cutoff|Norbuprenorphine cutoff
C4070650|T201|COMP|78865-3|LNC|Naltrexol cutoff|Naltrexol cutoff
C4070651|T201|COMP|78864-6|LNC|Naloxone cutoff|Naloxone cutoff
C4070652|T201|COMP|78863-8|LNC|Naloxol cutoff|Naloxol cutoff
C4070653|T201|COMP|78862-0|LNC|Naloxol|Naloxol
C4070654|T201|COMP|78861-2|LNC|Morphine|Morphine
C4070655|T201|COMP|78860-4|LNC|Mirtazapine cutoff|Mirtazapine cutoff
C4070656|T201|COMP|78859-6|LNC|Mirtazapine|Mirtazapine
C4070657|T201|COMP|78858-8|LNC|Methcathinone|Methcathinone
C4070658|T201|COMP|78857-0|LNC|Methadone|Methadone
C4070659|T201|COMP|78856-2|LNC|Meprobamate|Meprobamate
C4070660|T201|COMP|78855-4|LNC|M-chlorophenylpiperazine|M-chlorophenylpiperazine
C4070661|T201|COMP|78854-7|LNC|M-chlorophenylpiperazine|M-chlorophenylpiperazine
C4070662|T201|COMP|78853-9|LNC|M-chlorophenylpiperazine|M-chlorophenylpiperazine
C4070663|T201|COMP|78852-1|LNC|M-chlorophenylpiperazine|M-chlorophenylpiperazine
C4070664|T201|COMP|78851-3|LNC|M-chlorophenylpiperazine|M-chlorophenylpiperazine
C4070665|T201|COMP|78850-5|LNC|JWH-250 5-hydroxypentyl cutoff|JWH-250 5-hydroxypentyl cutoff
C4070666|T201|COMP|78849-7|LNC|JWH-210 5-hydroxypentyl cutoff|JWH-210 5-hydroxypentyl cutoff
C4070667|T201|COMP|78848-9|LNC|JWH-210 5-Hydroxypentyl|JWH-210 5-Hydroxypentyl
C4070668|T201|COMP|78847-1|LNC|JWH-210 5-carboxypentyl cutoff|JWH-210 5-carboxypentyl cutoff
C4070669|T201|COMP|78846-3|LNC|JWH-200 6-Hydroxyindole cutoff|JWH-200 6-Hydroxyindole cutoff
C4070670|T201|COMP|78845-5|LNC|JWH-200 6-Hydroxyindole|JWH-200 6-Hydroxyindole
C4070671|T201|COMP|78844-8|LNC|JWH-200 4-Hydroxyindole cutoff|JWH-200 4-Hydroxyindole cutoff
C4070672|T201|COMP|78843-0|LNC|JWH-200 4-Hydroxyindole|JWH-200 4-Hydroxyindole
C4070685|T201|COMP|79649-0|LNC|Homocysteine cysteine disulfide/Creatinine|Homocysteine cysteine disulfide/Creatinine
C4070686|T201|COMP|79647-4|LNC|Beta-ureidoisobutyrate/Creatinine|Beta-ureidoisobutyrate/Creatinine
C4070687|T201|COMP|79646-6|LNC|Delta aminolevulinate|Delta aminolevulinate
C4070688|T201|COMP|79645-8|LNC|L-serine/Creatinine|L-serine/Creatinine
C4070689|T201|COMP|79490-9|LNC|3,4-Dihydroxyhydrocinnamate/Creatinine|3,4-Dihydroxyhydrocinnamate/Creatinine
C4070690|T201|COMP|79489-1|LNC|Salicylurate|Salicylurate
C4070691|T201|COMP|79488-3|LNC|3,4-Dihydroxybutyrate|3,4-Dihydroxybutyrate
C4070692|T201|COMP|79487-5|LNC|Lactyl lactate/Creatinine|Lactyl lactate/Creatinine
C4070693|T201|COMP|79486-7|LNC|3,5-Dihydroxybenzoate/Creatinine|3,5-Dihydroxybenzoate/Creatinine
C4070694|T201|COMP|79485-9|LNC|4-Hydroxyvalerate/Creatinine|4-Hydroxyvalerate/Creatinine
C4070695|T201|COMP|79257-2|LNC|Methylenedioxyamphetamine cutoff|Methylenedioxyamphetamine cutoff
C4070696|T201|COMP|79256-4|LNC|Carisoprodol+Meprobamate cutoff|Carisoprodol+Meprobamate cutoff
C4070697|T201|COMP|79255-6|LNC|oxyCODONE cutoff|oxyCODONE cutoff
C4070698|T201|COMP|79254-9|LNC|LORazepam cutoff|LORazepam cutoff
C4070699|T201|COMP|79253-1|LNC|Oxazepam cutoff|Oxazepam cutoff
C4070711|T201|COMP|79228-3|LNC|amLODIPine|amLODIPine
C4070712|T201|COMP|79227-5|LNC|Amobarbital|Amobarbital
C4070713|T201|COMP|79226-7|LNC|ARIPiprazole|ARIPiprazole
C4070714|T201|COMP|79225-9|LNC|Barbital|Barbital
C4070715|T201|COMP|79224-2|LNC|Baclofen|Baclofen
C4070716|T201|COMP|79183-0|LNC|First name|First name
C4070717|T201|COMP|79182-2|LNC|RNA polymerase III Ab.IgG|RNA polymerase III Ab.IgG
C4070718|T201|COMP|79181-4|LNC|Somatotropin^15M post XXX challenge|Somatotropin^15M post XXX challenge
C4070719|T201|COMP|79180-6|LNC|Somatotropin^45M post XXX challenge|Somatotropin^45M post XXX challenge
C4070720|T201|COMP|79179-8|LNC|Somatotropin^75M post XXX challenge|Somatotropin^75M post XXX challenge
C4070721|T201|COMP|78982-6|LNC|D-3-phosphoglycerate dehydrogenase|D-3-phosphoglycerate dehydrogenase
C4070723|T201|COMP|78918-0|LNC|7-Hydroxyquetiapine|7-Hydroxyquetiapine
C4070724|T201|COMP|78917-2|LNC|Cells.FGFR1 gene rearrangements/Cells counted|Cells.FGFR1 gene rearrangements/Cells counted
C4070725|T201|COMP|78916-4|LNC|FGFR1 gene rearrangements|FGFR1 gene rearrangements
C4070726|T201|COMP|78915-6|LNC|FGFR1 gene rearrangements|FGFR1 gene rearrangements
C4070731|T201|COMP|78842-2|LNC|JWH-122 5-hydroxypentyl cutoff|JWH-122 5-hydroxypentyl cutoff
C4070732|T201|COMP|78841-4|LNC|JWH-122 5-hydroxypentyl|JWH-122 5-hydroxypentyl
C4070733|T201|COMP|78840-6|LNC|JWH-081 5-hydroxypentyl cutoff|JWH-081 5-hydroxypentyl cutoff
C4070734|T201|COMP|78839-8|LNC|JWH-073 butanoate cutoff|JWH-073 butanoate cutoff
C4070735|T201|COMP|78838-0|LNC|JWH-073 4-hydroxybutyl cutoff|JWH-073 4-hydroxybutyl cutoff
C4070736|T201|COMP|78837-2|LNC|JWH-018 pentanoate cutoff|JWH-018 pentanoate cutoff
C4070737|T201|COMP|78836-4|LNC|JWH-018 5-hydroxypentyl cutoff|JWH-018 5-hydroxypentyl cutoff
C4070738|T201|COMP|78835-6|LNC|Imipramine cutoff|Imipramine cutoff
C4070739|T201|COMP|78834-9|LNC|Hydroxylurasidone cutoff|Hydroxylurasidone cutoff
C4070740|T201|COMP|78833-1|LNC|Hydroxylurasidone|Hydroxylurasidone
C4070741|T201|COMP|78832-3|LNC|Hydroxybupropion cutoff|Hydroxybupropion cutoff
C4070742|T201|COMP|78831-5|LNC|Hydroxybupropion|Hydroxybupropion
C4070743|T201|COMP|78830-7|LNC|HYDROcodone|HYDROcodone
C4070744|T201|COMP|78829-9|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C4070745|T201|COMP|78828-1|LNC|fentaNYL|fentaNYL
C4070746|T201|COMP|78827-3|LNC|fentaNYL cutoff|fentaNYL cutoff
C4070747|T201|COMP|78826-5|LNC|Ethyl acetate|Ethyl acetate
C4070748|T201|COMP|78825-7|LNC|Ecgonine methyl ester|Ecgonine methyl ester
C4070749|T201|COMP|78824-0|LNC|DULoxetine cutoff|DULoxetine cutoff
C4070750|T201|COMP|78823-2|LNC|DULoxetine|DULoxetine
C4070751|T201|COMP|78822-4|LNC|Doxepin cutoff|Doxepin cutoff
C4070752|T201|COMP|78821-6|LNC|Desipramine cutoff|Desipramine cutoff
C4070753|T201|COMP|78820-8|LNC|Cyclobenzaprine cutoff|Cyclobenzaprine cutoff
C4070754|T201|COMP|78819-0|LNC|clomiPRAMINE cutoff|clomiPRAMINE cutoff
C4070755|T201|COMP|78818-2|LNC|Citalopram cutoff|Citalopram cutoff
C4070756|T201|COMP|78817-4|LNC|Cathinone|Cathinone
C4070757|T201|COMP|78816-6|LNC|Carisoprodol+Meprobamate|Carisoprodol+Meprobamate
C4070758|T201|COMP|78815-8|LNC|Carisoprodol|Carisoprodol
C4070769|T201|COMP|79382-8|LNC|Campylobacter coli+jejuni+lari fusA gene|Campylobacter coli+jejuni+lari fusA gene
C4070770|T201|COMP|79381-0|LNC|Gastrointestinal pathogens panel|Gastrointestinal pathogens panel
C4070771|T201|COMP|79380-2|LNC|HIV 1 RNA+proviral DNA|HIV 1 RNA+proviral DNA
C4070772|T201|COMP|79144-2|LNC|Methcathinone|Methcathinone
C4070773|T201|COMP|79143-4|LNC|Mercury|Mercury
C4070774|T201|COMP|79142-6|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C4070775|T201|COMP|79141-8|LNC|Cathinone|Cathinone
C4070776|T201|COMP|79140-0|LNC|Carisoprodol+Meprobamate|Carisoprodol+Meprobamate
C4070777|T201|COMP|79139-2|LNC|Buprenorphine|Buprenorphine
C4070778|T201|COMP|79138-4|LNC|Buprenorphine|Buprenorphine
C4070779|T201|COMP|79137-6|LNC|Benzylpiperazine|Benzylpiperazine
C4070780|T201|COMP|79136-8|LNC|Acepromazine|Acepromazine
C4070782|T201|COMP|78814-1|LNC|Cannabicyclohexanol cutoff|Cannabicyclohexanol cutoff
C4070783|T201|COMP|78813-3|LNC|Cannabicyclohexanol|Cannabicyclohexanol
C4070784|T201|COMP|78812-5|LNC|buPROPion cutoff|buPROPion cutoff
C4070785|T201|COMP|78811-7|LNC|Buprenorphine cutoff|Buprenorphine cutoff
C4070786|T201|COMP|78810-9|LNC|Beryllium|Beryllium
C4070787|T201|COMP|78809-1|LNC|Benzylpiperazine|Benzylpiperazine
C4070788|T201|COMP|78808-3|LNC|Benzodiazepines|Benzodiazepines
C4070789|T201|COMP|78807-5|LNC|Barium|Barium
C4070790|T201|COMP|78806-7|LNC|Alminoprofen|Alminoprofen
C4070791|T201|COMP|78805-9|LNC|Barium|Barium
C4070792|T201|COMP|78804-2|LNC|Barbital|Barbital
C4070793|T201|COMP|78803-4|LNC|Barbital|Barbital
C4070794|T201|COMP|78802-6|LNC|Baclofen|Baclofen
C4070795|T201|COMP|78801-8|LNC|Atropine|Atropine
C4070796|T201|COMP|78800-0|LNC|Atropine|Atropine
C4070797|T201|COMP|78799-4|LNC|Atenolol|Atenolol
C4070798|T201|COMP|78798-6|LNC|Atenolol|Atenolol
C4070799|T201|COMP|78797-8|LNC|Atazanavir^trough|Atazanavir^trough
C4070800|T201|COMP|78796-0|LNC|Atazanavir|Atazanavir
C4070801|T201|COMP|78795-2|LNC|Arsenic|Arsenic
C4070802|T201|COMP|78794-5|LNC|ARIPiprazole|ARIPiprazole
C4070803|T201|COMP|78793-7|LNC|ARIPiprazole|ARIPiprazole
C4070804|T201|COMP|78792-9|LNC|Anakinra|Anakinra
C4070805|T201|COMP|78790-3|LNC|Amphetamine|Amphetamine
C4070806|T201|COMP|78789-5|LNC|Amoxapine|Amoxapine
C4070807|T201|COMP|78788-7|LNC|amLODIPine|amLODIPine
C4070808|T201|COMP|78787-9|LNC|amLODIPine|amLODIPine
C4070809|T201|COMP|78786-1|LNC|Amitriptyline|Amitriptyline
C4070810|T201|COMP|78785-3|LNC|Amitriptyline|Amitriptyline
C4070811|T201|COMP|78784-6|LNC|Amiodarone|Amiodarone
C4070812|T201|COMP|78783-8|LNC|AM-2201 4-hydroxypentyl cutoff|AM-2201 4-hydroxypentyl cutoff
C4070813|T201|COMP|78782-0|LNC|Aluminum|Aluminum
C4070814|T201|COMP|78781-2|LNC|ALPRAZolam cutoff|ALPRAZolam cutoff
C4070815|T201|COMP|78779-6|LNC|Alizapride|Alizapride
C4070816|T201|COMP|78778-8|LNC|Alfentanil|Alfentanil
C4070817|T201|COMP|78777-0|LNC|Alfentanil|Alfentanil
C4070818|T201|COMP|78776-2|LNC|Acepromazine|Acepromazine
C4070819|T201|COMP|78775-4|LNC|Acenocoumarol|Acenocoumarol
C4070820|T201|COMP|78774-7|LNC|Acenocoumarol|Acenocoumarol
C4070821|T201|COMP|78773-9|LNC|Abacavir|Abacavir
C4070822|T201|COMP|78772-1|LNC|Abacavir|Abacavir
C4070823|T201|COMP|78771-3|LNC|9-Hydroxyrisperidone|9-Hydroxyrisperidone
C4070832|T201|COMP|78762-2|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C4070833|T201|COMP|78761-4|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C4070834|T201|COMP|78760-6|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C4070835|T201|COMP|78759-8|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C4070836|T201|COMP|78758-0|LNC|4-Hydroxymidazolam|4-Hydroxymidazolam
C4070837|T201|COMP|78757-2|LNC|2-Oxo-3-Hydroxy-Lysergate diethylamide|2-Oxo-3-Hydroxy-Lysergate diethylamide
C4070838|T201|COMP|78756-4|LNC|2-Oxo-3-Hydroxy-Lysergate diethylamide|2-Oxo-3-Hydroxy-Lysergate diethylamide
C4070839|T201|COMP|78755-6|LNC|1-Hydroxymidazolam|1-Hydroxymidazolam
C4070840|T201|COMP|78754-9|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C4070841|T201|COMP|78753-1|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C4070842|T201|COMP|78752-3|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C4070843|T201|COMP|78751-5|LNC|11-Hydroxy delta-9 tetrahydrocannabinol|11-Hydroxy delta-9 tetrahydrocannabinol
C4070844|T201|COMP|78750-7|LNC|Hepatitis E virus RNA|Hepatitis E virus RNA
C4070845|T201|COMP|78749-9|LNC|Glycolate|Glycolate
C4070846|T201|COMP|78748-1|LNC|Hemoglobin pattern|Hemoglobin pattern
C4070849|T201|COMP|78743-2|LNC|Steroid fractions interpretation|Steroid fractions interpretation
C4070850|T201|COMP|78742-4|LNC|Yeast|Yeast
C4070851|T201|COMP|78741-6|LNC|Pathologic casts|Pathologic casts
C4070852|T201|COMP|78740-8|LNC|Pathologic casts|Pathologic casts
C4070853|T201|COMP|78739-0|LNC|Platelet aggregation.ristocetin induced^low dose|Platelet aggregation.ristocetin induced^low dose
C4070887|T201|COMP|78702-8|LNC|Multiple drug resistant gram negative organism|Multiple drug resistant gram negative organism
C4070888|T201|COMP|78701-0|LNC|Ulmus crassifolia Ab.IgE|Ulmus crassifolia Ab.IgE
C4070890|T201|COMP|78699-6|LNC|Liver fibrosis score panel|Liver fibrosis score panel
C4070891|T201|COMP|78698-8|LNC|Liver fibrosis score panel|Liver fibrosis score panel
C4070892|T201|COMP|78697-0|LNC|Olea europaea Ab.IgG|Olea europaea Ab.IgG
C4070893|T201|COMP|78696-2|LNC|Selenium|Selenium
C4070894|T201|COMP|78695-4|LNC|Guanine/Creatinine|Guanine/Creatinine
C4070895|T201|COMP|78694-7|LNC|Dihydroorotate/Creatinine|Dihydroorotate/Creatinine
C4070896|T201|COMP|78693-9|LNC|Dihydrothymine/Creatinine|Dihydrothymine/Creatinine
C4070897|T201|COMP|78692-1|LNC|Pseudouridine/Creatinine|Pseudouridine/Creatinine
C4070898|T201|COMP|78691-3|LNC|Guanosine/Creatinine|Guanosine/Creatinine
C4070899|T201|COMP|78690-5|LNC|5-hydroxymethyluracil/Creatinine|5-hydroxymethyluracil/Creatinine
C4070900|T201|COMP|78689-7|LNC|Adenylosuccinate/Creatinine|Adenylosuccinate/Creatinine
C4070903|T201|COMP|78686-3|LNC|Platelet aggregation.ristocetin induced^high dose|Platelet aggregation.ristocetin induced^high dose
C4070904|T201|COMP|78685-5|LNC|Platelet aggregation.collagen induced|Platelet aggregation.collagen induced
C4070986|T201|COMP|78537-8|LNC|Urea nitrogen^4H dwell specimen|Urea nitrogen^4H dwell specimen
C4070987|T201|COMP|78536-0|LNC|Urea nitrogen^2H dwell specimen|Urea nitrogen^2H dwell specimen
C4070988|T201|COMP|78535-2|LNC|Glucose^4H dwell specimen|Glucose^4H dwell specimen
C4070989|T201|COMP|78534-5|LNC|Glucose^2H dwell specimen|Glucose^2H dwell specimen
C4070990|T201|COMP|78533-7|LNC|Creatinine^4H dwell specimen|Creatinine^4H dwell specimen
C4070991|T201|COMP|78532-9|LNC|Creatinine^2H dwell specimen|Creatinine^2H dwell specimen
C4070992|T201|COMP|78531-1|LNC|Vesicular stomatitis Indiana virus RNA|Vesicular stomatitis Indiana virus RNA
C4070993|T201|COMP|78530-3|LNC|Vesicular stomatitis New Jersey virus RNA|Vesicular stomatitis New Jersey virus RNA
C4070994|T201|COMP|78529-5|LNC|Adenovirus Ag|Adenovirus Ag
C4070996|T201|COMP|78527-9|LNC|Platelet aggregation.collagen induced^5 ug/mL|Platelet aggregation.collagen induced^5 ug/mL
C4070997|T201|COMP|78526-1|LNC|Platelet aggregation.collagen induced^1.25 ug/mL|Platelet aggregation.collagen induced^1.25 ug/mL
C4070999|T201|COMP|78524-6|LNC|Platelet aggregation.EPINEPHrine induced^6 umol/L|Platelet aggregation.EPINEPHrine induced^6 umol/L
C4071005|T201|COMP|78518-8|LNC|Cholesterol|Cholesterol
C4071006|T201|COMP|78517-0|LNC|Renin^2H post XXX challenge|Renin^2H post XXX challenge
C4071007|T201|COMP|78516-2|LNC|Lactose^45M post dose lactose PO|Lactose^45M post dose lactose PO
C4071008|T201|COMP|78515-4|LNC|Lactose^15M post dose lactose PO|Lactose^15M post dose lactose PO
C4071044|T201|COMP|78445-4|LNC|Cytomegalovirus Ab.IgG avidity|Cytomegalovirus Ab.IgG avidity
C4071045|T201|COMP|78444-7|LNC|Hepatitis A virus Ab.IgG+IgM|Hepatitis A virus Ab.IgG+IgM
C4071046|T201|COMP|78442-1|LNC|Bilirubin.non-glucuronidated|Bilirubin.non-glucuronidated
C4071047|T201|COMP|78441-3|LNC|Bilirubin.glucuronidated|Bilirubin.glucuronidated
C4071048|T201|COMP|78440-5|LNC|Risperidone trough & 9-Hydroxyrisperidone panel|Risperidone trough & 9-Hydroxyrisperidone panel
C4071049|T201|COMP|78439-7|LNC|Phenytoin free & total trough panel|Phenytoin free & total trough panel
C4071050|T201|COMP|78438-9|LNC|Sertraline trough & Norsertraline panel|Sertraline trough & Norsertraline panel
C4071052|T201|COMP|78436-3|LNC|Primidone & PHENobarbital trough panel|Primidone & PHENobarbital trough panel
C4071053|T201|COMP|78435-5|LNC|Mirtazapine trough & Normirtazapine panel|Mirtazapine trough & Normirtazapine panel
C4071091|T201|COMP|78384-5|LNC|Cat dander native (nFel d) 1 Ab.IgE|Cat dander native (nFel d) 1 Ab.IgE
C4071093|T201|COMP|78382-9|LNC|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C4071096|T201|COMP|78379-5|LNC|Epipregnanolone|Epipregnanolone
C4071097|T201|COMP|78378-7|LNC|PON1 gene.c.575A>G|PON1 gene.c.575A>G
C4071098|T201|COMP|78377-9|LNC|Epipregnanolone|Epipregnanolone
C4071099|T201|COMP|78376-1|LNC|Epipregnanolone|Epipregnanolone
C4071101|T201|COMP|78374-6|LNC|Dermatophagoides farinae native (nDer f) 2 Ab.IgE|Dermatophagoides farinae native (nDer f) 2 Ab.IgE
C4071106|T201|COMP|78368-8|LNC|Parrot serum proteins+feathers+droppings Ab.IgG|Parrot serum proteins+feathers+droppings Ab.IgG
C4071107|T201|COMP|78367-0|LNC|Pigeon serum proteins+feathers+droppings Ab.IgG|Pigeon serum proteins+feathers+droppings Ab.IgG
C4071108|T201|COMP|78366-2|LNC|Goose feather Ab.IgG|Goose feather Ab.IgG
C4071110|T201|COMP|78364-7|LNC|Amphetamine cutoff|Amphetamine cutoff
C4071111|T201|COMP|78363-9|LNC|Norhydrocodone|Norhydrocodone
C4071112|T201|COMP|78362-1|LNC|Imipramine+Desipramine^trough|Imipramine+Desipramine^trough
C4071113|T201|COMP|78361-3|LNC|Fatty acid & triglyceride panel|Fatty acid & triglyceride panel
C4071114|T201|COMP|78360-5|LNC|Acyl CoA dehydrogenases|Acyl CoA dehydrogenases
C4071116|T201|COMP|78358-9|LNC|Acyl CoA dehydrogenases|Acyl CoA dehydrogenases
C4071117|T201|COMP|78357-1|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C4071118|T201|COMP|78356-3|LNC|Bacteria identified|Bacteria identified
C4071119|T201|COMP|78355-5|LNC|Lymphocytes.abnormal|Lymphocytes.abnormal
C4071121|T201|COMP|78353-0|LNC|Hexadecadienoate|Hexadecadienoate
C4071122|T201|COMP|78352-2|LNC|Vaccenate|Vaccenate
C4071123|T201|COMP|78351-4|LNC|Tetradecadienoate|Tetradecadienoate
C4071124|T201|COMP|78350-6|LNC|Decenoate|Decenoate
C4071125|T201|COMP|78349-8|LNC|Lauroleate|Lauroleate
C4071126|T201|COMP|78348-0|LNC|Docosapentaenate w6|Docosapentaenate w6
C4071127|T201|COMP|78347-2|LNC|Docosapentaenate w3|Docosapentaenate w3
C4071128|T201|COMP|78346-4|LNC|Hexadecenoate|Hexadecenoate
C4071129|T201|COMP|78345-6|LNC|Docosenoate|Docosenoate
C4071130|T201|COMP|78344-9|LNC|Fatty acid panel.comprehensive C8-C26|Fatty acid panel.comprehensive C8-C26
C4071131|T201|COMP|78343-1|LNC|Cells.MYB gene deletion/Cells counted|Cells.MYB gene deletion/Cells counted
C4071132|T201|COMP|78342-3|LNC|MYB gene deletion|MYB gene deletion
C4071189|T201|COMP|78245-8|LNC|MYB gene deletion|MYB gene deletion
C4071196|T201|COMP|78238-3|LNC|Chromosome 3 copy number/nucleus|Chromosome 3 copy number/nucleus
C4071197|T201|COMP|78237-5|LNC|Chromosome 8 copy number/nucleus|Chromosome 8 copy number/nucleus
C4071198|T201|COMP|78236-7|LNC|Cells.IGH gene rearrangements/Cells counted|Cells.IGH gene rearrangements/Cells counted
C4071199|T201|COMP|78235-9|LNC|Cells.PDGFRB gene rearrangements/Cells counted|Cells.PDGFRB gene rearrangements/Cells counted
C4071200|T201|COMP|78234-2|LNC|Cells.MLL gene rearrangements/Cells counted|Cells.MLL gene rearrangements/Cells counted
C4071201|T201|COMP|78233-4|LNC|Cells.ALK gene rearrangements/Cells counted|Cells.ALK gene rearrangements/Cells counted
C4071202|T201|COMP|78232-6|LNC|Cells.BCL2 gene rearrangements/Cells counted|Cells.BCL2 gene rearrangements/Cells counted
C4071203|T201|COMP|78231-8|LNC|Cells.TRA+TRD gene rearrangements/Cells counted|Cells.TRA+TRD gene rearrangements/Cells counted
C4071204|T201|COMP|78230-0|LNC|Cells.RARA gene rearrangements/Cells counted|Cells.RARA gene rearrangements/Cells counted
C4071205|T201|COMP|78229-2|LNC|Cells.MYC gene rearrangements/Cells counted|Cells.MYC gene rearrangements/Cells counted
C4071206|T201|COMP|78228-4|LNC|IGH gene rearrangements|IGH gene rearrangements
C4071207|T201|COMP|78227-6|LNC|PDGFRB gene rearrangements|PDGFRB gene rearrangements
C4071208|T201|COMP|78226-8|LNC|MLL gene rearrangements|MLL gene rearrangements
C4071209|T201|COMP|78225-0|LNC|BCL2 gene rearrangements|BCL2 gene rearrangements
C4071210|T201|COMP|78224-3|LNC|RARA gene rearrangements|RARA gene rearrangements
C4071211|T201|COMP|78223-5|LNC|TRA+TRD gene rearrangements|TRA+TRD gene rearrangements
C4071212|T201|COMP|78222-7|LNC|MYC gene rearrangements|MYC gene rearrangements
C4071213|T201|COMP|78218-5|LNC|BCL2 gene rearrangements|BCL2 gene rearrangements
C4071214|T201|COMP|78217-7|LNC|RARA gene rearrangements|RARA gene rearrangements
C4071215|T201|COMP|78216-9|LNC|TRA+TRD gene rearrangements|TRA+TRD gene rearrangements
C4071216|T201|COMP|78215-1|LNC|MYC gene rearrangements|MYC gene rearrangements
C4071217|T201|COMP|78214-4|LNC|Cells.CCND1 gene duplication/Cells counted|Cells.CCND1 gene duplication/Cells counted
C4071218|T201|COMP|78213-6|LNC|Cells.BCL6 gene rearrangements/Cells counted|Cells.BCL6 gene rearrangements/Cells counted
C4071221|T201|COMP|78210-2|LNC|ALK gene rearrangements|ALK gene rearrangements
C4071222|T201|COMP|78209-4|LNC|CCND1 gene duplication|CCND1 gene duplication
C4071223|T201|COMP|78208-6|LNC|BCL6 gene rearrangements|BCL6 gene rearrangements
C4071224|T201|COMP|78207-8|LNC|9q34 chromosome region deletion|9q34 chromosome region deletion
C4071225|T201|COMP|78206-0|LNC|4q12 chromosome region rearrangements|4q12 chromosome region rearrangements
C4071226|T201|COMP|78205-2|LNC|ALK gene rearrangements|ALK gene rearrangements
C4071227|T201|COMP|78204-5|LNC|CCND1 gene duplication|CCND1 gene duplication
C4071228|T201|COMP|78203-7|LNC|BCL6 gene rearrangements|BCL6 gene rearrangements
C4071229|T201|COMP|78202-9|LNC|9q34 chromosome region deletion|9q34 chromosome region deletion
C4071230|T201|COMP|78201-1|LNC|4q12 chromosome region rearrangements|4q12 chromosome region rearrangements
C4071231|T201|COMP|78200-3|LNC|Resource identifier|Resource identifier
C4071345|T201|COMP|78221-9|LNC|IGH gene rearrangements|IGH gene rearrangements
C4071346|T201|COMP|78220-1|LNC|PDGFRB gene rearrangements|PDGFRB gene rearrangements
C4071347|T201|COMP|78219-3|LNC|MLL gene rearrangements|MLL gene rearrangements
C4071389|T201|COMP|78047-8|LNC|Cortisol^24H post XXX challenge|Cortisol^24H post XXX challenge
C4071393|T201|COMP|78043-7|LNC|Gene mutations tested for|Gene mutations tested for
C4071394|T201|COMP|78012-2|LNC|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C4071401|T201|COMP|79618-5|LNC|L-serine|L-serine
C4071402|T201|COMP|79617-7|LNC|Glycylproline|Glycylproline
C4071403|T201|COMP|79616-9|LNC|S-beta aminoisobutyrate|S-beta aminoisobutyrate
C4071404|T201|COMP|79615-1|LNC|R-beta aminoisobutyrate|R-beta aminoisobutyrate
C4071405|T201|COMP|79614-4|LNC|N-monomethylarginine|N-monomethylarginine
C4071407|T201|COMP|79612-8|LNC|L-homoarginine|L-homoarginine
C4071410|T201|COMP|79347-1|LNC|Sulfate.total/Creatinine|Sulfate.total/Creatinine
C4071411|T201|COMP|79346-3|LNC|Alpha-aminoadipic semialdehyde/Creatinine|Alpha-aminoadipic semialdehyde/Creatinine
C4071414|T201|COMP|79343-0|LNC|Dimethylacetals pattern|Dimethylacetals pattern
C4071416|T201|COMP|79160-8|LNC|Cold agglutinin panel|Cold agglutinin panel
C4071417|T201|COMP|79159-0|LNC|Cold agglutinin^24H post incubation|Cold agglutinin^24H post incubation
C4071418|T201|COMP|79158-2|LNC|Cold agglutinin^1H post incubation|Cold agglutinin^1H post incubation
C4071419|T201|COMP|79157-4|LNC|Cold agglutinin^1H post incubation|Cold agglutinin^1H post incubation
C4071420|T201|COMP|79156-6|LNC|Cold agglutinin^1H post incubation|Cold agglutinin^1H post incubation
C4071452|T201|COMP|79383-6|LNC|Salmonella sp rpoD gene|Salmonella sp rpoD gene
C4071495|T201|COMP|77959-5|LNC|Yellow fever virus ns5 gene|Yellow fever virus ns5 gene
C4071496|T201|COMP|77670-8|LNC|Gastrin^pre XXX challenge|Gastrin^pre XXX challenge
C4071497|T201|COMP|78042-9|LNC|Vendor FISH product name|Vendor FISH product name
C4071498|T201|COMP|78041-1|LNC|FISH probe target locus|FISH probe target locus
C4071499|T201|COMP|78040-3|LNC|FISH probe target gene|FISH probe target gene
C4071565|T201|COMP|76136-1|LNC|Lactulose^post XXX g sugar solution PO|Lactulose^post XXX g sugar solution PO
C4071567|T201|COMP|76134-6|LNC|Sucrose^post XXX g sugar solution PO|Sucrose^post XXX g sugar solution PO
C4071568|T201|COMP|76133-8|LNC|Sugar absorption test panel|Sugar absorption test panel
C4071631|T201|COMP|75940-7|LNC|Potassium|Potassium
C4071638|T201|COMP|75928-2|LNC|Hemoglobin|Hemoglobin
C4071655|T201|COMP|74533-1|LNC|Fatty acid oxidation panel|Fatty acid oxidation panel
C4071752|T201|COMP|60840-6|LNC|Base excess|Base excess
C4071755|T201|COMP|78791-1|LNC|Amprenavir^trough|Amprenavir^trough
C4071756|T201|COMP|7873-3|LNC|Echovirus NOS Ab|Echovirus NOS Ab
C4071757|T201|COMP|78443-9|LNC|carBAMazepine 10,11-Epoxide^trough|carBAMazepine 10,11-Epoxide^trough
C4071758|T201|COMP|77191-5|LNC|Human epididymis protein 4|Human epididymis protein 4
C4082220|T201|COMP|4107-9|LNC|Acyclovir|Acyclovir
C4082221|T201|COMP|4123-6|LNC|Amoxicillin|Amoxicillin
C4082222|T201|COMP|4132-7|LNC|Atenolol|Atenolol
C4082223|T201|COMP|4133-5|LNC|Atropine|Atropine
C4082224|T201|COMP|4150-9|LNC|Caffeine|Caffeine
C4082225|T201|COMP|4170-7|LNC|Cephalexin|Cephalexin
C4082226|T201|COMP|4186-3|LNC|Ciprofloxacin|Ciprofloxacin
C4082227|T201|COMP|4187-1|LNC|CISplatin|CISplatin
C4082228|T201|COMP|4189-7|LNC|Clindamycin|Clindamycin
C4082229|T201|COMP|4199-6|LNC|Codeine|Codeine
C4082230|T201|COMP|4212-7|LNC|Desipramine|Desipramine
C4082231|T201|COMP|4222-6|LNC|Digoxin|Digoxin
C4082232|T201|COMP|4281-2|LNC|Ibuprofen|Ibuprofen
C4082233|T201|COMP|4300-0|LNC|Lithium|Lithium
C4082234|T201|COMP|4307-5|LNC|Meperidine|Meperidine
C4082235|T201|COMP|4318-2|LNC|Methadone|Methadone
C4082236|T201|COMP|4331-5|LNC|Metoprolol|Metoprolol
C4082237|T201|COMP|4337-2|LNC|Morphine|Morphine
C4082238|T201|COMP|4370-3|LNC|oxyCODONE|oxyCODONE
C4082239|T201|COMP|4445-3|LNC|Tobramycin|Tobramycin
C4082240|T201|COMP|4459-4|LNC|Vancomycin|Vancomycin
C4082241|T201|COMP|4460-2|LNC|Verapamil|Verapamil
C4082242|T201|COMP|4461-0|LNC|Warfarin|Warfarin
C4082867|T201|COMP|32589-4|LNC|Gabapentin|Gabapentin
C4255034|T201|COMP|81250-3|LNC|Simple variant panel|Simple variant panel
C4255038|T201|COMP|81959-9|LNC|Public health laboratory ask at order entry panel|Public health laboratory ask at order entry panel
C4255111|T201|COMP|81303-0|LNC|HGVS version|HGVS version
C4255112|T201|COMP|81297-4|LNC|Structural variant panel|Structural variant panel
C4255115|T201|COMP|81291-7|LNC|Structural variant ISCN name|Structural variant ISCN name
C4255116|T201|COMP|81290-9|LNC|Genomic DNA change|Genomic DNA change
C4255159|T201|COMP|81878-1|LNC|Subtelomere analysis|Subtelomere analysis
C4255246|T201|COMP|81750-2|LNC|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript
C4255285|T201|COMP|81263-6|LNC|Complex variant type|Complex variant type
C4255286|T201|COMP|81262-8|LNC|Complex variant HGVS name|Complex variant HGVS name
C4255287|T201|COMP|81259-4|LNC|Associated phenotype|Associated phenotype
C4255288|T201|COMP|81258-6|LNC|Sample variant allelic frequency|Sample variant allelic frequency
C4255290|T201|COMP|81251-1|LNC|Complex variant panel|Complex variant panel
C4255299|T201|COMP|81857-5|LNC|GDAP1 gene targeted mutation analysis|GDAP1 gene targeted mutation analysis
C4255301|T201|COMP|82155-3|LNC|Genomic structural variant copy number|Genomic structural variant copy number
C4255303|T201|COMP|82154-6|LNC|Genomic structural variant name|Genomic structural variant name
C4255336|T201|COMP|62327-2|LNC|Post-discharge provider practice address|Post-discharge provider practice address
C4255337|T201|COMP|62326-4|LNC|Post-discharge provider practice name|Post-discharge provider practice name
C4255338|T201|COMP|62325-6|LNC|Post-discharge provider practice ID|Post-discharge provider practice ID
C4255339|T201|COMP|62323-1|LNC|Post-discharge provider ID|Post-discharge provider ID
C4255358|T201|COMP|80688-5|LNC|HIV 1 RNA tropism|HIV 1 RNA tropism
C4255382|T201|COMP|81139-8|LNC|CYP3A4 gene targeted mutation analysis|CYP3A4 gene targeted mutation analysis
C4255430|T201|COMP|80687-7|LNC|CYP1A2 gene targeted mutation analysis|CYP1A2 gene targeted mutation analysis
C4255431|T201|COMP|80686-9|LNC|CYP2C9 gene targeted mutation analysis|CYP2C9 gene targeted mutation analysis
C4255442|T201|COMP|81247-9|LNC|Master HL7 genetic variant reporting panel|Master HL7 genetic variant reporting panel
C4255472|T201|COMP|82117-3|LNC|Medication usage implications panel|Medication usage implications panel
C4255475|T201|COMP|82115-7|LNC|dbSNP version|dbSNP version
C4255498|T201|COMP|82118-1|LNC|Pharmacogenomics result panel|Pharmacogenomics result panel
C4255505|T201|COMP|82120-7|LNC|Allelic phase|Allelic phase
C4255506|T201|COMP|82121-5|LNC|Allelic read depth|Allelic read depth
C4255511|T201|COMP|81868-2|LNC|PRNP gene targeted mutation analysis|PRNP gene targeted mutation analysis
C4264627|T201|COMP|82024-1|LNC|Phadiatop Infant Ab.IgE.RAST class|Phadiatop Infant Ab.IgE.RAST class
C4264632|T201|COMP|81785-8|LNC|Duck feather Ab.IgG|Duck feather Ab.IgG
C4264633|T201|COMP|81774-2|LNC|Actin.smooth muscle Ab.IgG|Actin.smooth muscle Ab.IgG
C4264634|T201|COMP|80823-8|LNC|Zika virus Ab.IgM|Zika virus Ab.IgM
C4264640|T201|COMP|81627-2|LNC|Methotrexate diglutamate|Methotrexate diglutamate
C4264641|T201|COMP|80636-4|LNC|Alpha-amanitin|Alpha-amanitin
C4264643|T201|COMP|80588-7|LNC|Influenza virus A M gene|Influenza virus A M gene
C4264677|T201|COMP|82258-5|LNC|Subtelomere analysis|Subtelomere analysis
C4264678|T201|COMP|82257-7|LNC|SRY gene deletion|SRY gene deletion
C4264680|T201|COMP|82255-1|LNC|Marker & derivative chromosome analysis|Marker & derivative chromosome analysis
C4264681|T201|COMP|82254-4|LNC|Marker & derivative chromosome analysis|Marker & derivative chromosome analysis
C4264682|T201|COMP|82253-6|LNC|JAG1 gene deletion|JAG1 gene deletion
C4264683|T201|COMP|82252-8|LNC|Constitutive heterochromatin analysis|Constitutive heterochromatin analysis
C4264686|T201|COMP|82249-4|LNC|Chromosome region 8q23.3-24.13 deletion|Chromosome region 8q23.3-24.13 deletion
C4264687|T201|COMP|82248-6|LNC|Chromosome region 7q11.23 deletion|Chromosome region 7q11.23 deletion
C4264688|T201|COMP|82247-8|LNC|Chromosome region 7q11.23 deletion|Chromosome region 7q11.23 deletion
C4264689|T201|COMP|82246-0|LNC|Chromosome region 22q11.2 deletion+duplication|Chromosome region 22q11.2 deletion+duplication
C4264690|T201|COMP|82245-2|LNC|Chromosome region 22q11.2 deletion+duplication|Chromosome region 22q11.2 deletion+duplication
C4264691|T201|COMP|82244-5|LNC|Chromosome region 1p36 deletion|Chromosome region 1p36 deletion
C4264692|T201|COMP|82243-7|LNC|Chromosome region 17p13.3 deletion|Chromosome region 17p13.3 deletion
C4264693|T201|COMP|82242-9|LNC|Chromosome region 17p13.3 deletion|Chromosome region 17p13.3 deletion
C4264694|T201|COMP|82241-1|LNC|Chromosome region 17p11.2 deletion|Chromosome region 17p11.2 deletion
C4264695|T201|COMP|82240-3|LNC|Chromosome region 16p13.3 deletion|Chromosome region 16p13.3 deletion
C4264696|T201|COMP|82239-5|LNC|Chromosome region 16p13.3 deletion|Chromosome region 16p13.3 deletion
C4264697|T201|COMP|82238-7|LNC|Chromosome region 15q11-13 deletion+duplication|Chromosome region 15q11-13 deletion+duplication
C4264709|T201|COMP|82213-0|LNC|Sapovirus genogroups I+II+IV+V RNA|Sapovirus genogroups I+II+IV+V RNA
C4264710|T201|COMP|82212-2|LNC|Rotavirus A RNA|Rotavirus A RNA
C4264711|T201|COMP|82211-4|LNC|Norovirus genogroup I+II RNA|Norovirus genogroup I+II RNA
C4264712|T201|COMP|82210-6|LNC|Astrovirus subtypes 1-8 RNA|Astrovirus subtypes 1-8 RNA
C4264713|T201|COMP|82209-8|LNC|Adenovirus 40+41 DNA|Adenovirus 40+41 DNA
C4264714|T201|COMP|82208-0|LNC|Giardia lamblia DNA|Giardia lamblia DNA
C4264715|T201|COMP|82207-2|LNC|Entamoeba histolytica DNA|Entamoeba histolytica DNA
C4264716|T201|COMP|82206-4|LNC|Cyclospora cayetanensis DNA|Cyclospora cayetanensis DNA
C4264717|T201|COMP|82205-6|LNC|Cryptosporidium sp DNA|Cryptosporidium sp DNA
C4264718|T201|COMP|82204-9|LNC|Escherichia coli O157 DNA|Escherichia coli O157 DNA
C4264719|T201|COMP|82203-1|LNC|Escherichia coli Stx1+Stx2 toxin stx1+stx2 genes|Escherichia coli Stx1+Stx2 toxin stx1+stx2 genes
C4264720|T201|COMP|82202-3|LNC|Yersinia enterocolitica DNA|Yersinia enterocolitica DNA
C4264721|T201|COMP|82201-5|LNC|Vibrio cholerae DNA|Vibrio cholerae DNA
C4264722|T201|COMP|82200-7|LNC|Vibrio cholerae+parahaemolyticus+vulnificus DNA|Vibrio cholerae+parahaemolyticus+vulnificus DNA
C4264723|T201|COMP|82199-1|LNC|Salmonella enterica+bongori DNA|Salmonella enterica+bongori DNA
C4264724|T201|COMP|82198-3|LNC|Plesiomonas shigelloides DNA|Plesiomonas shigelloides DNA
C4264726|T201|COMP|82196-7|LNC|Campylobacter coli+jejuni+upsaliensis DNA|Campylobacter coli+jejuni+upsaliensis DNA
C4264727|T201|COMP|82195-9|LNC|Gastrointestinal pathogens DNA & RNA panel|Gastrointestinal pathogens DNA & RNA panel
C4264728|T201|COMP|82194-2|LNC|Enterovirus RNA|Enterovirus RNA
C4264729|T201|COMP|82193-4|LNC|Parechovirus A RNA|Parechovirus A RNA
C4264730|T201|COMP|82192-6|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C4264731|T201|COMP|82191-8|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C4264732|T201|COMP|82190-0|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C4264733|T201|COMP|82189-2|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C4264734|T201|COMP|82188-4|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C4264735|T201|COMP|82187-6|LNC|Streptococcus pneumoniae DNA|Streptococcus pneumoniae DNA
C4264736|T201|COMP|82186-8|LNC|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C4264737|T201|COMP|82185-0|LNC|Neisseria meningitidis DNA|Neisseria meningitidis DNA
C4264738|T201|COMP|82184-3|LNC|Listeria monocytogenes DNA|Listeria monocytogenes DNA
C4264739|T201|COMP|82183-5|LNC|Haemophilus influenzae DNA|Haemophilus influenzae DNA
C4264740|T201|COMP|82182-7|LNC|Escherichia coli K1 DNA|Escherichia coli K1 DNA
C4264741|T201|COMP|82181-9|LNC|Cryptococcus gattii+neoformans DNA|Cryptococcus gattii+neoformans DNA
C4264742|T201|COMP|82180-1|LNC|Meningitis+Encephalitis pathogens DNA & RNA panel|Meningitis+Encephalitis pathogens DNA & RNA panel
C4264744|T201|COMP|82178-5|LNC|Chlamydophila pneumoniae DNA|Chlamydophila pneumoniae DNA
C4264745|T201|COMP|82177-7|LNC|Mycoplasma pneumoniae DNA|Mycoplasma pneumoniae DNA
C4264746|T201|COMP|82176-9|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C4264747|T201|COMP|82175-1|LNC|Rhinovirus+Enterovirus RNA|Rhinovirus+Enterovirus RNA
C4264748|T201|COMP|82174-4|LNC|Parainfluenza virus 4 RNA|Parainfluenza virus 4 RNA
C4264749|T201|COMP|82173-6|LNC|Parainfluenza virus 3 RNA|Parainfluenza virus 3 RNA
C4264750|T201|COMP|82172-8|LNC|Parainfluenza virus 2 RNA|Parainfluenza virus 2 RNA
C4264751|T201|COMP|82171-0|LNC|Parainfluenza virus 1 RNA|Parainfluenza virus 1 RNA
C4264752|T201|COMP|82170-2|LNC|Influenza virus B RNA|Influenza virus B RNA
C4264753|T201|COMP|82169-4|LNC|Influenza virus A H3 RNA|Influenza virus A H3 RNA
C4264754|T201|COMP|82168-6|LNC|Influenza virus A H1 2009 pandemic RNA|Influenza virus A H1 2009 pandemic RNA
C4264755|T201|COMP|82167-8|LNC|Influenza virus A H1 RNA|Influenza virus A H1 RNA
C4264756|T201|COMP|82166-0|LNC|Influenza virus A RNA|Influenza virus A RNA
C4264757|T201|COMP|82162-9|LNC|Human coronavirus NL63 RNA|Human coronavirus NL63 RNA
C4264758|T201|COMP|82161-1|LNC|Human coronavirus HKU1 RNA|Human coronavirus HKU1 RNA
C4264759|T201|COMP|82160-3|LNC|Adenovirus DNA|Adenovirus DNA
C4264760|T201|COMP|82159-5|LNC|Respiratory pathogens DNA & RNA panel|Respiratory pathogens DNA & RNA panel
C4264777|T201|COMP|82140-5|LNC|MYD88 gene.p.Leu265Pro targeted mutation analysis|MYD88 gene.p.Leu265Pro targeted mutation analysis
C4264779|T201|COMP|82138-9|LNC|GJB2 gene.c.35delG targeted mutation analysis|GJB2 gene.c.35delG targeted mutation analysis
C4264780|T201|COMP|82137-1|LNC|FGFR3 gene.p.Gly380Arg targeted mutation analysis|FGFR3 gene.p.Gly380Arg targeted mutation analysis
C4264782|T201|COMP|82135-5|LNC|Respiratory pathogens DNA & RNA tested for|Respiratory pathogens DNA & RNA tested for
C4264783|T201|COMP|82134-8|LNC|Respiratory pathogens DNA & RNA tested for|Respiratory pathogens DNA & RNA tested for
C4264790|T201|COMP|82127-2|LNC|Respiratory pathogens DNA & RNA identified|Respiratory pathogens DNA & RNA identified
C4264792|T201|COMP|82125-6|LNC|Respiratory pathogens DNA & RNA tested for|Respiratory pathogens DNA & RNA tested for
C4264795|T201|COMP|82122-3|LNC|Variant coding system|Variant coding system
C4264796|T201|COMP|82119-9|LNC|COSMIC structural variant|COSMIC structural variant
C4264797|T201|COMP|82116-5|LNC|Medication usage suggestion|Medication usage suggestion
C4264836|T201|COMP|82075-3|LNC|(Beef+Chicken+Pork) Ab.IgE.RAST class|(Beef+Chicken+Pork) Ab.IgE.RAST class
C4264876|T201|COMP|82029-0|LNC|Olea europaea native (nOle e) 1 Ab.IgE.RAST class|Olea europaea native (nOle e) 1 Ab.IgE.RAST class
C4264877|T201|COMP|82028-2|LNC|Elaeagnus angustifolia Ab.IgE.RAST class|Elaeagnus angustifolia Ab.IgE.RAST class
C4264878|T201|COMP|82027-4|LNC|Ulmus crassifolia Ab.IgE.RAST class|Ulmus crassifolia Ab.IgE.RAST class
C4264879|T201|COMP|82026-6|LNC|Bromelin MUXF3 Ab.IgE.RAST class|Bromelin MUXF3 Ab.IgE.RAST class
C4264880|T201|COMP|82025-8|LNC|Epinephelus lanceolatus Ab.IgE.RAST class|Epinephelus lanceolatus Ab.IgE.RAST class
C4264881|T201|COMP|82023-3|LNC|Phadiatop Ab.IgE.RAST class|Phadiatop Ab.IgE.RAST class
C4264882|T201|COMP|82022-5|LNC|Galactose-alpha-1,3-galactose Ab.IgE.RAST class|Galactose-alpha-1,3-galactose Ab.IgE.RAST class
C4264884|T201|COMP|82020-9|LNC|Aspergillus flavus Ab.IgE.RAST class|Aspergillus flavus Ab.IgE.RAST class
C4264885|T201|COMP|82019-1|LNC|Termamyl Ab.IgE.RAST class|Termamyl Ab.IgE.RAST class
C4264886|T201|COMP|82018-3|LNC|Lipolase Ab.IgE.RAST class|Lipolase Ab.IgE.RAST class
C4264887|T201|COMP|82017-5|LNC|Latex recombinant (rHev b) 11 Ab.IgE.RAST class|Latex recombinant (rHev b) 11 Ab.IgE.RAST class
C4264888|T201|COMP|82016-7|LNC|Latex recombinant (rHev b) 9 Ab.IgE.RAST class|Latex recombinant (rHev b) 9 Ab.IgE.RAST class
C4264889|T201|COMP|82011-8|LNC|Latex recombinant (rHev b) 3 Ab.IgE.RAST class|Latex recombinant (rHev b) 3 Ab.IgE.RAST class
C4264890|T201|COMP|82010-0|LNC|Latex recombinant (rHev b) 1 Ab.IgE.RAST class|Latex recombinant (rHev b) 1 Ab.IgE.RAST class
C4264892|T201|COMP|82008-4|LNC|Polistes dominulus Ab.IgE.RAST class|Polistes dominulus Ab.IgE.RAST class
C4264894|T201|COMP|82006-8|LNC|House dust Bencard Ab.IgE.RAST class|House dust Bencard Ab.IgE.RAST class
C4264897|T201|COMP|82003-5|LNC|Dioscorea batatas Ab.IgE.RAST class|Dioscorea batatas Ab.IgE.RAST class
C4264902|T201|COMP|81998-7|LNC|Glycine max native (nGly m) 6 Ab.IgE.RAST class|Glycine max native (nGly m) 6 Ab.IgE.RAST class
C4264903|T201|COMP|81997-9|LNC|Glycine max native (nGly m) 5 Ab.IgE.RAST class|Glycine max native (nGly m) 5 Ab.IgE.RAST class
C4264919|T201|COMP|81981-3|LNC|Conalbumin native (nGal d) 3 Ab.IgE.RAST class|Conalbumin native (nGal d) 3 Ab.IgE.RAST class
C4264920|T201|COMP|81980-5|LNC|Cat recombinant (rFel d) 1 Ab.IgE.RAST class|Cat recombinant (rFel d) 1 Ab.IgE.RAST class
C4264921|T201|COMP|81979-7|LNC|Cat recombinant (rFel d) 4 Ab.IgE.RAST class|Cat recombinant (rFel d) 4 Ab.IgE.RAST class
C4264922|T201|COMP|81978-9|LNC|Horse recombinant (rEqu c) 1 Ab.IgE.RAST class|Horse recombinant (rEqu c) 1 Ab.IgE.RAST class
C4264923|T201|COMP|81977-1|LNC|Dog recombinant (rCan f) 5 Ab.IgE.RAST class|Dog recombinant (rCan f) 5 Ab.IgE.RAST class
C4264924|T201|COMP|81976-3|LNC|Dog recombinant (rCan f) 2 Ab.IgE.RAST class|Dog recombinant (rCan f) 2 Ab.IgE.RAST class
C4264925|T201|COMP|81975-5|LNC|Dog recombinant (rCan f) 1 Ab.IgE.RAST class|Dog recombinant (rCan f) 1 Ab.IgE.RAST class
C4264929|T201|COMP|81971-4|LNC|Pholcodine Ab.IgE.RAST class|Pholcodine Ab.IgE.RAST class
C4264930|T201|COMP|81970-6|LNC|Codeine Ab.IgE.RAST class|Codeine Ab.IgE.RAST class
C4264933|T201|COMP|81967-2|LNC|Salsola kali native (nSal k) 1 Ab.IgE.RAST class|Salsola kali native (nSal k) 1 Ab.IgE.RAST class
C4264939|T201|COMP|81961-5|LNC|Chamaecyparis obtusa Ab.IgE.RAST class|Chamaecyparis obtusa Ab.IgE.RAST class
C4264940|T201|COMP|81960-7|LNC|Olea europaea native (nOle e) 7 Ab.IgE.RAST class|Olea europaea native (nOle e) 7 Ab.IgE.RAST class
C4264993|T201|COMP|81893-0|LNC|Patient satisfaction with healthcare delivery|Patient satisfaction with healthcare delivery
C4265001|T201|COMP|81884-9|LNC|NIPA1 gene & REEP1 gene full mutation analysis|NIPA1 gene & REEP1 gene full mutation analysis
C4265002|T201|COMP|81883-1|LNC|CNBP gene CCTG repeat analysis|CNBP gene CCTG repeat analysis
C4265003|T201|COMP|81882-3|LNC|TSC2 gene & PKD1 gene deletion+duplication|TSC2 gene & PKD1 gene deletion+duplication
C4265010|T201|COMP|81874-0|LNC|SLC12A3 gene full mutation analysis|SLC12A3 gene full mutation analysis
C4265021|T201|COMP|81862-5|LNC|Karyotype^post mitogen stimulation|Karyotype^post mitogen stimulation
C4265022|T201|COMP|81861-7|LNC|Karyotype|Karyotype
C4265024|T201|COMP|81859-1|LNC|GRN gene full mutation analysis|GRN gene full mutation analysis
C4265026|T201|COMP|81856-7|LNC|FMR1 gene CGG repeat analysis|FMR1 gene CGG repeat analysis
C4265027|T201|COMP|81855-9|LNC|DMPK gene CTG repeat analysis|DMPK gene CTG repeat analysis
C4265029|T201|COMP|81853-4|LNC|Chromosome 15 & 16 & 22 aneuploidy|Chromosome 15 & 16 & 22 aneuploidy
C4265030|T201|COMP|81852-6|LNC|Chromosome region 7q11.23 deletion+duplication|Chromosome region 7q11.23 deletion+duplication
C4265035|T201|COMP|81847-6|LNC|C9orf72 gene GGGGCC repeat analysis|C9orf72 gene GGGGCC repeat analysis
C4265036|T201|COMP|81842-7|LNC|BCKDHB gene targeted mutation analysis|BCKDHB gene targeted mutation analysis
C4265037|T201|COMP|81841-9|LNC|MLC1 gene targeted mutation analysis|MLC1 gene targeted mutation analysis
C4265038|T201|COMP|81840-1|LNC|POMGNT1 gene full mutation analysis|POMGNT1 gene full mutation analysis
C4265039|T201|COMP|81839-3|LNC|CLN8 gene targeted mutation analysis|CLN8 gene targeted mutation analysis
C4265040|T201|COMP|81838-5|LNC|PEX1 gene targeted mutation analysis|PEX1 gene targeted mutation analysis
C4265041|T201|COMP|81837-7|LNC|GRHPR gene targeted mutation analysis|GRHPR gene targeted mutation analysis
C4265042|T201|COMP|81836-9|LNC|CTSK gene targeted mutation analysis|CTSK gene targeted mutation analysis
C4265043|T201|COMP|81835-1|LNC|PEX7 gene targeted mutation analysis|PEX7 gene targeted mutation analysis
C4265044|T201|COMP|81834-4|LNC|SLC17A5 gene full mutation analysis|SLC17A5 gene full mutation analysis
C4265045|T201|COMP|81833-6|LNC|ALDH3A2 gene full mutation analysis|ALDH3A2 gene full mutation analysis
C4265046|T201|COMP|81832-8|LNC|SLC26A2 gene targeted mutation analysis|SLC26A2 gene targeted mutation analysis
C4265047|T201|COMP|81831-0|LNC|LAMB3 gene targeted mutation analysis|LAMB3 gene targeted mutation analysis
C4265048|T201|COMP|81830-2|LNC|AGL gene targeted mutation analysis|AGL gene targeted mutation analysis
C4265049|T201|COMP|81829-4|LNC|SDHA gene full mutation analysis|SDHA gene full mutation analysis
C4265050|T201|COMP|81828-6|LNC|SLC37A4 gene targeted mutation analysis|SLC37A4 gene targeted mutation analysis
C4265051|T201|COMP|81827-8|LNC|CNGB3 gene targeted mutation analysis|CNGB3 gene targeted mutation analysis
C4265052|T201|COMP|81826-0|LNC|HGD gene targeted mutation analysis|HGD gene targeted mutation analysis
C4265053|T201|COMP|81825-2|LNC|MAN2B1 gene targeted mutation analysis|MAN2B1 gene targeted mutation analysis
C4265054|T201|COMP|81824-5|LNC|SLC12A6 gene targeted mutation analysis|SLC12A6 gene targeted mutation analysis
C4265055|T201|COMP|81823-7|LNC|SACS gene targeted mutation analysis|SACS gene targeted mutation analysis
C4265056|T201|COMP|81822-9|LNC|BBS10 gene targeted mutation analysis|BBS10 gene targeted mutation analysis
C4265057|T201|COMP|81821-1|LNC|RMRP gene targeted mutation analysis|RMRP gene targeted mutation analysis
C4265058|T201|COMP|81820-3|LNC|ASS1 gene targeted mutation analysis|ASS1 gene targeted mutation analysis
C4265059|T201|COMP|81819-5|LNC|CLN5 gene targeted mutation analysis|CLN5 gene targeted mutation analysis
C4265060|T201|COMP|81818-7|LNC|PMM2 gene targeted mutation analysis|PMM2 gene targeted mutation analysis
C4265061|T201|COMP|81817-9|LNC|MPI gene targeted mutation analysis|MPI gene targeted mutation analysis
C4265062|T201|COMP|81816-1|LNC|OPA3 gene targeted mutation analysis|OPA3 gene targeted mutation analysis
C4265063|T201|COMP|81815-3|LNC|CTNS gene targeted mutation analysis|CTNS gene targeted mutation analysis
C4265064|T201|COMP|81814-6|LNC|HSD17B4 gene targeted mutation analysis|HSD17B4 gene targeted mutation analysis
C4265065|T201|COMP|81813-8|LNC|F11 gene targeted mutation analysis|F11 gene targeted mutation analysis
C4265066|T201|COMP|81812-0|LNC|TPP1 gene targeted mutation analysis|TPP1 gene targeted mutation analysis
C4265067|T201|COMP|81811-2|LNC|3-Hydroxydecanoylcarnitine (C10-OH)|3-Hydroxydecanoylcarnitine (C10-OH)
C4265068|T201|COMP|81810-4|LNC|3-Hydroxydecanoylcarnitine (C10-OH)/creatinine|3-Hydroxydecanoylcarnitine (C10-OH)/creatinine
C4265069|T201|COMP|81809-6|LNC|3-Hydroxydodecanoylcarnitine (C12-OH)/Creatinine|3-Hydroxydodecanoylcarnitine (C12-OH)/Creatinine
C4265070|T201|COMP|81808-8|LNC|Androstenetriol/Creatinine|Androstenetriol/Creatinine
C4265071|T201|COMP|81807-0|LNC|Alpha cortol/Creatinine|Alpha cortol/Creatinine
C4265072|T201|COMP|81806-2|LNC|Alpha cortolone/Creatinine|Alpha cortolone/Creatinine
C4265073|T201|COMP|81801-3|LNC|16-Alpha hydroxydehydroepiandrosterone/Creatinine|16-Alpha hydroxydehydroepiandrosterone/Creatinine
C4265074|T201|COMP|81800-5|LNC|16-Ketoandrostenediol/Creatinine|16-Ketoandrostenediol/Creatinine
C4265075|T201|COMP|81799-9|LNC|16-Alpha hydroxypregnenolone/Creatinine|16-Alpha hydroxypregnenolone/Creatinine
C4265076|T201|COMP|81798-1|LNC|Pregnanediolone/Creatinine|Pregnanediolone/Creatinine
C4265077|T201|COMP|81797-3|LNC|11-Dehydrotetrahydrocorticosterone/Creatinine|11-Dehydrotetrahydrocorticosterone/Creatinine
C4265078|T201|COMP|81796-5|LNC|Tetrahydrocorticosterone/Creatinine|Tetrahydrocorticosterone/Creatinine
C4265079|T201|COMP|81795-7|LNC|Tetrahydrocortisone/Creatinine|Tetrahydrocortisone/Creatinine
C4265080|T201|COMP|81794-0|LNC|Tetrahydrocortisol/Creatinine|Tetrahydrocortisol/Creatinine
C4265081|T201|COMP|81793-2|LNC|Tetrahydrodeoxycortisol/Creatinine|Tetrahydrodeoxycortisol/Creatinine
C4265083|T201|COMP|81791-6|LNC|Malus domestica recombinant (rMal d) 3 Ab.IgE|Malus domestica recombinant (rMal d) 3 Ab.IgE
C4265084|T201|COMP|81790-8|LNC|Juglans regia recombinant (rJug r) 1 Ab.IgE|Juglans regia recombinant (rJug r) 1 Ab.IgE
C4265085|T201|COMP|81789-0|LNC|Juglans regia recombinant (rJug r) 3 Ab.IgE|Juglans regia recombinant (rJug r) 3 Ab.IgE
C4265086|T201|COMP|81788-2|LNC|Corylus avellana recombinant (rCor a) 14 Ab.IgE|Corylus avellana recombinant (rCor a) 14 Ab.IgE
C4265087|T201|COMP|81787-4|LNC|Myeloperoxidase Ab.IgG|Myeloperoxidase Ab.IgG
C4265088|T201|COMP|81786-6|LNC|Chemokine (C-C motif) ligand 17|Chemokine (C-C motif) ligand 17
C4265089|T201|COMP|81784-1|LNC|Canary droppings Ab.IgG|Canary droppings Ab.IgG
C4265090|T201|COMP|81783-3|LNC|Chicken feather Ab.IgG|Chicken feather Ab.IgG
C4265091|T201|COMP|81777-5|LNC|Nonanoylcarnitine (C9)/Creatinine|Nonanoylcarnitine (C9)/Creatinine
C4265092|T201|COMP|81776-7|LNC|Ureidopropionate/Creatinine|Ureidopropionate/Creatinine
C4265093|T201|COMP|81775-9|LNC|Epipregnanolone/Creatinine|Epipregnanolone/Creatinine
C4265094|T201|COMP|81773-4|LNC|Amyloid A|Amyloid A
C4265095|T201|COMP|81772-6|LNC|Dermatophagoides pteronyssinus Ab.IgG|Dermatophagoides pteronyssinus Ab.IgG
C4265096|T201|COMP|81771-8|LNC|Myeloperoxidase Ab.IgG|Myeloperoxidase Ab.IgG
C4265097|T201|COMP|81770-0|LNC|Tiglylcarnitine (C5:1)/Creatinine|Tiglylcarnitine (C5:1)/Creatinine
C4265098|T201|COMP|81769-2|LNC|Adipoylcarnitine (C6-DC)/Creatinine|Adipoylcarnitine (C6-DC)/Creatinine
C4265099|T201|COMP|81768-4|LNC|U1 small nuclear ribonucleoprotein 70kD Ab.IgG|U1 small nuclear ribonucleoprotein 70kD Ab.IgG
C4265100|T201|COMP|81767-6|LNC|Eicosatrienoate|Eicosatrienoate
C4265101|T201|COMP|81766-8|LNC|Eicosatrienoate|Eicosatrienoate
C4265102|T201|COMP|81765-0|LNC|Docosatrienoate|Docosatrienoate
C4265103|T201|COMP|81764-3|LNC|Docosatrienoate|Docosatrienoate
C4265104|T201|COMP|81763-5|LNC|Phytanate & pristanate panel|Phytanate & pristanate panel
C4265107|T201|COMP|81760-1|LNC|Lymphocyte proliferation.anti-CD3.maximum/CD45|Lymphocyte proliferation.anti-CD3.maximum/CD45
C4265108|T201|COMP|81752-8|LNC|Chromosome region 1q21 duplication|Chromosome region 1q21 duplication
C4265110|T201|COMP|81749-4|LNC|Chromosome region 13q14 deletion|Chromosome region 13q14 deletion
C4265112|T201|COMP|81747-8|LNC|Chromosome region 6q22 rearrangements|Chromosome region 6q22 rearrangements
C4265113|T201|COMP|81746-0|LNC|Chromosome region 17p13.1 deletion|Chromosome region 17p13.1 deletion
C4265114|T201|COMP|81744-5|LNC|Submitter's laboratory test method|Submitter's laboratory test method
C4265115|T201|COMP|81743-7|LNC|Th-To Ab|Th-To Ab
C4265116|T201|COMP|81742-9|LNC|Th-To Ab|Th-To Ab
C4265117|T201|COMP|81741-1|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C4265118|T201|COMP|81740-3|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C4265119|T201|COMP|81739-5|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C4265120|T201|COMP|81738-7|LNC|RNA polymerase III RP155 Ab|RNA polymerase III RP155 Ab
C4265121|T201|COMP|81737-9|LNC|RNA polymerase III RP11 Ab|RNA polymerase III RP11 Ab
C4265122|T201|COMP|81736-1|LNC|RNA polymerase III Ab|RNA polymerase III Ab
C4265123|T201|COMP|81735-3|LNC|Ribosomal P Ab|Ribosomal P Ab
C4265124|T201|COMP|81734-6|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C4265125|T201|COMP|81733-8|LNC|PM-SCL-75 Ab|PM-SCL-75 Ab
C4265126|T201|COMP|81732-0|LNC|PM-SCL-100 Ab|PM-SCL-100 Ab
C4265127|T201|COMP|81731-2|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C4265128|T201|COMP|81730-4|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C4265129|T201|COMP|81729-6|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C4265130|T201|COMP|81728-8|LNC|Neuronal nuclear Ab|Neuronal nuclear Ab
C4265131|T201|COMP|81727-0|LNC|Mitochondria M2-3E Ab|Mitochondria M2-3E Ab
C4265132|T201|COMP|81726-2|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C4265133|T201|COMP|81725-4|LNC|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C4265134|T201|COMP|81724-7|LNC|Glomerular basement membrane Ab|Glomerular basement membrane Ab
C4265135|T201|COMP|81723-9|LNC|Ganglioside GT1b Ab.IgM|Ganglioside GT1b Ab.IgM
C4265136|T201|COMP|81722-1|LNC|Ganglioside GT1b Ab.IgG+IgM|Ganglioside GT1b Ab.IgG+IgM
C4265137|T201|COMP|81721-3|LNC|Ganglioside GM2 Ab.IgG+IgM|Ganglioside GM2 Ab.IgG+IgM
C4265138|T201|COMP|81720-5|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C4265139|T201|COMP|81719-7|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C4265140|T201|COMP|81718-9|LNC|Ganglioside GM1 Ab.IgG+IgM|Ganglioside GM1 Ab.IgG+IgM
C4265141|T201|COMP|81717-1|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C4265142|T201|COMP|81716-3|LNC|DNA double strand Ab|DNA double strand Ab
C4265143|T201|COMP|81715-5|LNC|Centromere protein B Ab|Centromere protein B Ab
C4265144|T201|COMP|81714-8|LNC|Centromere protein A Ab|Centromere protein A Ab
C4265145|T201|COMP|81713-0|LNC|Actin.smooth muscle Ab|Actin.smooth muscle Ab
C4265146|T201|COMP|81712-2|LNC|Actin.filamentous Ab|Actin.filamentous Ab
C4265147|T201|COMP|81711-4|LNC|Microsatellite instability marker panel|Microsatellite instability marker panel
C4265148|T201|COMP|81710-6|LNC|PTEN gene|PTEN gene
C4265149|T201|COMP|81709-8|LNC|Microsatellite markers exhibiting instability|Microsatellite markers exhibiting instability
C4265151|T201|COMP|81707-2|LNC|Dissection technique|Dissection technique
C4265153|T201|COMP|81705-6|LNC|Serine-threonine protein kinase B-raf|Serine-threonine protein kinase B-raf
C4265154|T201|COMP|81704-9|LNC|Microsatellite instability marker D17S250|Microsatellite instability marker D17S250
C4265155|T201|COMP|81703-1|LNC|Microsatellite instability marker D5S346|Microsatellite instability marker D5S346
C4265156|T201|COMP|81702-3|LNC|Microsatellite instability marker D2S123|Microsatellite instability marker D2S123
C4265157|T201|COMP|81701-5|LNC|Microsatellite instability marker MONO27|Microsatellite instability marker MONO27
C4265158|T201|COMP|81700-7|LNC|Microsatellite instability marker NR24|Microsatellite instability marker NR24
C4265159|T201|COMP|81699-1|LNC|Microsatellite instability marker NR21|Microsatellite instability marker NR21
C4265160|T201|COMP|81698-3|LNC|Microsatellite instability marker BAT26|Microsatellite instability marker BAT26
C4265161|T201|COMP|81697-5|LNC|Microsatellite instability marker BAT25|Microsatellite instability marker BAT25
C4265162|T201|COMP|81696-7|LNC|Microsatellite instability markers assessed|Microsatellite instability markers assessed
C4265163|T201|COMP|81695-9|LNC|Microsatellite instability|Microsatellite instability
C4265164|T201|COMP|81694-2|LNC|Mismatch repair endonuclease PMS2|Mismatch repair endonuclease PMS2
C4265165|T201|COMP|81693-4|LNC|DNA mismatch repair protein Msh6|DNA mismatch repair protein Msh6
C4265166|T201|COMP|81692-6|LNC|DNA mismatch repair protein Msh2|DNA mismatch repair protein Msh2
C4265167|T201|COMP|81691-8|LNC|DNA mismatch repair protein Mlh1|DNA mismatch repair protein Mlh1
C4265168|T201|COMP|81690-0|LNC|Legionella longbeachae 1 & 2 DNA|Legionella longbeachae 1 & 2 DNA
C4265169|T201|COMP|81689-2|LNC|Hendra virus RNA|Hendra virus RNA
C4265170|T201|COMP|81688-4|LNC|Barmah forest virus RNA|Barmah forest virus RNA
C4265182|T201|COMP|81658-7|LNC|Suspected organism|Suspected organism
C4265183|T201|COMP|81657-9|LNC|Salmonella sp spaO gene|Salmonella sp spaO gene
C4265184|T201|COMP|81656-1|LNC|Campylobacter coli+jejuni tuf gene|Campylobacter coli+jejuni tuf gene
C4265185|T201|COMP|81655-3|LNC|Respiratory pathogens DNA & RNA identified|Respiratory pathogens DNA & RNA identified
C4265186|T201|COMP|81654-6|LNC|Repiratory pathogens DNA & RNA|Repiratory pathogens DNA & RNA
C4265188|T201|COMP|81652-0|LNC|HIV 2 RNA|HIV 2 RNA
C4265189|T201|COMP|81651-2|LNC|Murray Valley Encephalitis virus RNA|Murray Valley Encephalitis virus RNA
C4265190|T201|COMP|81650-4|LNC|West Nile virus Kunjin strain RNA|West Nile virus Kunjin strain RNA
C4265191|T201|COMP|81649-6|LNC|Cryptococcus sp rRNA gene|Cryptococcus sp rRNA gene
C4265192|T201|COMP|81648-8|LNC|Clostridium botulinum toxin G botG gene|Clostridium botulinum toxin G botG gene
C4265193|T201|COMP|81647-0|LNC|Clostridium botulinum toxin F botF gene|Clostridium botulinum toxin F botF gene
C4265194|T201|COMP|81646-2|LNC|Clostridium botulinum toxin E botE gene|Clostridium botulinum toxin E botE gene
C4265195|T201|COMP|81645-4|LNC|Clostridium botulinum toxin D botD gene|Clostridium botulinum toxin D botD gene
C4265196|T201|COMP|81644-7|LNC|Clostridium botulinum toxin C botC gene|Clostridium botulinum toxin C botC gene
C4265199|T201|COMP|81641-3|LNC|HIV 2 Ab|HIV 2 Ab
C4265200|T201|COMP|81640-5|LNC|Erythrocytes|Erythrocytes
C4265201|T201|COMP|81639-7|LNC|Heparin dose response slope|Heparin dose response slope
C4265204|T201|COMP|81632-2|LNC|Immunoglobulin light chains panel|Immunoglobulin light chains panel
C4265205|T201|COMP|81631-4|LNC|Methotrexate polyglutamates|Methotrexate polyglutamates
C4265206|T201|COMP|81630-6|LNC|Methotrexate polyglutamates 1-5 & total panel|Methotrexate polyglutamates 1-5 & total panel
C4265207|T201|COMP|81629-8|LNC|Gamma hydroxybutyrate|Gamma hydroxybutyrate
C4265208|T201|COMP|81628-0|LNC|Methotrexate monoglutamate|Methotrexate monoglutamate
C4265209|T201|COMP|81626-4|LNC|Methotrexate triglutamate|Methotrexate triglutamate
C4265210|T201|COMP|81625-6|LNC|Methotrexate tetraglutamate|Methotrexate tetraglutamate
C4265211|T201|COMP|81624-9|LNC|Methotrexate pentaglutamate|Methotrexate pentaglutamate
C4265212|T201|COMP|81623-1|LNC|Calcium oxalate|Calcium oxalate
C4265213|T201|COMP|81622-3|LNC|Hydroxyapatite|Hydroxyapatite
C4265214|T201|COMP|81621-5|LNC|Herpes simplex virus 1 & 2 Ab.IgG panel|Herpes simplex virus 1 & 2 Ab.IgG panel
C4265215|T201|COMP|81620-7|LNC|Differential panel|Differential panel
C4265342|T201|COMP|81439-2|LNC|Human papilloma virus 31+33 DNA|Human papilloma virus 31+33 DNA
C4265347|T201|COMP|81430-1|LNC|Lactate dehydrogenase|Lactate dehydrogenase
C4265348|T201|COMP|81429-3|LNC|Bismuth|Bismuth
C4265349|T201|COMP|81428-5|LNC|Influenza virus A H7 Eurasia RNA|Influenza virus A H7 Eurasia RNA
C4265355|T201|COMP|81422-8|LNC|GATA1 gene exon 2 targeted mutation analysis|GATA1 gene exon 2 targeted mutation analysis
C4265356|T201|COMP|81421-0|LNC|Saccharomyces cerevisiae Ab.IgG|Saccharomyces cerevisiae Ab.IgG
C4265357|T201|COMP|81420-2|LNC|KRAS & NRAS gene targeted mutation analysis|KRAS & NRAS gene targeted mutation analysis
C4265398|T201|COMP|81805-4|LNC|Allo-tetrahydrocorticosterone/Creatinine|Allo-tetrahydrocorticosterone/Creatinine
C4265399|T201|COMP|81804-7|LNC|Allo-tetrahydrocortisol/Creatinine|Allo-tetrahydrocortisol/Creatinine
C4265400|T201|COMP|81803-9|LNC|Beta cortolone/Creatinine|Beta cortolone/Creatinine
C4265403|T201|COMP|81638-9|LNC|Clotting time|Clotting time
C4265404|T201|COMP|81637-1|LNC|Glucose meter to reference method correlation|Glucose meter to reference method correlation
C4265421|T201|COMP|82165-2|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C4265422|T201|COMP|82164-5|LNC|Human coronavirus OC43 RNA|Human coronavirus OC43 RNA
C4265423|T201|COMP|82163-7|LNC|Human coronavirus 229E RNA|Human coronavirus 229E RNA
C4265427|T201|COMP|82015-9|LNC|Latex recombinant (rHev b) 8 Ab.IgE.RAST class|Latex recombinant (rHev b) 8 Ab.IgE.RAST class
C4265428|T201|COMP|82014-2|LNC|Latex recombinant (rHev b) 6.02 Ab.IgE.RAST class|Latex recombinant (rHev b) 6.02 Ab.IgE.RAST class
C4265429|T201|COMP|82013-4|LNC|Latex recombinant (rHev b) 6.01 Ab.IgE.RAST class|Latex recombinant (rHev b) 6.01 Ab.IgE.RAST class
C4265430|T201|COMP|82012-6|LNC|Latex recombinant (rHev b) 5 Ab.IgE.RAST class|Latex recombinant (rHev b) 5 Ab.IgE.RAST class
C4265431|T201|COMP|81846-8|LNC|C9orf72 gene GGGGCC repeat analysis|C9orf72 gene GGGGCC repeat analysis
C4265432|T201|COMP|81845-0|LNC|PALB2 gene full mutation analysis|PALB2 gene full mutation analysis
C4265433|T201|COMP|81844-3|LNC|IVD gene full mutation analysis|IVD gene full mutation analysis
C4265434|T201|COMP|81843-5|LNC|GALC gene targeted mutation analysis|GALC gene targeted mutation analysis
C4265435|T201|COMP|81782-5|LNC|Phleum pratense Ab.IgG|Phleum pratense Ab.IgG
C4265436|T201|COMP|81781-7|LNC|Saccharopine|Saccharopine
C4265437|T201|COMP|81780-9|LNC|Tetradecenoylcarnitine (C14:1)/Creatinine|Tetradecenoylcarnitine (C14:1)/Creatinine
C4265460|T201|COMP|81759-3|LNC|Lymphocyte proliferation.anti-CD28.maximum/CD45|Lymphocyte proliferation.anti-CD28.maximum/CD45
C4265461|T201|COMP|81758-5|LNC|Lymphocyte proliferation.anti-CD28.maximum/CD3|Lymphocyte proliferation.anti-CD28.maximum/CD3
C4265463|T201|COMP|81756-9|LNC|Lymphocyte proliferation.anti-CD3.maximum/CD3|Lymphocyte proliferation.anti-CD3.maximum/CD3
C4265465|T201|COMP|81754-4|LNC|Nortapentadol|Nortapentadol
C4265466|T201|COMP|81753-6|LNC|Somatotropin^1.75H post dose arginine+insulin|Somatotropin^1.75H post dose arginine+insulin
C4265500|T201|COMP|81328-7|LNC|Cytomegalovirus|Cytomegalovirus
C4265501|T201|COMP|81327-9|LNC|Influenza virus B Victoria lineage RNA|Influenza virus B Victoria lineage RNA
C4265502|T201|COMP|81326-1|LNC|Human RNase P RNA|Human RNase P RNA
C4265503|T201|COMP|81325-3|LNC|Influenza virus B Yamagata lineage RNA|Influenza virus B Yamagata lineage RNA
C4265504|T201|COMP|81324-6|LNC|Glucose tolerance 2H gestational panel|Glucose tolerance 2H gestational panel
C4265505|T201|COMP|81323-8|LNC|Urine collection associated observations panel|Urine collection associated observations panel
C4265506|T201|COMP|81322-0|LNC|Glucan 1,4 alpha glucosidase|Glucan 1,4 alpha glucosidase
C4265507|T201|COMP|81321-2|LNC|Influenza virus A H5 Asian RNA|Influenza virus A H5 Asian RNA
C4265508|T201|COMP|81320-4|LNC|Influenza virus A H5 Asian RNA|Influenza virus A H5 Asian RNA
C4265509|T201|COMP|81319-6|LNC|Spermatozoa.progressive|Spermatozoa.progressive
C4265510|T201|COMP|81318-8|LNC|Spermatozoa.normal morphology|Spermatozoa.normal morphology
C4265511|T201|COMP|81317-0|LNC|Additional pathological findings|Additional pathological findings
C4265512|T201|COMP|81316-2|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C4265513|T201|COMP|81315-4|LNC|Lactase|Lactase
C4265514|T201|COMP|81314-7|LNC|Palatinase|Palatinase
C4265515|T201|COMP|81313-9|LNC|Cryoglobulin.complement C3|Cryoglobulin.complement C3
C4265516|T201|COMP|81312-1|LNC|Cryoglobulin.IgM|Cryoglobulin.IgM
C4265517|T201|COMP|81311-3|LNC|Cryoglobulin.IgA|Cryoglobulin.IgA
C4265518|T201|COMP|81310-5|LNC|Carbonic anhydrase 2 Ab|Carbonic anhydrase 2 Ab
C4265519|T201|COMP|81309-7|LNC|Influenza virus B RNA|Influenza virus B RNA
C4265520|T201|COMP|81308-9|LNC|Influenza virus A RNA|Influenza virus A RNA
C4265521|T201|COMP|81307-1|LNC|Influenza virus A H7 Eurasia RNA|Influenza virus A H7 Eurasia RNA
C4265522|T201|COMP|81306-3|LNC|Variables that apply to the overall study|Variables that apply to the overall study
C4265523|T201|COMP|81305-5|LNC|Influenza virus A H1 2009 pandemic RNA|Influenza virus A H1 2009 pandemic RNA
C4265524|T201|COMP|81304-8|LNC|Structural variant analysis method|Structural variant analysis method
C4265525|T201|COMP|81302-2|LNC|Structural variant inner start-end|Structural variant inner start-end
C4265526|T201|COMP|81301-4|LNC|Structural variant outer start-end|Structural variant outer start-end
C4265527|T201|COMP|81300-6|LNC|Structural variant|Structural variant
C4265528|T201|COMP|81299-0|LNC|Structural variant reported arrCGH|Structural variant reported arrCGH
C4265529|T201|COMP|81298-2|LNC|Structural variant cytogenetic location|Structural variant cytogenetic location
C4265530|T201|COMP|81294-1|LNC|Genetic form configuration controls|Genetic form configuration controls
C4265531|T201|COMP|81293-3|LNC|Range(s) of DNA sequences examined|Range(s) of DNA sequences examined
C4265532|T201|COMP|81292-5|LNC|Simple variant|Simple variant
C4265533|T201|COMP|81289-1|LNC|Structural variant|Structural variant
C4265534|T201|COMP|81288-3|LNC|Precision of boundaries|Precision of boundaries
C4265535|T201|COMP|81287-5|LNC|Structural variant reported start-end|Structural variant reported start-end
C4265536|T201|COMP|81286-7|LNC|Structural variant|Structural variant
C4265538|T201|COMP|81284-2|LNC|Malignant cells/100 cells|Malignant cells/100 cells
C4265539|T201|COMP|81283-4|LNC|Spermatozoa.nonprogressive|Spermatozoa.nonprogressive
C4265540|T201|COMP|81282-6|LNC|Spermatozoa.motile|Spermatozoa.motile
C4265541|T201|COMP|81281-8|LNC|Heparin dose response panel|Heparin dose response panel
C4265542|T201|COMP|81280-0|LNC|Differential panel|Differential panel
C4265543|T201|COMP|81279-2|LNC|Meperidine & Normeperidine panel|Meperidine & Normeperidine panel
C4265544|T201|COMP|81278-4|LNC|Meperidine & Normeperidine panel|Meperidine & Normeperidine panel
C4265545|T201|COMP|81277-6|LNC|Fentanyl & Norfentanyl panel|Fentanyl & Norfentanyl panel
C4265546|T201|COMP|81276-8|LNC|Doxepin & Nordoxepin panel|Doxepin & Nordoxepin panel
C4265547|T201|COMP|81275-0|LNC|Fentanyl & Norfentanyl panel|Fentanyl & Norfentanyl panel
C4265548|T201|COMP|81274-3|LNC|Doxepin & Nordoxepin panel|Doxepin & Nordoxepin panel
C4265549|T201|COMP|81273-5|LNC|Fentanyl & Norfentanyl panel|Fentanyl & Norfentanyl panel
C4265550|T201|COMP|81272-7|LNC|Cell Count & Differential panel|Cell Count & Differential panel
C4265553|T201|COMP|81261-0|LNC|Complex variant name|Complex variant name
C4265554|T201|COMP|81260-2|LNC|Complex variant|Complex variant
C4265555|T201|COMP|81257-8|LNC|CIGAR|CIGAR
C4265556|T201|COMP|81256-0|LNC|COSMIC simple variant|COSMIC simple variant
C4265557|T201|COMP|81255-2|LNC|dbSNP|dbSNP
C4265558|T201|COMP|81254-5|LNC|Genomic allele start-end|Genomic allele start-end
C4265559|T201|COMP|81253-7|LNC|Simple variant name|Simple variant name
C4265560|T201|COMP|81252-9|LNC|Simple variant|Simple variant
C4265561|T201|COMP|81249-5|LNC|Default genomic reference sequence coding system|Default genomic reference sequence coding system
C4265564|T201|COMP|81234-7|LNC|Varicella zoster virus Ab.IgG & IgM panel|Varicella zoster virus Ab.IgG & IgM panel
C4265565|T201|COMP|81233-9|LNC|Influenza virus types A & B & subtypes panel|Influenza virus types A & B & subtypes panel
C4265566|T201|COMP|81232-1|LNC|Supersaturation panel|Supersaturation panel
C4265567|T201|COMP|81231-3|LNC|Protein fractions panel|Protein fractions panel
C4265581|T201|COMP|81212-3|LNC|Clomipramine & norclomipramine panel|Clomipramine & norclomipramine panel
C4265582|T201|COMP|81211-5|LNC|Amitriptyline & nortriptyline panel|Amitriptyline & nortriptyline panel
C4265583|T201|COMP|81210-7|LNC|Clomipramine & norclomipramine panel|Clomipramine & norclomipramine panel
C4265584|T201|COMP|81209-9|LNC|Clomipramine & norclomipramine panel|Clomipramine & norclomipramine panel
C4265585|T201|COMP|81208-1|LNC|Amitriptyline & nortriptyline panel|Amitriptyline & nortriptyline panel
C4265586|T201|COMP|81207-3|LNC|Amitriptyline & nortriptyline panel|Amitriptyline & nortriptyline panel
C4265588|T201|COMP|81205-7|LNC|Cryoglobulin IgA & IgG & IgM & C3 panel|Cryoglobulin IgA & IgG & IgM & C3 panel
C4265591|T201|COMP|81201-6|LNC|Phospholipase A2 receptor Ab.IgG|Phospholipase A2 receptor Ab.IgG
C4265593|T201|COMP|81199-2|LNC|Beta-ureidopropionase|Beta-ureidopropionase
C4265600|T201|COMP|81190-1|LNC|Histologic type|Histologic type
C4265601|T201|COMP|81185-1|LNC|Non-regional lymph nodes positive|Non-regional lymph nodes positive
C4265603|T201|COMP|81183-6|LNC|Distance of tumor from closest distal margin|Distance of tumor from closest distal margin
C4265604|T201|COMP|81182-8|LNC|Distance of tumor from closest proximal margin|Distance of tumor from closest proximal margin
C4265605|T201|COMP|81181-0|LNC|Serosal surface involvement|Serosal surface involvement
C4265606|T201|COMP|81180-2|LNC|Growth pattern|Growth pattern
C4265607|T201|COMP|81179-4|LNC|Histologic type|Histologic type
C4265608|T201|COMP|81178-6|LNC|Tissue block description and site|Tissue block description and site
C4265609|T201|COMP|81177-8|LNC|Serosal classification|Serosal classification
C4265611|T201|COMP|81175-2|LNC|Distance of tumor from closest margin|Distance of tumor from closest margin
C4265612|T201|COMP|81174-5|LNC|Tumor type|Tumor type
C4265613|T201|COMP|81173-7|LNC|Duodenum length|Duodenum length
C4265614|T201|COMP|81172-9|LNC|Esophagus length|Esophagus length
C4265615|T201|COMP|81171-1|LNC|Stomach.lesser curvature|Stomach.lesser curvature
C4265616|T201|COMP|81170-3|LNC|Stomach.greater curvature|Stomach.greater curvature
C4265629|T201|COMP|81157-0|LNC|Ubiquinone 10.reduced|Ubiquinone 10.reduced
C4265630|T201|COMP|81156-2|LNC|Ubiquinone 10.reduced/Ubiquinone 10|Ubiquinone 10.reduced/Ubiquinone 10
C4265631|T201|COMP|81155-4|LNC|Islet cell 512 Ab|Islet cell 512 Ab
C4265632|T201|COMP|81154-7|LNC|Dengue & Chikungunya & Zika virus panel|Dengue & Chikungunya & Zika virus panel
C4265635|T201|COMP|81151-3|LNC|Dengue virus 1+2+3+4 5' UTR RNA|Dengue virus 1+2+3+4 5' UTR RNA
C4265636|T201|COMP|81150-5|LNC|Dengue virus 1+2+3+4 5' UTR RNA|Dengue virus 1+2+3+4 5' UTR RNA
C4265637|T201|COMP|81149-7|LNC|Zika virus envelope (E) gene|Zika virus envelope (E) gene
C4265638|T201|COMP|81148-9|LNC|Zika virus envelope (E) gene|Zika virus envelope (E) gene
C4265639|T201|COMP|81147-1|LNC|Specimen source identification|Specimen source identification
C4265640|T201|COMP|81146-3|LNC|CYP3A4 & CYP3A5 gene targeted mutation analysis|CYP3A4 & CYP3A5 gene targeted mutation analysis
C4265641|T201|COMP|81144-8|LNC|Cerium|Cerium
C4265642|T201|COMP|81143-0|LNC|Galactokinase|Galactokinase
C4265643|T201|COMP|81142-2|LNC|PTPN22 gene.c.1858C>T|PTPN22 gene.c.1858C>T
C4265644|T201|COMP|81141-4|LNC|Spermatozoa motility|Spermatozoa motility
C4265645|T201|COMP|81140-6|LNC|CYP3A5 gene targeted mutation analysis|CYP3A5 gene targeted mutation analysis
C4265646|T201|COMP|81138-0|LNC|Spermatozoa.aggregated|Spermatozoa.aggregated
C4265654|T201|COMP|81125-7|LNC|Platelet aggregation.ristocetin inhibitor|Platelet aggregation.ristocetin inhibitor
C4265655|T201|COMP|81124-0|LNC|Coagulation factor V inhibitor|Coagulation factor V inhibitor
C4265656|T201|COMP|81123-2|LNC|Coagulation factor VII inhibitor|Coagulation factor VII inhibitor
C4265657|T201|COMP|81122-4|LNC|HIV 1 RNA reverse transcriptase & protease gene|HIV 1 RNA reverse transcriptase & protease gene
C4265658|T201|COMP|81121-6|LNC|Murray Valley encephalitis virus Ab|Murray Valley encephalitis virus Ab
C4265659|T201|COMP|81120-8|LNC|Barmah forest virus Ab|Barmah forest virus Ab
C4265660|T201|COMP|81119-0|LNC|Epstein Barr virus capsid Ab.IgG avidity|Epstein Barr virus capsid Ab.IgG avidity
C4265661|T201|COMP|81118-2|LNC|Legionella sp Ab.IgM|Legionella sp Ab.IgM
C4265662|T201|COMP|81117-4|LNC|Ross river virus RNA|Ross river virus RNA
C4265663|T201|COMP|81116-6|LNC|Hepatitis C virus core Ab+Ag|Hepatitis C virus core Ab+Ag
C4265664|T201|COMP|81115-8|LNC|Murray Valley encephalitis virus Ab|Murray Valley encephalitis virus Ab
C4265665|T201|COMP|81114-1|LNC|Murray Valley encephalitis virus Ab.IgM|Murray Valley encephalitis virus Ab.IgM
C4265666|T201|COMP|81113-3|LNC|Murray Valley encephalitis virus Ab.IgM|Murray Valley encephalitis virus Ab.IgM
C4265667|T201|COMP|81112-5|LNC|Murray Valley encephalitis virus Ab.IgG|Murray Valley encephalitis virus Ab.IgG
C4265668|T201|COMP|81111-7|LNC|Murray Valley encephalitis virus Ab.IgG|Murray Valley encephalitis virus Ab.IgG
C4265669|T201|COMP|81110-9|LNC|Leptospira weilii serovar Topaz Ab|Leptospira weilii serovar Topaz Ab
C4265670|T201|COMP|81109-1|LNC|Leptospira interrogans serovar Zanoni Ab|Leptospira interrogans serovar Zanoni Ab
C4265671|T201|COMP|81108-3|LNC|Leptospira interrogans serovar Szwajizak Ab|Leptospira interrogans serovar Szwajizak Ab
C4265672|T201|COMP|81107-5|LNC|Leptospira interrogans serovar Shermani Ab|Leptospira interrogans serovar Shermani Ab
C4265673|T201|COMP|81106-7|LNC|Leptospira interrogans serovar Robinsoni Ab|Leptospira interrogans serovar Robinsoni Ab
C4265674|T201|COMP|81105-9|LNC|Leptospira interrogans serovar Panama Ab|Leptospira interrogans serovar Panama Ab
C4265675|T201|COMP|81104-2|LNC|Leptospira interrogans serovar Medanensis Ab|Leptospira interrogans serovar Medanensis Ab
C4265676|T201|COMP|81103-4|LNC|Leptospira interrogans serovar Kremastos Ab|Leptospira interrogans serovar Kremastos Ab
C4265677|T201|COMP|81102-6|LNC|Leptospira interrogans serovar Cynopteri Ab|Leptospira interrogans serovar Cynopteri Ab
C4265678|T201|COMP|81101-8|LNC|Leptospira interrogans serovar Copenhageni Ab|Leptospira interrogans serovar Copenhageni Ab
C4265679|T201|COMP|81100-0|LNC|Leptospira interrogans serovar Celledoni Ab|Leptospira interrogans serovar Celledoni Ab
C4265680|T201|COMP|81099-4|LNC|Leptospira interrogans serovar Bulgarica Ab|Leptospira interrogans serovar Bulgarica Ab
C4265681|T201|COMP|81098-6|LNC|Leptospira borgpetersenii serovar Arborea Ab|Leptospira borgpetersenii serovar Arborea Ab
C4265682|T201|COMP|81097-8|LNC|West Nile virus Kunjin strain Ab|West Nile virus Kunjin strain Ab
C4265683|T201|COMP|81096-0|LNC|West Nile virus Kunjin strain Ab.IgM|West Nile virus Kunjin strain Ab.IgM
C4265776|T201|COMP|80982-2|LNC|Phytanoyl CoA hydroxlase|Phytanoyl CoA hydroxlase
C4265777|T201|COMP|80981-4|LNC|N,N-dimethylarginine|N,N-dimethylarginine
C4265778|T201|COMP|80980-6|LNC|Frataxin|Frataxin
C4265779|T201|COMP|80979-8|LNC|Frataxin|Frataxin
C4265784|T201|COMP|80974-9|LNC|Sulfamethoxazole.free|Sulfamethoxazole.free
C4265785|T201|COMP|80973-1|LNC|Trimethoprim.free|Trimethoprim.free
C4265786|T201|COMP|80972-3|LNC|Amikacin.free|Amikacin.free
C4265787|T201|COMP|80971-5|LNC|Gentamicin.free|Gentamicin.free
C4265788|T201|COMP|80970-7|LNC|Lithium.free|Lithium.free
C4265789|T201|COMP|80969-9|LNC|Methotrexate.free|Methotrexate.free
C4265790|T201|COMP|80968-1|LNC|Teicoplanin.free|Teicoplanin.free
C4265791|T201|COMP|80967-3|LNC|Theophylline.free|Theophylline.free
C4265792|T201|COMP|80966-5|LNC|Tobramycin.free|Tobramycin.free
C4265793|T201|COMP|80965-7|LNC|Topiramate.free|Topiramate.free
C4265794|T201|COMP|80964-0|LNC|Acetaminophen.free|Acetaminophen.free
C4265795|T201|COMP|80963-2|LNC|Salicylates.free|Salicylates.free
C4265796|T201|COMP|80962-4|LNC|ceFAZolin.free|ceFAZolin.free
C4265797|T201|COMP|80961-6|LNC|Cefotaxime.free|Cefotaxime.free
C4265798|T201|COMP|80960-8|LNC|cefTAZidime.free|cefTAZidime.free
C4265799|T201|COMP|80959-0|LNC|Glucose^1.5H post meal|Glucose^1.5H post meal
C4265800|T201|COMP|80958-2|LNC|Fractional excretion of magnesium|Fractional excretion of magnesium
C4265801|T201|COMP|80957-4|LNC|cefTRIAXone.free|cefTRIAXone.free
C4265835|T201|COMP|80912-9|LNC|Gadolinium|Gadolinium
C4265842|T201|COMP|80892-3|LNC|Heparin.unfractionated|Heparin.unfractionated
C4265899|T201|COMP|80832-9|LNC|Protein|Protein
C4265900|T201|COMP|80831-1|LNC|Pepsin A Panel|Pepsin A Panel
C4265902|T201|COMP|80829-5|LNC|Pepsin A+Pepsinogen A|Pepsin A+Pepsinogen A
C4265903|T201|COMP|80828-7|LNC|Pepsin A+Pepsinogen A|Pepsin A+Pepsinogen A
C4265905|T201|COMP|80826-1|LNC|Zika virus envelope (E) gene|Zika virus envelope (E) gene
C4265906|T201|COMP|80825-3|LNC|Zika virus envelope (E) gene|Zika virus envelope (E) gene
C4265907|T201|COMP|80824-6|LNC|Zika virus Ab.IgM|Zika virus Ab.IgM
C4265908|T201|COMP|80822-0|LNC|Zika virus Ab.Neut|Zika virus Ab.Neut
C4265909|T201|COMP|80821-2|LNC|Zika virus Ab.Neut|Zika virus Ab.Neut
C4265987|T201|COMP|80738-8|LNC|TPMT gene targeted mutation analysis|TPMT gene targeted mutation analysis
C4265988|T201|COMP|80737-0|LNC|Calculated panel reactive antibody|Calculated panel reactive antibody
C4265999|T201|COMP|80725-5|LNC|Trichomonas sp|Trichomonas sp
C4266000|T201|COMP|80724-8|LNC|Non-liquefied volume/Volume.total|Non-liquefied volume/Volume.total
C4266001|T201|COMP|80723-0|LNC|B-cell CD27 & IgD subsets|B-cell CD27 & IgD subsets
C4266007|T201|COMP|80717-2|LNC|B-cell CD27 & IgD subsets panel|B-cell CD27 & IgD subsets panel
C4266008|T201|COMP|80716-4|LNC|T-cell activated (CD38+HLA-DR+) subsets panel|T-cell activated (CD38+HLA-DR+) subsets panel
C4266009|T201|COMP|80715-6|LNC|FSHR gene targeted mutation analysis|FSHR gene targeted mutation analysis
C4266010|T201|COMP|80714-9|LNC|Cells.TCR gamma delta/100 Cells.CD3|Cells.TCR gamma delta/100 Cells.CD3
C4266011|T201|COMP|80713-1|LNC|Cells.TCR alpha beta/100 Cells.CD3|Cells.TCR alpha beta/100 Cells.CD3
C4266012|T201|COMP|80712-3|LNC|Cells.CD38+HLA-DR+/100 Cells.CD3+CD8+|Cells.CD38+HLA-DR+/100 Cells.CD3+CD8+
C4266013|T201|COMP|80711-5|LNC|Cells.CD38+HLA-DR+/100 Cells.CD3+CD4+|Cells.CD38+HLA-DR+/100 Cells.CD3+CD4+
C4266014|T201|COMP|80710-7|LNC|Cells.CD27-IgD+/100 Cells.CD19+CD20+|Cells.CD27-IgD+/100 Cells.CD19+CD20+
C4266015|T201|COMP|80709-9|LNC|Cells.CD27-CD45RA+/100 Cells.CD3+CD4+|Cells.CD27-CD45RA+/100 Cells.CD3+CD4+
C4266016|T201|COMP|80708-1|LNC|Cells.CD27-CD45RA-/100 Cells.CD3+CD4+|Cells.CD27-CD45RA-/100 Cells.CD3+CD4+
C4266017|T201|COMP|80707-3|LNC|Cells.CD27+IgD+/100 Cells.CD19+CD20+|Cells.CD27+IgD+/100 Cells.CD19+CD20+
C4266018|T201|COMP|80706-5|LNC|Cells.CD27+IgD-/100 Cells.CD19+CD20+|Cells.CD27+IgD-/100 Cells.CD19+CD20+
C4266019|T201|COMP|80705-7|LNC|Cells.CD27+CD45RA+/100 Cells.CD3+CD8+|Cells.CD27+CD45RA+/100 Cells.CD3+CD8+
C4266020|T201|COMP|80704-0|LNC|Cells.CD27+CD45RA+/100 Cells.CD3+CD4+|Cells.CD27+CD45RA+/100 Cells.CD3+CD4+
C4266021|T201|COMP|80703-2|LNC|Cells.CD27+CD45RA-/100 Cells.CD3+CD8+|Cells.CD27+CD45RA-/100 Cells.CD3+CD8+
C4266022|T201|COMP|80702-4|LNC|Cells.CD27+CD45RA-/100 Cells.CD3+CD4+|Cells.CD27+CD45RA-/100 Cells.CD3+CD4+
C4266023|T201|COMP|80701-6|LNC|Cells.CD27-/100 Cells.CD3+CD8+|Cells.CD27-/100 Cells.CD3+CD8+
C4266024|T201|COMP|80700-8|LNC|Cells.CD25+CD127-/100 cells.CD3+CD4+|Cells.CD25+CD127-/100 cells.CD3+CD4+
C4266025|T201|COMP|80699-2|LNC|Cells.CD4-CD8-/100 Cells.CD3+TCR alpha beta+|Cells.CD4-CD8-/100 Cells.CD3+TCR alpha beta+
C4266026|T201|COMP|80698-4|LNC|Viable CD34 cells/100 cells.CD34|Viable CD34 cells/100 cells.CD34
C4266027|T201|COMP|80697-6|LNC|Mycophenolate acyl-glucuronide|Mycophenolate acyl-glucuronide
C4266028|T201|COMP|80696-8|LNC|2-Chlorovinyl arsonous acid|2-Chlorovinyl arsonous acid
C4266029|T201|COMP|80695-0|LNC|HIV 1 proviral DNA genotype|HIV 1 proviral DNA genotype
C4266030|T201|COMP|80694-3|LNC|HIV 1 proviral DNA genotype|HIV 1 proviral DNA genotype
C4266033|T201|COMP|80684-4|LNC|Campylobacter coli+jejuni+lari 16S rRNA|Campylobacter coli+jejuni+lari 16S rRNA
C4266034|T201|COMP|80683-6|LNC|Giardia lamblia 18S rRNA|Giardia lamblia 18S rRNA
C4266035|T201|COMP|80682-8|LNC|Entamoeba histolytica 18S rRNA|Entamoeba histolytica 18S rRNA
C4266037|T201|COMP|80680-2|LNC|Vibrio cholerae toxin ctxA gene|Vibrio cholerae toxin ctxA gene
C4266038|T201|COMP|80679-4|LNC|Escherichia coli Stx1+Stx2 toxin stx1+stx2 genes|Escherichia coli Stx1+Stx2 toxin stx1+stx2 genes
C4266039|T201|COMP|80678-6|LNC|Salmonella sp invA+fliC genes|Salmonella sp invA+fliC genes
C4266040|T201|COMP|80677-8|LNC|Escherichia coli enterotoxigenic eltA+estB genes|Escherichia coli enterotoxigenic eltA+estB genes
C4266041|T201|COMP|80676-0|LNC|Escherichia coli O157 rfbE gene|Escherichia coli O157 rfbE gene
C4266042|T201|COMP|80675-2|LNC|Rotavirus A VP6 gene|Rotavirus A VP6 gene
C4266043|T201|COMP|80674-5|LNC|Adenovirus 40+41 fiber protein gene|Adenovirus 40+41 fiber protein gene
C4266054|T201|COMP|80663-8|LNC|4-Hydroxy 3-Nitrophenylacetate|4-Hydroxy 3-Nitrophenylacetate
C4266055|T201|COMP|80658-8|LNC|Activated clotting time|Activated clotting time
C4266056|T201|COMP|80657-0|LNC|Hemoglobin Q/Hemoglobin.total|Hemoglobin Q/Hemoglobin.total
C4266057|T201|COMP|80656-2|LNC|Hemoglobin Hope/Hemoglobin.total|Hemoglobin Hope/Hemoglobin.total
C4266058|T201|COMP|80655-4|LNC|Hemoglobin G-Philadelphia/Hemoglobin.total|Hemoglobin G-Philadelphia/Hemoglobin.total
C4266059|T201|COMP|80654-7|LNC|Spermatozoa.progressive.grade 1+2/100 spermatozoa|Spermatozoa.progressive.grade 1+2/100 spermatozoa
C4266060|T201|COMP|80653-9|LNC|Spermatozoa.normal chromatin/100 spermatozoa|Spermatozoa.normal chromatin/100 spermatozoa
C4266061|T201|COMP|80652-1|LNC|Everolimus|Everolimus
C4266062|T201|COMP|80651-3|LNC|Voriconazole N-oxide|Voriconazole N-oxide
C4266063|T201|COMP|80650-5|LNC|Tin|Tin
C4266064|T201|COMP|80649-7|LNC|Tetramethylenedisulfotetramine|Tetramethylenedisulfotetramine
C4266065|T201|COMP|80648-9|LNC|N-monodesmethyl bedaquiline|N-monodesmethyl bedaquiline
C4266066|T201|COMP|80647-1|LNC|Monoethyl methylphosphonate|Monoethyl methylphosphonate
C4266067|T201|COMP|80646-3|LNC|Monocyclohexyl methylphosphonate|Monocyclohexyl methylphosphonate
C4266068|T201|COMP|80645-5|LNC|Maprotiline+Normaprotiline|Maprotiline+Normaprotiline
C4266069|T201|COMP|80644-8|LNC|Isopropyl methylphosphonate|Isopropyl methylphosphonate
C4266070|T201|COMP|80643-0|LNC|Gadolinium|Gadolinium
C4266071|T201|COMP|80642-2|LNC|Floxacillin.free|Floxacillin.free
C4266072|T201|COMP|80641-4|LNC|Dothiepin+nordothiepin|Dothiepin+nordothiepin
C4266073|T201|COMP|80640-6|LNC|Disopyramide+Nordisopyramide|Disopyramide+Nordisopyramide
C4266074|T201|COMP|80639-8|LNC|Gamma-amanitin|Gamma-amanitin
C4266075|T201|COMP|80638-0|LNC|Beta-amanitin|Beta-amanitin
C4266076|T201|COMP|80637-2|LNC|Bedaquiline|Bedaquiline
C4266077|T201|COMP|80635-6|LNC|Aldicarb sulfoxide|Aldicarb sulfoxide
C4266078|T201|COMP|80634-9|LNC|Aldicarb sulfone|Aldicarb sulfone
C4266079|T201|COMP|80633-1|LNC|Aldicarb|Aldicarb
C4266080|T201|COMP|80632-3|LNC|2-Methylpropyl methylphosphonate|2-Methylpropyl methylphosphonate
C4266081|T201|COMP|80631-5|LNC|1,3-Dimethylbenzene+1,4-Dimethylbenzene|1,3-Dimethylbenzene+1,4-Dimethylbenzene
C4266082|T201|COMP|80630-7|LNC|1,2-Dichloroethane|1,2-Dichloroethane
C4266083|T201|COMP|80629-9|LNC|1,2,2-Trimethylpropyl methylphosphonate|1,2,2-Trimethylpropyl methylphosphonate
C4266084|T201|COMP|80628-1|LNC|1,1'-Sulfonylbis-2-Methylthioethane|1,1'-Sulfonylbis-2-Methylthioethane
C4266085|T201|COMP|80627-3|LNC|Coagulation factor X activated inhibitor|Coagulation factor X activated inhibitor
C4266087|T201|COMP|80625-7|LNC|Zika virus Ab.Neut^2nd specimen|Zika virus Ab.Neut^2nd specimen
C4266088|T201|COMP|80624-0|LNC|Zika virus Ab.Neut^1st specimen|Zika virus Ab.Neut^1st specimen
C4266089|T201|COMP|80623-2|LNC|Zika virus Ab.Neut^2nd specimen|Zika virus Ab.Neut^2nd specimen
C4266090|T201|COMP|80622-4|LNC|Zika virus Ab.Neut^1st specimen|Zika virus Ab.Neut^1st specimen
C4266091|T201|COMP|80621-6|LNC|Zika virus Ab.Neut|Zika virus Ab.Neut
C4266092|T201|COMP|80620-8|LNC|Zika virus Ab.Neut|Zika virus Ab.Neut
C4266093|T201|COMP|80619-0|LNC|Zika virus Ab.IgM|Zika virus Ab.IgM
C4266094|T201|COMP|80618-2|LNC|Zika virus Ab.IgM|Zika virus Ab.IgM
C4266095|T201|COMP|80617-4|LNC|Cefuroxime.free|Cefuroxime.free
C4266098|T201|COMP|80614-1|LNC|Baclofen|Baclofen
C4266099|T201|COMP|80613-3|LNC|Bicarbonate|Bicarbonate
C4266100|T201|COMP|80612-5|LNC|B Ab.IgG|B Ab.IgG
C4266101|T201|COMP|80611-7|LNC|Phosphate|Phosphate
C4266102|T201|COMP|80610-9|LNC|A Ab.IgG|A Ab.IgG
C4266103|T201|COMP|80609-1|LNC|Linezolid|Linezolid
C4266104|T201|COMP|80608-3|LNC|Cefuroxime|Cefuroxime
C4266105|T201|COMP|80607-5|LNC|14-Hydroxyclarithromycin|14-Hydroxyclarithromycin
C4266106|T201|COMP|80606-7|LNC|14-Hydroxyclarithromycin|14-Hydroxyclarithromycin
C4266107|T201|COMP|80605-9|LNC|Desacetylrifampicin|Desacetylrifampicin
C4266108|T201|COMP|80604-2|LNC|Desacetylrifampicin|Desacetylrifampicin
C4266109|T201|COMP|80603-4|LNC|Coagulation factor XI inhibitor|Coagulation factor XI inhibitor
C4266110|T201|COMP|80602-6|LNC|Respiratory pathogens identified|Respiratory pathogens identified
C4266113|T201|COMP|80599-4|LNC|Bordetella holmesii fumC gene|Bordetella holmesii fumC gene
C4266114|T201|COMP|80598-6|LNC|Respiratory syncytial virus B F gene|Respiratory syncytial virus B F gene
C4266115|T201|COMP|80597-8|LNC|Respiratory syncytial virus A 5' UTR RNA|Respiratory syncytial virus A 5' UTR RNA
C4266116|T201|COMP|80596-0|LNC|Rhinovirus 5' UTR RNA|Rhinovirus 5' UTR RNA
C4266117|T201|COMP|80595-2|LNC|Parainfluenza virus 4 P gene|Parainfluenza virus 4 P gene
C4266118|T201|COMP|80594-5|LNC|Parainfluenza virus 3 NP gene|Parainfluenza virus 3 NP gene
C4266119|T201|COMP|80593-7|LNC|Parainfluenza virus 2 L gene|Parainfluenza virus 2 L gene
C4266120|T201|COMP|80592-9|LNC|Parainfluenza virus 1 F gene|Parainfluenza virus 1 F gene
C4266121|T201|COMP|80591-1|LNC|Influenza virus B NS gene|Influenza virus B NS gene
C4266122|T201|COMP|80590-3|LNC|Influenza virus A H3 HA gene|Influenza virus A H3 HA gene
C4266123|T201|COMP|80589-5|LNC|Influenza virus A H1 HA gene|Influenza virus A H1 HA gene
C4266124|T201|COMP|80587-9|LNC|Human metapneumovirus A+B L+N genes|Human metapneumovirus A+B L+N genes
C4266125|T201|COMP|80586-1|LNC|Adenovirus hexon gene|Adenovirus hexon gene
C4266129|T201|COMP|80581-2|LNC|Incubation date & time range|Incubation date & time range
C4266140|T201|COMP|80561-4|LNC|cycloSPORINE|cycloSPORINE
C4266141|T201|COMP|80560-6|LNC|Citalopram|Citalopram
C4266142|T201|COMP|80559-8|LNC|Clarithromycin|Clarithromycin
C4266143|T201|COMP|80558-0|LNC|Amitriptyline|Amitriptyline
C4266144|T201|COMP|80557-2|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C4266145|T201|COMP|80556-4|LNC|cloZAPine|cloZAPine
C4266146|T201|COMP|80555-6|LNC|Diamorphine|Diamorphine
C4266147|T201|COMP|80554-9|LNC|Zopiclone|Zopiclone
C4266148|T201|COMP|80553-1|LNC|Voriconazole|Voriconazole
C4266149|T201|COMP|80552-3|LNC|Trimethoprim|Trimethoprim
C4266150|T201|COMP|80551-5|LNC|Tetrahydrocannabinol|Tetrahydrocannabinol
C4266151|T201|COMP|80550-7|LNC|Tacrolimus|Tacrolimus
C4266152|T201|COMP|80549-9|LNC|Sulfamethoxazole|Sulfamethoxazole
C4266153|T201|COMP|80548-1|LNC|Sirolimus|Sirolimus
C4266154|T201|COMP|80547-3|LNC|Rilpivirine|Rilpivirine
C4266155|T201|COMP|80546-5|LNC|rifAMPin|rifAMPin
C4266156|T201|COMP|80545-7|LNC|Posaconazole|Posaconazole
C4266157|T201|COMP|80544-0|LNC|Nortriptyline|Nortriptyline
C4266158|T201|COMP|80543-2|LNC|Norclozapine|Norclozapine
C4266159|T201|COMP|80542-4|LNC|Norcitalopram|Norcitalopram
C4266160|T201|COMP|80541-6|LNC|Nicotine|Nicotine
C4266161|T201|COMP|80540-8|LNC|Moxifloxacin|Moxifloxacin
C4266162|T201|COMP|80539-0|LNC|Morphine|Morphine
C4266163|T201|COMP|80538-2|LNC|Methylphenidate|Methylphenidate
C4266164|T201|COMP|80537-4|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C4266165|T201|COMP|80536-6|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C4266166|T201|COMP|80535-8|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C4266167|T201|COMP|80534-1|LNC|Methylenedioxyamphetamine|Methylenedioxyamphetamine
C4266168|T201|COMP|80533-3|LNC|Methamphetamine|Methamphetamine
C4266169|T201|COMP|80532-5|LNC|Methadone|Methadone
C4266170|T201|COMP|80531-7|LNC|Itraconazole|Itraconazole
C4266171|T201|COMP|80530-9|LNC|Fluconazole|Fluconazole
C4266172|T201|COMP|80529-1|LNC|Everolimus|Everolimus
C4266182|T201|COMP|80518-4|LNC|Clostridium baratii toxin F bont gene|Clostridium baratii toxin F bont gene
C4266184|T201|COMP|80516-8|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C4266185|T201|COMP|80515-0|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C4266205|T201|COMP|81246-1|LNC|HIV 2 RNA panel|HIV 2 RNA panel
C4266209|T201|COMP|81189-3|LNC|Tumor regression^post preoperative therapy|Tumor regression^post preoperative therapy
C4266211|T201|COMP|81187-7|LNC|Non-regional lymph nodes examined|Non-regional lymph nodes examined
C4266212|T201|COMP|81186-9|LNC|Cancer pathology panel|Cancer pathology panel
C4266222|T201|COMP|80662-0|LNC|Specimen volume|Specimen volume
C4266223|T201|COMP|80661-2|LNC|Color|Color
C4266224|T201|COMP|80660-4|LNC|Strongyloides sp Ab.IgG|Strongyloides sp Ab.IgG
C4266225|T201|COMP|80659-6|LNC|Activated clotting time|Activated clotting time
C4266226|T201|COMP|80376-7|LNC|Rotavirus & Adenovirus Ag panel|Rotavirus & Adenovirus Ag panel
C4266235|T201|COMP|80894-9|LNC|2-Methyltyrosine/Creatinine|2-Methyltyrosine/Creatinine
C4266254|T201|COMP|80690-1|LNC|HIV 1 proviral DNA tropism|HIV 1 proviral DNA tropism
C4266307|T201|COMP|69755-7|LNC|Bordetella pertussis.pertussis toxin Ab.IgG|Bordetella pertussis.pertussis toxin Ab.IgG
C4266310|T201|COMP|62324-9|LNC|Post-discharge provider name|Post-discharge provider name
C4283774|T201|COMP|82773-3|LNC|Lab result time reported|Lab result time reported
C4283776|T201|COMP|82955-6|LNC|HEDIS 2017 Value Sets|HEDIS 2017 Value Sets
C4283972|T201|COMP|82314-6|LNC|Specimen sent to CDC|Specimen sent to CDC
C4284219|T201|COMP|83006-7|LNC|Deletion-duplication overall interpretation|Deletion-duplication overall interpretation
C4284221|T201|COMP|83007-5|LNC|COSMIC version|COSMIC version
C4284333|T201|COMP|83005-9|LNC|Variant category|Variant category
C4284363|T201|COMP|82436-7|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C4284364|T201|COMP|82416-9|LNC|Histone Ab|Histone Ab
C4284365|T201|COMP|82428-4|LNC|Nucleosome Ab|Nucleosome Ab
C4284366|T201|COMP|82406-0|LNC|Ganglioside GM3 Ab.IgM|Ganglioside GM3 Ab.IgM
C4284384|T201|COMP|82959-8|LNC|HEDIS 2017-2020 Value Set - FOBT|HEDIS 2017-2020 Value Set - FOBT
C4284386|T201|COMP|82960-6|LNC|HEDIS 2017, 2018 Value Set - Group A Strep Tests|HEDIS 2017, 2018 Value Set - Group A Strep Tests
C4284540|T201|COMP|85093-3|LNC|Crystal casts|Crystal casts
C4284541|T201|COMP|85052-9|LNC|Ceftobiprole|Ceftobiprole
C4284543|T201|COMP|84924-0|LNC|Purkinje cell cytoplasmic type 1 Ab|Purkinje cell cytoplasmic type 1 Ab
C4284544|T201|COMP|84882-0|LNC|Histologic type|Histologic type
C4284663|T201|COMP|82446-6|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C4284664|T201|COMP|82429-2|LNC|Nucleosome Ab|Nucleosome Ab
C4284680|T201|COMP|84413-4|LNC|Genotype display name|Genotype display name
C4284722|T201|COMP|85069-3|LNC|Lab test method|Lab test method
C4284764|T201|COMP|82956-4|LNC|HEDIS 2017-2020 Value Set - FIT-DNA|HEDIS 2017-2020 Value Set - FIT-DNA
C4284771|T201|COMP|82962-2|LNC|HEDIS 2017, 2018 Value Set - Serum Potassium|HEDIS 2017, 2018 Value Set - Serum Potassium
C4284784|T201|COMP|82772-5|LNC|Lab result date reported|Lab result date reported
C4284786|T201|COMP|82785-7|LNC|Lab order date|Lab order date
C4284788|T201|COMP|84414-2|LNC|Haplotype name|Haplotype name
C4284868|T201|COMP|83140-4|LNC|17-Hydroxypregnenetriol|17-Hydroxypregnenetriol
C4284869|T201|COMP|83132-1|LNC|Pregnanolone|Pregnanolone
C4284870|T201|COMP|83094-3|LNC|Digoxin|Digoxin
C4284871|T201|COMP|83086-9|LNC|Choriogonadotropin|Choriogonadotropin
C4284929|T201|COMP|83008-3|LNC|ClinVar version|ClinVar version
C4284971|T201|COMP|85147-7|LNC|Programmed cell death ligand 1 by clone 22C3|Programmed cell death ligand 1 by clone 22C3
C4284974|T201|COMP|84928-1|LNC|N-methyl-D-aspartate receptor subunit 1 Ab|N-methyl-D-aspartate receptor subunit 1 Ab
C4284975|T201|COMP|84886-1|LNC|Satellite nodules|Satellite nodules
C4285014|T201|COMP|83120-6|LNC|Thyroxine|Thyroxine
C4285017|T201|COMP|83078-6|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C4285021|T201|COMP|82996-0|LNC|Mi-2 beta Ab.IgG|Mi-2 beta Ab.IgG
C4285022|T201|COMP|82988-7|LNC|N-methyl-D-aspartate receptor Ab.IgG|N-methyl-D-aspartate receptor Ab.IgG
C4285024|T201|COMP|82935-8|LNC|Oxazepam^trough|Oxazepam^trough
C4285025|T201|COMP|82924-2|LNC|Pl-7 Ab.IgG|Pl-7 Ab.IgG
C4285026|T201|COMP|82915-0|LNC|Fibrillarin Ab.IgG|Fibrillarin Ab.IgG
C4285027|T201|COMP|82885-5|LNC|Meta methylhippurate|Meta methylhippurate
C4285028|T201|COMP|82877-2|LNC|Cytochrome C oxidase|Cytochrome C oxidase
C4285034|T201|COMP|82730-3|LNC|GlycA|GlycA
C4285035|T201|COMP|82719-6|LNC|Enfuvirtide|Enfuvirtide
C4285045|T201|COMP|82576-0|LNC|Cyclic citrullinated peptide Ab.IgA|Cyclic citrullinated peptide Ab.IgA
C4285181|T201|COMP|85085-9|LNC|Nuclear Ab.IgG pattern.centrosomal|Nuclear Ab.IgG pattern.centrosomal
C4285183|T201|COMP|84904-2|LNC|Gleason score at positive margin|Gleason score at positive margin
C4285196|T201|COMP|82526-5|LNC|6-Beta naltrexol|6-Beta naltrexol
C4285197|T201|COMP|82518-2|LNC|IVD gene targeted mutation analysis|IVD gene targeted mutation analysis
C4285199|T201|COMP|82505-9|LNC|3-Hydroxyglutarate|3-Hydroxyglutarate
C4285200|T201|COMP|82497-9|LNC|TRBV6 gene segments/TRBV gene segments.total|TRBV6 gene segments/TRBV gene segments.total
C4285201|T201|COMP|82489-6|LNC|TRBV15 gene segments/TRBV gene segments.total|TRBV15 gene segments/TRBV gene segments.total
C4285203|T201|COMP|82452-4|LNC|U1 small nuclear ribonucleoprotein C Ab|U1 small nuclear ribonucleoprotein C Ab
C4285204|T201|COMP|82442-5|LNC|SUMO-activating enzyme subunit 2 Ab|SUMO-activating enzyme subunit 2 Ab
C4285205|T201|COMP|82394-8|LNC|Fibrillarin Ab|Fibrillarin Ab
C4285207|T201|COMP|82373-2|LNC|Buprenorphine|Buprenorphine
C4285209|T201|COMP|82302-1|LNC|Campylobacter sp|Campylobacter sp
C4285211|T201|COMP|82382-3|LNC|Sofosbuvir|Sofosbuvir
C4285212|T201|COMP|80375-9|LNC|Norovirus Ag|Norovirus Ag
C4285254|T201|COMP|85101-4|LNC|BRAF gene.p.Val600Glu|BRAF gene.p.Val600Glu
C4285256|T201|COMP|85051-1|LNC|Telavancin|Telavancin
C4285257|T201|COMP|84931-5|LNC|Gamma aminobutyrate B receptor Ab|Gamma aminobutyrate B receptor Ab
C4285258|T201|COMP|84894-5|LNC|Dimension|Dimension
C4285309|T201|COMP|84889-5|LNC|Extramural vein invasion|Extramural vein invasion
C4285397|T201|COMP|83125-5|LNC|Triiodothyronine|Triiodothyronine
C4285398|T201|COMP|83088-5|LNC|Cortisol|Cortisol
C4285399|T201|COMP|83081-0|LNC|Borrelia burgdorferi Ab.IgG+IgM|Borrelia burgdorferi Ab.IgG+IgM
C4285400|T201|COMP|83073-7|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C4285405|T201|COMP|82982-0|LNC|Exocrine pancreas Ab.IgA+IgG|Exocrine pancreas Ab.IgA+IgG
C4285406|T201|COMP|82974-7|LNC|O-nortramadol|O-nortramadol
C4285408|T201|COMP|82936-6|LNC|Signal recognition particle Ab.IgG|Signal recognition particle Ab.IgG
C4285409|T201|COMP|82925-9|LNC|PM-SCL-100 Ab.IgG|PM-SCL-100 Ab.IgG
C4285410|T201|COMP|82891-3|LNC|Para methylhippurate|Para methylhippurate
C4285435|T201|COMP|83111-5|LNC|Prolactin|Prolactin
C4285436|T201|COMP|83102-4|LNC|IgE|IgE
C4285437|T201|COMP|83060-4|LNC|NRAS gene|NRAS gene
C4285440|T201|COMP|82972-1|LNC|Butabarbital|Butabarbital
C4285441|T201|COMP|82964-8|LNC|Cannabidiol|Cannabidiol
C4285442|T201|COMP|82926-7|LNC|Phospholipase A2 receptor Ab.IgG|Phospholipase A2 receptor Ab.IgG
C4285443|T201|COMP|82917-6|LNC|Bromperidol^trough|Bromperidol^trough
C4285444|T201|COMP|82880-6|LNC|Escitalopram+norescitalopram|Escitalopram+norescitalopram
C4285445|T201|COMP|82872-3|LNC|A little n W little j Ab|A little n W little j Ab
C4285454|T201|COMP|83011-7|LNC|Haplotype definition panel|Haplotype definition panel
C4285488|T201|COMP|82884-8|LNC|MAOA gene.upstream VNTR repeats|MAOA gene.upstream VNTR repeats
C4285489|T201|COMP|82876-4|LNC|Complement C1 esterase inhibitor|Complement C1 esterase inhibitor
C4285503|T201|COMP|83071-1|LNC|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3
C4285504|T201|COMP|82600-8|LNC|Oncorhynchus keta roe Ab.IgE.RAST class|Oncorhynchus keta roe Ab.IgE.RAST class
C4285505|T201|COMP|82587-7|LNC|Leukocytes|Leukocytes
C4285508|T201|COMP|82541-4|LNC|Cetuximab Ab.IgE|Cetuximab Ab.IgE
C4285512|T201|COMP|82506-7|LNC|Oligosaccharides pattern|Oligosaccharides pattern
C4285513|T201|COMP|82475-5|LNC|Borrelia miyamotoi (glpQ) gene|Borrelia miyamotoi (glpQ) gene
C4285514|T201|COMP|82467-2|LNC|riTUXimab|riTUXimab
C4285515|T201|COMP|82459-9|LNC|Gadus chalcogrammus roe Ab.IgE.RAST class|Gadus chalcogrammus roe Ab.IgE.RAST class
C4285516|T201|COMP|82413-6|LNC|Ganglioside GT1a Ab.IgM|Ganglioside GT1a Ab.IgM
C4285521|T201|COMP|82780-8|LNC|Borrelia miyamotoi flaB gene|Borrelia miyamotoi flaB gene
C4285522|T201|COMP|82771-7|LNC|Lab test location performed|Lab test location performed
C4285530|T201|COMP|82602-4|LNC|Latex recombinant (rHev b) 10 Ab.IgE.RAST class|Latex recombinant (rHev b) 10 Ab.IgE.RAST class
C4285535|T201|COMP|82495-3|LNC|TRBV9 gene segments/TRBV gene segments.total|TRBV9 gene segments/TRBV gene segments.total
C4285536|T201|COMP|82486-2|LNC|TRBV19 gene segments/TRBV gene segments.total|TRBV19 gene segments/TRBV gene segments.total
C4285537|T201|COMP|82451-6|LNC|U1 small nuclear ribonucleoprotein A Ab|U1 small nuclear ribonucleoprotein A Ab
C4285538|T201|COMP|82441-7|LNC|SUMO-activating enzyme subunit 2 Ab|SUMO-activating enzyme subunit 2 Ab
C4285539|T201|COMP|82303-9|LNC|Escherichia coli O157|Escherichia coli O157
C4285540|T201|COMP|82866-5|LNC|Allo-pregnanediolone|Allo-pregnanediolone
C4285544|T201|COMP|82957-2|LNC|HEDIS 2017, 2018 Value Set - Chlamydia Tests|HEDIS 2017, 2018 Value Set - Chlamydia Tests
C4285566|T201|COMP|83137-0|LNC|OJ Ab.IgG|OJ Ab.IgG
C4285567|T201|COMP|83130-5|LNC|11-Deoxytetrahydrocorticosterone/Creatinine|11-Deoxytetrahydrocorticosterone/Creatinine
C4285568|T201|COMP|83092-7|LNC|Creatine kinase.MB|Creatine kinase.MB
C4285569|T201|COMP|83085-1|LNC|Carcinoembryonic Ag|Carcinoembryonic Ag
C4285570|T201|COMP|83077-8|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C4285573|T201|COMP|82994-5|LNC|MDA5 Ab.IgG|MDA5 Ab.IgG
C4285574|T201|COMP|82986-1|LNC|Contactin-associated protein 2 Ab.IgG|Contactin-associated protein 2 Ab.IgG
C4285575|T201|COMP|82978-8|LNC|Leucine-rich glioma-inactivated protein 1 Ab.IgG|Leucine-rich glioma-inactivated protein 1 Ab.IgG
C4285577|T201|COMP|82939-0|LNC|Genetic variant details|Genetic variant details
C4285578|T201|COMP|82931-7|LNC|Nuclear pore protein gp210 Ab.IgG|Nuclear pore protein gp210 Ab.IgG
C4285580|T201|COMP|82888-9|LNC|Ortho methylhippurate/Creatinine|Ortho methylhippurate/Creatinine
C4285583|T201|COMP|82399-7|LNC|Ganglioside GD2 Ab.IgG|Ganglioside GD2 Ab.IgG
C4285584|T201|COMP|82391-4|LNC|Centromere protein B Ab|Centromere protein B Ab
C4285587|T201|COMP|82335-1|LNC|Cytokines panel|Cytokines panel
C4285588|T201|COMP|82224-7|LNC|Ribose-5-phosphate isomerase|Ribose-5-phosphate isomerase
C4285589|T201|COMP|82216-3|LNC|3-Hydroxyisobutyrate dehydrogenase|3-Hydroxyisobutyrate dehydrogenase
C4285592|T201|COMP|82386-4|LNC|2-Methylcitrate|2-Methylcitrate
C4285614|T201|COMP|82738-6|LNC|DOPamine receptor D2 long Ab.IgG|DOPamine receptor D2 long Ab.IgG
C4285615|T201|COMP|82731-1|LNC|Zika virus Ab.IgM|Zika virus Ab.IgM
C4285624|T201|COMP|82603-2|LNC|Latex recombinant (rHev b) 2 Ab.IgE|Latex recombinant (rHev b) 2 Ab.IgE
C4285626|T201|COMP|82584-4|LNC|Dicarboxyhexenoylcarnitine (C6:1-DC)/Creatinine|Dicarboxyhexenoylcarnitine (C6:1-DC)/Creatinine
C4285629|T201|COMP|82538-0|LNC|CALR gene exon 9 full mutation analysis|CALR gene exon 9 full mutation analysis
C4285633|T201|COMP|82479-7|LNC|TRBV30 gene segment/TRBV gene segments.total|TRBV30 gene segment/TRBV gene segments.total
C4285634|T201|COMP|82472-2|LNC|Borrelia garinii+afzelii (oppA1) gene|Borrelia garinii+afzelii (oppA1) gene
C4285635|T201|COMP|82464-9|LNC|Mosquitoes tested|Mosquitoes tested
C4285636|T201|COMP|82422-7|LNC|Ks Ab|Ks Ab
C4285637|T201|COMP|82410-2|LNC|Ganglioside GQ1b Ab.IgG+IgM|Ganglioside GQ1b Ab.IgG+IgM
C4285638|T201|COMP|82396-3|LNC|Ganglioside GD1a Ab.IgG+IgM|Ganglioside GD1a Ab.IgG+IgM
C4285657|T201|COMP|82218-9|LNC|3-Methylcrotonyl-CoA carboxylase|3-Methylcrotonyl-CoA carboxylase
C4285659|T201|COMP|82383-1|LNC|Dengue virus 2+4 RNA|Dengue virus 2+4 RNA
C4285660|T201|COMP|80374-2|LNC|Adenovirus & Norovirus & Rotavirus Ag panel|Adenovirus & Norovirus & Rotavirus Ag panel
C4285662|T201|COMP|78433-0|LNC|Soluble liver Ab.IgG|Soluble liver Ab.IgG
C4297024|T201|COMP|83326-9|LNC|HIV 1 RNA genotype & phenotype|HIV 1 RNA genotype & phenotype
C4297025|T201|COMP|83056-2|LNC|Programmed cell death ligand 1 by clone 28-8|Programmed cell death ligand 1 by clone 28-8
C4297026|T201|COMP|82431-8|LNC|Platelet-derived growth factor receptor Ab|Platelet-derived growth factor receptor Ab
C4297028|T201|COMP|82225-4|LNC|Ribose-5-phosphate isomerase|Ribose-5-phosphate isomerase
C4297030|T201|COMP|85094-1|LNC|Escitalopram & norescitalopram panel|Escitalopram & norescitalopram panel
C4297034|T201|COMP|82723-8|LNC|Cocaine+Benzoylecgonine+Cocaethylene|Cocaine+Benzoylecgonine+Cocaethylene
C4297058|T201|COMP|85269-9|LNC|X-linked adrenoleukodystrophy|X-linked adrenoleukodystrophy
C4297134|T201|COMP|85149-3|LNC|Programmed cell death ligand 1 by clone SP142|Programmed cell death ligand 1 by clone SP142
C4297135|T201|COMP|85148-5|LNC|Programmed cell death ligand 1 by clone 28-8|Programmed cell death ligand 1 by clone 28-8
C4297138|T201|COMP|85100-6|LNC|FLT3 gene internal tandem duplication|FLT3 gene internal tandem duplication
C4297139|T201|COMP|85099-0|LNC|Norescitalopram|Norescitalopram
C4297140|T201|COMP|85098-2|LNC|Nitisinone|Nitisinone
C4297141|T201|COMP|85096-6|LNC|Myoglobin casts|Myoglobin casts
C4297142|T201|COMP|85095-8|LNC|D-3-phosphoglycerate dehydrogenase Ab.IgG|D-3-phosphoglycerate dehydrogenase Ab.IgG
C4297143|T201|COMP|85092-5|LNC|Autoimmune liver diseases Ab.IgG panel|Autoimmune liver diseases Ab.IgG panel
C4297144|T201|COMP|85091-7|LNC|HBA2 gene alpha 3.7kb triplication|HBA2 gene alpha 3.7kb triplication
C4297147|T201|COMP|85088-3|LNC|Maprotiline & normaprotiline panel|Maprotiline & normaprotiline panel
C4297148|T201|COMP|85087-5|LNC|Hexanoate|Hexanoate
C4297149|T201|COMP|85086-7|LNC|Elastase Ab.IgG|Elastase Ab.IgG
C4297150|T201|COMP|85084-2|LNC|Nuclear Ab.IgG pattern.coarse speckled|Nuclear Ab.IgG pattern.coarse speckled
C4297151|T201|COMP|85083-4|LNC|Nuclear Ab.IgG pattern.homogeneous|Nuclear Ab.IgG pattern.homogeneous
C4297152|T201|COMP|85082-6|LNC|Nuclear Ab.IgG pattern.nuclear membrane pores|Nuclear Ab.IgG pattern.nuclear membrane pores
C4297153|T201|COMP|85081-8|LNC|Nuclear Ab.IgG pattern.multiple nuclear dots|Nuclear Ab.IgG pattern.multiple nuclear dots
C4297154|T201|COMP|85080-0|LNC|Nuclear Ab.IgG pattern.nucleolar|Nuclear Ab.IgG pattern.nucleolar
C4297155|T201|COMP|85079-2|LNC|Nuclear Ab.IgG pattern.other|Nuclear Ab.IgG pattern.other
C4297157|T201|COMP|85068-5|LNC|Estradiol^post dose dexamethasone|Estradiol^post dose dexamethasone
C4297159|T201|COMP|85066-9|LNC|Estradiol^post dose lutropin|Estradiol^post dose lutropin
C4297160|T201|COMP|85065-1|LNC|Estradiol^post dose follitropin|Estradiol^post dose follitropin
C4297168|T201|COMP|85048-7|LNC|Micafungin|Micafungin
C4297173|T201|COMP|84927-3|LNC|Glial nuclear type 1 Ab|Glial nuclear type 1 Ab
C4297174|T201|COMP|84926-5|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C4297175|T201|COMP|84925-7|LNC|Purkinje cell cytoplasmic type 2 Ab|Purkinje cell cytoplasmic type 2 Ab
C4297176|T201|COMP|84923-2|LNC|Purkinje cell cytoplasmic type 1 Ab|Purkinje cell cytoplasmic type 1 Ab
C4297177|T201|COMP|84922-4|LNC|Cells.chromosome 7 monosomy/Cells counted|Cells.chromosome 7 monosomy/Cells counted
C4297181|T201|COMP|84913-3|LNC|Cells.chromosome 12 trisomy/Cells counted|Cells.chromosome 12 trisomy/Cells counted
C4297183|T201|COMP|84908-3|LNC|Cancer pathology panel|Cancer pathology panel
C4297184|T201|COMP|84907-5|LNC|Cancer pathology panel|Cancer pathology panel
C4297185|T201|COMP|84906-7|LNC|Bladder neck involvement|Bladder neck involvement
C4297186|T201|COMP|84905-9|LNC|Margin involvement|Margin involvement
C4297187|T201|COMP|84903-4|LNC|Extraprostatic extension extent|Extraprostatic extension extent
C4297188|T201|COMP|84902-6|LNC|Extraprostatic extension site|Extraprostatic extension site
C4297189|T201|COMP|84901-8|LNC|Other nodule plane|Other nodule plane
C4297190|T201|COMP|84900-0|LNC|Other nodule quadrant|Other nodule quadrant
C4297191|T201|COMP|84899-4|LNC|Other nodules greater than 10mm in diameter|Other nodules greater than 10mm in diameter
C4297192|T201|COMP|84898-6|LNC|Dominant nodule plane|Dominant nodule plane
C4297193|T201|COMP|84897-8|LNC|Dominant nodule quadrant|Dominant nodule quadrant
C4297194|T201|COMP|84896-0|LNC|Lymph node(s)|Lymph node(s)
C4297195|T201|COMP|84895-2|LNC|Seminal vesicles|Seminal vesicles
C4297197|T201|COMP|84892-9|LNC|Residual tumor classification|Residual tumor classification
C4297198|T201|COMP|84891-1|LNC|Response to neoadjuvant therapy|Response to neoadjuvant therapy
C4297199|T201|COMP|84885-3|LNC|Surgical margin tumor involvement.circumferential|Surgical margin tumor involvement.circumferential
C4297200|T201|COMP|84884-6|LNC|Distal &or proximal margin involvement|Distal &or proximal margin involvement
C4297201|T201|COMP|84883-8|LNC|Deepest extent of tumor invasion|Deepest extent of tumor invasion
C4297202|T201|COMP|84881-2|LNC|Polyps|Polyps
C4297204|T201|COMP|84879-6|LNC|Tumor perforation|Tumor perforation
C4297208|T201|COMP|84873-9|LNC|Myelin oligodendrocyte glycoprotein Ab.IgG|Myelin oligodendrocyte glycoprotein Ab.IgG
C4297209|T201|COMP|84872-1|LNC|Epstein Barr virus nuclear 1 Ab.IgG|Epstein Barr virus nuclear 1 Ab.IgG
C4297210|T201|COMP|84871-3|LNC|Epstein Barr virus capsid p18 Ab.IgG|Epstein Barr virus capsid p18 Ab.IgG
C4297283|T201|COMP|84919-0|LNC|Chromosome 21 aneuploidy|Chromosome 21 aneuploidy
C4297284|T201|COMP|84918-2|LNC|Chromosome X aneuploidy|Chromosome X aneuploidy
C4297285|T201|COMP|84917-4|LNC|Chromosome Y aneuploidy|Chromosome Y aneuploidy
C4297409|T201|COMP|85037-0|LNC|HIV 1 & 2 Ab & HIV 1 p24 Ag panel|HIV 1 & 2 Ab & HIV 1 p24 Ag panel
C4297428|T201|COMP|84890-3|LNC|Distant metastases confirmed by histology|Distant metastases confirmed by histology
C4297429|T201|COMP|84888-7|LNC|Intramural vein invasion|Intramural vein invasion
C4297430|T201|COMP|84887-9|LNC|Apical lymph node involvement|Apical lymph node involvement
C4298161|T201|COMP|83327-7|LNC|HIV 1 RNA phenotype|HIV 1 RNA phenotype
C4298162|T201|COMP|83325-1|LNC|HIV 1 RNA genotype|HIV 1 RNA genotype
C4298165|T201|COMP|83321-0|LNC|Pathology report.intraoperative observation|Pathology report.intraoperative observation
C4298211|T201|COMP|83139-6|LNC|17-Hydroxypregnenetriol/Creatinine|17-Hydroxypregnenetriol/Creatinine
C4298212|T201|COMP|83138-8|LNC|17-Hydroxypregnenetriol|17-Hydroxypregnenetriol
C4298213|T201|COMP|83136-2|LNC|Allo-pregnanediol/Creatinine|Allo-pregnanediol/Creatinine
C4298214|T201|COMP|83135-4|LNC|Allo-pregnanediolone/Creatinine|Allo-pregnanediolone/Creatinine
C4298215|T201|COMP|83133-9|LNC|Pregnanolone/Creatinine|Pregnanolone/Creatinine
C4298216|T201|COMP|83131-3|LNC|Pregnanolone|Pregnanolone
C4298217|T201|COMP|83127-1|LNC|Triiodothyronine.free|Triiodothyronine.free
C4298218|T201|COMP|83126-3|LNC|Triiodothyronine.free|Triiodothyronine.free
C4298219|T201|COMP|83124-8|LNC|Triiodothyronine|Triiodothyronine
C4298220|T201|COMP|83123-0|LNC|Toxoplasma gondii Ab.IgG+IgM|Toxoplasma gondii Ab.IgG+IgM
C4298221|T201|COMP|83122-2|LNC|Thyroxine.free|Thyroxine.free
C4298222|T201|COMP|83121-4|LNC|Thyroxine.free|Thyroxine.free
C4298223|T201|COMP|83119-8|LNC|Thyroxine|Thyroxine
C4298224|T201|COMP|83112-3|LNC|Prostate specific Ag|Prostate specific Ag
C4298225|T201|COMP|83110-7|LNC|Progesterone|Progesterone
C4298226|T201|COMP|83109-9|LNC|Progesterone|Progesterone
C4298227|T201|COMP|83108-1|LNC|Natriuretic peptide.B prohormone N-Terminal|Natriuretic peptide.B prohormone N-Terminal
C4298228|T201|COMP|83107-3|LNC|Natriuretic peptide.B prohormone N-Terminal|Natriuretic peptide.B prohormone N-Terminal
C4298229|T201|COMP|83106-5|LNC|Myoglobin|Myoglobin
C4298230|T201|COMP|83105-7|LNC|Mullerian inhibiting substance|Mullerian inhibiting substance
C4298231|T201|COMP|83104-0|LNC|Mullerian inhibiting substance|Mullerian inhibiting substance
C4298232|T201|COMP|83103-2|LNC|Lutropin|Lutropin
C4298233|T201|COMP|83101-6|LNC|HIV 1+2 Ab & HIV1 p24 Ag panel|HIV 1+2 Ab & HIV1 p24 Ag panel
C4298234|T201|COMP|83100-8|LNC|Hepatitis B virus core Ab.IgG+IgM|Hepatitis B virus core Ab.IgG+IgM
C4298235|T201|COMP|83099-2|LNC|Galectin 3|Galectin 3
C4298236|T201|COMP|83098-4|LNC|Follitropin|Follitropin
C4298237|T201|COMP|83097-6|LNC|Estradiol|Estradiol
C4298238|T201|COMP|83096-8|LNC|Estradiol|Estradiol
C4298239|T201|COMP|83095-0|LNC|Epstein Barr virus capsid+early Ab.IgG|Epstein Barr virus capsid+early Ab.IgG
C4298240|T201|COMP|83093-5|LNC|Digoxin|Digoxin
C4298241|T201|COMP|83091-9|LNC|Cortisol|Cortisol
C4298242|T201|COMP|83090-1|LNC|Cortisol|Cortisol
C4298243|T201|COMP|83089-3|LNC|Cortisol|Cortisol
C4298244|T201|COMP|83087-7|LNC|Clostridioides difficile glutamate dehydrogenase|Clostridioides difficile glutamate dehydrogenase
C4298245|T201|COMP|83084-4|LNC|Cancer Ag 19-9|Cancer Ag 19-9
C4298246|T201|COMP|83083-6|LNC|Cancer Ag 15-3|Cancer Ag 15-3
C4298247|T201|COMP|83082-8|LNC|Cancer Ag 125|Cancer Ag 125
C4298248|T201|COMP|83080-2|LNC|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C4298249|T201|COMP|83079-4|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C4298250|T201|COMP|83076-0|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C4298251|T201|COMP|83075-2|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C4298252|T201|COMP|83074-5|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C4298254|T201|COMP|83065-3|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C4298255|T201|COMP|83064-6|LNC|Calcium.ionized|Calcium.ionized
C4298256|T201|COMP|83063-8|LNC|PTEN gene|PTEN gene
C4298257|T201|COMP|83062-0|LNC|PIK3CA gene|PIK3CA gene
C4298258|T201|COMP|83061-2|LNC|BRAF gene|BRAF gene
C4298259|T201|COMP|83059-6|LNC|KRAS gene|KRAS gene
C4298260|T201|COMP|83058-8|LNC|Nucleoprotein expression|Nucleoprotein expression
C4298261|T201|COMP|83057-0|LNC|Programmed cell death ligand 1 by clone SP142|Programmed cell death ligand 1 by clone SP142
C4298266|T201|COMP|83118-0|LNC|Thyroperoxidase Ab.IgG|Thyroperoxidase Ab.IgG
C4298267|T201|COMP|83117-2|LNC|Thyroglobulin Ab.IgG|Thyroglobulin Ab.IgG
C4298268|T201|COMP|83116-4|LNC|Testosterone|Testosterone
C4298269|T201|COMP|83115-6|LNC|Testosterone|Testosterone
C4298270|T201|COMP|83113-1|LNC|Prostate specific Ag.free|Prostate specific Ag.free
C4298271|T201|COMP|83055-4|LNC|Programmed cell death ligand 1 by clone 28-8|Programmed cell death ligand 1 by clone 28-8
C4298272|T201|COMP|83054-7|LNC|Programmed cell death ligand 1 by clone 22C3|Programmed cell death ligand 1 by clone 22C3
C4298273|T201|COMP|83052-1|LNC|Programmed cell death ligand 1 by clone 22C3|Programmed cell death ligand 1 by clone 22C3
C4298293|T201|COMP|83010-9|LNC|Medication usage suggestion|Medication usage suggestion
C4298294|T201|COMP|83009-1|LNC|Genetic variation effect on high-risk allele|Genetic variation effect on high-risk allele
C4298295|T201|COMP|83004-2|LNC|Glutamate decarboxylase 65 Ab.IgG|Glutamate decarboxylase 65 Ab.IgG
C4298296|T201|COMP|83003-4|LNC|Recoverin Ab.IgG|Recoverin Ab.IgG
C4298297|T201|COMP|83002-6|LNC|Zinc finger protein of the cerebellum 4 Ab.IgG|Zinc finger protein of the cerebellum 4 Ab.IgG
C4298298|T201|COMP|83001-8|LNC|Glial nuclear type 1 Ab.IgG|Glial nuclear type 1 Ab.IgG
C4298299|T201|COMP|83000-0|LNC|Titin Ab.IgG|Titin Ab.IgG
C4298300|T201|COMP|82999-4|LNC|Purkinje cell cytoplasmic type Tr Ab.IgG|Purkinje cell cytoplasmic type Tr Ab.IgG
C4298301|T201|COMP|82998-6|LNC|Dense fine speckled 70 protein Ab.IgG|Dense fine speckled 70 protein Ab.IgG
C4298302|T201|COMP|82997-8|LNC|Mi-2 alpha Ab.IgG|Mi-2 alpha Ab.IgG
C4298303|T201|COMP|82995-2|LNC|TIF1-gamma Ab.IgG|TIF1-gamma Ab.IgG
C4298304|T201|COMP|82993-7|LNC|MJ Ab.IgG|MJ Ab.IgG
C4298305|T201|COMP|82992-9|LNC|SUMO-activating enzyme subunit 1 Ab.IgG|SUMO-activating enzyme subunit 1 Ab.IgG
C4298306|T201|COMP|82991-1|LNC|Phospholipase A2 receptor Ab.IgG|Phospholipase A2 receptor Ab.IgG
C4298307|T201|COMP|82989-5|LNC|Dipeptidyl aminopeptidase-like protein 6 Ab.IgG|Dipeptidyl aminopeptidase-like protein 6 Ab.IgG
C4298309|T201|COMP|82985-3|LNC|Leucine-rich glioma-inactivated protein 1 Ab.IgG|Leucine-rich glioma-inactivated protein 1 Ab.IgG
C4298310|T201|COMP|82984-6|LNC|Gamma aminobutyrate B receptor Ab.IgG|Gamma aminobutyrate B receptor Ab.IgG
C4298311|T201|COMP|82983-8|LNC|Ma+Ta Ab.IgG|Ma+Ta Ab.IgG
C4298312|T201|COMP|82981-2|LNC|N-methyl-D-aspartate receptor Ab.IgG|N-methyl-D-aspartate receptor Ab.IgG
C4298313|T201|COMP|82979-6|LNC|Contactin-associated protein 2 Ab.IgG|Contactin-associated protein 2 Ab.IgG
C4298314|T201|COMP|82977-0|LNC|Gamma aminobutyrate B receptor Ab.IgG|Gamma aminobutyrate B receptor Ab.IgG
C4298315|T201|COMP|82976-2|LNC|Dipeptidyl aminopeptidase-like protein 6 Ab.IgG|Dipeptidyl aminopeptidase-like protein 6 Ab.IgG
C4298316|T201|COMP|82975-4|LNC|Desmosome Ab.IgG|Desmosome Ab.IgG
C4298317|T201|COMP|82973-9|LNC|Amobarbital|Amobarbital
C4298318|T201|COMP|82971-3|LNC|Butalbital|Butalbital
C4298319|T201|COMP|82970-5|LNC|PHENobarbital|PHENobarbital
C4298320|T201|COMP|82969-7|LNC|PENTobarbital|PENTobarbital
C4298321|T201|COMP|82968-9|LNC|Secobarbital|Secobarbital
C4298322|T201|COMP|82967-1|LNC|Amphetamine|Amphetamine
C4298323|T201|COMP|82966-3|LNC|Methamphetamine|Methamphetamine
C4298324|T201|COMP|82965-5|LNC|Methylenedioxyethylamphetamine|Methylenedioxyethylamphetamine
C4298337|T201|COMP|82938-2|LNC|Smith extractable nuclear D Ab.IgG|Smith extractable nuclear D Ab.IgG
C4298339|T201|COMP|82934-1|LNC|clonazePAM^trough|clonazePAM^trough
C4298341|T201|COMP|82932-5|LNC|sp100 Ab.IgG|sp100 Ab.IgG
C4298342|T201|COMP|82928-3|LNC|Mitochondria M2 Ab.IgG|Mitochondria M2 Ab.IgG
C4298343|T201|COMP|82923-4|LNC|PML Ab.IgG|PML Ab.IgG
C4298344|T201|COMP|82921-8|LNC|Liver cytosol Ab.IgG|Liver cytosol Ab.IgG
C4298345|T201|COMP|82920-0|LNC|Legionella pneumophila Ab.IgA|Legionella pneumophila Ab.IgA
C4298346|T201|COMP|82919-2|LNC|Ku Ab.IgG|Ku Ab.IgG
C4298347|T201|COMP|82918-4|LNC|Jo-1 extractable nuclear Ab.IgG|Jo-1 extractable nuclear Ab.IgG
C4298348|T201|COMP|82916-8|LNC|Flurazepam^trough|Flurazepam^trough
C4298349|T201|COMP|82914-3|LNC|Dothiepin^trough|Dothiepin^trough
C4298350|T201|COMP|82913-5|LNC|Centromere protein B Ab.IgG|Centromere protein B Ab.IgG
C4298351|T201|COMP|82911-9|LNC|Vascular endothelial growth factor D|Vascular endothelial growth factor D
C4298352|T201|COMP|82910-1|LNC|Thromboxane beta 2|Thromboxane beta 2
C4298353|T201|COMP|82909-3|LNC|Tetrahydrocortisol/5-alpha tetrahydrocortisol|Tetrahydrocortisol/5-alpha tetrahydrocortisol
C4298354|T201|COMP|82908-5|LNC|Tetrahydrocortisol/5-alpha tetrahydrocortisol|Tetrahydrocortisol/5-alpha tetrahydrocortisol
C4298358|T201|COMP|82904-4|LNC|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript
C4298360|T201|COMP|82902-8|LNC|Somatotropin^15M pre XXX challenge|Somatotropin^15M pre XXX challenge
C4298368|T201|COMP|82893-9|LNC|Penfluridol|Penfluridol
C4298369|T201|COMP|82892-1|LNC|Para methylhippurate/Creatinine|Para methylhippurate/Creatinine
C4298372|T201|COMP|82887-1|LNC|Ortho methylhippurate|Ortho methylhippurate
C4298373|T201|COMP|82886-3|LNC|Meta methylhippurate/Creatinine|Meta methylhippurate/Creatinine
C4298374|T201|COMP|82883-0|LNC|Lysosomal acid lipase|Lysosomal acid lipase
C4298375|T201|COMP|82882-2|LNC|Etiocholanolone/Androsterone|Etiocholanolone/Androsterone
C4298376|T201|COMP|82881-4|LNC|Etiocholanolone/Androsterone|Etiocholanolone/Androsterone
C4298379|T201|COMP|82875-6|LNC|Campylobacter jejuni Ab.IgA|Campylobacter jejuni Ab.IgA
C4298380|T201|COMP|82874-9|LNC|Calprotectin|Calprotectin
C4298381|T201|COMP|82873-1|LNC|Brallobarbital|Brallobarbital
C4298382|T201|COMP|82871-5|LNC|Adenosine diphosphate|Adenosine diphosphate
C4298383|T201|COMP|82870-7|LNC|A little u super little b Ab|A little u super little b Ab
C4298387|T201|COMP|82860-8|LNC|11-Deoxytetrahydrocorticosterone|11-Deoxytetrahydrocorticosterone
C4298388|T201|COMP|82859-0|LNC|11-Deoxytetrahydrocorticosterone|11-Deoxytetrahydrocorticosterone
C4298389|T201|COMP|82858-2|LNC|11-Deoxytetrahydrocorticosterone|11-Deoxytetrahydrocorticosterone
C4298402|T201|COMP|82845-9|LNC|Campylobacter jejuni Ab.IgA & IgG & IgM panel|Campylobacter jejuni Ab.IgA & IgG & IgM panel
C4298404|T201|COMP|82842-6|LNC|Liver kidney microsomal Ab.IgG|Liver kidney microsomal Ab.IgG
C4298405|T201|COMP|82841-8|LNC|PCNA extractable nuclear Ab.IgG|PCNA extractable nuclear Ab.IgG
C4298406|T201|COMP|82840-0|LNC|Mitochondria Ab.IgG|Mitochondria Ab.IgG
C4298417|T201|COMP|82812-9|LNC|Sodium|Sodium
C4298427|T201|COMP|82799-8|LNC|Spatial clot growth analysis panel|Spatial clot growth analysis panel
C4298428|T201|COMP|82798-0|LNC|Clot formation lag time|Clot formation lag time
C4298429|T201|COMP|82797-2|LNC|Clot growth.initial|Clot growth.initial
C4298430|T201|COMP|82796-4|LNC|Clot growth.stationary|Clot growth.stationary
C4298431|T201|COMP|82795-6|LNC|Clot growth|Clot growth
C4298432|T201|COMP|82794-9|LNC|Clot formation.spontaneous|Clot formation.spontaneous
C4298433|T201|COMP|82793-1|LNC|Clot size^30M post incubation|Clot size^30M post incubation
C4298434|T201|COMP|82792-3|LNC|Clot density|Clot density
C4298436|T201|COMP|82781-6|LNC|Borrelia miyamotoi flaB gene|Borrelia miyamotoi flaB gene
C4298439|T201|COMP|82768-3|LNC|Lab order priority|Lab order priority
C4298447|T201|COMP|82748-5|LNC|Erythrocytes.Babesia sp infected/100 erythrocytes|Erythrocytes.Babesia sp infected/100 erythrocytes
C4298448|T201|COMP|82747-7|LNC|Babesia microti Ab.IgG|Babesia microti Ab.IgG
C4298449|T201|COMP|82746-9|LNC|Varicella zoster virus strain|Varicella zoster virus strain
C4298453|T201|COMP|82740-2|LNC|Lysoganglioside GM1 Ab.IgG|Lysoganglioside GM1 Ab.IgG
C4298454|T201|COMP|82739-4|LNC|DOPamine receptor D1 Ab.IgG|DOPamine receptor D1 Ab.IgG
C4298455|T201|COMP|82737-8|LNC|Beta tubulin Ab.IgG|Beta tubulin Ab.IgG
C4298461|T201|COMP|82722-0|LNC|Potassium|Potassium
C4298462|T201|COMP|82721-2|LNC|Intravenous lipid emulsion|Intravenous lipid emulsion
C4298463|T201|COMP|82720-4|LNC|Natural killer cell cytotoxicity panel|Natural killer cell cytotoxicity panel
C4298510|T201|COMP|82660-2|LNC|Glutamate decarboxylase Ab|Glutamate decarboxylase Ab
C4298511|T201|COMP|82659-4|LNC|Thyrotropin receptor Ab|Thyrotropin receptor Ab
C4298512|T201|COMP|82658-6|LNC|Glutamate decarboxylase Ab|Glutamate decarboxylase Ab
C4298569|T201|COMP|83072-9|LNC|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C4298570|T201|COMP|83070-3|LNC|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3
C4298571|T201|COMP|83069-5|LNC|Zika virus non-structural protein 1 Ab.IgG|Zika virus non-structural protein 1 Ab.IgG
C4298585|T201|COMP|82613-1|LNC|Apis mellifera recombinant (rApi m) 10 Ab.IgE|Apis mellifera recombinant (rApi m) 10 Ab.IgE
C4298591|T201|COMP|82604-0|LNC|Latex recombinant (rHev b) 2 Ab.IgE.RAST class|Latex recombinant (rHev b) 2 Ab.IgE.RAST class
C4298592|T201|COMP|82601-6|LNC|Latex recombinant (rHev b) 10 Ab.IgE|Latex recombinant (rHev b) 10 Ab.IgE
C4298593|T201|COMP|82599-2|LNC|Oncorhynchus keta roe Ab.IgE|Oncorhynchus keta roe Ab.IgE
C4298595|T201|COMP|82597-6|LNC|Chromosome painting analysis|Chromosome painting analysis
C4298599|T201|COMP|82588-5|LNC|Erythrocytes|Erythrocytes
C4298600|T201|COMP|82586-9|LNC|Nucleated cells|Nucleated cells
C4298601|T201|COMP|82585-1|LNC|Dicarboxyhexenoylcarnitine (C6:1-DC)|Dicarboxyhexenoylcarnitine (C6:1-DC)
C4298602|T201|COMP|82583-6|LNC|Triticum aestivum native (nTri a) 19+20+21 Ab.IgE|Triticum aestivum native (nTri a) 19+20+21 Ab.IgE
C4298608|T201|COMP|82575-2|LNC|Urobilinogen|Urobilinogen
C4298609|T201|COMP|82574-5|LNC|Staphylococcus aureus enterotoxin E Ab.IgE|Staphylococcus aureus enterotoxin E Ab.IgE
C4298611|T201|COMP|82572-9|LNC|Betula verrucosa recombinant (rBet v) 6 Ab.IgE|Betula verrucosa recombinant (rBet v) 6 Ab.IgE
C4298612|T201|COMP|82571-1|LNC|Coryphaena hippurus Ab.IgE.RAST class|Coryphaena hippurus Ab.IgE.RAST class
C4298613|T201|COMP|82570-3|LNC|Coryphaena hippurus Ab.IgE|Coryphaena hippurus Ab.IgE
C4298632|T201|COMP|82544-8|LNC|Dog recombinant (rCan f) 4 Ab.IgE.RAST class|Dog recombinant (rCan f) 4 Ab.IgE.RAST class
C4298633|T201|COMP|82543-0|LNC|Dog recombinant (rCan f) 4 Ab.IgE|Dog recombinant (rCan f) 4 Ab.IgE
C4298634|T201|COMP|82542-2|LNC|Cetuximab Ab.IgE.RAST class|Cetuximab Ab.IgE.RAST class
C4298637|T201|COMP|82537-2|LNC|RAF1 gene full mutation analysis|RAF1 gene full mutation analysis
C4298638|T201|COMP|82536-4|LNC|SOS1 gene full mutation analysis|SOS1 gene full mutation analysis
C4298639|T201|COMP|82535-6|LNC|KRAS gene full mutation analysis|KRAS gene full mutation analysis
C4298640|T201|COMP|82534-9|LNC|CASR gene full mutation analysis|CASR gene full mutation analysis
C4298641|T201|COMP|82527-3|LNC|6-Beta naltrexol/Creatinine|6-Beta naltrexol/Creatinine
C4298642|T201|COMP|82524-0|LNC|6-Beta naltrexol|6-Beta naltrexol
C4298643|T201|COMP|82523-2|LNC|Grazoprevir|Grazoprevir
C4298644|T201|COMP|82522-4|LNC|Simeprevir|Simeprevir
C4298645|T201|COMP|82521-6|LNC|Paritaprevir|Paritaprevir
C4298646|T201|COMP|82520-8|LNC|Velpatasvir|Velpatasvir
C4298647|T201|COMP|82519-0|LNC|Dengue virus 1+3 & 2+4 panel|Dengue virus 1+3 & 2+4 panel
C4298648|T201|COMP|82517-4|LNC|LAMA3 gene targeted mutation analysis|LAMA3 gene targeted mutation analysis
C4298649|T201|COMP|82516-6|LNC|LAMC2 gene targeted mutation analysis|LAMC2 gene targeted mutation analysis
C4298650|T201|COMP|82515-8|LNC|NBN gene targeted mutation analysis|NBN gene targeted mutation analysis
C4298651|T201|COMP|82513-3|LNC|Hepatitis C virus genotype 3|Hepatitis C virus genotype 3
C4298652|T201|COMP|82512-5|LNC|Hepatitis C virus genotype 1|Hepatitis C virus genotype 1
C4298654|T201|COMP|82509-1|LNC|Gamma interferon.negative control|Gamma interferon.negative control
C4298672|T201|COMP|82508-3|LNC|Ethyl sulfate|Ethyl sulfate
C4298673|T201|COMP|82507-5|LNC|Oligosaccharides pattern|Oligosaccharides pattern
C4298674|T201|COMP|82504-2|LNC|Glutarate|Glutarate
C4298675|T201|COMP|82503-4|LNC|Methylsuccinate|Methylsuccinate
C4298676|T201|COMP|82502-6|LNC|Ethylmalonate|Ethylmalonate
C4298677|T201|COMP|82501-8|LNC|TRBV2 gene segments/TRBV gene segments.total|TRBV2 gene segments/TRBV gene segments.total
C4298678|T201|COMP|82500-0|LNC|TRBV3-1 gene segment/TRBV gene segments.total|TRBV3-1 gene segment/TRBV gene segments.total
C4298679|T201|COMP|82499-5|LNC|TRBV4 gene segments/TRBV gene segments.total|TRBV4 gene segments/TRBV gene segments.total
C4298680|T201|COMP|82498-7|LNC|TRBV5 gene segments/TRBV gene segments.total|TRBV5 gene segments/TRBV gene segments.total
C4298681|T201|COMP|82496-1|LNC|TRBV7 gene segments/TRBV gene segments.total|TRBV7 gene segments/TRBV gene segments.total
C4298682|T201|COMP|82494-6|LNC|TRBV10 gene segments/TRBV gene segments.total|TRBV10 gene segments/TRBV gene segments.total
C4298683|T201|COMP|82493-8|LNC|TRBV11 gene segments/TRBV gene segments.total|TRBV11 gene segments/TRBV gene segments.total
C4298684|T201|COMP|82492-0|LNC|TRBV12 gene segments/TRBV gene segments.total|TRBV12 gene segments/TRBV gene segments.total
C4298685|T201|COMP|82491-2|LNC|TRBV13 gene segments/TRBV gene segments.total|TRBV13 gene segments/TRBV gene segments.total
C4298686|T201|COMP|82490-4|LNC|TRBV14 gene segments/TRBV gene segments.total|TRBV14 gene segments/TRBV gene segments.total
C4298687|T201|COMP|82488-8|LNC|TRBV16 gene segments/TRBV gene segments.total|TRBV16 gene segments/TRBV gene segments.total
C4298688|T201|COMP|82487-0|LNC|TRBV18 gene segments/TRBV gene segments.total|TRBV18 gene segments/TRBV gene segments.total
C4298689|T201|COMP|82485-4|LNC|TRBV20-1 gene segment/TRBV gene segments.total|TRBV20-1 gene segment/TRBV gene segments.total
C4298690|T201|COMP|82484-7|LNC|TRBV24-1 gene segment/TRBV gene segments.total|TRBV24-1 gene segment/TRBV gene segments.total
C4298691|T201|COMP|82483-9|LNC|TRBV25 gene segments/TRBV gene segments.total|TRBV25 gene segments/TRBV gene segments.total
C4298692|T201|COMP|82482-1|LNC|TRBV27 gene segment/TRBV gene segments.total|TRBV27 gene segment/TRBV gene segments.total
C4298693|T201|COMP|82481-3|LNC|TRBV28 gene segment/TRBV gene segments.total|TRBV28 gene segment/TRBV gene segments.total
C4298694|T201|COMP|82480-5|LNC|TRBV29 gene segments/TRBV gene segments.total|TRBV29 gene segments/TRBV gene segments.total
C4298695|T201|COMP|82478-9|LNC|3-Hydroxydecenoylcarnitine (C10:1-OH)|3-Hydroxydecenoylcarnitine (C10:1-OH)
C4298696|T201|COMP|82477-1|LNC|Erythrocyte sedimentation rate|Erythrocyte sedimentation rate
C4298697|T201|COMP|82476-3|LNC|Borrelia miyamotoi (glpQ) gene|Borrelia miyamotoi (glpQ) gene
C4298698|T201|COMP|82474-8|LNC|Borrelia mayonii (oppA1) gene|Borrelia mayonii (oppA1) gene
C4298699|T201|COMP|82473-0|LNC|Borrelia mayonii (oppA1) gene|Borrelia mayonii (oppA1) gene
C4298700|T201|COMP|82471-4|LNC|Borrelia garinii+afzelii (oppA1) gene|Borrelia garinii+afzelii (oppA1) gene
C4298701|T201|COMP|82470-6|LNC|Etanercept|Etanercept
C4298702|T201|COMP|82469-8|LNC|Etanercept Ab|Etanercept Ab
C4298703|T201|COMP|82468-0|LNC|Edoxaban|Edoxaban
C4298704|T201|COMP|82466-4|LNC|riTUXimab Ab|riTUXimab Ab
C4298705|T201|COMP|82465-6|LNC|Mosquito identified|Mosquito identified
C4298706|T201|COMP|82463-1|LNC|Aluminum|Aluminum
C4298707|T201|COMP|82462-3|LNC|Silver|Silver
C4298708|T201|COMP|82461-5|LNC|Influenza virus A & B & H1 2009 pandemic RNA|Influenza virus A & B & H1 2009 pandemic RNA
C4298709|T201|COMP|82458-1|LNC|Gadus chalcogrammus roe Ab.IgE|Gadus chalcogrammus roe Ab.IgE
C4298710|T201|COMP|82457-3|LNC|Human papilloma virus 16 & 18+45 E6+E7 mRNA panel|Human papilloma virus 16 & 18+45 E6+E7 mRNA panel
C4298711|T201|COMP|82456-5|LNC|Human papilloma virus 16 E6+E7 mRNA|Human papilloma virus 16 E6+E7 mRNA
C4298712|T201|COMP|82455-7|LNC|Ganglioside Ab panel|Ganglioside Ab panel
C4298713|T201|COMP|82454-0|LNC|Ganglioside Ab panel|Ganglioside Ab panel
C4298714|T201|COMP|82453-2|LNC|Zo ab|Zo ab
C4298715|T201|COMP|82450-8|LNC|U1 small nuclear ribonucleoprotein 70kD Ab|U1 small nuclear ribonucleoprotein 70kD Ab
C4298716|T201|COMP|82449-0|LNC|Titin Ab|Titin Ab
C4298717|T201|COMP|82448-2|LNC|TIF1-gamma Ab|TIF1-gamma Ab
C4298718|T201|COMP|82447-4|LNC|Sulfatide Ab.IgM|Sulfatide Ab.IgM
C4298719|T201|COMP|82445-8|LNC|Sulfatide Ab|Sulfatide Ab
C4298720|T201|COMP|82444-1|LNC|Glial nuclear type 1 ab|Glial nuclear type 1 ab
C4298721|T201|COMP|82440-9|LNC|SUMO-activating enzyme subunit 1 Ab|SUMO-activating enzyme subunit 1 Ab
C4298722|T201|COMP|82439-1|LNC|SUMO-activating enzyme subunit 1 Ab|SUMO-activating enzyme subunit 1 Ab
C4298723|T201|COMP|82432-6|LNC|Platelet-derived growth factor receptor Ab|Platelet-derived growth factor receptor Ab
C4298724|T201|COMP|82430-0|LNC|OJ Ab|OJ Ab
C4298725|T201|COMP|82426-8|LNC|MJ Ab|MJ Ab
C4298726|T201|COMP|82425-0|LNC|MJ Ab|MJ Ab
C4298727|T201|COMP|82424-3|LNC|MDA5 Ab|MDA5 Ab
C4298728|T201|COMP|82423-5|LNC|Ma+Ta Ab|Ma+Ta Ab
C4298729|T201|COMP|82421-9|LNC|Ks Ab|Ks Ab
C4298730|T201|COMP|82418-5|LNC|Human upstream binding factor Ab|Human upstream binding factor Ab
C4298731|T201|COMP|82417-7|LNC|Human upstream binding factor Ab|Human upstream binding factor Ab
C4298732|T201|COMP|82415-1|LNC|Ha Ab|Ha Ab
C4298733|T201|COMP|82414-4|LNC|Ha Ab|Ha Ab
C4298734|T201|COMP|82411-0|LNC|Ganglioside GT1a Ab.IgG|Ganglioside GT1a Ab.IgG
C4298735|T201|COMP|82409-4|LNC|Ganglioside GM4 Ab.IgM|Ganglioside GM4 Ab.IgM
C4298736|T201|COMP|82402-9|LNC|Ganglioside GD3 Ab.IgG|Ganglioside GD3 Ab.IgG
C4298737|T201|COMP|82401-1|LNC|Ganglioside GD2 Ab.IgM|Ganglioside GD2 Ab.IgM
C4298738|T201|COMP|82400-3|LNC|Ganglioside GD2 Ab.IgG+IgM|Ganglioside GD2 Ab.IgG+IgM
C4298739|T201|COMP|82398-9|LNC|Ganglioside GD1b Ab.IgG+IgM|Ganglioside GD1b Ab.IgG+IgM
C4298740|T201|COMP|82397-1|LNC|Ganglioside GD1a Ab.IgM|Ganglioside GD1a Ab.IgM
C4298741|T201|COMP|82395-5|LNC|Ganglioside GD1a Ab.IgG|Ganglioside GD1a Ab.IgG
C4298742|T201|COMP|82393-0|LNC|Fibrillarin Ab|Fibrillarin Ab
C4298743|T201|COMP|82392-2|LNC|Ej Ab|Ej Ab
C4298744|T201|COMP|82390-6|LNC|Centromere protein A Ab|Centromere protein A Ab
C4298749|T201|COMP|82379-9|LNC|Daclatasvir|Daclatasvir
C4298750|T201|COMP|82378-1|LNC|Ombitasvir|Ombitasvir
C4298751|T201|COMP|82377-3|LNC|Ledipasvir|Ledipasvir
C4298752|T201|COMP|82376-5|LNC|Elbasvir|Elbasvir
C4298753|T201|COMP|82375-7|LNC|Norbuprenorphine|Norbuprenorphine
C4298754|T201|COMP|82374-0|LNC|Norbuprenorphine|Norbuprenorphine
C4298755|T201|COMP|82372-4|LNC|Buprenorphine|Buprenorphine
C4298756|T201|COMP|82371-6|LNC|Norbuprenorphine|Norbuprenorphine
C4298757|T201|COMP|82370-8|LNC|Norbuprenorphine|Norbuprenorphine
C4298758|T201|COMP|82369-0|LNC|Buprenorphine|Buprenorphine
C4298759|T201|COMP|82368-2|LNC|Thyroid secretory capacity|Thyroid secretory capacity
C4298760|T201|COMP|82367-4|LNC|Peripheral deiodinase activity|Peripheral deiodinase activity
C4298767|T201|COMP|82354-2|LNC|Human papilloma virus 16 & 18+45 E6+E7 mRNA|Human papilloma virus 16 & 18+45 E6+E7 mRNA
C4298781|T201|COMP|82334-4|LNC|Interleukin 17A|Interleukin 17A
C4298782|T201|COMP|82309-6|LNC|Basis for allelic phase|Basis for allelic phase
C4298783|T201|COMP|82306-2|LNC|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C4298784|T201|COMP|82305-4|LNC|Gastrointestinal pathogens panel|Gastrointestinal pathogens panel
C4298785|T201|COMP|82304-7|LNC|Plesiomonas shigelloides|Plesiomonas shigelloides
C4298786|T201|COMP|82301-3|LNC|Salmonella sp|Salmonella sp
C4298787|T201|COMP|82300-5|LNC|Shigella sp|Shigella sp
C4298788|T201|COMP|82299-9|LNC|Escherichia coli shiga-like toxin 1+2|Escherichia coli shiga-like toxin 1+2
C4298789|T201|COMP|82298-1|LNC|Yersinia enterocolitica|Yersinia enterocolitica
C4298790|T201|COMP|82223-9|LNC|Cystathionine beta synthase|Cystathionine beta synthase
C4298791|T201|COMP|82222-1|LNC|Amylo-alpha-1,6-glucosidase|Amylo-alpha-1,6-glucosidase
C4298792|T201|COMP|82221-3|LNC|Alpha-methylacyl CoA racemase|Alpha-methylacyl CoA racemase
C4298793|T201|COMP|82220-5|LNC|Alkyl-dihydroxyacetonephosphate synthase|Alkyl-dihydroxyacetonephosphate synthase
C4298794|T201|COMP|82219-7|LNC|3-Methylglutaconyl-CoA hydratase|3-Methylglutaconyl-CoA hydratase
C4298795|T201|COMP|82217-1|LNC|3-Hydroxyisobutyryl-CoA hydrolase|3-Hydroxyisobutyryl-CoA hydrolase
C4298800|T201|COMP|82869-9|LNC|6-Thioguanine & 6-methylmercaptopurine panel|6-Thioguanine & 6-methylmercaptopurine panel
C4298801|T201|COMP|82868-1|LNC|Allo-pregnanediolone|Allo-pregnanediolone
C4298802|T201|COMP|82867-3|LNC|Allo-pregnanediolone|Allo-pregnanediolone
C4298809|T201|COMP|82408-6|LNC|Ganglioside GM4 Ab.IgG+IgM|Ganglioside GM4 Ab.IgG+IgM
C4298810|T201|COMP|82407-8|LNC|Ganglioside GM4 Ab.IgG|Ganglioside GM4 Ab.IgG
C4298811|T201|COMP|82404-5|LNC|Ganglioside GD3 Ab.IgM|Ganglioside GD3 Ab.IgM
C4298815|T201|COMP|82385-6|LNC|Methylmalonate|Methylmalonate
C4298816|T201|COMP|82384-9|LNC|Dengue virus 1+3 RNA|Dengue virus 1+3 RNA
C4298820|T201|COMP|82528-1|LNC|VHL gene full mutation analysis|VHL gene full mutation analysis
C4298864|T201|COMP|82438-3|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C4298865|T201|COMP|82437-5|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C4298866|T201|COMP|82435-9|LNC|RNA polymerase III Ab|RNA polymerase III Ab
C4298867|T201|COMP|82434-2|LNC|Ribosomal Ab|Ribosomal Ab
C4298868|T201|COMP|82433-4|LNC|Proteinase 3 Ab|Proteinase 3 Ab
C4298869|T201|COMP|82427-6|LNC|Myeloperoxidase Ab|Myeloperoxidase Ab
C4298870|T201|COMP|82420-1|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C4298871|T201|COMP|82419-3|LNC|Intrinsic factor Ab|Intrinsic factor Ab
C4298872|T201|COMP|82412-8|LNC|Ganglioside GT1a Ab.IgG+IgM|Ganglioside GT1a Ab.IgG+IgM
C4298873|T201|COMP|82403-7|LNC|Ganglioside GD3 Ab.IgG+IgM|Ganglioside GD3 Ab.IgG+IgM
C4298874|T201|COMP|82405-2|LNC|Ganglioside GM3 Ab.IgG+IgM|Ganglioside GM3 Ab.IgG+IgM
C4318511|T201|COMP|85346-5|LNC|Tissue blocks examined|Tissue blocks examined
C4318512|T201|COMP|85348-1|LNC|Procedure used to obtain tumor specimen|Procedure used to obtain tumor specimen
C4318516|T201|COMP|85363-0|LNC|21-Hydroxylase Ab|21-Hydroxylase Ab
C4318526|T201|COMP|85779-7|LNC|Neisseria meningitidis DNA|Neisseria meningitidis DNA
C4318539|T201|COMP|85424-0|LNC|Imipenem+Relebactam|Imipenem+Relebactam
C4318540|T201|COMP|85426-5|LNC|Meropenem|Meropenem
C4318541|T201|COMP|85428-1|LNC|Penicillin|Penicillin
C4318670|T201|COMP|85478-6|LNC|Influenza virus B RNA|Influenza virus B RNA
C4318672|T201|COMP|85487-7|LNC|S little c super 1 Ag|S little c super 1 Ag
C4318673|T201|COMP|85488-5|LNC|S little c super 2 Ag|S little c super 2 Ag
C4318675|T201|COMP|85497-6|LNC|cloZAPine N-oxide|cloZAPine N-oxide
C4318676|T201|COMP|85499-2|LNC|Bacterial carbapenem resistance blaKPC gene|Bacterial carbapenem resistance blaKPC gene
C4318677|T201|COMP|85505-6|LNC|Rh.presumptive|Rh.presumptive
C4318678|T201|COMP|85507-2|LNC|PIK3CA gene targeted mutation analysis|PIK3CA gene targeted mutation analysis
C4318679|T201|COMP|85509-8|LNC|KRAS gene targeted mutation analysis|KRAS gene targeted mutation analysis
C4318780|T201|COMP|85625-2|LNC|Kidney failure 5Y risk|Kidney failure 5Y risk
C4318781|T201|COMP|85627-8|LNC|Haemophilus influenzae hpd gene|Haemophilus influenzae hpd gene
C4318792|T201|COMP|85679-9|LNC|Haemophilus influenzae bex gene|Haemophilus influenzae bex gene
C4318793|T201|COMP|85680-7|LNC|Haemophilus influenzae ecs gene|Haemophilus influenzae ecs gene
C4318794|T201|COMP|85686-4|LNC|HIV 1 Ab|HIV 1 Ab
C4318796|T201|COMP|85690-6|LNC|Rubella virus genotype|Rubella virus genotype
C4318866|T201|COMP|85737-5|LNC|Bombay phenotype|Bombay phenotype
C4318867|T201|COMP|85739-1|LNC|Bombay phenotype|Bombay phenotype
C4318868|T201|COMP|85741-7|LNC|Streptococcus pneumoniae Danish serotype 4 DNA|Streptococcus pneumoniae Danish serotype 4 DNA
C4318869|T201|COMP|85746-6|LNC|Streptococcus pneumoniae Danish serotype 14 DNA|Streptococcus pneumoniae Danish serotype 14 DNA
C4318873|T201|COMP|85765-6|LNC|Staphylococcus aureus DNA|Staphylococcus aureus DNA
C4318874|T201|COMP|85767-2|LNC|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C4318875|T201|COMP|85774-8|LNC|Klebsiella oxytoca DNA|Klebsiella oxytoca DNA
C4318876|T201|COMP|85776-3|LNC|Proteus sp DNA|Proteus sp DNA
C4318877|T201|COMP|85777-1|LNC|Serratia marcescens DNA|Serratia marcescens DNA
C4318878|T201|COMP|85788-8|LNC|Bacterial carbapenem resistance blaKPC gene|Bacterial carbapenem resistance blaKPC gene
C4318879|T201|COMP|85790-4|LNC|Cells.CD3+CD8+CD45RO+|Cells.CD3+CD8+CD45RO+
C4318880|T201|COMP|85791-2|LNC|Cells.CD3+CD4+CD45RO+/100 cells.CD3|Cells.CD3+CD4+CD45RO+/100 cells.CD3
C4318881|T201|COMP|85797-9|LNC|Neisseria meningitidis serogroup DNA panel|Neisseria meningitidis serogroup DNA panel
C4318882|T201|COMP|85798-7|LNC|Measles virus N gene|Measles virus N gene
C4318883|T201|COMP|85800-1|LNC|Mumps virus SH gene|Mumps virus SH gene
C4318884|T201|COMP|85807-6|LNC|Mumps virus genotype|Mumps virus genotype
C4318885|T201|COMP|85808-4|LNC|Mumps virus RNA & SH gene panel|Mumps virus RNA & SH gene panel
C4318887|T201|COMP|85818-3|LNC|Clot formation+Clotting time|Clot formation+Clotting time
C4318888|T201|COMP|85824-1|LNC|Bacterial carbapenem resistance blaIMP gene|Bacterial carbapenem resistance blaIMP gene
C4318893|T201|COMP|85837-3|LNC|Bacterial beta-lactam resistance ESBL blaPER gene|Bacterial beta-lactam resistance ESBL blaPER gene
C4318962|T201|COMP|85954-6|LNC|Streptococcus pneumoniae Danish serotype 1 Ab.IgG|Streptococcus pneumoniae Danish serotype 1 Ab.IgG
C4318967|T201|COMP|86620-2|LNC|Bacterial methicillin resistance mecA+mecC genes|Bacterial methicillin resistance mecA+mecC genes
C4318968|T201|COMP|86621-0|LNC|Bacterial methicillin resistance mecC gene|Bacterial methicillin resistance mecC gene
C4318974|T201|COMP|85973-6|LNC|Streptococcus pneumoniae Danish serotype 12F Ab|Streptococcus pneumoniae Danish serotype 12F Ab
C4319031|T201|COMP|85990-0|LNC|Streptococcus pneumoniae Danish serotype 14 Ab|Streptococcus pneumoniae Danish serotype 14 Ab
C4319039|T201|COMP|86019-7|LNC|Streptococcus pneumoniae Danish serotype 19F Ab|Streptococcus pneumoniae Danish serotype 19F Ab
C4319055|T201|COMP|86079-1|LNC|Streptococcus pneumoniae Danish serotype 3 Ab|Streptococcus pneumoniae Danish serotype 3 Ab
C4319061|T201|COMP|86107-0|LNC|Streptococcus pneumoniae Danish serotype 4 Ab.IgG|Streptococcus pneumoniae Danish serotype 4 Ab.IgG
C4319115|T201|COMP|86108-8|LNC|Streptococcus pneumoniae Danish serotype 4 Ab.IgG|Streptococcus pneumoniae Danish serotype 4 Ab.IgG
C4319116|T201|COMP|86110-4|LNC|Streptococcus pneumoniae Danish serotype 4 Ab.IgG|Streptococcus pneumoniae Danish serotype 4 Ab.IgG
C4319117|T201|COMP|86226-8|LNC|Codeine|Codeine
C4319118|T201|COMP|86228-4|LNC|Ethyl sulfate|Ethyl sulfate
C4319121|T201|COMP|86515-4|LNC|Chikungunya virus RNA|Chikungunya virus RNA
C4319122|T201|COMP|86517-0|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C4319123|T201|COMP|86716-8|LNC|Actinobacillus pleuropneumoniae DNA|Actinobacillus pleuropneumoniae DNA
C4319124|T201|COMP|86718-4|LNC|Actinobacillus pleuropneumoniae serotype 3 Ab|Actinobacillus pleuropneumoniae serotype 3 Ab
C4319129|T201|COMP|86130-2|LNC|Streptococcus pneumoniae Danish serotype 5 Ab.IgG|Streptococcus pneumoniae Danish serotype 5 Ab.IgG
C4319134|T201|COMP|86150-0|LNC|Streptococcus pneumoniae Danish serotype 8 Ab.IgG|Streptococcus pneumoniae Danish serotype 8 Ab.IgG
C4319138|T201|COMP|86163-3|LNC|Streptococcus pneumoniae Danish serotype 9N Ab|Streptococcus pneumoniae Danish serotype 9N Ab
C4319139|T201|COMP|86165-8|LNC|Streptococcus pneumoniae Danish serotype 9N Ab|Streptococcus pneumoniae Danish serotype 9N Ab
C4319145|T201|COMP|86191-4|LNC|Eutylone|Eutylone
C4319146|T201|COMP|86197-1|LNC|Pentylone|Pentylone
C4319147|T201|COMP|86198-9|LNC|Neisseria meningitidis serogroup Y synF gene|Neisseria meningitidis serogroup Y synF gene
C4319198|T201|COMP|86200-3|LNC|Porcine epidemic diarrhea virus|Porcine epidemic diarrhea virus
C4319200|T201|COMP|86207-8|LNC|Porcine epidemic diarrhea virus Ab.IgG|Porcine epidemic diarrhea virus Ab.IgG
C4319211|T201|COMP|86217-7|LNC|Rotavirus A VP6 capsid protein|Rotavirus A VP6 capsid protein
C4319212|T201|COMP|86219-3|LNC|Porcine epidemic diarrhea virus Ab.IgG|Porcine epidemic diarrhea virus Ab.IgG
C4319213|T201|COMP|86221-9|LNC|Bacterial colistin resistance mcr-1 gene|Bacterial colistin resistance mcr-1 gene
C4319214|T201|COMP|86234-2|LNC|Neisseria meningitidis serogroup A sacB gene|Neisseria meningitidis serogroup A sacB gene
C4319215|T201|COMP|86236-7|LNC|Neisseria meningitidis serogroup C synE gene|Neisseria meningitidis serogroup C synE gene
C4319217|T201|COMP|86271-4|LNC|Transferrin.gastrointestinal|Transferrin.gastrointestinal
C4319227|T201|COMP|86317-5|LNC|Influenza virus A H1 2009 pandemic RNA|Influenza virus A H1 2009 pandemic RNA
C4319228|T201|COMP|86319-1|LNC|Staphylococcus aureus|Staphylococcus aureus
C4319229|T201|COMP|86325-8|LNC|Bordetella pertussis+parapertussis ptxS1 gene|Bordetella pertussis+parapertussis ptxS1 gene
C4319230|T201|COMP|86327-4|LNC|Bordetella parapertussis IS1001 DNA|Bordetella parapertussis IS1001 DNA
C4319285|T201|COMP|86328-2|LNC|Adenovirus 21 DNA|Adenovirus 21 DNA
C4319286|T201|COMP|86334-0|LNC|Adenovirus 3 DNA|Adenovirus 3 DNA
C4319288|T201|COMP|86342-3|LNC|Streptococcus pneumoniae Danish serotype 6A+6B Ab|Streptococcus pneumoniae Danish serotype 6A+6B Ab
C4319315|T201|COMP|86458-7|LNC|Brucella sp Ab|Brucella sp Ab
C4319371|T201|COMP|85298-8|LNC|Body structure included in specimen|Body structure included in specimen
C4319374|T201|COMP|85537-9|LNC|Mycoplasma hyosynoviae 16S rRNA gene|Mycoplasma hyosynoviae 16S rRNA gene
C4319387|T201|COMP|86542-8|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C4319388|T201|COMP|86544-4|LNC|Herpes virus 7 DNA|Herpes virus 7 DNA
C4319389|T201|COMP|86545-1|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C4319393|T201|COMP|86564-2|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C4319394|T201|COMP|86565-9|LNC|Influenza virus A Ag|Influenza virus A Ag
C4319395|T201|COMP|86567-5|LNC|Influenza virus A Ab.IgM|Influenza virus A Ab.IgM
C4319396|T201|COMP|86575-8|LNC|Measles virus RNA|Measles virus RNA
C4319397|T201|COMP|86577-4|LNC|Measles virus RNA|Measles virus RNA
C4319398|T201|COMP|86588-1|LNC|Rabies virus RNA|Rabies virus RNA
C4319399|T201|COMP|86590-7|LNC|Streptococcus pneumoniae Ag|Streptococcus pneumoniae Ag
C4319400|T201|COMP|86592-3|LNC|Varicella zoster virus Ag|Varicella zoster virus Ag
C4319401|T201|COMP|86605-3|LNC|Alpha hydroxytriazolam/Creatinine|Alpha hydroxytriazolam/Creatinine
C4319402|T201|COMP|86607-9|LNC|Cocaine/Creatinine|Cocaine/Creatinine
C4319403|T201|COMP|86609-5|LNC|Noroxymorphone/Creatinine|Noroxymorphone/Creatinine
C4319447|T201|COMP|85762-3|LNC|Blood pathogens panel|Blood pathogens panel
C4319448|T201|COMP|85764-9|LNC|Staphylococcus sp DNA|Staphylococcus sp DNA
C4319455|T201|COMP|85281-4|LNC|Intratumoral lymphocytic response|Intratumoral lymphocytic response
C4319458|T201|COMP|85290-5|LNC|Surgical margin tumor involvement|Surgical margin tumor involvement
C4319459|T201|COMP|85302-8|LNC|Growth pattern of DCIS|Growth pattern of DCIS
C4319462|T201|COMP|85311-9|LNC|Extent of anterior margin carcinoma involvement|Extent of anterior margin carcinoma involvement
C4319463|T201|COMP|85312-7|LNC|Extent of inferior margin carcinoma involvement|Extent of inferior margin carcinoma involvement
C4319464|T201|COMP|85314-3|LNC|Extent of medial margin carcinoma involvement|Extent of medial margin carcinoma involvement
C4319465|T201|COMP|85325-9|LNC|Cells.progesterone receptor/100 cells|Cells.progesterone receptor/100 cells
C4319466|T201|COMP|85327-5|LNC|Foci|Foci
C4319467|T201|COMP|85329-1|LNC|Cells.estrogen receptor/100 cells|Cells.estrogen receptor/100 cells
C4319468|T201|COMP|85335-8|LNC|DCIS.additional dimension 2|DCIS.additional dimension 2
C4319469|T201|COMP|85337-4|LNC|Estrogen receptor Ag|Estrogen receptor Ag
C4319474|T201|COMP|86667-3|LNC|Level of tumor invasion|Level of tumor invasion
C4319475|T201|COMP|86669-9|LNC|Mitotic figures|Mitotic figures
C4319477|T201|COMP|86696-2|LNC|Rotavirus B RNA|Rotavirus B RNA
C4319478|T201|COMP|86704-4|LNC|Lawsonia intracellularis RNA|Lawsonia intracellularis RNA
C4319479|T201|COMP|86705-1|LNC|Lawsonia intracellularis Ab|Lawsonia intracellularis Ab
C4319480|T201|COMP|86710-1|LNC|Porcine epidemic diarrhea virus RNA|Porcine epidemic diarrhea virus RNA
C4319481|T201|COMP|86726-7|LNC|Erysipelothrix rhusiopathiae DNA|Erysipelothrix rhusiopathiae DNA
C4319482|T201|COMP|86732-5|LNC|Leptospira sp identified|Leptospira sp identified
C4319483|T201|COMP|86734-1|LNC|Porcine parvovirus Ab|Porcine parvovirus Ab
C4319485|T201|COMP|86742-4|LNC|Growth phase|Growth phase
C4319489|T201|COMP|86860-4|LNC|Dengue virus 1 Ab.Neut|Dengue virus 1 Ab.Neut
C4319924|T201|COMP|85299-6|LNC|Serine-threonine protein kinase B-raf V600E|Serine-threonine protein kinase B-raf V600E
C4321527|T201|COMP|86243-3|LNC|Color|Color
C4321539|T201|COMP|85930-6|LNC|Date specimen sent to CDC|Date specimen sent to CDC
C4482452|T201|COMP|82743-6|LNC|Cells.CD8+CD45RA+|Cells.CD8+CD45RA+
C4482453|T201|COMP|82744-4|LNC|Cells.CD8+CD45RA+/100 cells.CD8|Cells.CD8+CD45RA+/100 cells.CD8
C4482614|T201|COMP|85316-8|LNC|Extent of superior margin carcinoma involvement|Extent of superior margin carcinoma involvement
C4482616|T201|COMP|85317-6|LNC|DCIS.max dimension|DCIS.max dimension
C4482618|T201|COMP|85318-4|LNC|HER2|HER2
C4482619|T201|COMP|85319-2|LNC|HER2|HER2
C4482620|T201|COMP|85296-2|LNC|Tumor budding|Tumor budding
C4482621|T201|COMP|85297-0|LNC|Tumor buds|Tumor buds
C4482624|T201|COMP|85300-2|LNC|Mitotic rate|Mitotic rate
C4482634|T201|COMP|85536-1|LNC|Mycoplasma hyopneumoniae DNA|Mycoplasma hyopneumoniae DNA
C4482635|T201|COMP|85538-7|LNC|Mycoplasma hyorhinis 16S rRNA gene|Mycoplasma hyorhinis 16S rRNA gene
C4482653|T201|COMP|85843-1|LNC|Bacterial beta-lactam resistance AmpC blaFOX gene|Bacterial beta-lactam resistance AmpC blaFOX gene
C4482667|T201|COMP|85761-5|LNC|Klebsiella pneumoniae DNA|Klebsiella pneumoniae DNA
C4482669|T201|COMP|85763-1|LNC|Listeria monocytogenes DNA|Listeria monocytogenes DNA
C4482688|T201|COMP|85275-6|LNC|Adjacent structure invaded by tumor|Adjacent structure invaded by tumor
C4482694|T201|COMP|85279-8|LNC|Excised length|Excised length
C4482697|T201|COMP|85282-2|LNC|Mucinous fraction|Mucinous fraction
C4482699|T201|COMP|85283-0|LNC|Organ tumor is adherent to|Organ tumor is adherent to
C4482701|T201|COMP|85284-8|LNC|Peritumoral lymphocytic response|Peritumoral lymphocytic response
C4482703|T201|COMP|85285-5|LNC|Polyp in which invasive carcinoma arose|Polyp in which invasive carcinoma arose
C4482704|T201|COMP|85286-3|LNC|Promoter methylation testing method|Promoter methylation testing method
C4482708|T201|COMP|85289-7|LNC|Signet ring cells/100 cells|Signet ring cells/100 cells
C4482711|T201|COMP|85291-3|LNC|Surgical margin tumor involvement.deep|Surgical margin tumor involvement.deep
C4482712|T201|COMP|85292-1|LNC|Surgical margin tumor involvement.distant|Surgical margin tumor involvement.distant
C4482713|T201|COMP|85293-9|LNC|Surgical margin tumor involvement.mesenteric|Surgical margin tumor involvement.mesenteric
C4482715|T201|COMP|85294-7|LNC|Surgical margin tumor involvement.mucosal|Surgical margin tumor involvement.mucosal
C4482716|T201|COMP|85295-4|LNC|Surgical margin tumor involvement.proximal|Surgical margin tumor involvement.proximal
C4482717|T201|COMP|85301-0|LNC|Adjacent structure invaded by tumor|Adjacent structure invaded by tumor
C4482719|T201|COMP|85303-6|LNC|Body structure of origin|Body structure of origin
C4482731|T201|COMP|85310-1|LNC|Estrogen receptor fluorescence intensity|Estrogen receptor fluorescence intensity
C4482735|T201|COMP|85313-5|LNC|Extent of lateral margin carcinoma involvement|Extent of lateral margin carcinoma involvement
C4482738|T201|COMP|85315-0|LNC|Extent of posterior margin carcinoma involvement|Extent of posterior margin carcinoma involvement
C4482740|T201|COMP|85320-0|LNC|Foci|Foci
C4482741|T201|COMP|85321-8|LNC|Glandular differentiation|Glandular differentiation
C4482742|T201|COMP|85322-6|LNC|Adjacent structure invaded by tumor|Adjacent structure invaded by tumor
C4482743|T201|COMP|85323-4|LNC|Response to neoadjuvant therapy|Response to neoadjuvant therapy
C4482744|T201|COMP|85326-7|LNC|Tissue blocks positive for DCIS|Tissue blocks positive for DCIS
C4482748|T201|COMP|85330-9|LNC|Cells.Ki-67 nuclear Ag/100 cells|Cells.Ki-67 nuclear Ag/100 cells
C4482749|T201|COMP|85331-7|LNC|Progesterone receptor fluorescence intensity|Progesterone receptor fluorescence intensity
C4482751|T201|COMP|85332-5|LNC|Radial position within breast|Radial position within breast
C4482753|T201|COMP|85333-3|LNC|DCIS.additional dimension 1|DCIS.additional dimension 1
C4482755|T201|COMP|85334-1|LNC|Surgical margin DCIS involvement|Surgical margin DCIS involvement
C4482758|T201|COMP|85336-6|LNC|DCIS intraductal extension|DCIS intraductal extension
C4482760|T201|COMP|85338-2|LNC|Lobular carcinoma in situ|Lobular carcinoma in situ
C4482761|T201|COMP|85339-0|LNC|Progesterone receptor Ag|Progesterone receptor Ag
C4482762|T201|COMP|85340-8|LNC|DCIS necrosis|DCIS necrosis
C4482764|T201|COMP|85341-6|LNC|Pathology report reviewed|Pathology report reviewed
C4482766|T201|COMP|85342-4|LNC|Lymph node site of origin|Lymph node site of origin
C4482768|T201|COMP|85343-2|LNC|Lymph nodes with macrometastases|Lymph nodes with macrometastases
C4482770|T201|COMP|85344-0|LNC|Lymph nodes with micrometastases|Lymph nodes with micrometastases
C4482771|T201|COMP|85345-7|LNC|Dermal lymph-vascular invasion|Dermal lymph-vascular invasion
C4482774|T201|COMP|85347-3|LNC|Sentinel lymph nodes examined|Sentinel lymph nodes examined
C4482777|T201|COMP|85349-9|LNC|Lymph node response to neoadjuvant therapy|Lymph node response to neoadjuvant therapy
C4482778|T201|COMP|85350-7|LNC|Extranodal extension of carcinoma|Extranodal extension of carcinoma
C4482780|T201|COMP|85351-5|LNC|Lymph node metastatic deposit.max dimension|Lymph node metastatic deposit.max dimension
C4482782|T201|COMP|85352-3|LNC|Lymph nodes with isolated tumor cells|Lymph nodes with isolated tumor cells
C4482790|T201|COMP|85358-0|LNC|Phosphatidylserine-prothrombin complex Ab.IgM|Phosphatidylserine-prothrombin complex Ab.IgM
C4482791|T201|COMP|85359-8|LNC|Phosphatidylserine-prothrombin complex Ab.IgG|Phosphatidylserine-prothrombin complex Ab.IgG
C4482795|T201|COMP|85361-4|LNC|HIV 1+2 RNA|HIV 1+2 RNA
C4482797|T201|COMP|85362-2|LNC|Mycobacterium tuberculosis complex DNA|Mycobacterium tuberculosis complex DNA
C4482799|T201|COMP|85364-8|LNC|Muscarinic acetylcholine receptor M3 Ab|Muscarinic acetylcholine receptor M3 Ab
C4482800|T201|COMP|85365-5|LNC|Neutrophil membrane Ab|Neutrophil membrane Ab
C4482802|T201|COMP|85366-3|LNC|Neutrophil membrane Ab.IgM|Neutrophil membrane Ab.IgM
C4482804|T201|COMP|85367-1|LNC|Neutrophil membrane Ab.IgG|Neutrophil membrane Ab.IgG
C4482806|T201|COMP|85368-9|LNC|HIV 1+2 RNA|HIV 1+2 RNA
C4482807|T201|COMP|85369-7|LNC|Neutrophils|Neutrophils
C4482819|T201|COMP|85379-6|LNC|Purine/pyrimidine|Purine/pyrimidine
C4482845|T201|COMP|85780-5|LNC|Pseudomonas aeruginosa DNA|Pseudomonas aeruginosa DNA
C4482846|T201|COMP|85781-3|LNC|Candida albicans DNA|Candida albicans DNA
C4482855|T201|COMP|85380-4|LNC|HIV immunoassay testing algorithm interpretation|HIV immunoassay testing algorithm interpretation
C4482857|T201|COMP|85381-2|LNC|Isavuconazole|Isavuconazole
C4482858|T201|COMP|85382-0|LNC|Osmolarity|Osmolarity
C4482859|T201|COMP|85383-8|LNC|EGFR gene.c.2369C>T actual/normal|EGFR gene.c.2369C>T actual/normal
C4482861|T201|COMP|85384-6|LNC|Amisulpride|Amisulpride
C4482901|T201|COMP|85421-6|LNC|Bacterial identification & susceptibility panel|Bacterial identification & susceptibility panel
C4482903|T201|COMP|85422-4|LNC|ceFAZolin|ceFAZolin
C4482905|T201|COMP|85423-2|LNC|Eravacycline|Eravacycline
C4482907|T201|COMP|85425-7|LNC|Lefamulin|Lefamulin
C4482909|T201|COMP|85427-3|LNC|Meropenem+Vaborbactam|Meropenem+Vaborbactam
C4482911|T201|COMP|85429-9|LNC|Penicillin|Penicillin
C4482959|T201|COMP|85477-8|LNC|Influenza virus A RNA|Influenza virus A RNA
C4482960|T201|COMP|85479-4|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C4482969|T201|COMP|85485-1|LNC|B little g super little b Ag|B little g super little b Ag
C4482971|T201|COMP|85486-9|LNC|B little g super little c Ag|B little g super little c Ag
C4482987|T201|COMP|85496-8|LNC|Streptococcus pneumoniae serotype|Streptococcus pneumoniae serotype
C4482988|T201|COMP|85498-4|LNC|Bacterial carbapenem resistance blaIMP gene|Bacterial carbapenem resistance blaIMP gene
C4482990|T201|COMP|85500-7|LNC|Bacterial carbapenem resistance blaNDM gene|Bacterial carbapenem resistance blaNDM gene
C4482991|T201|COMP|85501-5|LNC|Bacterial carbapenem resistance blaVIM gene|Bacterial carbapenem resistance blaVIM gene
C4482992|T201|COMP|85502-3|LNC|Bacterial carbapenem resistance genes panel|Bacterial carbapenem resistance genes panel
C4482994|T201|COMP|85503-1|LNC|Bacterial carbapenem resistance blaOXA-48 gene|Bacterial carbapenem resistance blaOXA-48 gene
C4482996|T201|COMP|85504-9|LNC|ABO group.presumptive|ABO group.presumptive
C4482999|T201|COMP|85506-4|LNC|PTEN gene targeted mutation analysis|PTEN gene targeted mutation analysis
C4483000|T201|COMP|85508-0|LNC|Satellite nodules|Satellite nodules
C4483001|T201|COMP|85510-6|LNC|NRAS gene targeted mutation analysis|NRAS gene targeted mutation analysis
C4483002|T201|COMP|85511-4|LNC|BRAF gene targeted mutation analysis|BRAF gene targeted mutation analysis
C4483003|T201|COMP|85512-2|LNC|Hepatitis D virus RNA|Hepatitis D virus RNA
C4483004|T201|COMP|85513-0|LNC|Hepatitis D virus RNA|Hepatitis D virus RNA
C4483013|T201|COMP|85526-2|LNC|Influenza virus D PB2 gene|Influenza virus D PB2 gene
C4483019|T201|COMP|85532-0|LNC|Influenza virus A whole genome|Influenza virus A whole genome
C4483041|T201|COMP|85553-6|LNC|Mycoplasma flocculare 16S rRNA gene|Mycoplasma flocculare 16S rRNA gene
C4483072|T201|COMP|85582-5|LNC|Chikungunya virus RNA+Dengue virus RNA|Chikungunya virus RNA+Dengue virus RNA
C4483074|T201|COMP|85583-3|LNC|Chikungunya virus RNA|Chikungunya virus RNA
C4483075|T201|COMP|85584-1|LNC|Dengue virus RNA|Dengue virus RNA
C4483117|T201|COMP|85621-1|LNC|Zika virus RNA|Zika virus RNA
C4483118|T201|COMP|85622-9|LNC|Zika virus RNA|Zika virus RNA
C4483119|T201|COMP|85623-7|LNC|Zika virus RNA|Zika virus RNA
C4483120|T201|COMP|85624-5|LNC|Kidney failure 2Y risk|Kidney failure 2Y risk
C4483123|T201|COMP|85626-0|LNC|Kidney failure 2Y & 5Y risk panel|Kidney failure 2Y & 5Y risk panel
C4483126|T201|COMP|85628-6|LNC|Neisseria meningitidis sodC gene|Neisseria meningitidis sodC gene
C4483186|T201|COMP|85678-1|LNC|Haemophilus influenzae acs gene|Haemophilus influenzae acs gene
C4483190|T201|COMP|85681-5|LNC|Haemophilus influenzae dcs gene|Haemophilus influenzae dcs gene
C4483192|T201|COMP|85682-3|LNC|Haemophilus influenzae ccs gene|Haemophilus influenzae ccs gene
C4483194|T201|COMP|85683-1|LNC|Haemophilus influenzae bcs gene|Haemophilus influenzae bcs gene
C4483196|T201|COMP|85684-9|LNC|Bordetella pertussis.pertussis toxin Ab.IgG|Bordetella pertussis.pertussis toxin Ab.IgG
C4483198|T201|COMP|85685-6|LNC|Mycoplasma hyopneumoniae P146 gene|Mycoplasma hyopneumoniae P146 gene
C4483200|T201|COMP|85688-0|LNC|Streptococcus pneumoniae lytA gene|Streptococcus pneumoniae lytA gene
C4483238|T201|COMP|85738-3|LNC|Bombay phenotype|Bombay phenotype
C4483239|T201|COMP|85740-9|LNC|Streptococcus pneumoniae Danish serotype 5 DNA|Streptococcus pneumoniae Danish serotype 5 DNA
C4483242|T201|COMP|85742-5|LNC|Streptococcus pneumoniae Danish serotype 3 DNA|Streptococcus pneumoniae Danish serotype 3 DNA
C4483244|T201|COMP|85743-3|LNC|Streptococcus pneumoniae Danish serotype 23F DNA|Streptococcus pneumoniae Danish serotype 23F DNA
C4483246|T201|COMP|85744-1|LNC|Streptococcus pneumoniae Danish serotype 2 DNA|Streptococcus pneumoniae Danish serotype 2 DNA
C4483248|T201|COMP|85745-8|LNC|Streptococcus pneumoniae Danish serotype 19F DNA|Streptococcus pneumoniae Danish serotype 19F DNA
C4483251|T201|COMP|85747-4|LNC|Streptococcus pneumoniae Danish serotype 1 DNA|Streptococcus pneumoniae Danish serotype 1 DNA
C4483256|T201|COMP|85750-8|LNC|Streptococcus pneumoniae Danish serotype 23A DNA|Streptococcus pneumoniae Danish serotype 23A DNA
C4483258|T201|COMP|85751-6|LNC|Streptococcus pneumoniae Danish serotype 16F DNA|Streptococcus pneumoniae Danish serotype 16F DNA
C4483274|T201|COMP|85760-7|LNC|Streptococcus pneumoniae Danish serotype 19A DNA|Streptococcus pneumoniae Danish serotype 19A DNA
C4483276|T201|COMP|85766-4|LNC|Streptococcus sp DNA|Streptococcus sp DNA
C4483277|T201|COMP|85768-0|LNC|Streptococcus pneumoniae DNA|Streptococcus pneumoniae DNA
C4483278|T201|COMP|85769-8|LNC|Streptococcus pyogenes DNA|Streptococcus pyogenes DNA
C4483279|T201|COMP|85770-6|LNC|Acinetobacter baumannii DNA|Acinetobacter baumannii DNA
C4483280|T201|COMP|85771-4|LNC|Enterobacteriaceae DNA|Enterobacteriaceae DNA
C4483282|T201|COMP|85772-2|LNC|Enterobacter cloacae complex DNA|Enterobacter cloacae complex DNA
C4483284|T201|COMP|85773-0|LNC|Escherichia coli DNA|Escherichia coli DNA
C4483285|T201|COMP|85775-5|LNC|Enterococcus sp DNA|Enterococcus sp DNA
C4483287|T201|COMP|85778-9|LNC|Haemophilus influenzae DNA|Haemophilus influenzae DNA
C4483288|T201|COMP|85782-1|LNC|Candida glabrata DNA|Candida glabrata DNA
C4483289|T201|COMP|85783-9|LNC|Candida krusei DNA|Candida krusei DNA
C4483290|T201|COMP|85784-7|LNC|Candida parapsilosis DNA|Candida parapsilosis DNA
C4483291|T201|COMP|85785-4|LNC|Candida tropicalis DNA|Candida tropicalis DNA
C4483292|T201|COMP|85786-2|LNC|Bacterial methicillin resistance mecA gene|Bacterial methicillin resistance mecA gene
C4483293|T201|COMP|85787-0|LNC|Bacterial vancomycin resistance vanA+vanB genes|Bacterial vancomycin resistance vanA+vanB genes
C4483294|T201|COMP|85789-6|LNC|Cells.CD3+CD8+CD45RO+/100 cells.CD3|Cells.CD3+CD8+CD45RO+/100 cells.CD3
C4483297|T201|COMP|85792-0|LNC|Cells.CD3+CD4+CD45RO+|Cells.CD3+CD4+CD45RO+
C4483298|T201|COMP|85793-8|LNC|Specimen source subject|Specimen source subject
C4483302|T201|COMP|85795-3|LNC|Rubella virus E1 gene & genotype panel|Rubella virus E1 gene & genotype panel
C4483304|T201|COMP|85796-1|LNC|Rubella virus E1 gene|Rubella virus E1 gene
C4483309|T201|COMP|85801-9|LNC|Influenza virus B Yamagata lineage Ag|Influenza virus B Yamagata lineage Ag
C4483311|T201|COMP|85802-7|LNC|Influenza virus A H1 Ag|Influenza virus A H1 Ag
C4483312|T201|COMP|85803-5|LNC|Influenza virus A H3 Ag|Influenza virus A H3 Ag
C4483313|T201|COMP|85804-3|LNC|Influenza virus A H5 Ag|Influenza virus A H5 Ag
C4483315|T201|COMP|85805-0|LNC|Influenza virus A H7 Ag|Influenza virus A H7 Ag
C4483317|T201|COMP|85806-8|LNC|Measles virus RNA & N gene panel|Measles virus RNA & N gene panel
C4483323|T201|COMP|85810-0|LNC|Adenovirus serotype DNA panel|Adenovirus serotype DNA panel
C4483338|T201|COMP|85821-7|LNC|Influenza Virus B Victoria lineage Ag|Influenza Virus B Victoria lineage Ag
C4483342|T201|COMP|85823-3|LNC|Bacterial carbapenem resistance blaGES gene|Bacterial carbapenem resistance blaGES gene
C4483350|T201|COMP|85829-0|LNC|Bacterial carbapenem resistance blaSPM gene|Bacterial carbapenem resistance blaSPM gene
C4483351|T201|COMP|85830-8|LNC|Bacterial carbapenem resistance blaVIM gene|Bacterial carbapenem resistance blaVIM gene
C4483352|T201|COMP|85831-6|LNC|Bacterial beta-lactam resistance ESBL blaBEL gene|Bacterial beta-lactam resistance ESBL blaBEL gene
C4483356|T201|COMP|85833-2|LNC|Bacterial carbapenem resistance blaGIM gene|Bacterial carbapenem resistance blaGIM gene
C4483360|T201|COMP|85836-5|LNC|Bacterial beta-lactam resistance ESBL blaGES gene|Bacterial beta-lactam resistance ESBL blaGES gene
C4483363|T201|COMP|85838-1|LNC|Bacterial beta-lactam resistance ESBL blaSHV gene|Bacterial beta-lactam resistance ESBL blaSHV gene
C4483365|T201|COMP|85839-9|LNC|Bacterial beta-lactam resistance ESBL blaTEM gene|Bacterial beta-lactam resistance ESBL blaTEM gene
C4483367|T201|COMP|85840-7|LNC|Bacterial beta-lactam resistance ESBL blaVEB gene|Bacterial beta-lactam resistance ESBL blaVEB gene
C4483369|T201|COMP|85841-5|LNC|Bacterial beta-lactam resistance AmpC blaACC gene|Bacterial beta-lactam resistance AmpC blaACC gene
C4483402|T201|COMP|85904-1|LNC|Cancer pathology panel|Cancer pathology panel
C4483403|T201|COMP|85905-8|LNC|Cancer pathology panel|Cancer pathology panel
C4483415|T201|COMP|85952-0|LNC|Streptococcus pneumoniae Danish serotype 1 Ab|Streptococcus pneumoniae Danish serotype 1 Ab
C4483416|T201|COMP|85953-8|LNC|Streptococcus pneumoniae Danish serotype 1 Ab|Streptococcus pneumoniae Danish serotype 1 Ab
C4483418|T201|COMP|85955-3|LNC|Streptococcus pneumoniae Danish serotype 1 Ab.IgG|Streptococcus pneumoniae Danish serotype 1 Ab.IgG
C4483448|T201|COMP|85956-1|LNC|Streptococcus pneumoniae Danish serotype 1 Ab.IgG|Streptococcus pneumoniae Danish serotype 1 Ab.IgG
C4483449|T201|COMP|85957-9|LNC|Streptococcus pneumoniae Danish serotype 1 Ab.IgG|Streptococcus pneumoniae Danish serotype 1 Ab.IgG
C4483460|T201|COMP|85971-0|LNC|Streptococcus pneumoniae Danish serotype 12F Ab|Streptococcus pneumoniae Danish serotype 12F Ab
C4483461|T201|COMP|85972-8|LNC|Streptococcus pneumoniae Danish serotype 12F Ab|Streptococcus pneumoniae Danish serotype 12F Ab
C4483470|T201|COMP|85989-2|LNC|Streptococcus pneumoniae Danish serotype 14 Ab|Streptococcus pneumoniae Danish serotype 14 Ab
C4483496|T201|COMP|86020-5|LNC|Streptococcus pneumoniae Danish serotype 19F Ab|Streptococcus pneumoniae Danish serotype 19F Ab
C4483506|T201|COMP|86038-7|LNC|Streptococcus pneumoniae Danish serotype 2 Ab.IgG|Streptococcus pneumoniae Danish serotype 2 Ab.IgG
C4483508|T201|COMP|86039-5|LNC|Streptococcus pneumoniae Danish serotype 2 Ab.IgG|Streptococcus pneumoniae Danish serotype 2 Ab.IgG
C4483524|T201|COMP|86059-3|LNC|Streptococcus pneumoniae Danish serotype 23F Ab|Streptococcus pneumoniae Danish serotype 23F Ab
C4483525|T201|COMP|86060-1|LNC|Streptococcus pneumoniae Danish serotype 23F Ab|Streptococcus pneumoniae Danish serotype 23F Ab
C4483539|T201|COMP|86078-3|LNC|Streptococcus pneumoniae Danish serotype 3 Ab|Streptococcus pneumoniae Danish serotype 3 Ab
C4483541|T201|COMP|86080-9|LNC|Streptococcus pneumoniae Danish serotype 3 Ab.IgG|Streptococcus pneumoniae Danish serotype 3 Ab.IgG
C4483543|T201|COMP|86081-7|LNC|Streptococcus pneumoniae Danish serotype 3 Ab.IgG|Streptococcus pneumoniae Danish serotype 3 Ab.IgG
C4483544|T201|COMP|86082-5|LNC|Streptococcus pneumoniae Danish serotype 3 Ab.IgG|Streptococcus pneumoniae Danish serotype 3 Ab.IgG
C4483545|T201|COMP|86083-3|LNC|Streptococcus pneumoniae Danish serotype 3 Ab.IgG|Streptococcus pneumoniae Danish serotype 3 Ab.IgG
C4483562|T201|COMP|86105-4|LNC|Streptococcus pneumoniae Danish serotype 4 Ab|Streptococcus pneumoniae Danish serotype 4 Ab
C4483564|T201|COMP|86106-2|LNC|Streptococcus pneumoniae Danish serotype 4 Ab|Streptococcus pneumoniae Danish serotype 4 Ab
C4483566|T201|COMP|86109-6|LNC|Streptococcus pneumoniae Danish serotype 4 Ab.IgG|Streptococcus pneumoniae Danish serotype 4 Ab.IgG
C4483569|T201|COMP|86222-7|LNC|Lipoprotein.alpha 3|Lipoprotein.alpha 3
C4483571|T201|COMP|86223-5|LNC|Acetyl norfentanyl|Acetyl norfentanyl
C4483573|T201|COMP|86224-3|LNC|ALPRAZolam/Creatinine|ALPRAZolam/Creatinine
C4483575|T201|COMP|86225-0|LNC|clonazePAM/Creatinine|clonazePAM/Creatinine
C4483577|T201|COMP|86227-6|LNC|Dihydrocodeine|Dihydrocodeine
C4483587|T201|COMP|86502-2|LNC|Varicella zoster virus strain DNA|Varicella zoster virus strain DNA
C4483588|T201|COMP|86503-0|LNC|Streptococcus pneumoniae serotype DNA|Streptococcus pneumoniae serotype DNA
C4483590|T201|COMP|86516-2|LNC|Coxsackievirus A Ab|Coxsackievirus A Ab
C4483591|T201|COMP|86518-8|LNC|Ebola virus RNA|Ebola virus RNA
C4483592|T201|COMP|86519-6|LNC|European tick borne encephalitis virus RNA|European tick borne encephalitis virus RNA
C4483598|T201|COMP|86715-0|LNC|Actinobacillus pleuropneumoniae Ab|Actinobacillus pleuropneumoniae Ab
C4483600|T201|COMP|86717-6|LNC|Actinobacillus pleuropneumoniae serotype 1 Ab|Actinobacillus pleuropneumoniae serotype 1 Ab
C4483601|T201|COMP|86719-2|LNC|Actinobacillus pleuropneumoniae serotype 5 Ab|Actinobacillus pleuropneumoniae serotype 5 Ab
C4483615|T201|COMP|86129-4|LNC|Streptococcus pneumoniae Danish serotype 5 Ab.IgG|Streptococcus pneumoniae Danish serotype 5 Ab.IgG
C4483627|T201|COMP|86143-5|LNC|Streptococcus pneumoniae Danish serotype 8 Ab|Streptococcus pneumoniae Danish serotype 8 Ab
C4483628|T201|COMP|86144-3|LNC|Streptococcus pneumoniae Danish serotype 8 Ab|Streptococcus pneumoniae Danish serotype 8 Ab
C4483629|T201|COMP|86145-0|LNC|Streptococcus pneumoniae Danish serotype 8 Ab|Streptococcus pneumoniae Danish serotype 8 Ab
C4483630|T201|COMP|86146-8|LNC|Streptococcus pneumoniae Danish serotype 8 Ab|Streptococcus pneumoniae Danish serotype 8 Ab
C4483631|T201|COMP|86147-6|LNC|Streptococcus pneumoniae Danish serotype 8 Ab.IgG|Streptococcus pneumoniae Danish serotype 8 Ab.IgG
C4483633|T201|COMP|86148-4|LNC|Streptococcus pneumoniae Danish serotype 8 Ab.IgG|Streptococcus pneumoniae Danish serotype 8 Ab.IgG
C4483634|T201|COMP|86149-2|LNC|Streptococcus pneumoniae Danish serotype 8 Ab.IgG|Streptococcus pneumoniae Danish serotype 8 Ab.IgG
C4483643|T201|COMP|86162-5|LNC|Streptococcus pneumoniae Danish serotype 9N Ab|Streptococcus pneumoniae Danish serotype 9N Ab
C4483645|T201|COMP|86164-1|LNC|Streptococcus pneumoniae Danish serotype 9N Ab|Streptococcus pneumoniae Danish serotype 9N Ab
C4483662|T201|COMP|86190-6|LNC|Zika virus RNA|Zika virus RNA
C4483664|T201|COMP|86192-2|LNC|4-Methylethcathinone|4-Methylethcathinone
C4483665|T201|COMP|86193-0|LNC|Pentedrone|Pentedrone
C4483666|T201|COMP|86194-8|LNC|3,4-Dimethylmethcathinone|3,4-Dimethylmethcathinone
C4483667|T201|COMP|86195-5|LNC|4-Ethylmethcathinone|4-Ethylmethcathinone
C4483669|T201|COMP|86196-3|LNC|Alpha pyrrolidinovalerophenone|Alpha pyrrolidinovalerophenone
C4483671|T201|COMP|86199-7|LNC|Rotavirus A Ag|Rotavirus A Ag
C4483674|T201|COMP|86202-9|LNC|Porcine epidemic diarrhea virus|Porcine epidemic diarrhea virus
C4483675|T201|COMP|86203-7|LNC|Lawsonia intracellularis Ag|Lawsonia intracellularis Ag
C4483677|T201|COMP|86204-5|LNC|Porcine deltacoronavirus|Porcine deltacoronavirus
C4483678|T201|COMP|86205-2|LNC|Whole exome sequence analysis|Whole exome sequence analysis
C4483679|T201|COMP|86206-0|LNC|Whole genome sequence analysis|Whole genome sequence analysis
C4483707|T201|COMP|86509-7|LNC|Varicella zoster virus clade|Varicella zoster virus clade
C4483709|T201|COMP|86510-5|LNC|Adenovirus DNA|Adenovirus DNA
C4483710|T201|COMP|86511-3|LNC|Adenovirus DNA|Adenovirus DNA
C4483711|T201|COMP|86512-1|LNC|Adenovirus DNA|Adenovirus DNA
C4483712|T201|COMP|86513-9|LNC|Adenovirus Ab.IgM|Adenovirus Ab.IgM
C4483713|T201|COMP|86514-7|LNC|Chikungunya virus RNA|Chikungunya virus RNA
C4483722|T201|COMP|86216-9|LNC|Porcine epidemic diarrhea virus Ab.Neut|Porcine epidemic diarrhea virus Ab.Neut
C4483725|T201|COMP|86218-5|LNC|Transmissible gastroenteritis virus RNA|Transmissible gastroenteritis virus RNA
C4483726|T201|COMP|86220-1|LNC|Bacterial carbapenem resistance blaOXA-48 gene|Bacterial carbapenem resistance blaOXA-48 gene
C4483728|T201|COMP|86229-2|LNC|HYDROcodone|HYDROcodone
C4483729|T201|COMP|86230-0|LNC|HYDROmorphone|HYDROmorphone
C4483730|T201|COMP|86231-8|LNC|Midazolam/Creatinine|Midazolam/Creatinine
C4483732|T201|COMP|86232-6|LNC|Norsufentanil|Norsufentanil
C4483733|T201|COMP|86233-4|LNC|HIV 1 Ab|HIV 1 Ab
C4483735|T201|COMP|86235-9|LNC|Neisseria meningitidis serogroup B synD gene|Neisseria meningitidis serogroup B synD gene
C4483738|T201|COMP|86237-5|LNC|Neisseria meningitidis serogroup w135 synG gene|Neisseria meningitidis serogroup w135 synG gene
C4483739|T201|COMP|86238-3|LNC|Neisseria meningitidis serogroup X xcbB gene|Neisseria meningitidis serogroup X xcbB gene
C4483741|T201|COMP|86239-1|LNC|Cells.chromosome 3 monosomy/cells counted|Cells.chromosome 3 monosomy/cells counted
C4483743|T201|COMP|86240-9|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C4483744|T201|COMP|86241-7|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C4483745|T201|COMP|86242-5|LNC|Color|Color
C4483756|T201|COMP|86285-4|LNC|Erythrocyte deformability|Erythrocyte deformability
C4483779|T201|COMP|86316-7|LNC|Human RNase P RNA|Human RNase P RNA
C4483780|T201|COMP|86318-3|LNC|Influenza Virus B Yamagata lineage Ag|Influenza Virus B Yamagata lineage Ag
C4483781|T201|COMP|86320-9|LNC|Zika virus Ab.Neut|Zika virus Ab.Neut
C4483782|T201|COMP|86321-7|LNC|Zika virus Ab.Neut|Zika virus Ab.Neut
C4483783|T201|COMP|86322-5|LNC|Enterovirus|Enterovirus
C4483784|T201|COMP|86323-3|LNC|Enterovirus Ag|Enterovirus Ag
C4483785|T201|COMP|86324-1|LNC|Coliform bacteria|Coliform bacteria
C4483787|T201|COMP|86326-6|LNC|Bordetella holmesii hIS1001 DNA|Bordetella holmesii hIS1001 DNA
C4483791|T201|COMP|86329-0|LNC|Adenovirus 16 DNA|Adenovirus 16 DNA
C4483793|T201|COMP|86330-8|LNC|Adenovirus 11 DNA|Adenovirus 11 DNA
C4483795|T201|COMP|86331-6|LNC|Adenovirus 14 DNA|Adenovirus 14 DNA
C4483797|T201|COMP|86332-4|LNC|Adenovirus 7 DNA|Adenovirus 7 DNA
C4483799|T201|COMP|86333-2|LNC|Adenovirus 4 DNA|Adenovirus 4 DNA
C4483804|T201|COMP|86337-3|LNC|Virus identified|Virus identified
C4483805|T201|COMP|86338-1|LNC|Streptococcus pneumoniae Danish serotype 6A+6B Ab|Streptococcus pneumoniae Danish serotype 6A+6B Ab
C4483904|T201|COMP|86453-8|LNC|O-nortramadol|O-nortramadol
C4483905|T201|COMP|86454-6|LNC|N-nortramadol|N-nortramadol
C4483906|T201|COMP|86455-3|LNC|Brucella sp Ab|Brucella sp Ab
C4483907|T201|COMP|86456-1|LNC|Brucella sp Ab|Brucella sp Ab
C4483908|T201|COMP|86457-9|LNC|Brucella sp Ab|Brucella sp Ab
C4483909|T201|COMP|86459-5|LNC|Brucella sp Ab|Brucella sp Ab
C4483915|T201|COMP|86465-2|LNC|AST to platelet ratio index|AST to platelet ratio index
C4483951|T201|COMP|86520-4|LNC|Hantavirus RNA|Hantavirus RNA
C4483952|T201|COMP|86536-0|LNC|Hantavirus RNA|Hantavirus RNA
C4483953|T201|COMP|86537-8|LNC|Hantavirus RNA|Hantavirus RNA
C4483954|T201|COMP|86538-6|LNC|Hantavirus RNA|Hantavirus RNA
C4483955|T201|COMP|86539-4|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C4483956|T201|COMP|86540-2|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C4483957|T201|COMP|86541-0|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C4483958|T201|COMP|86543-6|LNC|Herpes virus 6 DNA|Herpes virus 6 DNA
C4483959|T201|COMP|86546-9|LNC|Herpes virus 8 DNA|Herpes virus 8 DNA
C4483960|T201|COMP|86547-7|LNC|HIV 2 RNA|HIV 2 RNA
C4483961|T201|COMP|86548-5|LNC|HIV 2 RNA|HIV 2 RNA
C4483962|T201|COMP|86549-3|LNC|HIV 2 RNA|HIV 2 RNA
C4483963|T201|COMP|86550-1|LNC|HTLV I+II RNA|HTLV I+II RNA
C4483975|T201|COMP|86559-2|LNC|Human bocavirus DNA|Human bocavirus DNA
C4483976|T201|COMP|86560-0|LNC|Human papilloma virus 16 DNA|Human papilloma virus 16 DNA
C4483978|T201|COMP|86562-6|LNC|Human papilloma virus 18 DNA|Human papilloma virus 18 DNA
C4483980|T201|COMP|86566-7|LNC|Influenza virus A Ab.IgG|Influenza virus A Ab.IgG
C4483981|T201|COMP|86568-3|LNC|Influenza virus A RNA|Influenza virus A RNA
C4483982|T201|COMP|86569-1|LNC|Influenza virus A RNA|Influenza virus A RNA
C4483983|T201|COMP|86570-9|LNC|Influenza virus B Ab.IgM|Influenza virus B Ab.IgM
C4483984|T201|COMP|86571-7|LNC|Influenza virus B RNA|Influenza virus B RNA
C4483985|T201|COMP|86572-5|LNC|Influenza virus B RNA|Influenza virus B RNA
C4483986|T201|COMP|86573-3|LNC|JC virus DNA|JC virus DNA
C4483987|T201|COMP|86574-1|LNC|Marburg virus RNA|Marburg virus RNA
C4483988|T201|COMP|86576-6|LNC|Measles virus RNA|Measles virus RNA
C4483989|T201|COMP|86578-2|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C4483990|T201|COMP|86579-0|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C4483991|T201|COMP|86580-8|LNC|Mumps virus RNA|Mumps virus RNA
C4483992|T201|COMP|86581-6|LNC|Neisseria meningitidis|Neisseria meningitidis
C4483993|T201|COMP|86582-4|LNC|Parechovirus A RNA|Parechovirus A RNA
C4483994|T201|COMP|86586-5|LNC|Parechovirus A RNA|Parechovirus A RNA
C4483995|T201|COMP|86587-3|LNC|Rabies virus Ab.IgG|Rabies virus Ab.IgG
C4483996|T201|COMP|86589-9|LNC|Rubella virus RNA|Rubella virus RNA
C4483997|T201|COMP|86591-5|LNC|Toscana virus RNA|Toscana virus RNA
C4483999|T201|COMP|86593-1|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C4484000|T201|COMP|86594-9|LNC|Zika virus RNA|Zika virus RNA
C4484003|T201|COMP|86604-6|LNC|Alfentanil/Creatinine|Alfentanil/Creatinine
C4484006|T201|COMP|86606-1|LNC|Cocaethylene/Creatinine|Cocaethylene/Creatinine
C4484009|T201|COMP|86608-7|LNC|Norcodeine/Creatinine|Norcodeine/Creatinine
C4484012|T201|COMP|86610-3|LNC|SUFentanil/Creatinine|SUFentanil/Creatinine
C4484014|T201|COMP|86611-1|LNC|Chromosome analysis|Chromosome analysis
C4484037|T201|COMP|86666-5|LNC|Location within lymph node|Location within lymph node
C4484042|T201|COMP|86688-9|LNC|Rotavirus C|Rotavirus C
C4484043|T201|COMP|86689-7|LNC|Rotavirus A|Rotavirus A
C4484044|T201|COMP|86690-5|LNC|Rotavirus C RNA|Rotavirus C RNA
C4484046|T201|COMP|86691-3|LNC|Rotavirus B RNA|Rotavirus B RNA
C4484048|T201|COMP|86692-1|LNC|Rotavirus A RNA|Rotavirus A RNA
C4484054|T201|COMP|86697-0|LNC|Rotavirus A RNA|Rotavirus A RNA
C4484055|T201|COMP|86698-8|LNC|Porcine epidemic diarrhea virus RNA|Porcine epidemic diarrhea virus RNA
C4484056|T201|COMP|86699-6|LNC|Rotavirus C RNA|Rotavirus C RNA
C4484057|T201|COMP|86700-2|LNC|Rotavirus C RNA|Rotavirus C RNA
C4484058|T201|COMP|86701-0|LNC|Rotavirus A RNA|Rotavirus A RNA
C4484059|T201|COMP|86702-8|LNC|Rotavirus B RNA|Rotavirus B RNA
C4484060|T201|COMP|86703-6|LNC|Porcine respiratory coronavirus RNA|Porcine respiratory coronavirus RNA
C4484063|T201|COMP|86709-3|LNC|Lawsonia intracellularis RNA|Lawsonia intracellularis RNA
C4484064|T201|COMP|86711-9|LNC|Porcine deltacoronavirus Ag|Porcine deltacoronavirus Ag
C4484066|T201|COMP|86712-7|LNC|Bacterial carbapenem resistance blaOXA gene|Bacterial carbapenem resistance blaOXA gene
C4484067|T201|COMP|86720-0|LNC|Actinobacillus pleuropneumoniae serotype 7 Ab|Actinobacillus pleuropneumoniae serotype 7 Ab
C4484070|T201|COMP|86722-6|LNC|Actinobacillus suis DNA|Actinobacillus suis DNA
C4484072|T201|COMP|86723-4|LNC|Actinobacillus suis DNA|Actinobacillus suis DNA
C4484073|T201|COMP|86724-2|LNC|Erysipelothrix rhusiopathiae|Erysipelothrix rhusiopathiae
C4484074|T201|COMP|86725-9|LNC|Erysipelothrix rhusiopathiae Ag|Erysipelothrix rhusiopathiae Ag
C4484076|T201|COMP|86727-5|LNC|Erysipelothrix sp strain 2 DNA|Erysipelothrix sp strain 2 DNA
C4484078|T201|COMP|86728-3|LNC|Erysipelothrix tonsillarum DNA|Erysipelothrix tonsillarum DNA
C4484080|T201|COMP|86729-1|LNC|Haemophilus parasuis DNA|Haemophilus parasuis DNA
C4484084|T201|COMP|86731-7|LNC|Leptospira sp DNA|Leptospira sp DNA
C4484085|T201|COMP|86733-3|LNC|Porcine parvovirus|Porcine parvovirus
C4484086|T201|COMP|86735-8|LNC|Porcine parvovirus DNA|Porcine parvovirus DNA
C4484088|T201|COMP|86736-6|LNC|Porcine parvovirus type 1 DNA|Porcine parvovirus type 1 DNA
C4484090|T201|COMP|86737-4|LNC|Toxoplasma gondii Ag|Toxoplasma gondii Ag
C4484092|T201|COMP|86738-2|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C4484093|T201|COMP|86739-0|LNC|Streptococcus suis DNA|Streptococcus suis DNA
C4484095|T201|COMP|86740-8|LNC|Streptococcus suis Ag|Streptococcus suis Ag
C4484096|T201|COMP|86741-6|LNC|Porcine parvovirus type 2 DNA|Porcine parvovirus type 2 DNA
C4484098|T201|COMP|86743-2|LNC|Surgical margin tumor involvement.deep|Surgical margin tumor involvement.deep
C4484108|T201|COMP|86857-0|LNC|Flavivirus Ab.Neut|Flavivirus Ab.Neut
C4484110|T201|COMP|86858-8|LNC|Dengue virus 2 Ab.Neut|Dengue virus 2 Ab.Neut
C4484112|T201|COMP|86859-6|LNC|Dengue virus 3 Ab.Neut|Dengue virus 3 Ab.Neut
C4484115|T201|COMP|86861-2|LNC|Dengue virus 4 Ab.Neut|Dengue virus 4 Ab.Neut
C4484116|T201|COMP|86862-0|LNC|Dengue virus 4 Ab.Neut|Dengue virus 4 Ab.Neut
C4484117|T201|COMP|86863-8|LNC|Dengue virus 3 Ab.Neut|Dengue virus 3 Ab.Neut
C4484118|T201|COMP|86864-6|LNC|Dengue virus 2 Ab.Neut|Dengue virus 2 Ab.Neut
C4484119|T201|COMP|86865-3|LNC|Dengue virus 1 Ab.Neut|Dengue virus 1 Ab.Neut
C4521405|T201|COMP|87527-8|LNC|Fasting duration|Fasting duration
C4521427|T201|COMP|87623-5|LNC|HEDIS 2018 Value Set - Depression Screen|HEDIS 2018 Value Set - Depression Screen
C4522082|T201|COMP|87396-8|LNC|GenBank accession number|GenBank accession number
C4522117|T201|COMP|86504-8|LNC|These questions three panel|These questions three panel
C4522179|T201|COMP|87625-0|LNC|HEDIS 2018 Value Sets|HEDIS 2018 Value Sets
C4531425|T201|COMP|85039-6|LNC|JAK2 gene.p.Val617Phe mutant/normal|JAK2 gene.p.Val617Phe mutant/normal
C4531492|T201|COMP|86895-0|LNC|Adalimumab Ab|Adalimumab Ab
C4531493|T201|COMP|86896-8|LNC|inFLIXimab|inFLIXimab
C4531494|T201|COMP|86897-6|LNC|inFLIXimab Ab|inFLIXimab Ab
C4531495|T201|COMP|86898-4|LNC|Vedolizumab|Vedolizumab
C4531496|T201|COMP|86899-2|LNC|Vedolizumab Ab|Vedolizumab Ab
C4531898|T201|COMP|86894-3|LNC|Adalimumab|Adalimumab
C4531899|T201|COMP|86900-8|LNC|Plasma cells.monotypic population|Plasma cells.monotypic population
C4531938|T201|COMP|86925-5|LNC|Lawsonia intracellularis Ab|Lawsonia intracellularis Ab
C4531943|T201|COMP|86928-9|LNC|Porcine epidemic diarrhea virus whole genome|Porcine epidemic diarrhea virus whole genome
C4531945|T201|COMP|86929-7|LNC|Lawsonia intracellularis Ab/Negative control|Lawsonia intracellularis Ab/Negative control
C4531947|T201|COMP|86930-5|LNC|Carbapenemase|Carbapenemase
C4531948|T201|COMP|86931-3|LNC|Metanephrine, Normetanephrine & Creatinine panel|Metanephrine, Normetanephrine & Creatinine panel
C4531981|T201|COMP|86950-3|LNC|Thymus Ab.IgG|Thymus Ab.IgG
C4531983|T201|COMP|86951-1|LNC|Lipoprotein associated phospholipase A2|Lipoprotein associated phospholipase A2
C4531988|T201|COMP|86954-5|LNC|Foreign material|Foreign material
C4532113|T201|COMP|87570-8|LNC|Narasin|Narasin
C4532114|T201|COMP|87571-6|LNC|Fumonisin B3|Fumonisin B3
C4532115|T201|COMP|87572-4|LNC|Fumonisin B2|Fumonisin B2
C4532116|T201|COMP|87573-2|LNC|Fumonisin B1|Fumonisin B1
C4532117|T201|COMP|87574-0|LNC|Ergovaline|Ergovaline
C4532118|T201|COMP|87575-7|LNC|Ergotamine|Ergotamine
C4532119|T201|COMP|87576-5|LNC|Ergosine|Ergosine
C4532120|T201|COMP|87577-3|LNC|Ergocryptine|Ergocryptine
C4532121|T201|COMP|87578-1|LNC|Ergocristine|Ergocristine
C4532122|T201|COMP|87663-1|LNC|Disulfoton|Disulfoton
C4532123|T201|COMP|87664-9|LNC|Dimethoate|Dimethoate
C4532124|T201|COMP|87665-6|LNC|Dieldrin|Dieldrin
C4532125|T201|COMP|87666-4|LNC|Diazinon|Diazinon
C4532126|T201|COMP|87667-2|LNC|Alpha benzene hexachloride|Alpha benzene hexachloride
C4532128|T201|COMP|87668-0|LNC|Aldrin|Aldrin
C4532129|T201|COMP|87669-8|LNC|Chlorinated hydrocarbon panel|Chlorinated hydrocarbon panel
C4532131|T201|COMP|87670-6|LNC|Carbamate panel|Carbamate panel
C4532133|T201|COMP|87671-4|LNC|Cholecalciferol|Cholecalciferol
C4532134|T201|COMP|87672-2|LNC|Tocopherol+tocotrienol|Tocopherol+tocotrienol
C4532139|T201|COMP|87708-4|LNC|Beta-2-Microglobulin^post dialysis|Beta-2-Microglobulin^post dialysis
C4532140|T201|COMP|87709-2|LNC|Virus identified|Virus identified
C4532213|T201|COMP|87321-6|LNC|Escherichia coli enterotoxigenic sta gene|Escherichia coli enterotoxigenic sta gene
C4532215|T201|COMP|87322-4|LNC|Escherichia coli enterotoxigenic stb gene|Escherichia coli enterotoxigenic stb gene
C4532217|T201|COMP|87323-2|LNC|Porcine circovirus type 1 DNA|Porcine circovirus type 1 DNA
C4532219|T201|COMP|87379-4|LNC|Cannabinol|Cannabinol
C4532220|T201|COMP|87380-2|LNC|Escherichia coli Stx2e toxin stx2e gene|Escherichia coli Stx2e toxin stx2e gene
C4532222|T201|COMP|87381-0|LNC|Porcine Adenovirus Ab|Porcine Adenovirus Ab
C4532223|T201|COMP|87382-8|LNC|Porcine cytomegalovirus DNA|Porcine cytomegalovirus DNA
C4532227|T201|COMP|87429-7|LNC|Cortisol AM & PM panel|Cortisol AM & PM panel
C4532231|T201|COMP|87431-3|LNC|Herpes simplex virus 1 & 2 DNA panel|Herpes simplex virus 1 & 2 DNA panel
C4532232|T201|COMP|87432-1|LNC|Mycophenolate & mycophenolate glucuronide panel|Mycophenolate & mycophenolate glucuronide panel
C4532234|T201|COMP|87486-7|LNC|PB-22 3-carboxyindole|PB-22 3-carboxyindole
C4532236|T201|COMP|87487-5|LNC|MAB-CHMINACA butanoate|MAB-CHMINACA butanoate
C4532238|T201|COMP|87488-3|LNC|AM694 N-5-hydroxypentyl|AM694 N-5-hydroxypentyl
C4532240|T201|COMP|87489-1|LNC|AKB48 N-pentanoate|AKB48 N-pentanoate
C4532242|T201|COMP|87490-9|LNC|ADB-PINACA pentanoate|ADB-PINACA pentanoate
C4532244|T201|COMP|87491-7|LNC|ADBICA N-4-hydroxypentyl|ADBICA N-4-hydroxypentyl
C4532246|T201|COMP|87492-5|LNC|AB-PINACA pentanoate|AB-PINACA pentanoate
C4532248|T201|COMP|87493-3|LNC|AB-FUBINACA oxobutanoate|AB-FUBINACA oxobutanoate
C4532250|T201|COMP|87550-0|LNC|Haloperidol & haloperidol.reduced panel|Haloperidol & haloperidol.reduced panel
C4532254|T201|COMP|87552-6|LNC|IgA & IgA subclass 1 & IgA subclass 2 panel|IgA & IgA subclass 1 & IgA subclass 2 panel
C4532268|T201|COMP|87305-9|LNC|Clostridium perfringens cpb2 gene|Clostridium perfringens cpb2 gene
C4532270|T201|COMP|87306-7|LNC|Clostridium perfringens cpe gene|Clostridium perfringens cpe gene
C4532272|T201|COMP|87307-5|LNC|Clostridium perfringens etx gene|Clostridium perfringens etx gene
C4532280|T201|COMP|87390-1|LNC|Porcine sapelovirus RNA|Porcine sapelovirus RNA
C4532282|T201|COMP|87391-9|LNC|Porcine teschovirus RNA|Porcine teschovirus RNA
C4532284|T201|COMP|87392-7|LNC|Porcine teschovirus RNA|Porcine teschovirus RNA
C4532285|T201|COMP|87393-5|LNC|Salmonella sp Ab/Positive control|Salmonella sp Ab/Positive control
C4532287|T201|COMP|87394-3|LNC|Salmonella sp DNA|Salmonella sp DNA
C4532288|T201|COMP|87395-0|LNC|West Nile virus RNA|West Nile virus RNA
C4532289|T201|COMP|87941-1|LNC|Bacteria identified|Bacteria identified
C4532290|T201|COMP|87942-9|LNC|Bacteria identified|Bacteria identified
C4532291|T201|COMP|87943-7|LNC|Bacteria identified|Bacteria identified
C4532292|T201|COMP|87944-5|LNC|Bacteria identified|Bacteria identified
C4532293|T201|COMP|87945-2|LNC|Borrelia sp identified|Borrelia sp identified
C4532294|T201|COMP|87946-0|LNC|Borrelia sp identified|Borrelia sp identified
C4532295|T201|COMP|87947-8|LNC|Borrelia sp DNA|Borrelia sp DNA
C4532296|T201|COMP|87948-6|LNC|Clostridium botulinum|Clostridium botulinum
C4532482|T201|COMP|87241-6|LNC|Bacillus atrophaeus|Bacillus atrophaeus
C4532483|T201|COMP|87242-4|LNC|Geobacillus stearothermophilus|Geobacillus stearothermophilus
C4532505|T201|COMP|87275-4|LNC|Borrelia afzelii+burgdorferi+garinii Ab.IgG|Borrelia afzelii+burgdorferi+garinii Ab.IgG
C4532509|T201|COMP|87277-0|LNC|Borrelia afzelii+burgdorferi+garinii Ab.IgM|Borrelia afzelii+burgdorferi+garinii Ab.IgM
C4532517|T201|COMP|87282-0|LNC|Brachyspira hyodysenteriae DNA|Brachyspira hyodysenteriae DNA
C4532519|T201|COMP|87283-8|LNC|Brachyspira hampsonii DNA|Brachyspira hampsonii DNA
C4532521|T201|COMP|87284-6|LNC|Brachyspira hyodysenteriae DNA|Brachyspira hyodysenteriae DNA
C4532522|T201|COMP|87285-3|LNC|Brachyspira pilosicoli DNA|Brachyspira pilosicoli DNA
C4532543|T201|COMP|87304-2|LNC|Clostridium perfringens cpa gene|Clostridium perfringens cpa gene
C4532549|T201|COMP|87313-3|LNC|Clostridium perfringens iota toxin DNA|Clostridium perfringens iota toxin DNA
C4532551|T201|COMP|87314-1|LNC|Encephalomyocarditis virus|Encephalomyocarditis virus
C4532552|T201|COMP|87315-8|LNC|Encephalomyocarditis virus RNA|Encephalomyocarditis virus RNA
C4532554|T201|COMP|87316-6|LNC|Enterovirus G RNA|Enterovirus G RNA
C4532556|T201|COMP|87317-4|LNC|Escherichia coli|Escherichia coli
C4532557|T201|COMP|87318-2|LNC|Escherichia coli eaeA gene|Escherichia coli eaeA gene
C4532558|T201|COMP|87319-0|LNC|Escherichia coli enteroaggregative astA gene|Escherichia coli enteroaggregative astA gene
C4532560|T201|COMP|87324-0|LNC|Porcine circovirus type 2|Porcine circovirus type 2
C4532561|T201|COMP|87325-7|LNC|Porcine circovirus type 2 Ab|Porcine circovirus type 2 Ab
C4532563|T201|COMP|87326-5|LNC|Porcine circovirus type 2 Ab.IgG|Porcine circovirus type 2 Ab.IgG
C4532565|T201|COMP|87327-3|LNC|Porcine circovirus type 2 Ab.IgG+IgM|Porcine circovirus type 2 Ab.IgG+IgM
C4532567|T201|COMP|87328-1|LNC|Porcine circovirus type 2 Ab.IgG+IgM|Porcine circovirus type 2 Ab.IgG+IgM
C4532568|T201|COMP|87329-9|LNC|Porcine circovirus type 2 Ab.IgG/Positive control|Porcine circovirus type 2 Ab.IgG/Positive control
C4532570|T201|COMP|87330-7|LNC|Porcine Circovirus type 2 Ab.Neut|Porcine Circovirus type 2 Ab.Neut
C4532572|T201|COMP|87331-5|LNC|Porcine circovirus type 2 Ab/Negative control|Porcine circovirus type 2 Ab/Negative control
C4532574|T201|COMP|87332-3|LNC|Porcine circovirus type 2 Ag|Porcine circovirus type 2 Ag
C4532576|T201|COMP|87334-9|LNC|Porcine circovirus type 2 DNA|Porcine circovirus type 2 DNA
C4532578|T201|COMP|87335-6|LNC|Porcine circovirus type 2 DNA|Porcine circovirus type 2 DNA
C4532579|T201|COMP|87336-4|LNC|Porcine circovirus type 2 DNA|Porcine circovirus type 2 DNA
C4532580|T201|COMP|87337-2|LNC|Porcine circovirus type 2 RFLP pattern|Porcine circovirus type 2 RFLP pattern
C4532582|T201|COMP|87338-0|LNC|Porcine circovirus type 2 strain identified|Porcine circovirus type 2 strain identified
C4532584|T201|COMP|87339-8|LNC|Porcine circovirus type 2a DNA|Porcine circovirus type 2a DNA
C4532586|T201|COMP|87340-6|LNC|Porcine circovirus type 2b DNA|Porcine circovirus type 2b DNA
C4532588|T201|COMP|87341-4|LNC|Pseudorabies virus|Pseudorabies virus
C4532589|T201|COMP|87342-2|LNC|Pseudorabies virus DNA|Pseudorabies virus DNA
C4532594|T201|COMP|87345-5|LNC|Senecavirus A|Senecavirus A
C4532595|T201|COMP|87346-3|LNC|Senecavirus A Ab|Senecavirus A Ab
C4532597|T201|COMP|87347-1|LNC|Senecavirus A Ab.IgG/Positive control|Senecavirus A Ab.IgG/Positive control
C4532599|T201|COMP|87348-9|LNC|Senecavirus A RNA|Senecavirus A RNA
C4532601|T201|COMP|87350-5|LNC|Senecavirus A RNA|Senecavirus A RNA
C4532602|T201|COMP|87351-3|LNC|Senecavirus A RNA|Senecavirus A RNA
C4532603|T201|COMP|87352-1|LNC|Senecavirus A whole genome|Senecavirus A whole genome
C4532621|T201|COMP|87361-2|LNC|Toxoplasma gondii Ab/Negative control|Toxoplasma gondii Ab/Negative control
C4532627|T201|COMP|87364-6|LNC|Haemophilus parasuis Ab/Positive control|Haemophilus parasuis Ab/Positive control
C4532633|T201|COMP|87367-9|LNC|Erysipelothrix rhusiopathiae Ab/Positive control|Erysipelothrix rhusiopathiae Ab/Positive control
C4532637|T201|COMP|87369-5|LNC|Lawsonia intracellularis VNTR pattern|Lawsonia intracellularis VNTR pattern
C4532639|T201|COMP|87370-3|LNC|Escherichia coli fasA gene|Escherichia coli fasA gene
C4532641|T201|COMP|87371-1|LNC|Escherichia coli fedF gene|Escherichia coli fedF gene
C4532643|T201|COMP|87372-9|LNC|Escherichia coli FimF41a gene|Escherichia coli FimF41a gene
C4532645|T201|COMP|87373-7|LNC|Escherichia coli K88 DNA|Escherichia coli K88 DNA
C4532647|T201|COMP|87374-5|LNC|Escherichia coli K99 DNA|Escherichia coli K99 DNA
C4532649|T201|COMP|87375-2|LNC|Escherichia coli paa gene|Escherichia coli paa gene
C4532651|T201|COMP|87376-0|LNC|Escherichia coli Stx1 toxin stx1 gene|Escherichia coli Stx1 toxin stx1 gene
C4532653|T201|COMP|87377-8|LNC|Escherichia coli Stx2 toxin stx2 gene|Escherichia coli Stx2 toxin stx2 gene
C4532655|T201|COMP|87378-6|LNC|Tubular extraction rate/1.73 sq M|Tubular extraction rate/1.73 sq M
C4532657|T201|COMP|87384-4|LNC|Porcine parainfluenza virus 1 HN gene|Porcine parainfluenza virus 1 HN gene
C4532659|T201|COMP|87385-1|LNC|Porcine parainfluenza virus 1 F gene|Porcine parainfluenza virus 1 F gene
C4532661|T201|COMP|87386-9|LNC|Porcine parainfluenza virus 1 RNA|Porcine parainfluenza virus 1 RNA
C4532663|T201|COMP|87387-7|LNC|Porcine parainfluenza virus 1 RNA|Porcine parainfluenza virus 1 RNA
C4532664|T201|COMP|87388-5|LNC|Porcine sapelovirus|Porcine sapelovirus
C4532665|T201|COMP|87389-3|LNC|Porcine sapelovirus RNA|Porcine sapelovirus RNA
C4532666|T201|COMP|87397-6|LNC|Clostridium perfringens cpb gene|Clostridium perfringens cpb gene
C4532668|T201|COMP|87398-4|LNC|Brachyspira sp DNA|Brachyspira sp DNA
C4532670|T201|COMP|87399-2|LNC|Porcine teschovirus|Porcine teschovirus
C4532671|T201|COMP|87400-8|LNC|Brachyspira sp Ag|Brachyspira sp Ag
C4532673|T201|COMP|87401-6|LNC|Brachyspira pilosicoli DNA|Brachyspira pilosicoli DNA
C4532674|T201|COMP|87402-4|LNC|Escherichia coli aidA-I gene|Escherichia coli aidA-I gene
C4532676|T201|COMP|87403-2|LNC|Platelet aggregation.ristocetin induced^750 ug/mL|Platelet aggregation.ristocetin induced^750 ug/mL
C4532677|T201|COMP|87404-0|LNC|Certolizumab|Certolizumab
C4532678|T201|COMP|87405-7|LNC|Certolizumab Ab|Certolizumab Ab
C4532680|T201|COMP|87406-5|LNC|Golimumab|Golimumab
C4532681|T201|COMP|87407-3|LNC|Golimumab Ab|Golimumab Ab
C4532683|T201|COMP|87408-1|LNC|Ustekinumab|Ustekinumab
C4532684|T201|COMP|87409-9|LNC|Ustekinumab Ab|Ustekinumab Ab
C4532686|T201|COMP|87410-7|LNC|Thymidine synthase activity interpretation|Thymidine synthase activity interpretation
C4532688|T201|COMP|87411-5|LNC|Brachyspira hyodysenteriae DNA|Brachyspira hyodysenteriae DNA
C4532689|T201|COMP|87412-3|LNC|Brachyspira sp nox gene|Brachyspira sp nox gene
C4532691|T201|COMP|87413-1|LNC|Brachyspira sp|Brachyspira sp
C4532696|T201|COMP|87417-2|LNC|Cytolethal distending toxin B & Vinculin Ab panel|Cytolethal distending toxin B & Vinculin Ab panel
C4532698|T201|COMP|87418-0|LNC|Cytolethal distending toxin B Ab|Cytolethal distending toxin B Ab
C4532700|T201|COMP|87419-8|LNC|Cytolethal distending toxin B+Vinculin Ab|Cytolethal distending toxin B+Vinculin Ab
C4532702|T201|COMP|87420-6|LNC|Vinculin Ab|Vinculin Ab
C4532703|T201|COMP|87421-4|LNC|Glucose^pre-meal|Glucose^pre-meal
C4532704|T201|COMP|87422-2|LNC|Glucose^post meal|Glucose^post meal
C4532705|T201|COMP|87423-0|LNC|Borrelia burgdorferi Ab.IgG & IgM panel|Borrelia burgdorferi Ab.IgG & IgM panel
C4532706|T201|COMP|87424-8|LNC|Cytomegalovirus Ab.IgG & IgM Panel|Cytomegalovirus Ab.IgG & IgM Panel
C4532707|T201|COMP|87426-3|LNC|Inhibin A & B panel|Inhibin A & B panel
C4532709|T201|COMP|87427-1|LNC|Neutrophil cytoplasmic Ab panel|Neutrophil cytoplasmic Ab panel
C4532711|T201|COMP|87428-9|LNC|Drugs of abuse screen W Reflex confirm panel|Drugs of abuse screen W Reflex confirm panel
C4532713|T201|COMP|87433-9|LNC|Hemoglobin.free & oxyhemoglobin panel|Hemoglobin.free & oxyhemoglobin panel
C4532715|T201|COMP|87434-7|LNC|Protein & creatinine panel|Protein & creatinine panel
C4532717|T201|COMP|87435-4|LNC|Coccidioides immitis Ab.IgG & IgM panel|Coccidioides immitis Ab.IgG & IgM panel
C4532719|T201|COMP|87436-2|LNC|Chromosome X & Y aneuploidy|Chromosome X & Y aneuploidy
C4532720|T201|COMP|87437-0|LNC|Oxyhemoglobin|Oxyhemoglobin
C4532721|T201|COMP|87438-8|LNC|Dengue virus 1+2+3+4 & Zika virus Ab.IgA+IgG+IgM|Dengue virus 1+2+3+4 & Zika virus Ab.IgA+IgG+IgM
C4532723|T201|COMP|87439-6|LNC|Zika virus Ab.IgA+IgG+IgM|Zika virus Ab.IgA+IgG+IgM
C4532725|T201|COMP|87440-4|LNC|Dengue virus 1+2+3+4 Ab.IgA+IgG+IgM|Dengue virus 1+2+3+4 Ab.IgA+IgG+IgM
C4532729|T201|COMP|87442-0|LNC|Turbidity|Turbidity
C4532730|T201|COMP|87443-8|LNC|Hardness|Hardness
C4532731|T201|COMP|87444-6|LNC|Electrical conductivity|Electrical conductivity
C4532732|T201|COMP|87445-3|LNC|Fungus|Fungus
C4532733|T201|COMP|87446-1|LNC|Zinc|Zinc
C4532734|T201|COMP|87447-9|LNC|Vanadium|Vanadium
C4532735|T201|COMP|87448-7|LNC|Vanadium|Vanadium
C4532736|T201|COMP|87449-5|LNC|Sulfur|Sulfur
C4532737|T201|COMP|87450-3|LNC|Sulfur|Sulfur
C4532738|T201|COMP|87451-1|LNC|Sodium|Sodium
C4532739|T201|COMP|87452-9|LNC|Sodium|Sodium
C4532740|T201|COMP|87453-7|LNC|Selenium|Selenium
C4532741|T201|COMP|87454-5|LNC|Potassium|Potassium
C4532742|T201|COMP|87455-2|LNC|Potassium|Potassium
C4532743|T201|COMP|87456-0|LNC|Phosphate|Phosphate
C4532744|T201|COMP|87457-8|LNC|Phosphate|Phosphate
C4532745|T201|COMP|87458-6|LNC|Particle diameter.mean|Particle diameter.mean
C4532747|T201|COMP|87459-4|LNC|Nitrite|Nitrite
C4532748|T201|COMP|87460-2|LNC|Nitrite|Nitrite
C4532749|T201|COMP|87461-0|LNC|Nitrate|Nitrate
C4532750|T201|COMP|87462-8|LNC|Nitrate|Nitrate
C4532751|T201|COMP|87463-6|LNC|Nickel|Nickel
C4532752|T201|COMP|87464-4|LNC|Monensin|Monensin
C4532753|T201|COMP|87465-1|LNC|Monensin|Monensin
C4532754|T201|COMP|87466-9|LNC|Molybdenum|Molybdenum
C4532755|T201|COMP|87467-7|LNC|Manganese|Manganese
C4532756|T201|COMP|87468-5|LNC|Manganese|Manganese
C4532757|T201|COMP|87469-3|LNC|Magnesium|Magnesium
C4532758|T201|COMP|87470-1|LNC|Magnesium|Magnesium
C4532759|T201|COMP|87471-9|LNC|Iron|Iron
C4532760|T201|COMP|87472-7|LNC|Copper|Copper
C4532761|T201|COMP|87473-5|LNC|Cobalt|Cobalt
C4532762|T201|COMP|87474-3|LNC|Chromium|Chromium
C4532763|T201|COMP|87475-0|LNC|Chloride|Chloride
C4532764|T201|COMP|87476-8|LNC|Chloride|Chloride
C4532765|T201|COMP|87477-6|LNC|Calcium|Calcium
C4532766|T201|COMP|87478-4|LNC|Cadmium|Cadmium
C4532767|T201|COMP|87479-2|LNC|Boron|Boron
C4532768|T201|COMP|87480-0|LNC|Bone ash/Bone.total|Bone ash/Bone.total
C4532770|T201|COMP|87481-8|LNC|Arsenic|Arsenic
C4532771|T201|COMP|87482-6|LNC|Aluminum|Aluminum
C4532772|T201|COMP|87483-4|LNC|Aluminum|Aluminum
C4532773|T201|COMP|87484-2|LNC|BB-22 3-carboxyindole|BB-22 3-carboxyindole
C4532775|T201|COMP|87485-9|LNC|ADBICA N-pentanoate|ADBICA N-pentanoate
C4532777|T201|COMP|87494-1|LNC|AB-CHMINACA hydroxycyclohexyl|AB-CHMINACA hydroxycyclohexyl
C4532779|T201|COMP|87495-8|LNC|AB-CHMINACA butanoate|AB-CHMINACA butanoate
C4532781|T201|COMP|87496-6|LNC|Gabapentin|Gabapentin
C4532782|T201|COMP|87497-4|LNC|Meperidine|Meperidine
C4532783|T201|COMP|87498-2|LNC|3-Methoxytyramine.free/Creatinine|3-Methoxytyramine.free/Creatinine
C4532785|T201|COMP|87499-0|LNC|3-Methoxytyramine.free|3-Methoxytyramine.free
C4532841|T201|COMP|87546-8|LNC|Dengue virus Ab.IgG & IgM panel|Dengue virus Ab.IgG & IgM panel
C4532850|T201|COMP|87554-2|LNC|Epstein Barr virus Ab panel|Epstein Barr virus Ab panel
C4532854|T201|COMP|87556-7|LNC|Thyroglobulin & thyroperoxidase Ab panel|Thyroglobulin & thyroperoxidase Ab panel
C4532856|T201|COMP|87557-5|LNC|Protein S Ag & protein S Ag.free panel|Protein S Ag & protein S Ag.free panel
C4532858|T201|COMP|87558-3|LNC|Anaplasma phagocytophilum groEL gene|Anaplasma phagocytophilum groEL gene
C4532860|T201|COMP|87559-1|LNC|Ehrlichia chaffeensis groEL gene|Ehrlichia chaffeensis groEL gene
C4532862|T201|COMP|87560-9|LNC|Ehrlichia canis+ewingii groEL gene|Ehrlichia canis+ewingii groEL gene
C4532864|T201|COMP|87561-7|LNC|Ehrlichia muris eauclairensis groEL gene|Ehrlichia muris eauclairensis groEL gene
C4532866|T201|COMP|87562-5|LNC|Ammonia nitrogen|Ammonia nitrogen
C4532867|T201|COMP|87563-3|LNC|Antimony|Antimony
C4532868|T201|COMP|87564-1|LNC|Zearalenone|Zearalenone
C4532869|T201|COMP|87565-8|LNC|Zearalenol|Zearalenol
C4532870|T201|COMP|87566-6|LNC|Deoxynivalenol|Deoxynivalenol
C4532871|T201|COMP|87567-4|LNC|T-2 toxin|T-2 toxin
C4532872|T201|COMP|87568-2|LNC|Ochratoxin A|Ochratoxin A
C4532873|T201|COMP|87569-0|LNC|Nivalenol|Nivalenol
C4532874|T201|COMP|87579-9|LNC|Ergocornine|Ergocornine
C4532875|T201|COMP|87580-7|LNC|Aflatoxin M1|Aflatoxin M1
C4532876|T201|COMP|87581-5|LNC|Aflatoxin G2|Aflatoxin G2
C4532877|T201|COMP|87582-3|LNC|Aflatoxin G1|Aflatoxin G1
C4532878|T201|COMP|87583-1|LNC|Aflatoxin B2|Aflatoxin B2
C4532879|T201|COMP|87584-9|LNC|Aflatoxin B1|Aflatoxin B1
C4532880|T201|COMP|87585-6|LNC|Virginiamycin|Virginiamycin
C4532881|T201|COMP|87586-4|LNC|Tylvalosin|Tylvalosin
C4532882|T201|COMP|87587-2|LNC|Tylosin|Tylosin
C4532883|T201|COMP|87588-0|LNC|Tilmicosin|Tilmicosin
C4532884|T201|COMP|87589-8|LNC|Tiamulin|Tiamulin
C4532885|T201|COMP|87590-6|LNC|Tetracycline|Tetracycline
C4532886|T201|COMP|87591-4|LNC|Sulfathiazole|Sulfathiazole
C4532887|T201|COMP|87592-2|LNC|Sulfamethazine|Sulfamethazine
C4532888|T201|COMP|87593-0|LNC|Salinomycin|Salinomycin
C4532889|T201|COMP|87594-8|LNC|Penicillin|Penicillin
C4532890|T201|COMP|87595-5|LNC|Oxytetracycline|Oxytetracycline
C4532891|T201|COMP|87596-3|LNC|Nicotine|Nicotine
C4532892|T201|COMP|87597-1|LNC|Lincomycin|Lincomycin
C4532893|T201|COMP|87598-9|LNC|Lasalocid|Lasalocid
C4532894|T201|COMP|87599-7|LNC|Florfenicol|Florfenicol
C4532895|T201|COMP|87600-3|LNC|Chlortetracycline|Chlortetracycline
C4532896|T201|COMP|87601-1|LNC|Carbadox|Carbadox
C4532897|T201|COMP|87602-9|LNC|Bambermycins|Bambermycins
C4532898|T201|COMP|87603-7|LNC|Bacitracin zinc|Bacitracin zinc
C4532899|T201|COMP|87604-5|LNC|Ampicillin|Ampicillin
C4532900|T201|COMP|87605-2|LNC|Warfarin|Warfarin
C4532901|T201|COMP|87606-0|LNC|Diphacinone|Diphacinone
C4532902|T201|COMP|87607-8|LNC|Difethialone|Difethialone
C4532903|T201|COMP|87608-6|LNC|Difenacoum|Difenacoum
C4532904|T201|COMP|87609-4|LNC|Dicoumarol|Dicoumarol
C4532905|T201|COMP|87610-2|LNC|Chlorophacinone|Chlorophacinone
C4532906|T201|COMP|87611-0|LNC|Bromadiolone|Bromadiolone
C4532907|T201|COMP|87612-8|LNC|Brodifacoum|Brodifacoum
C4532908|T201|COMP|87613-6|LNC|Urea|Urea
C4532909|T201|COMP|87614-4|LNC|Thallium|Thallium
C4532910|T201|COMP|87615-1|LNC|Sulfate|Sulfate
C4532911|T201|COMP|87616-9|LNC|Gossypol|Gossypol
C4532912|T201|COMP|87617-7|LNC|Ethylene glycol|Ethylene glycol
C4532913|T201|COMP|87618-5|LNC|Cyanide|Cyanide
C4532914|T201|COMP|87619-3|LNC|Barium|Barium
C4532915|T201|COMP|87620-1|LNC|Candida auris ITS2 gene|Candida auris ITS2 gene
C4532917|T201|COMP|87621-9|LNC|Bordetella parapertussis IS1001 DNA|Bordetella parapertussis IS1001 DNA
C4532918|T201|COMP|87622-7|LNC|Zika virus Ab.IgM|Zika virus Ab.IgM
C4532919|T201|COMP|87624-3|LNC|HEDIS 2018 Value Set - Alcohol Screening|HEDIS 2018 Value Set - Alcohol Screening
C4532924|T201|COMP|87630-0|LNC|Mevinphos|Mevinphos
C4532925|T201|COMP|87631-8|LNC|Mexacarbate|Mexacarbate
C4532926|T201|COMP|87632-6|LNC|Toxaphene|Toxaphene
C4532927|T201|COMP|87633-4|LNC|Phorate|Phorate
C4532928|T201|COMP|87634-2|LNC|Aldicarb|Aldicarb
C4532929|T201|COMP|87635-9|LNC|Aldicarb sulfone|Aldicarb sulfone
C4532930|T201|COMP|87636-7|LNC|Crufomate|Crufomate
C4532931|T201|COMP|87637-5|LNC|Fenchlorphos|Fenchlorphos
C4532932|T201|COMP|87644-1|LNC|Ethoprop|Ethoprop
C4532933|T201|COMP|87645-8|LNC|Dechlorane|Dechlorane
C4532934|T201|COMP|87646-6|LNC|Methyl parathion|Methyl parathion
C4532935|T201|COMP|87647-4|LNC|Methoxychlor|Methoxychlor
C4532936|T201|COMP|87648-2|LNC|Malathion|Malathion
C4532937|T201|COMP|87649-0|LNC|Lindane|Lindane
C4532938|T201|COMP|87650-8|LNC|Methomyl|Methomyl
C4532939|T201|COMP|87651-6|LNC|2,3,5-trimethylphenyl methylcarbamate|2,3,5-trimethylphenyl methylcarbamate
C4532941|T201|COMP|87652-4|LNC|Isofenphos|Isofenphos
C4532942|T201|COMP|87653-2|LNC|Hexachlorobenzene|Hexachlorobenzene
C4532943|T201|COMP|87654-0|LNC|Heptachlor|Heptachlor
C4532944|T201|COMP|87655-7|LNC|Heptachlor epoxide|Heptachlor epoxide
C4532945|T201|COMP|87656-5|LNC|Carbofuran|Carbofuran
C4532946|T201|COMP|87657-3|LNC|Fenthion|Fenthion
C4532947|T201|COMP|87658-1|LNC|Famphur|Famphur
C4532948|T201|COMP|87659-9|LNC|Parathion|Parathion
C4532949|T201|COMP|87660-7|LNC|Endrin|Endrin
C4532950|T201|COMP|87661-5|LNC|Endosulfan I|Endosulfan I
C4532952|T201|COMP|87662-3|LNC|Fonofos|Fonofos
C4532953|T201|COMP|87673-0|LNC|Retinal+retinol+retinoic acid|Retinal+retinol+retinoic acid
C4533007|T201|COMP|87767-0|LNC|Primidone/Creatinine|Primidone/Creatinine
C4533009|T201|COMP|87768-8|LNC|Rufinamide/Creatinine|Rufinamide/Creatinine
C4533011|T201|COMP|87769-6|LNC|tiaGABine/Creatinine|tiaGABine/Creatinine
C4533013|T201|COMP|87770-4|LNC|Topiramate/Creatinine|Topiramate/Creatinine
C4533022|T201|COMP|88129-2|LNC|Respiratory pathogens panel|Respiratory pathogens panel
C4533023|T201|COMP|88130-0|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C4533024|T201|COMP|88131-8|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C4533025|T201|COMP|88132-6|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C4533026|T201|COMP|88195-3|LNC|Influenza virus B RNA|Influenza virus B RNA
C4533027|T201|COMP|88196-1|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C4533028|T201|COMP|88197-9|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C4533029|T201|COMP|88198-7|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C4533030|T201|COMP|88258-9|LNC|Escherichia coli oppA gene|Escherichia coli oppA gene
C4533031|T201|COMP|88259-7|LNC|Gram negative bacteria identified|Gram negative bacteria identified
C4533032|T201|COMP|88260-5|LNC|Gram negative blood culture panel|Gram negative blood culture panel
C4533041|T201|COMP|87710-0|LNC|Rotavirus C VP7 gene|Rotavirus C VP7 gene
C4533043|T201|COMP|87711-8|LNC|Rotavirus B VP7 gene|Rotavirus B VP7 gene
C4533045|T201|COMP|87712-6|LNC|Rotavirus A VP7 gene|Rotavirus A VP7 gene
C4533047|T201|COMP|87713-4|LNC|Rotavirus A VP4 gene|Rotavirus A VP4 gene
C4533049|T201|COMP|87714-2|LNC|Influenza virus A M gene|Influenza virus A M gene
C4533050|T201|COMP|87715-9|LNC|Influenza virus A HA gene|Influenza virus A HA gene
C4533052|T201|COMP|87716-7|LNC|Influenza virus A NA gene|Influenza virus A NA gene
C4533061|T201|COMP|87722-5|LNC|Complement C1q.functional|Complement C1q.functional
C4533063|T201|COMP|87723-3|LNC|Complement C3.functional|Complement C3.functional
C4533065|T201|COMP|87724-1|LNC|Complement C7.functional|Complement C7.functional
C4533067|T201|COMP|87725-8|LNC|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C4533068|T201|COMP|87726-6|LNC|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C4533069|T201|COMP|87727-4|LNC|Complement C9.functional|Complement C9.functional
C4533071|T201|COMP|87728-2|LNC|Appearance|Appearance
C4533073|T201|COMP|87730-8|LNC|HBA1 & HBA2 gene full mutation analysis|HBA1 & HBA2 gene full mutation analysis
C4533075|T201|COMP|87731-6|LNC|KIT gene exon 17 targeted mutation analysis|KIT gene exon 17 targeted mutation analysis
C4533077|T201|COMP|87732-4|LNC|KIT gene exon 13 targeted mutation analysis|KIT gene exon 13 targeted mutation analysis
C4533079|T201|COMP|87733-2|LNC|KIT gene exon 8 targeted mutation analysis|KIT gene exon 8 targeted mutation analysis
C4533081|T201|COMP|87734-0|LNC|cefTAZidime+Avibactam|cefTAZidime+Avibactam
C4533082|T201|COMP|87735-7|LNC|Ceftolozane+Tazobactam|Ceftolozane+Tazobactam
C4533084|T201|COMP|87737-3|LNC|3,4,5-trimethylphenyl methylcarbamate|3,4,5-trimethylphenyl methylcarbamate
C4533091|T201|COMP|87742-3|LNC|Adalimumab Ab|Adalimumab Ab
C4533092|T201|COMP|87743-1|LNC|Bufencarb|Bufencarb
C4533094|T201|COMP|87744-9|LNC|Carbaryl|Carbaryl
C4533095|T201|COMP|87745-6|LNC|Carbophenothion|Carbophenothion
C4533096|T201|COMP|87746-4|LNC|Chlordane|Chlordane
C4533097|T201|COMP|87747-2|LNC|Chlorpyrifos|Chlorpyrifos
C4533098|T201|COMP|87748-0|LNC|Coumaphos|Coumaphos
C4533099|T201|COMP|87749-8|LNC|Crotoxyphos|Crotoxyphos
C4533100|T201|COMP|87750-6|LNC|Dichlorvos|Dichlorvos
C4533101|T201|COMP|87751-4|LNC|Endosulfan II|Endosulfan II
C4533103|T201|COMP|87752-2|LNC|O-Ethyl O-(p-nitrophenyl) phenylphosphonothionate|O-Ethyl O-(p-nitrophenyl) phenylphosphonothionate
C4533104|T201|COMP|87753-0|LNC|Propoxur|Propoxur
C4533105|T201|COMP|87754-8|LNC|Terbufos|Terbufos
C4533106|T201|COMP|87755-5|LNC|Clostridioides difficile BI-NAP1-027 strain DNA|Clostridioides difficile BI-NAP1-027 strain DNA
C4533110|T201|COMP|87757-1|LNC|Platelet glycoprotein IV Ab|Platelet glycoprotein IV Ab
C4533112|T201|COMP|87758-9|LNC|Naegleria fowleri DNA|Naegleria fowleri DNA
C4533115|T201|COMP|87760-5|LNC|N-Nortramadol/Creatinine|N-Nortramadol/Creatinine
C4533117|T201|COMP|87761-3|LNC|Atomoxetine/Creatinine|Atomoxetine/Creatinine
C4533119|T201|COMP|87762-1|LNC|Methcathinone/Creatinine|Methcathinone/Creatinine
C4533121|T201|COMP|87763-9|LNC|Ezogabine/Creatinine|Ezogabine/Creatinine
C4533123|T201|COMP|87764-7|LNC|Pregabalin/Creatinine|Pregabalin/Creatinine
C4533124|T201|COMP|87765-4|LNC|levETIRAcetam/Creatinine|levETIRAcetam/Creatinine
C4533126|T201|COMP|87766-2|LNC|10-Hydroxycarbazepine/Creatinine|10-Hydroxycarbazepine/Creatinine
C4533128|T201|COMP|87771-2|LNC|Zonisamide/Creatinine|Zonisamide/Creatinine
C4533130|T201|COMP|87772-0|LNC|lamoTRIgine/Creatinine|lamoTRIgine/Creatinine
C4533132|T201|COMP|87773-8|LNC|Baclofen/Creatinine|Baclofen/Creatinine
C4533134|T201|COMP|87774-6|LNC|tiZANidine/Creatinine|tiZANidine/Creatinine
C4533136|T201|COMP|87775-3|LNC|Metaxalone/Creatinine|Metaxalone/Creatinine
C4533138|T201|COMP|87776-1|LNC|Zaleplon/Creatinine|Zaleplon/Creatinine
C4533140|T201|COMP|87777-9|LNC|8-Hydroxyloxapine/Creatinine|8-Hydroxyloxapine/Creatinine
C4533142|T201|COMP|87778-7|LNC|Molindone/Creatinine|Molindone/Creatinine
C4533144|T201|COMP|87779-5|LNC|Pimozide/Creatinine|Pimozide/Creatinine
C4533146|T201|COMP|87780-3|LNC|Ziprasidone/Creatinine|Ziprasidone/Creatinine
C4533148|T201|COMP|87781-1|LNC|ARIPiprazole/Creatinine|ARIPiprazole/Creatinine
C4533150|T201|COMP|87782-9|LNC|Diclofenac/Creatinine|Diclofenac/Creatinine
C4533152|T201|COMP|87783-7|LNC|Ketoprofen/Creatinine|Ketoprofen/Creatinine
C4533154|T201|COMP|87784-5|LNC|Naproxen/Creatinine|Naproxen/Creatinine
C4533156|T201|COMP|87785-2|LNC|Oxaprozin/Creatinine|Oxaprozin/Creatinine
C4533158|T201|COMP|87786-0|LNC|Bupivacaine/Creatinine|Bupivacaine/Creatinine
C4533160|T201|COMP|87787-8|LNC|guaiFENesin/Creatinine|guaiFENesin/Creatinine
C4533162|T201|COMP|87788-6|LNC|Milnacipran/Creatinine|Milnacipran/Creatinine
C4533164|T201|COMP|87789-4|LNC|Theophylline/Creatinine|Theophylline/Creatinine
C4533166|T201|COMP|87790-2|LNC|Carbadox|Carbadox
C4533167|T201|COMP|87791-0|LNC|Carbadox|Carbadox
C4533168|T201|COMP|87792-8|LNC|Cefovecin|Cefovecin
C4533169|T201|COMP|87793-6|LNC|Nitrofurazone|Nitrofurazone
C4533170|T201|COMP|87794-4|LNC|Furazolidone|Furazolidone
C4533171|T201|COMP|87795-1|LNC|Ormetoprim+Sulfadimethoxine|Ormetoprim+Sulfadimethoxine
C4533172|T201|COMP|87796-9|LNC|Sulfathiazole|Sulfathiazole
C4533173|T201|COMP|87797-7|LNC|Sulfathiazole|Sulfathiazole
C4533174|T201|COMP|87798-5|LNC|Tulathromycin|Tulathromycin
C4533175|T201|COMP|87799-3|LNC|Sulfadimethoxine|Sulfadimethoxine
C4533176|T201|COMP|87800-9|LNC|Pradofloxacin|Pradofloxacin
C4533177|T201|COMP|87801-7|LNC|Ormetoprim+Sulfadimethoxine|Ormetoprim+Sulfadimethoxine
C4533178|T201|COMP|87802-5|LNC|Sulfachloropyridazine|Sulfachloropyridazine
C4533179|T201|COMP|87803-3|LNC|Sulfadimethoxine|Sulfadimethoxine
C4533180|T201|COMP|87804-1|LNC|Sulfachloropyridazine|Sulfachloropyridazine
C4533181|T201|COMP|87805-8|LNC|Methylphenidate|Methylphenidate
C4533182|T201|COMP|87806-6|LNC|Methylphenidate|Methylphenidate
C4533183|T201|COMP|87807-4|LNC|Naloxone|Naloxone
C4533184|T201|COMP|87808-2|LNC|chlordiazePOXIDE|chlordiazePOXIDE
C4533185|T201|COMP|87809-0|LNC|Benzoylecgonine|Benzoylecgonine
C4533186|T201|COMP|87810-8|LNC|Methylenedioxymethamphetamine|Methylenedioxymethamphetamine
C4533187|T201|COMP|87811-6|LNC|Meprobamate|Meprobamate
C4533188|T201|COMP|87812-4|LNC|Flunitrazepam|Flunitrazepam
C4533189|T201|COMP|87813-2|LNC|Flurazepam|Flurazepam
C4533190|T201|COMP|87814-0|LNC|Midazolam|Midazolam
C4533191|T201|COMP|87815-7|LNC|fentaNYL|fentaNYL
C4533192|T201|COMP|87816-5|LNC|6-Monoacetylmorphine|6-Monoacetylmorphine
C4533193|T201|COMP|87817-3|LNC|Propoxyphene|Propoxyphene
C4533194|T201|COMP|87818-1|LNC|Tapentadol|Tapentadol
C4533195|T201|COMP|87819-9|LNC|Tapentadol|Tapentadol
C4533196|T201|COMP|87820-7|LNC|Zolpidem|Zolpidem
C4533197|T201|COMP|87821-5|LNC|Zolpidem|Zolpidem
C4533198|T201|COMP|87822-3|LNC|Naltrexone|Naltrexone
C4533199|T201|COMP|87823-1|LNC|Naltrexone|Naltrexone
C4533200|T201|COMP|87824-9|LNC|6-Beta naltrexol|6-Beta naltrexol
C4533201|T201|COMP|87826-4|LNC|t(11;18)(q21;q21)(BIRC3,MALT1) fusion transcript|t(11;18)(q21;q21)(BIRC3,MALT1) fusion transcript
C4533202|T201|COMP|87827-2|LNC|Casts|Casts
C4533203|T201|COMP|87828-0|LNC|Crystals|Crystals
C4533204|T201|COMP|87829-8|LNC|Bacteria|Bacteria
C4533205|T201|COMP|87830-6|LNC|Epithelial cells|Epithelial cells
C4533206|T201|COMP|87831-4|LNC|Yeast|Yeast
C4533207|T201|COMP|87832-2|LNC|Fibroblast growth factor 21.intact|Fibroblast growth factor 21.intact
C4533209|T201|COMP|87833-0|LNC|Protein.monoclonal band 3|Protein.monoclonal band 3
C4533210|T201|COMP|87834-8|LNC|Protein.monoclonal band 2|Protein.monoclonal band 2
C4533211|T201|COMP|87835-5|LNC|Protein.monoclonal|Protein.monoclonal
C4533319|T201|COMP|87923-9|LNC|Rickettsia conorii Ab.IgM|Rickettsia conorii Ab.IgM
C4533320|T201|COMP|87924-7|LNC|Rickettsia conorii Ab.IgG|Rickettsia conorii Ab.IgG
C4533321|T201|COMP|87926-2|LNC|Epithelial cells|Epithelial cells
C4533322|T201|COMP|87927-0|LNC|Bacterial susceptibility panel|Bacterial susceptibility panel
C4533323|T201|COMP|87928-8|LNC|Macroscopic observation|Macroscopic observation
C4533324|T201|COMP|87929-6|LNC|Bacteria identified|Bacteria identified
C4533325|T201|COMP|87930-4|LNC|Bacteria identified|Bacteria identified
C4533326|T201|COMP|87931-2|LNC|Bacteria identified|Bacteria identified
C4533327|T201|COMP|87932-0|LNC|Bacteria identified|Bacteria identified
C4533328|T201|COMP|87933-8|LNC|Bacteria identified|Bacteria identified
C4533329|T201|COMP|87934-6|LNC|Bacteria identified|Bacteria identified
C4533330|T201|COMP|87935-3|LNC|Bacteria identified|Bacteria identified
C4533331|T201|COMP|87936-1|LNC|Bacteria identified|Bacteria identified
C4533332|T201|COMP|87937-9|LNC|Bacteria identified|Bacteria identified
C4533333|T201|COMP|87938-7|LNC|Bacteria identified|Bacteria identified
C4533334|T201|COMP|87939-5|LNC|Bacteria identified|Bacteria identified
C4533335|T201|COMP|87940-3|LNC|Bacteria identified|Bacteria identified
C4533336|T201|COMP|87949-4|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C4533337|T201|COMP|87950-2|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C4533338|T201|COMP|87951-0|LNC|Escherichia coli eaeA gene|Escherichia coli eaeA gene
C4533339|T201|COMP|87952-8|LNC|Helicobacter pylori|Helicobacter pylori
C4533340|T201|COMP|87953-6|LNC|Helicobacter pylori|Helicobacter pylori
C4533341|T201|COMP|87954-4|LNC|Bacteria identified|Bacteria identified
C4533342|T201|COMP|87955-1|LNC|Bacteria identified|Bacteria identified
C4533343|T201|COMP|87956-9|LNC|Legionella sp identified|Legionella sp identified
C4533344|T201|COMP|87957-7|LNC|Legionella sp identified|Legionella sp identified
C4533345|T201|COMP|87958-5|LNC|Neisseria meningitidis|Neisseria meningitidis
C4533346|T201|COMP|87959-3|LNC|Adenovirus Ag|Adenovirus Ag
C4533347|T201|COMP|87960-1|LNC|Enterovirus RNA|Enterovirus RNA
C4533348|T201|COMP|87961-9|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C4533349|T201|COMP|87962-7|LNC|HIV 1 subtype|HIV 1 subtype
C4533350|T201|COMP|87963-5|LNC|HIV 1 RNA tropism|HIV 1 RNA tropism
C4533351|T201|COMP|87964-3|LNC|Respiratory pathogens panel|Respiratory pathogens panel
C4533363|T201|COMP|87976-7|LNC|Fungus identified|Fungus identified
C4533364|T201|COMP|87977-5|LNC|Fungus identified|Fungus identified
C4533365|T201|COMP|87978-3|LNC|Fungus identified|Fungus identified
C4533366|T201|COMP|87979-1|LNC|Fungus identified|Fungus identified
C4533367|T201|COMP|87980-9|LNC|Fungus identified|Fungus identified
C4533368|T201|COMP|87981-7|LNC|Fungus identified|Fungus identified
C4533369|T201|COMP|87982-5|LNC|Toxoplasma gondii|Toxoplasma gondii
C4533370|T201|COMP|87983-3|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C4533371|T201|COMP|87984-1|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C4533372|T201|COMP|87985-8|LNC|Trichinella spiralis DNA|Trichinella spiralis DNA
C4533374|T201|COMP|87986-6|LNC|Leishmania sp identified|Leishmania sp identified
C4533375|T201|COMP|87987-4|LNC|Leishmania sp identified|Leishmania sp identified
C4533376|T201|COMP|87988-2|LNC|Acanthamoeba sp DNA|Acanthamoeba sp DNA
C4533377|T201|COMP|87989-0|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C4533378|T201|COMP|87990-8|LNC|Acanthamoeba sp identified|Acanthamoeba sp identified
C4533379|T201|COMP|87991-6|LNC|Acanthamoeba sp identified|Acanthamoeba sp identified
C4533380|T201|COMP|87992-4|LNC|Onchocerca sp Ab.IgG|Onchocerca sp Ab.IgG
C4533381|T201|COMP|87993-2|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C4533382|T201|COMP|87994-0|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C4533383|T201|COMP|87995-7|LNC|Strongyloides sp identified|Strongyloides sp identified
C4533385|T201|COMP|87996-5|LNC|Fasciola hepatica Ab|Fasciola hepatica Ab
C4533386|T201|COMP|87997-3|LNC|Trypanosoma cruzi Ab.IgM|Trypanosoma cruzi Ab.IgM
C4533387|T201|COMP|87998-1|LNC|Amoeba identified|Amoeba identified
C4533391|T201|COMP|88002-1|LNC|Kanamycin 2.5 ug/mL|Kanamycin 2.5 ug/mL
C4533396|T201|COMP|88005-4|LNC|Glutarylcarnitine (C5-DC)/Acetylcarnitine (C2)|Glutarylcarnitine (C5-DC)/Acetylcarnitine (C2)
C4533398|T201|COMP|88006-2|LNC|Octanoylcarnitine (C8)/Carnitine.free (C0)|Octanoylcarnitine (C8)/Carnitine.free (C0)
C4533401|T201|COMP|88008-8|LNC|Palmitoylcarnitine (C16)/Carnitine.free (C0)|Palmitoylcarnitine (C16)/Carnitine.free (C0)
C4533403|T201|COMP|88009-6|LNC|Palmitoylcarnitine (C16)/Acetylcarnitine (C2)|Palmitoylcarnitine (C16)/Acetylcarnitine (C2)
C4533408|T201|COMP|88012-0|LNC|Sialate.lipid bound/Creatinine|Sialate.lipid bound/Creatinine
C4533411|T201|COMP|88014-6|LNC|Octanoylcarnitine (C8)/Carnitine.free (C0)|Octanoylcarnitine (C8)/Carnitine.free (C0)
C4533412|T201|COMP|88015-3|LNC|Palmitoylcarnitine (C16)/Acetylcarnitine (C2)|Palmitoylcarnitine (C16)/Acetylcarnitine (C2)
C4533413|T201|COMP|88016-1|LNC|Glutarylcarnitine (C5-DC)/Acetylcarnitine (C2)|Glutarylcarnitine (C5-DC)/Acetylcarnitine (C2)
C4533414|T201|COMP|88017-9|LNC|Glutarylcarnitine (C5-DC)/Propionylcarnitine (C3)|Glutarylcarnitine (C5-DC)/Propionylcarnitine (C3)
C4533416|T201|COMP|88018-7|LNC|Alanine/Lysine|Alanine/Lysine
C4533418|T201|COMP|88019-5|LNC|N-acetylgalactosamine-6-sulfatase|N-acetylgalactosamine-6-sulfatase
C4533422|T201|COMP|88022-9|LNC|5-fluoro PB-22 3-carboxyindole|5-fluoro PB-22 3-carboxyindole
C4533424|T201|COMP|88023-7|LNC|XLR-11 N-(4-hydroxypentyl)|XLR-11 N-(4-hydroxypentyl)
C4533426|T201|COMP|88024-5|LNC|Palmitoylcarnitine (C16)/Carnitine.free (C0)|Palmitoylcarnitine (C16)/Carnitine.free (C0)
C4533428|T201|COMP|88026-0|LNC|Glutarylcarnitine (C5-DC)/Propionylcarnitine (C3)|Glutarylcarnitine (C5-DC)/Propionylcarnitine (C3)
C4533429|T201|COMP|88027-8|LNC|Rh group Ag|Rh group Ag
C4533431|T201|COMP|88032-8|LNC|Organophosphate panel|Organophosphate panel
C4533441|T201|COMP|88038-5|LNC|H little y Ab|H little y Ab
C4533443|T201|COMP|88039-3|LNC|little p phenotype|little p phenotype
C4533445|T201|COMP|88041-9|LNC|little p phenotype|little p phenotype
C4533446|T201|COMP|88042-7|LNC|little p phenotype|little p phenotype
C4533447|T201|COMP|88043-5|LNC|P super little k Ab|P super little k Ab
C4533449|T201|COMP|88044-3|LNC|P super little k Ab|P super little k Ab
C4533450|T201|COMP|88045-0|LNC|P super little k Ab|P super little k Ab
C4533451|T201|COMP|88046-8|LNC|P super little k Ag|P super little k Ag
C4533453|T201|COMP|88047-6|LNC|P super little k Ag|P super little k Ag
C4533454|T201|COMP|88048-4|LNC|P super little k Ag|P super little k Ag
C4533455|T201|COMP|88049-2|LNC|P2 phenotype|P2 phenotype
C4533456|T201|COMP|88050-0|LNC|P2 phenotype|P2 phenotype
C4533457|T201|COMP|88051-8|LNC|P2 phenotype|P2 phenotype
C4533458|T201|COMP|88052-6|LNC|Cells.CD4-CD8-CD45R+TCR alpha beta+/100 cells.CD3|Cells.CD4-CD8-CD45R+TCR alpha beta+/100 cells.CD3
C4533460|T201|COMP|88053-4|LNC|Cells.CD4-CD8-CD45R+TCR alpha beta+|Cells.CD4-CD8-CD45R+TCR alpha beta+
C4533462|T201|COMP|88054-2|LNC|Lipopolysaccharide binding protein|Lipopolysaccharide binding protein
C4533463|T201|COMP|88055-9|LNC|Liver fibrosis score|Liver fibrosis score
C4533464|T201|COMP|88056-7|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C4533466|T201|COMP|88059-1|LNC|Acetaminophen|Acetaminophen
C4533467|T201|COMP|88064-1|LNC|Porcine epidemic diarrhea virus S1 gene|Porcine epidemic diarrhea virus S1 gene
C4533501|T201|COMP|88106-0|LNC|Parathyrin.intact|Parathyrin.intact
C4533504|T201|COMP|88110-2|LNC|OXcarbazepine^trough|OXcarbazepine^trough
C4533505|T201|COMP|88111-0|LNC|Gentamicin^random post extended interval dosing|Gentamicin^random post extended interval dosing
C4533506|T201|COMP|88112-8|LNC|Aspartate aminotransferase|Aspartate aminotransferase
C4533507|T201|COMP|88113-6|LNC|Erythrocytes|Erythrocytes
C4533508|T201|COMP|88114-4|LNC|Leukocytes|Leukocytes
C4533509|T201|COMP|88115-1|LNC|Round cells|Round cells
C4533510|T201|COMP|88116-9|LNC|Escherichia coli gene panel|Escherichia coli gene panel
C4533523|T201|COMP|88125-0|LNC|Escherichia coli enterotoxigenic gene panel|Escherichia coli enterotoxigenic gene panel
C4533525|T201|COMP|88127-6|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C4533526|T201|COMP|88128-4|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C4533527|T201|COMP|88133-4|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C4533528|T201|COMP|88134-2|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C4533529|T201|COMP|88135-9|LNC|Varicella zoster virus|Varicella zoster virus
C4533530|T201|COMP|88136-7|LNC|Varicella zoster virus|Varicella zoster virus
C4533531|T201|COMP|88137-5|LNC|Respiratory pathogens panel|Respiratory pathogens panel
C4533532|T201|COMP|88138-3|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C4533533|T201|COMP|88139-1|LNC|Bacteria identified|Bacteria identified
C4533534|T201|COMP|88140-9|LNC|Tropheryma whippelii DNA|Tropheryma whippelii DNA
C4533535|T201|COMP|88141-7|LNC|Bacteria identified|Bacteria identified
C4533536|T201|COMP|88142-5|LNC|Bacteria identified|Bacteria identified
C4533537|T201|COMP|88143-3|LNC|Fungus identified|Fungus identified
C4533554|T201|COMP|88160-7|LNC|Microsporidia DNA|Microsporidia DNA
C4533556|T201|COMP|88161-5|LNC|Toxoplasma gondii|Toxoplasma gondii
C4533557|T201|COMP|88162-3|LNC|Acanthamoeba sp identified|Acanthamoeba sp identified
C4533558|T201|COMP|88163-1|LNC|Acanthamoeba sp DNA|Acanthamoeba sp DNA
C4533559|T201|COMP|88164-9|LNC|Toxoplasma gondii DNA|Toxoplasma gondii DNA
C4533560|T201|COMP|88165-6|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C4533561|T201|COMP|88166-4|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C4533562|T201|COMP|88167-2|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C4533563|T201|COMP|88168-0|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C4533572|T201|COMP|88177-1|LNC|Coxiella burnetii DNA|Coxiella burnetii DNA
C4533573|T201|COMP|88178-9|LNC|Coxiella burnetii DNA|Coxiella burnetii DNA
C4533574|T201|COMP|88179-7|LNC|Wuchereria bancrofti+Brugia malayi Ab.IgG4|Wuchereria bancrofti+Brugia malayi Ab.IgG4
C4533576|T201|COMP|88180-5|LNC|Wuchereria bancrofti+Brugia malayi Ab.IgG3|Wuchereria bancrofti+Brugia malayi Ab.IgG3
C4533578|T201|COMP|88181-3|LNC|Wuchereria bancrofti+Brugia malayi Ab.IgG2|Wuchereria bancrofti+Brugia malayi Ab.IgG2
C4533580|T201|COMP|88182-1|LNC|Wuchereria bancrofti+Brugia malayi Ab.IgG1|Wuchereria bancrofti+Brugia malayi Ab.IgG1
C4533582|T201|COMP|88183-9|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C4533583|T201|COMP|88184-7|LNC|IgG+IgM.porcine|IgG+IgM.porcine
C4533585|T201|COMP|88185-4|LNC|IgG+IgM.porcine|IgG+IgM.porcine
C4533586|T201|COMP|88186-2|LNC|Ebola & Marburg virus RNA panel|Ebola & Marburg virus RNA panel
C4533588|T201|COMP|88187-0|LNC|Influenza virus A subtype|Influenza virus A subtype
C4533589|T201|COMP|88188-8|LNC|Dengue virus 1+2+3+4 RNA|Dengue virus 1+2+3+4 RNA
C4533590|T201|COMP|88189-6|LNC|Dengue virus 1+2+3+4 RNA|Dengue virus 1+2+3+4 RNA
C4533591|T201|COMP|88190-4|LNC|Crimean-Congo hemorrhagic fever virus Ab.IgM|Crimean-Congo hemorrhagic fever virus Ab.IgM
C4533593|T201|COMP|88191-2|LNC|Crimean-Congo hemorrhagic fever virus Ab.IgG|Crimean-Congo hemorrhagic fever virus Ab.IgG
C4533595|T201|COMP|88192-0|LNC|Crimean-Congo hemorrhagic fever virus RNA|Crimean-Congo hemorrhagic fever virus RNA
C4533597|T201|COMP|88193-8|LNC|Influenza virus A RNA|Influenza virus A RNA
C4533598|T201|COMP|88194-6|LNC|Influenza virus B Ag|Influenza virus B Ag
C4533599|T201|COMP|88199-5|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C4533600|T201|COMP|88200-1|LNC|Influenza virus identified|Influenza virus identified
C4533601|T201|COMP|88201-9|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C4533602|T201|COMP|88202-7|LNC|Respiratory syncytial virus B RNA|Respiratory syncytial virus B RNA
C4533603|T201|COMP|88203-5|LNC|Dengue virus 1 & 2 & 3 & 4 RNA|Dengue virus 1 & 2 & 3 & 4 RNA
C4533604|T201|COMP|88204-3|LNC|Respiratory syncytial virus A RNA|Respiratory syncytial virus A RNA
C4533605|T201|COMP|88205-0|LNC|Lymphocytic choriomeningitis virus Ab.IgM|Lymphocytic choriomeningitis virus Ab.IgM
C4533606|T201|COMP|88206-8|LNC|Lymphocytic choriomeningitis virus Ab.IgG|Lymphocytic choriomeningitis virus Ab.IgG
C4533607|T201|COMP|88207-6|LNC|Lymphocytic choriomeningitis virus RNA|Lymphocytic choriomeningitis virus RNA
C4533608|T201|COMP|88208-4|LNC|Parainfluenza virus 1 RNA|Parainfluenza virus 1 RNA
C4533609|T201|COMP|88209-2|LNC|Parainfluenza virus 2 RNA|Parainfluenza virus 2 RNA
C4533610|T201|COMP|88210-0|LNC|Parainfluenza virus 3 RNA|Parainfluenza virus 3 RNA
C4533611|T201|COMP|88211-8|LNC|Rabies virus Ag|Rabies virus Ag
C4533612|T201|COMP|88212-6|LNC|HIV 1 proviral DNA|HIV 1 proviral DNA
C4533613|T201|COMP|88213-4|LNC|Rhinovirus RNA|Rhinovirus RNA
C4533614|T201|COMP|88214-2|LNC|Rabies virus RNA|Rabies virus RNA
C4533615|T201|COMP|88215-9|LNC|Rabies virus RNA|Rabies virus RNA
C4533616|T201|COMP|88216-7|LNC|Hantavirus puumala RNA|Hantavirus puumala RNA
C4533618|T201|COMP|88217-5|LNC|Parechovirus RNA|Parechovirus RNA
C4533619|T201|COMP|88218-3|LNC|Parechovirus RNA|Parechovirus RNA
C4533620|T201|COMP|88219-1|LNC|Parechovirus RNA|Parechovirus RNA
C4533621|T201|COMP|88220-9|LNC|Hantavirus puumala RNA|Hantavirus puumala RNA
C4533622|T201|COMP|88221-7|LNC|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C4533623|T201|COMP|88222-5|LNC|Human metapneumovirus Ag|Human metapneumovirus Ag
C4533624|T201|COMP|88223-3|LNC|Francisella sp DNA|Francisella sp DNA
C4533626|T201|COMP|88224-1|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C4533627|T201|COMP|88225-8|LNC|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C4533628|T201|COMP|88226-6|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C4533629|T201|COMP|88227-4|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C4533630|T201|COMP|88228-2|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C4533631|T201|COMP|88229-0|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C4533632|T201|COMP|88230-8|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C4533634|T201|COMP|88232-4|LNC|Trypanosoma cruzi DNA|Trypanosoma cruzi DNA
C4533635|T201|COMP|88233-2|LNC|Babesia sp DNA|Babesia sp DNA
C4533638|T201|COMP|88236-5|LNC|Bacteria identified|Bacteria identified
C4533646|T201|COMP|88244-9|LNC|Acinetobacter sp (rpsA) gene|Acinetobacter sp (rpsA) gene
C4533647|T201|COMP|88245-6|LNC|Bacterial carbapenem resistance blaIMP gene|Bacterial carbapenem resistance blaIMP gene
C4533648|T201|COMP|88246-4|LNC|Bacterial carbapenem resistance blaKPC gene|Bacterial carbapenem resistance blaKPC gene
C4533649|T201|COMP|88247-2|LNC|Bacterial carbapenem resistance blaNDM gene|Bacterial carbapenem resistance blaNDM gene
C4533650|T201|COMP|88248-0|LNC|Bacterial carbapenem resistance blaOXA gene|Bacterial carbapenem resistance blaOXA gene
C4533651|T201|COMP|88249-8|LNC|Bacterial carbapenem resistance blaVIM gene|Bacterial carbapenem resistance blaVIM gene
C4533652|T201|COMP|88250-6|LNC|Bacterial cephalosporin resistance blaCTX-M gene|Bacterial cephalosporin resistance blaCTX-M gene
C4533653|T201|COMP|88251-4|LNC|Bacterial methicillin resistance mecA gene|Bacterial methicillin resistance mecA gene
C4533654|T201|COMP|88252-2|LNC|Bacterial vancomycin resistance vanA gene|Bacterial vancomycin resistance vanA gene
C4533655|T201|COMP|88253-0|LNC|Bacterial vancomycin resistance vanB gene|Bacterial vancomycin resistance vanB gene
C4533656|T201|COMP|88254-8|LNC|Citrobacter sp (ompA+mrkC) genes|Citrobacter sp (ompA+mrkC) genes
C4533657|T201|COMP|88255-5|LNC|Enterobacter sp (gyrB+metB) genes|Enterobacter sp (gyrB+metB) genes
C4533658|T201|COMP|88256-3|LNC|Enterococcus faecalis hsp60 gene|Enterococcus faecalis hsp60 gene
C4533659|T201|COMP|88257-1|LNC|Enterococcus faecium hsp60 gene|Enterococcus faecium hsp60 gene
C4533660|T201|COMP|88261-3|LNC|Gram positive bacteria identified|Gram positive bacteria identified
C4533661|T201|COMP|88262-1|LNC|Gram positive blood culture panel|Gram positive blood culture panel
C4533662|T201|COMP|88263-9|LNC|Klebsiella oxytoca (ompA) gene|Klebsiella oxytoca (ompA) gene
C4533663|T201|COMP|88264-7|LNC|Klebsiella pneumoniae yggE gene|Klebsiella pneumoniae yggE gene
C4533664|T201|COMP|88265-4|LNC|Listeria sp (tuf) gene|Listeria sp (tuf) gene
C4533665|T201|COMP|88266-2|LNC|Mycobacterium sp rRNA|Mycobacterium sp rRNA
C4533666|T201|COMP|88267-0|LNC|Proteus sp (atpD) gene|Proteus sp (atpD) gene
C4533667|T201|COMP|88268-8|LNC|Pseudomonas aeruginosa (sodA) gene|Pseudomonas aeruginosa (sodA) gene
C4533668|T201|COMP|88269-6|LNC|Staphylococcus aureus gyrB gene|Staphylococcus aureus gyrB gene
C4533669|T201|COMP|88270-4|LNC|Staphylococcus epidermidis hsp60 gene|Staphylococcus epidermidis hsp60 gene
C4533670|T201|COMP|88271-2|LNC|Staphylococcus lugdunensis sodA gene|Staphylococcus lugdunensis sodA gene
C4533671|T201|COMP|88272-0|LNC|Staphylococcus sp tuf gene|Staphylococcus sp tuf gene
C4533672|T201|COMP|88273-8|LNC|Streptococcus agalactiae hsp60 gene|Streptococcus agalactiae hsp60 gene
C4533673|T201|COMP|88274-6|LNC|Streptococcus anginosus group gyrB gene|Streptococcus anginosus group gyrB gene
C4533674|T201|COMP|88275-3|LNC|Streptococcus pneumoniae gryB gene|Streptococcus pneumoniae gryB gene
C4533675|T201|COMP|88276-1|LNC|Streptococcus pyogenes hsp60 gene|Streptococcus pyogenes hsp60 gene
C4533676|T201|COMP|88277-9|LNC|Streptococcus sp tuf gene|Streptococcus sp tuf gene
C4554784|T201|COMP|89543-3|LNC|Laboratory ask at order entry panel|Laboratory ask at order entry panel
C4695133|T201|COMP|83128-9|LNC|Hepatitis E virus Ab.IgM|Hepatitis E virus Ab.IgM
C4695170|T201|COMP|87333-1|LNC|Porcine circovirus type 2 ORF2 gene|Porcine circovirus type 2 ORF2 gene
C4695172|T201|COMP|87349-7|LNC|Senecavirus A VP1 gene|Senecavirus A VP1 gene
C4695174|T201|COMP|87638-3|LNC|p,p'- Dichlorodiphenyldichloroethane|p,p'- Dichlorodiphenyldichloroethane
C4695176|T201|COMP|87639-1|LNC|Dichlorodiphenyltrichloroethane|Dichlorodiphenyltrichloroethane
C4695177|T201|COMP|87640-9|LNC|Dichlorodiphenyldichloroethylene|Dichlorodiphenyldichloroethylene
C4695178|T201|COMP|87641-7|LNC|o,p'- Dichlorodiphenyltrichloroethane|o,p'- Dichlorodiphenyltrichloroethane
C4695179|T201|COMP|87642-5|LNC|o,p'- Dichlorodiphenyldichloroethylene|o,p'- Dichlorodiphenyldichloroethylene
C4695181|T201|COMP|87643-3|LNC|o,p'- Dichlorodiphenyldichloroethane|o,p'- Dichlorodiphenyldichloroethane
C4695183|T201|COMP|88304-1|LNC|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C4695199|T201|COMP|88446-0|LNC|Hydrogen/Expired gas^20M post dose lactose PO|Hydrogen/Expired gas^20M post dose lactose PO
C4695209|T201|COMP|88603-6|LNC|Adenovirus Ag|Adenovirus Ag
C4695210|T201|COMP|88604-4|LNC|Human coronavirus HKU1 RNA|Human coronavirus HKU1 RNA
C4695211|T201|COMP|88605-1|LNC|Human coronavirus OC43 RNA|Human coronavirus OC43 RNA
C4695212|T201|COMP|88606-9|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C4695213|T201|COMP|88607-7|LNC|Human coronavirus 229E RNA|Human coronavirus 229E RNA
C4695214|T201|COMP|88608-5|LNC|Human coronavirus 229E RNA|Human coronavirus 229E RNA
C4695228|T201|COMP|88447-8|LNC|Liver fibrosis interpretation|Liver fibrosis interpretation
C4695230|T201|COMP|88448-6|LNC|Necroinflammatory activity interpretation|Necroinflammatory activity interpretation
C4695232|T201|COMP|88449-4|LNC|Coagulation factor IX activity actual/Normal|Coagulation factor IX activity actual/Normal
C4695233|T201|COMP|88724-0|LNC|Ganglioside GD1a Ab.IgG+IgM|Ganglioside GD1a Ab.IgG+IgM
C4695234|T201|COMP|88725-7|LNC|MDA5 Ab|MDA5 Ab
C4695235|T201|COMP|88726-5|LNC|Glial nuclear type 1 Ab|Glial nuclear type 1 Ab
C4695236|T201|COMP|88727-3|LNC|Recoverin Ab|Recoverin Ab
C4695237|T201|COMP|88728-1|LNC|Babesia microti Ab.IgG & IgM panel|Babesia microti Ab.IgG & IgM panel
C4695254|T201|COMP|88580-6|LNC|Burkholderia sp identified|Burkholderia sp identified
C4695255|T201|COMP|88581-4|LNC|Borrelia sp DNA|Borrelia sp DNA
C4695256|T201|COMP|88582-2|LNC|Bordetella sp identified|Bordetella sp identified
C4695257|T201|COMP|88583-0|LNC|Bordetella sp DNA|Bordetella sp DNA
C4695262|T201|COMP|88713-3|LNC|Phosphate|Phosphate
C4695263|T201|COMP|88714-1|LNC|Dehydroaripiprazole|Dehydroaripiprazole
C4695264|T201|COMP|88715-8|LNC|Norquetiapine|Norquetiapine
C4695265|T201|COMP|88716-6|LNC|Adenovirus A+B+C+D+E+F DNA|Adenovirus A+B+C+D+E+F DNA
C4695267|T201|COMP|88838-8|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4695269|T201|COMP|88839-6|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4695270|T201|COMP|88840-4|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4695271|T201|COMP|88841-2|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4695272|T201|COMP|88842-0|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4695273|T201|COMP|88883-4|LNC|Autoimmune connective tissue Ab panel|Autoimmune connective tissue Ab panel
C4695275|T201|COMP|88884-2|LNC|Fatty acid omega-3 & omega-6 panel|Fatty acid omega-3 & omega-6 panel
C4695277|T201|COMP|88885-9|LNC|Delafloxacin|Delafloxacin
C4695278|T201|COMP|88886-7|LNC|Telavancin|Telavancin
C4695279|T201|COMP|88887-5|LNC|Isavuconazole|Isavuconazole
C4695332|T201|COMP|88301-7|LNC|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C4695333|T201|COMP|88302-5|LNC|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C4695334|T201|COMP|88303-3|LNC|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C4695369|T201|COMP|88335-5|LNC|Predominant leukocyte identified|Predominant leukocyte identified
C4695372|T201|COMP|88337-1|LNC|Mite identified|Mite identified
C4695373|T201|COMP|88338-9|LNC|Coccal bacteria|Coccal bacteria
C4695375|T201|COMP|88339-7|LNC|Bacilliform bacteria|Bacilliform bacteria
C4695377|T201|COMP|88340-5|LNC|Mite|Mite
C4695378|T201|COMP|88341-3|LNC|Cerumen|Cerumen
C4695379|T201|COMP|88342-1|LNC|Malassezia sp|Malassezia sp
C4695380|T201|COMP|88343-9|LNC|Leukocytes|Leukocytes
C4695381|T201|COMP|88344-7|LNC|Intracellular bacteria|Intracellular bacteria
C4695383|T201|COMP|88345-4|LNC|Microscopic exam panel|Microscopic exam panel
C4695404|T201|COMP|88365-2|LNC|Glucose^pre-meal|Glucose^pre-meal
C4695422|T201|COMP|88375-1|LNC|Tildipirosin|Tildipirosin
C4695423|T201|COMP|88376-9|LNC|Gamithromycin|Gamithromycin
C4695424|T201|COMP|88377-7|LNC|Tildipirosin|Tildipirosin
C4695425|T201|COMP|88378-5|LNC|Gamithromycin|Gamithromycin
C4695524|T201|COMP|88439-5|LNC|Hydrogen/Expired gas^10M post dose fructose PO|Hydrogen/Expired gas^10M post dose fructose PO
C4695525|T201|COMP|88440-3|LNC|Hydrogen/Expired gas^10M post dose lactose PO|Hydrogen/Expired gas^10M post dose lactose PO
C4695526|T201|COMP|88441-1|LNC|Hydrogen/Expired gas^20M post dose fructose PO|Hydrogen/Expired gas^20M post dose fructose PO
C4695527|T201|COMP|88442-9|LNC|Hydrogen/Expired gas^40M post dose lactose PO|Hydrogen/Expired gas^40M post dose lactose PO
C4695528|T201|COMP|88443-7|LNC|Hydrogen/Expired gas^40M post dose fructose PO|Hydrogen/Expired gas^40M post dose fructose PO
C4695529|T201|COMP|88444-5|LNC|Hydrogen/Expired gas^50M post dose fructose PO|Hydrogen/Expired gas^50M post dose fructose PO
C4695530|T201|COMP|88445-2|LNC|Hydrogen/Expired gas^50M post dose lactose PO|Hydrogen/Expired gas^50M post dose lactose PO
C4695531|T201|COMP|88450-2|LNC|Babesia divergens+MO-1 strain 18S rRNA gene|Babesia divergens+MO-1 strain 18S rRNA gene
C4695533|T201|COMP|88451-0|LNC|Babesia duncani 18S rRNA gene|Babesia duncani 18S rRNA gene
C4695535|T201|COMP|88452-8|LNC|Babesia microti 18S rRNA gene|Babesia microti 18S rRNA gene
C4695538|T201|COMP|88454-4|LNC|Mumps virus Ab.IgG+IgM|Mumps virus Ab.IgG+IgM
C4695539|T201|COMP|88455-1|LNC|California encephalitis virus Ab.IgG & IgM panel|California encephalitis virus Ab.IgG & IgM panel
C4695541|T201|COMP|88456-9|LNC|California encephalitis virus Ab.IgG+IgM|California encephalitis virus Ab.IgG+IgM
C4695543|T201|COMP|88457-7|LNC|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C4695544|T201|COMP|88458-5|LNC|Mumps virus Ab.IgG & IgM panel|Mumps virus Ab.IgG & IgM panel
C4695552|T201|COMP|88462-7|LNC|Carbapenem|Carbapenem
C4695647|T201|COMP|88516-0|LNC|Gastrointestinal pathogens identified|Gastrointestinal pathogens identified
C4695651|T201|COMP|88519-4|LNC|KIT gene.c.2447A>T|KIT gene.c.2447A>T
C4695666|T201|COMP|88527-7|LNC|Respiratory syncytial virus identified|Respiratory syncytial virus identified
C4695667|T201|COMP|88528-5|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C4695668|T201|COMP|88529-3|LNC|Parainfluenza virus RNA|Parainfluenza virus RNA
C4695669|T201|COMP|88530-1|LNC|Parainfluenza virus 4 RNA|Parainfluenza virus 4 RNA
C4695670|T201|COMP|88531-9|LNC|Parainfluenza virus identified|Parainfluenza virus identified
C4695671|T201|COMP|88532-7|LNC|Human metapneumovirus Identified|Human metapneumovirus Identified
C4695673|T201|COMP|88533-5|LNC|Adenovirus DNA|Adenovirus DNA
C4695674|T201|COMP|88534-3|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C4695675|T201|COMP|88535-0|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C4695676|T201|COMP|88536-8|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C4695677|T201|COMP|88537-6|LNC|Enterovirus identified|Enterovirus identified
C4695678|T201|COMP|88538-4|LNC|Enterovirus RNA|Enterovirus RNA
C4695679|T201|COMP|88539-2|LNC|Adenovirus DNA|Adenovirus DNA
C4695680|T201|COMP|88540-0|LNC|Enterovirus RNA|Enterovirus RNA
C4695681|T201|COMP|88541-8|LNC|Adenovirus DNA|Adenovirus DNA
C4695682|T201|COMP|88542-6|LNC|HIV 1 RNA integrase gene mutations detected|HIV 1 RNA integrase gene mutations detected
C4695684|T201|COMP|88543-4|LNC|HIV 1 RNA protease gene mutations detected|HIV 1 RNA protease gene mutations detected
C4695688|T201|COMP|88545-9|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C4695689|T201|COMP|88546-7|LNC|Chlamydophila pneumoniae DNA|Chlamydophila pneumoniae DNA
C4695690|T201|COMP|88547-5|LNC|Chlamydophila pneumoniae DNA|Chlamydophila pneumoniae DNA
C4695691|T201|COMP|88548-3|LNC|Scedosporium apiospermum DNA|Scedosporium apiospermum DNA
C4695693|T201|COMP|88549-1|LNC|Scedosporium apiospermum DNA|Scedosporium apiospermum DNA
C4695694|T201|COMP|88550-9|LNC|Scedosporium apiospermum DNA|Scedosporium apiospermum DNA
C4695695|T201|COMP|88551-7|LNC|Scedosporium apiospermum DNA|Scedosporium apiospermum DNA
C4695696|T201|COMP|88552-5|LNC|Scedosporium prolificans DNA|Scedosporium prolificans DNA
C4695698|T201|COMP|88553-3|LNC|Scedosporium prolificans DNA|Scedosporium prolificans DNA
C4695699|T201|COMP|88554-1|LNC|Scedosporium prolificans DNA|Scedosporium prolificans DNA
C4695700|T201|COMP|88555-8|LNC|Galactomannan Ag|Galactomannan Ag
C4695701|T201|COMP|88556-6|LNC|Scedosporium prolificans DNA|Scedosporium prolificans DNA
C4695702|T201|COMP|88557-4|LNC|Scedosporium apiospermum DNA|Scedosporium apiospermum DNA
C4695703|T201|COMP|88558-2|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C4695704|T201|COMP|88559-0|LNC|Parainfluenza virus 2 RNA|Parainfluenza virus 2 RNA
C4695705|T201|COMP|88560-8|LNC|Parainfluenza virus 3 RNA|Parainfluenza virus 3 RNA
C4695706|T201|COMP|88561-6|LNC|Parainfluenza virus 4 RNA|Parainfluenza virus 4 RNA
C4695707|T201|COMP|88562-4|LNC|Parainfluenza virus RNA|Parainfluenza virus RNA
C4695708|T201|COMP|88563-2|LNC|Parainfluenza virus 1 RNA|Parainfluenza virus 1 RNA
C4695709|T201|COMP|88564-0|LNC|Cytomegalovirus|Cytomegalovirus
C4695710|T201|COMP|88565-7|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C4695711|T201|COMP|88566-5|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C4695712|T201|COMP|88567-3|LNC|Cytomegalovirus DNA|Cytomegalovirus DNA
C4695713|T201|COMP|88568-1|LNC|Influenza virus identified|Influenza virus identified
C4695714|T201|COMP|88569-9|LNC|Ocular pathogens panel|Ocular pathogens panel
C4695716|T201|COMP|88570-7|LNC|Acanthamoeba sp DNA|Acanthamoeba sp DNA
C4695717|T201|COMP|88571-5|LNC|Fetal monosomy X risk|Fetal monosomy X risk
C4695718|T201|COMP|88572-3|LNC|Fetal 22q11.2 deletion risk|Fetal 22q11.2 deletion risk
C4695719|T201|COMP|88573-1|LNC|Onchocerca sp Ab.IgG2|Onchocerca sp Ab.IgG2
C4695720|T201|COMP|88574-9|LNC|Onchocerca sp Ab.IgG3|Onchocerca sp Ab.IgG3
C4695721|T201|COMP|88575-6|LNC|Onchocerca sp Ab.IgG4|Onchocerca sp Ab.IgG4
C4695722|T201|COMP|88576-4|LNC|Bordetella holmesii hIS1001 DNA|Bordetella holmesii hIS1001 DNA
C4695723|T201|COMP|88577-2|LNC|Legionella pneumophila DNA|Legionella pneumophila DNA
C4695724|T201|COMP|88578-0|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C4695725|T201|COMP|88579-8|LNC|Mycoplasma pneumoniae DNA|Mycoplasma pneumoniae DNA
C4695726|T201|COMP|88584-8|LNC|Corynebacterium diphtheriae|Corynebacterium diphtheriae
C4695727|T201|COMP|88585-5|LNC|Legionella sp identified|Legionella sp identified
C4695728|T201|COMP|88586-3|LNC|Shigella sp identified|Shigella sp identified
C4695729|T201|COMP|88587-1|LNC|Legionella sp DNA|Legionella sp DNA
C4695730|T201|COMP|88588-9|LNC|Legionella sp DNA|Legionella sp DNA
C4695731|T201|COMP|88589-7|LNC|Clostridium botulinum toxin|Clostridium botulinum toxin
C4695732|T201|COMP|88590-5|LNC|Legionella pneumophila DNA|Legionella pneumophila DNA
C4695733|T201|COMP|88591-3|LNC|Scedosporium prolificans DNA|Scedosporium prolificans DNA
C4695734|T201|COMP|88592-1|LNC|Influenza virus B RNA|Influenza virus B RNA
C4695735|T201|COMP|88593-9|LNC|Human bocavirus DNA|Human bocavirus DNA
C4695736|T201|COMP|88594-7|LNC|Human coronavirus HKU1 RNA|Human coronavirus HKU1 RNA
C4695737|T201|COMP|88595-4|LNC|Respiratory syncytial virus A RNA|Respiratory syncytial virus A RNA
C4695738|T201|COMP|88596-2|LNC|Influenza virus B RNA|Influenza virus B RNA
C4695739|T201|COMP|88597-0|LNC|Respiratory syncytial virus B RNA|Respiratory syncytial virus B RNA
C4695740|T201|COMP|88598-8|LNC|Toscana virus RNA|Toscana virus RNA
C4695741|T201|COMP|88599-6|LNC|Influenza virus A RNA|Influenza virus A RNA
C4695742|T201|COMP|88600-2|LNC|Influenza virus A RNA|Influenza virus A RNA
C4695743|T201|COMP|88601-0|LNC|Influenza virus A & B RNA panel|Influenza virus A & B RNA panel
C4695745|T201|COMP|88602-8|LNC|Adenovirus Ag|Adenovirus Ag
C4695746|T201|COMP|88609-3|LNC|Human coronavirus 229E RNA|Human coronavirus 229E RNA
C4695747|T201|COMP|88610-1|LNC|Human coronavirus 229E RNA|Human coronavirus 229E RNA
C4695748|T201|COMP|88611-9|LNC|Human coronavirus HKU1 RNA|Human coronavirus HKU1 RNA
C4695749|T201|COMP|88612-7|LNC|Human coronavirus HKU1 RNA|Human coronavirus HKU1 RNA
C4695750|T201|COMP|88613-5|LNC|Human bocavirus DNA|Human bocavirus DNA
C4695751|T201|COMP|88614-3|LNC|Human coronavirus RNA|Human coronavirus RNA
C4695752|T201|COMP|88615-0|LNC|Human coronavirus NL63 RNA|Human coronavirus NL63 RNA
C4695753|T201|COMP|88616-8|LNC|Human coronavirus NL63 RNA|Human coronavirus NL63 RNA
C4695754|T201|COMP|88617-6|LNC|Human coronavirus NL63 RNA|Human coronavirus NL63 RNA
C4695755|T201|COMP|88618-4|LNC|Human coronavirus NL63 RNA|Human coronavirus NL63 RNA
C4695756|T201|COMP|88619-2|LNC|Human coronavirus OC43 RNA|Human coronavirus OC43 RNA
C4695757|T201|COMP|88620-0|LNC|Human coronavirus RNA|Human coronavirus RNA
C4695758|T201|COMP|88621-8|LNC|Human coronavirus OC43 RNA|Human coronavirus OC43 RNA
C4695759|T201|COMP|88622-6|LNC|Cytomegalovirus|Cytomegalovirus
C4695760|T201|COMP|88623-4|LNC|Cytomegalovirus|Cytomegalovirus
C4695761|T201|COMP|88624-2|LNC|Cytomegalovirus|Cytomegalovirus
C4695762|T201|COMP|88625-9|LNC|Cytomegalovirus|Cytomegalovirus
C4695763|T201|COMP|88626-7|LNC|Human coronavirus OC43 RNA|Human coronavirus OC43 RNA
C4695764|T201|COMP|88627-5|LNC|Human coronavirus RNA|Human coronavirus RNA
C4695765|T201|COMP|88628-3|LNC|Human coronavirus RNA|Human coronavirus RNA
C4695766|T201|COMP|88629-1|LNC|Chikungunya virus Ab.IgM|Chikungunya virus Ab.IgM
C4695767|T201|COMP|88630-9|LNC|Chikungunya virus Ab.IgG|Chikungunya virus Ab.IgG
C4695794|T201|COMP|88678-8|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C4695795|T201|COMP|88679-6|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C4695796|T201|COMP|88680-4|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C4695797|T201|COMP|88681-2|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C4695798|T201|COMP|88682-0|LNC|Leishmania sp Ab.IgM|Leishmania sp Ab.IgM
C4695799|T201|COMP|88683-8|LNC|Bacteria identified|Bacteria identified
C4695802|T201|COMP|88686-1|LNC|Fungus identified|Fungus identified
C4695803|T201|COMP|88687-9|LNC|Fungus identified|Fungus identified
C4695804|T201|COMP|88688-7|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C4695805|T201|COMP|88689-5|LNC|Pneumocystis jiroveci|Pneumocystis jiroveci
C4695806|T201|COMP|88690-3|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C4695807|T201|COMP|88691-1|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C4695815|T201|COMP|88697-8|LNC|Electrolytes & Osmolality panel|Electrolytes & Osmolality panel
C4695817|T201|COMP|88698-6|LNC|Protein fractions panel|Protein fractions panel
C4695818|T201|COMP|88699-4|LNC|Procainamide & N-acetylprocainamide panel|Procainamide & N-acetylprocainamide panel
C4695820|T201|COMP|88700-0|LNC|Babesia microti Ab.IgG & IgM|Babesia microti Ab.IgG & IgM
C4695821|T201|COMP|88701-8|LNC|Norovirus genogroups I & II RNA panel|Norovirus genogroups I & II RNA panel
C4695823|T201|COMP|88702-6|LNC|Systemic sclerosis panel|Systemic sclerosis panel
C4695825|T201|COMP|88703-4|LNC|Bedaquiline|Bedaquiline
C4695826|T201|COMP|88704-2|LNC|Bedaquiline|Bedaquiline
C4695827|T201|COMP|88705-9|LNC|Kanamycin 3.5 ug/mL|Kanamycin 3.5 ug/mL
C4695828|T201|COMP|88706-7|LNC|Linezolid 1.0 ug/mL|Linezolid 1.0 ug/mL
C4695830|T201|COMP|88707-5|LNC|Moxifloxacin 0.25 ug/mL|Moxifloxacin 0.25 ug/mL
C4695834|T201|COMP|88709-1|LNC|Albumin/Globulin|Albumin/Globulin
C4695835|T201|COMP|88710-9|LNC|Amylase.pancreatic|Amylase.pancreatic
C4695836|T201|COMP|88711-7|LNC|Beta-2-Microglobulin|Beta-2-Microglobulin
C4695837|T201|COMP|88712-5|LNC|Triacylglycerol lipase|Triacylglycerol lipase
C4695838|T201|COMP|88717-4|LNC|Candida sp identified|Candida sp identified
C4695839|T201|COMP|88718-2|LNC|Chlamydophila pneumoniae DNA|Chlamydophila pneumoniae DNA
C4695840|T201|COMP|88719-0|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA|Human coronavirus 229E+HKU1+NL63+OC43 RNA
C4695842|T201|COMP|88720-8|LNC|Mycoplasma pneumoniae DNA|Mycoplasma pneumoniae DNA
C4695843|T201|COMP|88721-6|LNC|Rhinovirus+enterovirus RNA|Rhinovirus+enterovirus RNA
C4695844|T201|COMP|88722-4|LNC|Streptococcus pneumoniae serotype|Streptococcus pneumoniae serotype
C4695845|T201|COMP|88723-2|LNC|Asialoganglioside GM1 Ab.IgG+IgM|Asialoganglioside GM1 Ab.IgG+IgM
C4695847|T201|COMP|88729-9|LNC|Ganglioside GQ1b Ab.IgG+IgM|Ganglioside GQ1b Ab.IgG+IgM
C4695848|T201|COMP|88730-7|LNC|Ganglioside GD1b Ab.IgG+IgM|Ganglioside GD1b Ab.IgG+IgM
C4695849|T201|COMP|88731-5|LNC|Ganglioside GM2 Ab.IgG+IgM|Ganglioside GM2 Ab.IgG+IgM
C4695850|T201|COMP|88732-3|LNC|Mi-2 alpha Ab|Mi-2 alpha Ab
C4695851|T201|COMP|88733-1|LNC|Mi-2 beta Ab|Mi-2 beta Ab
C4695852|T201|COMP|88734-9|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C4695853|T201|COMP|88735-6|LNC|PM-SCL-100 Ab|PM-SCL-100 Ab
C4695854|T201|COMP|88736-4|LNC|PM-SCL-75 Ab|PM-SCL-75 Ab
C4695855|T201|COMP|88737-2|LNC|RNA polymerase III RP11 Ab|RNA polymerase III RP11 Ab
C4695856|T201|COMP|88738-0|LNC|RNA polymerase III RP155 Ab|RNA polymerase III RP155 Ab
C4695857|T201|COMP|88739-8|LNC|TIF1-gamma Ab|TIF1-gamma Ab
C4695858|T201|COMP|88740-6|LNC|Titin Ab|Titin Ab
C4695859|T201|COMP|88741-4|LNC|U1 small nuclear ribonucleoprotein A Ab|U1 small nuclear ribonucleoprotein A Ab
C4695860|T201|COMP|88742-2|LNC|U1 small nuclear ribonucleoprotein C Ab|U1 small nuclear ribonucleoprotein C Ab
C4695861|T201|COMP|88743-0|LNC|Zinc finger protein of the cerebellum 4 Ab|Zinc finger protein of the cerebellum 4 Ab
C4695862|T201|COMP|88744-8|LNC|inv(2)(p21;p23)(EML4,ALK) fusion transcript|inv(2)(p21;p23)(EML4,ALK) fusion transcript
C4695863|T201|COMP|88745-5|LNC|Coccidioides immitis Ab.IgG & IgM panel|Coccidioides immitis Ab.IgG & IgM panel
C4695864|T201|COMP|88746-3|LNC|Toxoplasma gondii Ab.IgG & IgM panel|Toxoplasma gondii Ab.IgG & IgM panel
C4695997|T201|COMP|89327-1|LNC|Cells.CD3+CD8+CD27-CD45RO+CD62L-|Cells.CD3+CD8+CD27-CD45RO+CD62L-
C4695999|T201|COMP|89328-9|LNC|Cells.CD3+CD4+CD27-CD45RO+CD62L-|Cells.CD3+CD4+CD27-CD45RO+CD62L-
C4696001|T201|COMP|89329-7|LNC|Cells.CD3+CD4+CD27+CD45RO+CD62L+|Cells.CD3+CD4+CD27+CD45RO+CD62L+
C4696003|T201|COMP|89330-5|LNC|Cells.CD3+CD8+CD27+CD62L+|Cells.CD3+CD8+CD27+CD62L+
C4696005|T201|COMP|89331-3|LNC|Cells.CD3+CD4+CD27+CD62L+|Cells.CD3+CD4+CD27+CD62L+
C4696019|T201|COMP|89481-6|LNC|Gentamicin|Gentamicin
C4696021|T201|COMP|89482-4|LNC|Kanamycin|Kanamycin
C4696022|T201|COMP|89483-2|LNC|Capreomycin|Capreomycin
C4696023|T201|COMP|89484-0|LNC|Amikacin|Amikacin
C4696027|T201|COMP|89583-9|LNC|Cytomegalovirus Ag|Cytomegalovirus Ag
C4696028|T201|COMP|89584-7|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C4696046|T201|COMP|88892-5|LNC|Meropenem+Vaborbactam|Meropenem+Vaborbactam
C4696047|T201|COMP|88893-3|LNC|Coagulation tissue factor induced.PIVKA sensitive|Coagulation tissue factor induced.PIVKA sensitive
C4696048|T201|COMP|88894-1|LNC|Brivaracetam|Brivaracetam
C4696049|T201|COMP|88895-8|LNC|Perampanel|Perampanel
C4696050|T201|COMP|88896-6|LNC|Reboxetine|Reboxetine
C4696051|T201|COMP|88897-4|LNC|Adenovirus Ag|Adenovirus Ag
C4696052|T201|COMP|88898-2|LNC|Adenovirus|Adenovirus
C4696079|T201|COMP|89431-1|LNC|Cells.CD25/100 Cells.CD4|Cells.CD25/100 Cells.CD4
C4696100|T201|COMP|88835-4|LNC|Influenza virus A swine origin RNA|Influenza virus A swine origin RNA
C4696101|T201|COMP|88836-2|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4696102|T201|COMP|88837-0|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4696103|T201|COMP|88843-8|LNC|Metabolic panel.dialysis patient|Metabolic panel.dialysis patient
C4696105|T201|COMP|88844-6|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4696106|T201|COMP|88845-3|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4696107|T201|COMP|88846-1|LNC|Urinary cell count CNAMTS panel|Urinary cell count CNAMTS panel
C4696109|T201|COMP|88847-9|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4696110|T201|COMP|88848-7|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4696111|T201|COMP|88849-5|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4696112|T201|COMP|88850-3|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4696123|T201|COMP|88863-6|LNC|Lung cancer antibody panel|Lung cancer antibody panel
C4696125|T201|COMP|88864-4|LNC|Microbiology CNAMTS panel|Microbiology CNAMTS panel
C4696126|T201|COMP|88865-1|LNC|Chemical XXX|Chemical XXX
C4696128|T201|COMP|88866-9|LNC|Chemical XXX|Chemical XXX
C4696129|T201|COMP|88867-7|LNC|Chemical XXX|Chemical XXX
C4696130|T201|COMP|88868-5|LNC|Veterinary toxicology panel|Veterinary toxicology panel
C4696132|T201|COMP|88869-3|LNC|Veterinary toxicology panel|Veterinary toxicology panel
C4696139|T201|COMP|88873-5|LNC|Sympathomimetics|Sympathomimetics
C4696140|T201|COMP|88874-3|LNC|Mycobacterium tuberculosis complex DNA|Mycobacterium tuberculosis complex DNA
C4696141|T201|COMP|88875-0|LNC|Measles virus genotype A vaccine strain N gene|Measles virus genotype A vaccine strain N gene
C4696143|T201|COMP|88876-8|LNC|Measles virus genotype A vaccine strain N gene|Measles virus genotype A vaccine strain N gene
C4696144|T201|COMP|88880-0|LNC|Monocyte distribution width|Monocyte distribution width
C4696146|T201|COMP|88881-8|LNC|Smith extractable nuclear D Ab|Smith extractable nuclear D Ab
C4696147|T201|COMP|88882-6|LNC|Smith extractable nuclear B Ab|Smith extractable nuclear B Ab
C4696148|T201|COMP|88888-3|LNC|Pancreatic stone protein|Pancreatic stone protein
C4696149|T201|COMP|88889-1|LNC|Middle east respiratory syndrome coronavirus RNA|Middle east respiratory syndrome coronavirus RNA
C4696150|T201|COMP|88890-9|LNC|Parainfluenza virus 1+2+3+4 RNA|Parainfluenza virus 1+2+3+4 RNA
C4696152|T201|COMP|88891-7|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA|Human coronavirus 229E+HKU1+NL63+OC43 RNA
C4696154|T201|COMP|88899-0|LNC|Adenovirus|Adenovirus
C4696155|T201|COMP|88900-6|LNC|Adenovirus|Adenovirus
C4696156|T201|COMP|88901-4|LNC|Adenovirus|Adenovirus
C4696157|T201|COMP|88902-2|LNC|Adenovirus|Adenovirus
C4696158|T201|COMP|88903-0|LNC|Influenza virus B Ab.IgG|Influenza virus B Ab.IgG
C4696159|T201|COMP|88904-8|LNC|Influenza virus A Ag|Influenza virus A Ag
C4696160|T201|COMP|88905-5|LNC|Influenza virus B Ag|Influenza virus B Ag
C4696161|T201|COMP|88906-3|LNC|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C4696162|T201|COMP|88907-1|LNC|Parainfluenza virus 2 Ag|Parainfluenza virus 2 Ag
C4696163|T201|COMP|88908-9|LNC|Parainfluenza virus 3 Ag|Parainfluenza virus 3 Ag
C4696164|T201|COMP|88909-7|LNC|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C4696165|T201|COMP|88910-5|LNC|Taenia sp DNA|Taenia sp DNA
C4696167|T201|COMP|88911-3|LNC|Taenia solium larva DNA|Taenia solium larva DNA
C4696168|T201|COMP|88912-1|LNC|Taenia solium larva DNA|Taenia solium larva DNA
C4696169|T201|COMP|88913-9|LNC|Strongyloides stercoralis DNA|Strongyloides stercoralis DNA
C4696171|T201|COMP|88914-7|LNC|Acanthamoeba sp DNA|Acanthamoeba sp DNA
C4696172|T201|COMP|88915-4|LNC|Filaria DNA|Filaria DNA
C4696174|T201|COMP|88916-2|LNC|Leishmania sp DNA|Leishmania sp DNA
C4696175|T201|COMP|88917-0|LNC|Leishmania sp DNA|Leishmania sp DNA
C4696176|T201|COMP|88918-8|LNC|Filaria DNA|Filaria DNA
C4696177|T201|COMP|88919-6|LNC|Taenia solium larva Ab.IgG|Taenia solium larva Ab.IgG
C4696178|T201|COMP|88920-4|LNC|Taenia solium larva Ag|Taenia solium larva Ag
C4696179|T201|COMP|88921-2|LNC|Echinococcus granulosus Ab|Echinococcus granulosus Ab
C4696180|T201|COMP|88922-0|LNC|Actinomyces sp identified|Actinomyces sp identified
C4696181|T201|COMP|88923-8|LNC|1,3 beta glucan|1,3 beta glucan
C4696182|T201|COMP|88924-6|LNC|Microsporidia DNA|Microsporidia DNA
C4696183|T201|COMP|88925-3|LNC|Microsporidia DNA|Microsporidia DNA
C4696184|T201|COMP|88926-1|LNC|Histoplasma capsulatum DNA|Histoplasma capsulatum DNA
C4696185|T201|COMP|88927-9|LNC|Cryptosporidium sp DNA|Cryptosporidium sp DNA
C4696186|T201|COMP|88928-7|LNC|Cryptosporidium sp DNA|Cryptosporidium sp DNA
C4696243|T201|COMP|88966-7|LNC|Hyaline casts|Hyaline casts
C4696244|T201|COMP|88967-5|LNC|Leucine crystals|Leucine crystals
C4696245|T201|COMP|88968-3|LNC|Waxy casts|Waxy casts
C4696246|T201|COMP|88969-1|LNC|Tyrosine crystals|Tyrosine crystals
C4696247|T201|COMP|88970-9|LNC|Erythrocyte casts|Erythrocyte casts
C4696248|T201|COMP|88971-7|LNC|Mixed cellular casts|Mixed cellular casts
C4696249|T201|COMP|88972-5|LNC|Broad casts|Broad casts
C4696250|T201|COMP|88973-3|LNC|Crystals.amorphous|Crystals.amorphous
C4696251|T201|COMP|88974-1|LNC|Granular casts|Granular casts
C4696252|T201|COMP|88975-8|LNC|Fatty casts|Fatty casts
C4696253|T201|COMP|88976-6|LNC|Leukocyte casts|Leukocyte casts
C4696254|T201|COMP|88977-4|LNC|Epithelial casts|Epithelial casts
C4696256|T201|COMP|88979-0|LNC|Mucus|Mucus
C4696261|T201|COMP|88985-7|LNC|Alpha-amanitin+gamma-amanitin|Alpha-amanitin+gamma-amanitin
C4696262|T201|COMP|88986-5|LNC|Elvitegravir|Elvitegravir
C4696263|T201|COMP|88987-3|LNC|Maraviroc|Maraviroc
C4696264|T201|COMP|88988-1|LNC|Melperone|Melperone
C4696265|T201|COMP|88989-9|LNC|Perazine|Perazine
C4696266|T201|COMP|88990-7|LNC|Sertindole|Sertindole
C4696267|T201|COMP|88991-5|LNC|Zotepine|Zotepine
C4696268|T201|COMP|88992-3|LNC|Ustekinumab Ab|Ustekinumab Ab
C4696269|T201|COMP|88993-1|LNC|Acute kidney injury risk|Acute kidney injury risk
C4696271|T201|COMP|88994-9|LNC|Arachidonate/Fatty acids.C14-C24|Arachidonate/Fatty acids.C14-C24
C4696273|T201|COMP|88995-6|LNC|Docosahexaenoate/Fatty acids.C14-C24|Docosahexaenoate/Fatty acids.C14-C24
C4696275|T201|COMP|88996-4|LNC|Eicosapentaenoate/Arachidonate|Eicosapentaenoate/Arachidonate
C4696277|T201|COMP|88997-2|LNC|Eicosapentaenoate/Fatty acids.C14-C24|Eicosapentaenoate/Fatty acids.C14-C24
C4696283|T201|COMP|89000-4|LNC|Ethyl glucuronide|Ethyl glucuronide
C4696284|T201|COMP|89001-2|LNC|Cancer-associated gene Ab|Cancer-associated gene Ab
C4696285|T201|COMP|89002-0|LNC|GBU4-5 Ab|GBU4-5 Ab
C4696320|T201|COMP|89523-5|LNC|Ganglioside GT1b Ab.IgG|Ganglioside GT1b Ab.IgG
C4696321|T201|COMP|89524-3|LNC|Ganglioside GM2 Ab.IgM|Ganglioside GM2 Ab.IgM
C4696322|T201|COMP|89525-0|LNC|Ganglioside GM2 Ab.IgG|Ganglioside GM2 Ab.IgG
C4696323|T201|COMP|89526-8|LNC|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C4696334|T201|COMP|89003-8|LNC|HuD Ab|HuD Ab
C4696335|T201|COMP|89004-6|LNC|Melanoma-associated antigen A4 Ab|Melanoma-associated antigen A4 Ab
C4696337|T201|COMP|89005-3|LNC|NY-ESO-1 Ab|NY-ESO-1 Ab
C4696338|T201|COMP|89006-1|LNC|p53 Ab|p53 Ab
C4696339|T201|COMP|89007-9|LNC|SOX-2 Ab|SOX-2 Ab
C4696368|T201|COMP|89040-0|LNC|Rubella virus Ab|Rubella virus Ab
C4696369|T201|COMP|89041-8|LNC|Lung cancer antibody|Lung cancer antibody
C4696371|T201|COMP|89042-6|LNC|Eszopiclone|Eszopiclone
C4696372|T201|COMP|89043-4|LNC|Zopiclone-N-oxide|Zopiclone-N-oxide
C4696373|T201|COMP|89044-2|LNC|Basic metabolic & albumin panel|Basic metabolic & albumin panel
C4696583|T201|COMP|89272-9|LNC|Oxygen saturation^during apnea|Oxygen saturation^during apnea
C4696586|T201|COMP|89276-0|LNC|Oxygen saturation^W exercise|Oxygen saturation^W exercise
C4696587|T201|COMP|89277-8|LNC|Oxygen saturation^during anesthesia|Oxygen saturation^during anesthesia
C4696616|T201|COMP|89300-8|LNC|Tapentadol glucuronide|Tapentadol glucuronide
C4696617|T201|COMP|89301-6|LNC|oxyMORphone-3-glucuronide|oxyMORphone-3-glucuronide
C4696618|T201|COMP|89302-4|LNC|Noroxymorphone|Noroxymorphone
C4696619|T201|COMP|89303-2|LNC|Noroxycodone|Noroxycodone
C4696620|T201|COMP|89304-0|LNC|Norhydrocodone|Norhydrocodone
C4696621|T201|COMP|89305-7|LNC|Norbuprenorphine-3-glucuronide|Norbuprenorphine-3-glucuronide
C4696623|T201|COMP|89306-5|LNC|Nortapentadol|Nortapentadol
C4696624|T201|COMP|89307-3|LNC|Naloxone-3-glucuronide|Naloxone-3-glucuronide
C4696625|T201|COMP|89308-1|LNC|Morphine-6-glucuronide|Morphine-6-glucuronide
C4696626|T201|COMP|89309-9|LNC|HYDROmorphone-3-glucuronide|HYDROmorphone-3-glucuronide
C4696627|T201|COMP|89310-7|LNC|Codeine-6-glucuronide|Codeine-6-glucuronide
C4696628|T201|COMP|89311-5|LNC|Cells.CD3-CD45+/100 cells|Cells.CD3-CD45+/100 cells
C4696630|T201|COMP|89312-3|LNC|Cells.CD3+CD45+|Cells.CD3+CD45+
C4696631|T201|COMP|89313-1|LNC|Cells.CD3-CD45+|Cells.CD3-CD45+
C4696635|T201|COMP|89315-6|LNC|Cells.CD4+CD25+CD45RA+CD127Low+|Cells.CD4+CD25+CD45RA+CD127Low+
C4696637|T201|COMP|89316-4|LNC|Cells.CD4+CD25+CD45RO+CD127Low+|Cells.CD4+CD25+CD45RO+CD127Low+
C4696639|T201|COMP|89317-2|LNC|Cells.CD4+CD25-CD127+|Cells.CD4+CD25-CD127+
C4696641|T201|COMP|89318-0|LNC|Cells.CD25-CD127+/100 Cells.CD4|Cells.CD25-CD127+/100 Cells.CD4
C4696643|T201|COMP|89319-8|LNC|Cells.CD25+CD45RA+CD127Low+/100 Cells.CD4|Cells.CD25+CD45RA+CD127Low+/100 Cells.CD4
C4696645|T201|COMP|89320-6|LNC|Cells.CD25+CD45RO+CD127Low+/100 Cells.CD4|Cells.CD25+CD45RO+CD127Low+/100 Cells.CD4
C4696647|T201|COMP|89321-4|LNC|Buprenorphine-3-glucuronide|Buprenorphine-3-glucuronide
C4696649|T201|COMP|89322-2|LNC|Norbuprenorphine-3-glucuronide|Norbuprenorphine-3-glucuronide
C4696650|T201|COMP|89323-0|LNC|APOB gene targeted mutation analysis|APOB gene targeted mutation analysis
C4696652|T201|COMP|89324-8|LNC|Insulin.intact|Insulin.intact
C4696654|T201|COMP|89325-5|LNC|Cells.CD3+CD8+CD28+HLA DR+|Cells.CD3+CD8+CD28+HLA DR+
C4696656|T201|COMP|89326-3|LNC|Cells.CD3+CD4+CD28+HLA DR+|Cells.CD3+CD4+CD28+HLA DR+
C4696658|T201|COMP|89332-1|LNC|Cells.CD28+HLA DR+/100 Cells.CD3+CD8+|Cells.CD28+HLA DR+/100 Cells.CD3+CD8+
C4696660|T201|COMP|89333-9|LNC|Cells.CD28+HLA DR+/100 Cells.CD3+CD4+|Cells.CD28+HLA DR+/100 Cells.CD3+CD4+
C4696662|T201|COMP|89334-7|LNC|Cells.CD27-CD45RO+CD62L-CCR7-/100 Cells.CD3+CD8+|Cells.CD27-CD45RO+CD62L-CCR7-/100 Cells.CD3+CD8+
C4696664|T201|COMP|89335-4|LNC|Cells.CD27+CD45RO+CD62L+CCR7+/100 Cells.CD3+CD8+|Cells.CD27+CD45RO+CD62L+CCR7+/100 Cells.CD3+CD8+
C4696666|T201|COMP|89336-2|LNC|Cells.CD45RO/100 Cells.CD3+CD8+|Cells.CD45RO/100 Cells.CD3+CD8+
C4696668|T201|COMP|89337-0|LNC|Cells.CD27-CD45RO+CD62L-CCR7-/100 Cells.CD3+CD4+|Cells.CD27-CD45RO+CD62L-CCR7-/100 Cells.CD3+CD4+
C4696670|T201|COMP|89338-8|LNC|Cells.CD27+CD45RO+CD62L+CCR7+/100 Cells.CD3+CD4+|Cells.CD27+CD45RO+CD62L+CCR7+/100 Cells.CD3+CD4+
C4696672|T201|COMP|89339-6|LNC|Cells.CD27+CD62L+/100 Cells.CD3+CD8+|Cells.CD27+CD62L+/100 Cells.CD3+CD8+
C4696674|T201|COMP|89340-4|LNC|Cells.CD27+CD62L+/100 Cells.CD3+CD4+|Cells.CD27+CD62L+/100 Cells.CD3+CD4+
C4696676|T201|COMP|89341-2|LNC|Cells.CD38+IgM+/100 Cells.CD19|Cells.CD38+IgM+/100 Cells.CD19
C4696678|T201|COMP|89342-0|LNC|Babesia sp 18S rRNA|Babesia sp 18S rRNA
C4696680|T201|COMP|89343-8|LNC|Cells.CD19+CD38+IgM-|Cells.CD19+CD38+IgM-
C4696682|T201|COMP|89344-6|LNC|Cells.CD38+IgM-/100 Cells.CD19|Cells.CD38+IgM-/100 Cells.CD19
C4696684|T201|COMP|89345-3|LNC|Cells.CD19+IgM+|Cells.CD19+IgM+
C4696685|T201|COMP|89346-1|LNC|Cells.IgM/100 Cells.CD19|Cells.IgM/100 Cells.CD19
C4696687|T201|COMP|89347-9|LNC|Cells.CD19+CD27+IgD-IgM+|Cells.CD19+CD27+IgD-IgM+
C4696689|T201|COMP|89348-7|LNC|Cells.CD27+IgD-IgM+/100 Cells.CD19|Cells.CD27+IgD-IgM+/100 Cells.CD19
C4696691|T201|COMP|89349-5|LNC|Cells.CD19+CD27+IgD-IgM-|Cells.CD19+CD27+IgD-IgM-
C4696693|T201|COMP|89350-3|LNC|Cells.CD27+IgD-IgM-/100 Cells.CD19|Cells.CD27+IgD-IgM-/100 Cells.CD19
C4696695|T201|COMP|89351-1|LNC|Cells.CD19+CD27+IgD+IgM+|Cells.CD19+CD27+IgD+IgM+
C4696697|T201|COMP|89352-9|LNC|Cells.CD27+IgD+IgM+/100 Cells.CD19|Cells.CD27+IgD+IgM+/100 Cells.CD19
C4696699|T201|COMP|89353-7|LNC|Cells.CD19+CD27+|Cells.CD19+CD27+
C4696701|T201|COMP|89354-5|LNC|Cells.CD19+CD21-|Cells.CD19+CD21-
C4696703|T201|COMP|89355-2|LNC|Cells.CD21-/100 Cells.CD19|Cells.CD21-/100 Cells.CD19
C4696705|T201|COMP|89356-0|LNC|Cells.CD21/100 Cells.CD19|Cells.CD21/100 Cells.CD19
C4696707|T201|COMP|89357-8|LNC|Cells.CD19+CD38+IgM+|Cells.CD19+CD38+IgM+
C4696709|T201|COMP|89358-6|LNC|Cells.CD27/100 Cells.CD19|Cells.CD27/100 Cells.CD19
C4696711|T201|COMP|89359-4|LNC|Hepatitis C virus Ab.IgG|Hepatitis C virus Ab.IgG
C4696712|T201|COMP|89360-2|LNC|Cells.CD45RA/100 Cells.CD4|Cells.CD45RA/100 Cells.CD4
C4696714|T201|COMP|89362-8|LNC|Cells.CD45RO/100 Cells.CD4|Cells.CD45RO/100 Cells.CD4
C4696716|T201|COMP|89363-6|LNC|Cholinesterase|Cholinesterase
C4696717|T201|COMP|89364-4|LNC|Hemoglobin.free|Hemoglobin.free
C4696718|T201|COMP|89365-1|LNC|HIV 1 & 2 Ab panel|HIV 1 & 2 Ab panel
C4696724|T201|COMP|89368-5|LNC|Zika virus non-structural protein 1 Ab.IgM panel|Zika virus non-structural protein 1 Ab.IgM panel
C4696726|T201|COMP|89369-3|LNC|Zika virus non-structural protein 1 Ab.IgM|Zika virus non-structural protein 1 Ab.IgM
C4696728|T201|COMP|89370-1|LNC|Zika virus non-structural protein 1 Ab.IgM|Zika virus non-structural protein 1 Ab.IgM
C4696733|T201|COMP|89373-5|LNC|Hepatitis A virus genotype|Hepatitis A virus genotype
C4696735|T201|COMP|89374-3|LNC|HIV 1 Ab|HIV 1 Ab
C4696877|T201|COMP|89480-8|LNC|Azithromycin|Azithromycin
C4696878|T201|COMP|89485-7|LNC|Clarithromycin|Clarithromycin
C4696879|T201|COMP|89486-5|LNC|Mycobacterial susceptibility panel|Mycobacterial susceptibility panel
C4696880|T201|COMP|89487-3|LNC|Fluoroquinolone|Fluoroquinolone
C4696881|T201|COMP|89488-1|LNC|Isoniazid|Isoniazid
C4696882|T201|COMP|89489-9|LNC|rifAMPin|rifAMPin
C4696883|T201|COMP|89490-7|LNC|Aminoglycoside|Aminoglycoside
C4696884|T201|COMP|89491-5|LNC|Ethambutol|Ethambutol
C4696892|T201|COMP|89500-3|LNC|Sulfatide Ab.IgG|Sulfatide Ab.IgG
C4696894|T201|COMP|89502-9|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C4696895|T201|COMP|89503-7|LNC|RNA polymerase III Ab|RNA polymerase III Ab
C4696896|T201|COMP|89504-5|LNC|Ribosomal Ab|Ribosomal Ab
C4696897|T201|COMP|89505-2|LNC|Proteinase 3 Ab|Proteinase 3 Ab
C4696898|T201|COMP|89506-0|LNC|Nucleosome Ab|Nucleosome Ab
C4696899|T201|COMP|89507-8|LNC|Myeloperoxidase Ab|Myeloperoxidase Ab
C4696900|T201|COMP|89508-6|LNC|Intrinsic factor Ab|Intrinsic factor Ab
C4696901|T201|COMP|89509-4|LNC|Ganglioside GT1a Ab.IgG+IgM|Ganglioside GT1a Ab.IgG+IgM
C4696902|T201|COMP|89510-2|LNC|Ganglioside GM3 Ab.IgM|Ganglioside GM3 Ab.IgM
C4696903|T201|COMP|89511-0|LNC|Ganglioside GM3 Ab.IgG+IgM|Ganglioside GM3 Ab.IgG+IgM
C4696904|T201|COMP|89512-8|LNC|Ganglioside GD3 Ab.IgG+IgM|Ganglioside GD3 Ab.IgG+IgM
C4696905|T201|COMP|89513-6|LNC|RNA polymerase III Ab|RNA polymerase III Ab
C4696906|T201|COMP|89514-4|LNC|Glomerular basement membrane Ab|Glomerular basement membrane Ab
C4696907|T201|COMP|89515-1|LNC|Ganglioside GT1b Ab.IgM|Ganglioside GT1b Ab.IgM
C4696908|T201|COMP|89516-9|LNC|Ganglioside GT1b Ab.IgG+IgM|Ganglioside GT1b Ab.IgG+IgM
C4696909|T201|COMP|89517-7|LNC|Ganglioside GM2 Ab.IgG+IgM|Ganglioside GM2 Ab.IgG+IgM
C4696910|T201|COMP|89518-5|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C4696911|T201|COMP|89519-3|LNC|Ganglioside GM1 Ab.IgG+IgM|Ganglioside GM1 Ab.IgG+IgM
C4696912|T201|COMP|89520-1|LNC|Actin.smooth muscle Ab|Actin.smooth muscle Ab
C4696913|T201|COMP|89521-9|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C4696914|T201|COMP|89522-7|LNC|Ganglioside GM3 Ab.IgG|Ganglioside GM3 Ab.IgG
C4696915|T201|COMP|89527-6|LNC|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C4696916|T201|COMP|89528-4|LNC|Nucleosome Ab|Nucleosome Ab
C4696917|T201|COMP|89529-2|LNC|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C4696918|T201|COMP|89530-0|LNC|Histone Ab|Histone Ab
C4696919|T201|COMP|89531-8|LNC|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C4696920|T201|COMP|89532-6|LNC|Sjogrens syndrome-A extractable nuclear 52kD Ab|Sjogrens syndrome-A extractable nuclear 52kD Ab
C4696921|T201|COMP|89533-4|LNC|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C4696922|T201|COMP|89534-2|LNC|Ribosomal P Ab|Ribosomal P Ab
C4696923|T201|COMP|89535-9|LNC|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C4696924|T201|COMP|89536-7|LNC|PM-SCL extractable nuclear Ab|PM-SCL extractable nuclear Ab
C4696925|T201|COMP|89537-5|LNC|PCNA extractable nuclear Ab|PCNA extractable nuclear Ab
C4696926|T201|COMP|89538-3|LNC|Neuronal nuclear type 2 Ab|Neuronal nuclear type 2 Ab
C4696927|T201|COMP|89539-1|LNC|Mitochondria M2 Ab|Mitochondria M2 Ab
C4696928|T201|COMP|89540-9|LNC|Ganglioside GM1 Ab.IgM|Ganglioside GM1 Ab.IgM
C4696929|T201|COMP|89541-7|LNC|Ganglioside GM1 Ab.IgG|Ganglioside GM1 Ab.IgG
C4696930|T201|COMP|89542-5|LNC|Centromere protein B Ab|Centromere protein B Ab
C4696958|T201|COMP|89575-5|LNC|Troponin T.cardiac|Troponin T.cardiac
C4696959|T201|COMP|89576-3|LNC|Troponin T.cardiac panel|Troponin T.cardiac panel
C4696961|T201|COMP|89577-1|LNC|Troponin I.cardiac panel|Troponin I.cardiac panel
C4696963|T201|COMP|89578-9|LNC|Troponin I.cardiac|Troponin I.cardiac
C4696964|T201|COMP|89579-7|LNC|Troponin I.cardiac|Troponin I.cardiac
C4696967|T201|COMP|89585-4|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C4696968|T201|COMP|89586-2|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C4696969|T201|COMP|89587-0|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C4696970|T201|COMP|89588-8|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C4696971|T201|COMP|89589-6|LNC|Varicella zoster virus Ag|Varicella zoster virus Ag
C4696972|T201|COMP|89590-4|LNC|Zika virus Ab.IgG|Zika virus Ab.IgG
C4696974|T201|COMP|89591-2|LNC|Zika virus Ab.IgM|Zika virus Ab.IgM
C4696975|T201|COMP|89592-0|LNC|Bartonella quintana DNA|Bartonella quintana DNA
C4696976|T201|COMP|89593-8|LNC|Bartonella sp DNA|Bartonella sp DNA
C4696977|T201|COMP|89594-6|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C4696978|T201|COMP|89595-3|LNC|Legionella pneumophila Ag|Legionella pneumophila Ag
C4696979|T201|COMP|89596-1|LNC|Listeria monocytogenes DNA|Listeria monocytogenes DNA
C4696980|T201|COMP|89597-9|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C4696981|T201|COMP|89598-7|LNC|Mycoplasma hominis DNA|Mycoplasma hominis DNA
C4696982|T201|COMP|89599-5|LNC|Toxoplasma gondii|Toxoplasma gondii
C4721465|T201|COMP|1307-8|LNC|D NOS Ab|D NOS Ab
C4721466|T201|COMP|1308-6|LNC|D NOS Ab|D NOS Ab
C4721467|T201|COMP|1310-2|LNC|D NOS Ag|D NOS Ag
C4721468|T201|COMP|1311-0|LNC|D NOS Ag|D NOS Ag
C4721469|T201|COMP|1312-8|LNC|D NOS Ag|D NOS Ag
C4721470|T201|COMP|1066-0|LNC|I NOS Ag|I NOS Ag
C4724106|T201|COMP|90431-8|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4724115|T201|COMP|90428-4|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4724291|T201|COMP|90763-4|LNC|HEDIS 2019-2020 Value Set - Chlamydia Tests|HEDIS 2019-2020 Value Set - Chlamydia Tests
C4724293|T201|COMP|90984-6|LNC|HEDIS 2019-2020 Value Set - PSA Test Exclusion|HEDIS 2019-2020 Value Set - PSA Test Exclusion
C4724295|T201|COMP|90766-7|LNC|HEDIS 2019 Value Sets|HEDIS 2019 Value Sets
C4724324|T201|COMP|90765-9|LNC|HEDIS 2019 Value Set - Rh|HEDIS 2019 Value Set - Rh
C4724346|T201|COMP|90056-3|LNC|Date and time lab result reported|Date and time lab result reported
C4724411|T201|COMP|90257-7|LNC|GLA gene full mutation analysis|GLA gene full mutation analysis
C4724482|T201|COMP|90777-4|LNC|HEDIS 2019 Value Set - Cytomegalovirus Antibody|HEDIS 2019 Value Set - Cytomegalovirus Antibody
C4724483|T201|COMP|90996-0|LNC|HEDIS 2019-2020 Value Set - Glucose Tests|HEDIS 2019-2020 Value Set - Glucose Tests
C4724485|T201|COMP|90997-8|LNC|HEDIS 2019-2020 Value Set - Group A Strep Tests|HEDIS 2019-2020 Value Set - Group A Strep Tests
C4724487|T201|COMP|90988-7|LNC|HEDIS 2019-2020 Value Set - HPV Tests|HEDIS 2019-2020 Value Set - HPV Tests
C4724489|T201|COMP|90983-8|LNC|HEDIS 2019-2020 Value Set - PSA Tests|HEDIS 2019-2020 Value Set - PSA Tests
C4724490|T201|COMP|90776-6|LNC|HEDIS 2019 Value Set - Rubella Antibody|HEDIS 2019 Value Set - Rubella Antibody
C4724491|T201|COMP|90986-1|LNC|HEDIS 2019 Value Set - Serum Potassium|HEDIS 2019 Value Set - Serum Potassium
C4724493|T201|COMP|90764-2|LNC|HEDIS 2019 Value Set - Toxoplasma Antibody|HEDIS 2019 Value Set - Toxoplasma Antibody
C4724494|T201|COMP|90989-5|LNC|HEDIS 2019 Value Set - Urine Protein Tests|HEDIS 2019 Value Set - Urine Protein Tests
C4724514|T201|COMP|90947-3|LNC|Pathology case identifier|Pathology case identifier
C4724567|T201|COMP|90101-7|LNC|Internal control result|Internal control result
C4724570|T201|COMP|90426-8|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4724571|T201|COMP|90427-6|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4724704|T201|COMP|90369-0|LNC|Sample collection timing related to drug dose|Sample collection timing related to drug dose
C4738069|T201|COMP|90993-7|LNC|Iothalamate clearance panel|Iothalamate clearance panel
C4738090|T201|COMP|90880-6|LNC|Arachis hypogaea recombinant (rAra h) 6 Ab.IgE|Arachis hypogaea recombinant (rAra h) 6 Ab.IgE
C4738153|T201|COMP|91105-7|LNC|Cholesterol.in LDL 1|Cholesterol.in LDL 1
C4738155|T201|COMP|91106-5|LNC|Cholesterol.in LDL 2|Cholesterol.in LDL 2
C4738157|T201|COMP|91107-3|LNC|Cholesterol.in LDL 3|Cholesterol.in LDL 3
C4738159|T201|COMP|91108-1|LNC|Cholesterol.in LDL 4|Cholesterol.in LDL 4
C4738161|T201|COMP|91109-9|LNC|Cholesterol.in LDL 5|Cholesterol.in LDL 5
C4738163|T201|COMP|91110-7|LNC|Cholesterol.in LDL 6|Cholesterol.in LDL 6
C4738165|T201|COMP|91111-5|LNC|Cholesterol.in LDL 7|Cholesterol.in LDL 7
C4738167|T201|COMP|91112-3|LNC|Cholesterol.in LDL 1|Cholesterol.in LDL 1
C4738168|T201|COMP|91113-1|LNC|Cholesterol.in LDL 2|Cholesterol.in LDL 2
C4738169|T201|COMP|91114-9|LNC|Cholesterol.in LDL 3|Cholesterol.in LDL 3
C4738170|T201|COMP|91115-6|LNC|Cholesterol.in LDL 4|Cholesterol.in LDL 4
C4738171|T201|COMP|91116-4|LNC|Cholesterol.in LDL 5|Cholesterol.in LDL 5
C4738172|T201|COMP|91117-2|LNC|Cholesterol.in LDL 6|Cholesterol.in LDL 6
C4738173|T201|COMP|91118-0|LNC|Cholesterol.in LDL 7|Cholesterol.in LDL 7
C4738175|T201|COMP|91120-6|LNC|Antithrombin|Antithrombin
C4738180|T201|COMP|91129-7|LNC|Clot strength.adenosine diphosphate induced|Clot strength.adenosine diphosphate induced
C4738182|T201|COMP|91130-5|LNC|Hantavirus RNA|Hantavirus RNA
C4738183|T201|COMP|91131-3|LNC|Rhinovirus RNA|Rhinovirus RNA
C4738184|T201|COMP|91132-1|LNC|Measles virus RNA|Measles virus RNA
C4738185|T201|COMP|91134-7|LNC|Sexually transmitted pathogens panel|Sexually transmitted pathogens panel
C4738187|T201|COMP|91135-4|LNC|Acanthocytes|Acanthocytes
C4738188|T201|COMP|91136-2|LNC|Lipoprotein metabolism panel|Lipoprotein metabolism panel
C4738190|T201|COMP|91137-0|LNC|ITPA gene.g.9330C>A|ITPA gene.g.9330C>A
C4738194|T201|COMP|90736-0|LNC|Cells.CD14-FLAER-/100 cells.CD33|Cells.CD14-FLAER-/100 cells.CD33
C4738196|T201|COMP|90737-8|LNC|Cells.CD24-FLAER-/100 cells.CD15|Cells.CD24-FLAER-/100 cells.CD15
C4738198|T201|COMP|90738-6|LNC|Erythrocytes.CD59 complete loss/100 Cells.235a|Erythrocytes.CD59 complete loss/100 Cells.235a
C4738202|T201|COMP|90740-2|LNC|Aggressive prostate cancer risk|Aggressive prostate cancer risk
C4738204|T201|COMP|90741-0|LNC|Parathyrin.1-84|Parathyrin.1-84
C4738206|T201|COMP|90742-8|LNC|Bovine Mullerian inhibiting substance|Bovine Mullerian inhibiting substance
C4738208|T201|COMP|90743-6|LNC|CYBB gene full & NCF1 gene c.75_76delGT analysis|CYBB gene full & NCF1 gene c.75_76delGT analysis
C4738290|T201|COMP|90992-9|LNC|Monoclonal gammopathy panel|Monoclonal gammopathy panel
C4738294|T201|COMP|90994-5|LNC|Iothalamate clearance|Iothalamate clearance
C4738295|T201|COMP|90995-2|LNC|Iothalamate clearance/Body surface area|Iothalamate clearance/Body surface area
C4738335|T201|COMP|90831-9|LNC|Leucine-rich glioma-inactivated protein 1 Ab|Leucine-rich glioma-inactivated protein 1 Ab
C4738336|T201|COMP|90832-7|LNC|Ma+Ta Ab|Ma+Ta Ab
C4738337|T201|COMP|90833-5|LNC|Ma+Ta Ab|Ma+Ta Ab
C4738338|T201|COMP|90834-3|LNC|Myelin Ab|Myelin Ab
C4738339|T201|COMP|90835-0|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C4738343|T201|COMP|90909-3|LNC|Arachidonate/Eicosapentaenoate|Arachidonate/Eicosapentaenoate
C4738345|T201|COMP|90910-1|LNC|Fatty acids.omega 6/Fatty acids.omega 3|Fatty acids.omega 6/Fatty acids.omega 3
C4738348|T201|COMP|90912-7|LNC|Eicosapentaenoate/Fatty acids.C14-C22|Eicosapentaenoate/Fatty acids.C14-C22
C4738350|T201|COMP|90913-5|LNC|Docosapentaenate w3/Fatty acids.C14-C22|Docosapentaenate w3/Fatty acids.C14-C22
C4738352|T201|COMP|90914-3|LNC|Docosahexaenoate/Fatty acids.C14-C22|Docosahexaenoate/Fatty acids.C14-C22
C4738354|T201|COMP|90915-0|LNC|Arachidonate+Linoleate/Fatty acids.C14-C22|Arachidonate+Linoleate/Fatty acids.C14-C22
C4738356|T201|COMP|90916-8|LNC|Arachidonate/Fatty acids.C14-C22|Arachidonate/Fatty acids.C14-C22
C4738358|T201|COMP|90917-6|LNC|Linoleate/Fatty acids.C14-C22|Linoleate/Fatty acids.C14-C22
C4738360|T201|COMP|90918-4|LNC|Fatty acid omega-3 & omega-6 panel|Fatty acid omega-3 & omega-6 panel
C4738365|T201|COMP|1045-4|LNC|H NOS Ab|H NOS Ab
C4738366|T201|COMP|1046-2|LNC|H NOS Ab|H NOS Ab
C4738367|T201|COMP|1047-0|LNC|H NOS Ab|H NOS Ab
C4738368|T201|COMP|1061-1|LNC|I NOS Ab|I NOS Ab
C4738369|T201|COMP|1062-9|LNC|I NOS Ab|I NOS Ab
C4738370|T201|COMP|1063-7|LNC|I NOS Ab|I NOS Ab
C4738374|T201|COMP|1127-0|LNC|L little e NOS Ab|L little e NOS Ab
C4738375|T201|COMP|1128-8|LNC|L little e NOS Ab|L little e NOS Ab
C4738376|T201|COMP|1238-5|LNC|M NOS Ab|M NOS Ab
C4738377|T201|COMP|1239-3|LNC|M NOS Ab|M NOS Ab
C4738378|T201|COMP|1240-1|LNC|M NOS Ab|M NOS Ab
C4738379|T201|COMP|1241-9|LNC|M NOS Ag|M NOS Ag
C4738380|T201|COMP|1242-7|LNC|M NOS Ag|M NOS Ag
C4738381|T201|COMP|1243-5|LNC|M NOS Ag|M NOS Ag
C4738383|T201|COMP|1262-5|LNC|N NOS Ab|N NOS Ab
C4738384|T201|COMP|1263-3|LNC|N NOS Ab|N NOS Ab
C4738385|T201|COMP|1264-1|LNC|N NOS Ab|N NOS Ab
C4738386|T201|COMP|1265-8|LNC|N NOS Ag|N NOS Ag
C4738387|T201|COMP|1266-6|LNC|N NOS Ag|N NOS Ag
C4738388|T201|COMP|1267-4|LNC|N NOS Ag|N NOS Ag
C4738389|T201|COMP|1280-7|LNC|P NOS Ab|P NOS Ab
C4738390|T201|COMP|1281-5|LNC|P NOS Ab|P NOS Ab
C4738391|T201|COMP|1282-3|LNC|P NOS Ab|P NOS Ab
C4738396|T201|COMP|90920-0|LNC|Lysophosphatidylcholine(20:0)|Lysophosphatidylcholine(20:0)
C4738469|T201|COMP|90921-8|LNC|Lysophosphatidylcholine(22:0)|Lysophosphatidylcholine(22:0)
C4738478|T201|COMP|90822-8|LNC|CV2 Ab|CV2 Ab
C4738479|T201|COMP|90850-9|LNC|cefTAZidime 1.0 ug/mL|cefTAZidime 1.0 ug/mL
C4738481|T201|COMP|90851-7|LNC|GJB2 gene full mutation analysis|GJB2 gene full mutation analysis
C4738510|T201|COMP|90223-9|LNC|Neutrophils.immature/Neutrophils.total|Neutrophils.immature/Neutrophils.total
C4738512|T201|COMP|90224-7|LNC|Thyroxine & Thyroxine.free panel|Thyroxine & Thyroxine.free panel
C4738516|T201|COMP|90226-2|LNC|Nicotine & Cotinine panel|Nicotine & Cotinine panel
C4738517|T201|COMP|90237-9|LNC|Phenylacetylcarnitine (PheC2)|Phenylacetylcarnitine (PheC2)
C4738540|T201|COMP|90452-4|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C4738541|T201|COMP|90453-2|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C4738542|T201|COMP|90454-0|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C4738543|T201|COMP|90455-7|LNC|Influenza virus A & B RNA panel|Influenza virus A & B RNA panel
C4738544|T201|COMP|90456-5|LNC|Influenza virus A & B RNA panel|Influenza virus A & B RNA panel
C4738545|T201|COMP|90457-3|LNC|Influenza virus A & B RNA panel|Influenza virus A & B RNA panel
C4738546|T201|COMP|90458-1|LNC|Actinomyces sp identified|Actinomyces sp identified
C4738547|T201|COMP|90459-9|LNC|Yellow fever virus RNA|Yellow fever virus RNA
C4738548|T201|COMP|90460-7|LNC|Hepatitis E virus RNA|Hepatitis E virus RNA
C4738549|T201|COMP|90461-5|LNC|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C4738550|T201|COMP|90462-3|LNC|Zika virus RNA|Zika virus RNA
C4738551|T201|COMP|90463-1|LNC|Adenovirus DNA|Adenovirus DNA
C4738552|T201|COMP|90464-9|LNC|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C4738574|T201|COMP|90922-6|LNC|Lysophosphatidylcholine(24:0)|Lysophosphatidylcholine(24:0)
C4738576|T201|COMP|90923-4|LNC|Lysophosphatidylcholine(26:0)|Lysophosphatidylcholine(26:0)
C4738579|T201|COMP|90784-0|LNC|Cystinuria panel|Cystinuria panel
C4738595|T201|COMP|89964-1|LNC|Ziprasidone|Ziprasidone
C4738597|T201|COMP|89965-8|LNC|Trifluoperazine|Trifluoperazine
C4738598|T201|COMP|89966-6|LNC|Norquetiapine|Norquetiapine
C4738599|T201|COMP|89967-4|LNC|Norquetiapine|Norquetiapine
C4738600|T201|COMP|89968-2|LNC|Norolanzapine|Norolanzapine
C4738601|T201|COMP|89969-0|LNC|Norolanzapine|Norolanzapine
C4738602|T201|COMP|89970-8|LNC|Molindone|Molindone
C4738634|T201|COMP|90042-3|LNC|Borrelia sp DNA|Borrelia sp DNA
C4738635|T201|COMP|90043-1|LNC|t(14;20)(q32;q12)(IGH,MAFB) fusion transcript|t(14;20)(q32;q12)(IGH,MAFB) fusion transcript
C4738637|T201|COMP|90044-9|LNC|Epithelial cells.renal|Epithelial cells.renal
C4738638|T201|COMP|90045-6|LNC|Treatment history of specimen|Treatment history of specimen
C4738676|T201|COMP|90823-6|LNC|Dipeptidyl aminopeptidase-like protein 6 Ab|Dipeptidyl aminopeptidase-like protein 6 Ab
C4738826|T201|COMP|90360-9|LNC|Trimethylamine N-oxide|Trimethylamine N-oxide
C4738827|T201|COMP|90361-7|LNC|Chlamydia trachomatis L1 Ab.IgA|Chlamydia trachomatis L1 Ab.IgA
C4738843|T201|COMP|89643-1|LNC|Bacteria identified|Bacteria identified
C4738844|T201|COMP|89644-9|LNC|Bacteria identified|Bacteria identified
C4738848|T201|COMP|90327-8|LNC|Porcine circovirus type 2d DNA|Porcine circovirus type 2d DNA
C4738850|T201|COMP|90328-6|LNC|Porcine circovirus type 3 DNA|Porcine circovirus type 3 DNA
C4738852|T201|COMP|90797-2|LNC|Thyroxine^2H post dose levothyroxine|Thyroxine^2H post dose levothyroxine
C4738866|T201|COMP|89655-5|LNC|Virus identified|Virus identified
C4738867|T201|COMP|89656-3|LNC|Fungus identified|Fungus identified
C4738873|T201|COMP|89632-4|LNC|Toxoplasma gondii|Toxoplasma gondii
C4738875|T201|COMP|89633-2|LNC|Actinomyces sp identified|Actinomyces sp identified
C4738876|T201|COMP|89634-0|LNC|Actinomyces sp identified|Actinomyces sp identified
C4738878|T201|COMP|89640-7|LNC|Chlamydophila pneumoniae Ab.IgM|Chlamydophila pneumoniae Ab.IgM
C4738879|T201|COMP|89641-5|LNC|Chlamydophila pneumoniae Ab.IgG|Chlamydophila pneumoniae Ab.IgG
C4738880|T201|COMP|89642-3|LNC|Corynebacterium diphtheriae toxin Ab.IgG|Corynebacterium diphtheriae toxin Ab.IgG
C4738881|T201|COMP|90238-7|LNC|Salicylcarnitine|Salicylcarnitine
C4738883|T201|COMP|90236-1|LNC|Keratan sulfate|Keratan sulfate
C4738884|T201|COMP|89648-0|LNC|Chlamydia trachomatis|Chlamydia trachomatis
C4738885|T201|COMP|89653-0|LNC|Parainfluenza virus identified|Parainfluenza virus identified
C4738886|T201|COMP|89654-8|LNC|Parainfluenza virus identified|Parainfluenza virus identified
C4738889|T201|COMP|90246-0|LNC|Bacterial whole genome|Bacterial whole genome
C4738902|T201|COMP|90080-3|LNC|Bictegravir|Bictegravir
C4738903|T201|COMP|90247-8|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C4738921|T201|COMP|90048-0|LNC|Somatotropin binding protein|Somatotropin binding protein
C4738924|T201|COMP|90900-2|LNC|HIV 1 proviral DNA integrase gene|HIV 1 proviral DNA integrase gene
C4738931|T201|COMP|90039-9|LNC|ABO & Rh group^post transfusion reaction|ABO & Rh group^post transfusion reaction
C4738934|T201|COMP|90041-5|LNC|Collection setting|Collection setting
C4738948|T201|COMP|90888-9|LNC|Porcine circovirus type 3 DNA|Porcine circovirus type 3 DNA
C4738949|T201|COMP|90889-7|LNC|Porcine circovirus type 2 Ab.IgG|Porcine circovirus type 2 Ab.IgG
C4738956|T201|COMP|90002-7|LNC|Candida auris|Candida auris
C4738957|T201|COMP|90003-5|LNC|Acinetobacter sp identified|Acinetobacter sp identified
C4738959|T201|COMP|90323-7|LNC|Influenza virus A Ab/Positive control|Influenza virus A Ab/Positive control
C4738961|T201|COMP|90324-5|LNC|Mycoplasma hyopneumoniae DNA|Mycoplasma hyopneumoniae DNA
C4738962|T201|COMP|90836-8|LNC|Neuronal nuclear type 3 Ab|Neuronal nuclear type 3 Ab
C4738964|T201|COMP|90828-5|LNC|Glial nuclear type 1 Ab|Glial nuclear type 1 Ab
C4738967|T201|COMP|89971-6|LNC|8-Hydroxyloxapine|8-Hydroxyloxapine
C4738968|T201|COMP|89972-4|LNC|Loxapine|Loxapine
C4738969|T201|COMP|89973-2|LNC|7-Hydroxyfluphenazine|7-Hydroxyfluphenazine
C4738970|T201|COMP|89974-0|LNC|7-Hydroxyfluphenazine|7-Hydroxyfluphenazine
C4738977|T201|COMP|89992-2|LNC|Hydroxybupropion|Hydroxybupropion
C4738985|T201|COMP|90830-1|LNC|Leucine-rich glioma-inactivated protein 1 Ab|Leucine-rich glioma-inactivated protein 1 Ab
C4738999|T201|COMP|90886-3|LNC|Influenza virus B RNA|Influenza virus B RNA
C4739000|T201|COMP|90887-1|LNC|Porcine circovirus type 3 ORF2 gene|Porcine circovirus type 3 ORF2 gene
C4739003|T201|COMP|90890-5|LNC|Benzodiazepines panel|Benzodiazepines panel
C4739004|T201|COMP|90891-3|LNC|Estradiol^2H post XXX challenge|Estradiol^2H post XXX challenge
C4739005|T201|COMP|90892-1|LNC|Borrelia sp panel|Borrelia sp panel
C4739007|T201|COMP|90893-9|LNC|Borrelia burgdorferi bba64 gene|Borrelia burgdorferi bba64 gene
C4739009|T201|COMP|90894-7|LNC|Noroxymorphone|Noroxymorphone
C4739067|T201|COMP|89635-7|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C4739068|T201|COMP|89636-5|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C4739069|T201|COMP|89637-3|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C4739070|T201|COMP|89638-1|LNC|Nocardia sp identified|Nocardia sp identified
C4739071|T201|COMP|89639-9|LNC|Nocardia sp identified|Nocardia sp identified
C4739110|T201|COMP|89873-4|LNC|Unique identifier|Unique identifier
C4739125|T201|COMP|90902-8|LNC|HIV 1 RNA reverse transcriptase gene|HIV 1 RNA reverse transcriptase gene
C4739132|T201|COMP|90785-7|LNC|Cystinuria panel|Cystinuria panel
C4739135|T201|COMP|90779-0|LNC|Adalimumab Ab|Adalimumab Ab
C4739136|T201|COMP|90798-0|LNC|Thyroxine^3H post dose levothyroxine|Thyroxine^3H post dose levothyroxine
C4739137|T201|COMP|90749-3|LNC|4-Hydroxyatomoxetine|4-Hydroxyatomoxetine
C4739143|T201|COMP|90829-3|LNC|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C4739145|T201|COMP|89691-0|LNC|Pseudocasts|Pseudocasts
C4739159|T201|COMP|91138-8|LNC|ITPA gene.g.9381A>C|ITPA gene.g.9381A>C
C4739165|T201|COMP|89861-9|LNC|BRAF gene.p.Val600Lys|BRAF gene.p.Val600Lys
C4739181|T201|COMP|89975-7|LNC|Norclozapine|Norclozapine
C4739182|T201|COMP|89976-5|LNC|7-Hydroxychlorpromazine|7-Hydroxychlorpromazine
C4739183|T201|COMP|89977-3|LNC|7-Hydroxychlorpromazine|7-Hydroxychlorpromazine
C4739184|T201|COMP|89978-1|LNC|ARIPiprazole|ARIPiprazole
C4739185|T201|COMP|89979-9|LNC|Ziprasidone|Ziprasidone
C4739186|T201|COMP|89980-7|LNC|Thiothixene|Thiothixene
C4739187|T201|COMP|89981-5|LNC|QUEtiapine|QUEtiapine
C4739188|T201|COMP|89982-3|LNC|9-Hydroxyrisperidone|9-Hydroxyrisperidone
C4739189|T201|COMP|89983-1|LNC|OLANZapine|OLANZapine
C4739190|T201|COMP|89984-9|LNC|Molindone|Molindone
C4739191|T201|COMP|89985-6|LNC|ARIPiprazole|ARIPiprazole
C4739192|T201|COMP|89986-4|LNC|Vortioxetine|Vortioxetine
C4739193|T201|COMP|89987-2|LNC|Vortioxetine|Vortioxetine
C4739194|T201|COMP|89988-0|LNC|Vilazodone|Vilazodone
C4739195|T201|COMP|89989-8|LNC|Vilazodone|Vilazodone
C4739196|T201|COMP|89990-6|LNC|fluvoxaMINE|fluvoxaMINE
C4739197|T201|COMP|89991-4|LNC|Citalopram+Escitalopram|Citalopram+Escitalopram
C4739202|T201|COMP|90437-5|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4739204|T201|COMP|90438-3|LNC|Mycobacterium preliminary growth|Mycobacterium preliminary growth
C4739206|T201|COMP|90439-1|LNC|Atypical pneumonia pathogens panel|Atypical pneumonia pathogens panel
C4739208|T201|COMP|90440-9|LNC|BK virus+JC Virus DNA|BK virus+JC Virus DNA
C4739211|T201|COMP|90442-5|LNC|Coxiella burnetii aroE gene|Coxiella burnetii aroE gene
C4739229|T201|COMP|90924-2|LNC|BK virus DNA|BK virus DNA
C4739230|T201|COMP|90925-9|LNC|HBB gene full mutation analysis|HBB gene full mutation analysis
C4739231|T201|COMP|90926-7|LNC|MET gene amplification|MET gene amplification
C4739232|T201|COMP|90927-5|LNC|RET gene rearrangements|RET gene rearrangements
C4739233|T201|COMP|90975-4|LNC|Clomethiazole|Clomethiazole
C4739234|T201|COMP|90976-2|LNC|Opipramol|Opipramol
C4739235|T201|COMP|90977-0|LNC|Tianeptine|Tianeptine
C4739236|T201|COMP|90978-8|LNC|Vilazodone|Vilazodone
C4739237|T201|COMP|90979-6|LNC|Vortioxetine|Vortioxetine
C4739238|T201|COMP|90980-4|LNC|Meropenem+Vaborbactam|Meropenem+Vaborbactam
C4739248|T201|COMP|90425-0|LNC|Microorganism preliminary growth detection panel|Microorganism preliminary growth detection panel
C4739250|T201|COMP|90429-2|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4739251|T201|COMP|90430-0|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4739252|T201|COMP|90432-6|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4739253|T201|COMP|90433-4|LNC|Mycobacterium preliminary growth|Mycobacterium preliminary growth
C4739254|T201|COMP|90434-2|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4739255|T201|COMP|90435-9|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4739256|T201|COMP|90436-7|LNC|Microorganism preliminary growth|Microorganism preliminary growth
C4739277|T201|COMP|91133-9|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C4739286|T201|COMP|90227-0|LNC|Histoplasma capsulatum H & M Ab panel|Histoplasma capsulatum H & M Ab panel
C4739288|T201|COMP|90228-8|LNC|Extractable nuclear antigen Ab.IgG panel|Extractable nuclear antigen Ab.IgG panel
C4739290|T201|COMP|90229-6|LNC|Herpes simplex virus 1 & 2 Ab.IgG & IgM panel|Herpes simplex virus 1 & 2 Ab.IgG & IgM panel
C4739294|T201|COMP|90231-2|LNC|Thymoma & myasthenia gravis antibody panel|Thymoma & myasthenia gravis antibody panel
C4739296|T201|COMP|90232-0|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C4739299|T201|COMP|90250-2|LNC|Vanillylmandelate & Homovanillate panel|Vanillylmandelate & Homovanillate panel
C4739302|T201|COMP|90253-6|LNC|Measles virus Ab.IgG & IgM panel|Measles virus Ab.IgG & IgM panel
C4739303|T201|COMP|90254-4|LNC|Measles virus Ab.IgG & IgM panel|Measles virus Ab.IgG & IgM panel
C4739306|T201|COMP|90256-9|LNC|CFTR gene full mutation analysis|CFTR gene full mutation analysis
C4739308|T201|COMP|90258-5|LNC|LDLR gene full mutation analysis|LDLR gene full mutation analysis
C4739310|T201|COMP|90259-3|LNC|NAT2 gene full mutation analysis|NAT2 gene full mutation analysis
C4739312|T201|COMP|90260-1|LNC|Rickettsia spotted fever group Ab.IgG & IgM panel|Rickettsia spotted fever group Ab.IgG & IgM panel
C4739320|T201|COMP|90270-0|LNC|Bacteria identified|Bacteria identified
C4739321|T201|COMP|90271-8|LNC|Bacteria identified|Bacteria identified
C4739322|T201|COMP|90272-6|LNC|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C4739323|T201|COMP|90273-4|LNC|Bacteria identified|Bacteria identified
C4739324|T201|COMP|90274-2|LNC|Bacteria identified|Bacteria identified
C4739325|T201|COMP|90275-9|LNC|Gardnerella vaginalis|Gardnerella vaginalis
C4739326|T201|COMP|90276-7|LNC|Bacteria identified|Bacteria identified
C4739327|T201|COMP|90277-5|LNC|Bacteria identified|Bacteria identified
C4739328|T201|COMP|90278-3|LNC|Bacteria identified|Bacteria identified
C4739329|T201|COMP|90279-1|LNC|Bacteria identified|Bacteria identified
C4739330|T201|COMP|90280-9|LNC|Bacteria identified|Bacteria identified
C4739331|T201|COMP|90281-7|LNC|Bacteria identified|Bacteria identified
C4739333|T201|COMP|90283-3|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C4739334|T201|COMP|90284-1|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C4739335|T201|COMP|90285-8|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C4739336|T201|COMP|90286-6|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C4739337|T201|COMP|90287-4|LNC|Norovirus RNA|Norovirus RNA
C4739338|T201|COMP|90288-2|LNC|Norovirus Genogroup I RNA|Norovirus Genogroup I RNA
C4739339|T201|COMP|90289-0|LNC|Norovirus Genogroup II RNA|Norovirus Genogroup II RNA
C4739340|T201|COMP|90290-8|LNC|Alpha-1-Fetoprotein Ab|Alpha-1-Fetoprotein Ab
C4739342|T201|COMP|90291-6|LNC|Epithelial cell adhesion molecule Ab|Epithelial cell adhesion molecule Ab
C4739344|T201|COMP|90292-4|LNC|Liver cancer antibodies & Alpha-1-Fetoprotein|Liver cancer antibodies & Alpha-1-Fetoprotein
C4739348|T201|COMP|90294-0|LNC|Matrix metalloproteinases-9 Ab|Matrix metalloproteinases-9 Ab
C4739350|T201|COMP|90295-7|LNC|RalA Ab|RalA Ab
C4739353|T201|COMP|90297-3|LNC|Entamoeba histolytica Ab|Entamoeba histolytica Ab
C4739354|T201|COMP|90298-1|LNC|Entamoeba sp DNA|Entamoeba sp DNA
C4739355|T201|COMP|90299-9|LNC|Giardia sp DNA|Giardia sp DNA
C4739357|T201|COMP|90300-5|LNC|Helminth identified|Helminth identified
C4739358|T201|COMP|90301-3|LNC|Toxoplasma gondii|Toxoplasma gondii
C4739359|T201|COMP|90302-1|LNC|Trichomonas vaginalis DNA|Trichomonas vaginalis DNA
C4739360|T201|COMP|90303-9|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C4739361|T201|COMP|90903-6|LNC|HIV 1 RNA integrase gene|HIV 1 RNA integrase gene
C4739362|T201|COMP|90904-4|LNC|HIV 1 RNA protease gene|HIV 1 RNA protease gene
C4739363|T201|COMP|90905-1|LNC|ABO & Rh group|ABO & Rh group
C4739364|T201|COMP|90906-9|LNC|ABO & Rh group|ABO & Rh group
C4739371|T201|COMP|90304-7|LNC|Cells.CD3/100 lymphocytes|Cells.CD3/100 lymphocytes
C4739373|T201|COMP|89994-8|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C4739374|T201|COMP|89995-5|LNC|Trypanosoma cruzi Ab.IgG|Trypanosoma cruzi Ab.IgG
C4739375|T201|COMP|89996-3|LNC|Pneumocystis jiroveci DNA|Pneumocystis jiroveci DNA
C4739376|T201|COMP|89997-1|LNC|SUMF1 gene full mutation analysis|SUMF1 gene full mutation analysis
C4739378|T201|COMP|89998-9|LNC|Albumin/Creatinine|Albumin/Creatinine
C4739379|T201|COMP|89999-7|LNC|Albumin|Albumin
C4739380|T201|COMP|90000-1|LNC|Albumin|Albumin
C4739381|T201|COMP|90001-9|LNC|Staphylococcus aureus.methicillin resistant DNA|Staphylococcus aureus.methicillin resistant DNA
C4739382|T201|COMP|89871-8|LNC|Bilirubin|Bilirubin
C4739383|T201|COMP|89872-6|LNC|Bilirubin|Bilirubin
C4739386|T201|COMP|89645-6|LNC|Bartonella henselae DNA|Bartonella henselae DNA
C4739387|T201|COMP|89646-4|LNC|Bartonella quintana DNA|Bartonella quintana DNA
C4739388|T201|COMP|89647-2|LNC|Bartonella sp DNA|Bartonella sp DNA
C4739389|T201|COMP|89649-8|LNC|Coxiella burnetii DNA|Coxiella burnetii DNA
C4739390|T201|COMP|89650-6|LNC|Tropheryma whippelii DNA|Tropheryma whippelii DNA
C4739391|T201|COMP|89651-4|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C4739392|T201|COMP|89652-2|LNC|Human metapneumovirus Identified|Human metapneumovirus Identified
C4739463|T201|COMP|90804-6|LNC|Levothyroxine absorption|Levothyroxine absorption
C4739465|T201|COMP|90805-3|LNC|Vedolizumab^trough|Vedolizumab^trough
C4739468|T201|COMP|90885-5|LNC|Influenza virus D RNA|Influenza virus D RNA
C4739481|T201|COMP|90815-2|LNC|Amphiphysin Ab|Amphiphysin Ab
C4739482|T201|COMP|90816-0|LNC|Amphiphysin Ab|Amphiphysin Ab
C4739483|T201|COMP|90821-0|LNC|Contactin-associated protein 2 Ab|Contactin-associated protein 2 Ab
C4739491|T201|COMP|90824-4|LNC|Dipeptidyl aminopeptidase-like protein 6 Ab|Dipeptidyl aminopeptidase-like protein 6 Ab
C4739492|T201|COMP|90825-1|LNC|Gamma aminobutyrate B receptor Ab|Gamma aminobutyrate B receptor Ab
C4739493|T201|COMP|90826-9|LNC|Gamma aminobutyrate B receptor Ab|Gamma aminobutyrate B receptor Ab
C4739494|T201|COMP|90827-7|LNC|Glial nuclear type 1 Ab|Glial nuclear type 1 Ab
C4739499|T201|COMP|90841-8|LNC|Purkinje cell cytoplasmic type 1 Ab|Purkinje cell cytoplasmic type 1 Ab
C4739500|T201|COMP|90842-6|LNC|Purkinje cell cytoplasmic type 1 Ab|Purkinje cell cytoplasmic type 1 Ab
C4739501|T201|COMP|90843-4|LNC|Purkinje cell cytoplasmic type 2 Ab|Purkinje cell cytoplasmic type 2 Ab
C4739502|T201|COMP|90844-2|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C4739503|T201|COMP|91001-8|LNC|Myelin associated glycoprotein Ab.IgM|Myelin associated glycoprotein Ab.IgM
C4739514|T201|COMP|90799-8|LNC|Thyroxine^4H post dose levothyroxine|Thyroxine^4H post dose levothyroxine
C4739515|T201|COMP|90800-4|LNC|Thyroxine^6H post dose levothyroxine|Thyroxine^6H post dose levothyroxine
C4739522|T201|COMP|90448-2|LNC|Coccidioides sp Ab.IgM|Coccidioides sp Ab.IgM
C4739523|T201|COMP|90449-0|LNC|Norovirus genogroup I & II RNA|Norovirus genogroup I & II RNA
C4739553|T201|COMP|90801-2|LNC|Thyrotropin^6H post dose levothyroxine|Thyrotropin^6H post dose levothyroxine
C4739615|T201|COMP|90233-8|LNC|Dermatan sulfate|Dermatan sulfate
C4739632|T201|COMP|90320-3|LNC|Aichivirus C RNA|Aichivirus C RNA
C4739634|T201|COMP|90239-5|LNC|Suppression of tumorigenicity 2.soluble|Suppression of tumorigenicity 2.soluble
C4739636|T201|COMP|90240-3|LNC|Eculizumab|Eculizumab
C4739655|T201|COMP|90329-4|LNC|Porcine deltacoronavirus Ab.IgG/Positive control|Porcine deltacoronavirus Ab.IgG/Positive control
C4739657|T201|COMP|90330-2|LNC|Porcine parainfluenza virus 1 RNA|Porcine parainfluenza virus 1 RNA
C4739664|T201|COMP|90305-4|LNC|t(2;5)(p23;q35.1)(ALK,NPM1) fusion transcript|t(2;5)(p23;q35.1)(ALK,NPM1) fusion transcript
C4739665|T201|COMP|90306-2|LNC|Mycobacterium sp identified|Mycobacterium sp identified
C4739686|T201|COMP|90248-6|LNC|Myelin oligodendrocyte glycoprotein Ab.IgG1|Myelin oligodendrocyte glycoprotein Ab.IgG1
C4739701|T201|COMP|90234-6|LNC|Globotriaosylsphingosine|Globotriaosylsphingosine
C4739703|T201|COMP|90235-3|LNC|Heparan sulfate|Heparan sulfate
C4739707|T201|COMP|90325-2|LNC|Mycoplasma suis DNA|Mycoplasma suis DNA
C4739709|T201|COMP|90326-0|LNC|Porcine circovirus type 2d DNA|Porcine circovirus type 2d DNA
C4739756|T201|COMP|90339-3|LNC|Aspergillus sp DNA|Aspergillus sp DNA
C4739757|T201|COMP|90340-1|LNC|Aspergillus sp DNA|Aspergillus sp DNA
C4739766|T201|COMP|90362-5|LNC|Chlamydia trachomatis L1 Ab.IgG|Chlamydia trachomatis L1 Ab.IgG
C4739768|T201|COMP|90363-3|LNC|Chlamydia trachomatis L1 Ab.IgM|Chlamydia trachomatis L1 Ab.IgM
C4739770|T201|COMP|90364-1|LNC|Cholesterol.in LDL.small dense|Cholesterol.in LDL.small dense
C4739819|T201|COMP|90337-7|LNC|Cryptococcus sp rRNA gene|Cryptococcus sp rRNA gene
C4739820|T201|COMP|90338-5|LNC|Cryptococcus sp rRNA gene|Cryptococcus sp rRNA gene
C4739828|T201|COMP|90321-1|LNC|Aichivirus C RNA|Aichivirus C RNA
C4739829|T201|COMP|90322-9|LNC|Haemophilus parasuis serotype|Haemophilus parasuis serotype
C4739831|T201|COMP|90416-9|LNC|Lymphocyte subset & B-cell phenotyping panel|Lymphocyte subset & B-cell phenotyping panel
C4739835|T201|COMP|90418-5|LNC|BAFF-R Cells/100 cells.CD19|BAFF-R Cells/100 cells.CD19
C4739837|T201|COMP|90419-3|LNC|Apolipoprotein CIII-0/Apolipoprotein CIII-2|Apolipoprotein CIII-0/Apolipoprotein CIII-2
C4739841|T201|COMP|90421-9|LNC|Apolipoprotein CIII-1/Apolipoprotein CIII-2|Apolipoprotein CIII-1/Apolipoprotein CIII-2
C4739843|T201|COMP|90422-7|LNC|Cells.TACI/100 cells.CD19|Cells.TACI/100 cells.CD19
C4739872|T201|COMP|91121-4|LNC|Maltose binding protein Ab.IgE.RAST class|Maltose binding protein Ab.IgE.RAST class
C4739874|T201|COMP|91122-2|LNC|Maltose binding protein Ab.IgE|Maltose binding protein Ab.IgE
C4739884|T201|COMP|90443-3|LNC|Coxiella burnetii aroE gene|Coxiella burnetii aroE gene
C4739907|T201|COMP|90444-1|LNC|Diethylpropion|Diethylpropion
C4739908|T201|COMP|90445-8|LNC|ePHEDrine|ePHEDrine
C4739909|T201|COMP|90446-6|LNC|Pseudoephedrine|Pseudoephedrine
C4739910|T201|COMP|90447-4|LNC|Delafloxacin|Delafloxacin
C4739915|T201|COMP|90413-6|LNC|T-cell regulatory subsets panel|T-cell regulatory subsets panel
C4739917|T201|COMP|90414-4|LNC|B-cell phenotyping panel|B-cell phenotyping panel
C4739919|T201|COMP|90415-1|LNC|B-cell TACI & BAFF-R subsets panel|B-cell TACI & BAFF-R subsets panel
C4739921|T201|COMP|90423-5|LNC|Microorganism preliminary growth detection panel|Microorganism preliminary growth detection panel
C4739922|T201|COMP|90424-3|LNC|Microorganism preliminary growth detection panel|Microorganism preliminary growth detection panel
C4739937|T201|COMP|90845-9|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C4739938|T201|COMP|90846-7|LNC|Purkinje cell cytoplasmic type Tr Ab|Purkinje cell cytoplasmic type Tr Ab
C4739939|T201|COMP|90847-5|LNC|Zinc finger protein of the cerebellum 4 Ab|Zinc finger protein of the cerebellum 4 Ab
C4739941|T201|COMP|90849-1|LNC|Cefpodoxime 4.0 ug/mL|Cefpodoxime 4.0 ug/mL
C4739944|T201|COMP|90990-3|LNC|Protein.monoclonal isotype|Protein.monoclonal isotype
C4739948|T201|COMP|90450-8|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C4739949|T201|COMP|90451-6|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C4739950|T201|COMP|90837-6|LNC|Neuronal nuclear type 3 Ab|Neuronal nuclear type 3 Ab
C4739951|T201|COMP|90838-4|LNC|Neuronal nuclear type 3 Ab|Neuronal nuclear type 3 Ab
C4739952|T201|COMP|90839-2|LNC|N-methyl-D-aspartate receptor subunit 1 Ab|N-methyl-D-aspartate receptor subunit 1 Ab
C4739953|T201|COMP|90840-0|LNC|N-methyl-D-aspartate receptor subunit 1 Ab|N-methyl-D-aspartate receptor subunit 1 Ab
C4739954|T201|COMP|90817-8|LNC|Aquaporin 4 water channel Ab|Aquaporin 4 water channel Ab
C4739955|T201|COMP|90818-6|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C4739956|T201|COMP|90819-4|LNC|Aquaporin 4 water channel Ab.IgG|Aquaporin 4 water channel Ab.IgG
C4739957|T201|COMP|90820-2|LNC|Contactin-associated protein 2 Ab|Contactin-associated protein 2 Ab
C4739960|T201|COMP|90808-7|LNC|Candida krusei DNA|Candida krusei DNA
C4739961|T201|COMP|90809-5|LNC|Candida parapsilosis DNA|Candida parapsilosis DNA
C4739962|T201|COMP|90810-3|LNC|Candida tropicalis DNA|Candida tropicalis DNA
C4739964|T201|COMP|90806-1|LNC|Candida albicans DNA|Candida albicans DNA
C4739965|T201|COMP|90807-9|LNC|Candida glabrata DNA|Candida glabrata DNA
C4740006|T201|COMP|91139-6|LNC|Thiopurine methyltransferase activity panel|Thiopurine methyltransferase activity panel
C4740008|T201|COMP|91140-4|LNC|Brucella sp Ab.IgG & IgM panel|Brucella sp Ab.IgG & IgM panel
C4740009|T201|COMP|91141-2|LNC|Thiopurine methyltransferase|Thiopurine methyltransferase
C4740010|T201|COMP|91142-0|LNC|Thiopurine methyltransferase|Thiopurine methyltransferase
C4740011|T201|COMP|91143-8|LNC|Thiopurine methyltransferase|Thiopurine methyltransferase
C4740020|T201|COMP|91027-3|LNC|Buprenorphine-3-glucuronide|Buprenorphine-3-glucuronide
C4740021|T201|COMP|91028-1|LNC|Barbiturates|Barbiturates
C4740022|T201|COMP|91029-9|LNC|Cocaine+Benzoylecgonine|Cocaine+Benzoylecgonine
C4740023|T201|COMP|91030-7|LNC|Methadone+Metabolite|Methadone+Metabolite
C4740024|T201|COMP|91031-5|LNC|Methamphetamine+Methylenedioxymethamphetamine|Methamphetamine+Methylenedioxymethamphetamine
C4740026|T201|COMP|91032-3|LNC|oxyCODONE+Oxymorphone|oxyCODONE+Oxymorphone
C4740027|T201|COMP|91033-1|LNC|Methadone+Metabolite|Methadone+Metabolite
C4740028|T201|COMP|91034-9|LNC|Methamphetamine+Methylenedioxymethamphetamine|Methamphetamine+Methylenedioxymethamphetamine
C4740029|T201|COMP|91035-6|LNC|Phencyclidine|Phencyclidine
C4740030|T201|COMP|91036-4|LNC|Benzodiazepines|Benzodiazepines
C4740031|T201|COMP|91037-2|LNC|Methamphetamine+Methylenedioxymethamphetamine|Methamphetamine+Methylenedioxymethamphetamine
C4740032|T201|COMP|91038-0|LNC|Cocaine+Benzoylecgonine|Cocaine+Benzoylecgonine
C4740033|T201|COMP|91039-8|LNC|Methadone+Metabolite|Methadone+Metabolite
C4740034|T201|COMP|91040-6|LNC|Phencyclidine|Phencyclidine
C4740035|T201|COMP|91041-4|LNC|Cannabinoids|Cannabinoids
C4740036|T201|COMP|91042-2|LNC|Methamphetamine+Methylenedioxymethamphetamine|Methamphetamine+Methylenedioxymethamphetamine
C4740037|T201|COMP|91043-0|LNC|Opiates|Opiates
C4740038|T201|COMP|91044-8|LNC|oxyCODONE+Oxymorphone|oxyCODONE+Oxymorphone
C4740039|T201|COMP|91045-5|LNC|Methamphetamine+Methylenedioxymethamphetamine|Methamphetamine+Methylenedioxymethamphetamine
C4740040|T201|COMP|91046-3|LNC|Methadone+Metabolite|Methadone+Metabolite
C4740041|T201|COMP|91047-1|LNC|Barbiturates|Barbiturates
C4740042|T201|COMP|91048-9|LNC|Cannabinoids|Cannabinoids
C4740043|T201|COMP|91049-7|LNC|Cocaine+Benzoylecgonine|Cocaine+Benzoylecgonine
C4740044|T201|COMP|91050-5|LNC|Methadone+Metabolite|Methadone+Metabolite
C4740045|T201|COMP|91051-3|LNC|Methamphetamine+Methylenedioxymethamphetamine|Methamphetamine+Methylenedioxymethamphetamine
C4740046|T201|COMP|91052-1|LNC|Opiates|Opiates
C4740047|T201|COMP|91053-9|LNC|oxyCODONE+Oxymorphone|oxyCODONE+Oxymorphone
C4740048|T201|COMP|91054-7|LNC|Drugs of abuse panel|Drugs of abuse panel
C4740049|T201|COMP|91055-4|LNC|Drugs of abuse panel|Drugs of abuse panel
C4740050|T201|COMP|91056-2|LNC|Drugs of abuse panel|Drugs of abuse panel
C4740051|T201|COMP|91057-0|LNC|Tropheryma whippelii DNA|Tropheryma whippelii DNA
C4740052|T201|COMP|91058-8|LNC|Kingella kingae DNA|Kingella kingae DNA
C4740053|T201|COMP|91059-6|LNC|Kingella kingae DNA|Kingella kingae DNA
C4740054|T201|COMP|91060-4|LNC|Helicobacter pylori DNA|Helicobacter pylori DNA
C4740055|T201|COMP|91061-2|LNC|Helicobacter pylori DNA|Helicobacter pylori DNA
C4740056|T201|COMP|91062-0|LNC|Bacteria identified|Bacteria identified
C4740057|T201|COMP|91063-8|LNC|Bacteria identified|Bacteria identified
C4740058|T201|COMP|91064-6|LNC|Dengue virus NS1 Ag|Dengue virus NS1 Ag
C4740059|T201|COMP|91065-3|LNC|14-3-3 protein|14-3-3 protein
C4740060|T201|COMP|91066-1|LNC|Enterovirus RNA|Enterovirus RNA
C4740061|T201|COMP|91067-9|LNC|Enterovirus RNA|Enterovirus RNA
C4740062|T201|COMP|91068-7|LNC|Enterovirus RNA|Enterovirus RNA
C4740063|T201|COMP|91069-5|LNC|Enterovirus RNA|Enterovirus RNA
C4740064|T201|COMP|91070-3|LNC|Hepatitis A virus RNA|Hepatitis A virus RNA
C4740065|T201|COMP|91071-1|LNC|Hepatitis E virus RNA|Hepatitis E virus RNA
C4740066|T201|COMP|91072-9|LNC|Influenza virus A subtype|Influenza virus A subtype
C4740067|T201|COMP|91073-7|LNC|Human papilloma virus genotype|Human papilloma virus genotype
C4740068|T201|COMP|91074-5|LNC|Phlebovirus sp RNA|Phlebovirus sp RNA
C4740070|T201|COMP|91075-2|LNC|Rabies virus Ag|Rabies virus Ag
C4740071|T201|COMP|91076-0|LNC|Rabies virus Ag|Rabies virus Ag
C4740072|T201|COMP|91077-8|LNC|Measles virus RNA|Measles virus RNA
C4740073|T201|COMP|91078-6|LNC|Zika virus RNA|Zika virus RNA
C4740074|T201|COMP|91079-4|LNC|Zika virus RNA|Zika virus RNA
C4740075|T201|COMP|91080-2|LNC|Zika virus Ab.IgG|Zika virus Ab.IgG
C4740076|T201|COMP|91081-0|LNC|Candida sp DNA|Candida sp DNA
C4740077|T201|COMP|91082-8|LNC|Fungal 18S rRNA gene|Fungal 18S rRNA gene
C4740079|T201|COMP|91083-6|LNC|Fungal 18S rRNA gene|Fungal 18S rRNA gene
C4740080|T201|COMP|91084-4|LNC|Fungal 18S rRNA gene|Fungal 18S rRNA gene
C4740081|T201|COMP|91085-1|LNC|Fungal 18S rRNA gene|Fungal 18S rRNA gene
C4740082|T201|COMP|91086-9|LNC|Fungal BT2 gene|Fungal BT2 gene
C4740084|T201|COMP|91087-7|LNC|Fungal BT2 gene|Fungal BT2 gene
C4740085|T201|COMP|91088-5|LNC|Fungal BT2 gene|Fungal BT2 gene
C4740086|T201|COMP|91089-3|LNC|Fungal BT2 gene|Fungal BT2 gene
C4740087|T201|COMP|91090-1|LNC|Fungal ITS region|Fungal ITS region
C4740089|T201|COMP|91091-9|LNC|Fungal ITS region|Fungal ITS region
C4740090|T201|COMP|91092-7|LNC|Fungal ITS region|Fungal ITS region
C4740091|T201|COMP|91093-5|LNC|Fungal ITS region|Fungal ITS region
C4740152|T201|COMP|90465-6|LNC|3-(4-fluorobenzoyl)propionate|3-(4-fluorobenzoyl)propionate
C4740154|T201|COMP|90466-4|LNC|3-(4-fluorobenzoyl)propionate|3-(4-fluorobenzoyl)propionate
C4740155|T201|COMP|90467-2|LNC|Hydroxyaripiprazole|Hydroxyaripiprazole
C4740157|T201|COMP|90468-0|LNC|Hydroxyaripiprazole|Hydroxyaripiprazole
C4740158|T201|COMP|90469-8|LNC|Norfluvoxamine|Norfluvoxamine
C4740160|T201|COMP|90470-6|LNC|Norfluvoxamine|Norfluvoxamine
C4740161|T201|COMP|90471-4|LNC|9-Hydroxyrisperidone|9-Hydroxyrisperidone
C4740162|T201|COMP|90780-8|LNC|inFLIXimab Ab|inFLIXimab Ab
C4740163|T201|COMP|90781-6|LNC|N,N'-Dimethylarginine|N,N'-Dimethylarginine
C4740164|T201|COMP|90782-4|LNC|F2-Isoprostanes|F2-Isoprostanes
C4740165|T201|COMP|90783-2|LNC|F2-Isoprostanes/Creatinine|F2-Isoprostanes/Creatinine
C4740167|T201|COMP|90794-9|LNC|Vedolizumab & Vedolizumab Ab Panel|Vedolizumab & Vedolizumab Ab Panel
C4740169|T201|COMP|90795-6|LNC|Levothyroxine absorption panel|Levothyroxine absorption panel
C4740171|T201|COMP|90796-4|LNC|Thyroxine^1H post dose levothyroxine|Thyroxine^1H post dose levothyroxine
C4740172|T201|COMP|90750-1|LNC|O-Nortramadol|O-Nortramadol
C4740173|T201|COMP|90746-9|LNC|5-fluoro ADB-M7|5-fluoro ADB-M7
C4740175|T201|COMP|90747-7|LNC|MDMB-FUBINACA-M1|MDMB-FUBINACA-M1
C4740177|T201|COMP|90748-5|LNC|Atomoxetine|Atomoxetine
C4759679|T201|COMP|35188-2|LNC|Aldosterone^upright|Aldosterone^upright
C4759680|T201|COMP|35190-8|LNC|Androstenedione|Androstenedione
C4759916|T201|COMP|92551-1|LNC|C Ag inferred phenotype|C Ag inferred phenotype
C4759948|T201|COMP|92496-9|LNC|K Ag inferred phenotype|K Ag inferred phenotype
C4759949|T201|COMP|92489-4|LNC|little k Ag inferred phenotype|little k Ag inferred phenotype
C4759950|T201|COMP|92534-7|LNC|K Ag inferred phenotype|K Ag inferred phenotype
C4759951|T201|COMP|92527-1|LNC|little k Ag inferred phenotype|little k Ag inferred phenotype
C4760186|T201|COMP|92506-5|LNC|E Ag inferred phenotype|E Ag inferred phenotype
C4760187|T201|COMP|92490-2|LNC|little e Ag inferred phenotype|little e Ag inferred phenotype
C4760188|T201|COMP|92544-6|LNC|E Ag inferred phenotype|E Ag inferred phenotype
C4760189|T201|COMP|92528-9|LNC|little e Ag inferred phenotype|little e Ag inferred phenotype
C4760229|T201|COMP|92236-9|LNC|Lab observation result status|Lab observation result status
C4760232|T201|COMP|92237-7|LNC|Lab observation sub-type|Lab observation sub-type
C4760233|T201|COMP|92235-1|LNC|Lab order result status|Lab order result status
C4760235|T201|COMP|91672-6|LNC|ABCB1 gene targeted mutation analysis|ABCB1 gene targeted mutation analysis
C4760253|T201|COMP|92483-7|LNC|S Ag inferred phenotype|S Ag inferred phenotype
C4760254|T201|COMP|92488-6|LNC|little s Ag inferred phenotype|little s Ag inferred phenotype
C4760255|T201|COMP|92521-4|LNC|S Ag inferred phenotype|S Ag inferred phenotype
C4760256|T201|COMP|92526-3|LNC|little s Ag inferred phenotype|little s Ag inferred phenotype
C4760312|T201|COMP|93044-6|LNC|Level of evidence|Level of evidence
C4760456|T201|COMP|92491-0|LNC|little c Ag inferred phenotype|little c Ag inferred phenotype
C4760457|T201|COMP|92513-1|LNC|C Ag inferred phenotype|C Ag inferred phenotype
C4760458|T201|COMP|92529-7|LNC|little c Ag inferred phenotype|little c Ag inferred phenotype
C4760461|T201|COMP|92824-2|LNC|Source of population allelic frequency data|Source of population allelic frequency data
C4760462|T201|COMP|93047-9|LNC|Specimen condition|Specimen condition
C4760533|T201|COMP|92005-8|LNC|Spinal muscular atrophy newborn screening panel|Spinal muscular atrophy newborn screening panel
C5143163|T201|COMP|87925-4|LNC|Reagin Ab|Reagin Ab
C5143203|T201|COMP|90066-2|LNC|Corynebacterium sp identified|Corynebacterium sp identified
C5143204|T201|COMP|90067-0|LNC|Enterobacteriaceae identified|Enterobacteriaceae identified
C5143205|T201|COMP|90068-8|LNC|Gram negative bacilli identified|Gram negative bacilli identified
C5143206|T201|COMP|90069-6|LNC|Gram positive bacilli identified|Gram positive bacilli identified
C5143207|T201|COMP|90070-4|LNC|Gram positive catalase producing cocci identified|Gram positive catalase producing cocci identified
C5143209|T201|COMP|90072-0|LNC|Haemophilus sp & Neisseria sp identified|Haemophilus sp & Neisseria sp identified
C5143210|T201|COMP|90073-8|LNC|Lactobacillales identified|Lactobacillales identified
C5143211|T201|COMP|90075-3|LNC|Non-Enterobacteriaceae identified|Non-Enterobacteriaceae identified
C5143212|T201|COMP|90076-1|LNC|Staphylococcus sp identified|Staphylococcus sp identified
C5143213|T201|COMP|90077-9|LNC|Urinary pathogens identified|Urinary pathogens identified
C5143214|T201|COMP|90078-7|LNC|Yeast identified|Yeast identified
C5143215|T201|COMP|90100-9|LNC|Listeria sp identified|Listeria sp identified
C5143645|T201|COMP|91542-1|LNC|Myelin oligodendrocyte glycoprotein Ab|Myelin oligodendrocyte glycoprotein Ab
C5143646|T201|COMP|91543-9|LNC|Myelin oligodendrocyte glycoprotein Ab|Myelin oligodendrocyte glycoprotein Ab
C5143647|T201|COMP|91544-7|LNC|Myelin oligodendrocyte glycoprotein Ab|Myelin oligodendrocyte glycoprotein Ab
C5143648|T201|COMP|91545-4|LNC|Myelin oligodendrocyte glycoprotein Ab|Myelin oligodendrocyte glycoprotein Ab
C5143650|T201|COMP|91551-2|LNC|Other cells/100 leukocytes|Other cells/100 leukocytes
C5143655|T201|COMP|91556-1|LNC|Fibrin D-dimer DDU|Fibrin D-dimer DDU
C5143674|T201|COMP|91586-8|LNC|Coding system|Coding system
C5143677|T201|COMP|91590-0|LNC|Mycobacterium preliminary growth|Mycobacterium preliminary growth
C5143690|T201|COMP|91606-4|LNC|Clomipramine+Norclomipramine|Clomipramine+Norclomipramine
C5143744|T201|COMP|91664-3|LNC|Ambrosia deltoidea Ab.IgE|Ambrosia deltoidea Ab.IgE
C5143745|T201|COMP|91665-0|LNC|Ascorbate oxidase Ab.IgE|Ascorbate oxidase Ab.IgE
C5143746|T201|COMP|91666-8|LNC|Ascorbate oxidase Ab.IgE.RAST class|Ascorbate oxidase Ab.IgE.RAST class
C5143747|T201|COMP|91667-6|LNC|Aspergillus clavatus Ab|Aspergillus clavatus Ab
C5143748|T201|COMP|91668-4|LNC|Aspergillus oryzae Ab|Aspergillus oryzae Ab
C5143749|T201|COMP|91669-2|LNC|CYP3A7 gene targeted mutation analysis|CYP3A7 gene targeted mutation analysis
C5143750|T201|COMP|91670-0|LNC|Orexin-A|Orexin-A
C5143752|T201|COMP|91673-4|LNC|Cells.CD3+CD16+CD56+/100 cells|Cells.CD3+CD16+CD56+/100 cells
C5143753|T201|COMP|91674-2|LNC|Cells.CD3+CD16+CD56+|Cells.CD3+CD16+CD56+
C5143754|T201|COMP|91675-9|LNC|Giardia lamblia & Cryptosporidium parvum Ag panel|Giardia lamblia & Cryptosporidium parvum Ag panel
C5143755|T201|COMP|91676-7|LNC|Giardia lamblia Ag|Giardia lamblia Ag
C5143756|T201|COMP|91677-5|LNC|Cryptosporidium parvum Ag|Cryptosporidium parvum Ag
C5143757|T201|COMP|91678-3|LNC|Zika virus Ab.IgM|Zika virus Ab.IgM
C5143761|T201|COMP|91682-5|LNC|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C5143763|T201|COMP|91684-1|LNC|Histoplasma capsulatum H & M Ab panel|Histoplasma capsulatum H & M Ab panel
C5143764|T201|COMP|91685-8|LNC|Glutathione|Glutathione
C5143782|T201|COMP|91705-4|LNC|Corticotropin^5M pre 1 ug/kg CRH IV|Corticotropin^5M pre 1 ug/kg CRH IV
C5143783|T201|COMP|91706-2|LNC|Corticotropin^1M pre 1 ug/kg CRH IV|Corticotropin^1M pre 1 ug/kg CRH IV
C5143785|T201|COMP|91708-8|LNC|Corticotropin^10M post 1 ug/kg CRH IV|Corticotropin^10M post 1 ug/kg CRH IV
C5143786|T201|COMP|91709-6|LNC|Corticotropin^2M post 1 ug/kg CRH IV|Corticotropin^2M post 1 ug/kg CRH IV
C5143787|T201|COMP|91712-0|LNC|F5 gene.c.1691G>A|F5 gene.c.1691G>A
C5143832|T201|COMP|91761-7|LNC|Giardia sp Ag|Giardia sp Ag
C5143833|T201|COMP|91763-3|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C5143834|T201|COMP|91764-1|LNC|Nocardia sp identified|Nocardia sp identified
C5143835|T201|COMP|91765-8|LNC|Entamoeba sp DNA|Entamoeba sp DNA
C5143836|T201|COMP|91766-6|LNC|Entamoeba histolytica DNA|Entamoeba histolytica DNA
C5143837|T201|COMP|91767-4|LNC|Giardia sp DNA|Giardia sp DNA
C5143838|T201|COMP|91768-2|LNC|Ova & parasites identified|Ova & parasites identified
C5143839|T201|COMP|91769-0|LNC|Enterovirus RNA|Enterovirus RNA
C5143840|T201|COMP|91770-8|LNC|Enterovirus identified|Enterovirus identified
C5143841|T201|COMP|91771-6|LNC|Influenza virus A subtype|Influenza virus A subtype
C5143842|T201|COMP|91772-4|LNC|Influenza virus identified|Influenza virus identified
C5143843|T201|COMP|91773-2|LNC|Herpes simplex virus identified|Herpes simplex virus identified
C5143844|T201|COMP|91774-0|LNC|Varicella zoster virus Ag|Varicella zoster virus Ag
C5143845|T201|COMP|91775-7|LNC|Bordetella sp identified|Bordetella sp identified
C5143846|T201|COMP|91776-5|LNC|Mycoplasma sp.respiratory identified|Mycoplasma sp.respiratory identified
C5143847|T201|COMP|91777-3|LNC|Bordetella sp identified|Bordetella sp identified
C5143848|T201|COMP|91778-1|LNC|Human metapneumovirus identified|Human metapneumovirus identified
C5143849|T201|COMP|91779-9|LNC|Yeast identified|Yeast identified
C5143850|T201|COMP|91780-7|LNC|Measles virus|Measles virus
C5143851|T201|COMP|91781-5|LNC|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C5143852|T201|COMP|91782-3|LNC|Respiratory syncytial virus identified|Respiratory syncytial virus identified
C5143853|T201|COMP|91783-1|LNC|Cytomegalovirus|Cytomegalovirus
C5143854|T201|COMP|91784-9|LNC|Varicella zoster virus|Varicella zoster virus
C5143855|T201|COMP|91785-6|LNC|Respiratory syncytial virus identified|Respiratory syncytial virus identified
C5143856|T201|COMP|91786-4|LNC|Measles virus|Measles virus
C5143857|T201|COMP|91787-2|LNC|Mumps virus|Mumps virus
C5143858|T201|COMP|91788-0|LNC|Neisseria meningitidis|Neisseria meningitidis
C5143859|T201|COMP|91789-8|LNC|Haemophilus ducreyi|Haemophilus ducreyi
C5143860|T201|COMP|91790-6|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C5143861|T201|COMP|91791-4|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C5143862|T201|COMP|91792-2|LNC|Rubella virus RNA|Rubella virus RNA
C5143863|T201|COMP|91793-0|LNC|Rhinovirus RNA|Rhinovirus RNA
C5143864|T201|COMP|91794-8|LNC|Respiratory syncytial virus B RNA|Respiratory syncytial virus B RNA
C5143865|T201|COMP|91795-5|LNC|Respiratory syncytial virus A RNA|Respiratory syncytial virus A RNA
C5143866|T201|COMP|91796-3|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C5143867|T201|COMP|91797-1|LNC|Parvovirus B19 DNA|Parvovirus B19 DNA
C5143868|T201|COMP|91798-9|LNC|Parainfluenza virus RNA|Parainfluenza virus RNA
C5143869|T201|COMP|91799-7|LNC|Parainfluenza virus 4 RNA|Parainfluenza virus 4 RNA
C5143870|T201|COMP|91800-3|LNC|Parainfluenza virus 3 RNA|Parainfluenza virus 3 RNA
C5143871|T201|COMP|91801-1|LNC|Parainfluenza virus 2 RNA|Parainfluenza virus 2 RNA
C5143872|T201|COMP|91802-9|LNC|Parainfluenza virus 1 RNA|Parainfluenza virus 1 RNA
C5143873|T201|COMP|91803-7|LNC|Neisseria meningitidis DNA|Neisseria meningitidis DNA
C5143874|T201|COMP|91804-5|LNC|Mycoplasma pneumoniae DNA|Mycoplasma pneumoniae DNA
C5143875|T201|COMP|91805-2|LNC|Mycobacterium leprae DNA|Mycobacterium leprae DNA
C5143876|T201|COMP|91806-0|LNC|Mumps virus RNA|Mumps virus RNA
C5143877|T201|COMP|91807-8|LNC|Middle east respiratory syndrome coronavirus RNA|Middle east respiratory syndrome coronavirus RNA
C5143879|T201|COMP|91809-4|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C5143880|T201|COMP|91810-2|LNC|Human metapneumovirus Ag|Human metapneumovirus Ag
C5143881|T201|COMP|91811-0|LNC|Human bocavirus Ag|Human bocavirus Ag
C5143882|T201|COMP|91812-8|LNC|Fungus identified|Fungus identified
C5143883|T201|COMP|91813-6|LNC|Bordetella sp DNA|Bordetella sp DNA
C5143884|T201|COMP|91814-4|LNC|Bordetella sp Ag|Bordetella sp Ag
C5143885|T201|COMP|91815-1|LNC|Bordetella pertussis DNA|Bordetella pertussis DNA
C5143886|T201|COMP|91816-9|LNC|Bordetella parapertussis DNA|Bordetella parapertussis DNA
C5143887|T201|COMP|91817-7|LNC|Bordetella holmesii DNA|Bordetella holmesii DNA
C5143888|T201|COMP|91818-5|LNC|Bacteria identified|Bacteria identified
C5143889|T201|COMP|91819-3|LNC|Bacteria identified|Bacteria identified
C5143890|T201|COMP|91820-1|LNC|Adenovirus DNA|Adenovirus DNA
C5143891|T201|COMP|91821-9|LNC|Adenovirus Ag|Adenovirus Ag
C5143892|T201|COMP|91822-7|LNC|Adenovirus Ag|Adenovirus Ag
C5143893|T201|COMP|91823-5|LNC|Rubella virus RNA|Rubella virus RNA
C5143894|T201|COMP|91824-3|LNC|Pneumocystis jiroveci Ag|Pneumocystis jiroveci Ag
C5143895|T201|COMP|91825-0|LNC|Parechovirus RNA|Parechovirus RNA
C5143896|T201|COMP|91826-8|LNC|Ova & parasites identified|Ova & parasites identified
C5143897|T201|COMP|91827-6|LNC|Mycoplasma hominis DNA|Mycoplasma hominis DNA
C5143898|T201|COMP|91828-4|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C5143899|T201|COMP|91829-2|LNC|Mycobacterium tuberculosis DNA|Mycobacterium tuberculosis DNA
C5143900|T201|COMP|91830-0|LNC|Middle east respiratory syndrome coronavirus RNA|Middle east respiratory syndrome coronavirus RNA
C5143901|T201|COMP|91831-8|LNC|Human metapneumovirus Ag|Human metapneumovirus Ag
C5143902|T201|COMP|91832-6|LNC|Human bocavirus Ag|Human bocavirus Ag
C5143903|T201|COMP|91833-4|LNC|Herpes simplex virus Ag|Herpes simplex virus Ag
C5143904|T201|COMP|91834-2|LNC|Herpes simplex virus 2 Ag|Herpes simplex virus 2 Ag
C5143905|T201|COMP|91835-9|LNC|Herpes simplex virus 1 Ag|Herpes simplex virus 1 Ag
C5143906|T201|COMP|91836-7|LNC|Giardia sp DNA|Giardia sp DNA
C5143907|T201|COMP|91837-5|LNC|Francisella sp DNA|Francisella sp DNA
C5143908|T201|COMP|91838-3|LNC|Bordetella sp DNA|Bordetella sp DNA
C5143909|T201|COMP|91839-1|LNC|Bordetella sp Ag|Bordetella sp Ag
C5143910|T201|COMP|91840-9|LNC|Bordetella holmesii DNA|Bordetella holmesii DNA
C5143911|T201|COMP|91841-7|LNC|Adenovirus Ag|Adenovirus Ag
C5143912|T201|COMP|91842-5|LNC|Ureaplasma urealyticum DNA|Ureaplasma urealyticum DNA
C5143913|T201|COMP|91843-3|LNC|Ureaplasma parvum DNA|Ureaplasma parvum DNA
C5143914|T201|COMP|91844-1|LNC|Trichomonas vaginalis DNA|Trichomonas vaginalis DNA
C5143915|T201|COMP|91845-8|LNC|Trichomonas vaginalis|Trichomonas vaginalis
C5143916|T201|COMP|91846-6|LNC|Treponema pallidum DNA|Treponema pallidum DNA
C5143917|T201|COMP|91847-4|LNC|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C5143918|T201|COMP|91848-2|LNC|Mycoplasma hominis DNA|Mycoplasma hominis DNA
C5143919|T201|COMP|91849-0|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C5143921|T201|COMP|91851-6|LNC|Human papilloma virus genotype|Human papilloma virus genotype
C5143922|T201|COMP|91852-4|LNC|Human papilloma virus DNA|Human papilloma virus DNA
C5143924|T201|COMP|91854-0|LNC|Human papilloma virus 18 DNA|Human papilloma virus 18 DNA
C5143926|T201|COMP|91856-5|LNC|Human papilloma virus 16 DNA|Human papilloma virus 16 DNA
C5143927|T201|COMP|91857-3|LNC|Herpes simplex virus DNA|Herpes simplex virus DNA
C5143928|T201|COMP|91858-1|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C5143929|T201|COMP|91859-9|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C5143930|T201|COMP|91860-7|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C5143931|T201|COMP|91861-5|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C5143932|T201|COMP|91862-3|LNC|Bartonella sp DNA|Bartonella sp DNA
C5143933|T201|COMP|91863-1|LNC|Bartonella quintana DNA|Bartonella quintana DNA
C5143934|T201|COMP|91864-9|LNC|Bartonella henselae DNA|Bartonella henselae DNA
C5143935|T201|COMP|91865-6|LNC|Bacteria identified|Bacteria identified
C5143936|T201|COMP|91866-4|LNC|Bacteria identified|Bacteria identified
C5143937|T201|COMP|91867-2|LNC|Bordetella holmesii DNA|Bordetella holmesii DNA
C5143938|T201|COMP|91868-0|LNC|Bordetella parapertussis DNA|Bordetella parapertussis DNA
C5143939|T201|COMP|91869-8|LNC|Bordetella pertussis DNA|Bordetella pertussis DNA
C5143940|T201|COMP|91870-6|LNC|Bordetella sp Ag|Bordetella sp Ag
C5143941|T201|COMP|91871-4|LNC|Bordetella sp DNA|Bordetella sp DNA
C5143942|T201|COMP|91872-2|LNC|Bordetella sp identified|Bordetella sp identified
C5143943|T201|COMP|91873-0|LNC|Chlamydia trachomatis Ag|Chlamydia trachomatis Ag
C5143944|T201|COMP|91874-8|LNC|Mycoplasma genitalium DNA|Mycoplasma genitalium DNA
C5143945|T201|COMP|91875-5|LNC|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C5143946|T201|COMP|91876-3|LNC|Brucella sp Ab|Brucella sp Ab
C5143953|T201|COMP|91895-3|LNC|Bacterial strain|Bacterial strain
C5143954|T201|COMP|91896-1|LNC|Mycoplasma pneumoniae Ab|Mycoplasma pneumoniae Ab
C5143955|T201|COMP|91897-9|LNC|Doravirine|Doravirine
C5143956|T201|COMP|91898-7|LNC|Epizootic hemorrhagic disease virus RNA|Epizootic hemorrhagic disease virus RNA
C5144051|T201|COMP|92002-5|LNC|SMN1 gene|SMN1 gene
C5144052|T201|COMP|92004-1|LNC|Spinal muscular atrophy|Spinal muscular atrophy
C5144053|T201|COMP|92006-6|LNC|T-cell receptor excision circle|T-cell receptor excision circle
C5144054|T201|COMP|92007-4|LNC|T-cell receptor excision circle|T-cell receptor excision circle
C5144055|T201|COMP|92008-2|LNC|T-cell receptor excision circle|T-cell receptor excision circle
C5144069|T201|COMP|92024-9|LNC|Plazomicin^trough|Plazomicin^trough
C5144154|T201|COMP|92125-4|LNC|Streptococcus pneumoniae DNA|Streptococcus pneumoniae DNA
C5144155|T201|COMP|92126-2|LNC|Mycoplasma pneumoniae DNA|Mycoplasma pneumoniae DNA
C5144156|T201|COMP|92127-0|LNC|Haemophilus influenzae DNA|Haemophilus influenzae DNA
C5144157|T201|COMP|92128-8|LNC|Bordetella pertussis DNA|Bordetella pertussis DNA
C5144158|T201|COMP|92129-6|LNC|Bordetella parapertussis DNA|Bordetella parapertussis DNA
C5144159|T201|COMP|92130-4|LNC|Rhinovirus RNA|Rhinovirus RNA
C5144160|T201|COMP|92131-2|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C5144161|T201|COMP|92132-0|LNC|Enterovirus A+B+C RNA|Enterovirus A+B+C RNA
C5144162|T201|COMP|92133-8|LNC|Chlamydophila pneumoniae DNA|Chlamydophila pneumoniae DNA
C5144163|T201|COMP|92134-6|LNC|Human metapneumovirus RNA|Human metapneumovirus RNA
C5144164|T201|COMP|92135-3|LNC|Human bocavirus 1+2+3 DNA|Human bocavirus 1+2+3 DNA
C5144165|T201|COMP|92136-1|LNC|Adenovirus B+C+E DNA|Adenovirus B+C+E DNA
C5144166|T201|COMP|92137-9|LNC|Parainfluenza virus 4 RNA|Parainfluenza virus 4 RNA
C5144167|T201|COMP|92138-7|LNC|Parainfluenza virus 3 RNA|Parainfluenza virus 3 RNA
C5144168|T201|COMP|92139-5|LNC|Parainfluenza virus 2 RNA|Parainfluenza virus 2 RNA
C5144169|T201|COMP|92140-3|LNC|Parainfluenza virus 1 RNA|Parainfluenza virus 1 RNA
C5144170|T201|COMP|92141-1|LNC|Influenza virus B RNA|Influenza virus B RNA
C5144171|T201|COMP|92142-9|LNC|Influenza virus A RNA|Influenza virus A RNA
C5144172|T201|COMP|92143-7|LNC|Respiratory pathogens DNA & RNA panel|Respiratory pathogens DNA & RNA panel
C5144173|T201|COMP|92144-5|LNC|Moraxella catarrhalis DNA|Moraxella catarrhalis DNA
C5144174|T201|COMP|92145-2|LNC|Legionella pneumophila DNA|Legionella pneumophila DNA
C5144175|T201|COMP|92146-0|LNC|Human coronavirus 229E+NL63 RNA|Human coronavirus 229E+NL63 RNA
C5144176|T201|COMP|92147-8|LNC|Human coronavirus HKU1+OC43 RNA|Human coronavirus HKU1+OC43 RNA
C5144250|T201|COMP|92241-9|LNC|Vancomycin|Vancomycin
C5144251|T201|COMP|92242-7|LNC|Pyrazinamide|Pyrazinamide
C5144252|T201|COMP|92243-5|LNC|Microorganism resistance mutation tested for|Microorganism resistance mutation tested for
C5144255|T201|COMP|92246-8|LNC|Microorganism resistance mutation detected|Microorganism resistance mutation detected
C5144258|T201|COMP|92249-2|LNC|Microorganism gene tested for|Microorganism gene tested for
C5144259|T201|COMP|92250-0|LNC|Microorganism gene target region|Microorganism gene target region
C5144260|T201|COMP|92251-8|LNC|Microorganism gene detected|Microorganism gene detected
C5144261|T201|COMP|92252-6|LNC|Microorganism molecular resistance panel|Microorganism molecular resistance panel
C5144262|T201|COMP|92253-4|LNC|Microorganism identified|Microorganism identified
C5144264|T201|COMP|92255-9|LNC|Methicillin|Methicillin
C5144462|T201|COMP|92478-7|LNC|VS Ag inferred phenotype|VS Ag inferred phenotype
C5144463|T201|COMP|92479-5|LNC|V Ag inferred phenotype|V Ag inferred phenotype
C5144464|T201|COMP|92480-3|LNC|U Ag inferred phenotype|U Ag inferred phenotype
C5144465|T201|COMP|92481-1|LNC|S little c super 2 Ag inferred phenotype|S little c super 2 Ag inferred phenotype
C5144466|T201|COMP|92482-9|LNC|S little c super 1 Ag inferred phenotype|S little c super 1 Ag inferred phenotype
C5144467|T201|COMP|92484-5|LNC|N Ag inferred phenotype|N Ag inferred phenotype
C5144468|T201|COMP|92485-2|LNC|M Ag inferred phenotype|M Ag inferred phenotype
C5144469|T201|COMP|92486-0|LNC|LW super little b Ag inferred phenotype|LW super little b Ag inferred phenotype
C5144470|T201|COMP|92487-8|LNC|LW super little a Ag inferred phenotype|LW super little a Ag inferred phenotype
C5144471|T201|COMP|92492-8|LNC|L little u super little b Ag inferred phenotype|L little u super little b Ag inferred phenotype
C5144472|T201|COMP|92493-6|LNC|L little u super little a Ag inferred phenotype|L little u super little a Ag inferred phenotype
C5144473|T201|COMP|92494-4|LNC|K little p super little b Ag inferred phenotype|K little p super little b Ag inferred phenotype
C5144474|T201|COMP|92495-1|LNC|K little p super little a Ag inferred phenotype|K little p super little a Ag inferred phenotype
C5144475|T201|COMP|92497-7|LNC|J little s super little b Ag inferred phenotype|J little s super little b Ag inferred phenotype
C5144476|T201|COMP|92498-5|LNC|J little s super little a Ag inferred phenotype|J little s super little a Ag inferred phenotype
C5144477|T201|COMP|92499-3|LNC|J little o super little a Ag inferred phenotype|J little o super little a Ag inferred phenotype
C5144478|T201|COMP|92500-8|LNC|J little k super little b Ag inferred phenotype|J little k super little b Ag inferred phenotype
C5144479|T201|COMP|92501-6|LNC|J little k super little a Ag inferred phenotype|J little k super little a Ag inferred phenotype
C5144480|T201|COMP|92502-4|LNC|Hemoglobin S inferred|Hemoglobin S inferred
C5144481|T201|COMP|92503-2|LNC|H little y Ag inferred phenotype|H little y Ag inferred phenotype
C5144482|T201|COMP|92504-0|LNC|F little y super little b Ag inferred phenotype|F little y super little b Ag inferred phenotype
C5144483|T201|COMP|92505-7|LNC|F little y super little a Ag inferred phenotype|F little y super little a Ag inferred phenotype
C5144484|T201|COMP|92507-3|LNC|D little o super little b Ag inferred phenotype|D little o super little b Ag inferred phenotype
C5144485|T201|COMP|92508-1|LNC|D little o super little a Ag inferred phenotype|D little o super little a Ag inferred phenotype
C5144486|T201|COMP|92509-9|LNC|D little i super little b Ag inferred phenotype|D little i super little b Ag inferred phenotype
C5144487|T201|COMP|92510-7|LNC|D little i super little a Ag inferred phenotype|D little i super little a Ag inferred phenotype
C5144488|T201|COMP|92511-5|LNC|C little o super little b Ag inferred phenotype|C little o super little b Ag inferred phenotype
C5144489|T201|COMP|92512-3|LNC|C little o super little a Ag inferred phenotype|C little o super little a Ag inferred phenotype
C5144491|T201|COMP|92516-4|LNC|VS Ag inferred phenotype|VS Ag inferred phenotype
C5144492|T201|COMP|92517-2|LNC|V Ag inferred phenotype|V Ag inferred phenotype
C5144493|T201|COMP|92518-0|LNC|U Ag inferred phenotype|U Ag inferred phenotype
C5144494|T201|COMP|92519-8|LNC|S little c super 2 Ag inferred phenotype|S little c super 2 Ag inferred phenotype
C5144495|T201|COMP|92520-6|LNC|S little c super 1 Ag inferred phenotype|S little c super 1 Ag inferred phenotype
C5144496|T201|COMP|92522-2|LNC|N Ag inferred phenotype|N Ag inferred phenotype
C5144497|T201|COMP|92523-0|LNC|M Ag inferred phenotype|M Ag inferred phenotype
C5144498|T201|COMP|92524-8|LNC|LW super little b Ag inferred phenotype|LW super little b Ag inferred phenotype
C5144499|T201|COMP|92525-5|LNC|LW super little a Ag inferred phenotype|LW super little a Ag inferred phenotype
C5144500|T201|COMP|92530-5|LNC|L little u super little b Ag inferred phenotype|L little u super little b Ag inferred phenotype
C5144501|T201|COMP|92531-3|LNC|L little u super little a Ag inferred phenotype|L little u super little a Ag inferred phenotype
C5144502|T201|COMP|92532-1|LNC|K little p super little b Ag inferred phenotype|K little p super little b Ag inferred phenotype
C5144503|T201|COMP|92533-9|LNC|K little p super little a Ag inferred phenotype|K little p super little a Ag inferred phenotype
C5144504|T201|COMP|92535-4|LNC|J little s super little b Ag inferred phenotype|J little s super little b Ag inferred phenotype
C5144505|T201|COMP|92536-2|LNC|J little s super little a Ag inferred phenotype|J little s super little a Ag inferred phenotype
C5144506|T201|COMP|92537-0|LNC|J little o super little a Ag inferred phenotype|J little o super little a Ag inferred phenotype
C5144507|T201|COMP|92538-8|LNC|J little k super little b Ag inferred phenotype|J little k super little b Ag inferred phenotype
C5144508|T201|COMP|92539-6|LNC|J little k super little a Ag inferred phenotype|J little k super little a Ag inferred phenotype
C5144509|T201|COMP|92540-4|LNC|Hemoglobin S inferred|Hemoglobin S inferred
C5144510|T201|COMP|92541-2|LNC|H little y Ag inferred phenotype|H little y Ag inferred phenotype
C5144511|T201|COMP|92542-0|LNC|F little y super little b Ag inferred phenotype|F little y super little b Ag inferred phenotype
C5144512|T201|COMP|92543-8|LNC|F little y super little a Ag inferred phenotype|F little y super little a Ag inferred phenotype
C5144513|T201|COMP|92545-3|LNC|D little o super little b Ag inferred phenotype|D little o super little b Ag inferred phenotype
C5144514|T201|COMP|92546-1|LNC|D little o super little a Ag inferred phenotype|D little o super little a Ag inferred phenotype
C5144515|T201|COMP|92547-9|LNC|D little i super little b Ag inferred phenotype|D little i super little b Ag inferred phenotype
C5144516|T201|COMP|92548-7|LNC|D little i super little a Ag inferred phenotype|D little i super little a Ag inferred phenotype
C5144517|T201|COMP|92549-5|LNC|C little o super little b Ag inferred phenotype|C little o super little b Ag inferred phenotype
C5144518|T201|COMP|92550-3|LNC|C little o super little a Ag inferred phenotype|C little o super little a Ag inferred phenotype
C5144533|T201|COMP|92572-7|LNC|Sodium|Sodium
C5144534|T201|COMP|92577-6|LNC|Chlamydophila pneumoniae DNA|Chlamydophila pneumoniae DNA
C5144535|T201|COMP|92635-2|LNC|Leukocytes|Leukocytes
C5144536|T201|COMP|92636-0|LNC|APOL1 inferred genotype|APOL1 inferred genotype
C5144537|T201|COMP|92637-8|LNC|traZODone|traZODone
C5144538|T201|COMP|92638-6|LNC|Sertraline|Sertraline
C5144539|T201|COMP|92639-4|LNC|O-nortramadol|O-nortramadol
C5144540|T201|COMP|92640-2|LNC|M-chlorophenylpiperazine|M-chlorophenylpiperazine
C5144541|T201|COMP|92641-0|LNC|diphenhydrAMINE|diphenhydrAMINE
C5144542|T201|COMP|92642-8|LNC|Dextromethorphan|Dextromethorphan
C5144543|T201|COMP|92643-6|LNC|Cotinine|Cotinine
C5144544|T201|COMP|92644-4|LNC|Phentermine|Phentermine
C5144545|T201|COMP|92645-1|LNC|Citalopram|Citalopram
C5144546|T201|COMP|92646-9|LNC|Dextromethorphan|Dextromethorphan
C5144547|T201|COMP|92647-7|LNC|diphenhydrAMINE|diphenhydrAMINE
C5144548|T201|COMP|92648-5|LNC|Gabapentin|Gabapentin
C5144549|T201|COMP|92649-3|LNC|Naloxone|Naloxone
C5144550|T201|COMP|92650-1|LNC|PARoxetine|PARoxetine
C5144551|T201|COMP|92651-9|LNC|Pregabalin|Pregabalin
C5144552|T201|COMP|92652-7|LNC|Sertraline|Sertraline
C5144553|T201|COMP|92653-5|LNC|traZODone|traZODone
C5144554|T201|COMP|92654-3|LNC|9-hydroxyrisperidone|9-hydroxyrisperidone
C5144560|T201|COMP|92665-9|LNC|Growth and differentiation factor 15|Growth and differentiation factor 15
C5144562|T201|COMP|92667-5|LNC|Glucose^30M post dose cloNIDine|Glucose^30M post dose cloNIDine
C5144563|T201|COMP|92668-3|LNC|Glucose^1H post dose cloNIDine|Glucose^1H post dose cloNIDine
C5144564|T201|COMP|92669-1|LNC|Glucose^1.5H post dose cloNIDine|Glucose^1.5H post dose cloNIDine
C5144565|T201|COMP|92670-9|LNC|Glucose^2H post dose cloNIDine|Glucose^2H post dose cloNIDine
C5144566|T201|COMP|92671-7|LNC|Basement membrane zone BP180 & BP230 Ab.IgG panel|Basement membrane zone BP180 & BP230 Ab.IgG panel
C5144580|T201|COMP|92685-7|LNC|Trichomonas vaginalis DNA|Trichomonas vaginalis DNA
C5144581|T201|COMP|92686-5|LNC|Vibrio cholerae+parahaemolyticus+vulnificus DNA|Vibrio cholerae+parahaemolyticus+vulnificus DNA
C5144582|T201|COMP|92687-3|LNC|Giardia lamblia DNA|Giardia lamblia DNA
C5144583|T201|COMP|92688-1|LNC|Cryptosporidium parvum+hominis DNA|Cryptosporidium parvum+hominis DNA
C5144584|T201|COMP|92689-9|LNC|Entamoeba histolytica DNA|Entamoeba histolytica DNA
C5144585|T201|COMP|92690-7|LNC|Adenovirus 40+41 DNA|Adenovirus 40+41 DNA
C5144586|T201|COMP|92691-5|LNC|Astrovirus RNA|Astrovirus RNA
C5144587|T201|COMP|92692-3|LNC|Norovirus genogroup I+II RNA|Norovirus genogroup I+II RNA
C5144588|T201|COMP|92693-1|LNC|Rotavirus A RNA|Rotavirus A RNA
C5144589|T201|COMP|92694-9|LNC|Sapovirus genogroups I+II+IV+V RNA|Sapovirus genogroups I+II+IV+V RNA
C5144590|T201|COMP|92695-6|LNC|Gastrointestinal bacterial pathogens panel|Gastrointestinal bacterial pathogens panel
C5144591|T201|COMP|92696-4|LNC|Gastrointestinal viral pathogens panel|Gastrointestinal viral pathogens panel
C5144592|T201|COMP|92697-2|LNC|Gastrointestinal parasitic pathogens panel|Gastrointestinal parasitic pathogens panel
C5144593|T201|COMP|92698-0|LNC|Gardnerella vaginalis DNA|Gardnerella vaginalis DNA
C5144594|T201|COMP|92699-8|LNC|Candida sp DNA|Candida sp DNA
C5144595|T201|COMP|92700-4|LNC|Trichomonas vaginalis DNA|Trichomonas vaginalis DNA
C5144596|T201|COMP|92701-2|LNC|Staphylococcus aureus DNA|Staphylococcus aureus DNA
C5144598|T201|COMP|92703-8|LNC|Vaginal pathogens panel|Vaginal pathogens panel
C5144602|T201|COMP|92711-1|LNC|Lipoprotein.alpha.subparticle.small|Lipoprotein.alpha.subparticle.small
C5144603|T201|COMP|92712-9|LNC|Lipoprotein.beta.subparticle.very small-d|Lipoprotein.beta.subparticle.very small-d
C5144604|T201|COMP|92713-7|LNC|Lipoprotein.beta.subparticle.very small-c|Lipoprotein.beta.subparticle.very small-c
C5144605|T201|COMP|92714-5|LNC|Lipoprotein.beta.subparticle.very small-b|Lipoprotein.beta.subparticle.very small-b
C5144606|T201|COMP|92715-2|LNC|Lipoprotein.beta.subparticle.very small-a|Lipoprotein.beta.subparticle.very small-a
C5144607|T201|COMP|92716-0|LNC|Lipoprotein.beta.subparticle.large-b|Lipoprotein.beta.subparticle.large-b
C5144608|T201|COMP|92717-8|LNC|Lipoprotein.beta.subparticle.large-a|Lipoprotein.beta.subparticle.large-a
C5144609|T201|COMP|92718-6|LNC|Lipoprotein.broad beta.subparticle.small|Lipoprotein.broad beta.subparticle.small
C5144610|T201|COMP|92719-4|LNC|Lipoprotein.broad beta.subparticle.large|Lipoprotein.broad beta.subparticle.large
C5144611|T201|COMP|92720-2|LNC|Lipoprotein.pre-beta.subparticle.small|Lipoprotein.pre-beta.subparticle.small
C5144612|T201|COMP|92721-0|LNC|Lipoprotein.pre-beta.subparticle.medium|Lipoprotein.pre-beta.subparticle.medium
C5144613|T201|COMP|92722-8|LNC|Lipoprotein subparticle profile panel|Lipoprotein subparticle profile panel
C5144614|T201|COMP|92723-6|LNC|Yersinia enterocolitica DNA|Yersinia enterocolitica DNA
C5144616|T201|COMP|92726-9|LNC|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C5144617|T201|COMP|92727-7|LNC|Tacrolimus|Tacrolimus
C5144618|T201|COMP|92728-5|LNC|Tacrolimus^4H post dose|Tacrolimus^4H post dose
C5144619|T201|COMP|92729-3|LNC|Tacrolimus^2H post dose|Tacrolimus^2H post dose
C5144620|T201|COMP|92730-1|LNC|Tacrolimus^1H post dose|Tacrolimus^1H post dose
C5144621|T201|COMP|92731-9|LNC|Hepatitis C virus genotype|Hepatitis C virus genotype
C5144622|T201|COMP|92732-7|LNC|Codon &or region with poor sequence quality|Codon &or region with poor sequence quality
C5144623|T201|COMP|92733-5|LNC|Glecaprevir|Glecaprevir
C5144624|T201|COMP|92734-3|LNC|Voxilaprevir|Voxilaprevir
C5144625|T201|COMP|92735-0|LNC|Pibrentasvir|Pibrentasvir
C5144626|T201|COMP|92736-8|LNC|Cells.CD3+CD4+|Cells.CD3+CD4+
C5144630|T201|COMP|92740-0|LNC|Oxysterols panel|Oxysterols panel
C5144632|T201|COMP|92742-6|LNC|Iron.microscopic observation|Iron.microscopic observation
C5144637|T201|COMP|92747-5|LNC|Lyso-sphingomyelin|Lyso-sphingomyelin
C5144638|T201|COMP|92748-3|LNC|Lyso-sphingomyelin|Lyso-sphingomyelin
C5144639|T201|COMP|92749-1|LNC|Lyso-sphingomyelin|Lyso-sphingomyelin
C5144640|T201|COMP|92750-9|LNC|Glucopsychosine|Glucopsychosine
C5144641|T201|COMP|92751-7|LNC|Glucopsychosine|Glucopsychosine
C5144642|T201|COMP|92752-5|LNC|Glucopsychosine|Glucopsychosine
C5144643|T201|COMP|92754-1|LNC|Globotriaosylsphingosine|Globotriaosylsphingosine
C5144644|T201|COMP|92755-8|LNC|Cholestane-3-beta, 5-alpha, 6-beta triol|Cholestane-3-beta, 5-alpha, 6-beta triol
C5144645|T201|COMP|92756-6|LNC|Cholestane-3-beta, 5-alpha, 6-beta triol|Cholestane-3-beta, 5-alpha, 6-beta triol
C5144646|T201|COMP|92757-4|LNC|Cholestane-3-beta, 5-alpha, 6-beta triol|Cholestane-3-beta, 5-alpha, 6-beta triol
C5144647|T201|COMP|92758-2|LNC|7-Alpha,12-alpha dihydroxycholest-4-en-3-one|7-Alpha,12-alpha dihydroxycholest-4-en-3-one
C5144648|T201|COMP|92759-0|LNC|7-Alpha,12-alpha dihydroxycholest-4-en-3-one|7-Alpha,12-alpha dihydroxycholest-4-en-3-one
C5144649|T201|COMP|92760-8|LNC|7-Alpha,12-alpha dihydroxycholest-4-en-3-one|7-Alpha,12-alpha dihydroxycholest-4-en-3-one
C5144650|T201|COMP|92761-6|LNC|7-Alpha hydroxy-4-cholesten-3-one|7-Alpha hydroxy-4-cholesten-3-one
C5144651|T201|COMP|92762-4|LNC|7-Alpha hydroxy-4-cholesten-3-one|7-Alpha hydroxy-4-cholesten-3-one
C5144652|T201|COMP|92763-2|LNC|7-Alpha hydroxy-4-cholesten-3-one|7-Alpha hydroxy-4-cholesten-3-one
C5144653|T201|COMP|92764-0|LNC|7-Ketocholesterol|7-Ketocholesterol
C5144654|T201|COMP|92765-7|LNC|Adalimumab Ab.Neut|Adalimumab Ab.Neut
C5144656|T201|COMP|92767-3|LNC|Listeria sp DNA|Listeria sp DNA
C5144657|T201|COMP|92768-1|LNC|Candida albicans+glabrata+krusei+parapsilosis DNA|Candida albicans+glabrata+krusei+parapsilosis DNA
C5144658|T201|COMP|92769-9|LNC|Gram negative bacteria DNA|Gram negative bacteria DNA
C5144659|T201|COMP|92770-7|LNC|Streptococcus pyogenes DNA|Streptococcus pyogenes DNA
C5144660|T201|COMP|92771-5|LNC|Streptococcus pneumoniae DNA|Streptococcus pneumoniae DNA
C5144661|T201|COMP|92772-3|LNC|Streptococcus anginosus group DNA|Streptococcus anginosus group DNA
C5144662|T201|COMP|92773-1|LNC|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C5144663|T201|COMP|92774-9|LNC|Streptococcus sp DNA|Streptococcus sp DNA
C5144664|T201|COMP|92775-6|LNC|Staphylococcus lugdunensis DNA|Staphylococcus lugdunensis DNA
C5144665|T201|COMP|92776-4|LNC|Staphylococcus epidermidis DNA|Staphylococcus epidermidis DNA
C5144666|T201|COMP|92777-2|LNC|Staphylococcus aureus DNA|Staphylococcus aureus DNA
C5144667|T201|COMP|92778-0|LNC|Staphylococcus sp DNA|Staphylococcus sp DNA
C5144668|T201|COMP|92779-8|LNC|Micrococcus sp DNA|Micrococcus sp DNA
C5144669|T201|COMP|92780-6|LNC|Listeria monocytogenes DNA|Listeria monocytogenes DNA
C5144670|T201|COMP|92781-4|LNC|Lactobacillus sp DNA|Lactobacillus sp DNA
C5144671|T201|COMP|92782-2|LNC|Enterococcus faecium DNA|Enterococcus faecium DNA
C5144672|T201|COMP|92783-0|LNC|Enterococcus faecalis DNA|Enterococcus faecalis DNA
C5144673|T201|COMP|92784-8|LNC|Enterococcus sp DNA|Enterococcus sp DNA
C5144674|T201|COMP|92785-5|LNC|Cutibacterium acnes DNA|Cutibacterium acnes DNA
C5144675|T201|COMP|92786-3|LNC|Corynebacterium sp DNA|Corynebacterium sp DNA
C5144676|T201|COMP|92787-1|LNC|Bacillus subtilis group DNA|Bacillus subtilis group DNA
C5144677|T201|COMP|92788-9|LNC|Bacillus cereus group DNA|Bacillus cereus group DNA
C5144678|T201|COMP|92789-7|LNC|Gram positive blood culture panel|Gram positive blood culture panel
C5144679|T201|COMP|92790-5|LNC|Candida albicans DNA|Candida albicans DNA
C5144680|T201|COMP|92791-3|LNC|Candida auris DNA|Candida auris DNA
C5144681|T201|COMP|92792-1|LNC|Candida dubliniensis DNA|Candida dubliniensis DNA
C5144682|T201|COMP|92793-9|LNC|Candida famata DNA|Candida famata DNA
C5144683|T201|COMP|92794-7|LNC|Candida glabrata DNA|Candida glabrata DNA
C5144684|T201|COMP|92795-4|LNC|Candida guilliermondii DNA|Candida guilliermondii DNA
C5144685|T201|COMP|92796-2|LNC|Candida kefyr DNA|Candida kefyr DNA
C5144686|T201|COMP|92797-0|LNC|Candida krusei DNA|Candida krusei DNA
C5144687|T201|COMP|92798-8|LNC|Candida lusitaniae DNA|Candida lusitaniae DNA
C5144688|T201|COMP|92799-6|LNC|Candida parapsilosis DNA|Candida parapsilosis DNA
C5144689|T201|COMP|92800-2|LNC|Candida tropicalis DNA|Candida tropicalis DNA
C5144690|T201|COMP|92801-0|LNC|Cryptococcus gattii DNA|Cryptococcus gattii DNA
C5144691|T201|COMP|92802-8|LNC|Cryptococcus neoformans DNA|Cryptococcus neoformans DNA
C5144692|T201|COMP|92803-6|LNC|Fusarium sp DNA|Fusarium sp DNA
C5144693|T201|COMP|92804-4|LNC|Rhodotorula spp DNA|Rhodotorula spp DNA
C5144694|T201|COMP|92805-1|LNC|Blood fungal pathogens panel|Blood fungal pathogens panel
C5144695|T201|COMP|92806-9|LNC|Keratan sulfate/Creatinine|Keratan sulfate/Creatinine
C5144696|T201|COMP|92807-7|LNC|Rhinovirus+Enterovirus RNA|Rhinovirus+Enterovirus RNA
C5144697|T201|COMP|92808-5|LNC|Influenza virus A H3 RNA|Influenza virus A H3 RNA
C5144698|T201|COMP|92809-3|LNC|Influenza virus A H1 RNA|Influenza virus A H1 RNA
C5144699|T201|COMP|92810-1|LNC|Borrelia afzelii+burgdorferi+garinii Ab.IgG|Borrelia afzelii+burgdorferi+garinii Ab.IgG
C5144700|T201|COMP|92811-9|LNC|Borrelia afzelii+burgdorferi+garinii Ab.IgG index|Borrelia afzelii+burgdorferi+garinii Ab.IgG index
C5144701|T201|COMP|92812-7|LNC|Borrelia afzelii+burgdorferi+garinii Ab.IgG|Borrelia afzelii+burgdorferi+garinii Ab.IgG
C5144702|T201|COMP|92813-5|LNC|Borrelia afzelii+burgdorferi+garinii Ab.IgG|Borrelia afzelii+burgdorferi+garinii Ab.IgG
C5144703|T201|COMP|92814-3|LNC|Borrelia afzelii+burgdorferi+garinii Ab.IgG|Borrelia afzelii+burgdorferi+garinii Ab.IgG
C5144704|T201|COMP|92815-0|LNC|Borrelia afzelii+burgdorferi+garinii Ab.IgG panel|Borrelia afzelii+burgdorferi+garinii Ab.IgG panel
C5144705|T201|COMP|92816-8|LNC|Phencyclidine|Phencyclidine
C5144706|T201|COMP|92817-6|LNC|Glucose^30M post dose glucagon|Glucose^30M post dose glucagon
C5144707|T201|COMP|92818-4|LNC|Glucose^20M post dose glucagon|Glucose^20M post dose glucagon
C5144708|T201|COMP|92819-2|LNC|Glucose^10M post dose glucagon|Glucose^10M post dose glucagon
C5144709|T201|COMP|92820-0|LNC|Glucose post glucagon stimulation panel|Glucose post glucagon stimulation panel
C5144710|T201|COMP|92821-8|LNC|Allelic frequency|Allelic frequency
C5144711|T201|COMP|92822-6|LNC|Genomic coordinate system|Genomic coordinate system
C5144713|T201|COMP|92825-9|LNC|Renin^upright|Renin^upright
C5144714|T201|COMP|92826-7|LNC|Renin^supine|Renin^supine
C5144716|T201|COMP|92828-3|LNC|Adenovirus B+E DNA|Adenovirus B+E DNA
C5144717|T201|COMP|92829-1|LNC|Location of metastasis within sentinel lymph node|Location of metastasis within sentinel lymph node
C5144718|T201|COMP|92830-9|LNC|Sentinel lymph node extranodal extension|Sentinel lymph node extranodal extension
C5144719|T201|COMP|92831-7|LNC|Lymph nodes with metastasis|Lymph nodes with metastasis
C5144720|T201|COMP|92832-5|LNC|Sentinel lymph nodes with metastasis|Sentinel lymph nodes with metastasis
C5144721|T201|COMP|92833-3|LNC|Lymph nodes examined|Lymph nodes examined
C5144722|T201|COMP|92834-1|LNC|Tumor regression at peripheral margin|Tumor regression at peripheral margin
C5144723|T201|COMP|92835-8|LNC|Associated nevus|Associated nevus
C5144724|T201|COMP|92836-6|LNC|Desmoplastic melanoma|Desmoplastic melanoma
C5144725|T201|COMP|92837-4|LNC|Perineural invasion|Perineural invasion
C5144726|T201|COMP|92838-2|LNC|Satellite nodules|Satellite nodules
C5144728|T201|COMP|92843-2|LNC|FLT3 gene.p.Asp835 mutations|FLT3 gene.p.Asp835 mutations
C5144729|T201|COMP|92844-0|LNC|FLT3 gene internal tandem duplication/normal|FLT3 gene internal tandem duplication/normal
C5144730|T201|COMP|92845-7|LNC|Insulin resistance score|Insulin resistance score
C5144732|T201|COMP|92848-1|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C5144736|T201|COMP|92852-3|LNC|Adenovirus & Bocavirus DNA panel|Adenovirus & Bocavirus DNA panel
C5144737|T201|COMP|92853-1|LNC|Adenovirus & Bocavirus DNA panel|Adenovirus & Bocavirus DNA panel
C5144738|T201|COMP|92854-9|LNC|Adenovirus DNA|Adenovirus DNA
C5144739|T201|COMP|92855-6|LNC|Bordetella parapertussis IS1001 DNA|Bordetella parapertussis IS1001 DNA
C5144740|T201|COMP|92856-4|LNC|Bordetella parapertussis IS1001 DNA|Bordetella parapertussis IS1001 DNA
C5144747|T201|COMP|92863-0|LNC|Herpes simplex virus 1 & 2 DNA panel|Herpes simplex virus 1 & 2 DNA panel
C5144748|T201|COMP|92864-8|LNC|Herpes simplex virus 1 & 2 DNA panel|Herpes simplex virus 1 & 2 DNA panel
C5144749|T201|COMP|92865-5|LNC|Herpes simplex virus 1 & 2 DNA panel|Herpes simplex virus 1 & 2 DNA panel
C5144750|T201|COMP|92866-3|LNC|Herpes simplex virus 1 & 2 DNA panel|Herpes simplex virus 1 & 2 DNA panel
C5144751|T201|COMP|92867-1|LNC|Herpes simplex virus 1 & 2 DNA panel|Herpes simplex virus 1 & 2 DNA panel
C5144752|T201|COMP|92868-9|LNC|Herpes simplex virus 1 & 2 DNA panel|Herpes simplex virus 1 & 2 DNA panel
C5144753|T201|COMP|92869-7|LNC|Herpes simplex virus 1 & 2 DNA panel|Herpes simplex virus 1 & 2 DNA panel
C5144754|T201|COMP|92870-5|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C5144755|T201|COMP|92871-3|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C5144756|T201|COMP|92872-1|LNC|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C5144757|T201|COMP|92873-9|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C5144758|T201|COMP|92874-7|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C5144759|T201|COMP|92875-4|LNC|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C5144762|T201|COMP|92878-8|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA|Human coronavirus 229E+HKU1+NL63+OC43 RNA
C5144763|T201|COMP|92879-6|LNC|Human coronavirus 229E+HKU1+NL63+OC43 RNA|Human coronavirus 229E+HKU1+NL63+OC43 RNA
C5144766|T201|COMP|92882-0|LNC|Influenza virus A & B RNA panel|Influenza virus A & B RNA panel
C5144767|T201|COMP|92883-8|LNC|Parainfluenza virus 1+2+3+4 RNA|Parainfluenza virus 1+2+3+4 RNA
C5144768|T201|COMP|92884-6|LNC|Parainfluenza virus 1+2+3+4 RNA|Parainfluenza virus 1+2+3+4 RNA
C5144769|T201|COMP|92885-3|LNC|Rhinovirus+Enterovirus RNA|Rhinovirus+Enterovirus RNA
C5144770|T201|COMP|92886-1|LNC|Torque teno virus DNA|Torque teno virus DNA
C5144771|T201|COMP|92887-9|LNC|Torque teno virus DNA|Torque teno virus DNA
C5144772|T201|COMP|92888-7|LNC|Varicella zoster virus DNA|Varicella zoster virus DNA
C5144775|T201|COMP|92891-1|LNC|Coagulation tissue factor induced.INR goal|Coagulation tissue factor induced.INR goal
C5144776|T201|COMP|92896-0|LNC|Aldosterone|Aldosterone
C5144777|T201|COMP|92897-8|LNC|Aldosterone|Aldosterone
C5144779|T201|COMP|92899-4|LNC|Fetal chromosome region 11q23 deletion|Fetal chromosome region 11q23 deletion
C5144780|T201|COMP|92900-0|LNC|Fetal chromosome region 4p16 deletion|Fetal chromosome region 4p16 deletion
C5144782|T201|COMP|92902-6|LNC|Fetal chromosome region 8q24 deletion|Fetal chromosome region 8q24 deletion
C5144783|T201|COMP|92903-4|LNC|Fetal chromosome region 15q11 deletion|Fetal chromosome region 15q11 deletion
C5144784|T201|COMP|92904-2|LNC|N-nortramadol|N-nortramadol
C5144785|T201|COMP|92905-9|LNC|Chromosome 7 copy number/nucleus|Chromosome 7 copy number/nucleus
C5144786|T201|COMP|92906-7|LNC|MET gene copy number/nucleus|MET gene copy number/nucleus
C5144787|T201|COMP|92907-5|LNC|MET gene copy number/Chromosome 7 copy number|MET gene copy number/Chromosome 7 copy number
C5144809|T201|COMP|92929-9|LNC|Measles & Mumps & Rubella virus Ab.IgG panel|Measles & Mumps & Rubella virus Ab.IgG panel
C5144810|T201|COMP|92930-7|LNC|LPA gene.c.3947+467T>C|LPA gene.c.3947+467T>C
C5144811|T201|COMP|92931-5|LNC|LPA gene.c.5673A>G|LPA gene.c.5673A>G
C5144812|T201|COMP|92932-3|LNC|KIF6 gene.c.2155T>C|KIF6 gene.c.2155T>C
C5144813|T201|COMP|92933-1|LNC|9p21 g.22125503G>C|9p21 g.22125503G>C
C5144814|T201|COMP|92934-9|LNC|9p21 g.22124478A>G|9p21 g.22124478A>G
C5144815|T201|COMP|92935-6|LNC|4q25 g.111720761T>G|4q25 g.111720761T>G
C5144816|T201|COMP|92936-4|LNC|4q25 g.111710169C>T|4q25 g.111710169C>T
C5144817|T201|COMP|92937-2|LNC|Eslicarbazepine|Eslicarbazepine
C5144818|T201|COMP|92938-0|LNC|Catecholamines 3 panel|Catecholamines 3 panel
C5144821|T201|COMP|92946-3|LNC|Streptococcus pyogenes DNA|Streptococcus pyogenes DNA
C5144822|T201|COMP|92947-1|LNC|Streptococcus pyogenes DNA|Streptococcus pyogenes DNA
C5144823|T201|COMP|92948-9|LNC|Streptococcus pneumoniae DNA|Streptococcus pneumoniae DNA
C5144824|T201|COMP|92949-7|LNC|Streptococcus pneumoniae DNA|Streptococcus pneumoniae DNA
C5144825|T201|COMP|92950-5|LNC|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C5144826|T201|COMP|92951-3|LNC|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C5144827|T201|COMP|92952-1|LNC|Staphylococcus aureus DNA|Staphylococcus aureus DNA
C5144828|T201|COMP|92953-9|LNC|Staphylococcus aureus DNA|Staphylococcus aureus DNA
C5144829|T201|COMP|92954-7|LNC|Serratia marcescens DNA|Serratia marcescens DNA
C5144830|T201|COMP|92955-4|LNC|Serratia marcescens DNA|Serratia marcescens DNA
C5144831|T201|COMP|92956-2|LNC|Rhinovirus+Enterovirus RNA|Rhinovirus+Enterovirus RNA
C5144832|T201|COMP|92957-0|LNC|Respiratory syncytial virus RNA|Respiratory syncytial virus RNA
C5144833|T201|COMP|92958-8|LNC|Respiratory pathogens DNA & RNA panel|Respiratory pathogens DNA & RNA panel
C5144834|T201|COMP|92959-6|LNC|Pseudomonas aeruginosa DNA|Pseudomonas aeruginosa DNA
C5144835|T201|COMP|92960-4|LNC|Pseudomonas aeruginosa DNA|Pseudomonas aeruginosa DNA
C5144836|T201|COMP|92961-2|LNC|Proteus sp DNA|Proteus sp DNA
C5144837|T201|COMP|92962-0|LNC|Proteus sp DNA|Proteus sp DNA
C5144838|T201|COMP|92963-8|LNC|Parainfluenza virus RNA|Parainfluenza virus RNA
C5144839|T201|COMP|92964-6|LNC|Mycoplasma pneumoniae DNA|Mycoplasma pneumoniae DNA
C5144840|T201|COMP|92965-3|LNC|Moraxella catarrhalis DNA|Moraxella catarrhalis DNA
C5144841|T201|COMP|92966-1|LNC|Moraxella catarrhalis DNA|Moraxella catarrhalis DNA
C5144842|T201|COMP|92967-9|LNC|Middle East respiratory syndrome coronavirus RNA|Middle East respiratory syndrome coronavirus RNA
C5144843|T201|COMP|92968-7|LNC|Bacterial methicillin resistance mecA+mecC genes|Bacterial methicillin resistance mecA+mecC genes
C5144844|T201|COMP|92969-5|LNC|Legionella pneumophila DNA|Legionella pneumophila DNA
C5144845|T201|COMP|92970-3|LNC|Klebsiella pneumoniae DNA|Klebsiella pneumoniae DNA
C5144846|T201|COMP|92971-1|LNC|Klebsiella pneumoniae DNA|Klebsiella pneumoniae DNA
C5144847|T201|COMP|92972-9|LNC|Klebsiella oxytoca DNA|Klebsiella oxytoca DNA
C5144848|T201|COMP|92973-7|LNC|Klebsiella oxytoca DNA|Klebsiella oxytoca DNA
C5144849|T201|COMP|92974-5|LNC|Klebsiella aerogenes DNA|Klebsiella aerogenes DNA
C5144850|T201|COMP|92975-2|LNC|Klebsiella aerogenes DNA|Klebsiella aerogenes DNA
C5144851|T201|COMP|92976-0|LNC|Influenza virus B RNA|Influenza virus B RNA
C5144852|T201|COMP|92977-8|LNC|Influenza virus A RNA|Influenza virus A RNA
C5144853|T201|COMP|92978-6|LNC|Human Metapneumovirus RNA|Human Metapneumovirus RNA
C5144854|T201|COMP|92979-4|LNC|Human Coronavirus RNA|Human Coronavirus RNA
C5144855|T201|COMP|92980-2|LNC|Haemophilus influenzae DNA|Haemophilus influenzae DNA
C5144856|T201|COMP|92981-0|LNC|Haemophilus influenzae DNA|Haemophilus influenzae DNA
C5144857|T201|COMP|92982-8|LNC|Escherichia coli DNA|Escherichia coli DNA
C5144858|T201|COMP|92983-6|LNC|Escherichia coli DNA|Escherichia coli DNA
C5144859|T201|COMP|92984-4|LNC|Enterobacter cloacae complex DNA|Enterobacter cloacae complex DNA
C5144860|T201|COMP|92985-1|LNC|Enterobacter cloacae complex DNA|Enterobacter cloacae complex DNA
C5144861|T201|COMP|92986-9|LNC|Chlamydophila pneumoniae DNA|Chlamydophila pneumoniae DNA
C5144862|T201|COMP|92987-7|LNC|Adenovirus DNA|Adenovirus DNA
C5144863|T201|COMP|92988-5|LNC|Acinetobacter baumannii DNA|Acinetobacter baumannii DNA
C5144864|T201|COMP|92989-3|LNC|Acinetobacter baumannii DNA|Acinetobacter baumannii DNA
C5144865|T201|COMP|92990-1|LNC|F10 gene full mutation analysis|F10 gene full mutation analysis
C5144866|T201|COMP|92991-9|LNC|F13A1 gene & F13B gene full mutation analysis|F13A1 gene & F13B gene full mutation analysis
C5144868|T201|COMP|92993-5|LNC|PROCR gene full mutation analysis|PROCR gene full mutation analysis
C5144869|T201|COMP|92994-3|LNC|PROS1 gene full mutation analysis|PROS1 gene full mutation analysis
C5144870|T201|COMP|92995-0|LNC|THBD gene full mutation analysis|THBD gene full mutation analysis
C5144880|T201|COMP|93017-2|LNC|Plasma cells.abnormal marker pattern|Plasma cells.abnormal marker pattern
C5144881|T201|COMP|93018-0|LNC|Plasma cells.polyclonal|Plasma cells.polyclonal
C5144882|T201|COMP|93019-8|LNC|Plasma cells|Plasma cells
C5144883|T201|COMP|93020-6|LNC|Plasma cells.polyclonal/Plasma cells.total|Plasma cells.polyclonal/Plasma cells.total
C5144885|T201|COMP|93022-2|LNC|Multiple myeloma minimal residual disease panel|Multiple myeloma minimal residual disease panel
C5144903|T201|COMP|93045-3|LNC|Carbon monoxide|Carbon monoxide
C5144904|T201|COMP|93048-7|LNC|Reason for specimen rejection|Reason for specimen rejection
C5144912|T201|COMP|92753-3|LNC|Globotriaosylsphingosine|Globotriaosylsphingosine
C5144913|T201|COMP|92839-0|LNC|Breslow thickness|Breslow thickness
C5144917|T201|COMP|91900-1|LNC|Parasite|Parasite
C5200951|T201|COMP|35185-8|LNC|Aldosterone|Aldosterone
C5200952|T201|COMP|35186-6|LNC|Aldosterone|Aldosterone
C5200953|T201|COMP|35187-4|LNC|Aldosterone^supine|Aldosterone^supine
C5200954|T201|COMP|35189-0|LNC|Androstanolone|Androstanolone
C5200955|T201|COMP|35191-6|LNC|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C5200956|T201|COMP|35192-4|LNC|Bilirubin.non-glucuronidated|Bilirubin.non-glucuronidated
C5200957|T201|COMP|35193-2|LNC|Bilirubin|Bilirubin
C5200958|T201|COMP|35196-5|LNC|Calcidiol|Calcidiol
C5200959|T201|COMP|35202-1|LNC|Cortisol|Cortisol
C5200960|T201|COMP|35242-7|LNC|Creatinine|Creatinine
C5200961|T201|COMP|35204-7|LNC|Creatinine|Creatinine
C5200962|T201|COMP|35262-5|LNC|Creatinine|Creatinine
C5200963|T201|COMP|35208-8|LNC|Estrone|Estrone
C5200964|T201|COMP|66734-5|LNC|Glucagon|Glucagon
C5200965|T201|COMP|35237-7|LNC|carBAMazepine|carBAMazepine
C5200966|T201|COMP|35240-1|LNC|Ethanol|Ethanol
C5200985|T201|COMP|35194-0|LNC|Bilirubin|Bilirubin
C5200986|T201|COMP|35207-0|LNC|Estradiol|Estradiol
C5201097|T201|COMP|35246-8|LNC|Calcium|Calcium
C5201098|T201|COMP|35247-6|LNC|Calcium|Calcium
C5201099|T201|COMP|35248-4|LNC|Calcium|Calcium
C5201100|T201|COMP|35251-8|LNC|Creatinine|Creatinine
C5201101|T201|COMP|35254-2|LNC|Ammonia|Ammonia
C5201102|T201|COMP|35258-3|LNC|Calcium^^corrected for total protein|Calcium^^corrected for total protein
C5201103|T201|COMP|35261-7|LNC|Cortisol.free|Cortisol.free
C5201128|T201|COMP|42567-8|LNC|Calcium.ionized|Calcium.ionized
C5203189|T201|COMP|93904-1|LNC|Transfusion reaction panel|Transfusion reaction panel
C5203317|T201|COMP|93479-4|LNC|Observation interpretation|Observation interpretation
C5203361|T201|COMP|93936-3|LNC|little c Ag^during infancy|little c Ag^during infancy
C5203362|T201|COMP|93938-9|LNC|C Ag^during infancy|C Ag^during infancy
C5203363|T201|COMP|93944-7|LNC|little c Ag|little c Ag
C5203364|T201|COMP|93946-2|LNC|C Ag|C Ag
C5203366|T201|COMP|94141-9|LNC|HEDIS 2020 Value Set - Mammography|HEDIS 2020 Value Set - Mammography
C5203435|T201|COMP|93927-2|LNC|E Ag^post hematopoietic stem cell transplant|E Ag^post hematopoietic stem cell transplant
C5203535|T201|COMP|93928-0|LNC|C Ag^post hematopoietic stem cell transplant|C Ag^post hematopoietic stem cell transplant
C5203536|T201|COMP|93921-5|LNC|C Ag^post transfusion reaction|C Ag^post transfusion reaction
C5203537|T201|COMP|93919-9|LNC|little c Ag^post transfusion reaction|little c Ag^post transfusion reaction
C5203538|T201|COMP|93199-8|LNC|DPYD gene targeted mutation analysis|DPYD gene targeted mutation analysis
C5203539|T201|COMP|93943-9|LNC|little e Ag|little e Ag
C5203540|T201|COMP|93945-4|LNC|E Ag|E Ag
C5203541|T201|COMP|93935-5|LNC|little e Ag^during infancy|little e Ag^during infancy
C5203542|T201|COMP|93937-1|LNC|E Ag^during infancy|E Ag^during infancy
C5203543|T201|COMP|93920-7|LNC|E Ag^post transfusion reaction|E Ag^post transfusion reaction
C5203544|T201|COMP|93918-1|LNC|little e Ag^post transfusion reaction|little e Ag^post transfusion reaction
C5203588|T201|COMP|93912-4|LNC|CE Ag|CE Ag
C5203605|T201|COMP|94142-7|LNC|HEDIS 2020 Value Set - Urine Protein Tests|HEDIS 2020 Value Set - Urine Protein Tests
C5203616|T201|COMP|94138-5|LNC|HEDIS 2020 Value Set - BMI|HEDIS 2020 Value Set - BMI
C5203619|T201|COMP|94139-3|LNC|HEDIS 2020 Value Set - BMI percentile|HEDIS 2020 Value Set - BMI percentile
C5203621|T201|COMP|94140-1|LNC|HEDIS 2020 Value Set - CT Colonography|HEDIS 2020 Value Set - CT Colonography
C5203622|T201|COMP|94143-5|LNC|HEDIS 2020 Value Set - Diastolic Blood Pressure|HEDIS 2020 Value Set - Diastolic Blood Pressure
C5203624|T201|COMP|94144-3|LNC|HEDIS 2020 Value Set - Systolic Blood Pressure|HEDIS 2020 Value Set - Systolic Blood Pressure
C5203626|T201|COMP|94137-7|LNC|HEDIS 2020 Value Sets|HEDIS 2020 Value Sets
C5211430|T201|COMP|93085-9|LNC|Dirofilaria immitis Ab.IgG|Dirofilaria immitis Ab.IgG
C5211499|T201|COMP|93121-2|LNC|Gabapentin|Gabapentin
C5211621|T201|COMP|93190-7|LNC|HTR2A gene.c.614-2211T>C|HTR2A gene.c.614-2211T>C
C5211623|T201|COMP|93191-5|LNC|HTR2C gene.c.-759C>T|HTR2C gene.c.-759C>T
C5211624|T201|COMP|93192-3|LNC|HTR2C gene.c.551-3008C>G|HTR2C gene.c.551-3008C>G
C5211628|T201|COMP|93194-9|LNC|NUDT15 gene targeted mutation analysis|NUDT15 gene targeted mutation analysis
C5211632|T201|COMP|93196-4|LNC|Warfarin response genotype panel|Warfarin response genotype panel
C5211634|T201|COMP|93197-2|LNC|CYP4F2 gene.c.1297G>A|CYP4F2 gene.c.1297G>A
C5211636|T201|COMP|93198-0|LNC|10q23 g.94645745G>A|10q23 g.94645745G>A
C5211638|T201|COMP|93200-4|LNC|Ehlers-Danlos syndrome multigene analysis|Ehlers-Danlos syndrome multigene analysis
C5211640|T201|COMP|93201-2|LNC|Coronary heart disease multigene analysis|Coronary heart disease multigene analysis
C5211684|T201|COMP|93224-4|LNC|Coccidioides sp Ag|Coccidioides sp Ag
C5211686|T201|COMP|93225-1|LNC|Coccidioides sp Ag|Coccidioides sp Ag
C5211687|T201|COMP|93226-9|LNC|Coccidioides sp Ag|Coccidioides sp Ag
C5211688|T201|COMP|93227-7|LNC|Coccidioides sp Ag|Coccidioides sp Ag
C5211697|T201|COMP|93232-7|LNC|Imipenem+Relebactam|Imipenem+Relebactam
C5211698|T201|COMP|93233-5|LNC|Intercellular substance Ab.IgG|Intercellular substance Ab.IgG
C5211707|T201|COMP|93242-6|LNC|11-Ketotestosterone|11-Ketotestosterone
C5211708|T201|COMP|93243-4|LNC|11-Hydroxytestosterone|11-Hydroxytestosterone
C5211709|T201|COMP|93244-2|LNC|Complement Sc5b-9|Complement Sc5b-9
C5211792|T201|COMP|93313-5|LNC|Platelet glycoprotein disorder|Platelet glycoprotein disorder
C5211794|T201|COMP|93314-3|LNC|Platelet glycoprotein VI actual/normal|Platelet glycoprotein VI actual/normal
C5211796|T201|COMP|93315-0|LNC|Platelet CD49b actual/normal|Platelet CD49b actual/normal
C5211798|T201|COMP|93316-8|LNC|Platelet CD42b actual/normal|Platelet CD42b actual/normal
C5211800|T201|COMP|93317-6|LNC|Platelet CD42a actual/normal|Platelet CD42a actual/normal
C5211802|T201|COMP|93318-4|LNC|Platelet CD61 actual/normal|Platelet CD61 actual/normal
C5211804|T201|COMP|93319-2|LNC|Platelet CD41 actual/normal|Platelet CD41 actual/normal
C5211806|T201|COMP|93320-0|LNC|Platelet glycoprotein disorder panel|Platelet glycoprotein disorder panel
C5211808|T201|COMP|93321-8|LNC|PT mixing study panel|PT mixing study panel
C5211810|T201|COMP|93323-4|LNC|Tauroursodeoxycholate|Tauroursodeoxycholate
C5211811|T201|COMP|93324-2|LNC|Taurolithocholate|Taurolithocholate
C5211812|T201|COMP|93325-9|LNC|Taurohyodeoxycholate|Taurohyodeoxycholate
C5211814|T201|COMP|93326-7|LNC|Taurodeoxycholate|Taurodeoxycholate
C5211815|T201|COMP|93327-5|LNC|Taurocholate|Taurocholate
C5211816|T201|COMP|93328-3|LNC|Taurochenodeoxycholate|Taurochenodeoxycholate
C5211817|T201|COMP|93329-1|LNC|Hyodeoxycholate|Hyodeoxycholate
C5211819|T201|COMP|93330-9|LNC|Glycoursodeoxycholate|Glycoursodeoxycholate
C5211821|T201|COMP|93331-7|LNC|Glycolithocholate|Glycolithocholate
C5211822|T201|COMP|93332-5|LNC|Glycohyodeoxycholate|Glycohyodeoxycholate
C5211824|T201|COMP|93333-3|LNC|Glycodeoxycholate|Glycodeoxycholate
C5211825|T201|COMP|93334-1|LNC|Glycocholate|Glycocholate
C5211826|T201|COMP|93335-8|LNC|Glycochenodeoxycholate|Glycochenodeoxycholate
C5211827|T201|COMP|93336-6|LNC|Bile acid|Bile acid
C5211828|T201|COMP|93337-4|LNC|Chenodeoxycholate+Cholate/Bile acid.total|Chenodeoxycholate+Cholate/Bile acid.total
C5211830|T201|COMP|93338-2|LNC|Bile acid panel|Bile acid panel
C5211831|T201|COMP|93339-0|LNC|Thrombospondin type I domain-containing 7A Ab.IgG|Thrombospondin type I domain-containing 7A Ab.IgG
C5211839|T201|COMP|93345-7|LNC|Genetic variant effect on drug resistance|Genetic variant effect on drug resistance
C5211841|T201|COMP|93346-5|LNC|Genetic variant effect on drug sensitivity|Genetic variant effect on drug sensitivity
C5211849|T201|COMP|93350-7|LNC|Monocytes.HLA-DR/100 Monocytes|Monocytes.HLA-DR/100 Monocytes
C5211851|T201|COMP|93351-5|LNC|HLA-DR Ag|HLA-DR Ag
C5211852|T201|COMP|93352-3|LNC|Neutrophils.CD64/100 Neutrophils|Neutrophils.CD64/100 Neutrophils
C5211854|T201|COMP|93353-1|LNC|CD64 Ag|CD64 Ag
C5211855|T201|COMP|93354-9|LNC|Neutrophil CD64 & Monocyte HLA DR panel|Neutrophil CD64 & Monocyte HLA DR panel
C5211857|T201|COMP|93356-4|LNC|Cells.cytogenetic abnormality|Cells.cytogenetic abnormality
C5211861|T201|COMP|93358-0|LNC|Plasma cells.polyclonal/Cells counted|Plasma cells.polyclonal/Cells counted
C5211863|T201|COMP|93359-8|LNC|Monotypic plasma cell DNA ploidy|Monotypic plasma cell DNA ploidy
C5211865|T201|COMP|93360-6|LNC|Monotypic plasma cell DNA index|Monotypic plasma cell DNA index
C5211867|T201|COMP|93361-4|LNC|Plasma cells.monotypic.S phase/100 cells|Plasma cells.monotypic.S phase/100 cells
C5211869|T201|COMP|93362-2|LNC|Plasma cells.monotypic population|Plasma cells.monotypic population
C5211870|T201|COMP|93363-0|LNC|Plasma cell DNA content & proliferation panel|Plasma cell DNA content & proliferation panel
C5211872|T201|COMP|93364-8|LNC|Genetic variant diagnostic significance|Genetic variant diagnostic significance
C5211874|T201|COMP|93365-5|LNC|Genetic variant prognostic significance|Genetic variant prognostic significance
C5211876|T201|COMP|93366-3|LNC|Gene studied with no variant found|Gene studied with no variant found
C5211878|T201|COMP|93367-1|LNC|Variant of unknown significance|Variant of unknown significance
C5211879|T201|COMP|93368-9|LNC|Summary of interaction between genetic variants|Summary of interaction between genetic variants
C5211881|T201|COMP|93369-7|LNC|Krebs von den Lungen-6|Krebs von den Lungen-6
C5211884|T201|COMP|93371-3|LNC|von Willebrand factor cleaving protease activity|von Willebrand factor cleaving protease activity
C5211890|T201|COMP|93384-6|LNC|Serratia sp DNA|Serratia sp DNA
C5211892|T201|COMP|93385-3|LNC|Salmonella sp DNA|Salmonella sp DNA
C5211893|T201|COMP|93386-1|LNC|Pseudomonas aeruginosa DNA|Pseudomonas aeruginosa DNA
C5211894|T201|COMP|93387-9|LNC|Proteus mirabilis DNA|Proteus mirabilis DNA
C5211895|T201|COMP|93388-7|LNC|Neisseria meningitidis DNA|Neisseria meningitidis DNA
C5211896|T201|COMP|93389-5|LNC|Gram positive bacteria DNA|Gram positive bacteria DNA
C5211900|T201|COMP|93391-1|LNC|Stenotrophomonas maltophilia DNA|Stenotrophomonas maltophilia DNA
C5211901|T201|COMP|93392-9|LNC|Serratia marcescens DNA|Serratia marcescens DNA
C5211902|T201|COMP|93393-7|LNC|Proteus sp DNA|Proteus sp DNA
C5211903|T201|COMP|93394-5|LNC|Morganella morganii DNA|Morganella morganii DNA
C5211905|T201|COMP|93395-2|LNC|Klebsiella pneumoniae DNA|Klebsiella pneumoniae DNA
C5211906|T201|COMP|93396-0|LNC|Fusobacterium nucleatum DNA|Fusobacterium nucleatum DNA
C5211908|T201|COMP|93397-8|LNC|Haemophilus influenzae DNA|Haemophilus influenzae DNA
C5211909|T201|COMP|93398-6|LNC|Klebsiella oxytoca DNA|Klebsiella oxytoca DNA
C5211910|T201|COMP|93399-4|LNC|Fusobacterium necrophorum DNA|Fusobacterium necrophorum DNA
C5211914|T201|COMP|93401-8|LNC|Escherichia coli DNA|Escherichia coli DNA
C5211915|T201|COMP|93402-6|LNC|Cronobacter sakazakii DNA|Cronobacter sakazakii DNA
C5211917|T201|COMP|93403-4|LNC|Citrobacter sp DNA|Citrobacter sp DNA
C5211919|T201|COMP|93404-2|LNC|Enterobacter cloacae complex DNA|Enterobacter cloacae complex DNA
C5211920|T201|COMP|93405-9|LNC|Bacteroides fragilis DNA|Bacteroides fragilis DNA
C5211921|T201|COMP|93406-7|LNC|Acinetobacter baumannii DNA|Acinetobacter baumannii DNA
C5211922|T201|COMP|93407-5|LNC|Gram negative blood culture panel|Gram negative blood culture panel
C5211924|T201|COMP|93409-1|LNC|Platelet aggregation.epinephrine induced^5 umol/L|Platelet aggregation.epinephrine induced^5 umol/L
C5211925|T201|COMP|93410-9|LNC|Platelet aggregation.ristocetin induced^5 ug/mL|Platelet aggregation.ristocetin induced^5 ug/mL
C5211928|T201|COMP|93412-5|LNC|SLCO1B1 gene targeted mutation analysis|SLCO1B1 gene targeted mutation analysis
C5211938|T201|COMP|93418-2|LNC|(8;8)(q13;q21)(HEY1,NCOA2) fusion transcript|(8;8)(q13;q21)(HEY1,NCOA2) fusion transcript
C5211940|T201|COMP|93419-0|LNC|Alpha 1 antitrypsin fecal clearance panel|Alpha 1 antitrypsin fecal clearance panel
C5211942|T201|COMP|93420-8|LNC|APOA1 gene full mutation analysis|APOA1 gene full mutation analysis
C5211944|T201|COMP|93421-6|LNC|Glial fibrillary acidic protein Ab.IgG|Glial fibrillary acidic protein Ab.IgG
C5211946|T201|COMP|93422-4|LNC|Glial fibrillary acidic protein.alpha Ab.IgG|Glial fibrillary acidic protein.alpha Ab.IgG
C5211948|T201|COMP|93423-2|LNC|Glial fibrillary acidic protein Ab.IgG|Glial fibrillary acidic protein Ab.IgG
C5211949|T201|COMP|93424-0|LNC|Glial fibrillary acidic protein.alpha Ab.IgG|Glial fibrillary acidic protein.alpha Ab.IgG
C5211950|T201|COMP|93425-7|LNC|Gamma aminobutyrate B receptor Ab.IgG|Gamma aminobutyrate B receptor Ab.IgG
C5211951|T201|COMP|93426-5|LNC|Gamma aminobutyrate B receptor Ab.IgG|Gamma aminobutyrate B receptor Ab.IgG
C5211952|T201|COMP|93427-3|LNC|Gamma aminobutyrate B receptor Ab.IgG|Gamma aminobutyrate B receptor Ab.IgG
C5211953|T201|COMP|93428-1|LNC|Gamma aminobutyrate B receptor Ab.IgG|Gamma aminobutyrate B receptor Ab.IgG
C5211954|T201|COMP|93429-9|LNC|Blastomyces sp Ag|Blastomyces sp Ag
C5211956|T201|COMP|93430-7|LNC|Blastomyces sp Ag|Blastomyces sp Ag
C5211957|T201|COMP|93431-5|LNC|Blastomyces sp Ag|Blastomyces sp Ag
C5211958|T201|COMP|93432-3|LNC|Blastomyces sp Ag|Blastomyces sp Ag
C5211959|T201|COMP|93433-1|LNC|Busulfan^4H post busulfan infusion completion|Busulfan^4H post busulfan infusion completion
C5211960|T201|COMP|93434-9|LNC|Busulfan^2H post busulfan infusion completion|Busulfan^2H post busulfan infusion completion
C5211961|T201|COMP|93435-6|LNC|Busulfan^1H post busulfan infusion completion|Busulfan^1H post busulfan infusion completion
C5211963|T201|COMP|93437-2|LNC|Lurasidone|Lurasidone
C5211964|T201|COMP|93438-0|LNC|Herpes Simplex Virus 2 DNA|Herpes Simplex Virus 2 DNA
C5211965|T201|COMP|93439-8|LNC|Herpes Simplex Virus 1 DNA|Herpes Simplex Virus 1 DNA
C5211966|T201|COMP|93440-6|LNC|Herpes Simplex Virus 1 & 2 DNA Panel|Herpes Simplex Virus 1 & 2 DNA Panel
C5211969|T201|COMP|93450-5|LNC|Coagulation factor VIII Inhibitor|Coagulation factor VIII Inhibitor
C5211970|T201|COMP|93451-3|LNC|Nor-W-18+Nor-W-15|Nor-W-18+Nor-W-15
C5211972|T201|COMP|93452-1|LNC|W-19|W-19
C5211974|T201|COMP|93453-9|LNC|W-15|W-15
C5211976|T201|COMP|93454-7|LNC|W-18|W-18
C5211978|T201|COMP|93455-4|LNC|IC-26|IC-26
C5211980|T201|COMP|93456-2|LNC|MT-45|MT-45
C5211981|T201|COMP|93457-0|LNC|AH-8529|AH-8529
C5211983|T201|COMP|93458-8|LNC|AH-8533|AH-8533
C5211985|T201|COMP|93459-6|LNC|U-47700|U-47700
C5211986|T201|COMP|93460-4|LNC|AH-7921|AH-7921
C5211987|T201|COMP|93461-2|LNC|4-Methoxybutyrylfentanyl|4-Methoxybutyrylfentanyl
C5211989|T201|COMP|93462-0|LNC|Norcarfentanil|Norcarfentanil
C5211991|T201|COMP|93463-8|LNC|Ocfentanil|Ocfentanil
C5211992|T201|COMP|93464-6|LNC|4-Fluorofentanyl|4-Fluorofentanyl
C5211993|T201|COMP|93465-3|LNC|3-Methylfentanyl|3-Methylfentanyl
C5211994|T201|COMP|93466-1|LNC|Valerylfentanyl|Valerylfentanyl
C5211996|T201|COMP|93467-9|LNC|Butyrylfentanyl|Butyrylfentanyl
C5211997|T201|COMP|93468-7|LNC|Acrylfentanyl|Acrylfentanyl
C5211998|T201|COMP|93469-5|LNC|4-Fluorobutyrylfentanyl|4-Fluorobutyrylfentanyl
C5212000|T201|COMP|93470-3|LNC|Furanylfentanyl|Furanylfentanyl
C5212002|T201|COMP|93471-1|LNC|Acetyl norfentanyl|Acetyl norfentanyl
C5212003|T201|COMP|93472-9|LNC|4-Methylphenethylacetylfentanyl|4-Methylphenethylacetylfentanyl
C5212005|T201|COMP|93473-7|LNC|Beta hydroxythiofentanyl|Beta hydroxythiofentanyl
C5212006|T201|COMP|93474-5|LNC|Synthetic opioids panel|Synthetic opioids panel
C5212008|T201|COMP|93475-2|LNC|Busulfan clearance|Busulfan clearance
C5212010|T201|COMP|93476-0|LNC|Busulfan|Busulfan
C5212011|T201|COMP|93477-8|LNC|Busulfan given|Busulfan given
C5212013|T201|COMP|93478-6|LNC|Busulfan area under the curve panel|Busulfan area under the curve panel
C5212017|T201|COMP|93481-0|LNC|Cortisol^10M post 1 ug/kg CRH IV|Cortisol^10M post 1 ug/kg CRH IV
C5212018|T201|COMP|93482-8|LNC|Cortisol^1M pre 1 ug/kg CRH IV|Cortisol^1M pre 1 ug/kg CRH IV
C5212019|T201|COMP|93483-6|LNC|Cortisol^2M post 1 ug/kg CRH IV|Cortisol^2M post 1 ug/kg CRH IV
C5212020|T201|COMP|93484-4|LNC|Cortisol^5M pre 1 ug/kg CRH IV|Cortisol^5M pre 1 ug/kg CRH IV
C5212026|T201|COMP|93488-5|LNC|Guanidinoacetate|Guanidinoacetate
C5212032|T201|COMP|93494-3|LNC|Buprenorphine|Buprenorphine
C5212033|T201|COMP|93495-0|LNC|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine|2-Ethylidene-1,5-Dimethyl-3,3-Diphenylpyrrolidine
C5212034|T201|COMP|93496-8|LNC|Nortriptyline|Nortriptyline
C5212035|T201|COMP|93497-6|LNC|Moxifloxacin 3.0 ug/mL|Moxifloxacin 3.0 ug/mL
C5212037|T201|COMP|93498-4|LNC|Metabotropic glutamate receptor 1 Ab.IgG|Metabotropic glutamate receptor 1 Ab.IgG
C5212039|T201|COMP|93499-2|LNC|Metabotropic glutamate receptor 1 Ab.IgG|Metabotropic glutamate receptor 1 Ab.IgG
C5212040|T201|COMP|93500-7|LNC|Metabotropic glutamate receptor 1 Ab.IgG|Metabotropic glutamate receptor 1 Ab.IgG
C5212041|T201|COMP|93501-5|LNC|Metabotropic glutamate receptor 1 Ab.IgG|Metabotropic glutamate receptor 1 Ab.IgG
C5212042|T201|COMP|93502-3|LNC|N-methyl-D-aspartate receptor subunit 1 Ab.IgG|N-methyl-D-aspartate receptor subunit 1 Ab.IgG
C5212044|T201|COMP|93503-1|LNC|N-methyl-D-aspartate receptor subunit 1 Ab.IgG|N-methyl-D-aspartate receptor subunit 1 Ab.IgG
C5212045|T201|COMP|93504-9|LNC|Cholesterol crystals|Cholesterol crystals
C5212046|T201|COMP|93505-6|LNC|Heptacarboxylporphyrin I|Heptacarboxylporphyrin I
C5212047|T201|COMP|93506-4|LNC|Heptacarboxylporphyrin III|Heptacarboxylporphyrin III
C5212048|T201|COMP|93507-2|LNC|Hexacarboxylporphyrin I|Hexacarboxylporphyrin I
C5212049|T201|COMP|93508-0|LNC|Hexacarboxylporphyrin III|Hexacarboxylporphyrin III
C5212050|T201|COMP|93509-8|LNC|Pentacarboxylporphyrin I|Pentacarboxylporphyrin I
C5212051|T201|COMP|93510-6|LNC|Pentacarboxylporphyrin III|Pentacarboxylporphyrin III
C5212171|T201|COMP|93684-9|LNC|Ammonia|Ammonia
C5212172|T201|COMP|93685-6|LNC|Gas & CO & electrolytes panel|Gas & CO & electrolytes panel
C5212174|T201|COMP|93686-4|LNC|Psychosine|Psychosine
C5212175|T201|COMP|93687-2|LNC|Psychosine|Psychosine
C5212176|T201|COMP|93688-0|LNC|Psychosine|Psychosine
C5212177|T201|COMP|93689-8|LNC|Thrombospondin type I domain-containing 7A Ab.IgG|Thrombospondin type I domain-containing 7A Ab.IgG
C5212178|T201|COMP|93690-6|LNC|BRAF gene.p.Val600 mutations|BRAF gene.p.Val600 mutations
C5212180|T201|COMP|93691-4|LNC|Nonalcoholic steatohepatitis & fibrosis panel|Nonalcoholic steatohepatitis & fibrosis panel
C5212182|T201|COMP|93692-2|LNC|Nonalcoholic steatohepatitis score|Nonalcoholic steatohepatitis score
C5212184|T201|COMP|93693-0|LNC|Nonalcoholic steatohepatitis grade|Nonalcoholic steatohepatitis grade
C5212186|T201|COMP|93694-8|LNC|Nonalcoholic steatohepatitis interpretation|Nonalcoholic steatohepatitis interpretation
C5212188|T201|COMP|93695-5|LNC|Liver steatosis score|Liver steatosis score
C5212190|T201|COMP|93696-3|LNC|Liver steatosis grade|Liver steatosis grade
C5212192|T201|COMP|93697-1|LNC|Liver steatosis interpretation|Liver steatosis interpretation
C5212194|T201|COMP|93698-9|LNC|Gram negative bacterial resistance panel|Gram negative bacterial resistance panel
C5212198|T201|COMP|93700-3|LNC|Bacterial beta-lactam resistance AmpC blaDHA gene|Bacterial beta-lactam resistance AmpC blaDHA gene
C5212200|T201|COMP|93701-1|LNC|Bacterial colistin resistance mcr-2 gene|Bacterial colistin resistance mcr-2 gene
C5212202|T201|COMP|93702-9|LNC|Platelet aggregation.ristocetin induced^15 ug/mL|Platelet aggregation.ristocetin induced^15 ug/mL
C5212206|T201|COMP|93705-2|LNC|Ethyl sulfate & Ethyl glucuronide panel|Ethyl sulfate & Ethyl glucuronide panel
C5212208|T201|COMP|93706-0|LNC|Ethyl sulfate+Ethyl glucuronide|Ethyl sulfate+Ethyl glucuronide
C5212209|T201|COMP|93707-8|LNC|Porphyrin fractions panel|Porphyrin fractions panel
C5212210|T201|COMP|93708-6|LNC|Heptacarboxylporphyrin I/Creatinine|Heptacarboxylporphyrin I/Creatinine
C5212212|T201|COMP|93709-4|LNC|Hexacarboxylporphyrin I/Creatinine|Hexacarboxylporphyrin I/Creatinine
C5212214|T201|COMP|93710-2|LNC|Pentacarboxylporphyrin I/Creatinine|Pentacarboxylporphyrin I/Creatinine
C5212216|T201|COMP|93711-0|LNC|Epstein Barr virus Ab panel|Epstein Barr virus Ab panel
C5212217|T201|COMP|93712-8|LNC|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C5212218|T201|COMP|93713-6|LNC|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C5212219|T201|COMP|93714-4|LNC|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C5212220|T201|COMP|93715-1|LNC|Francisella tularensis Ab.IgG & IgM panel|Francisella tularensis Ab.IgG & IgM panel
C5212222|T201|COMP|93716-9|LNC|Francisella tularensis Ab.IgM|Francisella tularensis Ab.IgM
C5212223|T201|COMP|93717-7|LNC|Francisella tularensis Ab.IgG|Francisella tularensis Ab.IgG
C5212224|T201|COMP|93718-5|LNC|Francisella tularensis Ab.IgG & IgM|Francisella tularensis Ab.IgG & IgM
C5212226|T201|COMP|93719-3|LNC|traMADol|traMADol
C5212227|T201|COMP|93720-1|LNC|traMADol|traMADol
C5212228|T201|COMP|93721-9|LNC|O-Nortramadol|O-Nortramadol
C5212229|T201|COMP|93722-7|LNC|N-Nortramadol|N-Nortramadol
C5212232|T201|COMP|93724-3|LNC|Keratan sulfate|Keratan sulfate
C5212233|T201|COMP|93725-0|LNC|Heparan sulfate|Heparan sulfate
C5212234|T201|COMP|93727-6|LNC|Insulin^post meal|Insulin^post meal
C5212235|T201|COMP|93728-4|LNC|Copper|Copper
C5212236|T201|COMP|93729-2|LNC|Beta-2-Microglobulin/Creatinine|Beta-2-Microglobulin/Creatinine
C5212237|T201|COMP|93730-0|LNC|Testosterone|Testosterone
C5212238|T201|COMP|93731-8|LNC|Androstenedione|Androstenedione
C5212239|T201|COMP|93732-6|LNC|IgE|IgE
C5212240|T201|COMP|93733-4|LNC|Creatinine|Creatinine
C5212241|T201|COMP|93734-2|LNC|Creatinine|Creatinine
C5212242|T201|COMP|93735-9|LNC|Creatinine|Creatinine
C5212243|T201|COMP|93736-7|LNC|Creatinine panel|Creatinine panel
C5212244|T201|COMP|93737-5|LNC|Brassica oleracea var gongylodes Ab.IgE|Brassica oleracea var gongylodes Ab.IgE
C5212246|T201|COMP|93738-3|LNC|Brassica oleracea var botrytis cooked Ab.IgE|Brassica oleracea var botrytis cooked Ab.IgE
C5212248|T201|COMP|93739-1|LNC|Brassica oleracea var capitata f rubra Ab.IgE|Brassica oleracea var capitata f rubra Ab.IgE
C5212250|T201|COMP|93740-9|LNC|Allium schoenoprasum Ab.IgE|Allium schoenoprasum Ab.IgE
C5212252|T201|COMP|93741-7|LNC|Melissa officinalis Ab.IgE|Melissa officinalis Ab.IgE
C5212254|T201|COMP|93742-5|LNC|HTLV I & II Ab band pattern|HTLV I & II Ab band pattern
C5212255|T201|COMP|93743-3|LNC|HTLV I & II Ab.IgG band|HTLV I & II Ab.IgG band
C5212257|T201|COMP|93744-1|LNC|HTLV I & II Ab.IgG panel|HTLV I & II Ab.IgG panel
C5212259|T201|COMP|93745-8|LNC|HTLV I+II Ab.IgG|HTLV I+II Ab.IgG
C5212260|T201|COMP|93746-6|LNC|Protein catabolic rate|Protein catabolic rate
C5212261|T201|COMP|93747-4|LNC|Parainfluenza virus 1+2+3+4 Ab.IgG|Parainfluenza virus 1+2+3+4 Ab.IgG
C5212263|T201|COMP|93748-2|LNC|Fibrin monomer|Fibrin monomer
C5212264|T201|COMP|93749-0|LNC|Mumps virus N gene|Mumps virus N gene
C5212266|T201|COMP|93750-8|LNC|Mumps virus RNA & N gene panel|Mumps virus RNA & N gene panel
C5212268|T201|COMP|93751-6|LNC|Atypical porcine pestivirus RNA|Atypical porcine pestivirus RNA
C5212270|T201|COMP|93752-4|LNC|Atypical porcine pestivirus RNA|Atypical porcine pestivirus RNA
C5212271|T201|COMP|93753-2|LNC|Porcine cytomegalovirus DNA|Porcine cytomegalovirus DNA
C5212272|T201|COMP|93754-0|LNC|Encephalomyocarditis virus RNA|Encephalomyocarditis virus RNA
C5212273|T201|COMP|93755-7|LNC|Porcine circovirus type 3 DNA|Porcine circovirus type 3 DNA
C5212274|T201|COMP|93756-5|LNC|Mycoplasma hyorhinis Ab.IgG/Positive control|Mycoplasma hyorhinis Ab.IgG/Positive control
C5212278|T201|COMP|93758-1|LNC|Erysipelothrix sp|Erysipelothrix sp
C5212279|T201|COMP|93759-9|LNC|Influenza virus A PB2 gene|Influenza virus A PB2 gene
C5212281|T201|COMP|93760-7|LNC|Influenza virus A PB1 gene|Influenza virus A PB1 gene
C5212283|T201|COMP|93761-5|LNC|Influenza virus A PA gene|Influenza virus A PA gene
C5212285|T201|COMP|93762-3|LNC|Influenza virus A NP gene|Influenza virus A NP gene
C5212287|T201|COMP|93763-1|LNC|Influenza virus A NS1 gene|Influenza virus A NS1 gene
C5212289|T201|COMP|93764-9|LNC|Porcine astrovirus type 3 RNA|Porcine astrovirus type 3 RNA
C5212291|T201|COMP|93765-6|LNC|Trimethylamine N-oxide|Trimethylamine N-oxide
C5212292|T201|COMP|93766-4|LNC|Cryptococcus sp Ag|Cryptococcus sp Ag
C5212293|T201|COMP|93767-2|LNC|Eravacycline|Eravacycline
C5212294|T201|COMP|93768-0|LNC|Acarboxyprothrombin|Acarboxyprothrombin
C5212295|T201|COMP|93769-8|LNC|Choriogonadotropin.intact+Beta subunit|Choriogonadotropin.intact+Beta subunit
C5212296|T201|COMP|93770-6|LNC|Ceramide trihexoside|Ceramide trihexoside
C5212297|T201|COMP|93771-4|LNC|Calprotectin|Calprotectin
C5212298|T201|COMP|93772-2|LNC|4-hydroxyglutamate/Creatinine|4-hydroxyglutamate/Creatinine
C5212300|T201|COMP|93773-0|LNC|11-Deoxycortisol|11-Deoxycortisol
C5212301|T201|COMP|93774-8|LNC|Trans-cinnamoylglycine/Creatinine|Trans-cinnamoylglycine/Creatinine
C5212302|T201|COMP|93775-5|LNC|2-Octenoate/Creatinine|2-Octenoate/Creatinine
C5212304|T201|COMP|93776-3|LNC|Babesia duncani Ab.IgG|Babesia duncani Ab.IgG
C5212306|T201|COMP|93777-1|LNC|Human papilloma virus 16+18 E6+E7 mRNA|Human papilloma virus 16+18 E6+E7 mRNA
C5212308|T201|COMP|93778-9|LNC|Human papilloma virus 6+11 E6+E7 mRNA|Human papilloma virus 6+11 E6+E7 mRNA
C5212310|T201|COMP|93779-7|LNC|Large B-cell lymphoma and cell of origin|Large B-cell lymphoma and cell of origin
C5212312|T201|COMP|93780-5|LNC|Primary mediastinal large B-cell lymphoma|Primary mediastinal large B-cell lymphoma
C5212314|T201|COMP|93782-1|LNC|Large B-cell lymphoma|Large B-cell lymphoma
C5212316|T201|COMP|93783-9|LNC|Diffuse large B-cell lymphoma cell of origin|Diffuse large B-cell lymphoma cell of origin
C5212320|T201|COMP|93785-4|LNC|Large B-cell lymphoma classification panel|Large B-cell lymphoma classification panel
C5212322|T201|COMP|93786-2|LNC|Varicella zoster virus Ab.IgM+total|Varicella zoster virus Ab.IgM+total
C5212324|T201|COMP|93787-0|LNC|Lymphocytic choriomeningitis virus Ab.IgG+IgM|Lymphocytic choriomeningitis virus Ab.IgG+IgM
C5212325|T201|COMP|93788-8|LNC|F5 gene HR2 haplotype|F5 gene HR2 haplotype
C5212327|T201|COMP|93789-6|LNC|Time to microorganism growth detection|Time to microorganism growth detection
C5212329|T201|COMP|93790-4|LNC|Delafloxacin|Delafloxacin
C5212330|T201|COMP|93791-2|LNC|Glucose|Glucose
C5212331|T201|COMP|93792-0|LNC|Insulin sensitivity index|Insulin sensitivity index
C5212333|T201|COMP|93793-8|LNC|Insulin|Insulin
C5212334|T201|COMP|93794-6|LNC|Glucose tolerance & insulin sensitivity 2H panel|Glucose tolerance & insulin sensitivity 2H panel
C5212336|T201|COMP|93795-3|LNC|NOP56 gene.GGCCTG repeats|NOP56 gene.GGCCTG repeats
C5212338|T201|COMP|93796-1|LNC|MYCN gene amplification|MYCN gene amplification
C5212339|T201|COMP|93797-9|LNC|MYCN gene copy number/Chromosome 2 copy number|MYCN gene copy number/Chromosome 2 copy number
C5212341|T201|COMP|93798-7|LNC|MYCN gene copy number/nucleus|MYCN gene copy number/nucleus
C5212343|T201|COMP|93799-5|LNC|Chromosome 2 copy number/nucleus|Chromosome 2 copy number/nucleus
C5212345|T201|COMP|93800-1|LNC|1p chromosome deletion/1q chromosome deletion|1p chromosome deletion/1q chromosome deletion
C5212347|T201|COMP|93801-9|LNC|Chromosome 1 polysomy|Chromosome 1 polysomy
C5212349|T201|COMP|93802-7|LNC|19q chromosome deletion/19p chromosome deletion|19q chromosome deletion/19p chromosome deletion
C5212351|T201|COMP|93803-5|LNC|Chromosome 19 polysomy|Chromosome 19 polysomy
C5212353|T201|COMP|93804-3|LNC|Chromosome 12 copy number/nucleus|Chromosome 12 copy number/nucleus
C5212355|T201|COMP|93805-0|LNC|MDM2 gene copy number/nucleus|MDM2 gene copy number/nucleus
C5212357|T201|COMP|93806-8|LNC|EWSR1 gene rearrangements|EWSR1 gene rearrangements
C5212359|T201|COMP|93807-6|LNC|FOXO1 gene rearrangements|FOXO1 gene rearrangements
C5212361|T201|COMP|93808-4|LNC|MDM2 gene amplification|MDM2 gene amplification
C5212362|T201|COMP|93809-2|LNC|MDM2 gene copy number/Chromosome 12 copy number|MDM2 gene copy number/Chromosome 12 copy number
C5212364|T201|COMP|93810-0|LNC|SS18 gene rearrangements|SS18 gene rearrangements
C5212366|T201|COMP|93811-8|LNC|F9 gene full mutation analysis|F9 gene full mutation analysis
C5212368|T201|COMP|93812-6|LNC|1,3 beta glucan|1,3 beta glucan
C5212371|T201|COMP|93814-2|LNC|SERPINC1 gene full mutation analysis|SERPINC1 gene full mutation analysis
C5212373|T201|COMP|93815-9|LNC|PROC gene full mutation analysis|PROC gene full mutation analysis
C5212391|T201|COMP|93834-0|LNC|Coccidioides sp Ab.IgM|Coccidioides sp Ab.IgM
C5212392|T201|COMP|93835-7|LNC|Coccidioides sp Ab.IgM|Coccidioides sp Ab.IgM
C5212393|T201|COMP|93836-5|LNC|Coccidioides sp Ab.IgG|Coccidioides sp Ab.IgG
C5212394|T201|COMP|93837-3|LNC|Coccidioides sp Ab.IgG|Coccidioides sp Ab.IgG
C5212395|T201|COMP|93838-1|LNC|Histoplasma capsulatum Ab.IgM|Histoplasma capsulatum Ab.IgM
C5212396|T201|COMP|93839-9|LNC|Histoplasma capsulatum Ab.IgG|Histoplasma capsulatum Ab.IgG
C5212397|T201|COMP|93840-7|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C5212398|T201|COMP|93841-5|LNC|Epstein Barr virus DNA|Epstein Barr virus DNA
C5212399|T201|COMP|93842-3|LNC|HOGA1 gene full mutation analysis|HOGA1 gene full mutation analysis
C5212401|T201|COMP|93843-1|LNC|Primary hyperoxaluria multigene analysis|Primary hyperoxaluria multigene analysis
C5212403|T201|COMP|93844-9|LNC|UGT1A1 gene full mutation analysis|UGT1A1 gene full mutation analysis
C5212405|T201|COMP|93845-6|LNC|UGT1A1 gene.TA repeats & c.211G>A|UGT1A1 gene.TA repeats & c.211G>A
C5212407|T201|COMP|93846-4|LNC|Hemoglobin|Hemoglobin
C5212408|T201|COMP|93847-2|LNC|Aspergillus oryzae Ab.IgE|Aspergillus oryzae Ab.IgE
C5212411|T201|COMP|93850-6|LNC|Pretomanid|Pretomanid
C5212412|T201|COMP|93851-4|LNC|Delamanid|Delamanid
C5212415|T201|COMP|93853-0|LNC|N-Acetylgalactosamine-6-Sulfatase|N-Acetylgalactosamine-6-Sulfatase
C5212416|T201|COMP|93854-8|LNC|Gadolinium/Creatinine|Gadolinium/Creatinine
C5212418|T201|COMP|93855-5|LNC|Iothalamate|Iothalamate
C5212419|T201|COMP|93856-3|LNC|Enterovirus RNA|Enterovirus RNA
C5212420|T201|COMP|93858-9|LNC|Toxoplasma gondii Ab.IgG panel|Toxoplasma gondii Ab.IgG panel
C5212422|T201|COMP|93859-7|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C5212423|T201|COMP|93860-5|LNC|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C5212430|T201|COMP|93866-2|LNC|C4 nephritic factor|C4 nephritic factor
C5212431|T201|COMP|93867-0|LNC|Gamma aminobutyrate B receptor Ab|Gamma aminobutyrate B receptor Ab
C5212434|T201|COMP|93870-4|LNC|N-methyl-D-aspartate receptor subunit 1 Ab|N-methyl-D-aspartate receptor subunit 1 Ab
C5212435|T201|COMP|93871-2|LNC|Borrelia miyamotoi Ab.IgG+IgM|Borrelia miyamotoi Ab.IgG+IgM
C5212437|T201|COMP|93872-0|LNC|Tamoxifen metabolites pattern|Tamoxifen metabolites pattern
C5212439|T201|COMP|93873-8|LNC|Borrelia miyamotoi Ab.IgG|Borrelia miyamotoi Ab.IgG
C5212441|T201|COMP|93874-6|LNC|Borrelia miyamotoi Ab.IgM|Borrelia miyamotoi Ab.IgM
C5212443|T201|COMP|93875-3|LNC|Phosphohistone H3|Phosphohistone H3
C5212445|T201|COMP|93876-1|LNC|Ceramide risk score|Ceramide risk score
C5212447|T201|COMP|93877-9|LNC|N-Nervonoylsphingosine/N-Lignoceroylsphingosine|N-Nervonoylsphingosine/N-Lignoceroylsphingosine
C5212449|T201|COMP|93878-7|LNC|N-Stearoylsphingosine/N-Lignoceroylsphingosine|N-Stearoylsphingosine/N-Lignoceroylsphingosine
C5212451|T201|COMP|93879-5|LNC|N-Palmitoylsphingosine/N-Lignoceroylsphingosine|N-Palmitoylsphingosine/N-Lignoceroylsphingosine
C5212453|T201|COMP|93880-3|LNC|N-Nervonoylsphingosine|N-Nervonoylsphingosine
C5212455|T201|COMP|93881-1|LNC|N-Stearoylsphingosine|N-Stearoylsphingosine
C5212457|T201|COMP|93882-9|LNC|N-Palmitoylsphingosine|N-Palmitoylsphingosine
C5212458|T201|COMP|93883-7|LNC|Ceramide panel|Ceramide panel
C5212460|T201|COMP|93884-5|LNC|Methane/Expired gas^2H post dose carbohydrate|Methane/Expired gas^2H post dose carbohydrate
C5212461|T201|COMP|93885-2|LNC|Methane/Expired gas^1.5H post dose carbohydrate|Methane/Expired gas^1.5H post dose carbohydrate
C5212462|T201|COMP|93886-0|LNC|Methane/Expired gas^1H post dose carbohydrate|Methane/Expired gas^1H post dose carbohydrate
C5212463|T201|COMP|93887-8|LNC|Methane/Expired gas^45M post dose carbohydrate|Methane/Expired gas^45M post dose carbohydrate
C5212464|T201|COMP|93888-6|LNC|Methane/Expired gas^30M post dose carbohydrate|Methane/Expired gas^30M post dose carbohydrate
C5212465|T201|COMP|93889-4|LNC|Methane/Expired gas^15M post dose carbohydrate|Methane/Expired gas^15M post dose carbohydrate
C5212466|T201|COMP|93890-2|LNC|Methane/Expired gas^pre dose carbohydrate|Methane/Expired gas^pre dose carbohydrate
C5212467|T201|COMP|93891-0|LNC|Methane/Expired gas^post dose carbohydrate|Methane/Expired gas^post dose carbohydrate
C5212480|T201|COMP|93905-8|LNC|ABO group^during infancy|ABO group^during infancy
C5212481|T201|COMP|93906-6|LNC|ABO & Rh group^during infancy|ABO & Rh group^during infancy
C5212482|T201|COMP|93907-4|LNC|L little u 20 Ag|L little u 20 Ag
C5212484|T201|COMP|93908-2|LNC|A little u super little b Ag|A little u super little b Ag
C5212486|T201|COMP|93909-0|LNC|J little k3 Ag|J little k3 Ag
C5212488|T201|COMP|93910-8|LNC|F little y3 Ag|F little y3 Ag
C5212490|T201|COMP|93911-6|LNC|little c E Ag|little c E Ag
C5212492|T201|COMP|93913-2|LNC|VS Ag|VS Ag
C5212493|T201|COMP|93914-0|LNC|Blood group antigens panel|Blood group antigens panel
C5212495|T201|COMP|93915-7|LNC|Rh antigens & K Ag panel|Rh antigens & K Ag panel
C5212497|T201|COMP|93916-5|LNC|ABO & Rh group panel|ABO & Rh group panel
C5212498|T201|COMP|93917-3|LNC|K Ag^post transfusion reaction|K Ag^post transfusion reaction
C5212501|T201|COMP|93923-1|LNC|ABO & Rh group post transfusion reaction panel|ABO & Rh group post transfusion reaction panel
C5212503|T201|COMP|93924-9|LNC|K Ag^post hematopoietic stem cell transplant|K Ag^post hematopoietic stem cell transplant
C5212506|T201|COMP|93930-6|LNC|D Ag^post hematopoietic stem cell transplant|D Ag^post hematopoietic stem cell transplant
C5212507|T201|COMP|93931-4|LNC|ABO group^post hematopoietic stem cell transplant|ABO group^post hematopoietic stem cell transplant
C5212511|T201|COMP|93934-8|LNC|K Ag^during infancy|K Ag^during infancy
C5212512|T201|COMP|93939-7|LNC|Rh antigens & K Ag during infancy panel|Rh antigens & K Ag during infancy panel
C5212514|T201|COMP|93940-5|LNC|D Ag^during infancy|D Ag^during infancy
C5212515|T201|COMP|93941-3|LNC|ABO & Rh group during infancy panel|ABO & Rh group during infancy panel
C5212517|T201|COMP|93942-1|LNC|K Ag|K Ag
C5212518|T201|COMP|93947-0|LNC|Rh antigens & K Ag panel|Rh antigens & K Ag panel
C5212519|T201|COMP|93948-8|LNC|D Ag|D Ag
C5212520|T201|COMP|93949-6|LNC|ABO & Rh group panel|ABO & Rh group panel
C5212521|T201|COMP|93950-4|LNC|D variant Ag|D variant Ag
C5212523|T201|COMP|93951-2|LNC|Rh antigens & K Ag panel|Rh antigens & K Ag panel
C5212524|T201|COMP|93952-0|LNC|Metamyelocytes.neutrophilic/100 leukocytes|Metamyelocytes.neutrophilic/100 leukocytes
C5212525|T201|COMP|93953-8|LNC|Lymphocytes.villous|Lymphocytes.villous
C5212545|T201|COMP|93972-8|LNC|Acetaminophen-cysteine adduct|Acetaminophen-cysteine adduct
C5212547|T201|COMP|93973-6|LNC|Iohexol|Iohexol
C5212548|T201|COMP|93974-4|LNC|Iohexol|Iohexol
C5212549|T201|COMP|93975-1|LNC|Urea nitrogen^1H specimen|Urea nitrogen^1H specimen
C5212550|T201|COMP|93976-9|LNC|Chikungunya virus Ab.IgM & IgG panel|Chikungunya virus Ab.IgM & IgG panel
C5212552|T201|COMP|93977-7|LNC|Complement C2.functional|Complement C2.functional
C5212554|T201|COMP|93978-5|LNC|Complement C4.functional|Complement C4.functional
C5212556|T201|COMP|93979-3|LNC|Chikungunya virus Ab.IgG|Chikungunya virus Ab.IgG
C5212557|T201|COMP|93980-1|LNC|Iothalamate|Iothalamate
C5212558|T201|COMP|93981-9|LNC|Hydrogen/Expired gas^2H post dose carbohydrate|Hydrogen/Expired gas^2H post dose carbohydrate
C5212559|T201|COMP|93982-7|LNC|Hydrogen/Expired gas^1.5H post dose carbohydrate|Hydrogen/Expired gas^1.5H post dose carbohydrate
C5212560|T201|COMP|93983-5|LNC|Hydrogen/Expired gas^1H post dose carbohydrate|Hydrogen/Expired gas^1H post dose carbohydrate
C5212561|T201|COMP|93984-3|LNC|Hydrogen/Expired gas^45M post dose carbohydrate|Hydrogen/Expired gas^45M post dose carbohydrate
C5212562|T201|COMP|93985-0|LNC|Hydrogen/Expired gas^30M post dose carbohydrate|Hydrogen/Expired gas^30M post dose carbohydrate
C5212563|T201|COMP|93986-8|LNC|Hydrogen/Expired gas^15M post dose carbohydrate|Hydrogen/Expired gas^15M post dose carbohydrate
C5212564|T201|COMP|93987-6|LNC|Hydrogen/Expired gas^pre dose carbohydrate|Hydrogen/Expired gas^pre dose carbohydrate
C5212565|T201|COMP|93988-4|LNC|Hydrogen/Expired gas^post dose carbohydrate|Hydrogen/Expired gas^post dose carbohydrate
C5212566|T201|COMP|93989-2|LNC|Carbohydrate challenge panel|Carbohydrate challenge panel
C5212568|T201|COMP|93990-0|LNC|Osmolality^post 1H FFst|Osmolality^post 1H FFst
C5212569|T201|COMP|93991-8|LNC|Osmolality^post 2H FFst|Osmolality^post 2H FFst
C5212570|T201|COMP|93992-6|LNC|Osmolality^post 3H FFst|Osmolality^post 3H FFst
C5212571|T201|COMP|93993-4|LNC|Osmolality^post 4H FFst|Osmolality^post 4H FFst
C5212572|T201|COMP|93994-2|LNC|Osmolality^post 5H FFst|Osmolality^post 5H FFst
C5212573|T201|COMP|93995-9|LNC|Osmolality^post 6H FFst|Osmolality^post 6H FFst
C5212574|T201|COMP|93996-7|LNC|Osmolality^post 7H FFst|Osmolality^post 7H FFst
C5212575|T201|COMP|93997-5|LNC|Sodium^1H post dose vasopressin|Sodium^1H post dose vasopressin
C5212576|T201|COMP|93998-3|LNC|Potassium^1H post dose vasopressin|Potassium^1H post dose vasopressin
C5212577|T201|COMP|93999-1|LNC|Creatinine^1H post dose vasopressin|Creatinine^1H post dose vasopressin
C5212578|T201|COMP|94000-7|LNC|Chloride^1H post dose vasopressin|Chloride^1H post dose vasopressin
C5212579|T201|COMP|94001-5|LNC|Bicarbonate^1H post dose vasopressin|Bicarbonate^1H post dose vasopressin
C5212580|T201|COMP|94002-3|LNC|Anion Gap 3^1H post dose vasopressin|Anion Gap 3^1H post dose vasopressin
C5212581|T201|COMP|94003-1|LNC|Urea nitrogen^1H post dose vasopressin|Urea nitrogen^1H post dose vasopressin
C5212582|T201|COMP|94004-9|LNC|Osmolality^1H post dose vasopressin|Osmolality^1H post dose vasopressin
C5212583|T201|COMP|94005-6|LNC|Osmolality^1H post dose vasopressin|Osmolality^1H post dose vasopressin
C5212584|T201|COMP|94006-4|LNC|Sodium^2H post dose vasopressin|Sodium^2H post dose vasopressin
C5212585|T201|COMP|94007-2|LNC|Potassium^2H post dose vasopressin|Potassium^2H post dose vasopressin
C5212586|T201|COMP|94008-0|LNC|Creatinine^2H post dose vasopressin|Creatinine^2H post dose vasopressin
C5212587|T201|COMP|94009-8|LNC|Chloride^2H post dose vasopressin|Chloride^2H post dose vasopressin
C5212588|T201|COMP|94010-6|LNC|Bicarbonate^2H post dose vasopressin|Bicarbonate^2H post dose vasopressin
C5212589|T201|COMP|94011-4|LNC|Anion Gap 3^2H post dose vasopressin|Anion Gap 3^2H post dose vasopressin
C5212590|T201|COMP|94012-2|LNC|Urea nitrogen^2H post dose vasopressin|Urea nitrogen^2H post dose vasopressin
C5212591|T201|COMP|94013-0|LNC|Osmolality^2H post dose vasopressin|Osmolality^2H post dose vasopressin
C5212592|T201|COMP|94014-8|LNC|Osmolality^2H post dose vasopressin|Osmolality^2H post dose vasopressin
C5212593|T201|COMP|94040-3|LNC|Adenovirus A+B+C+D+E DNA|Adenovirus A+B+C+D+E DNA
C5212620|T201|COMP|94054-4|LNC|Bacterial katG gene drug resistance mutation|Bacterial katG gene drug resistance mutation
C5212622|T201|COMP|94055-1|LNC|Bacterial inhA gene drug resistance mutation|Bacterial inhA gene drug resistance mutation
C5212624|T201|COMP|94056-9|LNC|Bacterial fabG1 gene drug resistance mutation|Bacterial fabG1 gene drug resistance mutation
C5212626|T201|COMP|94057-7|LNC|Bacterial ahpC gene drug resistance mutation|Bacterial ahpC gene drug resistance mutation
C5212628|T201|COMP|94058-5|LNC|Bacterial embB gene drug resistance mutation|Bacterial embB gene drug resistance mutation
C5212630|T201|COMP|94059-3|LNC|Bacterial pncA gene drug resistance mutation|Bacterial pncA gene drug resistance mutation
C5212632|T201|COMP|94060-1|LNC|Bacterial gyrA gene drug resistance mutation|Bacterial gyrA gene drug resistance mutation
C5212634|T201|COMP|94061-9|LNC|Bacterial gidB gene drug resistance mutation|Bacterial gidB gene drug resistance mutation
C5212636|T201|COMP|94062-7|LNC|Bacterial rrs gene drug resistance mutation|Bacterial rrs gene drug resistance mutation
C5212638|T201|COMP|94063-5|LNC|Bacterial rpsL gene drug resistance mutation|Bacterial rpsL gene drug resistance mutation
C5212640|T201|COMP|94064-3|LNC|Bacterial eis gene drug resistance mutation|Bacterial eis gene drug resistance mutation
C5212642|T201|COMP|94065-0|LNC|Bacterial rpoB gene drug resistance mutation|Bacterial rpoB gene drug resistance mutation
C5212650|T201|COMP|94076-7|LNC|Mutations/Megabase|Mutations/Megabase
C5212652|T201|COMP|94077-5|LNC|Tumor mutation burden|Tumor mutation burden
C5212653|T201|COMP|94078-3|LNC|PDX1 gene full mutation analysis|PDX1 gene full mutation analysis
C5212655|T201|COMP|94079-1|LNC|TYMP gene full mutation analysis|TYMP gene full mutation analysis
C5212657|T201|COMP|94080-9|LNC|RRM2B gene full mutation analysis|RRM2B gene full mutation analysis
C5212663|T201|COMP|94087-4|LNC|Chromosome analysis|Chromosome analysis
C5212674|T201|COMP|94096-5|LNC|Collagen type VII Ab.IgG|Collagen type VII Ab.IgG
C5212676|T201|COMP|94097-3|LNC|Cytosolic 5'-nucleotidase 1A Ab.IgG|Cytosolic 5'-nucleotidase 1A Ab.IgG
C5212678|T201|COMP|94098-1|LNC|Dense fine speckled 70 protein Ab.IgG|Dense fine speckled 70 protein Ab.IgG
C5212679|T201|COMP|94099-9|LNC|Hantavirus Ab.IgM|Hantavirus Ab.IgM
C5212680|T201|COMP|94100-5|LNC|Hantavirus seoul Ab.IgM|Hantavirus seoul Ab.IgM
C5212682|T201|COMP|94101-3|LNC|Hantavirus seoul Ab.IgG|Hantavirus seoul Ab.IgG
C5212683|T201|COMP|94102-1|LNC|Epstein Barr virus early diffuse Ab.IgA|Epstein Barr virus early diffuse Ab.IgA
C5212685|T201|COMP|94103-9|LNC|Zolpidem phenyl-4-carboxylate|Zolpidem phenyl-4-carboxylate
C5212686|T201|COMP|94104-7|LNC|Zolpidem|Zolpidem
C5212687|T201|COMP|94105-4|LNC|Alpha hydroxytriazolam|Alpha hydroxytriazolam
C5212688|T201|COMP|94106-2|LNC|Temazepam glucuronide|Temazepam glucuronide
C5212689|T201|COMP|94107-0|LNC|Oxazepam glucuronide|Oxazepam glucuronide
C5212690|T201|COMP|94108-8|LNC|1-Hydroxymidazolam|1-Hydroxymidazolam
C5212691|T201|COMP|94109-6|LNC|LORazepam glucuronide|LORazepam glucuronide
C5212692|T201|COMP|94110-4|LNC|2-Hydroxyethylflurazepam|2-Hydroxyethylflurazepam
C5212694|T201|COMP|94111-2|LNC|7-Aminoflunitrazepam|7-Aminoflunitrazepam
C5212695|T201|COMP|94112-0|LNC|7-Aminoclonazepam|7-Aminoclonazepam
C5212696|T201|COMP|94113-8|LNC|Norclobazam|Norclobazam
C5212697|T201|COMP|94114-6|LNC|cloBAZam|cloBAZam
C5212698|T201|COMP|94115-3|LNC|Alpha hydroxyalprazolam glucuronide|Alpha hydroxyalprazolam glucuronide
C5212700|T201|COMP|94116-1|LNC|ALPRAZolam|ALPRAZolam
C5212701|T201|COMP|94117-9|LNC|Benzodiazepines panel|Benzodiazepines panel
C5212714|T201|COMP|94127-8|LNC|Clarity|Clarity
C5212717|T201|COMP|94129-4|LNC|Water deprivation challenge panel|Water deprivation challenge panel
C1624104|T201|COMP|41995-2|LNC|HbA1c|HbA1c
C1624104|T201|COMP|41995-2|LNC|A1c|A1c
C1624104|T201|COMP|41995-2|LNC|A1c|A1c
