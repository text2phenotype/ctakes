// CUI|TUI|CODE|VOCAB|TXT|PREF TEXT
C000002|T109|2|DICT2|Drug|Drug annotation from dict 2
C000004|T060|4|DICT2|Proc|Procedure annotation from dict 2