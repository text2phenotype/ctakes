C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C1306838|T047|224729007|SNOMEDCT_US|PROLIFERATIVE ARTHRITIS|PROLIFERATIVE ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0157913|T047|267887009|SNOMEDCT_US|RHEUMATOID ARTHRITIS AND OTHER INFLAMMATORY POLYARTHROPATHIES|RHEUMATOID ARTHRITIS AND OTHER INFLAMMATORY POLYARTHROPATHIES (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTYS SYNDROME|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTYS SYNDROME, UNSPECIFIED SITE|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH SPLENOADENOMEGALY AND LEUKOPENIA|FELTY'S SYNDROME (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHIES|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHIES (M05-M14)|POLYARTHRITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|RHEUMATOID VASCULITIS|RHEUMATOID VASCULITIS (DISORDER)
C0264747|T047|28381002|SNOMEDCT_US|RHEUMATOID PERICARDITIS|RHEUMATIC PERICARDITIS (DISORDER)
C0392469|T047|28880005|SNOMEDCT_US|RHEUMATOID CARDITIS|RHEUMATOID CARDITIS (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|SEROPOSITIVE RHEUMATOID ARTHRITIS|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0477541|T047|203730003|SNOMEDCT_US|OTHER SEROPOSITIVE RHEUMATOID ARTHRITIS|[X]OTHER SEROPOSITIVE RHEUMATOID ARTHRITIS (DISORDER)
C0489959|T047|195136004|SNOMEDCT_US|RHEUMATOID MYOCARDITIS|RHEUMATOID MYOCARDITIS (DISORDER)
C0494896|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0837507|T047||SNOMEDCT_US|FELTYS SYNDROME, MULTIPLE SITES
C0837511|T047||SNOMEDCT_US|FELTYS SYNDROME, HAND
C0837511|T047||SNOMEDCT_US|FELTYS SYNDROME, UNSPECIFIED HAND
C0837514|T047||SNOMEDCT_US|FELTYS SYNDROME, ANKLE AND FOOT
C0837537|T047||SNOMEDCT_US|RHEU ARTHRITIS MULT SITE W INVOLV OF ORGANS AND SYSTEMS
C0837537|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF MULTIPLE SITES WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0837541|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0837544|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0837546|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP SITE W INVOLV OF ORGANS AND SYSTEMS
C0837546|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0994344|T047|155621007|SNOMEDCT_US|RHEUMATOID LUNG DISEASE|RHEUMATOID LUNG (DISORDER)
C2889108|T047||SNOMEDCT_US|FELTYS SYNDROME, RIGHT SHOULDER
C2889109|T047||SNOMEDCT_US|FELTYS SYNDROME, LEFT SHOULDER
C2889110|T047||SNOMEDCT_US|FELTYS SYNDROME, UNSPECIFIED SHOULDER
C2889112|T047||SNOMEDCT_US|FELTYS SYNDROME, RIGHT ELBOW
C2889113|T047||SNOMEDCT_US|FELTYS SYNDROME, LEFT ELBOW
C2889114|T047||SNOMEDCT_US|FELTYS SYNDROME, CARPAL BONES
C2889116|T047||SNOMEDCT_US|FELTYS SYNDROME, RIGHT WRIST
C2889117|T047||SNOMEDCT_US|FELTYS SYNDROME, LEFT WRIST
C2889118|T047||SNOMEDCT_US|FELTYS SYNDROME, UNSPECIFIED WRIST
C2889119|T047||SNOMEDCT_US|FELTYS SYNDROME, METACARPUS AND PHALANGES
C2889120|T047||SNOMEDCT_US|FELTYS SYNDROME, RIGHT HAND
C2889121|T047||SNOMEDCT_US|FELTYS SYNDROME, LEFT HAND
C2889122|T047||SNOMEDCT_US|FELTYS SYNDROME, RIGHT HIP
C2889123|T047||SNOMEDCT_US|FELTYS SYNDROME, LEFT HIP
C2889126|T047||SNOMEDCT_US|FELTYS SYNDROME, RIGHT KNEE
C2889127|T047||SNOMEDCT_US|FELTYS SYNDROME, LEFT KNEE
C2889128|T047||SNOMEDCT_US|FELTYS SYNDROME, TARSUS, METATARSUS AND PHALANGES
C2889129|T047||SNOMEDCT_US|FELTYS SYNDROME, RIGHT ANKLE AND FOOT
C2889130|T047||SNOMEDCT_US|FELTYS SYNDROME, LEFT ANKLE AND FOOT
C2889131|T047||SNOMEDCT_US|FELTYS SYNDROME, UNSPECIFIED ANKLE AND FOOT
C2889132|T047|319841000119107|SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS (DISORDER)
C2889133|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP SITE
C2889133|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889134|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889135|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889135|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889136|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889136|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889137|T047||SNOMEDCT_US|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889137|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889138|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889139|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF R ELBOW
C2889139|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889140|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889140|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889141|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889141|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889142|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS, CARPAL BONES
C2889143|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF WRIST
C2889144|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF R WRIST
C2889144|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889145|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889145|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889146|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889146|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889147|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS, METACARPUS AND PHALANGES
C2889148|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF HAND
C2889149|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889149|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889150|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT HAND
C2889150|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889151|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP HAND
C2889151|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889152|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP HIP
C2889152|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF HIP
C2889152|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889153|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889153|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889154|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT HIP
C2889154|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889155|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF KNEE
C2889156|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889156|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889157|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889157|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889158|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889158|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889159|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS, TARSUS, METATARSUS AND PHALANGES
C2889160|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889161|T047||SNOMEDCT_US|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889161|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889162|T047||SNOMEDCT_US|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889162|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889163|T047||SNOMEDCT_US|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889163|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889164|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS MULT SITE
C2889164|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889165|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS
C2889165|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP SITE
C2889165|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889166|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889166|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889167|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889167|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889168|T047||SNOMEDCT_US|RHEU VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889168|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889168|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889169|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889170|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889170|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889171|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889171|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889172|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889172|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889173|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS, CARPAL BONES
C2889174|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF WRIST
C2889175|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889175|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889176|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889176|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889177|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889177|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889178|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS, METACARPUS AND PHALANGES
C2889179|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF HAND
C2889179|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP HAND
C2889179|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889180|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889180|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889181|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889182|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF HIP
C2889183|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889184|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889185|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP HIP
C2889185|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889186|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF KNEE
C2889187|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889187|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889188|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889189|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889189|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889190|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS, TARSUS, METATARSUS AND PHALANGES
C2889191|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889192|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889192|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889193|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889193|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889194|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889194|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889195|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS MULT SITE
C2889195|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889196|T047||SNOMEDCT_US|RHEUMATOID ENDOCARDITIS
C2889197|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS
C2889198|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP SITE
C2889198|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889199|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889200|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889200|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889201|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889201|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889202|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889202|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889203|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889204|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF R ELBOW
C2889204|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889205|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF L ELBOW
C2889205|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889206|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889206|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889207|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS, CARPAL BONES
C2889208|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF WRIST
C2889209|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF R WRIST
C2889209|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889210|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF L WRIST
C2889210|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889211|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889211|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889212|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS, METACARPUS AND PHALANGES
C2889213|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF HAND
C2889214|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889214|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889215|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT HAND
C2889215|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889216|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP HAND
C2889216|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889217|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP HIP
C2889217|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF HIP
C2889217|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889218|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889218|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889219|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT HIP
C2889219|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889220|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF KNEE
C2889221|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889221|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889222|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889222|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889223|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889223|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889224|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS, TARSUS, METATARSUS AND PHALANGES
C2889225|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889226|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889226|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889227|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889227|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889228|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889228|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889229|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS MULT SITE
C2889229|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889230|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS
C2889231|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP SITE
C2889231|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889232|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889233|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889233|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889234|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889234|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889235|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889235|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889236|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889237|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889238|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889239|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889239|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889240|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS, CARPAL BONES
C2889241|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF WRIST
C2889242|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889243|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889244|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889244|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889245|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS, METACARPUS AND PHALANGES
C2889246|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF HAND
C2889246|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP HAND
C2889246|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889247|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889248|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889249|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF HIP
C2889250|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889251|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889252|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP HIP
C2889252|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889253|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF KNEE
C2889254|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889255|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889256|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889256|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889257|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS, TARSUS, METATARSUS AND PHALANGES
C2889258|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889259|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889259|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889260|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889260|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889261|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889261|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889262|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889262|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889263|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS
C2889264|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP SITE
C2889264|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889265|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889266|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889266|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889267|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889267|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889268|T047||SNOMEDCT_US|RHEU POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889268|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889269|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889269|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889270|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889270|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889271|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889271|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889271|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889272|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS, CARPAL BONES
C2889273|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF WRIST
C2889274|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889274|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889275|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889275|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889276|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889276|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889277|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS, METACARPUS AND PHALANGES
C2889278|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF HAND
C2889279|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889279|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889280|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT HAND
C2889280|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889281|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP HAND
C2889281|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889282|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF HIP
C2889283|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889283|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889284|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY W RHEUMATOID ARTHRITIS OF LEFT HIP
C2889284|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889285|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY W RHEUMATOID ARTHRITIS OF UNSP HIP
C2889285|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889286|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF KNEE
C2889287|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889287|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889288|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889288|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889289|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889289|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889290|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS, TARSUS, METATARSUS AND PHALANGES
C2889291|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889292|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889292|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889293|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889293|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889294|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889294|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889295|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY W RHEUMATOID ARTHRITIS MULT SITE
C2889295|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889296|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889297|T047||SNOMEDCT_US|RHEU ARTHRITIS OF R SHOULDER W INVOLV OF ORGANS AND SYSTEMS
C2889297|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889298|T047||SNOMEDCT_US|RHEU ARTHRITIS OF L SHOULDER W INVOLV OF ORGANS AND SYSTEMS
C2889298|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889299|T047||SNOMEDCT_US|RHEU ARTHRIT OF UNSP SHOULDER W INVOLV OF ORGANS AND SYSTEMS
C2889299|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889300|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889301|T047||SNOMEDCT_US|RHEU ARTHRITIS OF R ELBOW W INVOLV OF ORGANS AND SYSTEMS
C2889301|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889302|T047||SNOMEDCT_US|RHEU ARTHRITIS OF L ELBOW W INVOLV OF ORGANS AND SYSTEMS
C2889302|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889303|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP ELBOW W INVOLV OF ORGANS AND SYSTEMS
C2889303|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889304|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF CARPAL BONES WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889305|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889306|T047||SNOMEDCT_US|RHEU ARTHRITIS OF R WRIST W INVOLV OF ORGANS AND SYSTEMS
C2889306|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889307|T047||SNOMEDCT_US|RHEU ARTHRITIS OF L WRIST W INVOLV OF ORGANS AND SYSTEMS
C2889307|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889308|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP WRIST W INVOLV OF ORGANS AND SYSTEMS
C2889308|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889309|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF METACARPUS AND PHALANGES WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889310|T047||SNOMEDCT_US|RHEU ARTHRITIS OF RIGHT HAND W INVOLV OF ORGANS AND SYSTEMS
C2889310|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889311|T047||SNOMEDCT_US|RHEU ARTHRITIS OF LEFT HAND W INVOLV OF ORGANS AND SYSTEMS
C2889311|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889312|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP HAND W INVOLV OF ORGANS AND SYSTEMS
C2889312|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889313|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889314|T047||SNOMEDCT_US|RHEU ARTHRITIS OF RIGHT HIP W INVOLV OF ORGANS AND SYSTEMS
C2889314|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889315|T047||SNOMEDCT_US|RHEU ARTHRITIS OF LEFT HIP W INVOLV OF ORGANS AND SYSTEMS
C2889315|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889316|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP HIP W INVOLV OF ORGANS AND SYSTEMS
C2889316|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889317|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889318|T047||SNOMEDCT_US|RHEU ARTHRITIS OF RIGHT KNEE W INVOLV OF ORGANS AND SYSTEMS
C2889318|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889319|T047||SNOMEDCT_US|RHEU ARTHRITIS OF LEFT KNEE W INVOLV OF ORGANS AND SYSTEMS
C2889319|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889320|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP KNEE W INVOLV OF ORGANS AND SYSTEMS
C2889320|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889321|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF TARSUS, METATARSUS AND PHALANGES WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889322|T047||SNOMEDCT_US|RHEU ARTHRIT OF RIGHT ANK/FT W INVOLV OF ORGANS AND SYSTEMS
C2889322|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889323|T047||SNOMEDCT_US|RHEU ARTHRITIS OF LEFT ANK/FT W INVOLV OF ORGANS AND SYSTEMS
C2889323|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889324|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP ANK/FT W INVOLV OF ORGANS AND SYSTEMS
C2889324|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889325|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889326|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF UNSP SITE W/O ORG/SYS INVOLV
C2889326|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SITE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889327|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889328|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF R SHOULDER W/O ORG/SYS INVOLV
C2889328|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889329|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF L SHOULDER W/O ORG/SYS INVOLV
C2889329|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889330|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF UNSP SHLDR W/O ORG/SYS INVOLV
C2889330|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889331|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889332|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF R ELBOW W/O ORG/SYS INVOLV
C2889332|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889333|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF L ELBOW W/O ORG/SYS INVOLV
C2889333|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889334|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF UNSP ELBOW W/O ORG/SYS INVOLV
C2889334|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889335|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889336|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF R WRIST W/O ORG/SYS INVOLV
C2889336|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889337|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF L WRIST W/O ORG/SYS INVOLV
C2889337|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889338|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF UNSP WRIST W/O ORG/SYS INVOLV
C2889338|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889339|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889340|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF R HAND W/O ORG/SYS INVOLV
C2889340|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889341|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF LEFT HAND W/O ORG/SYS INVOLV
C2889341|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889342|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF UNSP HAND W/O ORG/SYS INVOLV
C2889342|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889343|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889344|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF RIGHT HIP W/O ORG/SYS INVOLV
C2889344|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889345|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF LEFT HIP W/O ORG/SYS INVOLV
C2889345|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889346|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF UNSP HIP W/O ORG/SYS INVOLV
C2889346|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889347|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889348|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF R KNEE W/O ORG/SYS INVOLV
C2889348|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889349|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF LEFT KNEE W/O ORG/SYS INVOLV
C2889349|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889350|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF UNSP KNEE W/O ORG/SYS INVOLV
C2889350|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889351|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889352|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FCTR OF RIGHT ANK/FT W/O ORG/SYS INVOLV
C2889352|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889353|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF LEFT ANK/FT W/O ORG/SYS INVOLV
C2889353|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889354|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF UNSP ANK/FT W/O ORG/SYS INVOLV
C2889354|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889355|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR MULT SITE W/O ORG/SYS INVOLV
C2889355|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF MULTIPLE SITES WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889356|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP SITE
C2889356|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR
C2889356|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SITE
C2889357|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF SHOULDER
C2889358|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF R SHOULDER
C2889358|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT SHOULDER
C2889359|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF L SHOULDER
C2889359|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT SHOULDER
C2889360|T047||SNOMEDCT_US|OTH RHEU ARTHRITIS W RHEUMATOID FACTOR OF UNSP SHOULDER
C2889360|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SHOULDER
C2889361|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF ELBOW
C2889362|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT ELBOW
C2889362|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ELBOW
C2889363|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF LEFT ELBOW
C2889363|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ELBOW
C2889364|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF UNSP ELBOW
C2889364|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ELBOW
C2889365|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF WRIST
C2889366|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT WRIST
C2889366|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT WRIST
C2889367|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF LEFT WRIST
C2889367|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT WRIST
C2889368|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF UNSP WRIST
C2889368|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED WRIST
C2889369|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT HAND
C2889369|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HAND
C2889370|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HAND
C2889370|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HAND
C2889371|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP HAND
C2889371|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF HAND
C2889371|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HAND
C2889372|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF HIP
C2889373|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HIP
C2889373|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HIP
C2889374|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HIP
C2889374|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HIP
C2889375|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP HIP
C2889375|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HIP
C2889376|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF KNEE
C2889377|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT KNEE
C2889377|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT KNEE
C2889378|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT KNEE
C2889378|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT KNEE
C2889379|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP KNEE
C2889379|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED KNEE
C2889380|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF ANKLE AND FOOT
C2889381|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT ANK/FT
C2889381|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ANKLE AND FOOT
C2889382|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF LEFT ANK/FT
C2889382|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ANKLE AND FOOT
C2889383|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF UNSP ANK/FT
C2889383|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ANKLE AND FOOT
C2889384|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR MULT SITE
C2889384|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF MULTIPLE SITES
C2889385|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR
C2889385|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR, UNSPECIFIED
C3469320|T047||SNOMEDCT_US|FELTYS SYNDROME, ELBOW
C3469320|T047||SNOMEDCT_US|FELTYS SYNDROME, UNSPECIFIED ELBOW
C3469322|T047||SNOMEDCT_US|FELTYS SYNDROME, HIP
C3469322|T047||SNOMEDCT_US|FELTYS SYNDROME, UNSPECIFIED HIP
C3469323|T047||SNOMEDCT_US|FELTYS SYNDROME, KNEE
C3469323|T047||SNOMEDCT_US|FELTYS SYNDROME, UNSPECIFIED KNEE
C3469325|T047||SNOMEDCT_US|FELTYS SYNDROME, SHOULDER
C3469326|T047||SNOMEDCT_US|FELTYS SYNDROME, WRIST
C3714757|T047|410795001|SNOMEDCT_US|NOT THE SAME AS RA, ALTHOUGH CAN BE RELASSIFIED AS RA WHEN THEY HIT ADULTHOOD|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|RHEUMATOID ARTHRITIS, JUVENILE|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|UNSPECIFIED JUVENILE RHEUMATOID ARTHRITIS|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JRA|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|CHILDHOOD ARTHRITIS|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE RHEUMATOID ARTHRITIS |JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JRA - JUVENILE RHEUMATOID ARTHRITIS|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE RHEUMATOID ARTHRITIS NOS |JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE RHEUMATOID ARTHRITIS NOS|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE RHEUMATOID A.|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE SEROPOSITIVE ARTHRITIS|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|RHEUMATOID ARTHRITIS IN CHILDREN|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE RA|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE ARTHRITIS|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE RHEUMATOID ARTHRITIS (AQ)|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS |JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE; ARTHRITIS, RHEUMATOID|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|ARTHRITIS; JUVENILE, RHEUMATOID|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, JUVENILE|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C3714757|T047|410795001|SNOMEDCT_US|JUVENILE RHEUMATOID ARTHRITIS, NOS|JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREWS DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE STRUEMPELL DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS, RHEUMATOID|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREW DIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE STRUEMPELL DIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREWS DIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLITIS |ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANK SPOND|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLOARTHRITIDES, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLOARTHRITIDES|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLARTHRITIDES, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLARTHRITIS, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLOARTHRITIS, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLARTHRITIDES|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SPINE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLARTHRITIS ANKYLOPOIETICA|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREW'S DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREW DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE-STRUEMPELL DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS, ANKYLOSING [DISEASE/FINDING]|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLARTHRITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLOARTHRITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|DISEASE;BECHTEREWS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLITIS |ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS ANKYLOPOIETICA|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLOARTHRITIS ANKYLOPOIETICA|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BEKHTEREV'S DISEASE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|AS - ANKYLOSING SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|IDIOPATHIC ANKYLOSING SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE-STRUMPELL SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE STRÜMPELL SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ARTHRITIS; SPINE OR VERTEBRA, MARIE-STRÜMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ARTHRITIS; SPINE OR VERTEBRA, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE-STRÜMPELL; SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|MARIE-STRÜMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|STRÜMPELL-MARIE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|VON BECHTEREW|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|BECHTEREW|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, SPINE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID; SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPINE OR VERTEBRA; ARTHRITIS, MARIE-STRÜMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPINE OR VERTEBRA; ARTHRITIS, ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS; MARIE-STRÜMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS; ANKYLOPOIETICA|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS; ANKYLOSING|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS; RHEUMATOID|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOPOIETICA; SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING; SPONDYLITIS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, SPINE|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|ANKYLOSING SPONDYLITIS, NOS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SPINE, NOS|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|SPONDYLITIS, MARIE-STRUMPELL|ANKYLOSING SPONDYLITIS (DISORDER)
C0038013|T047|9631008|SNOMEDCT_US|RHEUMATIOID ARTHRITIS OF SPINE NOS|ANKYLOSING SPONDYLITIS (DISORDER)
C0409628|T047|201792002|SNOMEDCT_US|OTHER RHEUMATOID ARTHROPATHY WITH VISCERAL OR SYSTEMIC INVOLVEMENT |OTHER RHEUMATOID ARTHROPATHY WITH VISCERAL OR SYSTEMIC INVOLVEMENT (DISORDER)
C0409628|T047|201792002|SNOMEDCT_US|OTHER RHEUMATOID ARTHROPATHY WITH VISCERAL OR SYSTEMIC INVOLVEMENT|OTHER RHEUMATOID ARTHROPATHY WITH VISCERAL OR SYSTEMIC INVOLVEMENT (DISORDER)
C0409629|T047|201785007|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF INTERPHALANGEAL JOINT OF TOE|RHEUMATOID ARTHRITIS OF INTERPHALANGEAL JOINT OF TOE (DISORDER)
C0409629|T047|201785007|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF INTERPHALANGEAL JOINT OF TOE |RHEUMATOID ARTHRITIS OF INTERPHALANGEAL JOINT OF TOE (DISORDER)
C0409630|T047|201784006|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LESSER METATARSOPHALANGEAL JOINT|RHEUMATOID ARTHRITIS OF LESSER METATARSOPHALANGEAL JOINT (DISORDER)
C0409630|T047|201784006|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LESSER METATARSOPHALANGEAL JOINT |RHEUMATOID ARTHRITIS OF LESSER METATARSOPHALANGEAL JOINT (DISORDER)
C0409631|T047|201783000|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF 1ST METATARSOPHALANGEAL JOINT|RHEUMATOID ARTHRITIS OF FIRST METATARSOPHALANGEAL JOINT (DISORDER)
C0409631|T047|201783000|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF FIRST METATARSOPHALANGEAL JOINT|RHEUMATOID ARTHRITIS OF FIRST METATARSOPHALANGEAL JOINT (DISORDER)
C0409631|T047|201783000|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF FIRST METATARSOPHALANGEAL JOINT |RHEUMATOID ARTHRITIS OF FIRST METATARSOPHALANGEAL JOINT (DISORDER)
C0409632|T047|201782005|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF OTHER TARSAL JOINT|RHEUMATOID ARTHRITIS OF OTHER TARSAL JOINT (DISORDER)
C0409632|T047|201782005|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF OTHER TARSAL JOINT |RHEUMATOID ARTHRITIS OF OTHER TARSAL JOINT (DISORDER)
C0409633|T047|201781003|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF TALONAVICULAR JOINT|RHEUMATOID ARTHRITIS OF TALONAVICULAR JOINT (DISORDER)
C0409633|T047|201781003|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF TALONAVICULAR JOINT |RHEUMATOID ARTHRITIS OF TALONAVICULAR JOINT (DISORDER)
C0409634|T047|201780002|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SUBTALAR JOINT|RHEUMATOID ARTHRITIS OF SUBTALAR JOINT (DISORDER)
C0409634|T047|201780002|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SUBTALAR JOINT |RHEUMATOID ARTHRITIS OF SUBTALAR JOINT (DISORDER)
C0409635|T047|201779000|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ANKLE |RHEUMATOID ARTHRITIS OF ANKLE (DISORDER)
C0409635|T047|201779000|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ANKLE|RHEUMATOID ARTHRITIS OF ANKLE (DISORDER)
C0409635|T047|201779000|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ANKLE |RHEUMATOID ARTHRITIS OF ANKLE (DISORDER)
C0409637|T047|201777003|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF KNEE|RHEUMATOID ARTHRITIS OF KNEE (DISORDER)
C0409637|T047|201777003|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF KNEE |RHEUMATOID ARTHRITIS OF KNEE (DISORDER)
C0409637|T047|201777003|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF KNEE |RHEUMATOID ARTHRITIS OF KNEE (DISORDER)
C0409639|T047|201775006|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HIP|RHEUMATOID ARTHRITIS OF HIP (DISORDER)
C0409639|T047|201775006|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HIP |RHEUMATOID ARTHRITIS OF HIP (DISORDER)
C0409639|T047|201775006|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HIP |RHEUMATOID ARTHRITIS OF HIP (DISORDER)
C0409640|T047|201774005|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF DISTAL INTERPHALANGEAL JOINT OF FINGER|RHEUMATOID ARTHRITIS OF DISTAL INTERPHALANGEAL JOINT OF FINGER (DISORDER)
C0409640|T047|201774005|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF DISTAL INTERPHALANGEAL JOINT OF FINGER |RHEUMATOID ARTHRITIS OF DISTAL INTERPHALANGEAL JOINT OF FINGER (DISORDER)
C0409641|T047|201773004|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF PROXIMAL INTERPHALANGEAL JOINT OF FINGER|RHEUMATOID ARTHRITIS OF PROXIMAL INTERPHALANGEAL JOINT OF FINGER (DISORDER)
C0409641|T047|201773004|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF PROXIMAL INTERPHALANGEAL JOINT OF FINGER |RHEUMATOID ARTHRITIS OF PROXIMAL INTERPHALANGEAL JOINT OF FINGER (DISORDER)
C0409642|T047|201772009|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF METACARPOPHALANGEAL JOINT|RHEUMATOID ARTHRITIS OF METACARPOPHALANGEAL JOINT (DISORDER)
C0409642|T047|201772009|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF METACARPOPHALANGEAL JOINT |RHEUMATOID ARTHRITIS OF METACARPOPHALANGEAL JOINT (DISORDER)
C0409643|T047|201771002|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF WRIST|RHEUMATOID ARTHRITIS OF WRIST (DISORDER)
C0409643|T047|201771002|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF WRIST |RHEUMATOID ARTHRITIS OF WRIST (DISORDER)
C0409643|T047|201771002|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF WRIST |RHEUMATOID ARTHRITIS OF WRIST (DISORDER)
C0409645|T047|201769002|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ELBOW |RHEUMATOID ARTHRITIS OF ELBOW (DISORDER)
C0409645|T047|201769002|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ELBOW|RHEUMATOID ARTHRITIS OF ELBOW (DISORDER)
C0409645|T047|201769002|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ELBOW |RHEUMATOID ARTHRITIS OF ELBOW (DISORDER)
C0409646|T047|201768005|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ACROMIOCLAVICULAR JOINT|RHEUMATOID ARTHRITIS OF ACROMIOCLAVICULAR JOINT (DISORDER)
C0409646|T047|201768005|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ACROMIOCLAVICULAR JOINT |RHEUMATOID ARTHRITIS OF ACROMIOCLAVICULAR JOINT (DISORDER)
C0409647|T047|201767000|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF STERNOCLAVICULAR JOINT|RHEUMATOID ARTHRITIS OF STERNOCLAVICULAR JOINT (DISORDER)
C0409647|T047|201767000|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF STERNOCLAVICULAR JOINT |RHEUMATOID ARTHRITIS OF STERNOCLAVICULAR JOINT (DISORDER)
C0409648|T047|201766009|SNOMEDCT_US|RHEUMATOID ARTHRITIS SHOULDER |RHEUMATOID ARTHRITIS OF SHOULDER (DISORDER)
C0409648|T047|201766009|SNOMEDCT_US|RHEUMATOID ARTHRITIS SHOULDER|RHEUMATOID ARTHRITIS OF SHOULDER (DISORDER)
C0409648|T047|201766009|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SHOULDER|RHEUMATOID ARTHRITIS OF SHOULDER (DISORDER)
C0409648|T047|201766009|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SHOULDER |RHEUMATOID ARTHRITIS OF SHOULDER (DISORDER)
C0409650|T047|201764007|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF CERVICAL SPINE|RHEUMATOID ARTHRITIS OF CERVICAL SPINE (DISORDER)
C0409650|T047|201764007|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF CERVICAL SPINE |RHEUMATOID ARTHRITIS OF CERVICAL SPINE (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|SEROPOSITIVE RHEUMATOID ARTHRITIS|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|RHEUMATOID FACTOR POSITIVE |[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|RHEUMATOID FACTOR POSITIVE|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED |[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|SEROPOSITIVE RA|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|SEROPOSITIVE RHEUMATOID ARTHRITIS |[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, SEROPOSITIVE|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409651|T047|203746006|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, SEROPOSITIVE|[X]SEROPOSITIVE RHEUMATOID ARTHRITIS, UNSPECIFIED (DISORDER)
C0409652|T047|239792003|SNOMEDCT_US|SERONEGATIVE RHEUMATOID ARTHRITIS|SERONEGATIVE RHEUMATOID ARTHRITIS (DISORDER)
C0409652|T047|239792003|SNOMEDCT_US|SERONEGATIVE RHEUMATOID ARTHRITIS |SERONEGATIVE RHEUMATOID ARTHRITIS (DISORDER)
C0409652|T047|239792003|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, SERONEGATIVE|SERONEGATIVE RHEUMATOID ARTHRITIS (DISORDER)
C0409652|T047|239792003|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, SERONEGATIVE|SERONEGATIVE RHEUMATOID ARTHRITIS (DISORDER)
C0409657|T047|239795001|SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH MULTISYSTEM INVOLVEMENT|RHEUMATOID ARTHRITIS WITH MULTISYSTEM INVOLVEMENT (DISORDER)
C0409657|T047|239795001|SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH MULTISYSTEM INVOLVEMENT |RHEUMATOID ARTHRITIS WITH MULTISYSTEM INVOLVEMENT (DISORDER)
C0856832|T047||SNOMEDCT_US|MONOARTHRITIC RHEUMATOID ARTHRITIS
C0477541|T047|203730003|SNOMEDCT_US|OTHER SEROPOSITIVE RHEUMATOID ARTHRITIS|[X]OTHER SEROPOSITIVE RHEUMATOID ARTHRITIS (DISORDER)
C0477541|T047|203730003|SNOMEDCT_US|[X]OTHER SEROPOSITIVE RHEUMATOID ARTHRITIS|[X]OTHER SEROPOSITIVE RHEUMATOID ARTHRITIS (DISORDER)
C0477541|T047|203730003|SNOMEDCT_US|[X]OTHER SEROPOSITIVE RHEUMATOID ARTHRITIS |[X]OTHER SEROPOSITIVE RHEUMATOID ARTHRITIS (DISORDER)
C0494896|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0494896|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH SYSTEMIC INVOLVEMENT
C0494896|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH SYSTEMIC INVOLVEMENT
C0235762|T047||SNOMEDCT_US|ARTHRITIS RHEUMATOID AGGRAVATED
C0235762|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS AGGRAVATED
C0837691|T047||SNOMEDCT_US|JUV RHEUM ARTHRITIS NOS
C0837691|T047||SNOMEDCT_US|POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS, CHRONIC OR UNSPECIFIED
C0837691|T047||SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS OF MULTIPLE SITES
C0837691|T047||SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS MULTIPLE SITES
C0837691|T047||SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS OF MULTIPLE SITES 
C0263737|T047|86219005|SNOMEDCT_US|UVEITIS-RHEUMATOID ARTHRITIS SYNDROME|UVEITIS-RHEUMATOID ARTHRITIS SYNDROME (DISORDER)
C0263737|T047|86219005|SNOMEDCT_US|UVEITIS-RHEUMATOID ARTHRITIS SYNDROME |UVEITIS-RHEUMATOID ARTHRITIS SYNDROME (DISORDER)
C0157914|T047|111218008|SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH VISCERAL OR SYSTEMIC INVOLVEMENT|RHEUMATOID ARTHRITIS WITH OTHER VISCERAL OR SYSTEMIC INVOLVEMENT (DISORDER)
C0157914|T047|111218008|SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH OTHER VISCERAL OR SYSTEMIC INVOLVEMENT -RETIRED-|RHEUMATOID ARTHRITIS WITH OTHER VISCERAL OR SYSTEMIC INVOLVEMENT (DISORDER)
C0157914|T047|111218008|SNOMEDCT_US|SYST RHEUM ARTHRITIS NEC|RHEUMATOID ARTHRITIS WITH OTHER VISCERAL OR SYSTEMIC INVOLVEMENT (DISORDER)
C0157914|T047|111218008|SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH OTHER VISCERAL OR SYSTEMIC INVOLVEMENT |RHEUMATOID ARTHRITIS WITH OTHER VISCERAL OR SYSTEMIC INVOLVEMENT (DISORDER)
C0157914|T047|111218008|SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH OTHER VISCERAL OR SYSTEMIC INVOLVEMENT|RHEUMATOID ARTHRITIS WITH OTHER VISCERAL OR SYSTEMIC INVOLVEMENT (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR JUVENILE ARTHRITIS|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|OLIGOARTICULAR STILL DISEASE|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|OLIGOARTICULAR STILL'S DISEASE|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIART JUV RHEUM ARTHR|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSPECIFIED SITE|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS, UNSP SITE|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS |PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR JRA|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR JUVENILE CHRONIC RA|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS (AQ)|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|OLIGOARTICULAR JRA|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|OLIGOARTICULAR JUVENILE RHEUMATOID ARTHRITIS|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|JCA - PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR ONSET JUVENILE ARTHRITIS|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|PAUCIARTICULAR JUVENILE RHEUMATOID ARTHRITIS |PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|JUVENILE; ARTHRITIS, PAUCIARTICULAR|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0157917|T047|201809006|SNOMEDCT_US|ARTHRITIS; JUVENILE, PAUCIARTICULAR|PAUCIARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0409636|T047|201778008|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF TIBIOFIBULAR JOINT|RHEUMATOID ARTHRITIS OF TIBIOFIBULAR JOINT (DISORDER)
C0409636|T047|201778008|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF TIBIOFIBULAR JOINT |RHEUMATOID ARTHRITIS OF TIBIOFIBULAR JOINT (DISORDER)
C0409644|T047|201770001|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF DISTAL RADIOULNAR JOINT|RHEUMATOID ARTHRITIS OF DISTAL RADIOULNAR JOINT (DISORDER)
C0409644|T047|201770001|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF DISTAL RADIOULNAR JOINT |RHEUMATOID ARTHRITIS OF DISTAL RADIOULNAR JOINT (DISORDER)
C0409638|T047|201776007|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SACROILIAC JOINT|RHEUMATOID ARTHRITIS OF SACROILIAC JOINT (DISORDER)
C0409638|T047|201776007|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SACROILIAC JOINT |RHEUMATOID ARTHRITIS OF SACROILIAC JOINT (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|CAPLANS SYNDROME|RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|CAPLAN'S SYNDROME|RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|CAPLAN'S SYNDROME |RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|CAPLAN SYNDROME|RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|CAPLAN SYNDROMES|RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|CAPLAN SYNDROME [DISEASE/FINDING]|RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|RHEUMATOID PNEUMOCONIOSIS |RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|RHEUMATOID PNEUMOCONIOSIS|RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|CAPLAN (ETIOLOGY)|RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0006915|T047|398640008|SNOMEDCT_US|CAPLAN (MANIFESTATION)|RHEUMATOID PNEUMOCONIOSIS (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTYS SYNDROME|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|SYNDROME, FELTY'S|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTY'S SYNDROME|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTY SYNDROME|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTY'S SYNDROME |FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH SPLENOADENOMEGALY AND LEUKOPENIA|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTY'S SYNDROME, UNSPECIFIED SITE|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|SYNDROME, FELTY|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTY SYNDROME [DISEASE/FINDING]|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTY'S SYNDROME |FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|RHEUMATOID ARTHRITIS, LEUCOPENIA AND SPLENOMEGALY|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|RHEUMATOID ARTHRITIS, LEUKOPENIA AND SPLENOMEGALY|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|FELTY|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH SPLENOADENOMEGALY AND LEUKOPENIA|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH SPLENOADENOMEGALY AND LEUKOPENIA|FELTY'S SYNDROME (DISORDER)
C0015773|T047|57160007|SNOMEDCT_US|RHEUMATOID ARTHRITIS, LEUKOPENIA AND SPLENADENOMEGALY|FELTY'S SYNDROME (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|NODULE, RHEUMATOID|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|NODULES, RHEUMATOID|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID NODULE|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID NODULES|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID NODULOSIS|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID NODULE [DISEASE/FINDING]|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID NODULOSES|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID NODULE |RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|SUBCUTANEOUS RHEUMATOID NODULE|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID NODULE (MORPHOLOGIC ABNORMALITY)|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID NODULOSIS |RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|SUBCUTANEOUS RHEUMATOID NODULE |RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|NODE; RHEUMATOID|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|NODULE; RHEUMATOID|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID; NODE|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID; NODULE|RHEUMATOID NODULE (DISORDER)
C0035450|T047|201789001|SNOMEDCT_US|RHEUMATOID NODULE, NOS|RHEUMATOID NODULE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT ONSET STILL DISEASE|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT ONSET STILL'S DISEASE|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT-ONSET STILLS DISEASE|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILL DISEASE, ADULT ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILL'S DISEASE, ADULT ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILL'S DISEASE, ADULT-ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILLS DISEASE, ADULT-ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT-ONSET STILL'S DISEASE|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT-ONSET STILL DISEASE|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT ONSET STILL DIS|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILLS DIS ADULT ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT ONSET STILLS DIS|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILL DIS ADULT ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILL'S DISEASE ADULT ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT ONSET STILL'S DISEASE |ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|AOSD (ADULT ONSET STILL'S DISEASE)|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT STILL'S DISEASE|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILL'S DISEASE, ADULT-ONSET [DISEASE/FINDING]|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILL DISEASE, ADULT-ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT ONSET STILL'S DISEASE |ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|DISEASE; STILL'S ADULT ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILL'S ADULT ONSET; DISEASE|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|STILL; ADULT-ONSET|ADULT ONSET STILL'S DISEASE (DISORDER)
C0085253|T047|239920006|SNOMEDCT_US|ADULT-ONSET; STILL|ADULT ONSET STILL'S DISEASE (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS, RHEUMATOID|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS, UNSPECIFIED|RHEUMATOID ARTHRITIS (DISORDER)
# C0003873|T047|69896004|SNOMEDCT_US|RA|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RA (RHEUMATOID ARTHRITIS)|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS |RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|R ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RH ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS, RHEUMATOID [DISEASE/FINDING]|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS NOS |RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS NOS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID ARTHRITIS |RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS RHEUMATOID|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ATROPHIC ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|SYSTEMIC RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|CHRONIC RHEUMATIC ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATIC GOUT|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RA - RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHA - RHEUMATOID ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID DISEASE|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ATROPHIC; ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|RHEUMATOID; ARTHRITIS|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS; ATROPHIC|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS; RHEUMATOID|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS OR POLYARTHRITIS, ATROPHIC|RHEUMATOID ARTHRITIS (DISORDER)
C0003873|T047|69896004|SNOMEDCT_US|ARTHRITIS OR POLYARTHRITIS, RHEUMATIC|RHEUMATOID ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|CHRONIC ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|RHEUMATOID ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE ARTHRITIS, UNSPECIFIED|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE CHRONIC|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE CHRONIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE RHEUMATOID ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE IDIOPATHIC|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE ARTHRITIS |JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ENTHESITIS RELATED ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE OLIGOARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE SYSTEMIC|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE ENTHESITIS-RELATED ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE SYSTEMIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE PSORIATIC|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE PSORIATIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE ENTHESITIS-RELATED|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|OLIGOARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE RHEUMATOID|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ENTHESITIS-RELATED ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|PSORIATIC ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|SYSTEMIC ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS, JUVENILE [DISEASE/FINDING]|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JIA|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|POLYARTHRITIS, JUVENILE, RHEUMATOID FACTOR POSITIVE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|POLYARTHRITIS, JUVENILE, RHEUMATOID FACTOR NEGATIVE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JCA - JUVENILE CHRONIC ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE CHRONIC ARTHRITIS |JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE; ARTHRITIS|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS; JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE CHRONIC ARTHRITIS, POLYARTICULAR SEROPOSITIVE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS |JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS, POLYARTHRITIS, RHEUMATOID FACTOR POSITIVE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|IDIOPATHIC ARTHRITIS, JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C3495559|T047|410502007|SNOMEDCT_US|ARTHRITIS;JUVENILE|JUVENILE IDIOPATHIC ARTHRITIS (DISORDER)
C0409679|T047|399112009|SNOMEDCT_US|SERONEGATIVE ARTHRITIS|SERONEGATIVE ARTHRITIS (DISORDER)
C0409679|T047|399112009|SNOMEDCT_US|SERONEGATIVE ARTHRITIS |SERONEGATIVE ARTHRITIS (DISORDER)
C0409679|T047|399112009|SNOMEDCT_US|SERONEGATIVE POLYARTHRITIS|SERONEGATIVE ARTHRITIS (DISORDER)
C0409679|T047|399112009|SNOMEDCT_US|SERO NEGATIVE ARTHROPATHY|SERONEGATIVE ARTHRITIS (DISORDER)
C0409679|T047|399112009|SNOMEDCT_US|SERONEGATIVE ARTHRITIS NOS|SERONEGATIVE ARTHRITIS (DISORDER)
C0409679|T047|399112009|SNOMEDCT_US|SERONEGATIVE ARTHROPATHY|SERONEGATIVE ARTHRITIS (DISORDER)
C0409679|T047|399112009|SNOMEDCT_US|SERONEGATIVE ARTHRITIS [AMBIGUOUS]|SERONEGATIVE ARTHRITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|RHEUMATOID VASCULITIS|RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|RHEUMATOID VASCULITIS |RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|VASCULITIDES, RHEUMATOID|RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|VASCULITIS, RHEUMATOID|RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|RHEUMATOID VASCULITIDES|RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|RHEUMATOID VASCULITIS [DISEASE/FINDING]|RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|RHEUMATOID VASCULITIS |RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH VASCULITIS|RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|RHEUMATOID; VASCULITIS|RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|VASCULITIS; RHEUMATOID|RHEUMATOID VASCULITIS (DISORDER)
C0240903|T047|400054000|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH VASCULITIS|RHEUMATOID VASCULITIS (DISORDER)
C2200410|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF FINGERS
C2200410|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF FINGERS 
C2200418|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF TOES 
C2200418|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF TOES
C0427391|T047|165840002|SNOMEDCT_US|RHEUMATOID FACTOR NEGATIVE|RHEUMATOID FACTOR NEGATIVE (FINDING)
C0427391|T047|165840002|SNOMEDCT_US|NEGATIVE RHEUMATOID FACTOR|RHEUMATOID FACTOR NEGATIVE (FINDING)
C0427391|T047|165840002|SNOMEDCT_US|RHEUMATOID FACTOR NEGATIVE |RHEUMATOID FACTOR NEGATIVE (FINDING)
C0427391|T047|165840002|SNOMEDCT_US|RHEUMATIOD FACTOR NEGATIVE|RHEUMATOID FACTOR NEGATIVE (FINDING)
C0427391|T047|165840002|SNOMEDCT_US|RHEUMATOID FACTOR NEGATIVE |RHEUMATOID FACTOR NEGATIVE (FINDING)
C2200417|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS STEINBROCKER CLASSIFICATION (___0-IV)
C2200417|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS STEINBROCKER CLASSIFICATION (___0-IV) 
C2062580|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH ATLANTOAXIAL SUBLUXATION 
C2062580|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH ATLANTOAXIAL SUBLUXATION
C0085574|T047|202456000|SNOMEDCT_US|THIS IS A SLIGHTLY DIFFERENT BUT I THINK SHOULD SHOW UP IF YOU ARE ASKING ABOUT RA|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROM RHEUM-UNSPEC|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROMIC RHEUMATISM, UNSPECIFIED SITE|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROMIC RHEUMATISM SYNDROME|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROMIC RHEUMATISM NOS |PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROMIC RHEUMATISM NOS|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE |PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|HENCH - ROSENBERG SYNDROME|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROMIC RHEUMATISM, SITE UNSPECIFIED|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|HENCH-ROSENBERG SYNDROME|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROMIC RHEUMATISM |PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|PALINDROMIC; RHEUMATISM|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C0085574|T047|202456000|SNOMEDCT_US|RHEUMATISM; PALINDROMIC|PALINDROMIC RHEUMATISM OF UNSPECIFIED SITE (DISORDER)
C3469328|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS NODULE
C3469328|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS NODULE 
C0451843|T047|201788009|SNOMEDCT_US|RHEUMATOID BURSITIS|RHEUMATOID BURSITIS (DISORDER)
C0451843|T047|201788009|SNOMEDCT_US|RHEUMATOID BURSITIS, UNSPECIFIED SITE|RHEUMATOID BURSITIS (DISORDER)
C0451843|T047|201788009|SNOMEDCT_US|RHEUMATOID BURSITIS |RHEUMATOID BURSITIS (DISORDER)
C0451843|T047|201788009|SNOMEDCT_US|RHEUMATOID BURSITIS |RHEUMATOID BURSITIS (DISORDER)
C0451843|T047|201788009|SNOMEDCT_US|BURSITIS; RHEUMATOID|RHEUMATOID BURSITIS (DISORDER)
C0451843|T047|201788009|SNOMEDCT_US|RHEUMATOID; BURSITIS|RHEUMATOID BURSITIS (DISORDER)
C2889134|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889134|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF SHOULDER 
C2889138|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889138|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF ELBOW 
C2889143|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF WRIST
C2889143|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF WRIST 
C2889148|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF HAND
C2889148|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF HAND 
C2889152|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889152|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF HIP
C2889152|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP HIP
C2889152|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF HIP 
C2889155|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF KNEE
C2889155|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF KNEE 
C2889160|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889160|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT 
C2889168|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889168|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889168|T047||SNOMEDCT_US|RHEU VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889168|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF SHOULDER 
C2889169|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889169|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF ELBOW 
C2889174|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF WRIST
C2889174|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF WRIST 
C0564785|T047|287007001|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HAND JOINT|RHEUMATOID ARTHRITIS OF HAND JOINT (DISORDER)
C0564785|T047|287007001|SNOMEDCT_US|RHEUMATOID ARTHRITIS - HAND JOINT |RHEUMATOID ARTHRITIS OF HAND JOINT (DISORDER)
C0564785|T047|287007001|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HAND JOINT |RHEUMATOID ARTHRITIS OF HAND JOINT (DISORDER)
C0564785|T047|287007001|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HAND |RHEUMATOID ARTHRITIS OF HAND JOINT (DISORDER)
C0564785|T047|287007001|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HAND|RHEUMATOID ARTHRITIS OF HAND JOINT (DISORDER)
C0564785|T047|287007001|SNOMEDCT_US|RHEUMATOID ARTHRITIS - HAND JOINT|RHEUMATOID ARTHRITIS OF HAND JOINT (DISORDER)
C0564786|T047|156479006|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ANKLE AND/OR FOOT|RHEUMATOID ARTHRITIS - ANKLE/FOOT (DISORDER)
C0564786|T047|156479006|SNOMEDCT_US|RHEUMATOID ARTHRITIS - ANKLE AND/OR FOOT |RHEUMATOID ARTHRITIS - ANKLE/FOOT (DISORDER)
C0564786|T047|156479006|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ANKLE AND/OR FOOT |RHEUMATOID ARTHRITIS - ANKLE/FOOT (DISORDER)
C0564786|T047|156479006|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ANKLE AND FOOT |RHEUMATOID ARTHRITIS - ANKLE/FOOT (DISORDER)
C0564786|T047|156479006|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ANKLE AND FOOT|RHEUMATOID ARTHRITIS - ANKLE/FOOT (DISORDER)
C0564786|T047|156479006|SNOMEDCT_US|RHEUMATOID ARTHRITIS ANKLE AND FOOT|RHEUMATOID ARTHRITIS - ANKLE/FOOT (DISORDER)
C0564786|T047|156479006|SNOMEDCT_US|RHEUMATOID ARTHRITIS - ANKLE/FOOT |RHEUMATOID ARTHRITIS - ANKLE/FOOT (DISORDER)
C0564786|T047|156479006|SNOMEDCT_US|RHEUMATOID ARTHRITIS - ANKLE/FOOT|RHEUMATOID ARTHRITIS - ANKLE/FOOT (DISORDER)
C0564786|T047|156479006|SNOMEDCT_US|RHEUMATOID ARTHRITIS - ANKLE AND/OR FOOT|RHEUMATOID ARTHRITIS - ANKLE/FOOT (DISORDER)
C3508970|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS VERTEBRAE
C3508970|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS VERTEBRAE 
C3508971|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS MULTIPLE SITES
C3508971|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS MULTIPLE SITES 
C0265176|T047|7607008|SNOMEDCT_US|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0265176|T047|7607008|SNOMEDCT_US|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS |PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0265176|T047|7607008|SNOMEDCT_US|PERICARDITIS; RHEUMATOID ARTHRITIS (ETIOLOGY)|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0265176|T047|7607008|SNOMEDCT_US|PERICARDITIS; RHEUMATOID ARTHRITIS (MANIFESTATION)|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0265176|T047|7607008|SNOMEDCT_US|RHEUMATOID ARTHRITIS; PERICARDITIS (ETIOLOGY)|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0265176|T047|7607008|SNOMEDCT_US|RHEUMATOID ARTHRITIS; PERICARDITIS (MANIFESTATION)|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0265176|T047|7607008|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH PERICARDITIS (ETIOLOGY)|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0265176|T047|7607008|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH PERICARDITIS (MANIFESTATION)|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0265176|T047|7607008|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH PERICARDITIS (ETIOLOGY)|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0265176|T047|7607008|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH PERICARDITIS (MANIFESTATION)|PERICARDITIS SECONDARY TO RHEUMATOID ARTHRITIS (DISORDER)
C0564787|T047|156480009|SNOMEDCT_US|RHEUMATOID ARTHRITIS - OTHER JOINT|RHEUMATOID ARTHRITIS - OTHER JOINT (DISORDER)
C0564787|T047|156480009|SNOMEDCT_US|RHEUMATOID ARTHRITIS - OTHER JOINT |RHEUMATOID ARTHRITIS - OTHER JOINT (DISORDER)
C0409649|T047|201765008|SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS OF SPINE|OTHER RHEUMATOID ARTHRITIS OF SPINE (DISORDER)
C0409649|T047|201765008|SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS OF SPINE |OTHER RHEUMATOID ARTHRITIS OF SPINE (DISORDER)
C3836171|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE WITHOUT INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C3836171|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE WITHOUT INVOLVEMENT OF OTHER ORGANS AND SYSTEMS 
C3899278|T047||SNOMEDCT_US|EARLY RHEUMATOID ARTHRITIS
C0702102|T047|200958001|SNOMEDCT_US|ARTHRITIS MUTILANS|PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE (DISORDER)
C0702102|T047|200958001|SNOMEDCT_US|PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE|PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE (DISORDER)
C0702102|T047|200958001|SNOMEDCT_US|PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE |PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE (DISORDER)
C0702102|T047|200958001|SNOMEDCT_US|ARTHRITIS MUTILANS |PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE (DISORDER)
C0702102|T047|200958001|SNOMEDCT_US|MUTILANS; ARTHRITIS (ETIOLOGY)|PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE (DISORDER)
C0702102|T047|200958001|SNOMEDCT_US|MUTILANS; ARTHRITIS (MANIFESTATION)|PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE (DISORDER)
C0702102|T047|200958001|SNOMEDCT_US|ARTHRITIS; MUTILANS (ETIOLOGY)|PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE (DISORDER)
C0702102|T047|200958001|SNOMEDCT_US|ARTHRITIS; MUTILANS (MANIFESTATION)|PSORIATIC ARTHRITIS - DESTRUCTIVE TYPE (DISORDER)
C0409653|T047|239793008|SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH ORGAN / SYSTEM INVOLVEMENT|RHEUMATOID ARTHRITIS WITH ORGAN / SYSTEM INVOLVEMENT (DISORDER)
C0409653|T047|239793008|SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH ORGAN / SYSTEM INVOLVEMENT |RHEUMATOID ARTHRITIS WITH ORGAN / SYSTEM INVOLVEMENT (DISORDER)
C0477542|T047|203732006|SNOMEDCT_US|OTHER SPECIFIED RHEUMATOID ARTHRITIS|[X]OTHER SPECIFIED RHEUMATOID ARTHRITIS (DISORDER)
C0477542|T047|203732006|SNOMEDCT_US|OTHER SPECIFIED RHEUMATOID ARTHRITIS, UNSPECIFIED SITE|[X]OTHER SPECIFIED RHEUMATOID ARTHRITIS (DISORDER)
C0477542|T047|203732006|SNOMEDCT_US|[X]OTHER SPECIFIED RHEUMATOID ARTHRITIS|[X]OTHER SPECIFIED RHEUMATOID ARTHRITIS (DISORDER)
C0477542|T047|203732006|SNOMEDCT_US|[X]OTHER SPECIFIED RHEUMATOID ARTHRITIS |[X]OTHER SPECIFIED RHEUMATOID ARTHRITIS (DISORDER)
C0581345|T047|201791009|SNOMEDCT_US|FLARE OF RHEUMATOID ARTHRITIS|FLARE OF RHEUMATOID ARTHRITIS (DISORDER)
C0581345|T047|201791009|SNOMEDCT_US|FLARE OF RHEUMATOID ARTHRITIS |FLARE OF RHEUMATOID ARTHRITIS (DISORDER)
C0564784|T047|287006005|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF MULTIPLE JOINTS|RHEUMATOID ARTHRITIS OF MULTIPLE JOINTS (DISORDER)
C0564784|T047|287006005|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF MULTIPLE JOINTS |RHEUMATOID ARTHRITIS OF MULTIPLE JOINTS (DISORDER)
C0564784|T047|287006005|SNOMEDCT_US|RHEUMATOID ARTHRITIS - MULTIPLE JOINT |RHEUMATOID ARTHRITIS OF MULTIPLE JOINTS (DISORDER)
C0564784|T047|287006005|SNOMEDCT_US|RHEUMATOID ARTHRITIS - MULTIPLE JOINT|RHEUMATOID ARTHRITIS OF MULTIPLE JOINTS (DISORDER)
C0263741|T047|52661003|SNOMEDCT_US|EXTRA-ARTICULAR RHEUMATOID PROCESS |EXTRA-ARTICULAR RHEUMATOID PROCESS (DISORDER)
C0263741|T047|52661003|SNOMEDCT_US|EXTRA-ARTICULAR RHEUMATOID PROCESS|EXTRA-ARTICULAR RHEUMATOID PROCESS (DISORDER)
C0263741|T047|52661003|SNOMEDCT_US|EXTRA-ARTICULAR RHEUMATOID PROCESS, NOS|EXTRA-ARTICULAR RHEUMATOID PROCESS (DISORDER)
C0866632|T047||SNOMEDCT_US|ARTHRITIS OR POLYARTHITIS, CHRONIC RHEUMATIC
C1405320|T047||SNOMEDCT_US|POLYARTHRITIS; RHEUMATOID
C1405320|T047||SNOMEDCT_US|RHEUMATOID; POLYARTHRITIS
C1406307|T047||SNOMEDCT_US|RHEUMATOID\\SEE ALSO CONDITION
C0087031|T047|123246003|SNOMEDCT_US|STILL'S DISEASE|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE ONSET STILL DISEASE|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE ONSET STILLS DISEASE|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE-ONSET STILL'S DISEASE|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL DISEASE, JUVENILE ONSET|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL'S DISEASE, JUVENILE ONSET|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILLS DISEASE, JUVENILE-ONSET|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE-ONSET STILL DISEASE|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL DISEASE JUVENILE ONSET|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE ONSET STILL DIS|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE ONSET STILLS DIS|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILLS DIS JUVENILE ONSET|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL'S DISEASE -RETIRED-|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE ONSET STILL'S DISEASE |STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE STILL'S DISEASE|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE ONSET STILL'S DISEASE|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL DISEASE|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL'S DISEASE NOS|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL'S DISEASE - JUVENILE R.A|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL'S DISEASE |STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL'S DISEASE - JUVENILE RHEUMATOID ARTHRITIS |STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL'S DISEASE - JUVENILE RHEUMATOID ARTHRITIS|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|SYSTEMIC ONSET JUVENILE RHEUMATOID ARTHRITIS|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|SYSTEMIC JRA|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|SJRA|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|SYSTEMIC JUVENILE RHEUMATOID ARTHRITIS (AQ)|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|JUVENILE-ONSET STILLS DISEASE|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL DISEASE, JUVENILE-ONSET|STILL'S DISEASE (DISORDER)
C0087031|T047|123246003|SNOMEDCT_US|STILL'S DISEASE, JUVENILE-ONSET|STILL'S DISEASE (DISORDER)
C0421288|T047|148074006|SNOMEDCT_US|RHEUMATOLOGY DISORDER - JOINTS AFFECTED |RHEUMATOLOGY DISORDER - JOINTS AFFECTED (DISORDER)
C0421288|T047|148074006|SNOMEDCT_US|RHEUMATOLOGY DISORDER - JOINTS AFFECTED|RHEUMATOLOGY DISORDER - JOINTS AFFECTED (DISORDER)
C0421288|T047|148074006|SNOMEDCT_US|RHEUMATOLOGY DISORDER - JOINTS AFFECTED |RHEUMATOLOGY DISORDER - JOINTS AFFECTED (DISORDER)
C1998379|T047|427770001|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF TEMPOROMANDIBULAR JOINT |RHEUMATOID ARTHRITIS OF TEMPOROMANDIBULAR JOINT (DISORDER)
C1998379|T047|427770001|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF TEMPOROMANDIBULAR JOINT|RHEUMATOID ARTHRITIS OF TEMPOROMANDIBULAR JOINT (DISORDER)
C1998063|T047|429422002|SNOMEDCT_US|RHEUMATIC ARTHRITIS OF TEMPOROMANDIBULAR JOINT |RHEUMATIC ARTHRITIS OF TEMPOROMANDIBULAR JOINT (DISORDER)
C1998063|T047|429422002|SNOMEDCT_US|RHEUMATIC ARTHRITIS OF TEMPOROMANDIBULAR JOINT|RHEUMATIC ARTHRITIS OF TEMPOROMANDIBULAR JOINT (DISORDER)
C0585962|T047|201810001|SNOMEDCT_US|SEROPOSITIVE ERROSIVE RHEUMATOID ARTHRITIS |SEROPOSITIVE ERROSIVE RHEUMATOID ARTHRITIS (DISORDER)
C0585962|T047|201810001|SNOMEDCT_US|SEROPOSITIVE ERROSIVE RHEUMATOID ARTHRITIS|SEROPOSITIVE ERROSIVE RHEUMATOID ARTHRITIS (DISORDER)
C1304220|T047|402434001|SNOMEDCT_US|CUTANEOUS COMPLICATION OF RHEUMATOID DISEASE |CUTANEOUS COMPLICATION OF RHEUMATOID DISEASE (DISORDER)
C1304220|T047|402434001|SNOMEDCT_US|CUTANEOUS COMPLICATION OF RHEUMATOID DISEASE|CUTANEOUS COMPLICATION OF RHEUMATOID DISEASE (DISORDER)
C0409579|T047|14175009|SNOMEDCT_US|ARTICULAR RHEUMATIC FEVER|RHEUMATIC JOINT DISEASE (DISORDER)
C0409579|T047|14175009|SNOMEDCT_US|RHEUMATIC JOINT DISEASE|RHEUMATIC JOINT DISEASE (DISORDER)
C0409579|T047|14175009|SNOMEDCT_US|ARTHRITIS DUE TO RHEUMATIC FEVER|RHEUMATIC JOINT DISEASE (DISORDER)
C0409579|T047|14175009|SNOMEDCT_US|RHEUMATIC JOINT DISEASE |RHEUMATIC JOINT DISEASE (DISORDER)
C0409579|T047|14175009|SNOMEDCT_US|ARTICULAR RHEUMATIC FEVER, NOS|RHEUMATIC JOINT DISEASE (DISORDER)
C0409579|T047|14175009|SNOMEDCT_US|RHEUMATIC JOINT DISEASE, NOS|RHEUMATIC JOINT DISEASE (DISORDER)
C1304215|T047|402427003|SNOMEDCT_US|ACCELERATED RHEUMATOID NODULOSIS |ACCELERATED RHEUMATOID NODULOSIS (DISORDER)
C1304215|T047|402427003|SNOMEDCT_US|ACCELERATED RHEUMATOID NODULOSIS|ACCELERATED RHEUMATOID NODULOSIS (DISORDER)
C1997893|T047|429192004|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF FOOT|RHEUMATOID ARTHRITIS OF FOOT (DISORDER)
C1997893|T047|429192004|SNOMEDCT_US|RHEUMATOID ARTHRITIS OF FOOT |RHEUMATOID ARTHRITIS OF FOOT (DISORDER)
C1306838|T047|224729007|SNOMEDCT_US|PROLIFERATIVE ARTHRITIS|PROLIFERATIVE ARTHRITIS (DISORDER)
C1306838|T047|224729007|SNOMEDCT_US|PROLIFERATIVE ARTHRITIS |PROLIFERATIVE ARTHRITIS (DISORDER)
C1306838|T047|224729007|SNOMEDCT_US|PROLIFERATIVE ARTHRITIS, NOS|PROLIFERATIVE ARTHRITIS (DISORDER)
C0157913|T047|267887009|SNOMEDCT_US|RHEUMATOID ARTHRITIS AND OTHER INFLAMMATORY POLYARTHROPATHIES|RHEUMATOID ARTHRITIS AND OTHER INFLAMMATORY POLYARTHROPATHIES (DISORDER)
C0157913|T047|267887009|SNOMEDCT_US|RHEUMATOID ARTHRITIS AND OTHER INFLAMMATORY POLYARTHROPATHIES |RHEUMATOID ARTHRITIS AND OTHER INFLAMMATORY POLYARTHROPATHIES (DISORDER)
C0157919|T047|201812009|SNOMEDCT_US|OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHIES|OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY (DISORDER)
C0157919|T047|201812009|SNOMEDCT_US|OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY|OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY (DISORDER)
C0157919|T047|201812009|SNOMEDCT_US|INFLAMM POLYARTHROP NEC|OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY (DISORDER)
C0157919|T047|201812009|SNOMEDCT_US|OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY |OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY (DISORDER)
C0157919|T047|201812009|SNOMEDCT_US|OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY NOS |OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY (DISORDER)
C0157919|T047|201812009|SNOMEDCT_US|OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY NOS|OTHER SPECIFIED INFLAMMATORY POLYARTHROPATHY (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|POLYARTHRITIS|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|POLYARTHRITIDES|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHY|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHIES|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|POLYARTHRITIS, UNSPECIFIED|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|POLYARTHRITIS |POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMM POLYARTHROP NOS|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHIES (M05-M14)|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHY NOS|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHY NOS |POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|POLYARTHRITIS |POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|POLYARTHRITIS NOS|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|[X]INFLAMMATORY POLYARTHROPATHIES |POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHY |POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|POLYARTHROPATHY NOS -INFLAMMAT|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|[X]INFLAMMATORY POLYARTHROPATHIES|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|POLYARTICULAR ARTHRITIS|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY ARTHRITIS OF MULTIPLE JOINTS|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|UNSPECIFIED INFLAMMATORY POLYARTHROPATHY|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHY, NOS|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|POLYARTHRITIS, NOS|POLYARTHRITIS (DISORDER)
C0162323|T047|41397009|SNOMEDCT_US|INFLAMMATORY POLYARTHROPATHY OR POLYARTHRITIS NOS|POLYARTHRITIS (DISORDER)
C0409667|T047|201803007|SNOMEDCT_US|JUVENILE CHRONIC POLYARTHRITIS|POLYARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0409667|T047|201803007|SNOMEDCT_US|POLYARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS |POLYARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0409667|T047|201803007|SNOMEDCT_US|JUVENILE CHRONIC POLYARTHRITIS |POLYARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0409667|T047|201803007|SNOMEDCT_US|POLYARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS|POLYARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0409667|T047|201803007|SNOMEDCT_US|POLYARTICULAR JUVENILE ARTHRITIS|POLYARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0409667|T047|201803007|SNOMEDCT_US|JUVENILE CHRONIC POLYARTHRITIS, NOS|POLYARTICULAR ONSET JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHRONIC POSTRHEUMATIC ARTHROPATHY|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD]|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHRONIC POSTRHEUMATIC ARTHROPATHY |CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHRONIC POSTRHEUMATIC ARTHROPATHY -RETIRED-|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHR POSTRHEUM ARTHRITIS|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|JACCOUD SYNDROME|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHRONIC POSTRHEUMATIC ARTHROPATHY [JACCOUD], UNSPECIFIED SITE|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHRONIC POSTRHEUMATIC ARTHROPATHY, UNSPECIFIED SITE|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHRONIC POSTRHEUMATIC ARTHROPATHY |CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|NON-DEFORMING EROSIVE ARTHROPATHY|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHRONIC POST RHEUMATIC ARTHROPATHY|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|JACCOUD'S ARTHROPATHY|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|JACCOUD'S SYNDROME|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|JACCOUD'S DISEASE|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|JACCOUD'S ARTHRITIS|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|CHRONIC POST - RHEUMATIC ARTHROPATHY|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|JACCOUD'S SYNDROME |CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|ARTHROPATHY; JACCOUD|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|JACCOUD; ARTHROPATHY|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C0152084|T047|123247007|SNOMEDCT_US|JACCOUD|CHRONIC POSTRHEUMATIC ARTHROPATHY (DISORDER)
C3469325|T047||SNOMEDCT_US|FELTY'S SYNDROME, SHOULDER
C3469325|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS FELTY'S SYNDROME SHOULDER
C3469325|T047||SNOMEDCT_US|FELTY'S SYNDROME OF SHOULDER 
C3469325|T047||SNOMEDCT_US|FELTY'S SYNDROME OF SHOULDER
C3469320|T047||SNOMEDCT_US|FELTY'S SYNDROME, ELBOW
C3469320|T047||SNOMEDCT_US|FELTY'S SYNDROME, UNSPECIFIED ELBOW
C3469320|T047||SNOMEDCT_US|FELTY'S SYNDROME OF ELBOW
C3469320|T047||SNOMEDCT_US|FELTY'S SYNDROME OF ELBOW 
C3469320|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS FELTY'S SYNDROME ELBOW
C3469326|T047||SNOMEDCT_US|FELTY'S SYNDROME, WRIST
C3469326|T047||SNOMEDCT_US|FELTY'S SYNDROME OF WRIST
C3469326|T047||SNOMEDCT_US|FELTY'S SYNDROME OF WRIST 
C3469326|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS FELTY'S SYNDROME WRIST
C0837511|T047||SNOMEDCT_US|FELTY'S SYNDROME, HAND
C0837511|T047||SNOMEDCT_US|FELTY'S SYNDROME, UNSPECIFIED HAND
C0837511|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS FELTY'S SYNDROME HAND
C0837511|T047||SNOMEDCT_US|FELTY'S SYNDROME OF HAND 
C0837511|T047||SNOMEDCT_US|FELTY'S SYNDROME OF HAND
C3469322|T047||SNOMEDCT_US|FELTY'S SYNDROME, HIP
C3469322|T047||SNOMEDCT_US|FELTY'S SYNDROME, UNSPECIFIED HIP
C3469322|T047||SNOMEDCT_US|FELTY'S SYNDROME OF HIP 
C3469322|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS FELTY'S SYNDROME HIP
C3469322|T047||SNOMEDCT_US|FELTY'S SYNDROME OF HIP
C3469323|T047||SNOMEDCT_US|FELTY'S SYNDROME, UNSPECIFIED KNEE
C3469323|T047||SNOMEDCT_US|FELTY'S SYNDROME, KNEE
C3469323|T047||SNOMEDCT_US|FELTY'S SYNDROME OF KNEE
C3469323|T047||SNOMEDCT_US|FELTY'S SYNDROME OF KNEE 
C3469323|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS FELTY'S SYNDROME KNEE
C0837514|T047||SNOMEDCT_US|FELTY'S SYNDROME, ANKLE AND FOOT
C0837514|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS FELTY'S SYNDROME ANKLE AND FOOT
C0837514|T047||SNOMEDCT_US|FELTY'S SYNDROME OF ANKLE AND FOOT
C0837514|T047||SNOMEDCT_US|FELTY'S SYNDROME OF ANKLE AND FOOT 
C0837507|T047||SNOMEDCT_US|FELTY'S SYNDROME, MULTIPLE SITES
C0837507|T047||SNOMEDCT_US|FELTY'S SYNDROME OF MULTIPLE SITES 
C0837507|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS FELTY'S SYNDROME MULTIPLE SITES
C0837507|T047||SNOMEDCT_US|FELTY'S SYNDROME OF MULTIPLE SITES
C2936659|T047||SNOMEDCT_US|FAMILIAL FELTYS SYNDROME
C2936659|T047||SNOMEDCT_US|FELTY'S SYNDROME, FAMILIAL
C2936659|T047||SNOMEDCT_US|SYNDROME, FAMILIAL FELTY'S
C2936659|T047||SNOMEDCT_US|SYNDROME, FAMILIAL FELTY
C2936659|T047||SNOMEDCT_US|FELTY SYNDROME, FAMILIAL
C2936659|T047||SNOMEDCT_US|FAMILIAL FELTY'S SYNDROME
C2936659|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS, SPLENOMEGALY AND NEUTROPENIA
C2936659|T047||SNOMEDCT_US|FAMILIAL FELTY SYNDROME
C0234948|T047||SNOMEDCT_US|POLYARTHRITIS GENERALIZED
C0234948|T047||SNOMEDCT_US|POLYARTHRITIS GENERALISED
C0158024|T047||SNOMEDCT_US|UNSPECIFIED POLYARTHROPATHY OR POLYARTHRITIS INVOLVING OTHER SPECIFIED SITES
C0158024|T047||SNOMEDCT_US|POLYARTHRIT NOS-OTH SITE
C0158024|T047||SNOMEDCT_US|UNSPECIFIED POLYARTHROPATHY OR POLYARTHRITIS, OTHER SPECIFIED SITES
C0856585|T047||SNOMEDCT_US|POLYARTHROPATHY (EXCL RHEUMATOID ARTHRITIS)
C0856585|T047||SNOMEDCT_US|POLYARTHROPATHY (EXCLUDING RHEUMATOID ARTHRITIS)
C0018099|T047|90560007|SNOMEDCT_US|GOUT|GOUT (DISORDER)
C0018099|T047|90560007|SNOMEDCT_US|GOUT, UNSPECIFIED|GOUT (DISORDER)
C0018099|T047|90560007|SNOMEDCT_US|GOUT |GOUT (DISORDER)
C0018099|T047|90560007|SNOMEDCT_US|GOUT NOS|GOUT (DISORDER)
C0018099|T047|90560007|SNOMEDCT_US|GOUT [DISEASE/FINDING]|GOUT (DISORDER)
C0018099|T047|90560007|SNOMEDCT_US|GOUTS|GOUT (DISORDER)
C0018099|T047|90560007|SNOMEDCT_US|GOUT NOS |GOUT (DISORDER)
C0018099|T047|90560007|SNOMEDCT_US|GOUT |GOUT (DISORDER)
C0018099|T047|90560007|SNOMEDCT_US|GOUT; IN|GOUT (DISORDER)
C0018099|T047|90560007|SNOMEDCT_US|GOUT, NOS|GOUT (DISORDER)
C0494904|T047||SNOMEDCT_US|OTHER ARTHRITIS
C0409848|T047|201675001|SNOMEDCT_US|OTHER CRYSTAL ARTHROPATHIES|OTHER CRYSTAL ARTHROPATHIES OF UNSPECIFIED SITE (DISORDER)
C0409848|T047|201675001|SNOMEDCT_US|OTHER CRYSTAL ARTHROPATHY NOS |OTHER CRYSTAL ARTHROPATHIES OF UNSPECIFIED SITE (DISORDER)
C0409848|T047|201675001|SNOMEDCT_US|OTHER CRYSTAL ARTHROPATHIES |OTHER CRYSTAL ARTHROPATHIES OF UNSPECIFIED SITE (DISORDER)
C0409848|T047|201675001|SNOMEDCT_US|OTHER CRYSTAL ARTHROPATHIES OF UNSPECIFIED SITE |OTHER CRYSTAL ARTHROPATHIES OF UNSPECIFIED SITE (DISORDER)
C0409848|T047|201675001|SNOMEDCT_US|OTHER CRYSTAL ARTHROPATHY NOS|OTHER CRYSTAL ARTHROPATHIES OF UNSPECIFIED SITE (DISORDER)
C0409848|T047|201675001|SNOMEDCT_US|OTHER CRYSTAL ARTHROPATHIES OF UNSPECIFIED SITE|OTHER CRYSTAL ARTHROPATHIES OF UNSPECIFIED SITE (DISORDER)
C0494897|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS
C0694515|T047||SNOMEDCT_US|PSORIATIC AND ENTEROPATHIC ARTHROPATHIES
C0694516|T047||SNOMEDCT_US|JUVENILE ARTHRITIS IN DISEASES CLASSIFIED ELSEWHERE
C0694517|T047||SNOMEDCT_US|ARTHROPATHIES IN OTHER DISEASES CLASSIFIED ELSEWHERE
C2889385|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR, UNSPECIFIED
C2889385|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR
C2889493|T047||SNOMEDCT_US|ENTEROPATHIC ARTHROPATHIES
C2889493|T047||SNOMEDCT_US|ENTEROPATHIC ARTHROPATHY 
C2889493|T047||SNOMEDCT_US|ENTEROPATHIC ARTHROPATHY
C2919482|T047|445345005|SNOMEDCT_US|RS3PE - REMITTING SERONEGATIVE SYMMETRIC SYNOVITIS WITH PITTING EDEMA|RS3PE - REMITTING SERONEGATIVE SYMMETRIC SYNOVITIS WITH PITTING EDEMA
C2919482|T047|445345005|SNOMEDCT_US|REMITTING SERONEGATIVE SYMMETRICAL SYNOVITIS WITH PITTING EDEMA |RS3PE - REMITTING SERONEGATIVE SYMMETRIC SYNOVITIS WITH PITTING EDEMA
C2919482|T047|445345005|SNOMEDCT_US|RELAPSING SERONEGATIVE SYMMETRICAL SYNOVITIS WITH PITTING OEDEMA|RS3PE - REMITTING SERONEGATIVE SYMMETRIC SYNOVITIS WITH PITTING EDEMA
C2919482|T047|445345005|SNOMEDCT_US|RS3PE - REMITTING SERONEGATIVE SYMMETRIC SYNOVITIS WITH PITTING OEDEMA|RS3PE - REMITTING SERONEGATIVE SYMMETRIC SYNOVITIS WITH PITTING EDEMA
C2919482|T047|445345005|SNOMEDCT_US|REMITTING SERONEGATIVE SYMMETRICAL SYNOVITIS WITH PITTING EDEMA|RS3PE - REMITTING SERONEGATIVE SYMMETRIC SYNOVITIS WITH PITTING EDEMA
C2919482|T047|445345005|SNOMEDCT_US|REMITTING SERONEGATIVE SYMMETRICAL SYNOVITIS WITH PITTING OEDEMA|RS3PE - REMITTING SERONEGATIVE SYMMETRIC SYNOVITIS WITH PITTING EDEMA
C2919482|T047|445345005|SNOMEDCT_US|RELAPSING SERONEGATIVE SYMMETRICAL SYNOVITIS WITH PITTING EDEMA|RS3PE - REMITTING SERONEGATIVE SYMMETRIC SYNOVITIS WITH PITTING EDEMA
C2083208|T047||SNOMEDCT_US|POLYARTHRITIS OF MULTIPLE SITES 
C2083208|T047||SNOMEDCT_US|POLYARTHRITIS OF MULTIPLE SITES
C0268108|T047|68451005|SNOMEDCT_US|CHRONIC GOUT|CHRONIC GOUTY ARTHRITIS (DISORDER)
C0268108|T047|68451005|SNOMEDCT_US|GOUTY ARTHROPATHY CHRONIC |CHRONIC GOUTY ARTHRITIS (DISORDER)
C0268108|T047|68451005|SNOMEDCT_US|GOUTY ARTHROPATHY CHRONIC|CHRONIC GOUTY ARTHRITIS (DISORDER)
C0268108|T047|68451005|SNOMEDCT_US|CHRONIC GOUT |CHRONIC GOUTY ARTHRITIS (DISORDER)
C0268108|T047|68451005|SNOMEDCT_US|GOUT CHRONIC|CHRONIC GOUTY ARTHRITIS (DISORDER)
C0268108|T047|68451005|SNOMEDCT_US|CHRONIC GOUTY ARTHRITIS|CHRONIC GOUTY ARTHRITIS (DISORDER)
C0268108|T047|68451005|SNOMEDCT_US|CHRONIC GOUTY ARTHRITIS |CHRONIC GOUTY ARTHRITIS (DISORDER)
C2103075|T047||SNOMEDCT_US|AXIAL POLYARTICULAR INFLAMMATION 
C2103075|T047||SNOMEDCT_US|AXIAL POLYARTICULAR INFLAMMATION
C3495373|T047||SNOMEDCT_US|ARTHRITIS OF MULTIPLE SITES
C3495373|T047||SNOMEDCT_US|ARTHRITIS MULTIPLE SITES
C3495373|T047||SNOMEDCT_US|ARTHRITIS MULTIPLE SITES 
C0263721|T047|6211002|SNOMEDCT_US|POLYARTHRITIS ASSOCIATED WITH DISORDER CLASSIFIED ELSEWHERE|POLYARTHRITIS ASSOCIATED WITH ANOTHER DISORDER (DISORDER)
C0263721|T047|6211002|SNOMEDCT_US|POLYARTHRITIS ASSOCIATED WITH ANOTHER DISORDER |POLYARTHRITIS ASSOCIATED WITH ANOTHER DISORDER (DISORDER)
C0263721|T047|6211002|SNOMEDCT_US|POLYARTHRITIS ASSOCIATED WITH ANOTHER DISORDER|POLYARTHRITIS ASSOCIATED WITH ANOTHER DISORDER (DISORDER)
C1290689|T047|109663009|SNOMEDCT_US|ARTHRITIS OF TEMPOROMANDIBULAR JOINT AS PART OF POLYARTHRITIS |SYSTEMIC ARTHRITIS INCLUDING TEMPOROMANDIBULAR JOINT
C1290689|T047|109663009|SNOMEDCT_US|ARTHRITIS OF TEMPOROMANDIBULAR JOINT AS PART OF POLYARTHRITIS|SYSTEMIC ARTHRITIS INCLUDING TEMPOROMANDIBULAR JOINT
C1290689|T047|109663009|SNOMEDCT_US|SYSTEMIC ARTHRITIS INCLUDING TEMPOROMANDIBULAR JOINT|SYSTEMIC ARTHRITIS INCLUDING TEMPOROMANDIBULAR JOINT
C0409668|T047|239799007|SNOMEDCT_US|EARLY ONSET POLYARTICULAR JUVENILE CHRONIC ARTHRITIS|EARLY ONSET POLYARTICULAR JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0409668|T047|239799007|SNOMEDCT_US|EARLY ONSET POLYARTICULAR JUVENILE CHRONIC ARTHRITIS |EARLY ONSET POLYARTICULAR JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0263739|T047|1961000|SNOMEDCT_US|POLYARTICULAR JCA|CHRONIC POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0263739|T047|1961000|SNOMEDCT_US|POLYARTICULAR JUVENILE CHRONIC RA|CHRONIC POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0263739|T047|1961000|SNOMEDCT_US|CHRONIC POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS|CHRONIC POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0263739|T047|1961000|SNOMEDCT_US|CHRONIC POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS |CHRONIC POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0409669|T047|239800006|SNOMEDCT_US|LATE ONSET POLYARTICULAR JUVENILE CHRONIC ARTHRITIS|LATE ONSET POLYARTICULAR JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0409669|T047|239800006|SNOMEDCT_US|LATE ONSET POLYARTICULAR JUVENILE CHRONIC ARTHRITIS |LATE ONSET POLYARTICULAR JUVENILE CHRONIC ARTHRITIS (DISORDER)
C0409702|T047|239819001|SNOMEDCT_US|UNDIFFERENTIATED INFLAMMATORY OLIGOARTHRITIS|UNDIFFERENTIATED INFLAMMATORY OLIGOARTHRITIS (DISORDER)
C0409702|T047|239819001|SNOMEDCT_US|UNDIFFERENTIATED INFLAMMATORY OLIGOARTHRITIS |UNDIFFERENTIATED INFLAMMATORY OLIGOARTHRITIS (DISORDER)
C0263733|T047|44221002|SNOMEDCT_US|IDIOPATHIC POLYARTHRITIS|IDIOPATHIC POLYARTHRITIS (DISORDER)
C0263733|T047|44221002|SNOMEDCT_US|IDIOPATHIC POLYARTHRITIS |IDIOPATHIC POLYARTHRITIS (DISORDER)
C0311284|T047|190801003|SNOMEDCT_US|LIPOID DERMATOARTHRITIS|MULTICENTRIC RETICULOHISTIOCYTOSIS (DISORDER)
C0311284|T047|190801003|SNOMEDCT_US|LIPOID METABOLISM DISORDER LIPOID DERMATOARTHRITIS|MULTICENTRIC RETICULOHISTIOCYTOSIS (DISORDER)
C0311284|T047|190801003|SNOMEDCT_US|LIPOID DERMATOARTHRITIS |MULTICENTRIC RETICULOHISTIOCYTOSIS (DISORDER)
C0311284|T047|190801003|SNOMEDCT_US|MULTICENTRIC RETICULOHISTIOCYTOSIS|MULTICENTRIC RETICULOHISTIOCYTOSIS (DISORDER)
C0311284|T047|190801003|SNOMEDCT_US|MULTICENTRIC RETICULOHISTIOCYTOSIS |MULTICENTRIC RETICULOHISTIOCYTOSIS (DISORDER)
C0311284|T047|190801003|SNOMEDCT_US|NICOLAU-BALUS SYNDROME|MULTICENTRIC RETICULOHISTIOCYTOSIS (DISORDER)
C0311284|T047|190801003|SNOMEDCT_US|LIPOID DERMATOARTHRITIS |MULTICENTRIC RETICULOHISTIOCYTOSIS (DISORDER)
C1302753|T047|399964004|SNOMEDCT_US|CASE REPORTABLE, SO WILL LEAVE SINCE IT'S CLOSE|FIBROBLASTIC RHEUMATISM (DISORDER)
C1302753|T047|399964004|SNOMEDCT_US|FIBROBLASTIC RHEUMATISM|FIBROBLASTIC RHEUMATISM (DISORDER)
C1535016|T047|268053003|SNOMEDCT_US|POLYARTHROPATHY (& [INFLAMMATORY]) NOS |POLYARTHROPATHY (& [INFLAMMATORY]) NOS (DISORDER)
C1535016|T047|268053003|SNOMEDCT_US|POLYARTHROPATHY (& [INFLAMMATORY]) NOS|POLYARTHROPATHY (& [INFLAMMATORY]) NOS (DISORDER)
C3646092|T047||SNOMEDCT_US|SPONDYLOPATHY INFLAMMATORY MULTIPLE SITES SPINE
C3646092|T047||SNOMEDCT_US|SPONDYLOPATHY INFLAMMATORY MULTIPLE SITES SPINE 
C3687214|T047||SNOMEDCT_US|IMMUNE MEDIATED POLYARTHRITIS
C3687214|T047||SNOMEDCT_US|IMMUNE MEDIATED POLYARTHRITIS 
C1692871|T047|417373000|SNOMEDCT_US|INFLAMMATORY POLYARTHRITIS|INFLAMMATORY POLYARTHRITIS
C1692871|T047|417373000|SNOMEDCT_US|INFLAMMATORY; POLYARTHRITIS|INFLAMMATORY POLYARTHRITIS
C1692871|T047|417373000|SNOMEDCT_US|POLYARTHRITIS; INFLAMMATORY|INFLAMMATORY POLYARTHRITIS
C1692871|T047|417373000|SNOMEDCT_US|INFLAMMATORY POLYARTHRITIS, NOS|INFLAMMATORY POLYARTHRITIS
C1692872|T047|416956002|SNOMEDCT_US|UNDIFFERENTIATED INFLAMMATORY POLYARTHRITIS|UNDIFFERENTIATED INFLAMMATORY POLYARTHRITIS (DISORDER)
C1692872|T047|416956002|SNOMEDCT_US|UNDIFFERENTIATED INFLAMMATORY POLYARTHRITIS |UNDIFFERENTIATED INFLAMMATORY POLYARTHRITIS (DISORDER)
C0409252|T047|201972000|SNOMEDCT_US|ALLERGIC ARTHRITIS INVOLVING MULTIPLE SITES|ALLERGIC ARTHRITIS OF MULTIPLE SITES (DISORDER)
C0409252|T047|201972000|SNOMEDCT_US|ALLERGIC ARTHRITIS OF MULTIPLE SITES |ALLERGIC ARTHRITIS OF MULTIPLE SITES (DISORDER)
C0409252|T047|201972000|SNOMEDCT_US|ALLERGIC ARTHRITIS OF MULTIPLE SITES|ALLERGIC ARTHRITIS OF MULTIPLE SITES (DISORDER)
C0409252|T047|201972000|SNOMEDCT_US|ALLERG ARTHRITIS-MULT|ALLERGIC ARTHRITIS OF MULTIPLE SITES (DISORDER)
C0409252|T047|201972000|SNOMEDCT_US|ALLERGIC ARTHRITIS, MULTIPLE SITES|ALLERGIC ARTHRITIS OF MULTIPLE SITES (DISORDER)
C0409252|T047|201972000|SNOMEDCT_US|ALLERGIC ARTHRITIS OF MULTIPLE SITES |ALLERGIC ARTHRITIS OF MULTIPLE SITES (DISORDER)
C0157916|T047|75822003|SNOMEDCT_US|ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS|ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0157916|T047|75822003|SNOMEDCT_US|POLYART JUV RHEUM ARTHR|ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0157916|T047|75822003|SNOMEDCT_US|ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS |ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0157916|T047|75822003|SNOMEDCT_US|POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS, ACUTE|ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0157916|T047|75822003|SNOMEDCT_US|ACUTE POLYARTICULAR JUVENILE IDIOPATHIC ARTHRITIS |ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0157916|T047|75822003|SNOMEDCT_US|JUVENILE IDIOPATHIC ARTHRITIS, POLYARTICULAR ACUTE|ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0157916|T047|75822003|SNOMEDCT_US|ACUTE POLYARTICULAR JUVENILE IDIOPATHIC ARTHRITIS|ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0157916|T047|75822003|SNOMEDCT_US|ACUTE JUVENILE RHEUMATOID ARTHRITIS|ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C0157916|T047|75822003|SNOMEDCT_US|ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS [DUP] |ACUTE POLYARTICULAR JUVENILE RHEUMATOID ARTHRITIS (DISORDER)
C1827497|T047|422565003|SNOMEDCT_US|POST-INFECTIVE POLYARTHRITIS|REACTIVE ARTHRITIS OF MULTIPLE SITES
C1827497|T047|422565003|SNOMEDCT_US|REACTIVE ARTHRITIS OF MULTIPLE SITES|REACTIVE ARTHRITIS OF MULTIPLE SITES
C1827497|T047|422565003|SNOMEDCT_US|POST-INFECTIVE POLYARTHRITIS |REACTIVE ARTHRITIS OF MULTIPLE SITES
C0409703|T047|239821006|SNOMEDCT_US|SECONDARY INFLAMMATORY ARTHRITIS|SECONDARY INFLAMMATORY ARTHRITIS (DISORDER)
C0409703|T047|239821006|SNOMEDCT_US|SECONDARY INFLAMMATORY ARTHRITIS |SECONDARY INFLAMMATORY ARTHRITIS (DISORDER)
C2889165|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS
C2889165|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889165|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP SITE
C2889165|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS 
C2889179|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889179|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF HAND
C2889179|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP HAND
C2889179|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF HAND 
C2889182|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF HIP
C2889182|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF HIP 
C2889186|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF KNEE
C2889186|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF KNEE 
C2889195|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889195|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS MULT SITE
C2889195|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES 
C0264993|T047|399923009|SNOMEDCT_US|RHEUMATOID ARTERITIS|RHEUMATOID ARTERITIS (DISORDER)
C0264993|T047|399923009|SNOMEDCT_US|RHEUMATOID ARTERITIS |RHEUMATOID ARTERITIS (DISORDER)
C0343204|T047|239943002|SNOMEDCT_US|NECROTIZING RHEUMATOID VASCULITIS|NECROTIZING RHEUMATOID VASCULITIS (DISORDER)
C0343204|T047|239943002|SNOMEDCT_US|NECROTIZING RHEUMATOID VASCULITIS |NECROTIZING RHEUMATOID VASCULITIS (DISORDER)
C0343204|T047|239943002|SNOMEDCT_US|NECROTISING RHEUMATOID VASCULITIS|NECROTIZING RHEUMATOID VASCULITIS (DISORDER)
C0343204|T047|239943002|SNOMEDCT_US|NECROTIZING RHEUMATOID VASCULITIS |NECROTIZING RHEUMATOID VASCULITIS (DISORDER)
C0343202|T047|239941000|SNOMEDCT_US|NAILFOLD RHEUMATOID VASCULITIS|NAILFOLD RHEUMATOID VASCULITIS (DISORDER)
C0343202|T047|239941000|SNOMEDCT_US|NAILFOLD RHEUMATOID VASCULITIS |NAILFOLD RHEUMATOID VASCULITIS (DISORDER)
C0343203|T047|239942007|SNOMEDCT_US|SYSTEMIC RHEUMATOID VASCULITIS|SYSTEMIC RHEUMATOID VASCULITIS (DISORDER)
C0343203|T047|239942007|SNOMEDCT_US|SYSTEMIC RHEUMATOID VASCULITIS |SYSTEMIC RHEUMATOID VASCULITIS (DISORDER)
C1276120|T047|402433007|SNOMEDCT_US|BYWATER LESIONS|NAILFOLD/FINGER-PULP INFARCTS IN RHEUMATOID DISEASE (DISORDER)
C1276120|T047|402433007|SNOMEDCT_US|NAILFOLD/FINGER-PULP INFARCTS IN RHEUMATOID DISEASE |NAILFOLD/FINGER-PULP INFARCTS IN RHEUMATOID DISEASE (DISORDER)
C1276120|T047|402433007|SNOMEDCT_US|NAILFOLD/FINGER-PULP INFARCTS IN RHEUMATOID DISEASE|NAILFOLD/FINGER-PULP INFARCTS IN RHEUMATOID DISEASE (DISORDER)
C0392469|T047|28880005|SNOMEDCT_US|EDGE CASE - NOT A COMMONLY USED TERM BUT MORE LIKELY REFERS TO HEART LESIONS IN RHEUMATOID ARTHRITIS (RARE) THAN RHEUMATIC HEART DISEASE (IF IT WAS "RHEUMATIC CARDITIS" I WOULD ABSOLUTELY EXCLUDE)|RHEUMATOID CARDITIS (DISORDER)
C0392469|T047|28880005|SNOMEDCT_US|RHEUMATOID CARDITIS |RHEUMATOID CARDITIS (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|RHEUMATOID LUNG|RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|RHEUMATOID LUNG DISEASE|RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|RHEUMATOID LUNG |RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|RHEUMATOID LUNG DISEASE |RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|LUNG; RHEUMATOID (ETIOLOGY)|RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|LUNG; RHEUMATOID (MANIFESTATION)|RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH LUNG INVOLVEMENT (ETIOLOGY)|RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH LUNG INVOLVEMENT (MANIFESTATION)|RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|RHEUMATOID; LUNG (ETIOLOGY)|RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|RHEUMATOID; LUNG (MANIFESTATION)|RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH LUNG INVOLVEMENT (ETIOLOGY)|RHEUMATOID LUNG (DISORDER)
C0994344|T047|155621007|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH LUNG INVOLVEMENT (MANIFESTATION)|RHEUMATOID LUNG (DISORDER)
C0151379|T047|165839004|SNOMEDCT_US|RHEUMATOID FACTOR POSITIVE|RHEUMATOID FACTOR POSITIVE
C0151379|T047|165839004|SNOMEDCT_US|RHEUMATOID FACTOR POSITIVE |RHEUMATOID FACTOR POSITIVE
C3508972|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF SHOULDER
C3508972|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF SHOULDER 
C3508973|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF ELBOW
C3508973|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF ELBOW 
C3508974|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF WRIST
C3508974|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF WRIST 
C3508975|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF HAND
C3508975|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF HAND 
C3508976|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF HIP 
C3508976|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF HIP
C3508977|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF KNEE 
C3508977|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF KNEE
C3508978|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF ANKLE AND FOOT
C3508978|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF ANKLE AND FOOT 
C3508979|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF MULTIPLE SITES
C3508979|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE OF MULTIPLE SITES 
C3507373|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS 
C3507373|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS RF POSITIVE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0848642|T047||SNOMEDCT_US|SACROILITIS
C0837546|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0837546|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP SITE W INVOLV OF ORGANS AND SYSTEMS
C2889296|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889300|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889305|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0837541|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889313|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889317|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0837544|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0837537|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF MULTIPLE SITES WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C0837537|T047||SNOMEDCT_US|RHEU ARTHRITIS MULT SITE W INVOLV OF ORGANS AND SYSTEMS
C1384964|T047||SNOMEDCT_US|DISEASE (OR DISORDER); HEART, IN RHEUMATOID ARTHRITIS (ETIOLOGY)
C1384964|T047||SNOMEDCT_US|DISEASE (OR DISORDER); HEART, IN RHEUMATOID ARTHRITIS (MANIFESTATION)
C1388626|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH INVOLVEMENT OF ORGANS
C1388626|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH INVOLVEMENT OF ORGANS
C1388627|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH CARDITIS (ETIOLOGY)
C1388627|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH CARDITIS (MANIFESTATION)
C1388627|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH CARDITIS (ETIOLOGY)
C1388627|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH CARDITIS (MANIFESTATION)
C1388628|T047||SNOMEDCT_US|ENDOCARDITIS; RHEUMATOID ARTHRITIS (ETIOLOGY)
C1388628|T047||SNOMEDCT_US|ENDOCARDITIS; RHEUMATOID ARTHRITIS (MANIFESTATION)
C1388628|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS; ENDOCARDITIS (ETIOLOGY)
C1388628|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS; ENDOCARDITIS (MANIFESTATION)
C1388628|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH ENDOCARDITIS (ETIOLOGY)
C1388628|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH ENDOCARDITIS (MANIFESTATION)
C1388628|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH ENDOCARDITIS (ETIOLOGY)
C1388628|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH ENDOCARDITIS (MANIFESTATION)
C1388629|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH HEART INVOLVEMENT (ETIOLOGY)
C1388629|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH HEART INVOLVEMENT (MANIFESTATION)
C1388629|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH HEART INVOLVEMENT (ETIOLOGY)
C1388629|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH HEART INVOLVEMENT (MANIFESTATION)
C1388630|T047||SNOMEDCT_US|MYOCARDITIS; RHEUMATOID ARTHRITIS (ETIOLOGY)
C1388630|T047||SNOMEDCT_US|MYOCARDITIS; RHEUMATOID ARTHRITIS (MANIFESTATION)
C1388630|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS; MYOCARDITIS (ETIOLOGY)
C1388630|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS; MYOCARDITIS (MANIFESTATION)
C1388630|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH MYOCARDITIS (ETIOLOGY)
C1388630|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH MYOCARDITIS (MANIFESTATION)
C1388630|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH MYOCARDITIS (ETIOLOGY)
C1388630|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH MYOCARDITIS (MANIFESTATION)
C0343237|T047|193250002|SNOMEDCT_US|MYOPATHY DUE TO RHEUMATOID ARTHRITIS|MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0343237|T047|193250002|SNOMEDCT_US|MYOPATHY DUE TO RHEUMATOID ARTHRITIS |MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0343237|T047|193250002|SNOMEDCT_US|MYOPATHY; RHEUMATOID ARTHRITIS (ETIOLOGY)|MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0343237|T047|193250002|SNOMEDCT_US|MYOPATHY; RHEUMATOID ARTHRITIS (MANIFESTATION)|MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0343237|T047|193250002|SNOMEDCT_US|RHEUMATOID ARTHRITIS; MYOPATHY (ETIOLOGY)|MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0343237|T047|193250002|SNOMEDCT_US|RHEUMATOID ARTHRITIS; MYOPATHY (MANIFESTATION)|MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0343237|T047|193250002|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH MYOPATHY (ETIOLOGY)|MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0343237|T047|193250002|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH MYOPATHY (MANIFESTATION)|MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0343237|T047|193250002|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH MYOPATHY (ETIOLOGY)|MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0343237|T047|193250002|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH MYOPATHY (MANIFESTATION)|MYOPATHY DUE TO RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS |POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|POLYNEUROPATHY; RHEUMATOID ARTHRITIS (ETIOLOGY)|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|POLYNEUROPATHY; RHEUMATOID ARTHRITIS (MANIFESTATION)|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|RHEUMATOID ARTHRITIS; POLYNEUROPATHY (ETIOLOGY)|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|RHEUMATOID ARTHRITIS; POLYNEUROPATHY (MANIFESTATION)|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH POLYNEUROPATHY (ETIOLOGY)|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH POLYNEUROPATHY (MANIFESTATION)|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH POLYNEUROPATHY (ETIOLOGY)|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C0338555|T047|193180002|SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH POLYNEUROPATHY (MANIFESTATION)|POLYNEUROPATHY IN RHEUMATOID ARTHRITIS (DISORDER)
C1388632|T047||SNOMEDCT_US|RHEUMATOID; ARTHRITIS, WITH VISCERAL INVOLVEMENT
C1388632|T047||SNOMEDCT_US|ARTHRITIS; RHEUMATOID, WITH VISCERAL INVOLVEMENT
C1392056|T047||SNOMEDCT_US|50/50 IF THIS REFERS TO RHEUMATIC HEART DZ OR RA WITH CARDITIS
C1392056|T047||SNOMEDCT_US|CARDITIS; RHEUMATOID (MANIFESTATION)
C1392056|T047||SNOMEDCT_US|RHEUMATOID; CARDITIS (ETIOLOGY)
C1392056|T047||SNOMEDCT_US|RHEUMATOID; CARDITIS (MANIFESTATION)
C1399132|T047||SNOMEDCT_US|HEART; DISEASE, IN RHEUMATOID ARTHRITIS (ETIOLOGY)
C1399132|T047||SNOMEDCT_US|HEART; DISEASE, IN RHEUMATOID ARTHRITIS (MANIFESTATION)
C1404498|T047||SNOMEDCT_US|MYOCARDITIS; RHEUMATOID (ETIOLOGY)
C1404498|T047||SNOMEDCT_US|MYOCARDITIS; RHEUMATOID (MANIFESTATION)
C1404498|T047||SNOMEDCT_US|RHEUMATOID; MYOCARDITIS (ETIOLOGY)
C1404498|T047||SNOMEDCT_US|RHEUMATOID; MYOCARDITIS (MANIFESTATION)
C1406303|T047||SNOMEDCT_US|PERICARDITIS; RHEUMATOID (ETIOLOGY)
C1406303|T047||SNOMEDCT_US|PERICARDITIS; RHEUMATOID (MANIFESTATION)
C1406303|T047||SNOMEDCT_US|RHEUMATOID; PERICARDITIS (ETIOLOGY)
C1406303|T047||SNOMEDCT_US|RHEUMATOID; PERICARDITIS (MANIFESTATION)
C2889120|T047||SNOMEDCT_US|FELTY'S SYNDROME, RIGHT HAND
C2889121|T047||SNOMEDCT_US|FELTY'S SYNDROME, LEFT HAND
C2889129|T047||SNOMEDCT_US|FELTY'S SYNDROME, RIGHT ANKLE AND FOOT
C2889130|T047||SNOMEDCT_US|FELTY'S SYNDROME, LEFT ANKLE AND FOOT
C2889131|T047||SNOMEDCT_US|FELTY'S SYNDROME, UNSPECIFIED ANKLE AND FOOT
C2889310|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889310|T047||SNOMEDCT_US|RHEU ARTHRITIS OF RIGHT HAND W INVOLV OF ORGANS AND SYSTEMS
C2889311|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889311|T047||SNOMEDCT_US|RHEU ARTHRITIS OF LEFT HAND W INVOLV OF ORGANS AND SYSTEMS
C2889312|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889312|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP HAND W INVOLV OF ORGANS AND SYSTEMS
C2889322|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889322|T047||SNOMEDCT_US|RHEU ARTHRIT OF RIGHT ANK/FT W INVOLV OF ORGANS AND SYSTEMS
C2889323|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889323|T047||SNOMEDCT_US|RHEU ARTHRITIS OF LEFT ANK/FT W INVOLV OF ORGANS AND SYSTEMS
C2889324|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889324|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP ANK/FT W INVOLV OF ORGANS AND SYSTEMS
C2889132|T047|319841000119107|SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS (DISORDER)
C2889132|T047|319841000119107|SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS |RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS (DISORDER)
C1385071|T047||SNOMEDCT_US|DISEASE (OR DISORDER); LUNG, RHEUMATOID (DIFFUSE) (INTERSTITIAL) (ETIOLOGY)
C1385071|T047||SNOMEDCT_US|DISEASE (OR DISORDER); LUNG, RHEUMATOID (DIFFUSE) (INTERSTITIAL) (MANIFESTATION)
C1385071|T047||SNOMEDCT_US|LUNG; DISEASE, RHEUMATOID (DIFFUSE) (INTERSTITIAL) (ETIOLOGY)
C1385071|T047||SNOMEDCT_US|LUNG; DISEASE, RHEUMATOID (DIFFUSE) (INTERSTITIAL) (MANIFESTATION)
C1385163|T047||SNOMEDCT_US|DISEASE (OR DISORDER); RESPIRATORY, IN RHEUMATOID ARTHRITIS (ETIOLOGY)
C1385163|T047||SNOMEDCT_US|DISEASE (OR DISORDER); RESPIRATORY, IN RHEUMATOID ARTHRITIS (MANIFESTATION)
C1405189|T047||SNOMEDCT_US|PNEUMOCONIOSIS; RHEUMATOID (ETIOLOGY)
C1405189|T047||SNOMEDCT_US|PNEUMOCONIOSIS; RHEUMATOID (MANIFESTATION)
C1405189|T047||SNOMEDCT_US|RHEUMATOID; PNEUMOCONIOSIS (ETIOLOGY)
C1405189|T047||SNOMEDCT_US|RHEUMATOID; PNEUMOCONIOSIS (MANIFESTATION)
C1406187|T047||SNOMEDCT_US|RESPIRATORY; DISORDER, IN RHEUMATOID ARTHRITIS (ETIOLOGY)
C1406187|T047||SNOMEDCT_US|RESPIRATORY; DISORDER, IN RHEUMATOID ARTHRITIS (MANIFESTATION)
C3505955|T047||SNOMEDCT_US|RHEUMATOID NECROBIOTIC NODULE 
C3505955|T047||SNOMEDCT_US|RHEUMATOID NECROBIOTIC NODULE
C3505955|T047||SNOMEDCT_US|RHEUMATOID NODULE
C3505955|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS - NECROBIOTIC NODULE
C2889108|T047||SNOMEDCT_US|FELTY'S SYNDROME, RIGHT SHOULDER
C2889109|T047||SNOMEDCT_US|FELTY'S SYNDROME, LEFT SHOULDER
C2889110|T047||SNOMEDCT_US|FELTY'S SYNDROME, UNSPECIFIED SHOULDER
C2889112|T047||SNOMEDCT_US|FELTY'S SYNDROME, RIGHT ELBOW
C2889113|T047||SNOMEDCT_US|FELTY'S SYNDROME, LEFT ELBOW
C2889116|T047||SNOMEDCT_US|FELTY'S SYNDROME, RIGHT WRIST
C2889117|T047||SNOMEDCT_US|FELTY'S SYNDROME, LEFT WRIST
C2889118|T047||SNOMEDCT_US|FELTY'S SYNDROME, UNSPECIFIED WRIST
C2889122|T047||SNOMEDCT_US|FELTY'S SYNDROME, RIGHT HIP
C2889123|T047||SNOMEDCT_US|FELTY'S SYNDROME, LEFT HIP
C2889126|T047||SNOMEDCT_US|FELTY'S SYNDROME, RIGHT KNEE
C2889127|T047||SNOMEDCT_US|FELTY'S SYNDROME, LEFT KNEE
C2889133|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889133|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP SITE
C2889164|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889164|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS MULT SITE
C2889164|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES 
C2889135|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889135|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889136|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889136|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889137|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889137|T047||SNOMEDCT_US|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889139|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889139|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF R ELBOW
C2889140|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889140|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889141|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889141|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889144|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889144|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF R WRIST
C2889145|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889145|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889146|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889146|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889149|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889149|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889150|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889150|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT HAND
C2889151|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889151|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP HAND
C2889153|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889153|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889154|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889154|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT HIP
C2889156|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889156|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889157|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889157|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889158|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889158|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889161|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889161|T047||SNOMEDCT_US|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889162|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889162|T047||SNOMEDCT_US|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889163|T047||SNOMEDCT_US|RHEUMATOID LUNG DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889163|T047||SNOMEDCT_US|RHEU LUNG DISEASE W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889191|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889191|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT 
C2889166|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889166|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889167|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889167|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889170|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889170|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889171|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889171|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889172|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889172|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889175|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889175|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889176|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889176|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889177|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889177|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889180|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889180|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889181|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889183|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889184|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889185|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889185|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP HIP
C2889187|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889187|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889188|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889189|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889189|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889192|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889192|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889193|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889193|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889194|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889194|T047||SNOMEDCT_US|RHEUMATOID VASCULITIS W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889198|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889198|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP SITE
C2889199|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889199|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF SHOULDER 
C2889203|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889203|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF ELBOW 
C2889208|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF WRIST
C2889208|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF WRIST 
C2889213|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF HAND
C2889213|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF HAND 
C2889217|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF HIP
C2889217|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889217|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP HIP
C2889217|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF HIP 
C2889220|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF KNEE
C2889220|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF KNEE 
C2889225|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889225|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT 
C2889229|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889229|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS MULT SITE
C2889229|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES 
C2889200|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889200|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889201|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889201|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889202|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889202|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889204|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889204|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF R ELBOW
C2889205|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889205|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF L ELBOW
C2889206|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889206|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889209|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889209|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF R WRIST
C2889210|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889210|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF L WRIST
C2889211|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889211|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889214|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889214|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889215|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889215|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT HAND
C2889216|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889216|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP HAND
C2889218|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889218|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889219|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889219|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT HIP
C2889221|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889221|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889222|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889222|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889223|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889223|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889226|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889226|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889227|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889227|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889228|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889228|T047||SNOMEDCT_US|RHEU HEART DISEASE W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889231|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889231|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP SITE
C2889232|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889236|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889241|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF WRIST
C2889246|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF HAND
C2889246|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889246|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP HAND
C2889249|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF HIP
C2889253|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF KNEE
C2889258|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889262|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889262|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889233|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889233|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889234|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889234|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889235|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889235|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889237|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889238|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889239|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889239|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889242|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889243|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889244|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889244|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889247|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889248|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889250|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889251|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889252|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889252|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP HIP
C2889254|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889255|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889256|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889256|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889259|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889259|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889260|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889260|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889261|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889261|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889264|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SITE
C2889264|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP SITE
C2889265|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF SHOULDER
C2889271|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF ELBOW
C2889271|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW
C2889271|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP ELBOW
C2889273|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF WRIST
C2889278|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF HAND
C2889282|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF HIP
C2889286|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF KNEE
C2889291|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF ANKLE AND FOOT
C2889295|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF MULTIPLE SITES
C2889295|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY W RHEUMATOID ARTHRITIS MULT SITE
C2889266|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT SHOULDER
C2889266|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF R SHOULDER
C2889267|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT SHOULDER
C2889267|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF L SHOULDER
C2889268|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER
C2889268|T047||SNOMEDCT_US|RHEU POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP SHOULDER
C2889269|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889269|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT ELBOW
C2889270|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889270|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT ELBOW
C2889274|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889274|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT WRIST
C2889275|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889275|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT WRIST
C2889276|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST
C2889276|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP WRIST
C2889279|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889279|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT HAND
C2889280|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HAND
C2889280|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT HAND
C2889281|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HAND
C2889281|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP HAND
C2889283|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889283|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT HIP
C2889284|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT HIP
C2889284|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY W RHEUMATOID ARTHRITIS OF LEFT HIP
C2889285|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP
C2889285|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY W RHEUMATOID ARTHRITIS OF UNSP HIP
C2889287|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889287|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT KNEE
C2889288|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889288|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT KNEE
C2889289|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE
C2889289|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP KNEE
C2889292|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF RIGHT ANKLE AND FOOT
C2889292|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF RIGHT ANK/FT
C2889293|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF LEFT ANKLE AND FOOT
C2889293|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF LEFT ANK/FT
C2889294|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS OF UNSPECIFIED ANKLE AND FOOT
C2889294|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROP W RHEUMATOID ARTHRITIS OF UNSP ANK/FT
C2889297|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889297|T047||SNOMEDCT_US|RHEU ARTHRITIS OF R SHOULDER W INVOLV OF ORGANS AND SYSTEMS
C2889298|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889298|T047||SNOMEDCT_US|RHEU ARTHRITIS OF L SHOULDER W INVOLV OF ORGANS AND SYSTEMS
C2889299|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED SHOULDER WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889299|T047||SNOMEDCT_US|RHEU ARTHRIT OF UNSP SHOULDER W INVOLV OF ORGANS AND SYSTEMS
C2889301|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889301|T047||SNOMEDCT_US|RHEU ARTHRITIS OF R ELBOW W INVOLV OF ORGANS AND SYSTEMS
C2889302|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889302|T047||SNOMEDCT_US|RHEU ARTHRITIS OF L ELBOW W INVOLV OF ORGANS AND SYSTEMS
C2889303|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED ELBOW WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889303|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP ELBOW W INVOLV OF ORGANS AND SYSTEMS
C2889306|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889306|T047||SNOMEDCT_US|RHEU ARTHRITIS OF R WRIST W INVOLV OF ORGANS AND SYSTEMS
C2889307|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889307|T047||SNOMEDCT_US|RHEU ARTHRITIS OF L WRIST W INVOLV OF ORGANS AND SYSTEMS
C2889308|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED WRIST WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889308|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP WRIST W INVOLV OF ORGANS AND SYSTEMS
C2889314|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889314|T047||SNOMEDCT_US|RHEU ARTHRITIS OF RIGHT HIP W INVOLV OF ORGANS AND SYSTEMS
C2889315|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889315|T047||SNOMEDCT_US|RHEU ARTHRITIS OF LEFT HIP W INVOLV OF ORGANS AND SYSTEMS
C2889316|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED HIP WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889316|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP HIP W INVOLV OF ORGANS AND SYSTEMS
C2889318|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF RIGHT KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889318|T047||SNOMEDCT_US|RHEU ARTHRITIS OF RIGHT KNEE W INVOLV OF ORGANS AND SYSTEMS
C2889319|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF LEFT KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889319|T047||SNOMEDCT_US|RHEU ARTHRITIS OF LEFT KNEE W INVOLV OF ORGANS AND SYSTEMS
C2889320|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS OF UNSPECIFIED KNEE WITH INVOLVEMENT OF OTHER ORGANS AND SYSTEMS
C2889320|T047||SNOMEDCT_US|RHEU ARTHRITIS OF UNSP KNEE W INVOLV OF ORGANS AND SYSTEMS
C2889326|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SITE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889326|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF UNSP SITE W/O ORG/SYS INVOLV
C2889327|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889331|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889335|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889339|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889343|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889347|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889351|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889355|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF MULTIPLE SITES WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889355|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR MULT SITE W/O ORG/SYS INVOLV
C2889328|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889328|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF R SHOULDER W/O ORG/SYS INVOLV
C2889329|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889329|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF L SHOULDER W/O ORG/SYS INVOLV
C2889330|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SHOULDER WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889330|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF UNSP SHLDR W/O ORG/SYS INVOLV
C2889332|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889332|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF R ELBOW W/O ORG/SYS INVOLV
C2889333|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889333|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF L ELBOW W/O ORG/SYS INVOLV
C2889334|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ELBOW WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889334|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF UNSP ELBOW W/O ORG/SYS INVOLV
C2889336|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889336|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF R WRIST W/O ORG/SYS INVOLV
C2889337|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889337|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF L WRIST W/O ORG/SYS INVOLV
C2889338|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED WRIST WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889338|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF UNSP WRIST W/O ORG/SYS INVOLV
C2889340|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889340|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF R HAND W/O ORG/SYS INVOLV
C2889341|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889341|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF LEFT HAND W/O ORG/SYS INVOLV
C2889342|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HAND WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889342|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF UNSP HAND W/O ORG/SYS INVOLV
C2889344|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889344|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF RIGHT HIP W/O ORG/SYS INVOLV
C2889345|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889345|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF LEFT HIP W/O ORG/SYS INVOLV
C2889346|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HIP WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889346|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF UNSP HIP W/O ORG/SYS INVOLV
C2889348|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889348|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF R KNEE W/O ORG/SYS INVOLV
C2889349|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889349|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF LEFT KNEE W/O ORG/SYS INVOLV
C2889350|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED KNEE WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889350|T047||SNOMEDCT_US|RHEU ARTHRITIS W RHEU FACTOR OF UNSP KNEE W/O ORG/SYS INVOLV
C2889352|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889352|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FCTR OF RIGHT ANK/FT W/O ORG/SYS INVOLV
C2889353|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889353|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF LEFT ANK/FT W/O ORG/SYS INVOLV
C2889354|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ANKLE AND FOOT WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
C2889354|T047||SNOMEDCT_US|RHEU ARTHRIT W RHEU FACTOR OF UNSP ANK/FT W/O ORG/SYS INVOLV
C2889356|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR
C2889356|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SITE
C2889356|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP SITE
C2889357|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF SHOULDER
C2889361|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF ELBOW
C2889365|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF WRIST
C2889371|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF HAND
C2889371|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HAND
C2889371|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP HAND
C2889372|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF HIP
C2889376|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF KNEE
C2889380|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF ANKLE AND FOOT
C2889384|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF MULTIPLE SITES
C2889384|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR MULT SITE
C2889358|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT SHOULDER
C2889358|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF R SHOULDER
C2889359|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT SHOULDER
C2889359|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF L SHOULDER
C2889360|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED SHOULDER
C2889360|T047||SNOMEDCT_US|OTH RHEU ARTHRITIS W RHEUMATOID FACTOR OF UNSP SHOULDER
C2889362|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ELBOW
C2889362|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT ELBOW
C2889363|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ELBOW
C2889363|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF LEFT ELBOW
C2889364|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ELBOW
C2889364|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF UNSP ELBOW
C2889366|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT WRIST
C2889366|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT WRIST
C2889367|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT WRIST
C2889367|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF LEFT WRIST
C2889368|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED WRIST
C2889368|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF UNSP WRIST
C2889369|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HAND
C2889369|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT HAND
C2889370|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HAND
C2889370|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HAND
C2889373|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HIP
C2889373|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT HIP
C2889374|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HIP
C2889374|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT HIP
C2889375|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED HIP
C2889375|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP HIP
C2889377|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT KNEE
C2889377|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT KNEE
C2889378|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT KNEE
C2889378|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT KNEE
C2889379|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED KNEE
C2889379|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSP KNEE
C2889381|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF RIGHT ANKLE AND FOOT
C2889381|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF RIGHT ANK/FT
C2889382|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF LEFT ANKLE AND FOOT
C2889382|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF LEFT ANK/FT
C2889383|T047||SNOMEDCT_US|OTHER RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR OF UNSPECIFIED ANKLE AND FOOT
C2889383|T047||SNOMEDCT_US|OTH RHEUMATOID ARTHRITIS W RHEUMATOID FACTOR OF UNSP ANK/FT
C2889197|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS
C2889197|T047||SNOMEDCT_US|RHEUMATOID HEART DISEASE WITH RHEUMATOID ARTHRITIS 
C2889230|T047||SNOMEDCT_US|RHEUMATOID MYOPATHY WITH RHEUMATOID ARTHRITIS
C2889263|T047||SNOMEDCT_US|RHEUMATOID POLYNEUROPATHY WITH RHEUMATOID ARTHRITIS
C2889325|T047||SNOMEDCT_US|RHEUMATOID ARTHRITIS WITH RHEUMATOID FACTOR WITHOUT ORGAN OR SYSTEMS INVOLVEMENT
