// CUI|TUI|Text|preferredTerm
C0201838|T059|Albumin
C0202202|T059|Protein
C0201850|T059|alkaline phosphatase|Alkaline phosphatase measurement
C0201836|T059|ALT|Alanine aminotransferase measurement
C0201899|T059|AST|Aspartate aminotransferase measurement
C0201913|T059|bilirubin|Bilirubin, total measurement
C0036808|T059|Bilirubin, Indirect
C0858048|T059|Bilirubin, Direct
C0201973|T059|Total CK
C0523584|T059|CK-MB|Creatine kinase MB measurement
C0523584|T059|CKMB|Creatine kinase MB measurement
C0023508|T060|white count|White Blood Cell Count procedure
C0201803|T059|osmolality|Osmolality Measurement
C0017564|T060|GFR|Glomerular Filtration Rate
C0588466|T059|RBC, UA|Red blood cells urine (lab test)
C0000010|T059|WBC, UA|White blood cells urine (lab test)
C0201837|T201|A/G Ratio|Albumin/Globulin ratio
C0373670|T059|Lipase|Lipase measurement
C0033707|T059|Protime|Prothrombin time assay
C0525032|T059|INR|International Normalized Ratio
C1443182|T059|Calc|Calculated (procedure)
C00337443|T059|sodium|Sodium measurement
C00202194|T059|potassium|Potassium measurement
C00003074|T201|Anion Gap
C00202230|T059|TSH|Thyroid stimulating hormone measurement
C01171408|T059|LDL/HDL|High density/low density lipoprotein ratio measurement
C00518015|T059|hemoglobin|Hemoglobin measurement
C00032181|T059|platelet count|Platelet Count measurement
C00018935|T059|hematocrit|Hematocrit procedure
C00201657|T059|CRP|C-reactive protein measurement
C01535922|T059|procalcitonin|Procalcitonin measurement
C00202115|T059|lactate|Lactic acid measurement
C00202225|T059|free T4|T4 free measurement
C00201934|T059|cardiac enzymes|Cardiac enzymes measurement
C00337438|T059|glucose|Glucose measurement
C00201802|T059|specific gravity|Specific gravity measurement
C00200635|T059|lymphocytes|Lymphocyte Count measurement
C00005845|T059|BUN|Blood urea nitrogen measurement
C00201975|T059|creatinine|Creatinine measurement
C01305866|T060|weight|Weighing patient
C01305855|T201|BMI|Body mass index
000|T034|ALBUMIN [G/DL] IN SER/PLAS
3255-7|T034|Fibrinogen PPP-mCnc
14979-9|T034|aPTT Time PPP
3173-2|T034|aPTT Time Bld
34714-6|T034|INR Bld
6301-6|T034|INR PPP
5902-2|T034|PT Time PPP
3184-9|T034|ACT Time Bld
2276-4|T034|Ferritin SerPl-mCnc
2498-4|T034|Iron SerPl-mCnc
2500-7|T034|TIBC SerPl-mCnc
2501-5|T034|UIBC SerPl-mCnc
2571-8|T034|Trigl SerPl-mCnc
2085-9|T034|HDLc SerPl-mCnc
2093-3|T034|Cholest SerPl-mCnc
43396-1|T034|NonHDLc SerPl-mCnc
9830-1|T034|Cholest/HDLc SerPl-mRto
11054-4|T034|LDLc/HDLc SerPl-mRto
13457-7|T034|LDLc SerPl Calc-mCnc
18262-6|T034|LDLc SerPl Direct Assay-mCnc
2089-1|T034|LDLc SerPl-mCnc
13458-5|T034|VLDLc SerPl Calc-mCnc
2091-7|T034|VLDLc SerPl-mCnc
10834-0|T034|Globulin Ser Calc-mCnc
2336-6|T034|Globulin Ser-mCnc
1988-5|T034|CRP SerPl-mCnc
2458-8|T034|IgA Ser-mCnc
2465-3|T034|IgG Ser-mCnc
2472-9|T034|IgM Ser-mCnc
14338-8|T034|Prealb SerPl-mCnc
14957-5|T034|Microalbumin Ur-mCnc
14959-1|T034|Microalbumin/Creat Ur-mRto
1751-7|T034|Albumin SerPl-mCnc
1759-0|T034|Albumin/Glob SerPl-mRto
1959-6|T034|HCO3 Bld-sCnc
2823-3|T034|Potassium SerPl-sCnc
6298-4|T034|Potassium Bld-sCnc
2947-0|T034|Sodium Bld-sCnc
2951-2|T034|Sodium SerPl-sCnc
2069-3|T034|Chloride Bld-sCnc
2075-0|T034|Chloride SerPl-sCnc
10466-1|T034|Anion Gap3 SerPl-sCnc
33037-3|T034|Anion Gap SerPl-sCnc
1798-8|T034|Amylase SerPl-cCnc
3040-3|T034|Lipase SerPl-cCnc
2532-0|T034|LDH SerPl-cCnc
1742-6|T034|ALT SerPl-cCnc
6768-6|T034|ALP SerPl-cCnc
1920-8|T034|AST SerPl-cCnc
2157-6|T034|CK SerPl-cCnc
13969-1|T034|CK MB SerPl-mCnc
20569-0|T034|CK MB CFr SerPl
49136-5|T034|CK MB SerPl-Rto
2324-2|T034|GGT SerPl-cCnc
1989-3|T034|25(OH)D3 SerPl-mCnc
2132-9|T034|Vit B12 SerPl-mCnc
2284-8|T034|Folate SerPl-mCnc
2243-4|T034|Estradiol SerPl-mCnc
2986-8|T034|Testost SerPl-mCnc
19080-1|T034|HCG SerPl-aCnc
2106-3|T034|HCG Preg Ur Ql
2731-8|T034|PTH-Intact SerPl-mCnc
2842-3|T034|Prolactin SerPl-mCnc
11579-0|T034|TSH SerPl DL<=0.05 mIU/L-aCnc
11580-8|T034|TSH SerPl DL<=0.005 mIU/L-aCnc
3016-3|T034|TSH SerPl-aCnc
15067-2|T034|FSH SerPl-aCnc
10501-5|T034|LH SerPl-aCnc
3024-7|T034|T4 Free SerPl-mCnc
32215-6|T034|FTI SerPl-aCnc
3026-2|T034|T4 SerPl-mCnc
3050-2|T034|T3RU NFr SerPl
3051-0|T034|T3Free SerPl-mCnc
3053-6|T034|T3 SerPl-mCnc
1968-7|T034|Bilirub Direct SerPl-mCnc
1971-1|T034|Bilirub Indirect SerPl-mCnc
1975-2|T034|Bilirub SerPl-mCnc
1978-6|T034|Bilirub Ur-mCnc
3107-0|T034|Urobilinogen Ur-mCnc
5818-0|T034|Urobilinogen Ur Ql Strip
2161-8|T034|Creat Ur-mCnc
2160-0|T034|Creat SerPl-mCnc
38483-4|T034|Creat Bld-mCnc
3094-0|T034|BUN SerPl-mCnc
3097-3|T034|BUN/Creat SerPl-mRto
6299-2|T034|BUN Bld-mCnc
2965-2|T034|Sp Gr Ur
2349-9|T034|Glucose Ur Ql
27353-2|T034|Est. average glucose Bld gHb Est-mCnc
2339-0|T034|Glucose Bld-mCnc
2345-7|T034|Glucose SerPl-mCnc
2713-6|T034|SaO2% from pO2 Bld
11556-8|T034|pO2 Bld
2703-7|T034|pO2 BldA
11558-4|T034|pH Bld
2753-2|T034|pH SerPl
2744-1|T034|pH BldA
11557-6|T034|pCO2 Bld
2028-9|T034|CO2 SerPl-sCnc
20565-8|T034|CO2 Bld-sCnc
2019-8|T034|pCO2 BldA
11555-0|T034|Base excess Bld-sCnc
3084-1|T034|Urate SerPl-mCnc
10839-9|T034|Troponin I SerPl-mCnc
6598-7|T034|Troponin T SerPl-mCnc
30934-4|T034|BNP SerPl-mCnc
2857-1|T034|PSA SerPl-mCnc
2777-1|T034|Phosphate SerPl-mCnc
19123-9|T034|Magnesium SerPl-mCnc
2601-3|T034|Magnesium SerPl-sCnc
29265-6|T034|Calcium Album cor SerPl-sCnc
1994-3|T034|Ca-I Bld-sCnc
1995-0|T034|Ca-I SerPl-sCnc
2514-8|T034|Ketones Ur Ql Strip
33903-6|T034|Ketones Ur Ql
3390-2|T034|Benzodiaz Ur Ql
3377-9|T034|Barbiturates Ur Ql
18282-4|T034|Cannabinoids Ur Ql Scn
19659-2|T034|PCP Ur Ql Scn
3349-8|T034|Amphetamines Ur Ql
3879-4|T034|Opiates Ur Ql
3393-6|T034|BZE Ur Ql
11253-2|T034|Tacrolimus Bld-mCnc
5671-3|T034|Lead Bld-mCnc
56598-6|T034|EBV EA IgM Ser EIA-aCnc
5334-8|T034|RUBV IgG Ser EIA-aCnc
30167-1|T034|HPV I/H Risk 1 DNA Cervix Ql bDNA
48345-3|T034|HIV 1+O+2 Ab SerPl Ql
48346-1|T034|HIV 1+O+2 Ab SerPl-aCnc
5195-3|T034|HBV surface Ag Ser Ql
5196-1|T034|HBV surface Ag Ser Ql EIA
51656-7|T034|HCV Ab s/co Fld-Rto
5198-7|T034|HCV Ab Ser EIA-aCnc
21613-5|T034|C trach DNA XXX Ql PCR
42931-6|T034|C trach rRNA Ur Ql PCR
43304-5|T034|C trach rRNA XXX Ql PCR
50387-0|T034|C trach rRNA Cervix Ql PCR
53925-4|T034|C trach rRNA Urth Ql PCR
20507-0|T034|RPR Ser Ql
24111-7|T034|N gonorrhoea DNA XXX Ql PCR
43305-2|T034|N gonorrhoea rRNA XXX Ql PCR
50388-8|T034|N gonorrhoea rRNA Cervix Ql PCR
53927-0|T034|N gonorrhoea rRNA Urth Ql PCR
60256-5|T034|N gonorrhoea rRNA Ur Ql PCR
600-7|T034|Bacteria Bld Cult
624-7|T034|Bacteria Spt Resp Cult
630-4|T034|Bacteria Ur Cult
634-6|T034|Bacteria XXX Aerobe Cult
6462-6|T034|Bacteria Wnd Cult
6463-4|T034|Bacteria XXX Cult
10701-1|T034|O+P Stl Conc
35691-5|T034|Other microorganism DNA XXX Ql PCR
664-3|T034|Gram Stn XXX
30313-1|T034|Hgb BldA-mCnc
718-7|T034|Hgb Bld-mCnc
11282-1|T034|Total Cells Counted Bld
20570-8|T034|Hct VFr Bld
31100-1|T034|Hct VFr Bld Imped
4544-3|T034|Hct VFr Bld Auto
30341-2|T034|ESR Bld Qn
4537-7|T034|ESR Bld Qn Westrgrn
774-0|T034|Ovalocytes Bld Ql Smear
15150-6|T034|Anisocytosis Bld Ql Auto
702-1|T034|Anisocytosis Bld Ql Smear
15198-5|T034|Macrocytes Bld Ql Auto
738-5|T034|Macrocytes Bld Ql Smear
15199-3|T034|Microcytes Bld Ql Auto
741-9|T034|Microcytes Bld Ql Smear
18314-5|T034|Morphology Bld-Imp
10378-8|T034|Polychromasia Bld Ql Smear
15180-3|T034|Hypochromia Bld Ql Auto
728-6|T034|Hypochromia Bld Ql Smear
11125-2|T034|Plat morph Bld
6742-1|T034|RBC morph Bld
735-1|T034|Variant Lymphs NFr Bld Manual
26474-7|T034|Lymphocytes # Bld
26478-8|T034|Lymphocytes NFr Bld
731-0|T034|Lymphocytes # Bld Auto
736-9|T034|Lymphocytes NFr Bld Auto
737-7|T034|Lymphocytes NFr Bld Manual
769-0|T034|Neuts Seg NFr Bld Manual
26507-4|T034|Neuts Band # Bld
26508-2|T034|Neuts Band NFr Bld
764-1|T034|Neuts Band NFr Bld Manual
26499-4|T034|Neutrophils # Bld
26511-6|T034|Neutrophils NFr Bld
751-8|T034|Neutrophils # Bld Auto
770-8|T034|Neutrophils NFr Bld Auto
26444-0|T034|Basophils # Bld
30180-4|T034|Basophils NFr Bld
704-7|T034|Basophils # Bld Auto
706-2|T034|Basophils NFr Bld Auto
707-0|T034|Basophils NFr Bld Manual
26449-9|T034|Eosinophil # Bld
26450-7|T034|Eosinophil NFr Bld
711-2|T034|Eosinophil # Bld Auto
713-8|T034|Eosinophil NFr Bld Auto
714-6|T034|Eosinophil NFr Bld Manual
26464-8|T034|WBC # Bld
6690-2|T034|WBC # Bld Auto
30405-5|T034|WBC # Ur
26484-6|T034|Monocytes # Bld
26485-3|T034|Monocytes NFr Bld
5905-5|T034|Monocytes NFr Bld Auto
742-7|T034|Monocytes # Bld Auto
744-3|T034|Monocytes NFr Bld Manual
32623-1|T034|PMV Bld Auto
26515-7|T034|Platelet # Bld
777-3|T034|Platelet # Bld Auto
9317-9|T034|Platelet Bld Ql Smear
4679-7|T034|Retics/100 RBC NFr
789-8|T034|RBC # Bld Auto
798-9|T034|RBC # Ur Auto
17856-6|T034|Hgb A1c MFr Bld HPLC
4548-4|T034|Hgb A1c MFr Bld
30428-7|T034|MCV RBC
787-2|T034|MCV RBC Auto
785-6|T034|MCH RBC Qn Auto
786-4|T034|MCHC RBC Auto-mCnc
21000-5|T034|RDW RBC Auto
788-0|T034|RDW RBC Auto-Rto
10331-7|T034|Rh Bld
883-9|T034|ABO Group Bld
925-8|T034|Bld Prod Disposition BPU
933-2|T034|Bld Prod Typ BPU
934-0|T034|BPU ID
1003-3|T034|IAT Comp-Sp Reag SerPl Ql
1250-0|T034|Maj XM SerPl-Imp
882-1|T034|ABO+Rh Gp Bld
890-4|T034|Bld gp Ab Scn SerPl Ql
11572-5|T034|Rheumatoid fact Ser-aCnc
8061-4|T034|ANA Ser Ql
13362-9|T034|Collect duration Time Ur
19244-3|T034|Character Ur
31208-2|T034|Specimen source XXX
5767-9|T034|Appearance Ur
5778-6|T034|Color Ur
25162-9|T034|Hyaline Casts UrnS Ql Micro
5796-8|T034|Hyaline Casts #/area UrnS LPF
9842-6|T034|Casts #/area UrnS LPF
5769-5|T034|Bacteria #/area UrnS HPF
20453-7|T034|Epi Cells UrnS Ql Micro
5787-7|T034|Epi Cells #/area UrnS HPF
11277-1|T034|Squamous #/area UrnS HPF
12258-0|T034|Squamous UrnS Ql Micro
13945-1|T034|RBC #/area UrnS HPF
20409-9|T034|RBC # Ur Strip
33051-4|T034|RBC Ur Ql
5808-1|T034|RBC # UrnS HPF
20408-1|T034|WBC # Ur Strip
5821-4|T034|WBC #/area UrnS HPF
12454-5|T034|Amorph Urate Cry UrnS Ql Micro
8247-9|T034|Mucous Threads UrnS Ql Micro
5770-3|T034|Bilirub Ur Ql Strip
5792-7|T034|Glucose Ur Strip-mCnc
5794-3|T034|Hgb Ur Ql Strip
5797-6|T034|Ketones Ur Strip-mCnc
5799-2|T034|Leukocyte esterase Ur Ql Strip
5802-4|T034|Nitrite Ur Ql Strip
5803-2|T034|pH Ur Strip
5811-5|T034|Sp Gr Ur Strip
20454-5|T034|Prot Ur Ql Strip
2888-6|T034|Prot Ur-mCnc
5804-0|T034|Prot Ur Strip-mCnc
19161-9|T034|Urobilinogen Ur Strip-aCnc
20405-7|T034|Urobilinogen Ur Strip-mCnc
19763-2|T034|Specimen source Cvx/Vag Cyto
19764-0|T034|Stat of Adq Cvx/Vag Cyto-Imp
19767-3|T034|Cytologist Cvx/Vag Cyto
19769-9|T034|Pathologist Cvx/Vag Cyto
27045-4|T034|Microscopic Ur-Imp
47527-7|T034|Cytology Cvx/Vag Doc Thin Prep
19773-1|T034|Recom F/U Cvx/Vag Cyto
18928-2|T034|Gentamicin Susc Islt
20629-2|T034|Levofloxacin Susc Islt
23658-8|T034|Other Antibiotic Susc Islt
18998-5|T034|TMP SMX Susc Islt