C0001617|T121|N0000011309|NDFRT|ADRENAL CORTICOSTEROIDS|ADRENAL CORTEX HORMONES [CHEMICAL/INGREDIENT]
C0001947|T121|N0000029067|NDFRT|ALCOHOL DETERRENTS|[AD100] ALCOHOL DETERRENTS
C0002556|T121|N0000007853|NDFRT|AMINOGLYCOSIDES|AMINOGLYCOSIDES [CHEMICAL/INGREDIENT]
C0002667|T121|N0000007883|NDFRT|AMPHETAMINES|AMPHETAMINES [CHEMICAL/INGREDIENT]
C0002763|T121|N0000029152|NDFRT|CNS STIMULANTS|[CN800] CNS STIMULANTS
C0002771|T121|N0000029133|NDFRT|ANALGESICS|[CN100] ANALGESICS
C0002772|T121|N0000029136|NDFRT|OPIOID ANALGESICS|[CN101] OPIOID ANALGESICS
C0002932|T121|N0000029138|NDFRT|ANESTHETICS|[CN200] ANESTHETICS
C0003015|T121|N0000029130|NDFRT|ACE INHIBITORS|[CV800] ACE INHIBITORS
C0003138|T121|N0000029169|NDFRT|ANTACIDS|[GA100] ANTACIDS
C0003158|T121|N0000029099|NDFRT|ANTHELMINTICS|[AP200] ANTHELMINTICS
C0003191|T121|N0000029207|NDFRT|ANTIRHEUMATICS|[MS100] ANTIRHEUMATICS
C0003195|T121|N0000029121|NDFRT|ANTIARRHYTHMICS|[CV300] ANTIARRHYTHMICS
C0003216|T121|N0000029171|NDFRT|ANTIULCER AGENTS|[GA300] ANTIULCER AGENTS
C0003236|T121|N0000029093|NDFRT|ANTINEOPLASTIC ANTIBIOTICS|[AN200] ANTINEOPLASTIC ANTIBIOTICS
C0003280|T121|N0000029110|NDFRT|ANTICOAGULANTS|[BL110] ANTICOAGULANTS
C0003286|T121|N0000029145|NDFRT|ANTICONVULSANTS|[CN400] ANTICONVULSANTS
C0003289|T121|N0000029147|NDFRT|ANTIDEPRESSANTS|[CN600] ANTIDEPRESSANTS
C0003290|T121|N0000029148|NDFRT|TRICYCLIC ANTIDEPRESSANTS|[CN601] TRICYCLIC ANTIDEPRESSANTS
C0003292|T121|N0000029172|NDFRT|ANTIDIARRHEAL AGENTS|[GA208] ANTIDIARRHEAL AGENTS
C0003297|T121|N0000029175|NDFRT|ANTIEMETICS|[GA605] ANTIEMETICS
C0003308|T121|N0000029088|NDFRT|ANTIFUNGALS|[AM700] ANTIFUNGALS
C0003360|T121|N0000029071|NDFRT|ANTIHISTAMINES|[AH000] ANTIHISTAMINES
C0003367|T121||NDFRT|ANTILIPEMIC AGENTS
C0003374|T121|N0000029367|NDFRT|ANTIMALARIALS|[AP101] ANTIMALARIALS
C0003377|T121|N0000029094|NDFRT|ANTINEOPLASTICS,ANTIMETABOLITES|[AN300] ANTINEOPLASTICS,ANTIMETABOLITES
C0003392|T121|N0000029091|NDFRT|ANTINEOPLASTICS|[AN000] ANTINEOPLASTICS
C0003404|T121|N0000029097|NDFRT|ANTIPARASITICS|[AP000] ANTIPARASITICS
C0003405|T121|N0000029146|NDFRT|ANTIPARKINSON AGENTS|[CN500] ANTIPARKINSON AGENTS
C0003416|T121|N0000029098|NDFRT|ANTIPROTOZOALS|[AP100] ANTIPROTOZOALS
C0003419|T121|N0000029468|NDFRT|ANTIPYRETICS|[CN850] ANTIPYRETICS
C0003448|T121|N0000029084|NDFRT|ANTITUBERCULARS|[AM500] ANTITUBERCULARS
C0003451|T121|N0000029089|NDFRT|ANTIVIRALS|[AM800] ANTIVIRALS
C0003620|T121|N0000029396|NDFRT|APPETITE SUPPRESSANTS|[GA750] APPETITE SUPPRESSANTS
C0005367|T121|N0000007694|NDFRT|BICARBONATES|BICARBONATES [CHEMICAL/INGREDIENT]
C0006684|T121|N0000029119|NDFRT|CALCIUM CHANNEL BLOCKERS|[CV200] CALCIUM CHANNEL BLOCKERS
C0007220|T121|N0000029116|NDFRT|CARDIOVASCULAR MEDICATIONS|[CV000] CARDIOVASCULAR MEDICATIONS
C0007680|T121|N0000029132|NDFRT|CENTRAL NERVOUS SYSTEM MEDICATIONS|[CN000] CENTRAL NERVOUS SYSTEM MEDICATIONS
C0011427|T121|N0000011231|NDFRT|DENTIFRICES|DENTIFRICES [CHEMICAL/INGREDIENT]
C0011625|T121|N0000029154|NDFRT|DERMATOLOGICAL AGENTS|[DE000] DERMATOLOGICAL AGENTS
C0012237|T121|N0000029173|NDFRT|DIGESTANTS|[GA500] DIGESTANTS
C0012253|T121|N0000007534|NDFRT|DIGITALIS GLYCOSIDES|DIGITALIS GLYCOSIDES [CHEMICAL/INGREDIENT]
C0012798|T121|N0000029125|NDFRT|DIURETICS|[CV700] DIURETICS
C0012802|T121|N0000029126|NDFRT|THIAZIDES/RELATED DIURETICS|[CV701] THIAZIDES/RELATED DIURETICS
C0013973|T121|N0000029174|NDFRT|EMETICS|[GA600] EMETICS
C0013983|T121|N0000029370|NDFRT|EMOLLIENTS|[DE350] EMOLLIENTS
C0016018|T121|N0000029298|NDFRT|THROMBOLYTICS|[BL115] THROMBOLYTICS
C0017173|T121|N0000029168|NDFRT|GASTROINTESTINAL MEDICATIONS|[GA000] GASTROINTESTINAL MEDICATIONS
C0017710|T121|N0000175142|NDFRT|GLUCOCORTICOIDS|GLUCOCORTICOIDS [CHEMICAL/INGREDIENT]
C0018061|T121|N0000011199|NDFRT|GONADOTROPINS|GONADOTROPINS [CHEMICAL/INGREDIENT]
C0018100|T121|N0000029322|NDFRT|ANTIGOUT AGENTS|[MS400] ANTIGOUT AGENTS
C0018928|T121|N0000029113|NDFRT|BLOOD FORMATION PRODUCTS|[BL400] BLOOD FORMATION PRODUCTS
C0019006|T121|N0000029205|NDFRT|HEMODIALYSIS SOLUTIONS|[IR300] HEMODIALYSIS SOLUTIONS
C0019135|T121|N0000029111|NDFRT|HEPARIN ANTAGONISTS|[BL118] HEPARIN ANTAGONISTS
C0019590|T121|N0000029309|NDFRT|HISTAMINE ANTAGONISTS|[GA301] HISTAMINE ANTAGONISTS
C0020960|T121|N0000170864|NDFRT|IMMUNE SERUMS|IMMUNE SERA [CHEMICAL/INGREDIENT]
C0021027|T121|N0000007920|NDFRT|IMMUNOGLOBULINS|IMMUNOGLOBULINS [CHEMICAL/INGREDIENT]
C0021081|T121|N0000029316|NDFRT|IMMUNE SUPPRESSANTS|[IM600] IMMUNE SUPPRESSANTS
C0026160|T121|N0000029313|NDFRT|MINERALOCORTICOIDS|[HS052] MINERALOCORTICOIDS
C0026647|T121|N0000011404|NDFRT|MOUTHWASHES|MOUTHWASHES [CHEMICAL/INGREDIENT]
C0026698|T121|N0000029245|NDFRT|MUCOLYTICS|[RE400] MUCOLYTICS
C0027866|T121|N0000029362|NDFRT|NEUROMUSCULAR BLOCKING AGENTS|[MS300] NEUROMUSCULAR BLOCKING AGENTS
C0030094|T121|N0000029359|NDFRT|OXYTOCICS|[GU600] OXYTOCICS
C0030511|T121|N0000029107|NDFRT|PARASYMPATHOLYTICS|[AU350] PARASYMPATHOLYTICS
C0032016|T121|N0000011200|NDFRT|ANTERIOR PITUITARY|PITUITARY HORMONES, ANTERIOR [CHEMICAL/INGREDIENT]
C0032177|T121|N0000029299|NDFRT|PLATELET AGGREGATION INHIBITORS|[BL117] PLATELET AGGREGATION INHIBITORS
C0033306|T121|N0000029189|NDFRT|PROGESTINS|[HS800] PROGESTINS
C0033554|T121|N0000007706|NDFRT|PROSTAGLANDINS|PROSTAGLANDINS [CHEMICAL/INGREDIENT]
C0033613|T121|N0000029551|NDFRT|PROTECTIVE AGENTS|[AN700] PROTECTIVE AGENTS
C0036426|T121|N0000029285|NDFRT|SCLEROSING AGENTS|[CV600] SCLEROSING AGENTS
C0037250|T121|N0000029210|NDFRT|SKELETAL MUSCLE RELAXANTS|[MS200] SKELETAL MUSCLE RELAXANTS
C0039051|T121|N0000029105|NDFRT|SYMPATHOLYTICS|[AU200] SYMPATHOLYTICS
C0040125|T121|N0000029192|NDFRT|ANTITHYROID AGENTS|[HS852] ANTITHYROID AGENTS
C0040555|T121|N0000011209|NDFRT|TOXOIDS|TOXOIDS [CHEMICAL/INGREDIENT]
C0040615|T121|N0000029150|NDFRT|ANTIPSYCHOTICS|[CN700] ANTIPSYCHOTICS
C0042210|T121|N0000011210|NDFRT|VACCINES|VACCINES [CHEMICAL/INGREDIENT]
C0042398|T121|N0000029213|NDFRT|DECONGESTANTS,NASAL|[NT100] DECONGESTANTS,NASAL
C0085824|T121|N0000029112|NDFRT|ANTIHEMORRHAGICS|[BL116] ANTIHEMORRHAGICS
C0242859|T121|N0000029220|NDFRT|CONTACT LENS SOLUTIONS|[OP400] CONTACT LENS SOLUTIONS
C0242903|T121|N0000029139|NDFRT|ANESTHETICS,INHALATION|[CN201] ANESTHETICS,INHALATION
C0242937|T121|N0000029135|NDFRT|NON-OPIOID ANALGESICS|[CN103] NON-OPIOID ANALGESICS
C0280049|T121|N0000029295|NDFRT|EXTENDED SPECTRUM PENICILLINS|[AM113] EXTENDED SPECTRUM PENICILLINS
C0282090|T121|N0000029395|NDFRT|LAXATIVES|[GA209] LAXATIVES,OTHER
C0282090|T121|N0000029395|NDFRT|LAXATIVES,OTHER|[GA209] LAXATIVES,OTHER
C0282532|T121|N0000029092|NDFRT|ANTINEOPLASTICS,ALKYLATING AGENTS|[AN100] ANTINEOPLASTICS,ALKYLATING AGENTS
C0301470|T121|N0000029393|NDFRT|STOOL SOFTENER|[GA205] STOOL SOFTENER
C0302213|T121|N0000029346|NDFRT|LITHIUM SALTS|[CN750] LITHIUM SALTS
C0304317|T121|N0000029077|NDFRT|CEPHALOSPORIN 1ST GENERATION|[AM115] CEPHALOSPORIN 1ST GENERATION
C0304320|T121|N0000029079|NDFRT|CEPHALOSPORIN 3RD GENERATION|[AM117] CEPHALOSPORIN 3RD GENERATION
C0304412|T121|N0000029311|NDFRT|ANTIMUSCARINICS/ANTISPASMODICS|[GA800] ANTIMUSCARINICS/ANTISPASMODICS
C0304412|T121|N0000029311|NDFRT|ANTIMUSCARINICS/ANTISPASMODICS|[GA800] ANTIMUSCARINICS/ANTISPASMODICS
C0304450|T121|N0000029345|NDFRT|ANESTHETIC ADJUNCTS|[CN205] ANESTHETIC ADJUNCTS
C0304550|T121|N0000029389|NDFRT|BULK-FORMING LAXATIVES|[GA201] BULK-FORMING LAXATIVES
C0304551|T121|N0000029390|NDFRT|HYPEROSMOTIC LAXATIVES|[GA202] HYPEROSMOTIC LAXATIVES
C0304553|T121|N0000029392|NDFRT|STIMULANT LAXATIVES|[GA204] STIMULANT LAXATIVES
C0304599|T121|N0000029100|NDFRT|PEDICULICIDES|[AP300] PEDICULICIDES
C0304812|T121|N0000029188|NDFRT|PITUITARY|[HS700] PITUITARY
C0304951|T121|N0000029467|NDFRT|DIAGNOSTIC ANTIGENS|[DX300] DIAGNOSTIC ANTIGENS
C0305072|T121|N0000029284|NDFRT|HEAVY METAL ANTAGONISTS|[AD300] HEAVY METAL ANTAGONISTS
C0350167|T121|N0000029427|NDFRT|ANTIHYPERTENSIVES,OTHER|[CV490] ANTIHYPERTENSIVES,OTHER
C0353714|T121|N0000029204|NDFRT|PERITONEAL DIALYSIS SOLUTIONS|[IR200] PERITONEAL DIALYSIS SOLUTIONS
C0354100|T121|N0000029127|NDFRT|LOOP DIURETICS|[CV702] LOOP DIURETICS
C0354764|T121|N0000029357|NDFRT|BRONCHODILATORS,ANTICHOLINERGIC|[RE105] BRONCHODILATORS,ANTICHOLINERGIC
C0355335|T121|N0000029397|NDFRT|CENTRALLY-ACTING APPETITE SUPPRESSANTS|[GA751] CENTRALLY-ACTING APPETITE SUPPRESSANTS
C0355614|T121|N0000029300|NDFRT|ANTIMIGRAINE AGENTS|[CN105] ANTIMIGRAINE AGENTS
C0355824|T121|N0000029294|NDFRT|PENICILLINASE-RESISTANT PENICILLINS|[AM112] PENICILLINASE-RESISTANT PENICILLINS
C0358514|T121|N0000029164|NDFRT|DIAGNOSTIC AGENTS|[DX000] DIAGNOSTIC AGENTS
C0358587|T121|N0000029380|NDFRT|ALUMINUM/MAGNESIUM CONTAINING ANTACIDS|[GA103] ALUMINUM/MAGNESIUM CONTAINING ANTACIDS
C0360048|T121|N0000029166|NDFRT|RADIOPHARMACEUTICALS,DIAGNOSTIC|[DX200] RADIOPHARMACEUTICALS,DIAGNOSTIC
C0361823|T121|N0000029554|NDFRT|CEPHALOSPORIN 4TH GENERATION|[AM118] CEPHALOSPORIN 4TH GENERATION
C0486441|T121|N0000029115|NDFRT|BLOOD PRODUCTS,OTHER|[BL900] BLOOD PRODUCTS,OTHER
C0595375|T121|N0000029068|NDFRT|CYANIDE ANTIDOTES|[AD200] CYANIDE ANTIDOTES
C0682895|T121|N0000029353|NDFRT|MISCELLANEOUS AGENTS|[XX000] MISCELLANEOUS AGENTS
C0718581|T121|N0000029334|NDFRT|ANTIHISTAMINE/DECONGESTANT|[RE501] ANTIHISTAMINE/DECONGESTANT
C0721844|T121|N0000029466|NDFRT|MULTIVITAMINS WITH MINERALS|[VT802] MULTIVITAMINS WITH MINERALS
C0724138|T121|N0000029261|NDFRT|ANALGESICS,URINARY|[GU100] ANALGESICS,URINARY
C0724804|T121|N0000029124|NDFRT|PERIPHERAL VASODILATORS|[CV500] PERIPHERAL VASODILATORS
C0731742|T121|N0000029351|NDFRT|CNS STIMULANTS,OTHER|[CN809] CNS STIMULANTS,OTHER
C0876271|T121|N0000029262|NDFRT|ANTISPASMODICS,URINARY|[GU200] ANTISPASMODICS,URINARY
C0876271|T121|N0000029262|NDFRT|ANTISPASMODICS,URINARY|[GU200] ANTISPASMODICS,URINARY
C0973578|T121|N0000029209|NDFRT|ANTIRHEUMATICS,OTHER|[MS190] ANTIRHEUMATICS,OTHER
C0973585|T121|N0000029216|NDFRT|OPHTHALMIC AGENTS|[OP000] OPHTHALMIC AGENTS
C0973601|T121|N0000029223|NDFRT|ANESTHETICS,TOPICAL OPHTHALMIC|[OP700] ANESTHETICS,TOPICAL OPHTHALMIC
C0973654|T121|N0000029257|NDFRT|ENTERAL NUTRITION|[TN200] ENTERAL NUTRITION
C0973669|T121|N0000029274|NDFRT|VITAMINS,OTHER|[VT900] VITAMINS,OTHER
C0991617|T121|N0000029231|NDFRT|OTIC AGENTS|[OT000] OTIC AGENTS
C1136254|T121|N0000029074|NDFRT|ANTIMICROBIALS|[AM000] ANTIMICROBIALS
C1322965|T121|N0000029229|NDFRT|DENTURE ADHESIVES|[OR400] DENTURE ADHESIVES
C1533693|T121|N0000183553|NDFRT|QUINOLONES|[AM400] QUINOLONES
C1579312|T121|N0000029194|NDFRT|IMMUNOLOGICAL AGENTS|[IM000] IMMUNOLOGICAL AGENTS
C1579313|T121|N0000029352|NDFRT|IMMUNE STIMULANTS|[IM700] IMMUNE STIMULANTS
C1579337|T121|N0000029293|NDFRT|PENICILLINS,AMINO DERIVATIVES|[AM111] PENICILLINS,AMINO DERIVATIVES
C1579362|T121|N0000029425|NDFRT|ANTIDEPRESSANTS,OTHER|[CN609] ANTIDEPRESSANTS,OTHER
C1579395|T121|N0000029253|NDFRT|THERAPEUTIC NUTRIENTS/MINERALS/ELECTROLYTES|[TN000] THERAPEUTIC NUTRIENTS/MINERALS/ELECTROLYTES
C1579396|T121|N0000029358|NDFRT|ELECTROLYTES/MINERALS|[TN400] ELECTROLYTES/MINERALS
C1579411|T121|N0000029096|NDFRT|ANTINEOPLASTIC,OTHER|[AN900] ANTINEOPLASTIC,OTHER
C1579431|T121|N0000029186|NDFRT|ANTIHYPOGLYCEMICS|[HS503] ANTIHYPOGLYCEMICS
C1579434|T121|N0000029109|NDFRT|BLOOD PRODUCTS/MODIFIERS/VOLUME EXPANDERS|[BL000] BLOOD PRODUCTS/MODIFIERS/VOLUME EXPANDERS
C1629497|T121|N0000029114|NDFRT|BLOOD DERIVATIVES|[BL500] BLOOD DERIVATIVES
C1744619|T121|N0000029082|NDFRT|TETRACYCLINES|[AM250] TETRACYCLINES
C1874023|T121|N0000029325|NDFRT|ADRENERGICS,TOPICAL OPHTHALMIC|[OP103] ADRENERGICS,TOPICAL OPHTHALMIC
C1874153|T121|N0000029337|NDFRT|ALPHA BLOCKERS/RELATED|[CV150] ALPHA BLOCKERS/RELATED
C1874163|T121|N0000029378|NDFRT|ALUMINUM CONTAINING ANTACIDS|[GA101] ALUMINUM CONTAINING ANTACIDS
C1874176|T121|N0000029379|NDFRT|ALUMINUM/CALCIUM/MAGNESIUM CONTAINING ANTACIDS|[GA102] ALUMINUM/CALCIUM/MAGNESIUM CONTAINING ANTACIDS
C1874177|T121|N0000029381|NDFRT|ALUMINUM/MAGNESIUM/SODIUM BICARBONATE CONTAINING ANTACIDS|[GA104] ALUMINUM/MAGNESIUM/SODIUM BICARBONATE CONTAINING ANTACIDS
C1874187|T121|N0000029433|NDFRT|AMINO ACIDS/PROTEINS|[TN500] AMINO ACIDS/PROTEINS
C1874188|T121|N0000029447|NDFRT|AMINO ACIDS/PROTEINS,ORAL|[TN503] AMINO ACIDS/PROTEINS,ORAL
C1874189|T121|N0000029448|NDFRT|AMINO ACIDS/PROTEINS,OTHER|[TN509] AMINO ACIDS/PROTEINS,OTHER
C1874190|T121|N0000029446|NDFRT|AMINO ACIDS/PROTEINS,PARENTERAL,WITH ADDED ELECTROLYTES|[TN502] AMINO ACIDS/PROTEINS,PARENTERAL,WITH ADDED ELECTROLYTES
C1874191|T121|N0000029432|NDFRT|AMINO ACIDS/PROTEINS,PARENTERAL,WITHOUT ADDED ELECTROLYTES|[TN501] AMINO ACIDS/PROTEINS,PARENTERAL,WITHOUT ADDED ELECTROLYTES
C1874222|T121|N0000029350|NDFRT|AMPHETAMINE LIKE STIMULANTS|[CN802] AMPHETAMINE LIKE STIMULANTS
C1874237|T121|N0000029372|NDFRT|ANALGESICS,TOPICAL|[DE650] ANALGESICS,TOPICAL
C1874238|T121|N0000029356|NDFRT|ANALGESICS,TOPICAL OTIC|[OT400] ANALGESICS,TOPICAL OTIC
C1874239|T121|N0000029179|NDFRT|ANDROGENS/ANABOLICS|[HS100] ANDROGENS/ANABOLICS
C1874240|T121|N0000029215|NDFRT|ANESTHETICS,MUCOSAL|[NT300] ANESTHETICS,MUCOSAL
C1874242|T121|N0000029550|NDFRT|ANGIOTENSIN II INHIBITOR|[CV805] ANGIOTENSIN II INHIBITOR
C1874245|T121|N0000029388|NDFRT|ANTACIDS,OTHER|[GA199] ANTACIDS,OTHER
C1874247|T121|N0000029155|NDFRT|ANTI-INFECTIVE,TOPICAL|[DE100] ANTI-INFECTIVE,TOPICAL
C1874248|T121|N0000029218|NDFRT|ANTI-INFECTIVE,TOPICAL OPHTHALMIC|[OP200] ANTI-INFECTIVE,TOPICAL OPHTHALMIC
C1874249|T121|N0000029406|NDFRT|ANTI-INFECTIVE,TOPICAL OPHTHALMIC,OTHER|[OP219] ANTI-INFECTIVE,TOPICAL OPHTHALMIC,OTHER
C1874250|T121|N0000029232|NDFRT|ANTI-INFECTIVE,TOPICAL OTIC|[OT100] ANTI-INFECTIVE,TOPICAL OTIC
C1874251|T121|N0000029369|NDFRT|ANTI-INFECTIVE,TOPICAL,OTHER|[DE109] ANTI-INFECTIVE,TOPICAL,OTHER
C1874252|T121|N0000029344|NDFRT|ANTI-INFECTIVE/ANTI-INFLAMMATORY COMBINATIONS,TOPICAL|[DE250] ANTI-INFECTIVE/ANTI-INFLAMMATORY COMBINATIONS,TOPICAL
C1874253|T121|N0000029340|NDFRT|ANTI-INFECTIVE/ANTI-INFLAMMATORY COMBINATIONS,TOPICAL OPHTHALMIC|[OP350] ANTI-INFECTIVE/ANTI-INFLAMMATORY COMBINATIONS,TOPICAL OPHTHALMIC
C1874254|T121|N0000029341|NDFRT|ANTI-INFECTIVE/ANTI-INFLAMMATORY COMBINATIONS,TOPICAL OTIC|[OT250] ANTI-INFECTIVE/ANTI-INFLAMMATORY COMBINATIONS,TOPICAL OTIC
C1874255|T121|N0000029090|NDFRT|ANTI-INFECTIVES,OTHER|[AM900] ANTI-INFECTIVES,OTHER
C1874256|T121|N0000029407|NDFRT|ANTI-INFECTIVES,TOPICAL OTIC OTHER|[OT109] ANTI-INFECTIVES,TOPICAL OTIC OTHER
C1874257|T121|N0000029263|NDFRT|ANTI-INFECTIVES,VAGINAL|[GU300] ANTI-INFECTIVES,VAGINAL
C1874258|T121|N0000029239|NDFRT|ANTI-INFLAMMATORIES,INHALATION|[RE101] ANTI-INFLAMMATORIES,INHALATION
C1874259|T121|N0000029214|NDFRT|ANTI-INFLAMMATORIES,NASAL|[NT200] ANTI-INFLAMMATORIES,NASAL
C1874260|T121|N0000029249|NDFRT|ANTI-INFLAMMATORIES,RECTAL|[RS100] ANTI-INFLAMMATORIES,RECTAL
C1874261|T121|N0000029219|NDFRT|ANTI-INFLAMMATORIES,TOPICAL OPHTHALMIC|[OP300] ANTI-INFLAMMATORIES,TOPICAL OPHTHALMIC
C1874262|T121|N0000029233|NDFRT|ANTI-INFLAMMATORIES,TOPICAL OTIC|[OT200] ANTI-INFLAMMATORIES,TOPICAL OTIC
C1874263|T121|N0000029156|NDFRT|ANTI-INFLAMMATORY,TOPICAL|[DE200] ANTI-INFLAMMATORY,TOPICAL
C1874264|T121|N0000029373|NDFRT|ANTIACNE AGENTS|[DE750] ANTIACNE AGENTS
C1874265|T121|N0000029374|NDFRT|ANTIACNE AGENTS,SYSTEMIC|[DE751] ANTIACNE AGENTS,SYSTEMIC
C1874266|T121|N0000029375|NDFRT|ANTIACNE AGENTS,TOPICAL|[DE752] ANTIACNE AGENTS,TOPICAL
C1874268|T121|N0000029553|NDFRT|ANTIASTHMA,ANTILEUKOTRIENES|[RE108] ANTIASTHMA,ANTILEUKOTRIENES
C1874269|T121|N0000029242|NDFRT|ANTIASTHMA,OTHER|[RE109] ANTIASTHMA,OTHER
C1874270|T121|N0000029238|NDFRT|ANTIASTHMA/BRONCHODILATORS|[RE100] ANTIASTHMA/BRONCHODILATORS
C1874271|T121|N0000029302|NDFRT|ANTIBACTERIAL,TOPICAL|[DE101] ANTIBACTERIAL,TOPICAL
C1874272|T121|N0000029327|NDFRT|ANTIBACTERIALS,TOPICAL OPHTHALMIC|[OP210] ANTIBACTERIALS,TOPICAL OPHTHALMIC
C1874273|T121|N0000029331|NDFRT|ANTIBACTERIALS,TOPICAL OTIC|[OT101] ANTIBACTERIALS,TOPICAL OTIC
C1874278|T121|N0000029066|NDFRT|ANTIDOTES,DETERRENTS AND POISON CONTROL|[AD000] ANTIDOTES,DETERRENTS AND POISON CONTROL
C1874279|T121|N0000029069|NDFRT|ANTIDOTES,DETERRENTS,AND POISON CONTROL EXCHANGE RESINS|[AD400] ANTIDOTES,DETERRENTS,AND POISON CONTROL EXCHANGE RESINS
C1874280|T121|N0000029070|NDFRT|ANTIDOTES/DETERRENTS,OTHER|[AD900] ANTIDOTES/DETERRENTS,OTHER
C1874281|T121|N0000029303|NDFRT|ANTIFUNGAL,TOPICAL|[DE102] ANTIFUNGAL,TOPICAL
C1874282|T121|N0000029328|NDFRT|ANTIFUNGALS,TOPICAL OPHTHALMIC|[OP220] ANTIFUNGALS,TOPICAL OPHTHALMIC
C1874283|T121|N0000029332|NDFRT|ANTIFUNGALS,TOPICAL OTIC|[OT102] ANTIFUNGALS,TOPICAL OTIC
C1874284|T121|N0000029339|NDFRT|ANTIGLAUCOMA COMBINATIONS,TOPICAL OPHTHALMIC|[OP105] ANTIGLAUCOMA COMBINATIONS,TOPICAL OPHTHALMIC
C1874285|T121|N0000029217|NDFRT|ANTIGLAUCOMA MEDICATIONS|[OP100] ANTIGLAUCOMA MEDICATIONS
C1874286|T121|N0000029405|NDFRT|ANTIGLAUCOMA,OTHER|[OP109] ANTIGLAUCOMA,OTHER
C1874288|T121|N0000029414|NDFRT|ANTIHISTAMINE/ANTITUSSIVE|[RE507] ANTIHISTAMINE/ANTITUSSIVE
C1874289|T121|N0000029342|NDFRT|ANTIHISTAMINE/ANTITUSSIVE/ANALGESIC|[RE509] ANTIHISTAMINE/ANTITUSSIVE/ANALGESIC
C1874290|T121|N0000029415|NDFRT|ANTIHISTAMINE/ANTITUSSIVE/EXPECTORANT|[RE508] ANTIHISTAMINE/ANTITUSSIVE/EXPECTORANT
C1874291|T121|N0000029335|NDFRT|ANTIHISTAMINE/DECONGESTANT/ANTITUSSIVE|[RE502] ANTIHISTAMINE/DECONGESTANT/ANTITUSSIVE
C1874292|T121|N0000029413|NDFRT|ANTIHISTAMINE/DECONGESTANT/ANTITUSSIVE/ANALGESIC|[RE506] ANTIHISTAMINE/DECONGESTANT/ANTITUSSIVE/ANALGESIC
C1874293|T121|N0000029411|NDFRT|ANTIHISTAMINE/DECONGESTANT/ANTITUSSIVE/EXPECTORANT|[RE504] ANTIHISTAMINE/DECONGESTANT/ANTITUSSIVE/EXPECTORANT
C1874294|T121|N0000029412|NDFRT|ANTIHISTAMINE/DECONGESTANT/ANTITUSSIVE/EXPECTORANT/ANALGESIC|[RE505] ANTIHISTAMINE/DECONGESTANT/ANTITUSSIVE/EXPECTORANT/ANALGESIC
C1874295|T121|N0000029410|NDFRT|ANTIHISTAMINE/DECONGESTANT/EXPECTORANT|[RE503] ANTIHISTAMINE/DECONGESTANT/EXPECTORANT
C1874296|T121|N0000029290|NDFRT|ANTIHISTAMINES,ALKYLAMINE|[AH104] ANTIHISTAMINES,ALKYLAMINE
C1874297|T121|N0000029364|NDFRT|ANTIHISTAMINES,BUTYROPHENONE|[AH106] ANTIHISTAMINES,BUTYROPHENONE
C1874298|T121|N0000029288|NDFRT|ANTIHISTAMINES,ETHANOLAMINE|[AH102] ANTIHISTAMINES,ETHANOLAMINE
C1874299|T121|N0000029289|NDFRT|ANTIHISTAMINES,ETHYLENEDIAMINE|[AH103] ANTIHISTAMINES,ETHYLENEDIAMINE
C1874300|T121|N0000029555|NDFRT|ANTIHISTAMINES,NASAL|[NT400] ANTIHISTAMINES,NASAL
C1874301|T121|N0000029073|NDFRT|ANTIHISTAMINES,OTHER|[AH109] ANTIHISTAMINES,OTHER
C1874302|T121|N0000029072|NDFRT|ANTIHISTAMINES,PHENOTHIAZINE|[AH100] ANTIHISTAMINES,PHENOTHIAZINE
C1874303|T121|N0000029291|NDFRT|ANTIHISTAMINES,PIPERAZINE|[AH105] ANTIHISTAMINES,PIPERAZINE
C1874304|T121|N0000029365|NDFRT|ANTIHISTAMINES,PIPERIDINE|[AH107] ANTIHISTAMINES,PIPERIDINE
C1874305|T121|N0000029123|NDFRT|ANTIHYPERTENSIVE COMBINATIONS|[CV400] ANTIHYPERTENSIVE COMBINATIONS
C1874306|T121|N0000029319|NDFRT|ANTIMALARIALS,ANTIRHEUMATIC|[MS130] ANTIMALARIALS,ANTIRHEUMATIC
C1874307|T121|N0000029401|NDFRT|ANTIMUSCARINIC/ANTIPASMODIC COMBINATIONS|[GA802] ANTIMUSCARINIC/ANTIPASMODIC COMBINATIONS
C1874308|T121|N0000029095|NDFRT|ANTINEOPLASTIC ADJUVANTS|[AN400] ANTINEOPLASTIC ADJUVANTS
C1874309|T121|N0000029297|NDFRT|ANTINEOPLASTIC HORMONES|[AN500] ANTINEOPLASTIC HORMONES
C1874310|T121|N0000029347|NDFRT|ANTINEOPLASTIC RADIOPHARMACEUTICALS|[AN600] ANTINEOPLASTIC RADIOPHARMACEUTICALS
C1874311|T121|N0000029160|NDFRT|ANTINEOPLASTIC,TOPICAL|[DE600] ANTINEOPLASTIC,TOPICAL
C1874312|T121|N0000029101|NDFRT|ANTIPARASITICS,OTHER|[AP900] ANTIPARASITICS,OTHER
C1874313|T121|N0000029368|NDFRT|ANTIPROTOZOALS,OTHER|[AP109] ANTIPROTOZOALS,OTHER
C1874314|T121|N0000029162|NDFRT|ANTIPSORIATIC|[DE800] ANTIPSORIATIC
C1874315|T121|N0000029376|NDFRT|ANTIPSORIATICS,SYSTEMIC|[DE810] ANTIPSORIATICS,SYSTEMIC
C1874316|T121|N0000029377|NDFRT|ANTIPSORIATICS,TOPICAL|[DE820] ANTIPSORIATICS,TOPICAL
C1874317|T121|N0000029426|NDFRT|ANTIPSYCHOTICS,OTHER|[CN709] ANTIPSYCHOTICS,OTHER
C1874321|T121|N0000029102|NDFRT|ANTISEPTICS/DISINFECTANTS|[AS000] ANTISEPTICS/DISINFECTANTS
C1874322|T121|N0000029430|NDFRT|ANTISPASMODICS,URINARY,OTHER|[GU209] ANTISPASMODICS,URINARY,OTHER
C1874323|T121|N0000029416|NDFRT|ANTITUSSIVE/ANTIMUSCARINIC|[RE510] ANTITUSSIVE/ANTIMUSCARINIC
C1874324|T121|N0000029417|NDFRT|ANTITUSSIVE/BRONCHODILATOR|[RE511] ANTITUSSIVE/BRONCHODILATOR
C1874325|T121|N0000029244|NDFRT|ANTITUSSIVES/EXPECTORANTS|[RE300] ANTITUSSIVES/EXPECTORANTS
C1874326|T121|N0000029429|NDFRT|ANTIULCER AGENTS,OTHER|[GA309] ANTIULCER AGENTS,OTHER
C1874327|T121|N0000029197|NDFRT|ANTIVENINS/ANTITOXINS|[IM300] ANTIVENINS/ANTITOXINS
C1874328|T121|N0000029301|NDFRT|ANTIVERTIGO AGENTS|[CN550] ANTIVERTIGO AGENTS
C1874329|T121|N0000029304|NDFRT|ANTIVIRAL,TOPICAL|[DE103] ANTIVIRAL,TOPICAL
C1874330|T121|N0000029329|NDFRT|ANTIVIRALS,TOPICAL OPHTHALMIC|[OP230] ANTIVIRALS,TOPICAL OPHTHALMIC
C1874331|T121|N0000029399|NDFRT|APPETITE SUPPRESSANTS,OTHER|[GA759] APPETITE SUPPRESSANTS,OTHER
C1874402|T121|N0000029108|NDFRT|AUTONOMIC AGENTS,OTHER|[AU900] AUTONOMIC AGENTS,OTHER
C1874403|T121|N0000029103|NDFRT|AUTONOMIC MEDICATIONS|[AU000] AUTONOMIC MEDICATIONS
C1874444|T121|N0000029286|NDFRT|BARBITURIC ACID DERIVATIVE ANESTHETICS|[CN202] BARBITURIC ACID DERIVATIVE ANESTHETICS
C1874445|T121|N0000029140|NDFRT|BARBITURIC ACID DERIVATIVE SEDATIVES/HYPNOTICS|[CN301] BARBITURIC ACID DERIVATIVE SEDATIVES/HYPNOTICS
C1874525|T121|N0000029144|NDFRT|BENZODIAZEPINE DERIVATIVE SEDATIVES/HYPNOTICS|[CN302] BENZODIAZEPINE DERIVATIVE SEDATIVES/HYPNOTICS
C1874540|T121|N0000029118|NDFRT|BETA BLOCKERS/RELATED|[CV100] BETA BLOCKERS/RELATED
C1874542|T121|N0000029404|NDFRT|BETA-BLOCKERS,SYSTEMIC OPHTHALMIC|[OP107] BETA-BLOCKERS,SYSTEMIC OPHTHALMIC
C1874543|T121|N0000029323|NDFRT|BETA-BLOCKERS,TOPICAL OPHTHALMIC|[OP101] BETA-BLOCKERS,TOPICAL OPHTHALMIC
C1874545|T121|N0000029366|NDFRT|BETA-LACTAMS ANTIMICROBIALS,OTHER|[AM119] BETA-LACTAMS ANTIMICROBIALS,OTHER
C1874587|T121|N0000029183|NDFRT|BLOOD GLUCOSE REGULATION AGENTS|[HS500] BLOOD GLUCOSE REGULATION AGENTS
C1874620|T121|N0000029240|NDFRT|BRONCHODILATORS,SYMPATHOMIMETIC,INHALATION|[RE102] BRONCHODILATORS,SYMPATHOMIMETIC,INHALATION
C1874621|T121|N0000029241|NDFRT|BRONCHODILATORS,SYMPATHOMIMETIC,ORAL|[RE103] BRONCHODILATORS,SYMPATHOMIMETIC,ORAL
C1874622|T121|N0000029333|NDFRT|BRONCHODILATORS,XANTHINE-DERIVATIVE|[RE104] BRONCHODILATORS,XANTHINE-DERIVATIVE
C1874624|T121|N0000029398|NDFRT|BULKING AGENT,APPETITE SUPPRESSANTS|[GA752] BULKING AGENT,APPETITE SUPPRESSANTS
C1874663|T121|N0000029382|NDFRT|CALCIUM CONTAINING ANTACIDS|[GA105] CALCIUM CONTAINING ANTACIDS
C1874677|T121|N0000029383|NDFRT|CALCIUM/MAGNESIUM CONTAINING ANTACIDS|[GA106] CALCIUM/MAGNESIUM CONTAINING ANTACIDS
C1874718|T121|N0000029394|NDFRT|CARBON DIOXIDE-RELEASING LAXATIVES|[GA206] CARBON DIOXIDE-RELEASING LAXATIVES
C1874722|T121|N0000029128|NDFRT|CARBONIC ANHYDRASE INHIBITOR DIURETICS|[CV703] CARBONIC ANHYDRASE INHIBITOR DIURETICS
C1874723|T121|N0000029326|NDFRT|CARBONIC ANHYDRASE INHIBITORS,SYSTEMIC OPHTHALMIC|[OP140] CARBONIC ANHYDRASE INHIBITORS,SYSTEMIC OPHTHALMIC
C1874728|T121|N0000029131|NDFRT|CARDIOVASCULAR AGENTS,OTHER|[CV900] CARDIOVASCULAR AGENTS,OTHER
C1874730|T121|N0000029226|NDFRT|CARIOSTATICS,TOPICAL|[OR100] CARIOSTATICS,TOPICAL
C1874766|T121|N0000029078|NDFRT|CEPHALOSPORIN 2ND GENERATION|[AM116] CEPHALOSPORIN 2ND GENERATION
C1874769|T121|N0000029234|NDFRT|CERUMINOLYTICS|[OT300] CERUMINOLYTICS
C1874882|T121|N0000029153|NDFRT|CNS MEDICATIONS,OTHER|[CN900] CNS MEDICATIONS,OTHER
C1874910|T121|N0000029246|NDFRT|COLD REMEDIES,COMBINATIONS|[RE500] COLD REMEDIES,COMBINATIONS
C1874911|T121|N0000029423|NDFRT|COLD REMEDIES,OTHER|[RE599] COLD REMEDIES,OTHER
C1874923|T121|N0000029180|NDFRT|CONTRACEPTIVES,SYSTEMIC|[HS200] CONTRACEPTIVES,SYSTEMIC
C1874924|T121|N0000029264|NDFRT|CONTRACEPTIVES,VAGINAL/TOPICAL|[GU400] CONTRACEPTIVES,VAGINAL/TOPICAL
C1874925|T121|N0000029635|NDFRT|CONTRAST MEDIA, OTHER|[DX109] CONTRAST MEDIA, OTHER
C1874949|T121|N0000029321|NDFRT|CYTOTOXICS,ANTIRHEUMATIC|[MS150] CYTOTOXICS,ANTIRHEUMATIC
C1874952|T121|N0000029418|NDFRT|DECONGESTANT/ANTITUSSIVE|[RE512] DECONGESTANT/ANTITUSSIVE
C1874953|T121|N0000029421|NDFRT|DECONGESTANT/ANTITUSSIVE/ANALGESIC|[RE515] DECONGESTANT/ANTITUSSIVE/ANALGESIC
C1874954|T121|N0000029419|NDFRT|DECONGESTANT/ANTITUSSIVE/EXPECTORANT|[RE513] DECONGESTANT/ANTITUSSIVE/EXPECTORANT
C1874955|T121|N0000029420|NDFRT|DECONGESTANT/ANTITUSSIVE/EXPECTORANT/ANALGESIC|[RE514] DECONGESTANT/ANTITUSSIVE/EXPECTORANT/ANALGESIC
C1874956|T121|N0000029422|NDFRT|DECONGESTANT/EXPECTORANT|[RE516] DECONGESTANT/EXPECTORANT
C1874957|T121|N0000029243|NDFRT|DECONGESTANTS,SYSTEMIC|[RE200] DECONGESTANTS,SYSTEMIC
C1874958|T121|N0000029355|NDFRT|DECONGESTANTS,TOPICAL OPHTHALMIC|[OP800] DECONGESTANTS,TOPICAL OPHTHALMIC
C1874965|T121|N0000029225|NDFRT|DENTAL AND ORAL AGENTS,TOPICAL|[OR000] DENTAL AND ORAL AGENTS,TOPICAL
C1874966|T121|N0000029330|NDFRT|DENTAL AND ORAL AGENTS,TOPICAL,OTHER|[OR900] DENTAL AND ORAL AGENTS,TOPICAL,OTHER
C1874967|T121|N0000029227|NDFRT|DENTAL PROTECTANTS|[OR200] DENTAL PROTECTANTS
C1874968|T121|N0000029371|NDFRT|DEODORANTS/ANTIPERSPIRANTS,TOPICAL|[DE450] DEODORANTS/ANTIPERSPIRANTS,TOPICAL
C1874969|T121|N0000029428|NDFRT|DERMATOLOGICALS,SYSTEMIC,OTHER|[DE890] DERMATOLOGICALS,SYSTEMIC,OTHER
C1874970|T121|N0000029163|NDFRT|DERMATOLOGICALS,TOPICAL OTHER|[DE900] DERMATOLOGICALS,TOPICAL OTHER
C1875013|T121|N0000029167|NDFRT|DIAGNOSTICS,OTHER|[DX900] DIAGNOSTICS,OTHER
C1875040|T121|N0000029338|NDFRT|DIURETICS,OTHER|[CV709] DIURETICS,OTHER
C1875099|T121|N0000029435|NDFRT|ELECTROLYTES/MINERALS,COMBINATIONS|[TN490] ELECTROLYTES/MINERALS,COMBINATIONS
C1875100|T121|N0000029434|NDFRT|ELECTROLYTES/MINERALS,OTHER|[TN499] ELECTROLYTES/MINERALS,OTHER
C1875123|T121|N0000029081|NDFRT|ERYTHROMYCINS/MACROLIDES|[AM200] ERYTHROMYCINS/MACROLIDES
C1875126|T121|N0000029265|NDFRT|ESTROGENS,VAGINAL|[GU500] ESTROGENS,VAGINAL
C1875146|T121|N0000029221|NDFRT|EYE WASHES/LUBRICANTS|[OP500] EYE WASHES/LUBRICANTS
C1875167|T121|N0000029450|NDFRT|FOLIC ACID/LEUCOVORIN|[VT102] FOLIC ACID/LEUCOVORIN
C1875178|T121|N0000029176|NDFRT|GASTRIC MEDICATIONS,OTHER|[GA900] GASTRIC MEDICATIONS,OTHER
C1875185|T121|N0000029141|NDFRT|GENERAL ANESTHETICS,OTHER|[CN203] GENERAL ANESTHETICS,OTHER
C1875186|T121|N0000029266|NDFRT|GENITO-URINARY AGENTS,OTHER|[GU900] GENITO-URINARY AGENTS,OTHER
C1875187|T121|N0000029260|NDFRT|GENITOURINARY MEDICATIONS|[GU000] GENITOURINARY MEDICATIONS
C1875221|T121|N0000029208|NDFRT|GOLD COMPOUNDS,ANTIRHEUMATIC|[MS160] GOLD COMPOUNDS,ANTIRHEUMATIC
C1875232|T121|N0000029552|NDFRT|H. PYLORI AGENTS|[GA303] H. PYLORI AGENTS
C1875239|T121|N0000029549|NDFRT|HEMORRHOIDAL PREPARATIONS WITH STEROID|[RS202] HEMORRHOIDAL PREPARATIONS WITH STEROID
C1875240|T121|N0000029548|NDFRT|HEMORRHOIDAL PREPARATIONS WITHOUT STEROID|[RS201] HEMORRHOIDAL PREPARATIONS WITHOUT STEROID
C1875241|T121|N0000029250|NDFRT|HEMORRHOIDAL PREPARATIONS,RECTAL|[RS200] HEMORRHOIDAL PREPARATIONS,RECTAL
C1875248|T121|N0000029634|NDFRT|HERBS/ALTERNATIVE THERAPIES|[HA000] HERBS/ALTERNATIVE THERAPIES
C1875254|T121|N0000029177|NDFRT|HORMONES/SYNTHETICS/MODIFIERS|[HS000] HORMONES/SYNTHETICS/MODIFIERS
C1875255|T121|N0000029193|NDFRT|HORMONES/SYNTHETICS/MODIFIERS,OTHER|[HS900] HORMONES/SYNTHETICS/MODIFIERS,OTHER
C1875291|T121|N0000029307|NDFRT|IMAGING AGENTS (IN VIVO) RADIOPHARMACEUTICALS|[DX201] IMAGING AGENTS (IN VIVO) RADIOPHARMACEUTICALS
C1875294|T121|N0000029200|NDFRT|IMMUNOLOGICAL AGENTS,OTHER|[IM900] IMMUNOLOGICAL AGENTS,OTHER
C1875299|T121|N0000029558|NDFRT|INTRAPLEURAL AGENTS,OTHER|[IP900] INTRAPLEURAL AGENTS,OTHER
C1875300|T121|N0000029556|NDFRT|INTRAPLEURAL MEDICATIONS|[IP000] INTRAPLEURAL MEDICATIONS
C1875301|T121|N0000029557|NDFRT|INTRAPLEURAL SCLEROSING AGENTS|[IP100] INTRAPLEURAL SCLEROSING AGENTS
C1875309|T121|N0000029573|NDFRT|INVEST ANTI-NEOPLASTIC BONE,CONNECTIVE TISSUE,SKIN,BREAST|[IN200] INVEST ANTI-NEOPLASTIC BONE,CONNECTIVE TISSUE,SKIN,BREAST
C1875310|T121|N0000029575|NDFRT|INVEST ANTI-NEOPLASTIC DIGESTIVE ORGANS,PERITONEUM|[IN220] INVEST ANTI-NEOPLASTIC DIGESTIVE ORGANS,PERITONEUM
C1875311|T121|N0000029579|NDFRT|INVEST ANTI-NEOPLASTIC DRUGS LIP,ORAL CAVITY AND PHARYNX|[IN260] INVEST ANTI-NEOPLASTIC DRUGS LIP,ORAL CAVITY AND PHARYNX
C1875312|T121|N0000029580|NDFRT|INVEST ANTI-NEOPLASTIC DRUGS LYMPHATIC AND HEMAPOIETIC TISSUE|[IN270] INVEST ANTI-NEOPLASTIC DRUGS LYMPHATIC AND HEMAPOIETIC TISSUE
C1875313|T121|N0000029623|NDFRT|INVEST DRUGS FOR DIALYSIS AND VOLUME/ELECTROLYTE SUPPORT|[IN880] INVEST DRUGS FOR DIALYSIS AND VOLUME/ELECTROLYTE SUPPORT
C1875314|T121|N0000029597|NDFRT|INVEST DRUGS FOR PSYCHOSIS AND POST TRAMATIC STRESS DISORDER|[IN570] INVEST DRUGS FOR PSYCHOSIS AND POST TRAMATIC STRESS DISORDER
C1875315|T121|N0000029612|NDFRT|INVEST DRUGS PSORIASIS,ECZEMA,NON-INFECTIOUS DERMATITIS|[IN700] INVEST DRUGS PSORIASIS,ECZEMA,NON-INFECTIOUS DERMATITIS
C1875316|T121|N0000029584|NDFRT|INVEST HEMATOLOGIC DEFICIENCIES,HEMATOPOEITIC GROWTH FACTORS|[IN400] INVEST HEMATOLOGIC DEFICIENCIES,HEMATOPOEITIC GROWTH FACTORS
C1875317|T121|N0000029624|NDFRT|INVEST HORMONE THERAPY/REPLACEMENT ANDROGEN AND ANABOLIC|[IN900] INVEST HORMONE THERAPY/REPLACEMENT ANDROGEN AND ANABOLIC
C1875318|T121|N0000029625|NDFRT|INVEST HORMONE THERAPY/REPLACEMENT ESTROGENS AND PROGESTINS|[IN910] INVEST HORMONE THERAPY/REPLACEMENT ESTROGENS AND PROGESTINS
C1875319|T121|N0000029201|NDFRT|INVESTIGATIONAL AGENTS|[IN000] INVESTIGATIONAL AGENTS
C1875320|T121|N0000029588|NDFRT|INVESTIGATIONAL ANALGESICS|[IN500] INVESTIGATIONAL ANALGESICS
C1875321|T121|N0000029590|NDFRT|INVESTIGATIONAL ANESTHETICS|[IN510] INVESTIGATIONAL ANESTHETICS
C1875322|T121|N0000029602|NDFRT|INVESTIGATIONAL ANTI-ANGINA DRUGS|[IN600] INVESTIGATIONAL ANTI-ANGINA DRUGS
C1875323|T121|N0000029592|NDFRT|INVESTIGATIONAL ANTI-ANXIETY DRUGS|[IN520] INVESTIGATIONAL ANTI-ANXIETY DRUGS
C1875324|T121|N0000029559|NDFRT|INVESTIGATIONAL ANTI-BACTERIAL DRUGS|[IN100] INVESTIGATIONAL ANTI-BACTERIAL DRUGS
C1875325|T121|N0000029593|NDFRT|INVESTIGATIONAL ANTI-CONVULSANT DRUGS|[IN530] INVESTIGATIONAL ANTI-CONVULSANT DRUGS
C1875326|T121|N0000029595|NDFRT|INVESTIGATIONAL ANTI-DEPRESSANTS|[IN550] INVESTIGATIONAL ANTI-DEPRESSANTS
C1875327|T121|N0000029626|NDFRT|INVESTIGATIONAL ANTI-DIABETIC DRUGS|[IN920] INVESTIGATIONAL ANTI-DIABETIC DRUGS
C1875328|T121|N0000029619|NDFRT|INVESTIGATIONAL ANTI-DIARRHEAL DRUGS|[IN840] INVESTIGATIONAL ANTI-DIARRHEAL DRUGS
C1875329|T121|N0000029603|NDFRT|INVESTIGATIONAL ANTI-DYSRHYTHMIC DRUGS|[IN610] INVESTIGATIONAL ANTI-DYSRHYTHMIC DRUGS
C1875330|T121|N0000029566|NDFRT|INVESTIGATIONAL ANTI-FUNGAL DRUGS|[IN120] INVESTIGATIONAL ANTI-FUNGAL DRUGS
C1875331|T121|N0000029614|NDFRT|INVESTIGATIONAL ANTI-GLAUCOMA DRUGS|[IN720] INVESTIGATIONAL ANTI-GLAUCOMA DRUGS
C1875332|T121|N0000029605|NDFRT|INVESTIGATIONAL ANTI-HYPERTENSIVE DRUGS|[IN630] INVESTIGATIONAL ANTI-HYPERTENSIVE DRUGS
C1875333|T121|N0000029571|NDFRT|INVESTIGATIONAL ANTI-INFECTIVE DRUGS,OTHER|[IN170] INVESTIGATIONAL ANTI-INFECTIVE DRUGS,OTHER
C1875334|T121|N0000029620|NDFRT|INVESTIGATIONAL ANTI-NAUSEA AND ANTI-EMETIC DRUGS|[IN850] INVESTIGATIONAL ANTI-NAUSEA AND ANTI-EMETIC DRUGS
C1875335|T121|N0000029574|NDFRT|INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS CNS|[IN210] INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS CNS
C1875336|T121|N0000029577|NDFRT|INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS GENITOURINARY ORGANS|[IN240] INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS GENITOURINARY ORGANS
C1875337|T121|N0000029578|NDFRT|INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS INTRATHORACIC ORGANS|[IN250] INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS INTRATHORACIC ORGANS
C1875338|T121|N0000029576|NDFRT|INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS, GENE THERAPY|[IN230] INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS, GENE THERAPY
C1875339|T121|N0000029581|NDFRT|INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS,OTHER|[IN280] INVESTIGATIONAL ANTI-NEOPLASTIC DRUGS,OTHER
C1875340|T121|N0000029582|NDFRT|INVESTIGATIONAL ANTI-PARASITIC DRUGS|[IN300] INVESTIGATIONAL ANTI-PARASITIC DRUGS
C1875341|T121|N0000029585|NDFRT|INVESTIGATIONAL ANTI-THROMBOTIC DRUGS|[IN410] INVESTIGATIONAL ANTI-THROMBOTIC DRUGS
C1875342|T121|N0000029565|NDFRT|INVESTIGATIONAL ANTI-TUBERCULAR DRUGS|[IN110] INVESTIGATIONAL ANTI-TUBERCULAR DRUGS
C1875343|T121|N0000029567|NDFRT|INVESTIGATIONAL ANTI-VIRAL DRUGS HEPATITIS B|[IN130] INVESTIGATIONAL ANTI-VIRAL DRUGS HEPATITIS B
C1875344|T121|N0000029568|NDFRT|INVESTIGATIONAL ANTI-VIRAL DRUGS HEPATITIS C|[IN140] INVESTIGATIONAL ANTI-VIRAL DRUGS HEPATITIS C
C1875345|T121|N0000029569|NDFRT|INVESTIGATIONAL ANTI-VIRAL DRUGS HIV|[IN150] INVESTIGATIONAL ANTI-VIRAL DRUGS HIV
C1875346|T121|N0000029570|NDFRT|INVESTIGATIONAL ANTI-VIRAL DRUGS,OTHER|[IN160] INVESTIGATIONAL ANTI-VIRAL DRUGS,OTHER
C1875347|T121|N0000029606|NDFRT|INVESTIGATIONAL CONGESTIVE HEART FAILURE|[IN640] INVESTIGATIONAL CONGESTIVE HEART FAILURE
C1875348|T121|N0000029562|NDFRT|INVESTIGATIONAL DIAGNOSTIC AGENTS,GLUCOSE TESTING|[IN003] INVESTIGATIONAL DIAGNOSTIC AGENTS,GLUCOSE TESTING
C1875349|T121|N0000029560|NDFRT|INVESTIGATIONAL DIAGNOSTIC AGENTS,OTHER|[IN001] INVESTIGATIONAL DIAGNOSTIC AGENTS,OTHER
C1875350|T121|N0000029561|NDFRT|INVESTIGATIONAL DIAGNOSTIC AGENTS,SKIN TESTING|[IN002] INVESTIGATIONAL DIAGNOSTIC AGENTS,SKIN TESTING
C1875351|T121|N0000029608|NDFRT|INVESTIGATIONAL DRUGS FOR ALLERGY AND NASAL CONGESTION|[IN660] INVESTIGATIONAL DRUGS FOR ALLERGY AND NASAL CONGESTION
C1875352|T121|N0000029591|NDFRT|INVESTIGATIONAL DRUGS FOR ARTHRITIS AND GOUT|[IN515] INVESTIGATIONAL DRUGS FOR ARTHRITIS AND GOUT
C1875353|T121|N0000029610|NDFRT|INVESTIGATIONAL DRUGS FOR ASTHMA AND COPD|[IN670] INVESTIGATIONAL DRUGS FOR ASTHMA AND COPD
C1875354|T121|N0000029596|NDFRT|INVESTIGATIONAL DRUGS FOR CENTRAL AND PERIPHERAL NEUROPATHY|[IN560] INVESTIGATIONAL DRUGS FOR CENTRAL AND PERIPHERAL NEUROPATHY
C1875355|T121|N0000029616|NDFRT|INVESTIGATIONAL DRUGS FOR CONSTIPATION|[IN810] INVESTIGATIONAL DRUGS FOR CONSTIPATION
C1875356|T121|N0000029599|NDFRT|INVESTIGATIONAL DRUGS FOR DEMENTIA|[IN585] INVESTIGATIONAL DRUGS FOR DEMENTIA
C1875357|T121|N0000029604|NDFRT|INVESTIGATIONAL DRUGS FOR DYSLIPIDEMIAS|[IN620] INVESTIGATIONAL DRUGS FOR DYSLIPIDEMIAS
C1875358|T121|N0000029615|NDFRT|INVESTIGATIONAL DRUGS FOR DYSPEPSIA|[IN800] INVESTIGATIONAL DRUGS FOR DYSPEPSIA
C1875359|T121|N0000029618|NDFRT|INVESTIGATIONAL DRUGS FOR GASTROESOPHAGEAL REFLUX DISEASE|[IN830] INVESTIGATIONAL DRUGS FOR GASTROESOPHAGEAL REFLUX DISEASE
C1875360|T121|N0000029587|NDFRT|INVESTIGATIONAL DRUGS FOR HEMATOLOGIC DEFICIENCIES,OTHER|[IN430] INVESTIGATIONAL DRUGS FOR HEMATOLOGIC DEFICIENCIES,OTHER
C1875361|T121|N0000029630|NDFRT|INVESTIGATIONAL DRUGS FOR IMMUNOLOGIC DISEASES,OTHER|[IN960] INVESTIGATIONAL DRUGS FOR IMMUNOLOGIC DISEASES,OTHER
C1875362|T121|N0000029598|NDFRT|INVESTIGATIONAL DRUGS FOR MANIA AND BIPOLAR DISORDERS|[IN580] INVESTIGATIONAL DRUGS FOR MANIA AND BIPOLAR DISORDERS
C1875363|T121|N0000029589|NDFRT|INVESTIGATIONAL DRUGS FOR MUSCULOSKELETAL CONDITIONS,OTHER|[IN505] INVESTIGATIONAL DRUGS FOR MUSCULOSKELETAL CONDITIONS,OTHER
C1875364|T121|N0000029609|NDFRT|INVESTIGATIONAL DRUGS FOR NASAL/THROAT DISEASES,OTHER|[IN665] INVESTIGATIONAL DRUGS FOR NASAL/THROAT DISEASES,OTHER
C1875365|T121|N0000029583|NDFRT|INVESTIGATIONAL DRUGS FOR ORGAN TRANSPLANTATION|[IN350] INVESTIGATIONAL DRUGS FOR ORGAN TRANSPLANTATION
C1875366|T121|N0000029613|NDFRT|INVESTIGATIONAL DRUGS FOR OTHER DERMATOLOGICAL DISEASES|[IN710] INVESTIGATIONAL DRUGS FOR OTHER DERMATOLOGICAL DISEASES
C1875367|T121|N0000029621|NDFRT|INVESTIGATIONAL DRUGS FOR OTHER GASTROINTESTINAL DISEASES|[IN860] INVESTIGATIONAL DRUGS FOR OTHER GASTROINTESTINAL DISEASES
C1875368|T121|N0000029633|NDFRT|INVESTIGATIONAL DRUGS FOR OTHER INDICATIONS|[IN999] INVESTIGATIONAL DRUGS FOR OTHER INDICATIONS
C1875369|T121|N0000029622|NDFRT|INVESTIGATIONAL DRUGS FOR PANCREATIC ENZYME DEFICIENCY|[IN870] INVESTIGATIONAL DRUGS FOR PANCREATIC ENZYME DEFICIENCY
C1875370|T121|N0000029594|NDFRT|INVESTIGATIONAL DRUGS FOR PARKINSON'S DISEASE|[IN540] INVESTIGATIONAL DRUGS FOR PARKINSON'S DISEASE
C1875371|T121|N0000029617|NDFRT|INVESTIGATIONAL DRUGS FOR PEPTIC ULCER DISEASE|[IN820] INVESTIGATIONAL DRUGS FOR PEPTIC ULCER DISEASE
C1875372|T121|N0000029600|NDFRT|INVESTIGATIONAL DRUGS FOR PSYCHIATRIC DISEASE,OTHER|[IN590] INVESTIGATIONAL DRUGS FOR PSYCHIATRIC DISEASE,OTHER
C1875373|T121|N0000029611|NDFRT|INVESTIGATIONAL DRUGS FOR RESPIRATORY TRACT DISEASE,OTHER|[IN675] INVESTIGATIONAL DRUGS FOR RESPIRATORY TRACT DISEASE,OTHER
C1875374|T121|N0000029601|NDFRT|INVESTIGATIONAL DRUGS FOR SUBSTANCE ADDICTION TREATMENT|[IN595] INVESTIGATIONAL DRUGS FOR SUBSTANCE ADDICTION TREATMENT
C1875375|T121|N0000029632|NDFRT|INVESTIGATIONAL DRUGS FOR VITAMIN OR MINERAL DEFICIENCY|[IN980] INVESTIGATIONAL DRUGS FOR VITAMIN OR MINERAL DEFICIENCY
C1875376|T121|N0000029629|NDFRT|INVESTIGATIONAL GENE THERAPY|[IN950] INVESTIGATIONAL GENE THERAPY
C1875377|T121|N0000029627|NDFRT|INVESTIGATIONAL HORMONE THERAPY/REPLACEMENT, THYROID|[IN930] INVESTIGATIONAL HORMONE THERAPY/REPLACEMENT, THYROID
C1875378|T121|N0000029628|NDFRT|INVESTIGATIONAL HORMONE THERAPY/REPLACEMENT,OTHER|[IN940] INVESTIGATIONAL HORMONE THERAPY/REPLACEMENT,OTHER
C1875379|T121|N0000029607|NDFRT|INVESTIGATIONAL OTHER CARDIOVASCULAR DISEASES|[IN650] INVESTIGATIONAL OTHER CARDIOVASCULAR DISEASES
C1875380|T121|N0000029563|NDFRT|INVESTIGATIONAL PHARMACEUTICAL AIDS/REAGENTS|[IN004] INVESTIGATIONAL PHARMACEUTICAL AIDS/REAGENTS
C1875381|T121|N0000029564|NDFRT|INVESTIGATIONAL PROSTHETICS/SUPPLIES/DEVICES|[IN005] INVESTIGATIONAL PROSTHETICS/SUPPLIES/DEVICES
C1875382|T121|N0000029631|NDFRT|INVESTIGATIONAL THERAPEUTIC NUTRIENTS/MINERAL/ELECTROLYTES|[IN970] INVESTIGATIONAL THERAPEUTIC NUTRIENTS/MINERAL/ELECTROLYTES
C1875383|T121|N0000029586|NDFRT|INVESTIGATIONAL THROMBOLYTIC DRUGS|[IN420] INVESTIGATIONAL THROMBOLYTIC DRUGS
C1875384|T121|N0000029572|NDFRT|INVESTIGATIONAL VACCINES|[IN180] INVESTIGATIONAL VACCINES
C1875388|T121|N0000029306|NDFRT|IONIC CONTRAST MEDIA|[DX102] IONIC CONTRAST MEDIA
C1875396|T121|N0000029202|NDFRT|IRRIGATION/DIALYSIS SOLUTIONS|[IR000] IRRIGATION/DIALYSIS SOLUTIONS
C1875397|T121|N0000029431|NDFRT|IRRIGATION/DIALYSIS SOLUTIONS,OTHER|[IR900] IRRIGATION/DIALYSIS SOLUTIONS,OTHER
C1875408|T121|N0000029254|NDFRT|IV SOLUTIONS|[TN100] IV SOLUTIONS
C1875409|T121|N0000029256|NDFRT|IV SOLUTIONS WITH ELECTROLYTES|[TN102] IV SOLUTIONS WITH ELECTROLYTES
C1875410|T121|N0000029255|NDFRT|IV SOLUTIONS WITHOUT ELECTROLYTES|[TN101] IV SOLUTIONS WITHOUT ELECTROLYTES
C1875417|T121|N0000029159|NDFRT|KERATOLYTICS/CAUSTICS,TOPICAL|[DE500] KERATOLYTICS/CAUSTICS,TOPICAL
C1875434|T121|N0000029251|NDFRT|LAXATIVES,RECTAL|[RS300] LAXATIVES,RECTAL
C1875444|T121|N0000029258|NDFRT|LIPID SUPPLEMENTS|[TN300] LIPID SUPPLEMENTS
C1875449|T121|N0000029142|NDFRT|LOCAL ANESTHETICS,INJECTION|[CN204] LOCAL ANESTHETICS,INJECTION
C1875450|T121|N0000029161|NDFRT|LOCAL ANESTHETICS,TOPICAL|[DE700] LOCAL ANESTHETICS,TOPICAL
C1875454|T121|N0000029391|NDFRT|LUBRICANT LAXATIVES|[GA203] LUBRICANT LAXATIVES
C1875456|T121|N0000029384|NDFRT|MAGALDRATE CONTAINING ANTACIDS|[GA107] MAGALDRATE CONTAINING ANTACIDS
C1875461|T121|N0000029385|NDFRT|MAGNESIUM CONTAINING ANTACIDS|[GA108] MAGNESIUM CONTAINING ANTACIDS
C1875464|T121|N0000029386|NDFRT|MAGNESIUM/SODIUM BICARBONATE CONTAINING ANTACIDS|[GA109] MAGNESIUM/SODIUM BICARBONATE CONTAINING ANTACIDS
C1875486|T121|N0000029085|NDFRT|METHENAMINE SALTS ANTIMICROBIALS|[AM550] METHENAMINE SALTS ANTIMICROBIALS
C1875506|T121|N0000029324|NDFRT|MIOTICS,TOPICAL OPHTHALMIC|[OP102] MIOTICS,TOPICAL OPHTHALMIC
C1875508|T121|N0000029149|NDFRT|MONAMINE OXIDASE INHIBITOR ANTIDEPRESSANTS|[CN602] MONAMINE OXIDASE INHIBITOR ANTIDEPRESSANTS
C1875516|T121|N0000029211|NDFRT|MUSCULOSKELETAL AGENTS,OTHER|[MS900] MUSCULOSKELETAL AGENTS,OTHER
C1875517|T121|N0000029206|NDFRT|MUSCULOSKELETAL MEDICATIONS|[MS000] MUSCULOSKELETAL MEDICATIONS
C1875518|T121|N0000029222|NDFRT|MYDRIATICS/CYCLOPLEGICS,TOPICAL OPHTHALMIC|[OP600] MYDRIATICS/CYCLOPLEGICS,TOPICAL OPHTHALMIC
C1875521|T121|N0000029212|NDFRT|NASAL AND THROAT AGENTS,TOPICAL|[NT000] NASAL AND THROAT AGENTS,TOPICAL
C1875522|T121|N0000029336|NDFRT|NASAL AND THROAT,TOPICAL,OTHER|[NT900] NASAL AND THROAT,TOPICAL,OTHER
C1875539|T121|N0000029086|NDFRT|NITROFURANS ANTIMICROBIALS|[AM600] NITROFURANS ANTIMICROBIALS
C1875542|T121|N0000029343|NDFRT|NON-ANESTHETIC GASES|[RE600] NON-ANESTHETIC GASES
C1875543|T121|N0000029308|NDFRT|NON-IMAGING AGENTS RADIOPHARMACEUTICALS|[DX202] NON-IMAGING AGENTS RADIOPHARMACEUTICALS
C1875544|T121|N0000029305|NDFRT|NON-IONIC CONTRAST MEDIA|[DX101] NON-IONIC CONTRAST MEDIA
C1875545|T121|N0000029409|NDFRT|NON-OPIOID-CONTAINING ANTITUSSIVES/EXPECTORANTS|[RE302] NON-OPIOID-CONTAINING ANTITUSSIVES/EXPECTORANTS
C1875546|T121|N0000029137|NDFRT|NON-STEROIDAL ANTI-INFLAMMATORY ANALGESICS|[CN104] NON-STEROIDAL ANTI-INFLAMMATORY ANALGESICS
C1875547|T121|N0000029318|NDFRT|NONSALICYLATE NSAIS,ANTIRHEUMATIC|[MS102] NONSALICYLATE NSAIS,ANTIRHEUMATIC
C1875577|T121|N0000029224|NDFRT|OPHTHALMICS,OTHER|[OP900] OPHTHALMICS,OTHER
C1875578|T121|N0000029134|NDFRT|OPIOID ANTAGONIST ANALGESICS|[CN102] OPIOID ANTAGONIST ANALGESICS
C1875579|T121|N0000029408|NDFRT|OPIOID-CONTAINING ANTITUSSIVES/EXPECTORANTS|[RE301] OPIOID-CONTAINING ANTITUSSIVES/EXPECTORANTS
C1875585|T121|N0000029185|NDFRT|ORAL HYPOGLYCEMIC AGENTS,ORAL|[HS502] ORAL HYPOGLYCEMIC AGENTS,ORAL
C1875589|T121|N0000029354|NDFRT|OSMOTIC AGENTS,SYSTEMIC OPHTHALMIC|[OP160] OSMOTIC AGENTS,SYSTEMIC OPHTHALMIC
C1875591|T121|N0000029235|NDFRT|OTIC AGENTS,OTHER|[OT900] OTIC AGENTS,OTHER
C1875624|T121|N0000029106|NDFRT|PARASYMPATHOMIMETICS (CHOLINERGICS)|[AU300] PARASYMPATHOMIMETICS (CHOLINERGICS)
C1875631|T121|N0000029292|NDFRT|PENICILLIN-G RELATED PENICILLINS|[AM110] PENICILLIN-G RELATED PENICILLINS
C1875633|T121|N0000029076|NDFRT|PENICILLINS AND BETA-LACTAM ANTIMICROBIALS|[AM114] PENICILLINS AND BETA-LACTAM ANTIMICROBIALS
C1875643|T121|N0000029236|NDFRT|PHARMACEUTICAL AIDS/REAGENTS|[PH000] PHARMACEUTICAL AIDS/REAGENTS
C1875654|T121|N0000029151|NDFRT|PHENOTHIAZINE/RELATED ANTIPSYCHOTICS|[CN701] PHENOTHIAZINE/RELATED ANTIPSYCHOTICS
C1875688|T121|N0000029129|NDFRT|POTASSIUM SPARING/COMBINATIONS DIURETICS|[CV704] POTASSIUM SPARING/COMBINATIONS DIURETICS
C1875707|T121|N0000029310|NDFRT|PROTECTANTS,ULCER|[GA302] PROTECTANTS,ULCER
C1875717|T121|N0000029165|NDFRT|RADIOLOGICAL/CONTRAST MEDIA|[DX100] RADIOLOGICAL/CONTRAST MEDIA
C1875720|T121|N0000029248|NDFRT|RECTAL,LOCAL|[RS000] RECTAL,LOCAL
C1875721|T121|N0000029252|NDFRT|RECTAL,LOCAL OTHER|[RS900] RECTAL,LOCAL OTHER
C1875728|T121|N0000029247|NDFRT|RESPIRATORY AGENTS,OTHER|[RE900] RESPIRATORY AGENTS,OTHER
C1875729|T121|N0000029237|NDFRT|RESPIRATORY TRACT MEDICATIONS|[RE000] RESPIRATORY TRACT MEDICATIONS
C1875734|T121|N0000029317|NDFRT|SALICYLATES,ANTIRHEUMATIC|[MS101] SALICYLATES,ANTIRHEUMATIC
C1875739|T121|N0000029424|NDFRT|SEDATIVES/HYPNOTICS,OTHER|[CN309] SEDATIVES/HYPNOTICS,OTHER
C1875740|T121|N0000029143|NDFRT|SEDATIVES/HYPONTICS|[CN300] SEDATIVES/HYPONTICS
C1875761|T121|N0000029158|NDFRT|SOAPS/SHAMPOOS/SOAP-FREE CLEANSERS|[DE400] SOAPS/SHAMPOOS/SOAP-FREE CLEANSERS
C1875763|T121|N0000029387|NDFRT|SODIUM BICARBONATE CONTAINING ANTACIDS|[GA110] SODIUM BICARBONATE CONTAINING ANTACIDS
C1875793|T121|N0000029087|NDFRT|SULFONAMIDE/RELATED ANTIMICROBIALS|[AM650] SULFONAMIDE/RELATED ANTIMICROBIALS
C1875798|T121|N0000029157|NDFRT|SUN PROTECTANTS/SCREENS,TOPICAL|[DE300] SUN PROTECTANTS/SCREENS,TOPICAL
C1875809|T121|N0000029104|NDFRT|SYMPATHOMIMETICS (ADRENERGICS)|[AU100] SYMPATHOMIMETICS (ADRENERGICS)
C1875826|T121|N0000029259|NDFRT|THERAPEUTIC NUTRIENTS/MINERALS/ELECTROLYES,OTHER|[TN900] THERAPEUTIC NUTRIENTS/MINERALS/ELECTROLYES,OTHER
C1875830|T121|N0000029190|NDFRT|THYROID MODIFIERS|[HS850] THYROID MODIFIERS
C1875831|T121|N0000029191|NDFRT|THYROID SUPPLEMENTS|[HS851] THYROID SUPPLEMENTS
C1875852|T121|N0000029636|NDFRT|VACCINES/TOXOIDS, OTHER|[IM109] VACCINES/TOXOIDS, OTHER
C1875860|T121|N0000029456|NDFRT|VITAMIN B,OTHER|[VT109] VITAMIN B,OTHER
C1875861|T121|N0000029361|NDFRT|VITAMIN COMBINATIONS,OTHER|[VT809] VITAMIN COMBINATIONS,OTHER
C1875862|T121|N0000029462|NDFRT|VITAMIN D,OTHER|[VT509] VITAMIN D,OTHER
C1875863|T121|N0000029465|NDFRT|VITAMIN K,OTHER|[VT709] VITAMIN K,OTHER
C1875864|T121|N0000029273|NDFRT|VITAMINS,COMBINATIONS|[VT800] VITAMINS,COMBINATIONS
C1875865|T121|N0000029348|NDFRT|VOLUME EXPANDERS|[BL800] VOLUME EXPANDERS
C1950687|T121|N0000175986|NDFRT|DIRECT RENIN INHIBITOR|[CV806] DIRECT RENIN INHIBITOR
C2240799|T121|N0000175988|NDFRT|HYPOGLYCEMIC AGENTS,OTHER|[HS509] HYPOGLYCEMIC AGENTS,OTHER
C2365945|T121|N0000177916|NDFRT|VESICULAR MONOAMINE TRANSPORT TYPE 2 BLOCKER|[MS205] VESICULAR MONOAMINE TRANSPORT TYPE 2 BLOCKER
C2746010|T121|N0000029203|NDFRT|IRRIGATION SOLUTIONS|[IR100] IRRIGATION SOLUTIONS
C3537168|T121|N0000029120|NDFRT|ANTIANGINALS|[CV250] ANTIANGINALS
C3537192|T121|N0000175987|NDFRT|TUMOR NECROSIS FACTOR BLOCKER|[GA400] TUMOR NECROSIS FACTOR BLOCKER
C3714498|T121|N0000029443|NDFRT|PHOSPHORUS|[TN475] PHOSPHORUS
C3714501|T121|N0000029184|NDFRT|INSULIN|[HS501] INSULIN
C3714502|T121|N0000029454|NDFRT|RIBOFLAVIN|[VT106] RIBOFLAVIN
C3714503|T121|N0000029270|NDFRT|VITAMIN D|[VT500] VITAMIN D
C3714504|T121|N0000029460|NDFRT|DIHYDROTACHYSTEROL|[VT503] DIHYDROTACHYSTEROL
C3714601|T121|N0000029445|NDFRT|CITRATES|[TN478] CITRATES
C3714609|T121|N0000029458|NDFRT|CALCIFEDIOL|[VT501] CALCIFEDIOL
C3714610|T121|N0000029459|NDFRT|CALCITRIOL|[VT502] CALCITRIOL
C3714611|T121|N0000029437|NDFRT|CALCIUM|[TN420] CALCIUM
C3714612|T121|N0000029080|NDFRT|CHLORAMPHENICOL|[AM150] CHLORAMPHENICOL
C3714615|T121|N0000029181|NDFRT|ESTROGENS|[HS300] ESTROGENS
C3714616|T121|N0000029442|NDFRT|FLUORIDE|[TN470] FLUORIDE
C3714620|T121|N0000029296|NDFRT|LINCOMYCINS|[AM350] LINCOMYCINS
C3714621|T121|N0000029441|NDFRT|MAGNESIUM|[TN460] MAGNESIUM
C3714626|T121|N0000029451|NDFRT|NICOTINIC ACID|[VT103] NICOTINIC ACID
C3714629|T121|N0000029455|NDFRT|PANTOTHENIC ACID|[VT107] PANTOTHENIC ACID
C3714631|T121|N0000029187|NDFRT|PARATHYROID|[HS600] PARATHYROID
C3714633|T121|N0000029320|NDFRT|PENICILLAMINE|[MS140] PENICILLAMINE
C3714635|T121|N0000029315|NDFRT|POSTERIOR PITUITARY|[HS702] POSTERIOR PITUITARY
C3714637|T121|N0000029438|NDFRT|POTASSIUM|[TN430] POTASSIUM
C3714638|T121|N0000029452|NDFRT|PYRIDOXINE|[VT104] PYRIDOXINE
C3714642|T121|N0000029439|NDFRT|SODIUM|[TN440] SODIUM
C3714647|T121|N0000029457|NDFRT|VITAMIN B|[VT100] VITAMIN B
C3714648|T121|N0000029272|NDFRT|VITAMIN K|[VT700] VITAMIN K
C3714649|T121|N0000029267|NDFRT|VITAMINS|[VT000] VITAMINS
C3714650|T121|N0000029440|NDFRT|ZINC|[TN450] ZINC
C3714656|T121|N0000029268|NDFRT|VITAMIN A|[VT050] VITAMIN A
C3714687|T121|N0000029269|NDFRT|VITAMIN C|[VT400] VITAMIN C
C3714696|T121|N0000029461|NDFRT|ERGOCALCIFEROL|[VT504] ERGOCALCIFEROL
C3714701|T121|N0000029436|NDFRT|IRON|[TN410] IRON
C3714706|T121|N0000029463|NDFRT|MENADIOL|[VT701] MENADIOL
C3714737|T121|N0000029464|NDFRT|PHYTONADIONE|[VT702] PHYTONADIONE
C3714801|T121|N0000029449|NDFRT|CYANOCOBALAMIN|[VT101] CYANOCOBALAMIN
C3714802|T121|N0000029453|NDFRT|THIAMINE|[VT105] THIAMINE
C3714803|T121|N0000029271|NDFRT|VITAMIN E|[VT600] VITAMIN E
C3714835|T121|N0000029360|NDFRT|MULTIVITAMINS|[VT801] MULTIVITAMINS
