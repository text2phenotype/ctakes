// Index|Test name|Text|IsCorrect
0|Correct facility|CENTER FOR HEALTH EDUCATION AND DENTISTRY|True
1|Incorrect facility|CENTRE FOR HEALTH EDUCATION AND DENTISTRY|False