C3828565|T034|328661|MEDCIN|PHQ-9: TOTAL SCORE|PHQ-9: TOTAL SCORE (PROCEDURE)
C1718207|T034||MEDCIN|PHQ-9 INTERPRETATION
C1718207|T034||MEDCIN|PHQ-9 SCORE
C1718207|T034||MEDCIN|PHQ9 SCORE
C4283755|T034||MEDCIN|PATIENT HEALTH QUESTIONNAIRE NINE ITEM SCORE
C1718917|T034|328659|MEDCIN|PATIENT HEALTH QUESTIONNAIRE PHQ-9 ADMINISTRATION|PHQ-9 (PROCEDURE)
C4083201|T034||MEDCIN|PATIENT HEALTH QUESTIONNAIRE 9 ITEM
C3641315|T034||MEDCIN|PHQ-9 QUESTIONNAIRE QUESTION
C1715519|T034||MEDCIN|PATIENT HEALTH QUESTIONNAIRE 9 ITEM TOTAL SCORE:SCORE:PT:^PATIENT:QN:REPORTED.PHQ
C3828565|T034|328661|MEDCIN|PHQ01-TOTAL SCORE|PHQ-9: TOTAL SCORE (PROCEDURE)
C3828565|T034|328661|MEDCIN|PHQ-9 - TOTAL SCORE|PHQ-9: TOTAL SCORE (PROCEDURE)
C3828565|T034|328661|MEDCIN|PHQ0111|PHQ-9: TOTAL SCORE (PROCEDURE)
C3828565|T034|328661|MEDCIN|QUESTIONNAIRES PHQ-9 TOTAL SCORE|PHQ-9: TOTAL SCORE (PROCEDURE)
C3828565|T034|328661|MEDCIN|PHQ-9: TOTAL SCORE|PHQ-9: TOTAL SCORE (PROCEDURE)
C3828565|T034|328661|MEDCIN|PHQ-9: TOTAL SCORE |PHQ-9: TOTAL SCORE (PROCEDURE)
C1976603|T034|328660|MEDCIN|PHQ-9 QUICK DEPRESSION ASSESSMENT PANEL|PHQ-9: QUICK DEPRESSION ASSESSMENT PANEL (PROCEDURE)
C1976603|T034|328660|MEDCIN|QUESTIONNAIRES PHQ-9 QUICK DEPRESSION ASSESSMENT PANEL|PHQ-9: QUICK DEPRESSION ASSESSMENT PANEL (PROCEDURE)
C1976603|T034|328660|MEDCIN|PHQ-9: QUICK DEPRESSION ASSESSMENT PANEL |PHQ-9: QUICK DEPRESSION ASSESSMENT PANEL (PROCEDURE)
C1976603|T034|328660|MEDCIN|PHQ-9: QUICK DEPRESSION ASSESSMENT PANEL|PHQ-9: QUICK DEPRESSION ASSESSMENT PANEL (PROCEDURE)
C3641512|T034||MEDCIN|PHQ-9 - FEELING DOWN, DEPRESSED, OR HOPELESS
C3641512|T034||MEDCIN|PHQ01-FEELING DOWN DEPRESSED OR HOPELESS
C3641512|T034||MEDCIN|PHQ0102
C3641518|T034||MEDCIN|PHQ-9 - MOVING OR SPEAKING SLOWLY OR THE OPPOSITE BEING FIDGETY OR RESTLESS
C3641518|T034||MEDCIN|PHQ01-MOVING SLOWLY OR FIDGETY/RESTLESS
C3641518|T034||MEDCIN|PHQ0108
C3641514|T034||MEDCIN|PHQ-9 - FEELING TIRED OR HAVING LITTLE ENERGY
C3641514|T034||MEDCIN|PHQ0104
C3641514|T034||MEDCIN|PHQ01-FEELING TIRED OR LITTLE ENERGY
C3641515|T034||MEDCIN|PHQ-9 - POOR APPETITE OR OVEREATING
C3641515|T034||MEDCIN|PHQ0105
C3641515|T034||MEDCIN|PHQ01-POOR APPETITE OR OVEREATING
C3641516|T034||MEDCIN|PHQ-9 - FEELING BAD ABOUT YOURSELF
C3641516|T034||MEDCIN|PHQ01-FEELING BAD ABOUT YOURSELF
C3641516|T034||MEDCIN|PHQ0106
C3641511|T034||MEDCIN|PHQ-9 - LITTLE INTEREST OR PLEASURE IN DOING THINGS
C3641511|T034||MEDCIN|PHQ0101
C3641511|T034||MEDCIN|PHQ01-LITTLE INTEREST/PLEASURE IN THINGS
C3641520|T034||MEDCIN|PHQ01-DIFFICULT TO WORK/TAKE CARE THINGS
C3641520|T034||MEDCIN|PHQ-9 - HOW DIFFICULT HAVE PROBLEMS MADE IT FOR YOU TO WORK, TAKE CARE OF THINGS, OR GET ALONG WITH OTHER PEOPLE
C3641520|T034||MEDCIN|PHQ0110
C3641519|T034||MEDCIN|PHQ-9 - THOUGHTS THAT YOU WOULD BE BETTER OFF DEAD
C3641519|T034||MEDCIN|PHQ01-THOUGHTS YOU BE BETTER OFF DEAD
C3641519|T034||MEDCIN|PHQ0109
C3641513|T034||MEDCIN|PHQ-9 - TROUBLE FALLING OR STAYING ASLEEP, OR SLEEPING TOO MUCH
C3641513|T034||MEDCIN|PHQ01-TROUBLE FALLING OR STAYING ASLEEP
C3641513|T034||MEDCIN|PHQ0103
C3641517|T034||MEDCIN|PHQ-9 - TROUBLE CONCENTRATING ON THINGS
C3641517|T034||MEDCIN|PHQ01-TROUBLE CONCENTRATING ON THINGS
C3641517|T034||MEDCIN|PHQ0107
C1715519|T034||MEDCIN|PATIENT HEALTH QUESTIONNAIRE 9 ITEM (PHQ-9) TOTAL SCORE [REPORTED]
C1715519|T034||MEDCIN|PATIENT HEALTH QUESTIONNAIRE 9 ITEM TOTAL SCORE:SCORE:POINT IN TIME:^PATIENT:QUANTITATIVE:REPORTED.PHQ
C1715519|T034||MEDCIN|PATIENT HEALTH QUESTIONNAIRE 9 ITEM TOTAL SCORE:SCORE:PT:^PATIENT:QN:REPORTED.PHQ
