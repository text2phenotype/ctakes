C1515945|T098||CDC|AMERICAN INDIAN OR ALASKA NATIVE
C3261247|T098||CDC|AMERICAN INDIAN AND ALASKA NATIVE ALONE
C0078988|T098||CDC|ASIAN
C0003988|T098||CDC|ASIAN AMERICAN
C0438971|T098||CDC|OTHER ASIAN ETHNIC GROUP
C1524069|T098||CDC|ASIAN INDIAN
C3261249|T098||CDC|ASIAN ALONE
C0085756|T098||CDC|AFRICAN AMERICAN
C0005680|T098||CDC|BLACK RACE
C0027567|T098||CDC|AFRICAN RACE
C0085756|T098||CDC|AFRICAN AMERICAN
C0085756|T098||CDC|AFRICAN
C0085756|T098||CDC|BOTSWANAN
C0085756|T098||CDC|ETHIOPIAN
C0085756|T098||CDC|LIBERIAN
C0085756|T098||CDC|NAMIBIAN
C0085756|T098||CDC|NIGERIAN
C0085756|T098||CDC|ZAIREAN
C0085756|T098||CDC|BAHAMIAN
C0085756|T098||CDC|BARBADIAN
C0085756|T098||CDC|DOMINICA ISLANDER
C0085756|T098||CDC|DOMINICAN
C0085756|T098||CDC|HAITIAN
C0085756|T098||CDC|JAMAICAN
C0085756|T098||CDC|TOBAGOAN
C0085756|T098||CDC|TRINIDADIAN
C0085756|T098||CDC|WEST INDIAN
C1513907|T098||CDC|NATIVE HAWAIIAN OR OTHER PACIFIC ISLANDER
C1513907|T098||CDC|MELANESIAN
C1513907|T098||CDC|FIJIAN
C1513907|T098||CDC|NEW HEBRIDES
C1513907|T098||CDC|PAPUA NEW GUINEAN
C1513907|T098||CDC|SOLOMON ISLANDER
C1513907|T098||CDC|MICRONESIAN
C1513907|T098||CDC|CAROLINIAN
C1513907|T098||CDC|CHAMORRO
C1513907|T098||CDC|CHUUKESE
C1513907|T098||CDC|GUAMANIAN OR CHAMORRO
C1513907|T098||CDC|GUAMANIAN
C1513907|T098||CDC|KIRIBATI
C1513907|T098||CDC|KOSRAEAN
C1513907|T098||CDC|MARIANA ISLANDER
C1513907|T098||CDC|MARSHALLESE
C1513907|T098||CDC|PALAUAN
C1513907|T098||CDC|POHNPEIAN
C1513907|T098||CDC|SAIPANESE
C1513907|T098||CDC|YAPESE
C1513907|T098||CDC|OTHER PACIFIC ISLANDER
C1513907|T098||CDC|POLYNESIAN
C1513907|T098||CDC|NATIVE HAWAIIAN
C1513907|T098||CDC|SAMOAN
C1513907|T098||CDC|TAHITIAN
C1513907|T098||CDC|TOKELAUAN
C1513907|T098||CDC|TONGAN
C0043157|T098||CDC|CAUCASIANS
C0043157|T098||CDC|EUROPEAN
C0043157|T098||CDC|ARMENIAN
C0043157|T098||CDC|ENGLISH
C0043157|T098||CDC|FRENCH
C0043157|T098||CDC|GERMAN
C0043157|T098||CDC|IRISH
C0043157|T098||CDC|ITALIAN
C0043157|T098||CDC|POLISH
C0043157|T098||CDC|SCOTTISH
C0221786|T098||CDC|WHITE AMERICAN
C1535514|T098||CDC|EUROPEAN RACE
C0086409|T098||CDC|HISPANICS
C0086409|T098||CDC|CENTRAL AMERICAN
C0086409|T098||CDC|CANAL ZONE
C0086409|T098||CDC|CENTRAL AMERICAN INDIAN
C0086409|T098||CDC|COSTA RICAN
C0086409|T098||CDC|GUATEMALAN
C0086409|T098||CDC|HONDURAN
C0086409|T098||CDC|NICARAGUAN
C0086409|T098||CDC|PANAMANIAN
C0086409|T098||CDC|SALVADORAN
C0086409|T098||CDC|CUBAN
C0086409|T098||CDC|DOMINICAN
C0086409|T098||CDC|LATIN AMERICAN
C0086409|T098||CDC|MEXICAN
C0086409|T098||CDC|CHICANO
C0086409|T098||CDC|LA RAZA
C0086409|T098||CDC|MEXICAN AMERICAN INDIAN
C0086409|T098||CDC|MEXICAN AMERICAN
C0086409|T098||CDC|MEXICANO
C0086409|T098||CDC|PUERTO RICAN
C0086409|T098||CDC|SOUTH AMERICAN
C0086409|T098||CDC|ARGENTINEAN
C0086409|T098||CDC|BOLIVIAN
C0086409|T098||CDC|CHILEAN
C0086409|T098||CDC|COLOMBIAN
C0086409|T098||CDC|CRIOLLO
C0086409|T098||CDC|ECUADORIAN
C0086409|T098||CDC|PARAGUAYAN
C0086409|T098||CDC|PERUVIAN
C0086409|T098||CDC|SOUTH AMERICAN INDIAN
C0086409|T098||CDC|URUGUAYAN
C0086409|T098||CDC|VENEZUELAN
C0086409|T098||CDC|SPANIARD
C0086409|T098||CDC|ANDALUSIAN
C0086409|T098||CDC|ASTURIAN
C0086409|T098||CDC|BELEARIC ISLANDER
C0086409|T098||CDC|CANARIAN
C0086409|T098||CDC|CASTILLIAN
C0086409|T098||CDC|CATALONIAN
C0086409|T098||CDC|GALLEGO
C0086409|T098||CDC|SPANISH BASQUE
C0086409|T098||CDC|VALENCIAN
C3846650|T098||CDC|SPANISH,NOS; HISPANIC,NOS
C0019576|T098||CDC|HISPANIC AMERICANS
C1533017|T098||CDC|HISPANIC BLACK FINDING
C1533018|T098||CDC|HISPANIC BLACK RACIAL GROUP
C1533020|T098||CDC|HISPANIC WHITE FINDING
C1533021|T098||CDC|HISPANIC WHITE RACIAL GROUP
C1881927|T098||CDC|MULTIPLE HISPANIC
C2741637|T098||CDC|HISPANIC OR LATINO:FINDING:POINT IN TIME:^PATIENT:ORDINA
C3844642|T098||CDC|OTHER HISPANIC
C4036190|T098||CDC|YES, ANOTHER HISPANIC, LATINO-A, OR SPANISH ORIGIN
C3161701|T098||CDC|CULTURAL BACKGROUND ALASKAN NATIVE (___ %) 
C3161701|T098||CDC|CULTURAL BACKGROUND ALASKAN NATIVE (___ %)
C0002460|T098||CDC|AMERICAN INDIAN
C0002460|T098||CDC|AMERICAN INDIANS
C0002460|T098||CDC|INDIAN, AMERICAN
C0002460|T098||CDC|INDIANS, AMERICAN
C0002460|T098||CDC|RACEAMERICANINDIAN
C0002460|T098||CDC|AMERICAN INDIAN RACE 
C0002460|T098||CDC|AMERICAN INDIAN RACE
C0002460|T098||CDC|AMERINDIAN RACE
C0002460|T098||CDC|AMERINDIAN
C0002460|T098||CDC|INDIANS (AMERICAN)
C0002460|T098||CDC|AMERICAN INDIAN RACE (RACIAL GROUP)
C0682125|T098||CDC|ALASKA INDIAN
C0682125|T098||CDC|RACEALASKANNATIVE
C0682125|T098||CDC|RACEALASKANINDIAN
C0682125|T098||CDC|ALASKA NATIVE
C0682125|T098||CDC|ALASKA NATIVES
C0682125|T098||CDC|NATIVE ALASKANS
C0682125|T098||CDC|ALASKA INDIANS
C0152035|T098||CDC|CHINESE
C0152035|T098||CDC|CHINESE PEOPLE
C0152035|T098||CDC|CHINESE 
C0152035|T098||CDC|-- CHINESE
C1556094|T098||CDC|JAPANESE
C1556094|T098||CDC|RACE: JAPANESE 
C1556094|T098||CDC|RACE: JAPANESE
C1556094|T098||CDC|-- JAPANESE
C1556094|T098||CDC|JAPANESE 
C1556094|T098||CDC|JAPANESE RACE
C0238697|T098||CDC|SOUTHEAST ASIAN
C0238697|T098||CDC|SOUTH EAST ASIAN
C0238697|T098||CDC|SOUTH EAST ASIAN 
C0596476|T098||CDC|EAST INDIAN
C1556093|T098||CDC|FILIPINO
C1556093|T098||CDC|-- FILIPINO
C1556093|T098||CDC|FILIPINOS
C1556093|T098||CDC|FILIPINOS 
C1556093|T098||CDC|FILIPINO RACE
C0078988|T098||CDC|ASIAN
C0078988|T098||CDC|ASIANS
C0078988|T098||CDC|ORIENTAL
C0078988|T098||CDC|RACEASIAN
C0078988|T098||CDC|ASIAN RACE
C0078988|T098||CDC|RACE: ORIENTAL 
C0078988|T098||CDC|ASIAN RACE 
C0078988|T098||CDC|RACE: ORIENTAL
C0078988|T098||CDC|ORIENTAL 
C0078988|T098||CDC|ASIAN RACE (RACIAL GROUP)
C0438971|T098||CDC|OTHER ASIAN ETHNIC GROUP
C0438971|T098||CDC|OTHER ASIAN 
C0438971|T098||CDC|OTHER ASIAN ETHNIC GROUP 
C0438971|T098||CDC|OTHER ASIAN
C0438971|T098||CDC|-- OTHER ASIAN
C0870279|T098||CDC|CHINESE CULTURAL GROUPS
C0870754|T098||CDC|JAPANESE CULTURAL GROUPS
C0870776|T098||CDC|KOREAN CULTURAL GROUPS
C0871579|T098||CDC|VIETNAMESE CULTURAL GROUPS
C1510645|T098||CDC|SOUTH ASIAN CULTURAL GROUPS
C1510577|T098||CDC|SOUTHEAST ASIAN CULTURAL GROUPS
C1553332|T098||CDC|MALAGASY
C1553332|T098||CDC|MADAGASCAR
C1553332|T098||CDC|MADAGASCAR RACE
C1553322|T098||CDC|BURMESE
C1553322|T098||CDC|BURMESES
C0337900|T098||CDC|INDONESIAN
C0337900|T098||CDC|INDONESIANS
C0337900|T098||CDC|INDONESIANS 
C1556095|T098||CDC|KOREAN
C1556095|T098||CDC|RACE: KOREAN
C1556095|T098||CDC|RACE: KOREAN 
C1556095|T098||CDC|-- KOREAN
C1556095|T098||CDC|KOREANS
C1556095|T098||CDC|KOREANS 
C1556095|T098||CDC|KOREAN RACE
C0337910|T098||CDC|THAI
C0337910|T098||CDC|THAUS
C0337910|T098||CDC|THAIS (POPULATION GROUP)
C0337910|T098||CDC|THAIS
C0337910|T098||CDC|THAIS 
C1561452|T098||CDC|VIETNAMESE
C1561452|T098||CDC|VIETNAMESES
C1561452|T098||CDC|VIETNAMESE 
C1561452|T098||CDC|-- VIETNAMESE
C1561452|T098||CDC|VIETNAMESE RACE
C1553323|T098||CDC|CAMBODIAN
C1553323|T098||CDC|KAMPUCHEAN
C1553323|T098||CDC|CAMBODIANS
C0337894|T098||CDC|BHUTANESE
C0337894|T098||CDC|BHUTANESE 
C1556096|T098||CDC|TAIWANESE
C1556096|T098||CDC|TAIWANESE 
C1556096|T098||CDC|RACE - TAIWANESE
C1556107|T098||CDC|BANGLADESHI
C1556107|T098||CDC|BANGLADESHI RACE
C0425375|T098||CDC|PAKISTANI
C0425375|T098||CDC|RACE: PAKISTANI
C0425375|T098||CDC|RACE: PAKISTANI 
C0425375|T098||CDC|PAKISTANI RACE
C0240293|T098||CDC|MALAYSIAN
C0240293|T098||CDC|MALAYSIAN RACE
C1524069|T098||CDC|INDIAN
C1524069|T098||CDC|INDIAN (EAST INDIAN)
C1524069|T098||CDC|INDIAN 
C1524069|T098||CDC|INDIAN RACE 
C1524069|T098||CDC|INDIAN SUB-CONTINENT (NMO)
C1524069|T098||CDC|INDIAN RACE
C1524069|T098||CDC|INDIAN SUB-CONTINENT (NMO) 
C1524069|T098||CDC|ASIAN INDIAN
C1524069|T098||CDC|-- ASIAN INDIAN
C1524069|T098||CDC|INDIAN (EAST INDIAN) 
C1524069|T098||CDC|ASIAN INDIANS
C1524069|T098||CDC|INDIAN (RACIAL GROUP)
C1553324|T098||CDC|HMONG
C1553328|T098||CDC|IWO JIMAN
C1553328|T098||CDC|IWO JIMAN RACE
C1553325|T098||CDC|LAOTIAN
C1553325|T098||CDC|LAOTIAN RACE
C1553329|T098||CDC|MALDIVIAN
C1553329|T098||CDC|MALDIVIAN RACE
C1553330|T098||CDC|NEPALESE
C1553330|T098||CDC|NEPALESE RACE
C1553326|T098||CDC|OKINAWAN
C1553326|T098||CDC|OKINAWAN RACE
C1553331|T098||CDC|SINGAPOREAN
C1553331|T098||CDC|SINGAPOREAN RACE
C1553327|T098||CDC|SRI LANKAN
C1553327|T098||CDC|SRI LANKAN RACE
C0337893|T098||CDC|AINU
C0337893|T098||CDC|AINU 
C0337892|T098||CDC|MONGOLOID POPULATION
C0337892|T098||CDC|MONGOL 
C0337892|T098||CDC|MONGOLOID
C0337892|T098||CDC|MONGOLOID 
C0337892|T098||CDC|MONGOL
C0337892|T098||CDC|MONGOLOID RACE
C0337892|T098||CDC|ASIATIC RACE
C0337892|T098||CDC|ASIATIC RACES
C0337892|T098||CDC|MONGOLOID RACES
C0337892|T098||CDC|RACE, ASIATIC
C0337892|T098||CDC|RACE, MONGOLOID
C0337892|T098||CDC|RACES, ASIATIC
C0337892|T098||CDC|RACES, MONGOLOID
C0337892|T098||CDC|MONGOLOID, NOS
C0337920|T098||CDC|HAWAIIAN
C0337920|T098||CDC|HAWAIIAN POPULATION
C0337920|T098||CDC|NATIVE HAWAIIAN
C0337920|T098||CDC|-- NATIVE HAWAIIAN
C0337920|T098||CDC|HAWAIIAN, NATIVE
C0337920|T098||CDC|HAWAIIANS, NATIVE
C0337920|T098||CDC|NATIVE HAWAIIANS
C0337920|T098||CDC|HAWAIIANS
C0337920|T098||CDC|HAWAIIANS 
C0337920|T098||CDC|HAWAII NATIVES
C1519427|T098||CDC|SOUTH ASIANS
C1519427|T098||CDC|SOUTH ASIAN
C1709065|T098||CDC|MONGOLIAN
C1709065|T098||CDC|MONGOLIAN (RACE)
C0008121|T098||CDC|AMERICAN, CHINESE
C0008121|T098||CDC|AMERICANS, CHINESE
C0008121|T098||CDC|CHINESE AMERICAN
C0008121|T098||CDC|CHINESE AMERICANS
C0022343|T098||CDC|AMERICAN, JAPANESE
C0022343|T098||CDC|AMERICANS, JAPANESE
C0022343|T098||CDC|JAPANESE AMERICAN
C0022343|T098||CDC|JAPANESE AMERICANS
C0597918|T098||CDC|FILIPINO AMERICAN
C0597919|T098||CDC|INDOCHINESE AMERICAN
C0597920|T098||CDC|INDONESIAN AMERICAN
C0597921|T098||CDC|KOREAN AMERICAN
C0597921|T098||CDC|AMERICANS, KOREAN
C0597921|T098||CDC|AMERICAN, KOREAN
C0597921|T098||CDC|KOREAN AMERICANS
C0003988|T098||CDC|AMERICAN, ASIAN
C0003988|T098||CDC|AMERICANS, ASIAN
C0003988|T098||CDC|ASIAN AMERICAN
C0003988|T098||CDC|ASIAN-AMERICAN
C0085756|T098||CDC|AFRICAN AMERICAN
C0085756|T098||CDC|AMERICANS, AFRICAN
C0085756|T098||CDC|AFROAMERICAN
C0085756|T098||CDC|BLACK AMERICAN
C0085756|T098||CDC|RACEBLACKORAFRICANAMERICAN
C0085756|T098||CDC|AFRICAN AMERICANS
# C0085756|T098||CDC|BLACK
C0085756|T098||CDC|BLACK OR AFRICAN AMERICAN
C0085756|T098||CDC|BLACK OR AFRICAN-AMERICAN
C0085756|T098||CDC|AFRICAN-AMERICAN
C0085756|T098||CDC|BLACK/AFRICAN AMERICAN
C0085756|T098||CDC|AFRICAN AMERICAN 
C0085756|T098||CDC|BLACK POPULATIONS
C0085756|T098||CDC|AFRO AMERICAN
C0005680|T098||CDC|BLACK RACE
C0005680|T098||CDC|BLACKS
# C0005680|T098||CDC|BLACK
C0005680|T098||CDC|BLACK - ETHNIC GROUP 
C0005680|T098||CDC|BLACK - ETHNIC GROUP
C0027567|T098||CDC|AFRICAN
C0027567|T098||CDC|AFRICAN RACE 
C0027567|T098||CDC|AFRICAN RACE
# C0027567|T098||CDC|BLACK
C0027567|T098||CDC|AFRICAN RACE (RACIAL GROUP)
C1553338|T098||CDC|DOMINICAN
C1553338|T098||CDC|DOMINICA ISLANDER
C1553338|T098||CDC|DOMINICA ISLANDER RACE
C0239806|T098||CDC|HAITIAN
C0239806|T098||CDC|HAITIAN RACE
C0240072|T098||CDC|JAMAICAN
C1553339|T098||CDC|TOBAGOAN
C1553339|T098||CDC|TOBAGOAN RACE
C1553340|T098||CDC|TRINIDADIAN
C1553340|T098||CDC|TRINIDADIAN RACE
C0425373|T098||CDC|WEST INDIAN
C0425373|T098||CDC|RACE: WEST INDIAN
C0425373|T098||CDC|RACE: WEST INDIAN 
C0425373|T098||CDC|RACE: WEST INDIAN 
C0425373|T098||CDC|WEST INDIAN RACE
C1553336|T098||CDC|BAHAMIAN
C1553336|T098||CDC|BAHAMIAN RACE
C1553337|T098||CDC|BARBADIAN
C1553337|T098||CDC|BARBADIAN RACE
C2135340|T098||CDC|CULTURAL BACKGROUND AFRICAN AMERICAN 
C2135340|T098||CDC|CULTURAL BACKGROUND AFRICAN AMERICAN
C2135340|T098||CDC|THE CULTURAL BACKGROUND IS AFRICAN AMERICAN
C2135340|T098||CDC|SOCIAL HISTORY - CULTURAL BACKGROUND AFRICAN AMERICAN
C0422781|T098||CDC|BLACK - OTHER, MIXED
C0422781|T098||CDC|BLACK - OTHER, MIXED 
C0337824|T098||CDC|BLACK AFRICAN 
C0337824|T098||CDC|BLACK AFRICAN
C0337824|T098||CDC|BLACK AFRICAN, NOS
C0422771|T098||CDC|AFRICAN CARIBBEAN
C0422771|T098||CDC|BLACK CARIB
C0422771|T098||CDC|BLACK CARIBBEAN
C0422771|T098||CDC|BLACK CARIBBEAN 
C0422772|T098||CDC|BLACK, OTHER, NON-MIXED ORIGIN
C0422772|T098||CDC|BLACK, OTHER, NON-MIXED ORIGIN 
C1278528|T098||CDC|OTHER BLACK ETHNIC GROUP
C1278528|T098||CDC|OTHER BLACK ETHNIC GROUP 
C2135370|T098||CDC|RACIAL BACKGROUND BLACK 
C2135370|T098||CDC|RACIAL BACKGROUND BLACK
C1531522|T098||CDC|BLACK, NOT OF HISPANIC ORIGIN (RACIAL GROUP)
C1531522|T098||CDC|BLACK, NOT OF HISPANIC ORIGIN
C0239304|T098||CDC|ETHIOPIAN
C1556088|T098||CDC|LIBERIAN
C1556088|T098||CDC|LIBERIANS
C1556088|T098||CDC|LIBERIANS 
C1556088|T098||CDC|LIBERIAN RACE
C1553334|T098||CDC|NAMIBIAN
C1553334|T098||CDC|NAMIBIAN RACE
C1556089|T098||CDC|NIGERIAN
C1556089|T098||CDC|NIGERIANS
C1556089|T098||CDC|NIGERIANS 
C1556089|T098||CDC|NIGERIAN RACE
C1553335|T098||CDC|ZAIREAN
C1553335|T098||CDC|ZAIREAN RACE
C1553333|T098||CDC|BOTSWANAN
C1553333|T098||CDC|MOTSWANA
C1553333|T098||CDC|BOTSWANAN RACE
C1553351|T098||CDC|OTHER PACIFIC ISLANDER
C1553351|T098||CDC|-- OTHER PACIFIC ISLANDER
C0337924|T098||CDC|MELANESIAN
C0337924|T098||CDC|RACEPACIFICISLANDMELANESIAN
C0337924|T098||CDC|MELANESIAN, NOS
C0337924|T098||CDC|MELANESIANS
C0337924|T098||CDC|MELANESIANS 
C0337924|T098||CDC|MELANESIAN-PAPUAN
C0337924|T098||CDC|MELANESIAN 
C0240790|T098||CDC|POLYNESIAN
C0240790|T098||CDC|RACEPACIFICISLANDPOLYNESIAN
C0240790|T098||CDC|POLYNESIAN RACE 
C0240790|T098||CDC|POLYNESIAN RACE
C0240790|T098||CDC|POLYNESIAN, NOS
C0240790|T098||CDC|POLYNESIANS
C0240790|T098||CDC|POLYNESIANS 
C1556099|T098||CDC|MICRONESIAN
C1556099|T098||CDC|RACEPACIFICISLANDMICRONESIAN
C1556099|T098||CDC|MICRONESIAN RACE 
C1556099|T098||CDC|MICRONESIAN RACE
C1556099|T098||CDC|MICRONESIAN, NOS
C1556099|T098||CDC|MICRONESIANS
C1556099|T098||CDC|MICRONESIANS 
C0221786|T098||CDC|CAUCASIAN AMERICAN
C0221786|T098||CDC|WHITE AMERICAN
C0337815|T098||CDC|POLES
C0337815|T098||CDC|POLES 
C0337799|T098||CDC|CZECHS
C0337799|T098||CDC|CZECHS 
C1556085|T098||CDC|GERMAN
C1556085|T098||CDC|GERMANS
C1556085|T098||CDC|GERMANS 
C1556085|T098||CDC|GERMAN RACE
C0337800|T098||CDC|DANES
C0337800|T098||CDC|DANES 
C0337796|T098||CDC|BASQUES
C0337796|T098||CDC|BASQUES 
C0337806|T098||CDC|GREEK
C0337806|T098||CDC|GREEKS
C0337806|T098||CDC|GREEKS 
C1556083|T098||CDC|ENGLISH
C1556083|T098||CDC|ENGLISH 
C1556083|T098||CDC|ENGLISH RACE
C0337795|T098||CDC|AUSTRIANS
C0337795|T098||CDC|AUSTRIANS 
C1556087|T098||CDC|IRAQI
C1556087|T098||CDC|IRAQI 
C1556087|T098||CDC|IRAQI RACE
C0337811|T098||CDC|IRANI
C0337811|T098||CDC|IRANI 
C0337817|T098||CDC|SPANIARDS
C0337817|T098||CDC|SPANIARDS 
C0337817|T098||CDC|SPANIARD
C0337797|T098||CDC|BELGIANS
C0337797|T098||CDC|BELGIANS 
C0337801|T098||CDC|EGYPTIAN
C0337801|T098||CDC|EGYPTIANS
C0337801|T098||CDC|EGYPTIANS 
C0032730|T098||CDC|PORTUGUESE POPULATION
C0032730|T098||CDC|PORTUGUESE
C0032730|T098||CDC|PORTUGUESE 
C0337802|T098||CDC|ESTONIANS
C0337802|T098||CDC|ESTONIANS 
C0013331|T098||CDC|DUTCH POPULATION
C0013331|T098||CDC|DUTCH
C0013331|T098||CDC|DUTCH 
C0337809|T098||CDC|INDIANS (HINDI-SPEAKING)
C0337809|T098||CDC|INDIANS (HINDI-SPEAKING) 
C0337798|T098||CDC|BULGARIANS
C0337798|T098||CDC|BULGARIANS 
C0337821|T098||CDC|SERBS
C0337821|T098||CDC|SERBS 
C0241315|T098||CDC|SWISS
C0241315|T098||CDC|SWISS 
C0337816|T098||CDC|RUSSIAN
C0337816|T098||CDC|RUSSIANS
C0337816|T098||CDC|RUSSIANS 
C1556084|T098||CDC|FRENCH
C1556084|T098||CDC|FRENCH 
C1556084|T098||CDC|FRENCH RACE
C0337804|T098||CDC|GEORGIANS
C0337804|T098||CDC|GEORGIANS 
C0337820|T098||CDC|TRISTAN DA CUNHANS
C0337820|T098||CDC|TRISTAN DA CUNHANS 
C0337818|T098||CDC|SWEDES
C0337818|T098||CDC|SWEDES 
C0337808|T098||CDC|ICELANDERS
C0337808|T098||CDC|ICELANDERS 
C0337819|T098||CDC|SYRIAN
C0337819|T098||CDC|SYRIANS 
C0337819|T098||CDC|SYRIANS
C0337822|T098||CDC|SLOVAKS
C0337822|T098||CDC|SLOVAKS 
C0337812|T098||CDC|NORWEGIAN
C0337812|T098||CDC|NORWEGIANS
C0337812|T098||CDC|NORWEGIANS 
C0043114|T098||CDC|WELSH POPULATION
C0043114|T098||CDC|WELSH
C0043114|T098||CDC|WELSH 
C0337803|T098||CDC|FINNS
C0337803|T098||CDC|FINNS 
C1278525|T098||CDC|OTHER WHITE ETHNIC GROUP 
C1278525|T098||CDC|OTHER WHITE ETHNIC GROUP
C0043157|T098||CDC|CAUCASIANS
C0043157|T098||CDC|CAUCASIAN
C0043157|T098||CDC|RACEWHITE
C0043157|T098||CDC|CAUCASIAN (LIVING ORGANISM) 
C0043157|T098||CDC|WHITE - ETHNIC GROUP 
C0043157|T098||CDC|WHITE - ETHNIC GROUP
# C0043157|T098||CDC|WHITE
C0043157|T098||CDC|WHITE/CAUCASIAN
C0043157|T098||CDC|CAUCASIAN/WHITE
C0043157|T098||CDC|CAUCASIAN-WHITE
# C0043157|T098||CDC|WHITES
C0043157|T098||CDC|CAUCASOID
C0043157|T098||CDC|CAUCASIAN 
C0043157|T098||CDC|CAUCASIAN, NOS
C0043157|T098||CDC|CAUCASIAN 
C1278523|T098||CDC|WHITE BRITISH 
C1278523|T098||CDC|WHITE BRITISH
C1278524|T098||CDC|WHITE IRISH 
C1278524|T098||CDC|WHITE IRISH
C0870136|T098||CDC|ANGLOS
C0007457|T098||CDC|CAUCASOID RACE
C0007457|T098||CDC|WHITE RACE
C0007457|T098||CDC|RACIAL BACKGROUND CAUCASIAN
C0007457|T098||CDC|RACIAL BACKGROUND CAUCASIAN 
C0007457|T098||CDC|RACE: CAUCASIAN
C0007457|T098||CDC|CAUCASIAN RACE
C0007457|T098||CDC|RACE: CAUCASIAN (RACIAL GROUP)
C0007457|T098||CDC|RACE: CAUCASIAN 
C0007457|T098||CDC|RACE: WHITE
C0007457|T098||CDC|CAUCASOID
# C0007457|T098||CDC|WHITE
C0007457|T098||CDC|CAUCASIAN RACES
C0007457|T098||CDC|CAUCASOID RACES
C0007457|T098||CDC|RACE, CAUCASIAN
C0007457|T098||CDC|RACE, CAUCASOID
C0007457|T098||CDC|RACES, CAUCASIAN
C0007457|T098||CDC|RACES, CAUCASOID
C0007457|T098||CDC|CAUCASIAN
# C0007457|T098||CDC|WHITES
C0007457|T098||CDC|CAUCASIANS
C0007457|T098||CDC|OCCIDENTAL
C0007457|T098||CDC|CAUCASIAN (RACIAL GROUP)
C0239307|T098||CDC|EUROPEAN
C0239307|T098||CDC|EUROPEAN 
C0239307|T098||CDC|ETHNIC EUROPEAN
C0337794|T098||CDC|ARMENIAN
C0337794|T098||CDC|ARMENIANS
C0337794|T098||CDC|ARMENIANS 
C0087186|T098||CDC|IRISH
C0087186|T098||CDC|IRISH RACE
C0337810|T098||CDC|ITALIAN
C0337810|T098||CDC|ITALIANS
C0337810|T098||CDC|ITALIANS 
C0220896|T098||CDC|POLISH POPULATION
C0220896|T098||CDC|POLISH
C0240966|T098||CDC|SCOTTISH
C0240966|T098||CDC|SCOTTISH RACE
C1710263|T098||CDC|SWEDISH
C1710525|T098||CDC|UKRANIAN
C1711254|T098||CDC|FINNISH
C0019576|T098||CDC|AMERICAN, HISPANIC
C0019576|T098||CDC|AMERICANS, HISPANIC
C0019576|T098||CDC|AMERICANS, SPANISH
C0019576|T098||CDC|HISPANIC AMERICAN
C0019576|T098||CDC|HISPANIC AMERICANS
C0019576|T098||CDC|SPANISH AMERICAN
C0019576|T098||CDC|SPANISH AMERICANS
C1553379|T098||CDC|CUBAN
C1553379|T098||CDC|-- CUBAN
C3829110|T098||CDC|MEXICAN OR MEXICAN AMERICAN
C3828691|T098||CDC|OTHER HISPANIC OR LATINO(A)
C3161473|T098||CDC|SPANISH
C3161473|T098||CDC|SPANISH PERSON
C0086409|T098||CDC|HISPANIC
C0086409|T098||CDC|HISPANICS
C0086409|T098||CDC|HISPANIC OR LATINO
C0086409|T098||CDC|ETHNICITYHISPANIC
C0086409|T098||CDC|HISPANIC ORIGIN
C0086409|T098||CDC|SPANISH
C0086409|T098||CDC|HISPANIC POPULATIONS
C0086409|T098||CDC|HISPANICS OR LATINOS
C0086409|T098||CDC|LATINO POPULATION
C0086409|T098||CDC|SPANISH ORIGIN
C0086409|T098||CDC|HISPANIC (RACIAL GROUP)
C0025884|T098||CDC|AMERICAN, MEXICAN
C0025884|T098||CDC|AMERICANS, MEXICAN
C0025884|T098||CDC|CHICANO
C0025884|T098||CDC|MEXICAN AMERICAN
C0025884|T098||CDC|MEXICAN AMERICANS
C0025884|T098||CDC|CHICANOS
C0025884|T098||CDC|CHICANAS
C0025884|T098||CDC|CHICANA
C0010436|T098||CDC|AMERICANS, CUBAN
C0010436|T098||CDC|CUBAN AMERICAN
C0010436|T098||CDC|CUBAN AMERICANS
C0086528|T098||CDC|LATINO
C0086528|T098||CDC|LATINOS
C0034043|T098||CDC|PUERTO RICAN
C0034043|T098||CDC|PUERTORICAN
C0034043|T098||CDC|-- PUERTO RICAN
C0034043|T098||CDC|PUERTO RICANS
C0935556|T098||CDC|LATINOS/LATINAS
C1533018|T098||CDC|HISPANIC, BLACK (RACIAL GROUP)
C1533018|T098||CDC|HISPANIC, BLACK
C1533018|T098||CDC|HISPANIC BLACK RACIAL GROUP
C1533019|T098||CDC|HISPANIC, COLOR UNKNOWN (RACIAL GROUP)
C1533019|T098||CDC|HISPANIC, COLOR UNKNOWN
C1533019|T098||CDC|HISPANIC, COLOUR UNKNOWN
C1533021|T098||CDC|HISPANIC, WHITE (RACIAL GROUP)
C1533021|T098||CDC|HISPANIC, WHITE
C1533021|T098||CDC|HISPANIC WHITE RACIAL GROUP
C0425359|T098||CDC|SOUTH AMERICAN
C0425359|T098||CDC|-- SOUTH AMERICAN
C0240339|T098||CDC|MEXICAN
C0240339|T098||CDC|ETHNICITYHISPANICMEXICAN
C0240339|T098||CDC|-- MEXICAN
C0238914|T098||CDC|CENTRAL AMERICAN
C0238914|T098||CDC|ETHNICITYHISPANICCENTRALAMERICAN
C0238914|T098||CDC|-- CENTRAL AMERICAN
C1328872|T098||CDC|DOMINICAN
C1328872|T098||CDC|DOMINICAN - ETHNICITY
C1553378|T098||CDC|LATIN AMERICAN
C1881927|T098||CDC|MULTIPLE HISPANIC
C1880193|T098||CDC|CUBAN OR CUBAN AMERICAN
C2135343|T098||CDC|CULTURAL BACKGROUND HISPANIC 
C2135343|T098||CDC|THE CULTURAL BACKGROUND IS HISPANIC
C2135343|T098||CDC|CULTURAL BACKGROUND HISPANIC
C2741637|T098||CDC|HISPANIC OR LATINO:FINDING:POINT IN TIME:^PATIENT:ORDINAL
C2741637|T098||CDC|HISPANIC OR LATINO
C2741637|T098||CDC|HISPANIC OR LATINO:FIND:PT:^PATIENT:ORD
