C0032181|T034||LNC|BLOOD PLATELET COUNTS
C0005821|T034|MTHU008063|LNC|BLOOD PLATELETS|THROMBOCYTE (PLATELET)
C0200642|T034||LNC|PLATELET ESTIMATE
C1254925|T034||LNC|OPERATING ROOM MISC LABS: PLATELETS
C0032181|T034||LNC|BLOOD PLATELET COUNTS
C0032181|T034||LNC|BLOOD PLATELET NUMBERS
C0032181|T034||LNC|COUNT, BLOOD PLATELET
C0032181|T034||LNC|COUNT, PLATELET
C0032181|T034||LNC|COUNTS, BLOOD PLATELET
C0032181|T034||LNC|COUNTS, PLATELET
C0032181|T034||LNC|NUMBER, BLOOD PLATELET
C0032181|T034||LNC|NUMBER, PLATELET
C0032181|T034||LNC|NUMBERS, BLOOD PLATELET
C0032181|T034||LNC|NUMBERS, PLATELET
C0032181|T034||LNC|PLATELET COUNT
C0032181|T034||LNC|PLATELET COUNT, BLOOD
C0032181|T034||LNC|PLATELET COUNTS
C0032181|T034||LNC|PLATELET COUNTS, BLOOD
C0032181|T034||LNC|PLATELET NUMBER, BLOOD
C0032181|T034||LNC|PLATELET NUMBERS
C0032181|T034||LNC|PLATELET NUMBERS, BLOOD
C0032181|T034||LNC|PLATELETS
C0032181|T034||LNC|PLATELET COUNT 
C0032181|T034||LNC|PLATELET COUNT NOS 
C0032181|T034||LNC|PLATELET COUNT NOS
C0032181|T034||LNC|PLATELET COUNT 
C0032181|T034||LNC|PLAT
C0032181|T034||LNC|ANUCLEATED THROMBOCYTES
C0032181|T034||LNC|THROMBOCYTE COUNT
C0032181|T034||LNC|PLATELET NUMBER
C0032181|T034||LNC|BLOOD PLATELET COUNT
C0032181|T034||LNC|BLOOD PLATELET NUMBER
C0032181|T034||LNC|WHOLE BLOOD PLATELET COUNTS
C0032181|T034||LNC|PLT - PLATELET COUNT
C0032181|T034||LNC|PLATELET COUNT - OBSERVATION
C0032181|T034||LNC|PLATELET COUNT MEASUREMENT
C2082381|T034||LNC|PLASMA PLATELET COUNT
C2082381|T034||LNC|PLASMA PLATELET COUNT 
C0523117|T034||LNC|MANUAL PLATELET COUNT 
C0523117|T034||LNC|MANUAL PLATELET COUNT
C0523117|T034||LNC|PLATELET COUNT, BLOOD, MANUAL
C0523117|T034||LNC|PLATELET COUNT, BLOOD, MANUAL 
C1144713|T034||LNC|AUTOMATED PLATELET COUNT
C1144713|T034||LNC|AUTOMATED PLATELET COUNT 
C1144713|T034||LNC|BLOOD COUNT PLATELET AUTOMATED
C1144713|T034||LNC|PLATELET COUNT, AUTOMATED TEST
C1144713|T034||LNC|BLOOD COUNT; PLATELET, AUTOMATED
C0523118|T034||LNC|PLATELET COUNT, BLOOD, AUTOMATED
C0523118|T034||LNC|PLATELET COUNT, BLOOD, AUTOMATED 
C1294068|T034||LNC|PLATELET COUNT, REES-ECKER METHOD 
C1294068|T034||LNC|PLATELET COUNT, REES-ECKER METHOD
C0005821|T034|MTHU008063|LNC|THROMBOCYTE|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|BLOOD PLATELETS|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLATELET|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLATELET, BLOOD|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLATELETS, BLOOD|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|BLOOD PLATELET|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLATELETS|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLATELET |THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLT - PLATELET|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLT - PLATELETS|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLATELET |THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|THROMBOCYTE (PLATELET)|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|DEETJEN BODY|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|BIZZOZERO CORPUSCLE|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|THROMBOCYTES|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLATELET [DUP] |THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|PLATELETS (BLOOD)|THROMBOCYTE (PLATELET)
C0005821|T034|MTHU008063|LNC|RETICULOENDOTHELIAL SYSTEM, PLATELETS|THROMBOCYTE (PLATELET)
C1994889|T034|LP50307-5|LNC|PLATELETS AGRANULAR &#X7C; BLD-SER-PLAS|PLATELETS AGRANULAR &#X7C; BLD-SER-PLAS
C1994885|T034|LP51977-4|LNC|PLATELETS &#X7C; BODY FLUID|PLATELETS &#X7C; BODY FLUID
C1994891|T034|LP49896-1|LNC|PLATELETS LARGE &#X7C; BLD-SER-PLAS|PLATELETS LARGE &#X7C; BLD-SER-PLAS
C3700279|T034|LP181025-0|LNC|PLATELETS &#X7C; BLOOD CAPILLARY|PLATELETS &#X7C; BLOOD CAPILLARY
C1994893|T034|LP49928-2|LNC|PLATELETS SMALL &#X7C; BLD-SER-PLAS|PLATELETS SMALL &#X7C; BLD-SER-PLAS
C1994883|T034|LP41375-4|LNC|PLATELETS &#X7C; BLD-SER-PLAS|PLATELETS &#X7C; BLD-SER-PLAS
C3847483|T034|LP184163-6|LNC|PLATELETS &#X7C; PLATELET RICH PLASMA|PLATELETS &#X7C; PLATELET RICH PLASMA
