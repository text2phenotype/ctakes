//CUI|TUI|TTY|CODE|SAB|STR|PREF
C0078988|T098|LN|2028-9|LNC|carbon dioxide|carbon dioxide
C0078988|T098|MTH_LN|2028-9|LNC|carbon dioxide|carbon dioxide
C0078988|T098|OSN|2028-9|LNC|carbon dioxide|carbon dioxide
C0078988|T098|LC|2028-9|LNC|carbon dioxide|carbon dioxide
C0240790|T098|LN|2078-4|LNC|chloride|chloride
C0240790|T098|MTH_LN|2078-4|LNC|chloride|chloride
C0240790|T098|OSN|2078-4|LNC|chloride|chloride
C0240790|T098|LC|2078-4|LNC|chloride|chloride
C0337928|T098|LC|2091-7|LNC|VLDL cholesterol|VLDL cholesterol
C0337928|T098|MTH_LN|2091-7|LNC|VLDL cholesterol|VLDL cholesterol
C0337928|T098|LN|2091-7|LNC|VLDL cholesterol|VLDL cholesterol
C0337928|T098|OSN|2091-7|LNC|VLDL cholesterol|VLDL cholesterol
C0337928|T098|LC|2091-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0337928|T098|MTH_LN|2091-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0337928|T098|LN|2091-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0337928|T098|OSN|2091-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0337928|T098|LC|2091-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0337928|T098|MTH_LN|2091-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0337928|T098|LN|2091-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0337928|T098|OSN|2091-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0337928|T098|LC|2091-7|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0337928|T098|MTH_LN|2091-7|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0337928|T098|LN|2091-7|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0337928|T098|OSN|2091-7|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0337933|T098|LN|2082-6|LNC|cholesterol|cholesterol
C0337933|T098|MTH_LN|2082-6|LNC|cholesterol|cholesterol
C0337933|T098|OSN|2082-6|LNC|cholesterol|cholesterol
C0337933|T098|LC|2082-6|LNC|cholesterol|cholesterol
C0337933|T098|LN|2082-6|LNC|total cholesterol|total cholesterol
C0337933|T098|MTH_LN|2082-6|LNC|total cholesterol|total cholesterol
C0337933|T098|OSN|2082-6|LNC|total cholesterol|total cholesterol
C0337933|T098|LC|2082-6|LNC|total cholesterol|total cholesterol
C0337933|T098|LN|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C0337933|T098|MTH_LN|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C0337933|T098|OSN|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C0337933|T098|LC|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C0362890|T201|LN|702-1|LNC|Unequal sizered|Unequal sizered
C0362890|T201|MTH_LN|702-1|LNC|Unequal sizered|Unequal sizered
C0362890|T201|OSN|702-1|LNC|Unequal sizered|Unequal sizered
C0362890|T201|LC|702-1|LNC|Unequal sizered|Unequal sizered
C0362892|T201|LN|704-7|LNC|basophil count|basophil count
C0362892|T201|OSN|704-7|LNC|basophil count|basophil count
C0362892|T201|MTH_LN|704-7|LNC|basophil count|basophil count
C0362892|T201|LC|704-7|LNC|basophil count|basophil count
C0362893|T201|LN|705-4|LNC|basophil count|basophil count
C0362893|T201|OSN|705-4|LNC|basophil count|basophil count
C0362893|T201|MTH_LN|705-4|LNC|basophil count|basophil count
C0362893|T201|LC|705-4|LNC|basophil count|basophil count
C0362894|T201|LN|706-2|LNC|basophil count|basophil count
C0362894|T201|MTH_LN|706-2|LNC|basophil count|basophil count
C0362894|T201|OSN|706-2|LNC|basophil count|basophil count
C0362894|T201|LC|706-2|LNC|basophil count|basophil count
C0362895|T201|LN|707-0|LNC|basophil count|basophil count
C0362895|T201|MTH_LN|707-0|LNC|basophil count|basophil count
C0362895|T201|OSN|707-0|LNC|basophil count|basophil count
C0362895|T201|LC|707-0|LNC|basophil count|basophil count
C0362900|T201|LN|711-2|LNC|eosinophil count|eosinophil count
C0362900|T201|OSN|711-2|LNC|eosinophil count|eosinophil count
C0362900|T201|MTH_LN|711-2|LNC|eosinophil count|eosinophil count
C0362900|T201|LC|711-2|LNC|eosinophil count|eosinophil count
C0362900|T201|LN|711-2|LNC|eosinophil morphology|eosinophil morphology
C0362900|T201|OSN|711-2|LNC|eosinophil morphology|eosinophil morphology
C0362900|T201|MTH_LN|711-2|LNC|eosinophil morphology|eosinophil morphology
C0362900|T201|LC|711-2|LNC|eosinophil morphology|eosinophil morphology
C0362900|T201|LN|711-2|LNC|eosinophils|eosinophils
C0362900|T201|OSN|711-2|LNC|eosinophils|eosinophils
C0362900|T201|MTH_LN|711-2|LNC|eosinophils|eosinophils
C0362900|T201|LC|711-2|LNC|eosinophils|eosinophils
C0362901|T201|LN|712-0|LNC|eosinophil count|eosinophil count
C0362901|T201|OSN|712-0|LNC|eosinophil count|eosinophil count
C0362901|T201|MTH_LN|712-0|LNC|eosinophil count|eosinophil count
C0362901|T201|LC|712-0|LNC|eosinophil count|eosinophil count
C0362901|T201|LN|712-0|LNC|eosinophil morphology|eosinophil morphology
C0362901|T201|OSN|712-0|LNC|eosinophil morphology|eosinophil morphology
C0362901|T201|MTH_LN|712-0|LNC|eosinophil morphology|eosinophil morphology
C0362901|T201|LC|712-0|LNC|eosinophil morphology|eosinophil morphology
C0362901|T201|LN|712-0|LNC|eosinophils|eosinophils
C0362901|T201|OSN|712-0|LNC|eosinophils|eosinophils
C0362901|T201|MTH_LN|712-0|LNC|eosinophils|eosinophils
C0362901|T201|LC|712-0|LNC|eosinophils|eosinophils
C0362902|T201|LN|713-8|LNC|eosinophil count|eosinophil count
C0362902|T201|MTH_LN|713-8|LNC|eosinophil count|eosinophil count
C0362902|T201|OSN|713-8|LNC|eosinophil count|eosinophil count
C0362902|T201|LC|713-8|LNC|eosinophil count|eosinophil count
C0362902|T201|LN|713-8|LNC|eosinophil morphology|eosinophil morphology
C0362902|T201|MTH_LN|713-8|LNC|eosinophil morphology|eosinophil morphology
C0362902|T201|OSN|713-8|LNC|eosinophil morphology|eosinophil morphology
C0362902|T201|LC|713-8|LNC|eosinophil morphology|eosinophil morphology
C0362902|T201|LN|713-8|LNC|eosinophils|eosinophils
C0362902|T201|MTH_LN|713-8|LNC|eosinophils|eosinophils
C0362902|T201|OSN|713-8|LNC|eosinophils|eosinophils
C0362902|T201|LC|713-8|LNC|eosinophils|eosinophils
C0362903|T201|LN|714-6|LNC|eosinophil count|eosinophil count
C0362903|T201|MTH_LN|714-6|LNC|eosinophil count|eosinophil count
C0362903|T201|OSN|714-6|LNC|eosinophil count|eosinophil count
C0362903|T201|LC|714-6|LNC|eosinophil count|eosinophil count
C0362903|T201|LN|714-6|LNC|eosinophil morphology|eosinophil morphology
C0362903|T201|MTH_LN|714-6|LNC|eosinophil morphology|eosinophil morphology
C0362903|T201|OSN|714-6|LNC|eosinophil morphology|eosinophil morphology
C0362903|T201|LC|714-6|LNC|eosinophil morphology|eosinophil morphology
C0362903|T201|LN|714-6|LNC|eosinophils|eosinophils
C0362903|T201|MTH_LN|714-6|LNC|eosinophils|eosinophils
C0362903|T201|OSN|714-6|LNC|eosinophils|eosinophils
C0362903|T201|LC|714-6|LNC|eosinophils|eosinophils
C0362905|T201|LN|784-9|LNC|erythrocyte volume|erythrocyte volume
C0362905|T201|MTH_LN|784-9|LNC|erythrocyte volume|erythrocyte volume
C0362905|T201|OSN|784-9|LNC|erythrocyte volume|erythrocyte volume
C0362905|T201|LC|784-9|LNC|erythrocyte volume|erythrocyte volume
C0362905|T201|LN|784-9|LNC|mean corpuscular volume|mean corpuscular volume
C0362905|T201|MTH_LN|784-9|LNC|mean corpuscular volume|mean corpuscular volume
C0362905|T201|OSN|784-9|LNC|mean corpuscular volume|mean corpuscular volume
C0362905|T201|LC|784-9|LNC|mean corpuscular volume|mean corpuscular volume
C0362906|T201|LN|785-6|LNC|MCH|MCH
C0362906|T201|LC|785-6|LNC|MCH|MCH
C0362906|T201|MTH_LN|785-6|LNC|MCH|MCH
C0362906|T201|OSN|785-6|LNC|MCH|MCH
C0362906|T201|LN|785-6|LNC|mean corpuscular hemoglobin|mean corpuscular hemoglobin
C0362906|T201|LC|785-6|LNC|mean corpuscular hemoglobin|mean corpuscular hemoglobin
C0362906|T201|MTH_LN|785-6|LNC|mean corpuscular hemoglobin|mean corpuscular hemoglobin
C0362906|T201|OSN|785-6|LNC|mean corpuscular hemoglobin|mean corpuscular hemoglobin
C0362906|T201|LN|785-6|LNC|mean corpuscular haemoglobin|mean corpuscular haemoglobin
C0362906|T201|LC|785-6|LNC|mean corpuscular haemoglobin|mean corpuscular haemoglobin
C0362906|T201|MTH_LN|785-6|LNC|mean corpuscular haemoglobin|mean corpuscular haemoglobin
C0362906|T201|OSN|785-6|LNC|mean corpuscular haemoglobin|mean corpuscular haemoglobin
C0362907|T201|LN|786-4|LNC|MCH|MCH
C0362907|T201|MTH_LN|786-4|LNC|MCH|MCH
C0362907|T201|LC|786-4|LNC|MCH|MCH
C0362907|T201|OSN|786-4|LNC|MCH|MCH
C0362907|T201|LN|786-4|LNC|mean corpuscular hemoglobin|mean corpuscular hemoglobin
C0362907|T201|MTH_LN|786-4|LNC|mean corpuscular hemoglobin|mean corpuscular hemoglobin
C0362907|T201|LC|786-4|LNC|mean corpuscular hemoglobin|mean corpuscular hemoglobin
C0362907|T201|OSN|786-4|LNC|mean corpuscular hemoglobin|mean corpuscular hemoglobin
C0362907|T201|LN|786-4|LNC|mean corpuscular haemoglobin|mean corpuscular haemoglobin
C0362907|T201|MTH_LN|786-4|LNC|mean corpuscular haemoglobin|mean corpuscular haemoglobin
C0362907|T201|LC|786-4|LNC|mean corpuscular haemoglobin|mean corpuscular haemoglobin
C0362907|T201|OSN|786-4|LNC|mean corpuscular haemoglobin|mean corpuscular haemoglobin
C0362908|T201|LN|787-2|LNC|erythrocyte volume|erythrocyte volume
C0362908|T201|MTH_LN|787-2|LNC|erythrocyte volume|erythrocyte volume
C0362908|T201|LC|787-2|LNC|erythrocyte volume|erythrocyte volume
C0362908|T201|OSN|787-2|LNC|erythrocyte volume|erythrocyte volume
C0362908|T201|LN|787-2|LNC|mean corpuscular volume|mean corpuscular volume
C0362908|T201|MTH_LN|787-2|LNC|mean corpuscular volume|mean corpuscular volume
C0362908|T201|LC|787-2|LNC|mean corpuscular volume|mean corpuscular volume
C0362908|T201|OSN|787-2|LNC|mean corpuscular volume|mean corpuscular volume
// C0362919|T201|LN|798-9|LNC||
// C0362919|T201|OSN|798-9|LNC||
// C0362919|T201|MTH_LN|798-9|LNC||
// C0362919|T201|LC|798-9|LNC||
C0362919|T201|LN|798-9|LNC|occult|occult
C0362919|T201|OSN|798-9|LNC|occult|occult
C0362919|T201|MTH_LN|798-9|LNC|occult|occult
C0362919|T201|LC|798-9|LNC|occult|occult
// C0362920|T201|LN|799-7|LNC||
// C0362920|T201|OSN|799-7|LNC||
// C0362920|T201|MTH_LN|799-7|LNC||
// C0362920|T201|LC|799-7|LNC||
C0362920|T201|LN|799-7|LNC|occult|occult
C0362920|T201|OSN|799-7|LNC|occult|occult
C0362920|T201|MTH_LN|799-7|LNC|occult|occult
C0362920|T201|LC|799-7|LNC|occult|occult
C0362926|T201|LN|721-1|LNC|hemoglobin|hemoglobin
C0362926|T201|OSN|721-1|LNC|hemoglobin|hemoglobin
C0362926|T201|MTH_LN|721-1|LNC|hemoglobin|hemoglobin
C0362926|T201|LC|721-1|LNC|hemoglobin|hemoglobin
C0362930|T201|LN|725-2|LNC|Hemoglobin|Hemoglobin
C0362930|T201|MTH_LN|725-2|LNC|Hemoglobin|Hemoglobin
C0362930|T201|OSN|725-2|LNC|Hemoglobin|Hemoglobin
C0362930|T201|LC|725-2|LNC|Hemoglobin|Hemoglobin
C0362931|T201|LN|726-0|LNC|Hemoglobin|Hemoglobin
C0362931|T201|MTH_LN|726-0|LNC|Hemoglobin|Hemoglobin
C0362931|T201|OSN|726-0|LNC|Hemoglobin|Hemoglobin
C0362931|T201|LC|726-0|LNC|Hemoglobin|Hemoglobin
C0362947|T201|LN|731-0|LNC|lymphocyte count|lymphocyte count
C0362947|T201|OSN|731-0|LNC|lymphocyte count|lymphocyte count
C0362947|T201|MTH_LN|731-0|LNC|lymphocyte count|lymphocyte count
C0362947|T201|LC|731-0|LNC|lymphocyte count|lymphocyte count
C0362947|T201|LN|731-0|LNC|lymphocyte number|lymphocyte number
C0362947|T201|OSN|731-0|LNC|lymphocyte number|lymphocyte number
C0362947|T201|MTH_LN|731-0|LNC|lymphocyte number|lymphocyte number
C0362947|T201|LC|731-0|LNC|lymphocyte number|lymphocyte number
C0362947|T201|LN|731-0|LNC|lymphocyte counts|lymphocyte counts
C0362947|T201|OSN|731-0|LNC|lymphocyte counts|lymphocyte counts
C0362947|T201|MTH_LN|731-0|LNC|lymphocyte counts|lymphocyte counts
C0362947|T201|LC|731-0|LNC|lymphocyte counts|lymphocyte counts
C0362947|T201|LN|731-0|LNC|lymphocytes|lymphocytes
C0362947|T201|OSN|731-0|LNC|lymphocytes|lymphocytes
C0362947|T201|MTH_LN|731-0|LNC|lymphocytes|lymphocytes
C0362947|T201|LC|731-0|LNC|lymphocytes|lymphocytes
C0362947|T201|LN|731-0|LNC|numberslymphocytes|numberslymphocytes
C0362947|T201|OSN|731-0|LNC|numberslymphocytes|numberslymphocytes
C0362947|T201|MTH_LN|731-0|LNC|numberslymphocytes|numberslymphocytes
C0362947|T201|LC|731-0|LNC|numberslymphocytes|numberslymphocytes
C0362951|T201|LN|735-1|LNC|lymphocytes|lymphocytes
C0362951|T201|OSN|735-1|LNC|lymphocytes|lymphocytes
C0362951|T201|LC|735-1|LNC|lymphocytes|lymphocytes
C0362951|T201|MTH_LN|735-1|LNC|lymphocytes|lymphocytes
C0362951|T201|LN|735-1|LNC|lymphoid lineage|lymphoid lineage
C0362951|T201|OSN|735-1|LNC|lymphoid lineage|lymphoid lineage
C0362951|T201|LC|735-1|LNC|lymphoid lineage|lymphoid lineage
C0362951|T201|MTH_LN|735-1|LNC|lymphoid lineage|lymphoid lineage
C0362951|T201|LN|735-1|LNC|lymphocyte morphology|lymphocyte morphology
C0362951|T201|OSN|735-1|LNC|lymphocyte morphology|lymphocyte morphology
C0362951|T201|LC|735-1|LNC|lymphocyte morphology|lymphocyte morphology
C0362951|T201|MTH_LN|735-1|LNC|lymphocyte morphology|lymphocyte morphology
C0362952|T201|LN|736-9|LNC|lymphocyte count|lymphocyte count
C0362952|T201|MTH_LN|736-9|LNC|lymphocyte count|lymphocyte count
C0362952|T201|OSN|736-9|LNC|lymphocyte count|lymphocyte count
C0362952|T201|LC|736-9|LNC|lymphocyte count|lymphocyte count
C0362952|T201|LN|736-9|LNC|lymphocyte number|lymphocyte number
C0362952|T201|MTH_LN|736-9|LNC|lymphocyte number|lymphocyte number
C0362952|T201|OSN|736-9|LNC|lymphocyte number|lymphocyte number
C0362952|T201|LC|736-9|LNC|lymphocyte number|lymphocyte number
C0362952|T201|LN|736-9|LNC|lymphocyte counts|lymphocyte counts
C0362952|T201|MTH_LN|736-9|LNC|lymphocyte counts|lymphocyte counts
C0362952|T201|OSN|736-9|LNC|lymphocyte counts|lymphocyte counts
C0362952|T201|LC|736-9|LNC|lymphocyte counts|lymphocyte counts
C0362952|T201|LN|736-9|LNC|lymphocytes|lymphocytes
C0362952|T201|MTH_LN|736-9|LNC|lymphocytes|lymphocytes
C0362952|T201|OSN|736-9|LNC|lymphocytes|lymphocytes
C0362952|T201|LC|736-9|LNC|lymphocytes|lymphocytes
C0362952|T201|LN|736-9|LNC|numberslymphocytes|numberslymphocytes
C0362952|T201|MTH_LN|736-9|LNC|numberslymphocytes|numberslymphocytes
C0362952|T201|OSN|736-9|LNC|numberslymphocytes|numberslymphocytes
C0362952|T201|LC|736-9|LNC|numberslymphocytes|numberslymphocytes
C0362953|T201|LN|737-7|LNC|lymphocyte count|lymphocyte count
C0362953|T201|MTH_LN|737-7|LNC|lymphocyte count|lymphocyte count
C0362953|T201|OSN|737-7|LNC|lymphocyte count|lymphocyte count
C0362953|T201|LC|737-7|LNC|lymphocyte count|lymphocyte count
C0362953|T201|LN|737-7|LNC|lymphocyte number|lymphocyte number
C0362953|T201|MTH_LN|737-7|LNC|lymphocyte number|lymphocyte number
C0362953|T201|OSN|737-7|LNC|lymphocyte number|lymphocyte number
C0362953|T201|LC|737-7|LNC|lymphocyte number|lymphocyte number
C0362953|T201|LN|737-7|LNC|lymphocyte counts|lymphocyte counts
C0362953|T201|MTH_LN|737-7|LNC|lymphocyte counts|lymphocyte counts
C0362953|T201|OSN|737-7|LNC|lymphocyte counts|lymphocyte counts
C0362953|T201|LC|737-7|LNC|lymphocyte counts|lymphocyte counts
C0362953|T201|LN|737-7|LNC|lymphocytes|lymphocytes
C0362953|T201|MTH_LN|737-7|LNC|lymphocytes|lymphocytes
C0362953|T201|OSN|737-7|LNC|lymphocytes|lymphocytes
C0362953|T201|LC|737-7|LNC|lymphocytes|lymphocytes
C0362953|T201|LN|737-7|LNC|numberslymphocytes|numberslymphocytes
C0362953|T201|MTH_LN|737-7|LNC|numberslymphocytes|numberslymphocytes
C0362953|T201|OSN|737-7|LNC|numberslymphocytes|numberslymphocytes
C0362953|T201|LC|737-7|LNC|numberslymphocytes|numberslymphocytes
C0362955|T201|LN|739-3|LNC|granulocyte precursors|granulocyte precursors
C0362955|T201|OSN|739-3|LNC|granulocyte precursors|granulocyte precursors
C0362955|T201|MTH_LN|739-3|LNC|granulocyte precursors|granulocyte precursors
C0362955|T201|LC|739-3|LNC|granulocyte precursors|granulocyte precursors
C0362956|T201|LN|740-1|LNC|granulocyte precursors|granulocyte precursors
C0362956|T201|MTH_LN|740-1|LNC|granulocyte precursors|granulocyte precursors
C0362956|T201|OSN|740-1|LNC|granulocyte precursors|granulocyte precursors
C0362956|T201|LC|740-1|LNC|granulocyte precursors|granulocyte precursors
C0362958|T201|LN|742-7|LNC|monocyte number|monocyte number
C0362958|T201|OSN|742-7|LNC|monocyte number|monocyte number
C0362958|T201|MTH_LN|742-7|LNC|monocyte number|monocyte number
C0362958|T201|LC|742-7|LNC|monocyte number|monocyte number
C0362958|T201|LN|742-7|LNC|monocyte count|monocyte count
C0362958|T201|OSN|742-7|LNC|monocyte count|monocyte count
C0362958|T201|MTH_LN|742-7|LNC|monocyte count|monocyte count
C0362958|T201|LC|742-7|LNC|monocyte count|monocyte count
C0362960|T201|LN|5905-5|LNC|monocyte number|monocyte number
C0362960|T201|MTH_LN|5905-5|LNC|monocyte number|monocyte number
C0362960|T201|OSN|5905-5|LNC|monocyte number|monocyte number
C0362960|T201|LC|5905-5|LNC|monocyte number|monocyte number
C0362960|T201|LN|5905-5|LNC|monocyte count|monocyte count
C0362960|T201|MTH_LN|5905-5|LNC|monocyte count|monocyte count
C0362960|T201|OSN|5905-5|LNC|monocyte count|monocyte count
C0362960|T201|LC|5905-5|LNC|monocyte count|monocyte count
C0362961|T201|LN|744-3|LNC|monocyte number|monocyte number
C0362961|T201|MTH_LN|744-3|LNC|monocyte number|monocyte number
C0362961|T201|OSN|744-3|LNC|monocyte number|monocyte number
C0362961|T201|LC|744-3|LNC|monocyte number|monocyte number
C0362961|T201|LN|744-3|LNC|monocyte count|monocyte count
C0362961|T201|MTH_LN|744-3|LNC|monocyte count|monocyte count
C0362961|T201|OSN|744-3|LNC|monocyte count|monocyte count
C0362961|T201|LC|744-3|LNC|monocyte count|monocyte count
C0362965|T201|LN|748-4|LNC|myeloid leukocytes|myeloid leukocytes
C0362965|T201|OSN|748-4|LNC|myeloid leukocytes|myeloid leukocytes
C0362965|T201|MTH_LN|748-4|LNC|myeloid leukocytes|myeloid leukocytes
C0362965|T201|LC|748-4|LNC|myeloid leukocytes|myeloid leukocytes
C0362967|T201|LN|749-2|LNC|myeloid leukocytes|myeloid leukocytes
C0362967|T201|MTH_LN|749-2|LNC|myeloid leukocytes|myeloid leukocytes
C0362967|T201|OSN|749-2|LNC|myeloid leukocytes|myeloid leukocytes
C0362967|T201|LC|749-2|LNC|myeloid leukocytes|myeloid leukocytes
C0362968|T201|OSN|751-8|LNC|neutrophil counts|neutrophil counts
C0362968|T201|LN|751-8|LNC|neutrophil counts|neutrophil counts
C0362968|T201|MTH_LN|751-8|LNC|neutrophil counts|neutrophil counts
C0362968|T201|LC|751-8|LNC|neutrophil counts|neutrophil counts
C0362968|T201|OSN|751-8|LNC|neutrophil count|neutrophil count
C0362968|T201|LN|751-8|LNC|neutrophil count|neutrophil count
C0362968|T201|MTH_LN|751-8|LNC|neutrophil count|neutrophil count
C0362968|T201|LC|751-8|LNC|neutrophil count|neutrophil count
C0362968|T201|OSN|751-8|LNC|neutrophil|neutrophil
C0362968|T201|LN|751-8|LNC|neutrophil|neutrophil
C0362968|T201|MTH_LN|751-8|LNC|neutrophil|neutrophil
C0362968|T201|LC|751-8|LNC|neutrophil|neutrophil
C0362969|T201|LN|753-4|LNC|neutrophil counts|neutrophil counts
C0362969|T201|OSN|753-4|LNC|neutrophil counts|neutrophil counts
C0362969|T201|MTH_LN|753-4|LNC|neutrophil counts|neutrophil counts
C0362969|T201|LC|753-4|LNC|neutrophil counts|neutrophil counts
C0362969|T201|LN|753-4|LNC|neutrophil count|neutrophil count
C0362969|T201|OSN|753-4|LNC|neutrophil count|neutrophil count
C0362969|T201|MTH_LN|753-4|LNC|neutrophil count|neutrophil count
C0362969|T201|LC|753-4|LNC|neutrophil count|neutrophil count
C0362969|T201|LN|753-4|LNC|neutrophil|neutrophil
C0362969|T201|OSN|753-4|LNC|neutrophil|neutrophil
C0362969|T201|MTH_LN|753-4|LNC|neutrophil|neutrophil
C0362969|T201|LC|753-4|LNC|neutrophil|neutrophil
C0362987|T201|LN|770-8|LNC|neutrophil counts|neutrophil counts
C0362987|T201|MTH_LN|770-8|LNC|neutrophil counts|neutrophil counts
C0362987|T201|OSN|770-8|LNC|neutrophil counts|neutrophil counts
C0362987|T201|LC|770-8|LNC|neutrophil counts|neutrophil counts
C0362987|T201|LN|770-8|LNC|neutrophil count|neutrophil count
C0362987|T201|MTH_LN|770-8|LNC|neutrophil count|neutrophil count
C0362987|T201|OSN|770-8|LNC|neutrophil count|neutrophil count
C0362987|T201|LC|770-8|LNC|neutrophil count|neutrophil count
C0362987|T201|LN|770-8|LNC|neutrophil|neutrophil
C0362987|T201|MTH_LN|770-8|LNC|neutrophil|neutrophil
C0362987|T201|OSN|770-8|LNC|neutrophil|neutrophil
C0362987|T201|LC|770-8|LNC|neutrophil|neutrophil
C0362994|T201|OSN|777-3|LNC|platelet count|platelet count
C0362994|T201|LN|777-3|LNC|platelet count|platelet count
C0362994|T201|MTH_LN|777-3|LNC|platelet count|platelet count
C0362994|T201|LC|777-3|LNC|platelet count|platelet count
C0363494|T201|LN|1358-1|LNC|adrenocorticotropin|adrenocorticotropin
C0363494|T201|OSN|1358-1|LNC|adrenocorticotropin|adrenocorticotropin
C0363494|T201|MTH_LN|1358-1|LNC|adrenocorticotropin|adrenocorticotropin
C0363494|T201|LC|1358-1|LNC|adrenocorticotropin|adrenocorticotropin
C0363494|T201|LN|1358-1|LNC|ACTH|ACTH
C0363494|T201|OSN|1358-1|LNC|ACTH|ACTH
C0363494|T201|MTH_LN|1358-1|LNC|ACTH|ACTH
C0363494|T201|LC|1358-1|LNC|ACTH|ACTH
C0363496|T201|LN|1360-7|LNC|adrenocorticotropin|adrenocorticotropin
C0363496|T201|MTH_LN|1360-7|LNC|adrenocorticotropin|adrenocorticotropin
C0363496|T201|OSN|1360-7|LNC|adrenocorticotropin|adrenocorticotropin
C0363496|T201|LC|1360-7|LNC|adrenocorticotropin|adrenocorticotropin
C0363496|T201|LN|1360-7|LNC|ACTH|ACTH
C0363496|T201|MTH_LN|1360-7|LNC|ACTH|ACTH
C0363496|T201|OSN|1360-7|LNC|ACTH|ACTH
C0363496|T201|LC|1360-7|LNC|ACTH|ACTH
C0363499|T201|LN|1363-1|LNC|adrenocorticotropin|adrenocorticotropin
C0363499|T201|MTH_LN|1363-1|LNC|adrenocorticotropin|adrenocorticotropin
C0363499|T201|OSN|1363-1|LNC|adrenocorticotropin|adrenocorticotropin
C0363499|T201|LC|1363-1|LNC|adrenocorticotropin|adrenocorticotropin
C0363499|T201|LN|1363-1|LNC|ACTH|ACTH
C0363499|T201|MTH_LN|1363-1|LNC|ACTH|ACTH
C0363499|T201|OSN|1363-1|LNC|ACTH|ACTH
C0363499|T201|LC|1363-1|LNC|ACTH|ACTH
C0363501|T201|LN|1365-6|LNC|adrenocorticotropin|adrenocorticotropin
C0363501|T201|MTH_LN|1365-6|LNC|adrenocorticotropin|adrenocorticotropin
C0363501|T201|OSN|1365-6|LNC|adrenocorticotropin|adrenocorticotropin
C0363501|T201|LC|1365-6|LNC|adrenocorticotropin|adrenocorticotropin
C0363501|T201|LN|1365-6|LNC|ACTH|ACTH
C0363501|T201|MTH_LN|1365-6|LNC|ACTH|ACTH
C0363501|T201|OSN|1365-6|LNC|ACTH|ACTH
C0363501|T201|LC|1365-6|LNC|ACTH|ACTH
C0363617|T201|LN|1483-7|LNC|galactose|galactose
C0363617|T201|MTH_LN|1483-7|LNC|galactose|galactose
C0363617|T201|OSN|1483-7|LNC|galactose|galactose
C0363617|T201|LC|1483-7|LNC|galactose|galactose
C0363625|T201|LN|1491-0|LNC|glucose|glucose
C0363625|T201|MTH_LN|1491-0|LNC|glucose|glucose
C0363625|T201|OSN|1491-0|LNC|glucose|glucose
C0363625|T201|LC|1491-0|LNC|glucose|glucose
C0363626|T201|LN|1492-8|LNC|glucose|glucose
C0363626|T201|OSN|1492-8|LNC|glucose|glucose
C0363626|T201|MTH_LN|1492-8|LNC|glucose|glucose
C0363626|T201|LC|1492-8|LNC|glucose|glucose
C0363627|T201|LN|1493-6|LNC|glucose|glucose
C0363627|T201|OSN|1493-6|LNC|glucose|glucose
C0363627|T201|MTH_LN|1493-6|LNC|glucose|glucose
C0363627|T201|LC|1493-6|LNC|glucose|glucose
C0363628|T201|LN|1494-4|LNC|glucose|glucose
C0363628|T201|OSN|1494-4|LNC|glucose|glucose
C0363628|T201|MTH_LN|1494-4|LNC|glucose|glucose
C0363628|T201|LC|1494-4|LNC|glucose|glucose
C0363629|T201|LN|1495-1|LNC|glucose|glucose
C0363629|T201|OSN|1495-1|LNC|glucose|glucose
C0363629|T201|MTH_LN|1495-1|LNC|glucose|glucose
C0363629|T201|LC|1495-1|LNC|glucose|glucose
C0363631|T201|LN|1497-7|LNC|glucose|glucose
C0363631|T201|OSN|1497-7|LNC|glucose|glucose
C0363631|T201|MTH_LN|1497-7|LNC|glucose|glucose
C0363631|T201|LC|1497-7|LNC|glucose|glucose
C0363632|T201|LN|1498-5|LNC|glucose|glucose
C0363632|T201|MTH_LN|1498-5|LNC|glucose|glucose
C0363632|T201|OSN|1498-5|LNC|glucose|glucose
C0363632|T201|LC|1498-5|LNC|glucose|glucose
C0363633|T201|LN|1499-3|LNC|glucose|glucose
C0363633|T201|MTH_LN|1499-3|LNC|glucose|glucose
C0363633|T201|OSN|1499-3|LNC|glucose|glucose
C0363633|T201|LC|1499-3|LNC|glucose|glucose
C0363634|T201|LN|1500-8|LNC|glucose|glucose
C0363634|T201|MTH_LN|1500-8|LNC|glucose|glucose
C0363634|T201|OSN|1500-8|LNC|glucose|glucose
C0363634|T201|LC|1500-8|LNC|glucose|glucose
C0363635|T201|LN|1501-6|LNC|glucose|glucose
C0363635|T201|MTH_LN|1501-6|LNC|glucose|glucose
C0363635|T201|OSN|1501-6|LNC|glucose|glucose
C0363635|T201|LC|1501-6|LNC|glucose|glucose
C0363637|T201|LN|1503-2|LNC|glucose|glucose
C0363637|T201|MTH_LN|1503-2|LNC|glucose|glucose
C0363637|T201|OSN|1503-2|LNC|glucose|glucose
C0363637|T201|LC|1503-2|LNC|glucose|glucose
C0363638|T201|LN|1504-0|LNC|glucose|glucose
C0363638|T201|MTH_LN|1504-0|LNC|glucose|glucose
C0363638|T201|OSN|1504-0|LNC|glucose|glucose
C0363638|T201|LC|1504-0|LNC|glucose|glucose
C0363639|T201|LN|1505-7|LNC|glucose|glucose
C0363639|T201|MTH_LN|1505-7|LNC|glucose|glucose
C0363639|T201|OSN|1505-7|LNC|glucose|glucose
C0363639|T201|LC|1505-7|LNC|glucose|glucose
C0363640|T201|LN|1506-5|LNC|glucose|glucose
C0363640|T201|MTH_LN|1506-5|LNC|glucose|glucose
C0363640|T201|OSN|1506-5|LNC|glucose|glucose
C0363640|T201|LC|1506-5|LNC|glucose|glucose
C0363641|T201|LN|1507-3|LNC|glucose|glucose
C0363641|T201|MTH_LN|1507-3|LNC|glucose|glucose
C0363641|T201|OSN|1507-3|LNC|glucose|glucose
C0363641|T201|LC|1507-3|LNC|glucose|glucose
C0363643|T201|LN|1509-9|LNC|glucose|glucose
C0363643|T201|MTH_LN|1509-9|LNC|glucose|glucose
C0363643|T201|OSN|1509-9|LNC|glucose|glucose
C0363643|T201|LC|1509-9|LNC|glucose|glucose
C0363644|T201|MTH_LN|1510-7|LNC|glucose|glucose
C0363644|T201|LN|1510-7|LNC|glucose|glucose
C0363644|T201|OSN|1510-7|LNC|glucose|glucose
C0363644|T201|LC|1510-7|LNC|glucose|glucose
C0363645|T201|LN|1512-3|LNC|glucose|glucose
C0363645|T201|MTH_LN|1512-3|LNC|glucose|glucose
C0363645|T201|OSN|1512-3|LNC|glucose|glucose
C0363645|T201|LC|1512-3|LNC|glucose|glucose
C0363646|T201|LN|1513-1|LNC|glucose|glucose
C0363646|T201|MTH_LN|1513-1|LNC|glucose|glucose
C0363646|T201|OSN|1513-1|LNC|glucose|glucose
C0363646|T201|LC|1513-1|LNC|glucose|glucose
C0363647|T201|LN|1514-9|LNC|glucose|glucose
C0363647|T201|MTH_LN|1514-9|LNC|glucose|glucose
C0363647|T201|OSN|1514-9|LNC|glucose|glucose
C0363647|T201|LC|1514-9|LNC|glucose|glucose
C0363649|T201|LN|1516-4|LNC|glucose|glucose
C0363649|T201|MTH_LN|1516-4|LNC|glucose|glucose
C0363649|T201|OSN|1516-4|LNC|glucose|glucose
C0363649|T201|LC|1516-4|LNC|glucose|glucose
C0363650|T201|LN|1517-2|LNC|glucose|glucose
C0363650|T201|MTH_LN|1517-2|LNC|glucose|glucose
C0363650|T201|OSN|1517-2|LNC|glucose|glucose
C0363650|T201|LC|1517-2|LNC|glucose|glucose
C0363651|T201|LN|1518-0|LNC|glucose|glucose
C0363651|T201|MTH_LN|1518-0|LNC|glucose|glucose
C0363651|T201|OSN|1518-0|LNC|glucose|glucose
C0363651|T201|LC|1518-0|LNC|glucose|glucose
C0363653|T201|LN|1520-6|LNC|glucose|glucose
C0363653|T201|MTH_LN|1520-6|LNC|glucose|glucose
C0363653|T201|OSN|1520-6|LNC|glucose|glucose
C0363653|T201|LC|1520-6|LNC|glucose|glucose
C0363655|T201|LN|1522-2|LNC|glucose|glucose
C0363655|T201|MTH_LN|1522-2|LNC|glucose|glucose
C0363655|T201|OSN|1522-2|LNC|glucose|glucose
C0363655|T201|LC|1522-2|LNC|glucose|glucose
C0363656|T201|LN|1523-0|LNC|glucose|glucose
C0363656|T201|MTH_LN|1523-0|LNC|glucose|glucose
C0363656|T201|OSN|1523-0|LNC|glucose|glucose
C0363656|T201|LC|1523-0|LNC|glucose|glucose
C0363658|T201|LN|1525-5|LNC|glucose|glucose
C0363658|T201|MTH_LN|1525-5|LNC|glucose|glucose
C0363658|T201|OSN|1525-5|LNC|glucose|glucose
C0363658|T201|LC|1525-5|LNC|glucose|glucose
C0363659|T201|LN|1526-3|LNC|glucose|glucose
C0363659|T201|MTH_LN|1526-3|LNC|glucose|glucose
C0363659|T201|OSN|1526-3|LNC|glucose|glucose
C0363659|T201|LC|1526-3|LNC|glucose|glucose
C0363661|T201|MTH_LN|1528-9|LNC|glucose|glucose
C0363661|T201|LN|1528-9|LNC|glucose|glucose
C0363661|T201|OSN|1528-9|LNC|glucose|glucose
C0363661|T201|LC|1528-9|LNC|glucose|glucose
C0363662|T201|LN|1530-5|LNC|glucose|glucose
C0363662|T201|MTH_LN|1530-5|LNC|glucose|glucose
C0363662|T201|OSN|1530-5|LNC|glucose|glucose
C0363662|T201|LC|1530-5|LNC|glucose|glucose
C0363665|T201|LN|1533-9|LNC|glucose|glucose
C0363665|T201|MTH_LN|1533-9|LNC|glucose|glucose
C0363665|T201|OSN|1533-9|LNC|glucose|glucose
C0363665|T201|LC|1533-9|LNC|glucose|glucose
C0363666|T201|LN|1534-7|LNC|glucose|glucose
C0363666|T201|MTH_LN|1534-7|LNC|glucose|glucose
C0363666|T201|OSN|1534-7|LNC|glucose|glucose
C0363666|T201|LC|1534-7|LNC|glucose|glucose
C0363667|T201|LN|1535-4|LNC|glucose|glucose
C0363667|T201|MTH_LN|1535-4|LNC|glucose|glucose
C0363667|T201|OSN|1535-4|LNC|glucose|glucose
C0363667|T201|LC|1535-4|LNC|glucose|glucose
C0363668|T201|LN|1536-2|LNC|glucose|glucose
C0363668|T201|MTH_LN|1536-2|LNC|glucose|glucose
C0363668|T201|OSN|1536-2|LNC|glucose|glucose
C0363668|T201|LC|1536-2|LNC|glucose|glucose
C0363669|T201|LN|1537-0|LNC|glucose|glucose
C0363669|T201|MTH_LN|1537-0|LNC|glucose|glucose
C0363669|T201|OSN|1537-0|LNC|glucose|glucose
C0363669|T201|LC|1537-0|LNC|glucose|glucose
C0363671|T201|LN|1539-6|LNC|glucose|glucose
C0363671|T201|MTH_LN|1539-6|LNC|glucose|glucose
C0363671|T201|OSN|1539-6|LNC|glucose|glucose
C0363671|T201|LC|1539-6|LNC|glucose|glucose
C0363672|T201|LN|1540-4|LNC|glucose|glucose
C0363672|T201|MTH_LN|1540-4|LNC|glucose|glucose
C0363672|T201|OSN|1540-4|LNC|glucose|glucose
C0363672|T201|LC|1540-4|LNC|glucose|glucose
C0363674|T201|LN|1542-0|LNC|glucose|glucose
C0363674|T201|MTH_LN|1542-0|LNC|glucose|glucose
C0363674|T201|OSN|1542-0|LNC|glucose|glucose
C0363674|T201|LC|1542-0|LNC|glucose|glucose
C0363675|T201|LN|1543-8|LNC|glucose|glucose
C0363675|T201|MTH_LN|1543-8|LNC|glucose|glucose
C0363675|T201|OSN|1543-8|LNC|glucose|glucose
C0363675|T201|LC|1543-8|LNC|glucose|glucose
C0363678|T201|LN|1547-9|LNC|glucose|glucose
C0363678|T201|MTH_LN|1547-9|LNC|glucose|glucose
C0363678|T201|OSN|1547-9|LNC|glucose|glucose
C0363678|T201|LC|1547-9|LNC|glucose|glucose
C0363685|T201|LN|1554-5|LNC|glucose|glucose
C0363685|T201|MTH_LN|1554-5|LNC|glucose|glucose
C0363685|T201|OSN|1554-5|LNC|glucose|glucose
C0363685|T201|LC|1554-5|LNC|glucose|glucose
C0363686|T201|LN|1555-2|LNC|glucose|glucose
C0363686|T201|MTH_LN|1555-2|LNC|glucose|glucose
C0363686|T201|OSN|1555-2|LNC|glucose|glucose
C0363686|T201|LC|1555-2|LNC|glucose|glucose
C0363688|T201|LN|1557-8|LNC|glucose|glucose
C0363688|T201|MTH_LN|1557-8|LNC|glucose|glucose
C0363688|T201|OSN|1557-8|LNC|glucose|glucose
C0363688|T201|LC|1557-8|LNC|glucose|glucose
C0363688|T201|LN|1557-8|LNC|sugar when fasting|sugar when fasting
C0363688|T201|MTH_LN|1557-8|LNC|sugar when fasting|sugar when fasting
C0363688|T201|OSN|1557-8|LNC|sugar when fasting|sugar when fasting
C0363688|T201|LC|1557-8|LNC|sugar when fasting|sugar when fasting
C0363720|T201|LN|1588-3|LNC|luteinizing|luteinizing
C0363720|T201|OSN|1588-3|LNC|luteinizing|luteinizing
C0363720|T201|MTH_LN|1588-3|LNC|luteinizing|luteinizing
C0363720|T201|LC|1588-3|LNC|luteinizing|luteinizing
C0363720|T201|LN|1588-3|LNC|LH|LH
C0363720|T201|OSN|1588-3|LNC|LH|LH
C0363720|T201|MTH_LN|1588-3|LNC|LH|LH
C0363720|T201|LC|1588-3|LNC|LH|LH
C0363720|T201|LN|1588-3|LNC|luteinising|luteinising
C0363720|T201|OSN|1588-3|LNC|luteinising|luteinising
C0363720|T201|MTH_LN|1588-3|LNC|luteinising|luteinising
C0363720|T201|LC|1588-3|LNC|luteinising|luteinising
C0363724|T201|LN|1592-5|LNC|luteinizing|luteinizing
C0363724|T201|MTH_LN|1592-5|LNC|luteinizing|luteinizing
C0363724|T201|OSN|1592-5|LNC|luteinizing|luteinizing
C0363724|T201|LC|1592-5|LNC|luteinizing|luteinizing
C0363724|T201|LN|1592-5|LNC|LH|LH
C0363724|T201|MTH_LN|1592-5|LNC|LH|LH
C0363724|T201|OSN|1592-5|LNC|LH|LH
C0363724|T201|LC|1592-5|LNC|LH|LH
C0363724|T201|LN|1592-5|LNC|luteinising|luteinising
C0363724|T201|MTH_LN|1592-5|LNC|luteinising|luteinising
C0363724|T201|OSN|1592-5|LNC|luteinising|luteinising
C0363724|T201|LC|1592-5|LNC|luteinising|luteinising
C0363726|T201|LN|1594-1|LNC|luteinizing|luteinizing
C0363726|T201|MTH_LN|1594-1|LNC|luteinizing|luteinizing
C0363726|T201|OSN|1594-1|LNC|luteinizing|luteinizing
C0363726|T201|LC|1594-1|LNC|luteinizing|luteinizing
C0363726|T201|LN|1594-1|LNC|LH|LH
C0363726|T201|MTH_LN|1594-1|LNC|LH|LH
C0363726|T201|OSN|1594-1|LNC|LH|LH
C0363726|T201|LC|1594-1|LNC|LH|LH
C0363726|T201|LN|1594-1|LNC|luteinising|luteinising
C0363726|T201|MTH_LN|1594-1|LNC|luteinising|luteinising
C0363726|T201|OSN|1594-1|LNC|luteinising|luteinising
C0363726|T201|LC|1594-1|LNC|luteinising|luteinising
C0363728|T201|LN|1596-6|LNC|luteinizing|luteinizing
C0363728|T201|MTH_LN|1596-6|LNC|luteinizing|luteinizing
C0363728|T201|OSN|1596-6|LNC|luteinizing|luteinizing
C0363728|T201|LC|1596-6|LNC|luteinizing|luteinizing
C0363728|T201|LN|1596-6|LNC|LH|LH
C0363728|T201|MTH_LN|1596-6|LNC|LH|LH
C0363728|T201|OSN|1596-6|LNC|LH|LH
C0363728|T201|LC|1596-6|LNC|LH|LH
C0363728|T201|LN|1596-6|LNC|luteinising|luteinising
C0363728|T201|MTH_LN|1596-6|LNC|luteinising|luteinising
C0363728|T201|OSN|1596-6|LNC|luteinising|luteinising
C0363728|T201|LC|1596-6|LNC|luteinising|luteinising
C0363731|T201|LN|1599-0|LNC|luteinizing|luteinizing
C0363731|T201|MTH_LN|1599-0|LNC|luteinizing|luteinizing
C0363731|T201|OSN|1599-0|LNC|luteinizing|luteinizing
C0363731|T201|LC|1599-0|LNC|luteinizing|luteinizing
C0363731|T201|LN|1599-0|LNC|LH|LH
C0363731|T201|MTH_LN|1599-0|LNC|LH|LH
C0363731|T201|OSN|1599-0|LNC|LH|LH
C0363731|T201|LC|1599-0|LNC|LH|LH
C0363731|T201|LN|1599-0|LNC|luteinising|luteinising
C0363731|T201|MTH_LN|1599-0|LNC|luteinising|luteinising
C0363731|T201|OSN|1599-0|LNC|luteinising|luteinising
C0363731|T201|LC|1599-0|LNC|luteinising|luteinising
C0363783|T201|LN|1649-3|LNC|calcium|calcium
C0363783|T201|MTH_LN|1649-3|LNC|calcium|calcium
C0363783|T201|LC|1649-3|LNC|calcium|calcium
C0363783|T201|OSN|1649-3|LNC|calcium|calcium
C0363802|T201|LN|1668-3|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C0363802|T201|MTH_LN|1668-3|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C0363802|T201|OSN|1668-3|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C0363802|T201|LC|1668-3|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C0363802|T201|LN|1668-3|LNC|17-OHP|17-OHP
C0363802|T201|MTH_LN|1668-3|LNC|17-OHP|17-OHP
C0363802|T201|OSN|1668-3|LNC|17-OHP|17-OHP
C0363802|T201|LC|1668-3|LNC|17-OHP|17-OHP
C0363808|T201|LN|1674-1|LNC|corticosterone|corticosterone
C0363808|T201|MTH_LN|1674-1|LNC|corticosterone|corticosterone
C0363808|T201|OSN|1674-1|LNC|corticosterone|corticosterone
C0363808|T201|LC|1674-1|LNC|corticosterone|corticosterone
C0363813|T201|LN|1679-0|LNC|vitamin D metabolism|vitamin D metabolism
C0363813|T201|MTH_LN|1679-0|LNC|vitamin D metabolism|vitamin D metabolism
C0363813|T201|OSN|1679-0|LNC|vitamin D metabolism|vitamin D metabolism
C0363813|T201|LC|1679-0|LNC|vitamin D metabolism|vitamin D metabolism
C0363813|T201|LN|1679-0|LNC|calcifediol|calcifediol
C0363813|T201|MTH_LN|1679-0|LNC|calcifediol|calcifediol
C0363813|T201|OSN|1679-0|LNC|calcifediol|calcifediol
C0363813|T201|LC|1679-0|LNC|calcifediol|calcifediol
C0363813|T201|LN|1679-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C0363813|T201|MTH_LN|1679-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C0363813|T201|OSN|1679-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C0363813|T201|LC|1679-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C0363813|T201|LN|1679-0|LNC|calcidiol|calcidiol
C0363813|T201|MTH_LN|1679-0|LNC|calcidiol|calcidiol
C0363813|T201|OSN|1679-0|LNC|calcidiol|calcidiol
C0363813|T201|LC|1679-0|LNC|calcidiol|calcidiol
C0363813|T201|LN|1679-0|LNC|calcitriol|calcitriol
C0363813|T201|MTH_LN|1679-0|LNC|calcitriol|calcitriol
C0363813|T201|OSN|1679-0|LNC|calcitriol|calcitriol
C0363813|T201|LC|1679-0|LNC|calcitriol|calcitriol
C0363813|T201|LN|1679-0|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C0363813|T201|MTH_LN|1679-0|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C0363813|T201|OSN|1679-0|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C0363813|T201|LC|1679-0|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C0363813|T201|LN|1679-0|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C0363813|T201|MTH_LN|1679-0|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C0363813|T201|OSN|1679-0|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C0363813|T201|LC|1679-0|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C0363822|T201|LN|1688-1|LNC|vitamin b6|vitamin b6
C0363822|T201|MTH_LN|1688-1|LNC|vitamin b6|vitamin b6
C0363822|T201|OSN|1688-1|LNC|vitamin b6|vitamin b6
C0363822|T201|LC|1688-1|LNC|vitamin b6|vitamin b6
C0363822|T201|LN|1688-1|LNC|vitamin B metabolism|vitamin B metabolism
C0363822|T201|MTH_LN|1688-1|LNC|vitamin B metabolism|vitamin B metabolism
C0363822|T201|OSN|1688-1|LNC|vitamin B metabolism|vitamin B metabolism
C0363822|T201|LC|1688-1|LNC|vitamin B metabolism|vitamin B metabolism
C0363822|T201|LN|1688-1|LNC|B-vitamin metabolism|B-vitamin metabolism
C0363822|T201|MTH_LN|1688-1|LNC|B-vitamin metabolism|B-vitamin metabolism
C0363822|T201|OSN|1688-1|LNC|B-vitamin metabolism|B-vitamin metabolism
C0363822|T201|LC|1688-1|LNC|B-vitamin metabolism|B-vitamin metabolism
C0363851|T201|LN|1717-8|LNC|acylcarnitine|acylcarnitine
C0363851|T201|LC|1717-8|LNC|acylcarnitine|acylcarnitine
C0363851|T201|MTH_LN|1717-8|LNC|acylcarnitine|acylcarnitine
C0363851|T201|OSN|1717-8|LNC|acylcarnitine|acylcarnitine
C0363856|T201|LN|1722-8|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C0363856|T201|MTH_LN|1722-8|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C0363856|T201|OSN|1722-8|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C0363856|T201|LC|1722-8|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C0363856|T201|LN|1722-8|LNC|red cell adenosine deaminase activity|red cell adenosine deaminase activity
C0363856|T201|MTH_LN|1722-8|LNC|red cell adenosine deaminase activity|red cell adenosine deaminase activity
C0363856|T201|OSN|1722-8|LNC|red cell adenosine deaminase activity|red cell adenosine deaminase activity
C0363856|T201|LC|1722-8|LNC|red cell adenosine deaminase activity|red cell adenosine deaminase activity
C0363880|T201|LN|1746-7|LNC|CSF albumin|CSF albumin
C0363880|T201|MTH_LN|1746-7|LNC|CSF albumin|CSF albumin
C0363880|T201|OSN|1746-7|LNC|CSF albumin|CSF albumin
C0363880|T201|LC|1746-7|LNC|CSF albumin|CSF albumin
C0363880|T201|LN|1746-7|LNC|CSF albumin is belowlower limitnormal.|CSF albumin is belowlower limitnormal.
C0363880|T201|MTH_LN|1746-7|LNC|CSF albumin is belowlower limitnormal.|CSF albumin is belowlower limitnormal.
C0363880|T201|OSN|1746-7|LNC|CSF albumin is belowlower limitnormal.|CSF albumin is belowlower limitnormal.
C0363880|T201|LC|1746-7|LNC|CSF albumin is belowlower limitnormal.|CSF albumin is belowlower limitnormal.
C0363880|T201|LN|1746-7|LNC|CSF protein|CSF protein
C0363880|T201|MTH_LN|1746-7|LNC|CSF protein|CSF protein
C0363880|T201|OSN|1746-7|LNC|CSF protein|CSF protein
C0363880|T201|LC|1746-7|LNC|CSF protein|CSF protein
C0363885|T201|LN|1751-7|LNC|albumin|albumin
C0363885|T201|MTH_LN|1751-7|LNC|albumin|albumin
C0363885|T201|OSN|1751-7|LNC|albumin|albumin
C0363885|T201|LC|1751-7|LNC|albumin|albumin
C0363893|T201|LN|1759-0|LNC|albumin|albumin
C0363893|T201|OSN|1759-0|LNC|albumin|albumin
C0363893|T201|MTH_LN|1759-0|LNC|albumin|albumin
C0363893|T201|LC|1759-0|LNC|albumin|albumin
C0363895|T201|LN|1761-6|LNC|aldolase|aldolase
C0363895|T201|MTH_LN|1761-6|LNC|aldolase|aldolase
C0363895|T201|OSN|1761-6|LNC|aldolase|aldolase
C0363895|T201|LC|1761-6|LNC|aldolase|aldolase
C0363897|T201|LN|1763-2|LNC|aldosterone|aldosterone
C0363897|T201|MTH_LN|1763-2|LNC|aldosterone|aldosterone
C0363897|T201|OSN|1763-2|LNC|aldosterone|aldosterone
C0363897|T201|LC|1763-2|LNC|aldosterone|aldosterone
C0363911|T201|LN|1777-2|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363911|T201|MTH_LN|1777-2|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363911|T201|OSN|1777-2|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363911|T201|LC|1777-2|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363911|T201|LN|1777-2|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C0363911|T201|MTH_LN|1777-2|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C0363911|T201|OSN|1777-2|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C0363911|T201|LC|1777-2|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C0363911|T201|LN|1777-2|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C0363911|T201|MTH_LN|1777-2|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C0363911|T201|OSN|1777-2|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C0363911|T201|LC|1777-2|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C0363911|T201|LN|1777-2|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0363911|T201|MTH_LN|1777-2|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0363911|T201|OSN|1777-2|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0363911|T201|LC|1777-2|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0363912|T201|LN|1778-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363912|T201|MTH_LN|1778-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363912|T201|OSN|1778-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363912|T201|LC|1778-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0363912|T201|LN|1778-0|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C0363912|T201|MTH_LN|1778-0|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C0363912|T201|OSN|1778-0|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C0363912|T201|LC|1778-0|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C0363912|T201|LN|1778-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0363912|T201|MTH_LN|1778-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0363912|T201|OSN|1778-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0363912|T201|LC|1778-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0363968|T201|LN|1834-1|LNC|alpha-fetoprotein|alpha-fetoprotein
C0363968|T201|OSN|1834-1|LNC|alpha-fetoprotein|alpha-fetoprotein
C0363968|T201|MTH_LN|1834-1|LNC|alpha-fetoprotein|alpha-fetoprotein
C0363968|T201|LC|1834-1|LNC|alpha-fetoprotein|alpha-fetoprotein
C0363968|T201|LN|1834-1|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0363968|T201|OSN|1834-1|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0363968|T201|MTH_LN|1834-1|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0363968|T201|LC|1834-1|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0363968|T201|LN|1834-1|LNC|alpha fetoprotein|alpha fetoprotein
C0363968|T201|OSN|1834-1|LNC|alpha fetoprotein|alpha fetoprotein
C0363968|T201|MTH_LN|1834-1|LNC|alpha fetoprotein|alpha fetoprotein
C0363968|T201|LC|1834-1|LNC|alpha fetoprotein|alpha fetoprotein
C0363971|T201|LN|1836-6|LNC|retinol-binding protein|retinol-binding protein
C0363971|T201|MTH_LN|1836-6|LNC|retinol-binding protein|retinol-binding protein
C0363971|T201|OSN|1836-6|LNC|retinol-binding protein|retinol-binding protein
C0363971|T201|LC|1836-6|LNC|retinol-binding protein|retinol-binding protein
C0363974|T201|LN|1839-0|LNC|ammonia|ammonia
C0363974|T201|MTH_LN|1839-0|LNC|ammonia|ammonia
C0363974|T201|OSN|1839-0|LNC|ammonia|ammonia
C0363974|T201|LC|1839-0|LNC|ammonia|ammonia
C0363976|T201|LN|1841-6|LNC|ammonia|ammonia
C0363976|T201|MTH_LN|1841-6|LNC|ammonia|ammonia
C0363976|T201|OSN|1841-6|LNC|ammonia|ammonia
C0363976|T201|LC|1841-6|LNC|ammonia|ammonia
C0363983|T201|LN|1848-1|LNC|testosterone|testosterone
C0363983|T201|MTH_LN|1848-1|LNC|testosterone|testosterone
C0363983|T201|OSN|1848-1|LNC|testosterone|testosterone
C0363983|T201|LC|1848-1|LNC|testosterone|testosterone
C0363983|T201|LN|1848-1|LNC|androgen|androgen
C0363983|T201|MTH_LN|1848-1|LNC|androgen|androgen
C0363983|T201|OSN|1848-1|LNC|androgen|androgen
C0363983|T201|LC|1848-1|LNC|androgen|androgen
C0363989|T201|LN|1854-9|LNC|androstenedione|androstenedione
C0363989|T201|MTH_LN|1854-9|LNC|androstenedione|androstenedione
C0363989|T201|OSN|1854-9|LNC|androstenedione|androstenedione
C0363989|T201|LC|1854-9|LNC|androstenedione|androstenedione
C0363989|T201|LN|1854-9|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C0363989|T201|MTH_LN|1854-9|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C0363989|T201|OSN|1854-9|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C0363989|T201|LC|1854-9|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C0363989|T201|LN|1854-9|LNC|androstenolone|androstenolone
C0363989|T201|MTH_LN|1854-9|LNC|androstenolone|androstenolone
C0363989|T201|OSN|1854-9|LNC|androstenolone|androstenolone
C0363989|T201|LC|1854-9|LNC|androstenolone|androstenolone
C0363989|T201|LN|1854-9|LNC|DHEA|DHEA
C0363989|T201|MTH_LN|1854-9|LNC|DHEA|DHEA
C0363989|T201|OSN|1854-9|LNC|DHEA|DHEA
C0363989|T201|LC|1854-9|LNC|DHEA|DHEA
C0364019|T201|MTH_LN|1884-6|LNC|apolipoprotein|apolipoprotein
C0364019|T201|LN|1884-6|LNC|apolipoprotein|apolipoprotein
C0364019|T201|OSN|1884-6|LNC|apolipoprotein|apolipoprotein
C0364019|T201|LC|1884-6|LNC|apolipoprotein|apolipoprotein
C0364019|T201|MTH_LN|1884-6|LNC|apolipoprotein B|apolipoprotein B
C0364019|T201|LN|1884-6|LNC|apolipoprotein B|apolipoprotein B
C0364019|T201|OSN|1884-6|LNC|apolipoprotein B|apolipoprotein B
C0364019|T201|LC|1884-6|LNC|apolipoprotein B|apolipoprotein B
C0364019|T201|MTH_LN|1884-6|LNC|ApoB|ApoB
C0364019|T201|LN|1884-6|LNC|ApoB|ApoB
C0364019|T201|OSN|1884-6|LNC|ApoB|ApoB
C0364019|T201|LC|1884-6|LNC|ApoB|ApoB
C0364028|T201|LN|1893-7|LNC|arginine metabolism|arginine metabolism
C0364028|T201|MTH_LN|1893-7|LNC|arginine metabolism|arginine metabolism
C0364028|T201|OSN|1893-7|LNC|arginine metabolism|arginine metabolism
C0364028|T201|LC|1893-7|LNC|arginine metabolism|arginine metabolism
C0364028|T201|LN|1893-7|LNC|arginine|arginine
C0364028|T201|MTH_LN|1893-7|LNC|arginine|arginine
C0364028|T201|OSN|1893-7|LNC|arginine|arginine
C0364028|T201|LC|1893-7|LNC|arginine|arginine
C0364029|T201|LN|1894-5|LNC|arginine|arginine
C0364029|T201|MTH_LN|1894-5|LNC|arginine|arginine
C0364029|T201|OSN|1894-5|LNC|arginine|arginine
C0364029|T201|LC|1894-5|LNC|arginine|arginine
C0364030|T201|LN|1895-2|LNC|arginine|arginine
C0364030|T201|MTH_LN|1895-2|LNC|arginine|arginine
C0364030|T201|OSN|1895-2|LNC|arginine|arginine
C0364030|T201|LC|1895-2|LNC|arginine|arginine
C0364085|T201|LN|1952-1|LNC|beta-2-microglobulin|beta-2-microglobulin
C0364085|T201|OSN|1952-1|LNC|beta-2-microglobulin|beta-2-microglobulin
C0364085|T201|LC|1952-1|LNC|beta-2-microglobulin|beta-2-microglobulin
C0364085|T201|MTH_LN|1952-1|LNC|beta-2-microglobulin|beta-2-microglobulin
C0364085|T201|LN|1952-1|LNC|B2M|B2M
C0364085|T201|OSN|1952-1|LNC|B2M|B2M
C0364085|T201|LC|1952-1|LNC|B2M|B2M
C0364085|T201|MTH_LN|1952-1|LNC|B2M|B2M
C0364085|T201|LN|1952-1|LNC|beta2m|beta2m
C0364085|T201|OSN|1952-1|LNC|beta2m|beta2m
C0364085|T201|LC|1952-1|LNC|beta2m|beta2m
C0364085|T201|MTH_LN|1952-1|LNC|beta2m|beta2m
C0364085|T201|LN|1952-1|LNC|beta2 microglobulin|beta2 microglobulin
C0364085|T201|OSN|1952-1|LNC|beta2 microglobulin|beta2 microglobulin
C0364085|T201|LC|1952-1|LNC|beta2 microglobulin|beta2 microglobulin
C0364085|T201|MTH_LN|1952-1|LNC|beta2 microglobulin|beta2 microglobulin
C0364085|T201|LN|1952-1|LNC|beta2-m|beta2-m
C0364085|T201|OSN|1952-1|LNC|beta2-m|beta2-m
C0364085|T201|LC|1952-1|LNC|beta2-m|beta2-m
C0364085|T201|MTH_LN|1952-1|LNC|beta2-m|beta2-m
C0364097|T201|LN|1964-6|LNC|bicarbonate|bicarbonate
C0364097|T201|MTH_LN|1964-6|LNC|bicarbonate|bicarbonate
C0364097|T201|OSN|1964-6|LNC|bicarbonate|bicarbonate
C0364097|T201|LC|1964-6|LNC|bicarbonate|bicarbonate
C0364101|T201|LN|1968-7|LNC|bilirubin|bilirubin
C0364101|T201|MTH_LN|1968-7|LNC|bilirubin|bilirubin
C0364101|T201|OSN|1968-7|LNC|bilirubin|bilirubin
C0364101|T201|LC|1968-7|LNC|bilirubin|bilirubin
C0364101|T201|LN|1968-7|LNC|metabolism/homeostasis|metabolism/homeostasis
C0364101|T201|MTH_LN|1968-7|LNC|metabolism/homeostasis|metabolism/homeostasis
C0364101|T201|OSN|1968-7|LNC|metabolism/homeostasis|metabolism/homeostasis
C0364101|T201|LC|1968-7|LNC|metabolism/homeostasis|metabolism/homeostasis
C0364101|T201|LN|1968-7|LNC|Metabolism|Metabolism
C0364101|T201|MTH_LN|1968-7|LNC|Metabolism|Metabolism
C0364101|T201|OSN|1968-7|LNC|Metabolism|Metabolism
C0364101|T201|LC|1968-7|LNC|Metabolism|Metabolism
C0364101|T201|LN|1968-7|LNC|Laboratory|Laboratory
C0364101|T201|MTH_LN|1968-7|LNC|Laboratory|Laboratory
C0364101|T201|OSN|1968-7|LNC|Laboratory|Laboratory
C0364101|T201|LC|1968-7|LNC|Laboratory|Laboratory
C0364104|T201|LN|1971-1|LNC|bilirubin|bilirubin
C0364104|T201|MTH_LN|1971-1|LNC|bilirubin|bilirubin
C0364104|T201|OSN|1971-1|LNC|bilirubin|bilirubin
C0364104|T201|LC|1971-1|LNC|bilirubin|bilirubin
C0364108|T201|LN|1975-2|LNC|bilirubin|bilirubin
C0364108|T201|MTH_LN|1975-2|LNC|bilirubin|bilirubin
C0364108|T201|OSN|1975-2|LNC|bilirubin|bilirubin
C0364108|T201|LC|1975-2|LNC|bilirubin|bilirubin
C0364108|T201|LN|1975-2|LNC|total bilirubin|total bilirubin
C0364108|T201|MTH_LN|1975-2|LNC|total bilirubin|total bilirubin
C0364108|T201|OSN|1975-2|LNC|total bilirubin|total bilirubin
C0364108|T201|LC|1975-2|LNC|total bilirubin|total bilirubin
C0364108|T201|LN|1975-2|LNC|bili total|bili total
C0364108|T201|MTH_LN|1975-2|LNC|bili total|bili total
C0364108|T201|OSN|1975-2|LNC|bili total|bili total
C0364108|T201|LC|1975-2|LNC|bili total|bili total
C0364119|T201|MTH_LN|1986-9|LNC|C-peptide|C-peptide
C0364119|T201|LN|1986-9|LNC|C-peptide|C-peptide
C0364119|T201|OSN|1986-9|LNC|C-peptide|C-peptide
C0364119|T201|LC|1986-9|LNC|C-peptide|C-peptide
C0364119|T201|MTH_LN|1986-9|LNC|C peptide|C peptide
C0364119|T201|LN|1986-9|LNC|C peptide|C peptide
C0364119|T201|OSN|1986-9|LNC|C peptide|C peptide
C0364119|T201|LC|1986-9|LNC|C peptide|C peptide
C0364121|T201|LN|1988-5|LNC|CRP|CRP
C0364121|T201|MTH_LN|1988-5|LNC|CRP|CRP
C0364121|T201|OSN|1988-5|LNC|CRP|CRP
C0364121|T201|LC|1988-5|LNC|CRP|CRP
C0364121|T201|LN|1988-5|LNC|C-reactive protein|C-reactive protein
C0364121|T201|MTH_LN|1988-5|LNC|C-reactive protein|C-reactive protein
C0364121|T201|OSN|1988-5|LNC|C-reactive protein|C-reactive protein
C0364121|T201|LC|1988-5|LNC|C-reactive protein|C-reactive protein
C0364121|T201|LN|1988-5|LNC|C-peptide|C-peptide
C0364121|T201|MTH_LN|1988-5|LNC|C-peptide|C-peptide
C0364121|T201|OSN|1988-5|LNC|C-peptide|C-peptide
C0364121|T201|LC|1988-5|LNC|C-peptide|C-peptide
C0364121|T201|LN|1988-5|LNC|C peptide|C peptide
C0364121|T201|MTH_LN|1988-5|LNC|C peptide|C peptide
C0364121|T201|OSN|1988-5|LNC|C peptide|C peptide
C0364121|T201|LC|1988-5|LNC|C peptide|C peptide
C0364122|T201|LN|1989-3|LNC|vitamin D metabolism|vitamin D metabolism
C0364122|T201|MTH_LN|1989-3|LNC|vitamin D metabolism|vitamin D metabolism
C0364122|T201|LC|1989-3|LNC|vitamin D metabolism|vitamin D metabolism
C0364122|T201|OSN|1989-3|LNC|vitamin D metabolism|vitamin D metabolism
C0364122|T201|LN|1989-3|LNC|calcifediol|calcifediol
C0364122|T201|MTH_LN|1989-3|LNC|calcifediol|calcifediol
C0364122|T201|LC|1989-3|LNC|calcifediol|calcifediol
C0364122|T201|OSN|1989-3|LNC|calcifediol|calcifediol
C0364122|T201|LN|1989-3|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C0364122|T201|MTH_LN|1989-3|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C0364122|T201|LC|1989-3|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C0364122|T201|OSN|1989-3|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C0364122|T201|LN|1989-3|LNC|calcidiol|calcidiol
C0364122|T201|MTH_LN|1989-3|LNC|calcidiol|calcidiol
C0364122|T201|LC|1989-3|LNC|calcidiol|calcidiol
C0364122|T201|OSN|1989-3|LNC|calcidiol|calcidiol
C0364122|T201|LN|1989-3|LNC|calcitriol|calcitriol
C0364122|T201|MTH_LN|1989-3|LNC|calcitriol|calcitriol
C0364122|T201|LC|1989-3|LNC|calcitriol|calcitriol
C0364122|T201|OSN|1989-3|LNC|calcitriol|calcitriol
C0364122|T201|LN|1989-3|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C0364122|T201|MTH_LN|1989-3|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C0364122|T201|LC|1989-3|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C0364122|T201|OSN|1989-3|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C0364122|T201|LN|1989-3|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C0364122|T201|MTH_LN|1989-3|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C0364122|T201|LC|1989-3|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C0364122|T201|OSN|1989-3|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C0364127|T201|LN|1994-3|LNC|calcium|calcium
C0364127|T201|MTH_LN|1994-3|LNC|calcium|calcium
C0364127|T201|OSN|1994-3|LNC|calcium|calcium
C0364127|T201|LC|1994-3|LNC|calcium|calcium
C0364127|T201|LN|1994-3|LNC|calcium homeostasis|calcium homeostasis
C0364127|T201|MTH_LN|1994-3|LNC|calcium homeostasis|calcium homeostasis
C0364127|T201|OSN|1994-3|LNC|calcium homeostasis|calcium homeostasis
C0364127|T201|LC|1994-3|LNC|calcium homeostasis|calcium homeostasis
C0364128|T201|LN|1995-0|LNC|calcium|calcium
C0364128|T201|MTH_LN|1995-0|LNC|calcium|calcium
C0364128|T201|OSN|1995-0|LNC|calcium|calcium
C0364128|T201|LC|1995-0|LNC|calcium|calcium
C0364128|T201|LN|1995-0|LNC|calcium homeostasis|calcium homeostasis
C0364128|T201|MTH_LN|1995-0|LNC|calcium homeostasis|calcium homeostasis
C0364128|T201|OSN|1995-0|LNC|calcium homeostasis|calcium homeostasis
C0364128|T201|LC|1995-0|LNC|calcium homeostasis|calcium homeostasis
C0364129|T201|LN|1996-8|LNC|calcium|calcium
C0364129|T201|MTH_LN|1996-8|LNC|calcium|calcium
C0364129|T201|OSN|1996-8|LNC|calcium|calcium
C0364129|T201|LC|1996-8|LNC|calcium|calcium
C0364129|T201|LN|1996-8|LNC|calcium homeostasis|calcium homeostasis
C0364129|T201|MTH_LN|1996-8|LNC|calcium homeostasis|calcium homeostasis
C0364129|T201|OSN|1996-8|LNC|calcium homeostasis|calcium homeostasis
C0364129|T201|LC|1996-8|LNC|calcium homeostasis|calcium homeostasis
C0364133|T201|LN|2000-8|LNC|calcium|calcium
C0364133|T201|MTH_LN|2000-8|LNC|calcium|calcium
C0364133|T201|OSN|2000-8|LNC|calcium|calcium
C0364133|T201|LC|2000-8|LNC|calcium|calcium
C0364133|T201|LN|2000-8|LNC|calcium homeostasis|calcium homeostasis
C0364133|T201|MTH_LN|2000-8|LNC|calcium homeostasis|calcium homeostasis
C0364133|T201|OSN|2000-8|LNC|calcium homeostasis|calcium homeostasis
C0364133|T201|LC|2000-8|LNC|calcium homeostasis|calcium homeostasis
C0364151|T201|LN|2019-8|LNC|carbon dioxide|carbon dioxide
C0364151|T201|MTH_LN|2019-8|LNC|carbon dioxide|carbon dioxide
C0364151|T201|LC|2019-8|LNC|carbon dioxide|carbon dioxide
C0364151|T201|OSN|2019-8|LNC|carbon dioxide|carbon dioxide
C0364152|T201|LN|2020-6|LNC|carbon dioxide|carbon dioxide
C0364152|T201|MTH_LN|2020-6|LNC|carbon dioxide|carbon dioxide
C0364152|T201|LC|2020-6|LNC|carbon dioxide|carbon dioxide
C0364152|T201|OSN|2020-6|LNC|carbon dioxide|carbon dioxide
C0364153|T201|LN|2021-4|LNC|carbon dioxide|carbon dioxide
C0364153|T201|MTH_LN|2021-4|LNC|carbon dioxide|carbon dioxide
C0364153|T201|OSN|2021-4|LNC|carbon dioxide|carbon dioxide
C0364153|T201|LC|2021-4|LNC|carbon dioxide|carbon dioxide
C0364159|T201|LN|2027-1|LNC|carbon dioxide|carbon dioxide
C0364159|T201|MTH_LN|2027-1|LNC|carbon dioxide|carbon dioxide
C0364159|T201|OSN|2027-1|LNC|carbon dioxide|carbon dioxide
C0364159|T201|LC|2027-1|LNC|carbon dioxide|carbon dioxide
C0364160|T201|LN|2028-9|LNC|carbon dioxide|carbon dioxide
C0364160|T201|MTH_LN|2028-9|LNC|carbon dioxide|carbon dioxide
C0364160|T201|OSN|2028-9|LNC|carbon dioxide|carbon dioxide
C0364160|T201|LC|2028-9|LNC|carbon dioxide|carbon dioxide
C0364171|T201|LN|2039-6|LNC|carcinoembryonic antigen|carcinoembryonic antigen
C0364171|T201|MTH_LN|2039-6|LNC|carcinoembryonic antigen|carcinoembryonic antigen
C0364171|T201|OSN|2039-6|LNC|carcinoembryonic antigen|carcinoembryonic antigen
C0364171|T201|LC|2039-6|LNC|carcinoembryonic antigen|carcinoembryonic antigen
C0364171|T201|LN|2039-6|LNC|CEA|CEA
C0364171|T201|MTH_LN|2039-6|LNC|CEA|CEA
C0364171|T201|OSN|2039-6|LNC|CEA|CEA
C0364171|T201|LC|2039-6|LNC|CEA|CEA
C0364201|T201|LN|2069-3|LNC|chloride|chloride
C0364201|T201|MTH_LN|2069-3|LNC|chloride|chloride
C0364201|T201|OSN|2069-3|LNC|chloride|chloride
C0364201|T201|LC|2069-3|LNC|chloride|chloride
C0364201|T201|LN|2069-3|LNC|chloride homeostasis|chloride homeostasis
C0364201|T201|MTH_LN|2069-3|LNC|chloride homeostasis|chloride homeostasis
C0364201|T201|OSN|2069-3|LNC|chloride homeostasis|chloride homeostasis
C0364201|T201|LC|2069-3|LNC|chloride homeostasis|chloride homeostasis
C0364207|T201|LN|2075-0|LNC|chloride|chloride
C0364207|T201|MTH_LN|2075-0|LNC|chloride|chloride
C0364207|T201|OSN|2075-0|LNC|chloride|chloride
C0364207|T201|LC|2075-0|LNC|chloride|chloride
C0364207|T201|LN|2075-0|LNC|chloride homeostasis|chloride homeostasis
C0364207|T201|MTH_LN|2075-0|LNC|chloride homeostasis|chloride homeostasis
C0364207|T201|OSN|2075-0|LNC|chloride homeostasis|chloride homeostasis
C0364207|T201|LC|2075-0|LNC|chloride homeostasis|chloride homeostasis
C0364209|T201|LN|2077-6|LNC|sweat chloride|sweat chloride
C0364209|T201|MTH_LN|2077-6|LNC|sweat chloride|sweat chloride
C0364209|T201|OSN|2077-6|LNC|sweat chloride|sweat chloride
C0364209|T201|LC|2077-6|LNC|sweat chloride|sweat chloride
C0364210|T201|LN|2078-4|LNC|chloride|chloride
C0364210|T201|MTH_LN|2078-4|LNC|chloride|chloride
C0364210|T201|OSN|2078-4|LNC|chloride|chloride
C0364210|T201|LC|2078-4|LNC|chloride|chloride
C0364214|T201|LN|2082-6|LNC|cholesterol|cholesterol
C0364214|T201|MTH_LN|2082-6|LNC|cholesterol|cholesterol
C0364214|T201|OSN|2082-6|LNC|cholesterol|cholesterol
C0364214|T201|LC|2082-6|LNC|cholesterol|cholesterol
C0364214|T201|LN|2082-6|LNC|total cholesterol|total cholesterol
C0364214|T201|MTH_LN|2082-6|LNC|total cholesterol|total cholesterol
C0364214|T201|OSN|2082-6|LNC|total cholesterol|total cholesterol
C0364214|T201|LC|2082-6|LNC|total cholesterol|total cholesterol
C0364214|T201|LN|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C0364214|T201|MTH_LN|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C0364214|T201|OSN|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C0364214|T201|LC|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C0364221|T201|LC|2085-9|LNC|HDL cholesterol|HDL cholesterol
C0364221|T201|MTH_LN|2085-9|LNC|HDL cholesterol|HDL cholesterol
C0364221|T201|LN|2085-9|LNC|HDL cholesterol|HDL cholesterol
C0364221|T201|OSN|2085-9|LNC|HDL cholesterol|HDL cholesterol
C0364221|T201|LC|2085-9|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0364221|T201|MTH_LN|2085-9|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0364221|T201|LN|2085-9|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0364221|T201|OSN|2085-9|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0364221|T201|LC|2085-9|LNC|HDL-cholesterol|HDL-cholesterol
C0364221|T201|MTH_LN|2085-9|LNC|HDL-cholesterol|HDL-cholesterol
C0364221|T201|LN|2085-9|LNC|HDL-cholesterol|HDL-cholesterol
C0364221|T201|OSN|2085-9|LNC|HDL-cholesterol|HDL-cholesterol
C0364221|T201|LC|2085-9|LNC|high-density lipoprotein|high-density lipoprotein
C0364221|T201|MTH_LN|2085-9|LNC|high-density lipoprotein|high-density lipoprotein
C0364221|T201|LN|2085-9|LNC|high-density lipoprotein|high-density lipoprotein
C0364221|T201|OSN|2085-9|LNC|high-density lipoprotein|high-density lipoprotein
C0364221|T201|LC|2085-9|LNC|HDL|HDL
C0364221|T201|MTH_LN|2085-9|LNC|HDL|HDL
C0364221|T201|LN|2085-9|LNC|HDL|HDL
C0364221|T201|OSN|2085-9|LNC|HDL|HDL
C0364225|T201|MTH_LN|2089-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0364225|T201|LN|2089-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0364225|T201|OSN|2089-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0364225|T201|LC|2089-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0364225|T201|MTH_LN|2089-1|LNC|LDL|LDL
C0364225|T201|LN|2089-1|LNC|LDL|LDL
C0364225|T201|OSN|2089-1|LNC|LDL|LDL
C0364225|T201|LC|2089-1|LNC|LDL|LDL
C0364225|T201|MTH_LN|2089-1|LNC|LDL cholesterol|LDL cholesterol
C0364225|T201|LN|2089-1|LNC|LDL cholesterol|LDL cholesterol
C0364225|T201|OSN|2089-1|LNC|LDL cholesterol|LDL cholesterol
C0364225|T201|LC|2089-1|LNC|LDL cholesterol|LDL cholesterol
C0364225|T201|MTH_LN|2089-1|LNC|low-density lipoprotein|low-density lipoprotein
C0364225|T201|LN|2089-1|LNC|low-density lipoprotein|low-density lipoprotein
C0364225|T201|OSN|2089-1|LNC|low-density lipoprotein|low-density lipoprotein
C0364225|T201|LC|2089-1|LNC|low-density lipoprotein|low-density lipoprotein
C0364225|T201|MTH_LN|2089-1|LNC|beta-lipoproteins|beta-lipoproteins
C0364225|T201|LN|2089-1|LNC|beta-lipoproteins|beta-lipoproteins
C0364225|T201|OSN|2089-1|LNC|beta-lipoproteins|beta-lipoproteins
C0364225|T201|LC|2089-1|LNC|beta-lipoproteins|beta-lipoproteins
C0364225|T201|MTH_LN|2089-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0364225|T201|LN|2089-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0364225|T201|OSN|2089-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0364225|T201|LC|2089-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0364225|T201|MTH_LN|2089-1|LNC|LDL-C|LDL-C
C0364225|T201|LN|2089-1|LNC|LDL-C|LDL-C
C0364225|T201|OSN|2089-1|LNC|LDL-C|LDL-C
C0364225|T201|LC|2089-1|LNC|LDL-C|LDL-C
C0364227|T201|LC|2091-7|LNC|VLDL cholesterol|VLDL cholesterol
C0364227|T201|MTH_LN|2091-7|LNC|VLDL cholesterol|VLDL cholesterol
C0364227|T201|LN|2091-7|LNC|VLDL cholesterol|VLDL cholesterol
C0364227|T201|OSN|2091-7|LNC|VLDL cholesterol|VLDL cholesterol
C0364227|T201|LC|2091-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0364227|T201|MTH_LN|2091-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0364227|T201|LN|2091-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0364227|T201|OSN|2091-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0364227|T201|LC|2091-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0364227|T201|MTH_LN|2091-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0364227|T201|LN|2091-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0364227|T201|OSN|2091-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0364227|T201|LC|2091-7|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0364227|T201|MTH_LN|2091-7|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0364227|T201|LN|2091-7|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0364227|T201|OSN|2091-7|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0364238|T201|LN|2118-8|LNC|maternal chorionic gonadotropin|maternal chorionic gonadotropin
C0364238|T201|MTH_LN|2118-8|LNC|maternal chorionic gonadotropin|maternal chorionic gonadotropin
C0364238|T201|LC|2118-8|LNC|maternal chorionic gonadotropin|maternal chorionic gonadotropin
C0364238|T201|OSN|2118-8|LNC|maternal chorionic gonadotropin|maternal chorionic gonadotropin
C0364238|T201|LN|2118-8|LNC|maternal hCG|maternal hCG
C0364238|T201|MTH_LN|2118-8|LNC|maternal hCG|maternal hCG
C0364238|T201|LC|2118-8|LNC|maternal hCG|maternal hCG
C0364238|T201|OSN|2118-8|LNC|maternal hCG|maternal hCG
C0364238|T201|LN|2118-8|LNC|maternal screening|maternal screening
C0364238|T201|MTH_LN|2118-8|LNC|maternal screening|maternal screening
C0364238|T201|LC|2118-8|LNC|maternal screening|maternal screening
C0364238|T201|OSN|2118-8|LNC|maternal screening|maternal screening
C0364264|T201|LC|2132-9|LNC|vitamin B12|vitamin B12
C0364264|T201|MTH_LN|2132-9|LNC|vitamin B12|vitamin B12
C0364264|T201|OSN|2132-9|LNC|vitamin B12|vitamin B12
C0364264|T201|LN|2132-9|LNC|vitamin B12|vitamin B12
C0364264|T201|LC|2132-9|LNC|cobalamin|cobalamin
C0364264|T201|MTH_LN|2132-9|LNC|cobalamin|cobalamin
C0364264|T201|OSN|2132-9|LNC|cobalamin|cobalamin
C0364264|T201|LN|2132-9|LNC|cobalamin|cobalamin
C0364271|T201|LN|2139-4|LNC|corticosterone|corticosterone
C0364271|T201|MTH_LN|2139-4|LNC|corticosterone|corticosterone
C0364271|T201|LC|2139-4|LNC|corticosterone|corticosterone
C0364271|T201|OSN|2139-4|LNC|corticosterone|corticosterone
C0364273|T201|LC|2141-0|LNC|ACTH|ACTH
C0364273|T201|MTH_LN|2141-0|LNC|ACTH|ACTH
C0364273|T201|LN|2141-0|LNC|ACTH|ACTH
C0364273|T201|OSN|2141-0|LNC|ACTH|ACTH
C0364273|T201|LC|2141-0|LNC|corticotropin|corticotropin
C0364273|T201|MTH_LN|2141-0|LNC|corticotropin|corticotropin
C0364273|T201|LN|2141-0|LNC|corticotropin|corticotropin
C0364273|T201|OSN|2141-0|LNC|corticotropin|corticotropin
C0364273|T201|LC|2141-0|LNC|adrenocorticotropin|adrenocorticotropin
C0364273|T201|MTH_LN|2141-0|LNC|adrenocorticotropin|adrenocorticotropin
C0364273|T201|LN|2141-0|LNC|adrenocorticotropin|adrenocorticotropin
C0364273|T201|OSN|2141-0|LNC|adrenocorticotropin|adrenocorticotropin
C0364275|T201|LN|2143-6|LNC|cortisol|cortisol
C0364275|T201|MTH_LN|2143-6|LNC|cortisol|cortisol
C0364275|T201|OSN|2143-6|LNC|cortisol|cortisol
C0364275|T201|LC|2143-6|LNC|cortisol|cortisol
C0364275|T201|LN|2143-6|LNC|cortisol low|cortisol low
C0364275|T201|MTH_LN|2143-6|LNC|cortisol low|cortisol low
C0364275|T201|OSN|2143-6|LNC|cortisol low|cortisol low
C0364275|T201|LC|2143-6|LNC|cortisol low|cortisol low
C0364275|T201|LN|2143-6|LNC|to undetectable cortisol|to undetectable cortisol
C0364275|T201|MTH_LN|2143-6|LNC|to undetectable cortisol|to undetectable cortisol
C0364275|T201|OSN|2143-6|LNC|to undetectable cortisol|to undetectable cortisol
C0364275|T201|LC|2143-6|LNC|to undetectable cortisol|to undetectable cortisol
C0364290|T201|LN|2157-6|LNC|creatine phosphokinase|creatine phosphokinase
C0364290|T201|MTH_LN|2157-6|LNC|creatine phosphokinase|creatine phosphokinase
C0364290|T201|OSN|2157-6|LNC|creatine phosphokinase|creatine phosphokinase
C0364290|T201|LC|2157-6|LNC|creatine phosphokinase|creatine phosphokinase
C0364290|T201|LN|2157-6|LNC|CPK|CPK
C0364290|T201|MTH_LN|2157-6|LNC|CPK|CPK
C0364290|T201|OSN|2157-6|LNC|CPK|CPK
C0364290|T201|LC|2157-6|LNC|CPK|CPK
C0364290|T201|LN|2157-6|LNC|creatine kinase|creatine kinase
C0364290|T201|MTH_LN|2157-6|LNC|creatine kinase|creatine kinase
C0364290|T201|OSN|2157-6|LNC|creatine kinase|creatine kinase
C0364290|T201|LC|2157-6|LNC|creatine kinase|creatine kinase
C0364290|T201|LN|2157-6|LNC|CK|CK
C0364290|T201|MTH_LN|2157-6|LNC|CK|CK
C0364290|T201|OSN|2157-6|LNC|CK|CK
C0364290|T201|LC|2157-6|LNC|CK|CK
C0364294|T201|LC|2160-0|LNC|creatinine|creatinine
C0364294|T201|LN|2160-0|LNC|creatinine|creatinine
C0364294|T201|MTH_LN|2160-0|LNC|creatinine|creatinine
C0364294|T201|OSN|2160-0|LNC|creatinine|creatinine
C0364295|T201|LN|2161-8|LNC|creatinine|creatinine
C0364295|T201|MTH_LN|2161-8|LNC|creatinine|creatinine
C0364295|T201|OSN|2161-8|LNC|creatinine|creatinine
C0364295|T201|LC|2161-8|LNC|creatinine|creatinine
C0364295|T201|LN|2161-8|LNC|metabolism/homeostasis|metabolism/homeostasis
C0364295|T201|MTH_LN|2161-8|LNC|metabolism/homeostasis|metabolism/homeostasis
C0364295|T201|OSN|2161-8|LNC|metabolism/homeostasis|metabolism/homeostasis
C0364295|T201|LC|2161-8|LNC|metabolism/homeostasis|metabolism/homeostasis
C0364295|T201|LN|2161-8|LNC|Metabolism|Metabolism
C0364295|T201|MTH_LN|2161-8|LNC|Metabolism|Metabolism
C0364295|T201|OSN|2161-8|LNC|Metabolism|Metabolism
C0364295|T201|LC|2161-8|LNC|Metabolism|Metabolism
C0364295|T201|LN|2161-8|LNC|Laboratory|Laboratory
C0364295|T201|MTH_LN|2161-8|LNC|Laboratory|Laboratory
C0364295|T201|OSN|2161-8|LNC|Laboratory|Laboratory
C0364295|T201|LC|2161-8|LNC|Laboratory|Laboratory
C0364325|T201|LN|2191-5|LNC|dehydroepiandrosterone-sulfate|dehydroepiandrosterone-sulfate
C0364325|T201|MTH_LN|2191-5|LNC|dehydroepiandrosterone-sulfate|dehydroepiandrosterone-sulfate
C0364325|T201|OSN|2191-5|LNC|dehydroepiandrosterone-sulfate|dehydroepiandrosterone-sulfate
C0364325|T201|LC|2191-5|LNC|dehydroepiandrosterone-sulfate|dehydroepiandrosterone-sulfate
C0364327|T201|MTH_LN|2193-1|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C0364327|T201|LN|2193-1|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C0364327|T201|OSN|2193-1|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C0364327|T201|LC|2193-1|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C0364352|T201|LN|2218-6|LNC|catecholamine|catecholamine
C0364352|T201|MTH_LN|2218-6|LNC|catecholamine|catecholamine
C0364352|T201|OSN|2218-6|LNC|catecholamine|catecholamine
C0364352|T201|LC|2218-6|LNC|catecholamine|catecholamine
C0364352|T201|LN|2218-6|LNC|dopamine|dopamine
C0364352|T201|MTH_LN|2218-6|LNC|dopamine|dopamine
C0364352|T201|OSN|2218-6|LNC|dopamine|dopamine
C0364352|T201|LC|2218-6|LNC|dopamine|dopamine
C0364378|T201|LN|2243-4|LNC|estradiol|estradiol
C0364378|T201|LC|2243-4|LNC|estradiol|estradiol
C0364378|T201|MTH_LN|2243-4|LNC|estradiol|estradiol
C0364378|T201|OSN|2243-4|LNC|estradiol|estradiol
C0364378|T201|LN|2243-4|LNC|oestradiol|oestradiol
C0364378|T201|LC|2243-4|LNC|oestradiol|oestradiol
C0364378|T201|MTH_LN|2243-4|LNC|oestradiol|oestradiol
C0364378|T201|OSN|2243-4|LNC|oestradiol|oestradiol
C0364393|T201|LN|2258-2|LNC|estradiol|estradiol
C0364393|T201|MTH_LN|2258-2|LNC|estradiol|estradiol
C0364393|T201|OSN|2258-2|LNC|estradiol|estradiol
C0364393|T201|LC|2258-2|LNC|estradiol|estradiol
C0364393|T201|LN|2258-2|LNC|estrone|estrone
C0364393|T201|MTH_LN|2258-2|LNC|estrone|estrone
C0364393|T201|OSN|2258-2|LNC|estrone|estrone
C0364393|T201|LC|2258-2|LNC|estrone|estrone
C0364411|T201|LC|2276-4|LNC|ferritin|ferritin
C0364411|T201|MTH_LN|2276-4|LNC|ferritin|ferritin
C0364411|T201|LN|2276-4|LNC|ferritin|ferritin
C0364411|T201|OSN|2276-4|LNC|ferritin|ferritin
C0364417|T201|LN|2282-2|LNC|folate metabolism|folate metabolism
C0364417|T201|MTH_LN|2282-2|LNC|folate metabolism|folate metabolism
C0364417|T201|OSN|2282-2|LNC|folate metabolism|folate metabolism
C0364417|T201|LC|2282-2|LNC|folate metabolism|folate metabolism
C0364418|T201|LN|2283-0|LNC|folate metabolism|folate metabolism
C0364418|T201|MTH_LN|2283-0|LNC|folate metabolism|folate metabolism
C0364418|T201|OSN|2283-0|LNC|folate metabolism|folate metabolism
C0364418|T201|LC|2283-0|LNC|folate metabolism|folate metabolism
C0364419|T201|LC|2284-8|LNC|folate metabolism|folate metabolism
C0364419|T201|OSN|2284-8|LNC|folate metabolism|folate metabolism
C0364419|T201|LN|2284-8|LNC|folate metabolism|folate metabolism
C0364419|T201|MTH_LN|2284-8|LNC|folate metabolism|folate metabolism
C0364425|T201|LN|2290-5|LNC|luteinizing|luteinizing
C0364425|T201|OSN|2290-5|LNC|luteinizing|luteinizing
C0364425|T201|LC|2290-5|LNC|luteinizing|luteinizing
C0364425|T201|MTH_LN|2290-5|LNC|luteinizing|luteinizing
C0364425|T201|LN|2290-5|LNC|LH|LH
C0364425|T201|OSN|2290-5|LNC|LH|LH
C0364425|T201|LC|2290-5|LNC|LH|LH
C0364425|T201|MTH_LN|2290-5|LNC|LH|LH
C0364425|T201|LN|2290-5|LNC|luteinising|luteinising
C0364425|T201|OSN|2290-5|LNC|luteinising|luteinising
C0364425|T201|LC|2290-5|LNC|luteinising|luteinising
C0364425|T201|MTH_LN|2290-5|LNC|luteinising|luteinising
C0364444|T201|LN|2309-3|LNC|galactose|galactose
C0364444|T201|MTH_LN|2309-3|LNC|galactose|galactose
C0364444|T201|OSN|2309-3|LNC|galactose|galactose
C0364444|T201|LC|2309-3|LNC|galactose|galactose
C0364445|T201|LN|2310-1|LNC|galactose|galactose
C0364445|T201|MTH_LN|2310-1|LNC|galactose|galactose
C0364445|T201|OSN|2310-1|LNC|galactose|galactose
C0364445|T201|LC|2310-1|LNC|galactose|galactose
C0364459|T201|LN|2324-2|LNC|gamma-glutamyltransferase activity|gamma-glutamyltransferase activity
C0364459|T201|MTH_LN|2324-2|LNC|gamma-glutamyltransferase activity|gamma-glutamyltransferase activity
C0364459|T201|OSN|2324-2|LNC|gamma-glutamyltransferase activity|gamma-glutamyltransferase activity
C0364459|T201|LC|2324-2|LNC|gamma-glutamyltransferase activity|gamma-glutamyltransferase activity
C0364479|T201|LN|2339-0|LNC|glucose|glucose
C0364479|T201|MTH_LN|2339-0|LNC|glucose|glucose
C0364479|T201|OSN|2339-0|LNC|glucose|glucose
C0364479|T201|LC|2339-0|LNC|glucose|glucose
C0364480|T201|LN|2340-8|LNC|glucose|glucose
C0364480|T201|OSN|2340-8|LNC|glucose|glucose
C0364480|T201|LC|2340-8|LNC|glucose|glucose
C0364480|T201|MTH_LN|2340-8|LNC|glucose|glucose
C0364481|T201|LN|2341-6|LNC|glucose|glucose
C0364481|T201|MTH_LN|2341-6|LNC|glucose|glucose
C0364481|T201|OSN|2341-6|LNC|glucose|glucose
C0364481|T201|LC|2341-6|LNC|glucose|glucose
C0364482|T201|LN|2342-4|LNC|CSF glucose|CSF glucose
C0364482|T201|MTH_LN|2342-4|LNC|CSF glucose|CSF glucose
C0364482|T201|OSN|2342-4|LNC|CSF glucose|CSF glucose
C0364482|T201|LC|2342-4|LNC|CSF glucose|CSF glucose
C0364482|T201|LN|2342-4|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C0364482|T201|MTH_LN|2342-4|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C0364482|T201|OSN|2342-4|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C0364482|T201|LC|2342-4|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C0364490|T201|LC|2350-7|LNC|glucose|glucose
C0364490|T201|MTH_LN|2350-7|LNC|glucose|glucose
C0364490|T201|OSN|2350-7|LNC|glucose|glucose
C0364490|T201|LN|2350-7|LNC|glucose|glucose
C0364491|T201|LN|2351-5|LNC|glucose|glucose
C0364491|T201|MTH_LN|2351-5|LNC|glucose|glucose
C0364491|T201|OSN|2351-5|LNC|glucose|glucose
C0364491|T201|LC|2351-5|LNC|glucose|glucose
C0364496|T201|LN|2356-4|LNC|glucose-6-phosphate dehydrogenase in red|glucose-6-phosphate dehydrogenase in red
C0364496|T201|MTH_LN|2356-4|LNC|glucose-6-phosphate dehydrogenase in red|glucose-6-phosphate dehydrogenase in red
C0364496|T201|OSN|2356-4|LNC|glucose-6-phosphate dehydrogenase in red|glucose-6-phosphate dehydrogenase in red
C0364496|T201|LC|2356-4|LNC|glucose-6-phosphate dehydrogenase in red|glucose-6-phosphate dehydrogenase in red
C0364496|T201|LN|2356-4|LNC|G6PD in red|G6PD in red
C0364496|T201|MTH_LN|2356-4|LNC|G6PD in red|G6PD in red
C0364496|T201|OSN|2356-4|LNC|G6PD in red|G6PD in red
C0364496|T201|LC|2356-4|LNC|G6PD in red|G6PD in red
C0364498|T201|LN|2358-0|LNC|glucose-6-phosphate dehydrogenase|glucose-6-phosphate dehydrogenase
C0364498|T201|MTH_LN|2358-0|LNC|glucose-6-phosphate dehydrogenase|glucose-6-phosphate dehydrogenase
C0364498|T201|OSN|2358-0|LNC|glucose-6-phosphate dehydrogenase|glucose-6-phosphate dehydrogenase
C0364498|T201|LC|2358-0|LNC|glucose-6-phosphate dehydrogenase|glucose-6-phosphate dehydrogenase
C0364498|T201|LN|2358-0|LNC|G6PD|G6PD
C0364498|T201|MTH_LN|2358-0|LNC|G6PD|G6PD
C0364498|T201|OSN|2358-0|LNC|G6PD|G6PD
C0364498|T201|LC|2358-0|LNC|G6PD|G6PD
C0364500|T201|LN|2360-6|LNC|glucose-6-phosphate dehydrogenase in leukocytes|glucose-6-phosphate dehydrogenase in leukocytes
C0364500|T201|MTH_LN|2360-6|LNC|glucose-6-phosphate dehydrogenase in leukocytes|glucose-6-phosphate dehydrogenase in leukocytes
C0364500|T201|OSN|2360-6|LNC|glucose-6-phosphate dehydrogenase in leukocytes|glucose-6-phosphate dehydrogenase in leukocytes
C0364500|T201|LC|2360-6|LNC|glucose-6-phosphate dehydrogenase in leukocytes|glucose-6-phosphate dehydrogenase in leukocytes
C0364500|T201|LN|2360-6|LNC|G6PD in leukocytes|G6PD in leukocytes
C0364500|T201|MTH_LN|2360-6|LNC|G6PD in leukocytes|G6PD in leukocytes
C0364500|T201|OSN|2360-6|LNC|G6PD in leukocytes|G6PD in leukocytes
C0364500|T201|LC|2360-6|LNC|G6PD in leukocytes|G6PD in leukocytes
C0364598|T201|LN|2458-8|LNC|IgA|IgA
C0364598|T201|OSN|2458-8|LNC|IgA|IgA
C0364598|T201|LC|2458-8|LNC|IgA|IgA
C0364598|T201|MTH_LN|2458-8|LNC|IgA|IgA
C0364598|T201|LN|2458-8|LNC|immunoglobulin A|immunoglobulin A
C0364598|T201|OSN|2458-8|LNC|immunoglobulin A|immunoglobulin A
C0364598|T201|LC|2458-8|LNC|immunoglobulin A|immunoglobulin A
C0364598|T201|MTH_LN|2458-8|LNC|immunoglobulin A|immunoglobulin A
C0364605|T201|LN|2465-3|LNC|IgG|IgG
C0364605|T201|LC|2465-3|LNC|IgG|IgG
C0364605|T201|OSN|2465-3|LNC|IgG|IgG
C0364605|T201|MTH_LN|2465-3|LNC|IgG|IgG
C0364605|T201|LN|2465-3|LNC|gamma-globin expression|gamma-globin expression
C0364605|T201|LC|2465-3|LNC|gamma-globin expression|gamma-globin expression
C0364605|T201|OSN|2465-3|LNC|gamma-globin expression|gamma-globin expression
C0364605|T201|MTH_LN|2465-3|LNC|gamma-globin expression|gamma-globin expression
C0364605|T201|LN|2465-3|LNC|immunoglobulin G|immunoglobulin G
C0364605|T201|LC|2465-3|LNC|immunoglobulin G|immunoglobulin G
C0364605|T201|OSN|2465-3|LNC|immunoglobulin G|immunoglobulin G
C0364605|T201|MTH_LN|2465-3|LNC|immunoglobulin G|immunoglobulin G
C0364607|T201|LN|2467-9|LNC|IgG2|IgG2
C0364607|T201|MTH_LN|2467-9|LNC|IgG2|IgG2
C0364607|T201|OSN|2467-9|LNC|IgG2|IgG2
C0364607|T201|LC|2467-9|LNC|IgG2|IgG2
C0364612|T201|LN|2472-9|LNC|IgM|IgM
C0364612|T201|OSN|2472-9|LNC|IgM|IgM
C0364612|T201|MTH_LN|2472-9|LNC|IgM|IgM
C0364612|T201|LC|2472-9|LNC|IgM|IgM
C0364626|T201|LC|2484-4|LNC|insulin-like growth factor 1|insulin-like growth factor 1
C0364626|T201|MTH_LN|2484-4|LNC|insulin-like growth factor 1|insulin-like growth factor 1
C0364626|T201|LN|2484-4|LNC|insulin-like growth factor 1|insulin-like growth factor 1
C0364626|T201|OSN|2484-4|LNC|insulin-like growth factor 1|insulin-like growth factor 1
C0364626|T201|LC|2484-4|LNC|IGF1|IGF1
C0364626|T201|MTH_LN|2484-4|LNC|IGF1|IGF1
C0364626|T201|LN|2484-4|LNC|IGF1|IGF1
C0364626|T201|OSN|2484-4|LNC|IGF1|IGF1
C0364639|T201|LC|2498-4|LNC|iron|iron
C0364639|T201|MTH_LN|2498-4|LNC|iron|iron
C0364639|T201|LN|2498-4|LNC|iron|iron
C0364639|T201|OSN|2498-4|LNC|iron|iron
C0364641|T201|LC|2500-7|LNC|total iron binding capacity|total iron binding capacity
C0364641|T201|MTH_LN|2500-7|LNC|total iron binding capacity|total iron binding capacity
C0364641|T201|LN|2500-7|LNC|total iron binding capacity|total iron binding capacity
C0364641|T201|OSN|2500-7|LNC|total iron binding capacity|total iron binding capacity
C0364641|T201|LC|2500-7|LNC|iron homeostasis|iron homeostasis
C0364641|T201|MTH_LN|2500-7|LNC|iron homeostasis|iron homeostasis
C0364641|T201|LN|2500-7|LNC|iron homeostasis|iron homeostasis
C0364641|T201|OSN|2500-7|LNC|iron homeostasis|iron homeostasis
C0364643|T201|LN|2502-3|LNC|iron|iron
C0364643|T201|LC|2502-3|LNC|iron|iron
C0364643|T201|OSN|2502-3|LNC|iron|iron
C0364643|T201|MTH_LN|2502-3|LNC|iron|iron
C0364654|T201|LN|2513-0|LNC|ketone bodies|ketone bodies
C0364654|T201|MTH_LN|2513-0|LNC|ketone bodies|ketone bodies
C0364654|T201|OSN|2513-0|LNC|ketone bodies|ketone bodies
C0364654|T201|LC|2513-0|LNC|ketone bodies|ketone bodies
C0364659|T201|LN|2518-9|LNC|lactate|lactate
C0364659|T201|MTH_LN|2518-9|LNC|lactate|lactate
C0364659|T201|OSN|2518-9|LNC|lactate|lactate
C0364659|T201|LC|2518-9|LNC|lactate|lactate
C0364660|T201|LN|2519-7|LNC|lactate|lactate
C0364660|T201|MTH_LN|2519-7|LNC|lactate|lactate
C0364660|T201|OSN|2519-7|LNC|lactate|lactate
C0364660|T201|LC|2519-7|LNC|lactate|lactate
C0364661|T201|LN|2520-5|LNC|CSF lactate|CSF lactate
C0364661|T201|MTH_LN|2520-5|LNC|CSF lactate|CSF lactate
C0364661|T201|OSN|2520-5|LNC|CSF lactate|CSF lactate
C0364661|T201|LC|2520-5|LNC|CSF lactate|CSF lactate
C0364661|T201|LN|2520-5|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C0364661|T201|MTH_LN|2520-5|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C0364661|T201|OSN|2520-5|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C0364661|T201|LC|2520-5|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C0364661|T201|LN|2520-5|LNC|CSF lactic acid|CSF lactic acid
C0364661|T201|MTH_LN|2520-5|LNC|CSF lactic acid|CSF lactic acid
C0364661|T201|OSN|2520-5|LNC|CSF lactic acid|CSF lactic acid
C0364661|T201|LC|2520-5|LNC|CSF lactic acid|CSF lactic acid
C0364665|T201|LN|2524-7|LNC|lactate|lactate
C0364665|T201|MTH_LN|2524-7|LNC|lactate|lactate
C0364665|T201|OSN|2524-7|LNC|lactate|lactate
C0364665|T201|LC|2524-7|LNC|lactate|lactate
C0364674|T201|LN|2532-0|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0364674|T201|MTH_LN|2532-0|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0364674|T201|OSN|2532-0|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0364674|T201|LC|2532-0|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0364680|T201|LN|2537-9|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0364680|T201|MTH_LN|2537-9|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0364680|T201|OSN|2537-9|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0364680|T201|LC|2537-9|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0364693|T201|LN|2550-2|LNC|lactate|lactate
C0364693|T201|OSN|2550-2|LNC|lactate|lactate
C0364693|T201|LC|2550-2|LNC|lactate|lactate
C0364693|T201|MTH_LN|2550-2|LNC|lactate|lactate
C0364708|T201|MTH_LN|2093-3|LNC|cholesterol|cholesterol
C0364708|T201|LN|2093-3|LNC|cholesterol|cholesterol
C0364708|T201|OSN|2093-3|LNC|cholesterol|cholesterol
C0364708|T201|LC|2093-3|LNC|cholesterol|cholesterol
C0364708|T201|MTH_LN|2093-3|LNC|total cholesterol|total cholesterol
C0364708|T201|LN|2093-3|LNC|total cholesterol|total cholesterol
C0364708|T201|OSN|2093-3|LNC|total cholesterol|total cholesterol
C0364708|T201|LC|2093-3|LNC|total cholesterol|total cholesterol
C0364708|T201|MTH_LN|2093-3|LNC|cholesterol metabolism|cholesterol metabolism
C0364708|T201|LN|2093-3|LNC|cholesterol metabolism|cholesterol metabolism
C0364708|T201|OSN|2093-3|LNC|cholesterol metabolism|cholesterol metabolism
C0364708|T201|LC|2093-3|LNC|cholesterol metabolism|cholesterol metabolism
C0364712|T201|LN|2569-2|LNC|lipid metabolism|lipid metabolism
C0364712|T201|MTH_LN|2569-2|LNC|lipid metabolism|lipid metabolism
C0364712|T201|OSN|2569-2|LNC|lipid metabolism|lipid metabolism
C0364712|T201|LC|2569-2|LNC|lipid metabolism|lipid metabolism
C0364714|T201|LC|2571-8|LNC|triglyceride|triglyceride
C0364714|T201|MTH_LN|2571-8|LNC|triglyceride|triglyceride
C0364714|T201|LN|2571-8|LNC|triglyceride|triglyceride
C0364714|T201|OSN|2571-8|LNC|triglyceride|triglyceride
C0364714|T201|LC|2571-8|LNC|Tg|Tg
C0364714|T201|MTH_LN|2571-8|LNC|Tg|Tg
C0364714|T201|LN|2571-8|LNC|Tg|Tg
C0364714|T201|OSN|2571-8|LNC|Tg|Tg
C0364714|T201|LC|2571-8|LNC|triglycerides|triglycerides
C0364714|T201|MTH_LN|2571-8|LNC|triglycerides|triglycerides
C0364714|T201|LN|2571-8|LNC|triglycerides|triglycerides
C0364714|T201|OSN|2571-8|LNC|triglycerides|triglycerides
C0364714|T201|LC|2571-8|LNC|lipid metabolism|lipid metabolism
C0364714|T201|MTH_LN|2571-8|LNC|lipid metabolism|lipid metabolism
C0364714|T201|LN|2571-8|LNC|lipid metabolism|lipid metabolism
C0364714|T201|OSN|2571-8|LNC|lipid metabolism|lipid metabolism
C0364716|T201|LN|2572-6|LNC|enzyme/coenzyme activity|enzyme/coenzyme activity
C0364716|T201|MTH_LN|2572-6|LNC|enzyme/coenzyme activity|enzyme/coenzyme activity
C0364716|T201|OSN|2572-6|LNC|enzyme/coenzyme activity|enzyme/coenzyme activity
C0364716|T201|LC|2572-6|LNC|enzyme/coenzyme activity|enzyme/coenzyme activity
C0364716|T201|LN|2572-6|LNC|lipoprotein lipase activity|lipoprotein lipase activity
C0364716|T201|MTH_LN|2572-6|LNC|lipoprotein lipase activity|lipoprotein lipase activity
C0364716|T201|OSN|2572-6|LNC|lipoprotein lipase activity|lipoprotein lipase activity
C0364716|T201|LC|2572-6|LNC|lipoprotein lipase activity|lipoprotein lipase activity
C0364722|T201|LN|2578-3|LNC|luteinizing|luteinizing
C0364722|T201|MTH_LN|2578-3|LNC|luteinizing|luteinizing
C0364722|T201|OSN|2578-3|LNC|luteinizing|luteinizing
C0364722|T201|LC|2578-3|LNC|luteinizing|luteinizing
C0364722|T201|LN|2578-3|LNC|LH|LH
C0364722|T201|MTH_LN|2578-3|LNC|LH|LH
C0364722|T201|OSN|2578-3|LNC|LH|LH
C0364722|T201|LC|2578-3|LNC|LH|LH
C0364722|T201|LN|2578-3|LNC|luteinising|luteinising
C0364722|T201|MTH_LN|2578-3|LNC|luteinising|luteinising
C0364722|T201|OSN|2578-3|LNC|luteinising|luteinising
C0364722|T201|LC|2578-3|LNC|luteinising|luteinising
C0364723|T201|LN|2579-1|LNC|luteinizing|luteinizing
C0364723|T201|MTH_LN|2579-1|LNC|luteinizing|luteinizing
C0364723|T201|OSN|2579-1|LNC|luteinizing|luteinizing
C0364723|T201|LC|2579-1|LNC|luteinizing|luteinizing
C0364723|T201|LN|2579-1|LNC|LH|LH
C0364723|T201|MTH_LN|2579-1|LNC|LH|LH
C0364723|T201|OSN|2579-1|LNC|LH|LH
C0364723|T201|LC|2579-1|LNC|LH|LH
C0364723|T201|LN|2579-1|LNC|luteinising|luteinising
C0364723|T201|MTH_LN|2579-1|LNC|luteinising|luteinising
C0364723|T201|OSN|2579-1|LNC|luteinising|luteinising
C0364723|T201|LC|2579-1|LNC|luteinising|luteinising
C0364726|T201|LN|2582-5|LNC|luteinizing|luteinizing
C0364726|T201|OSN|2582-5|LNC|luteinizing|luteinizing
C0364726|T201|MTH_LN|2582-5|LNC|luteinizing|luteinizing
C0364726|T201|LC|2582-5|LNC|luteinizing|luteinizing
C0364726|T201|LN|2582-5|LNC|LH|LH
C0364726|T201|OSN|2582-5|LNC|LH|LH
C0364726|T201|MTH_LN|2582-5|LNC|LH|LH
C0364726|T201|LC|2582-5|LNC|LH|LH
C0364726|T201|LN|2582-5|LNC|luteinising|luteinising
C0364726|T201|OSN|2582-5|LNC|luteinising|luteinising
C0364726|T201|MTH_LN|2582-5|LNC|luteinising|luteinising
C0364726|T201|LC|2582-5|LNC|luteinising|luteinising
C0364727|T201|LN|2583-3|LNC|luteinizing|luteinizing
C0364727|T201|OSN|2583-3|LNC|luteinizing|luteinizing
C0364727|T201|MTH_LN|2583-3|LNC|luteinizing|luteinizing
C0364727|T201|LC|2583-3|LNC|luteinizing|luteinizing
C0364727|T201|LN|2583-3|LNC|LH|LH
C0364727|T201|OSN|2583-3|LNC|LH|LH
C0364727|T201|MTH_LN|2583-3|LNC|LH|LH
C0364727|T201|LC|2583-3|LNC|LH|LH
C0364727|T201|LN|2583-3|LNC|luteinising|luteinising
C0364727|T201|OSN|2583-3|LNC|luteinising|luteinising
C0364727|T201|MTH_LN|2583-3|LNC|luteinising|luteinising
C0364727|T201|LC|2583-3|LNC|luteinising|luteinising
C0364745|T201|MTH_LN|2601-3|LNC|magnesium|magnesium
C0364745|T201|LN|2601-3|LNC|magnesium|magnesium
C0364745|T201|OSN|2601-3|LNC|magnesium|magnesium
C0364745|T201|LC|2601-3|LNC|magnesium|magnesium
C0364745|T201|MTH_LN|2601-3|LNC|magnesium metabolism|magnesium metabolism
C0364745|T201|LN|2601-3|LNC|magnesium metabolism|magnesium metabolism
C0364745|T201|OSN|2601-3|LNC|magnesium metabolism|magnesium metabolism
C0364745|T201|LC|2601-3|LNC|magnesium metabolism|magnesium metabolism
C0364745|T201|MTH_LN|2601-3|LNC|magnesium homeostasis|magnesium homeostasis
C0364745|T201|LN|2601-3|LNC|magnesium homeostasis|magnesium homeostasis
C0364745|T201|OSN|2601-3|LNC|magnesium homeostasis|magnesium homeostasis
C0364745|T201|LC|2601-3|LNC|magnesium homeostasis|magnesium homeostasis
C0364840|T201|LC|2697-1|LNC|osteocalcin|osteocalcin
C0364840|T201|MTH_LN|2697-1|LNC|osteocalcin|osteocalcin
C0364840|T201|OSN|2697-1|LNC|osteocalcin|osteocalcin
C0364840|T201|LN|2697-1|LNC|osteocalcin|osteocalcin
C0364844|T201|LN|2701-1|LNC|oxalate|oxalate
C0364844|T201|MTH_LN|2701-1|LNC|oxalate|oxalate
C0364844|T201|OSN|2701-1|LNC|oxalate|oxalate
C0364844|T201|LC|2701-1|LNC|oxalate|oxalate
C0364846|T201|LN|19255-9|LNC|oxygen|oxygen
C0364846|T201|MTH_LN|19255-9|LNC|oxygen|oxygen
C0364846|T201|OSN|19255-9|LNC|oxygen|oxygen
C0364846|T201|LC|19255-9|LNC|oxygen|oxygen
C0364851|T201|LN|2708-6|LNC|oxygen|oxygen
C0364851|T201|LC|2708-6|LNC|oxygen|oxygen
C0364851|T201|MTH_LN|2708-6|LNC|oxygen|oxygen
C0364851|T201|OSN|2708-6|LNC|oxygen|oxygen
C0364852|T201|LN|2709-4|LNC|oxygen|oxygen
C0364852|T201|LC|2709-4|LNC|oxygen|oxygen
C0364852|T201|MTH_LN|2709-4|LNC|oxygen|oxygen
C0364852|T201|OSN|2709-4|LNC|oxygen|oxygen
C0364874|T201|LC|2731-8|LNC|parathyroid|parathyroid
C0364874|T201|MTH_LN|2731-8|LNC|parathyroid|parathyroid
C0364874|T201|LN|2731-8|LNC|parathyroid|parathyroid
C0364874|T201|OSN|2731-8|LNC|parathyroid|parathyroid
C0364874|T201|LC|2731-8|LNC|parathyroid physiology|parathyroid physiology
C0364874|T201|MTH_LN|2731-8|LNC|parathyroid physiology|parathyroid physiology
C0364874|T201|LN|2731-8|LNC|parathyroid physiology|parathyroid physiology
C0364874|T201|OSN|2731-8|LNC|parathyroid physiology|parathyroid physiology
C0364887|T201|LN|2744-1|LNC|acid-base homeostasis|acid-base homeostasis
C0364887|T201|LC|2744-1|LNC|acid-base homeostasis|acid-base homeostasis
C0364887|T201|MTH_LN|2744-1|LNC|acid-base homeostasis|acid-base homeostasis
C0364887|T201|OSN|2744-1|LNC|acid-base homeostasis|acid-base homeostasis
C0364888|T201|LN|2745-8|LNC|acid-base homeostasis|acid-base homeostasis
C0364888|T201|MTH_LN|2745-8|LNC|acid-base homeostasis|acid-base homeostasis
C0364888|T201|OSN|2745-8|LNC|acid-base homeostasis|acid-base homeostasis
C0364888|T201|LC|2745-8|LNC|acid-base homeostasis|acid-base homeostasis
C0364889|T201|LN|2746-6|LNC|acid-base homeostasis|acid-base homeostasis
C0364889|T201|LC|2746-6|LNC|acid-base homeostasis|acid-base homeostasis
C0364889|T201|MTH_LN|2746-6|LNC|acid-base homeostasis|acid-base homeostasis
C0364889|T201|OSN|2746-6|LNC|acid-base homeostasis|acid-base homeostasis
C0364896|T201|LN|2753-2|LNC|acid-base homeostasis|acid-base homeostasis
C0364896|T201|MTH_LN|2753-2|LNC|acid-base homeostasis|acid-base homeostasis
C0364896|T201|OSN|2753-2|LNC|acid-base homeostasis|acid-base homeostasis
C0364896|T201|LC|2753-2|LNC|acid-base homeostasis|acid-base homeostasis
C0364899|T201|LN|2756-5|LNC|acid-base homeostasis|acid-base homeostasis
C0364899|T201|LC|2756-5|LNC|acid-base homeostasis|acid-base homeostasis
C0364899|T201|MTH_LN|2756-5|LNC|acid-base homeostasis|acid-base homeostasis
C0364899|T201|OSN|2756-5|LNC|acid-base homeostasis|acid-base homeostasis
C0364906|T201|LN|2765-6|LNC|phenylalanine metabolism|phenylalanine metabolism
C0364906|T201|MTH_LN|2765-6|LNC|phenylalanine metabolism|phenylalanine metabolism
C0364906|T201|OSN|2765-6|LNC|phenylalanine metabolism|phenylalanine metabolism
C0364906|T201|LC|2765-6|LNC|phenylalanine metabolism|phenylalanine metabolism
C0364961|T201|LN|6298-4|LNC|potassium|potassium
C0364961|T201|MTH_LN|6298-4|LNC|potassium|potassium
C0364961|T201|OSN|6298-4|LNC|potassium|potassium
C0364961|T201|LC|6298-4|LNC|potassium|potassium
C0364961|T201|LN|6298-4|LNC|potassium homeostasis|potassium homeostasis
C0364961|T201|MTH_LN|6298-4|LNC|potassium homeostasis|potassium homeostasis
C0364961|T201|OSN|6298-4|LNC|potassium homeostasis|potassium homeostasis
C0364961|T201|LC|6298-4|LNC|potassium homeostasis|potassium homeostasis
C0364968|T201|LN|2823-3|LNC|potassium|potassium
C0364968|T201|MTH_LN|2823-3|LNC|potassium|potassium
C0364968|T201|OSN|2823-3|LNC|potassium|potassium
C0364968|T201|LC|2823-3|LNC|potassium|potassium
C0364968|T201|LN|2823-3|LNC|potassium homeostasis|potassium homeostasis
C0364968|T201|MTH_LN|2823-3|LNC|potassium homeostasis|potassium homeostasis
C0364968|T201|OSN|2823-3|LNC|potassium homeostasis|potassium homeostasis
C0364968|T201|LC|2823-3|LNC|potassium homeostasis|potassium homeostasis
C0364971|T201|LN|2828-2|LNC|potassium|potassium
C0364971|T201|MTH_LN|2828-2|LNC|potassium|potassium
C0364971|T201|OSN|2828-2|LNC|potassium|potassium
C0364971|T201|LC|2828-2|LNC|potassium|potassium
C0364972|T201|LN|2829-0|LNC|potassium|potassium
C0364972|T201|MTH_LN|2829-0|LNC|potassium|potassium
C0364972|T201|OSN|2829-0|LNC|potassium|potassium
C0364972|T201|LC|2829-0|LNC|potassium|potassium
C0365000|T201|LN|2857-1|LNC|Serum protein|Serum protein
C0365000|T201|MTH_LN|2857-1|LNC|Serum protein|Serum protein
C0365000|T201|OSN|2857-1|LNC|Serum protein|Serum protein
C0365000|T201|LC|2857-1|LNC|Serum protein|Serum protein
C0365000|T201|LN|2857-1|LNC|protein disease|protein disease
C0365000|T201|MTH_LN|2857-1|LNC|protein disease|protein disease
C0365000|T201|OSN|2857-1|LNC|protein disease|protein disease
C0365000|T201|LC|2857-1|LNC|protein disease|protein disease
C0365000|T201|LN|2857-1|LNC|protein|protein
C0365000|T201|MTH_LN|2857-1|LNC|protein|protein
C0365000|T201|OSN|2857-1|LNC|protein|protein
C0365000|T201|LC|2857-1|LNC|protein|protein
C0365000|T201|LN|2857-1|LNC|prostate-specific antigen|prostate-specific antigen
C0365000|T201|MTH_LN|2857-1|LNC|prostate-specific antigen|prostate-specific antigen
C0365000|T201|OSN|2857-1|LNC|prostate-specific antigen|prostate-specific antigen
C0365000|T201|LC|2857-1|LNC|prostate-specific antigen|prostate-specific antigen
C0365005|T201|LN|2862-1|LNC|albumin|albumin
C0365005|T201|MTH_LN|2862-1|LNC|albumin|albumin
C0365005|T201|OSN|2862-1|LNC|albumin|albumin
C0365005|T201|LC|2862-1|LNC|albumin|albumin
C0365014|T201|LN|2871-2|LNC|beta globulin|beta globulin
C0365014|T201|OSN|2871-2|LNC|beta globulin|beta globulin
C0365014|T201|MTH_LN|2871-2|LNC|beta globulin|beta globulin
C0365014|T201|LC|2871-2|LNC|beta globulin|beta globulin
C0365023|T201|LN|2880-3|LNC|CSF protein|CSF protein
C0365023|T201|MTH_LN|2880-3|LNC|CSF protein|CSF protein
C0365023|T201|OSN|2880-3|LNC|CSF protein|CSF protein
C0365023|T201|LC|2880-3|LNC|CSF protein|CSF protein
C0365023|T201|LN|2880-3|LNC|protein in csf|protein in csf
C0365023|T201|MTH_LN|2880-3|LNC|protein in csf|protein in csf
C0365023|T201|OSN|2880-3|LNC|protein in csf|protein in csf
C0365023|T201|LC|2880-3|LNC|protein in csf|protein in csf
C0365023|T201|LN|2880-3|LNC|Spinal fluid protein|Spinal fluid protein
C0365023|T201|MTH_LN|2880-3|LNC|Spinal fluid protein|Spinal fluid protein
C0365023|T201|OSN|2880-3|LNC|Spinal fluid protein|Spinal fluid protein
C0365023|T201|LC|2880-3|LNC|Spinal fluid protein|Spinal fluid protein
C0365023|T201|LN|2880-3|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C0365023|T201|MTH_LN|2880-3|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C0365023|T201|OSN|2880-3|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C0365023|T201|LC|2880-3|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C0365023|T201|LN|2880-3|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C0365023|T201|MTH_LN|2880-3|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C0365023|T201|OSN|2880-3|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C0365023|T201|LC|2880-3|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C0365023|T201|LN|2880-3|LNC|CSF total protein|CSF total protein
C0365023|T201|MTH_LN|2880-3|LNC|CSF total protein|CSF total protein
C0365023|T201|OSN|2880-3|LNC|CSF total protein|CSF total protein
C0365023|T201|LC|2880-3|LNC|CSF total protein|CSF total protein
C0365023|T201|LN|2880-3|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C0365023|T201|MTH_LN|2880-3|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C0365023|T201|OSN|2880-3|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C0365023|T201|LC|2880-3|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C0365029|T201|LN|2885-2|LNC|Serum protein|Serum protein
C0365029|T201|MTH_LN|2885-2|LNC|Serum protein|Serum protein
C0365029|T201|OSN|2885-2|LNC|Serum protein|Serum protein
C0365029|T201|LC|2885-2|LNC|Serum protein|Serum protein
C0365029|T201|LN|2885-2|LNC|protein disease|protein disease
C0365029|T201|MTH_LN|2885-2|LNC|protein disease|protein disease
C0365029|T201|OSN|2885-2|LNC|protein disease|protein disease
C0365029|T201|LC|2885-2|LNC|protein disease|protein disease
C0365029|T201|LN|2885-2|LNC|protein|protein
C0365029|T201|MTH_LN|2885-2|LNC|protein|protein
C0365029|T201|OSN|2885-2|LNC|protein|protein
C0365029|T201|LC|2885-2|LNC|protein|protein
C0365032|T201|LN|2888-6|LNC|Protein|Protein
C0365032|T201|MTH_LN|2888-6|LNC|Protein|Protein
C0365032|T201|OSN|2888-6|LNC|Protein|Protein
C0365032|T201|LC|2888-6|LNC|Protein|Protein
C0365034|T201|LN|2890-2|LNC|Protein|Protein
C0365034|T201|OSN|2890-2|LNC|Protein|Protein
C0365034|T201|MTH_LN|2890-2|LNC|Protein|Protein
C0365034|T201|LC|2890-2|LNC|Protein|Protein
C0365059|T201|LN|2915-7|LNC|renin|renin
C0365059|T201|MTH_LN|2915-7|LNC|renin|renin
C0365059|T201|OSN|2915-7|LNC|renin|renin
C0365059|T201|LC|2915-7|LNC|renin|renin
C0365059|T201|LN|2915-7|LNC|Suppressed renin activity|Suppressed renin activity
C0365059|T201|MTH_LN|2915-7|LNC|Suppressed renin activity|Suppressed renin activity
C0365059|T201|OSN|2915-7|LNC|Suppressed renin activity|Suppressed renin activity
C0365059|T201|LC|2915-7|LNC|Suppressed renin activity|Suppressed renin activity
C0365059|T201|LN|2915-7|LNC|renin activity|renin activity
C0365059|T201|MTH_LN|2915-7|LNC|renin activity|renin activity
C0365059|T201|OSN|2915-7|LNC|renin activity|renin activity
C0365059|T201|LC|2915-7|LNC|renin activity|renin activity
C0365086|T201|LN|2942-1|LNC|sex-binding globulin|sex-binding globulin
C0365086|T201|OSN|2942-1|LNC|sex-binding globulin|sex-binding globulin
C0365086|T201|MTH_LN|2942-1|LNC|sex-binding globulin|sex-binding globulin
C0365086|T201|LC|2942-1|LNC|sex-binding globulin|sex-binding globulin
C0365091|T201|LN|2947-0|LNC|sodium|sodium
C0365091|T201|MTH_LN|2947-0|LNC|sodium|sodium
C0365091|T201|OSN|2947-0|LNC|sodium|sodium
C0365091|T201|LC|2947-0|LNC|sodium|sodium
C0365091|T201|LN|2947-0|LNC|sodium homeostasis|sodium homeostasis
C0365091|T201|MTH_LN|2947-0|LNC|sodium homeostasis|sodium homeostasis
C0365091|T201|OSN|2947-0|LNC|sodium homeostasis|sodium homeostasis
C0365091|T201|LC|2947-0|LNC|sodium homeostasis|sodium homeostasis
C0365095|T201|LN|2951-2|LNC|sodium|sodium
C0365095|T201|MTH_LN|2951-2|LNC|sodium|sodium
C0365095|T201|OSN|2951-2|LNC|sodium|sodium
C0365095|T201|LC|2951-2|LNC|sodium|sodium
C0365095|T201|LN|2951-2|LNC|sodium homeostasis|sodium homeostasis
C0365095|T201|MTH_LN|2951-2|LNC|sodium homeostasis|sodium homeostasis
C0365095|T201|OSN|2951-2|LNC|sodium homeostasis|sodium homeostasis
C0365095|T201|LC|2951-2|LNC|sodium homeostasis|sodium homeostasis
C0365099|T201|LN|2955-3|LNC|sodium|sodium
C0365099|T201|MTH_LN|2955-3|LNC|sodium|sodium
C0365099|T201|OSN|2955-3|LNC|sodium|sodium
C0365099|T201|LC|2955-3|LNC|sodium|sodium
C0365100|T201|LN|2956-1|LNC|sodium|sodium
C0365100|T201|MTH_LN|2956-1|LNC|sodium|sodium
C0365100|T201|OSN|2956-1|LNC|sodium|sodium
C0365100|T201|LC|2956-1|LNC|sodium|sodium
C0365110|T201|LN|2966-0|LNC|osmolality|osmolality
C0365110|T201|MTH_LN|2966-0|LNC|osmolality|osmolality
C0365110|T201|OSN|2966-0|LNC|osmolality|osmolality
C0365110|T201|LC|2966-0|LNC|osmolality|osmolality
C0365110|T201|LN|2966-0|LNC|homeostasis|homeostasis
C0365110|T201|MTH_LN|2966-0|LNC|homeostasis|homeostasis
C0365110|T201|OSN|2966-0|LNC|homeostasis|homeostasis
C0365110|T201|LC|2966-0|LNC|homeostasis|homeostasis
C0365111|T201|MTH_LN|2965-2|LNC|osmolality|osmolality
C0365111|T201|LC|2965-2|LNC|osmolality|osmolality
C0365111|T201|LN|2965-2|LNC|osmolality|osmolality
C0365111|T201|OSN|2965-2|LNC|osmolality|osmolality
C0365111|T201|MTH_LN|2965-2|LNC|homeostasis|homeostasis
C0365111|T201|LC|2965-2|LNC|homeostasis|homeostasis
C0365111|T201|LN|2965-2|LNC|homeostasis|homeostasis
C0365111|T201|OSN|2965-2|LNC|homeostasis|homeostasis
C0365127|T201|LN|2982-7|LNC|taurine|taurine
C0365127|T201|MTH_LN|2982-7|LNC|taurine|taurine
C0365127|T201|OSN|2982-7|LNC|taurine|taurine
C0365127|T201|LC|2982-7|LNC|taurine|taurine
C0365135|T201|LC|2991-8|LNC|testosterone|testosterone
C0365135|T201|MTH_LN|2991-8|LNC|testosterone|testosterone
C0365135|T201|LN|2991-8|LNC|testosterone|testosterone
C0365135|T201|OSN|2991-8|LNC|testosterone|testosterone
C0365137|T201|LC|2986-8|LNC|testosterone|testosterone
C0365137|T201|MTH_LN|2986-8|LNC|testosterone|testosterone
C0365137|T201|LN|2986-8|LNC|testosterone|testosterone
C0365137|T201|OSN|2986-8|LNC|testosterone|testosterone
C0365157|T201|LN|3013-0|LNC|thyroglobulin|thyroglobulin
C0365157|T201|MTH_LN|3013-0|LNC|thyroglobulin|thyroglobulin
C0365157|T201|OSN|3013-0|LNC|thyroglobulin|thyroglobulin
C0365157|T201|LC|3013-0|LNC|thyroglobulin|thyroglobulin
C0365160|T201|LN|3016-3|LNC|thyroid stimulating|thyroid stimulating
C0365160|T201|MTH_LN|3016-3|LNC|thyroid stimulating|thyroid stimulating
C0365160|T201|OSN|3016-3|LNC|thyroid stimulating|thyroid stimulating
C0365160|T201|LC|3016-3|LNC|thyroid stimulating|thyroid stimulating
C0365160|T201|LN|3016-3|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C0365160|T201|MTH_LN|3016-3|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C0365160|T201|OSN|3016-3|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C0365160|T201|LC|3016-3|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C0365160|T201|LN|3016-3|LNC|TSH|TSH
C0365160|T201|MTH_LN|3016-3|LNC|TSH|TSH
C0365160|T201|OSN|3016-3|LNC|TSH|TSH
C0365160|T201|LC|3016-3|LNC|TSH|TSH
C0365160|T201|LN|3016-3|LNC|thyroid-stimulating|thyroid-stimulating
C0365160|T201|MTH_LN|3016-3|LNC|thyroid-stimulating|thyroid-stimulating
C0365160|T201|OSN|3016-3|LNC|thyroid-stimulating|thyroid-stimulating
C0365160|T201|LC|3016-3|LNC|thyroid-stimulating|thyroid-stimulating
C0365168|T201|MTH_LN|3024-7|LNC|thyroxine|thyroxine
C0365168|T201|LN|3024-7|LNC|thyroxine|thyroxine
C0365168|T201|OSN|3024-7|LNC|thyroxine|thyroxine
C0365168|T201|LC|3024-7|LNC|thyroxine|thyroxine
C0365168|T201|MTH_LN|3024-7|LNC|T4|T4
C0365168|T201|LN|3024-7|LNC|T4|T4
C0365168|T201|OSN|3024-7|LNC|T4|T4
C0365168|T201|LC|3024-7|LNC|T4|T4
C0365170|T201|MTH_LN|3026-2|LNC|thyroxine|thyroxine
C0365170|T201|LN|3026-2|LNC|thyroxine|thyroxine
C0365170|T201|OSN|3026-2|LNC|thyroxine|thyroxine
C0365170|T201|LC|3026-2|LNC|thyroxine|thyroxine
C0365170|T201|MTH_LN|3026-2|LNC|T4|T4
C0365170|T201|LN|3026-2|LNC|T4|T4
C0365170|T201|OSN|3026-2|LNC|T4|T4
C0365170|T201|LC|3026-2|LNC|T4|T4
C0365195|T201|MTH_LN|3051-0|LNC|thyroxine|thyroxine
C0365195|T201|LN|3051-0|LNC|thyroxine|thyroxine
C0365195|T201|OSN|3051-0|LNC|thyroxine|thyroxine
C0365195|T201|LC|3051-0|LNC|thyroxine|thyroxine
C0365195|T201|MTH_LN|3051-0|LNC|T4|T4
C0365195|T201|LN|3051-0|LNC|T4|T4
C0365195|T201|OSN|3051-0|LNC|T4|T4
C0365195|T201|LC|3051-0|LNC|T4|T4
C0365213|T201|LN|3069-2|LNC|tryptophan metabolism|tryptophan metabolism
C0365213|T201|MTH_LN|3069-2|LNC|tryptophan metabolism|tryptophan metabolism
C0365213|T201|OSN|3069-2|LNC|tryptophan metabolism|tryptophan metabolism
C0365213|T201|LC|3069-2|LNC|tryptophan metabolism|tryptophan metabolism
C0365223|T201|LN|3079-1|LNC|tyrosine|tyrosine
C0365223|T201|MTH_LN|3079-1|LNC|tyrosine|tyrosine
C0365223|T201|OSN|3079-1|LNC|tyrosine|tyrosine
C0365223|T201|LC|3079-1|LNC|tyrosine|tyrosine
C0365223|T201|LN|3079-1|LNC|tyrosine metabolism|tyrosine metabolism
C0365223|T201|MTH_LN|3079-1|LNC|tyrosine metabolism|tyrosine metabolism
C0365223|T201|OSN|3079-1|LNC|tyrosine metabolism|tyrosine metabolism
C0365223|T201|LC|3079-1|LNC|tyrosine metabolism|tyrosine metabolism
C0365228|T201|LC|3084-1|LNC|uric acid|uric acid
C0365228|T201|MTH_LN|3084-1|LNC|uric acid|uric acid
C0365228|T201|LN|3084-1|LNC|uric acid|uric acid
C0365228|T201|OSN|3084-1|LNC|uric acid|uric acid
C0365228|T201|LC|3084-1|LNC|purine|purine
C0365228|T201|MTH_LN|3084-1|LNC|purine|purine
C0365228|T201|LN|3084-1|LNC|purine|purine
C0365228|T201|OSN|3084-1|LNC|purine|purine
C0365230|T201|LC|3086-6|LNC|urate|urate
C0365230|T201|MTH_LN|3086-6|LNC|urate|urate
C0365230|T201|OSN|3086-6|LNC|urate|urate
C0365230|T201|LN|3086-6|LNC|urate|urate
C0365230|T201|LC|3086-6|LNC|uric acid|uric acid
C0365230|T201|MTH_LN|3086-6|LNC|uric acid|uric acid
C0365230|T201|OSN|3086-6|LNC|uric acid|uric acid
C0365230|T201|LN|3086-6|LNC|uric acid|uric acid
C0365231|T201|LN|3087-4|LNC|urate|urate
C0365231|T201|MTH_LN|3087-4|LNC|urate|urate
C0365231|T201|OSN|3087-4|LNC|urate|urate
C0365231|T201|LC|3087-4|LNC|urate|urate
C0365231|T201|LN|3087-4|LNC|uric acid|uric acid
C0365231|T201|MTH_LN|3087-4|LNC|uric acid|uric acid
C0365231|T201|OSN|3087-4|LNC|uric acid|uric acid
C0365231|T201|LC|3087-4|LNC|uric acid|uric acid
C0365237|T201|LN|6299-2|LNC|BUN|BUN
C0365237|T201|MTH_LN|6299-2|LNC|BUN|BUN
C0365237|T201|OSN|6299-2|LNC|BUN|BUN
C0365237|T201|LC|6299-2|LNC|BUN|BUN
C0365237|T201|LN|6299-2|LNC|urea nitrogen|urea nitrogen
C0365237|T201|MTH_LN|6299-2|LNC|urea nitrogen|urea nitrogen
C0365237|T201|OSN|6299-2|LNC|urea nitrogen|urea nitrogen
C0365237|T201|LC|6299-2|LNC|urea nitrogen|urea nitrogen
C0365240|T201|LC|3094-0|LNC|BUN|BUN
C0365240|T201|MTH_LN|3094-0|LNC|BUN|BUN
C0365240|T201|LN|3094-0|LNC|BUN|BUN
C0365240|T201|OSN|3094-0|LNC|BUN|BUN
C0365240|T201|LC|3094-0|LNC|urea nitrogen|urea nitrogen
C0365240|T201|MTH_LN|3094-0|LNC|urea nitrogen|urea nitrogen
C0365240|T201|LN|3094-0|LNC|urea nitrogen|urea nitrogen
C0365240|T201|OSN|3094-0|LNC|urea nitrogen|urea nitrogen
C0365243|T201|LN|3097-3|LNC|BUN|BUN
C0365243|T201|MTH_LN|3097-3|LNC|BUN|BUN
C0365243|T201|OSN|3097-3|LNC|BUN|BUN
C0365243|T201|LC|3097-3|LNC|BUN|BUN
C0365243|T201|LN|3097-3|LNC|urea nitrogen|urea nitrogen
C0365243|T201|MTH_LN|3097-3|LNC|urea nitrogen|urea nitrogen
C0365243|T201|OSN|3097-3|LNC|urea nitrogen|urea nitrogen
C0365243|T201|LC|3097-3|LNC|urea nitrogen|urea nitrogen
C0365245|T201|LN|3099-9|LNC|uridine diphosphate glucose-4-epimerase activity in|uridine diphosphate glucose-4-epimerase activity in
C0365245|T201|MTH_LN|3099-9|LNC|uridine diphosphate glucose-4-epimerase activity in|uridine diphosphate glucose-4-epimerase activity in
C0365245|T201|OSN|3099-9|LNC|uridine diphosphate glucose-4-epimerase activity in|uridine diphosphate glucose-4-epimerase activity in
C0365245|T201|LC|3099-9|LNC|uridine diphosphate glucose-4-epimerase activity in|uridine diphosphate glucose-4-epimerase activity in
C0365245|T201|LN|3099-9|LNC|UDP-glucose 4-epimerase activity activity in|UDP-glucose 4-epimerase activity activity in
C0365245|T201|MTH_LN|3099-9|LNC|UDP-glucose 4-epimerase activity activity in|UDP-glucose 4-epimerase activity activity in
C0365245|T201|OSN|3099-9|LNC|UDP-glucose 4-epimerase activity activity in|UDP-glucose 4-epimerase activity activity in
C0365245|T201|LC|3099-9|LNC|UDP-glucose 4-epimerase activity activity in|UDP-glucose 4-epimerase activity activity in
C0365253|T201|LC|3107-0|LNC|urobilinogen|urobilinogen
C0365253|T201|MTH_LN|3107-0|LNC|urobilinogen|urobilinogen
C0365253|T201|OSN|3107-0|LNC|urobilinogen|urobilinogen
C0365253|T201|LN|3107-0|LNC|urobilinogen|urobilinogen
C0365254|T201|LN|3108-8|LNC|urobilinogen|urobilinogen
C0365254|T201|MTH_LN|3108-8|LNC|urobilinogen|urobilinogen
C0365254|T201|OSN|3108-8|LNC|urobilinogen|urobilinogen
C0365254|T201|LC|3108-8|LNC|urobilinogen|urobilinogen
C0365255|T201|LN|3109-6|LNC|urobilinogen|urobilinogen
C0365255|T201|MTH_LN|3109-6|LNC|urobilinogen|urobilinogen
C0365255|T201|OSN|3109-6|LNC|urobilinogen|urobilinogen
C0365255|T201|LC|3109-6|LNC|urobilinogen|urobilinogen
C0365282|T201|LN|3137-7|LNC|body height|body height
C0365282|T201|MTH_LN|3137-7|LNC|body height|body height
C0365282|T201|LC|3137-7|LNC|body height|body height
C0365282|T201|OSN|3137-7|LNC|body height|body height
C0365282|T201|LN|3137-7|LNC|linear growth|linear growth
C0365282|T201|MTH_LN|3137-7|LNC|linear growth|linear growth
C0365282|T201|LC|3137-7|LNC|linear growth|linear growth
C0365282|T201|OSN|3137-7|LNC|linear growth|linear growth
C0365286|T201|LN|3141-9|LNC|weight|weight
C0365286|T201|LC|3141-9|LNC|weight|weight
C0365286|T201|OSN|3141-9|LNC|weight|weight
C0365286|T201|MTH_LN|3141-9|LNC|weight|weight
C0365286|T201|LN|3141-9|LNC|body weight|body weight
C0365286|T201|LC|3141-9|LNC|body weight|body weight
C0365286|T201|OSN|3141-9|LNC|body weight|body weight
C0365286|T201|MTH_LN|3141-9|LNC|body weight|body weight
C0365286|T201|LN|3141-9|LNC|habitus|habitus
C0365286|T201|LC|3141-9|LNC|habitus|habitus
C0365286|T201|OSN|3141-9|LNC|habitus|habitus
C0365286|T201|MTH_LN|3141-9|LNC|habitus|habitus
C0365392|T201|LN|3173-2|LNC|coagulation disorder|coagulation disorder
C0365392|T201|MTH_LN|3173-2|LNC|coagulation disorder|coagulation disorder
C0365392|T201|LC|3173-2|LNC|coagulation disorder|coagulation disorder
C0365392|T201|OSN|3173-2|LNC|coagulation disorder|coagulation disorder
C0365392|T201|LN|3173-2|LNC|partial thromboplastin time|partial thromboplastin time
C0365392|T201|MTH_LN|3173-2|LNC|partial thromboplastin time|partial thromboplastin time
C0365392|T201|LC|3173-2|LNC|partial thromboplastin time|partial thromboplastin time
C0365392|T201|OSN|3173-2|LNC|partial thromboplastin time|partial thromboplastin time
C0365392|T201|LN|3173-2|LNC|coagulation|coagulation
C0365392|T201|MTH_LN|3173-2|LNC|coagulation|coagulation
C0365392|T201|LC|3173-2|LNC|coagulation|coagulation
C0365392|T201|OSN|3173-2|LNC|coagulation|coagulation
C0365392|T201|LN|3173-2|LNC|Coagulationities|Coagulationities
C0365392|T201|MTH_LN|3173-2|LNC|Coagulationities|Coagulationities
C0365392|T201|LC|3173-2|LNC|Coagulationities|Coagulationities
C0365392|T201|OSN|3173-2|LNC|Coagulationities|Coagulationities
C0365392|T201|LN|3173-2|LNC|coagulation studies|coagulation studies
C0365392|T201|MTH_LN|3173-2|LNC|coagulation studies|coagulation studies
C0365392|T201|LC|3173-2|LNC|coagulation studies|coagulation studies
C0365392|T201|OSN|3173-2|LNC|coagulation studies|coagulation studies
C0365392|T201|LN|3173-2|LNC|clotting|clotting
C0365392|T201|MTH_LN|3173-2|LNC|clotting|clotting
C0365392|T201|LC|3173-2|LNC|clotting|clotting
C0365392|T201|OSN|3173-2|LNC|clotting|clotting
C0365531|T201|LN|3297-9|LNC|xenobiotic|xenobiotic
C0365531|T201|OSN|3297-9|LNC|xenobiotic|xenobiotic
C0365531|T201|MTH_LN|3297-9|LNC|xenobiotic|xenobiotic
C0365531|T201|LC|3297-9|LNC|xenobiotic|xenobiotic
C0365532|T201|LN|3298-7|LNC|xenobiotic|xenobiotic
C0365532|T201|MTH_LN|3298-7|LNC|xenobiotic|xenobiotic
C0365532|T201|OSN|3298-7|LNC|xenobiotic|xenobiotic
C0365532|T201|LC|3298-7|LNC|xenobiotic|xenobiotic
C0366000|T201|LN|3773-9|LNC|methadone test|methadone test
C0366000|T201|MTH_LN|3773-9|LNC|methadone test|methadone test
C0366000|T201|OSN|3773-9|LNC|methadone test|methadone test
C0366000|T201|LC|3773-9|LNC|methadone test|methadone test
C0366001|T201|LN|3774-7|LNC|methadone test|methadone test
C0366001|T201|MTH_LN|3774-7|LNC|methadone test|methadone test
C0366001|T201|OSN|3774-7|LNC|methadone test|methadone test
C0366001|T201|LC|3774-7|LNC|methadone test|methadone test
C0366002|T201|LN|3775-4|LNC|methadone test|methadone test
C0366002|T201|MTH_LN|3775-4|LNC|methadone test|methadone test
C0366002|T201|OSN|3775-4|LNC|methadone test|methadone test
C0366002|T201|LC|3775-4|LNC|methadone test|methadone test
C0366097|T201|LN|3870-3|LNC|xenobiotic|xenobiotic
C0366097|T201|MTH_LN|3870-3|LNC|xenobiotic|xenobiotic
C0366097|T201|OSN|3870-3|LNC|xenobiotic|xenobiotic
C0366097|T201|LC|3870-3|LNC|xenobiotic|xenobiotic
C0366711|T201|LN|4485-9|LNC|complement C3|complement C3
C0366711|T201|MTH_LN|4485-9|LNC|complement C3|complement C3
C0366711|T201|OSN|4485-9|LNC|complement C3|complement C3
C0366711|T201|LC|4485-9|LNC|complement C3|complement C3
C0366711|T201|LN|4485-9|LNC|C3|C3
C0366711|T201|MTH_LN|4485-9|LNC|C3|C3
C0366711|T201|OSN|4485-9|LNC|C3|C3
C0366711|T201|LC|4485-9|LNC|C3|C3
C0366711|T201|LN|4485-9|LNC|complement system|complement system
C0366711|T201|MTH_LN|4485-9|LNC|complement system|complement system
C0366711|T201|OSN|4485-9|LNC|complement system|complement system
C0366711|T201|LC|4485-9|LNC|complement system|complement system
C0366727|T201|LN|4498-2|LNC|complement system|complement system
C0366727|T201|MTH_LN|4498-2|LNC|complement system|complement system
C0366727|T201|OSN|4498-2|LNC|complement system|complement system
C0366727|T201|LC|4498-2|LNC|complement system|complement system
C0366727|T201|LN|4498-2|LNC|complement C4|complement C4
C0366727|T201|MTH_LN|4498-2|LNC|complement C4|complement C4
C0366727|T201|OSN|4498-2|LNC|complement C4|complement C4
C0366727|T201|LC|4498-2|LNC|complement C4|complement C4
C0366770|T201|LN|4537-7|LNC|erythrocyte|erythrocyte
C0366770|T201|MTH_LN|4537-7|LNC|erythrocyte|erythrocyte
C0366770|T201|OSN|4537-7|LNC|erythrocyte|erythrocyte
C0366770|T201|LC|4537-7|LNC|erythrocyte|erythrocyte
C0366770|T201|LN|4537-7|LNC|ESR|ESR
C0366770|T201|MTH_LN|4537-7|LNC|ESR|ESR
C0366770|T201|OSN|4537-7|LNC|ESR|ESR
C0366770|T201|LC|4537-7|LNC|ESR|ESR
// C0366770|T201|LN|4537-7|LNC||
// C0366770|T201|MTH_LN|4537-7|LNC||
// C0366770|T201|OSN|4537-7|LNC||
// C0366770|T201|LC|4537-7|LNC||
C0366770|T201|LN|4537-7|LNC|Raised erythrocyte|Raised erythrocyte
C0366770|T201|MTH_LN|4537-7|LNC|Raised erythrocyte|Raised erythrocyte
C0366770|T201|OSN|4537-7|LNC|Raised erythrocyte|Raised erythrocyte
C0366770|T201|LC|4537-7|LNC|Raised erythrocyte|Raised erythrocyte
C0366770|T201|LN|4537-7|LNC|Westergren|Westergren
C0366770|T201|MTH_LN|4537-7|LNC|Westergren|Westergren
C0366770|T201|OSN|4537-7|LNC|Westergren|Westergren
C0366770|T201|LC|4537-7|LNC|Westergren|Westergren
C0366777|T201|LN|4544-3|LNC|hematocrit|hematocrit
C0366777|T201|MTH_LN|4544-3|LNC|hematocrit|hematocrit
C0366777|T201|LC|4544-3|LNC|hematocrit|hematocrit
C0366777|T201|OSN|4544-3|LNC|hematocrit|hematocrit
C0366778|T201|LN|4545-0|LNC|hematocrit|hematocrit
C0366778|T201|MTH_LN|4545-0|LNC|hematocrit|hematocrit
C0366778|T201|LC|4545-0|LNC|hematocrit|hematocrit
C0366778|T201|OSN|4545-0|LNC|hematocrit|hematocrit
C0366779|T201|LN|4546-8|LNC|hemoglobin|hemoglobin
C0366779|T201|MTH_LN|4546-8|LNC|hemoglobin|hemoglobin
C0366779|T201|LC|4546-8|LNC|hemoglobin|hemoglobin
C0366779|T201|OSN|4546-8|LNC|hemoglobin|hemoglobin
C0366779|T201|LN|4546-8|LNC|hemoglobin A|hemoglobin A
C0366779|T201|MTH_LN|4546-8|LNC|hemoglobin A|hemoglobin A
C0366779|T201|LC|4546-8|LNC|hemoglobin A|hemoglobin A
C0366779|T201|OSN|4546-8|LNC|hemoglobin A|hemoglobin A
C0366781|T201|LN|4548-4|LNC|hemoglobin|hemoglobin
C0366781|T201|MTH_LN|4548-4|LNC|hemoglobin|hemoglobin
C0366781|T201|OSN|4548-4|LNC|hemoglobin|hemoglobin
C0366781|T201|LC|4548-4|LNC|hemoglobin|hemoglobin
C0366781|T201|LN|4548-4|LNC|hemoglobin A|hemoglobin A
C0366781|T201|MTH_LN|4548-4|LNC|hemoglobin A|hemoglobin A
C0366781|T201|OSN|4548-4|LNC|hemoglobin A|hemoglobin A
C0366781|T201|LC|4548-4|LNC|hemoglobin A|hemoglobin A
C0366781|T201|LN|4548-4|LNC|hemoglobin A1c|hemoglobin A1c
C0366781|T201|MTH_LN|4548-4|LNC|hemoglobin A1c|hemoglobin A1c
C0366781|T201|OSN|4548-4|LNC|hemoglobin A1c|hemoglobin A1c
C0366781|T201|LC|4548-4|LNC|hemoglobin A1c|hemoglobin A1c
C0366781|T201|LN|4548-4|LNC|glycosylated hemoglobin|glycosylated hemoglobin
C0366781|T201|MTH_LN|4548-4|LNC|glycosylated hemoglobin|glycosylated hemoglobin
C0366781|T201|OSN|4548-4|LNC|glycosylated hemoglobin|glycosylated hemoglobin
C0366781|T201|LC|4548-4|LNC|glycosylated hemoglobin|glycosylated hemoglobin
C0366781|T201|LN|4548-4|LNC|HbA1c|HbA1c
C0366781|T201|MTH_LN|4548-4|LNC|HbA1c|HbA1c
C0366781|T201|OSN|4548-4|LNC|HbA1c|HbA1c
C0366781|T201|LC|4548-4|LNC|HbA1c|HbA1c
C0366781|T201|LN|4548-4|LNC|glycated hemoglobin|glycated hemoglobin
C0366781|T201|MTH_LN|4548-4|LNC|glycated hemoglobin|glycated hemoglobin
C0366781|T201|OSN|4548-4|LNC|glycated hemoglobin|glycated hemoglobin
C0366781|T201|LC|4548-4|LNC|glycated hemoglobin|glycated hemoglobin
C0366784|T201|LN|4551-8|LNC|hemoglobin|hemoglobin
C0366784|T201|MTH_LN|4551-8|LNC|hemoglobin|hemoglobin
C0366784|T201|LC|4551-8|LNC|hemoglobin|hemoglobin
C0366784|T201|OSN|4551-8|LNC|hemoglobin|hemoglobin
C0366784|T201|LN|4551-8|LNC|hemoglobin A|hemoglobin A
C0366784|T201|MTH_LN|4551-8|LNC|hemoglobin A|hemoglobin A
C0366784|T201|LC|4551-8|LNC|hemoglobin A|hemoglobin A
C0366784|T201|OSN|4551-8|LNC|hemoglobin A|hemoglobin A
C0366785|T201|LN|4552-6|LNC|hemoglobin|hemoglobin
C0366785|T201|MTH_LN|4552-6|LNC|hemoglobin|hemoglobin
C0366785|T201|LC|4552-6|LNC|hemoglobin|hemoglobin
C0366785|T201|OSN|4552-6|LNC|hemoglobin|hemoglobin
C0366785|T201|LN|4552-6|LNC|hemoglobin A|hemoglobin A
C0366785|T201|MTH_LN|4552-6|LNC|hemoglobin A|hemoglobin A
C0366785|T201|LC|4552-6|LNC|hemoglobin A|hemoglobin A
C0366785|T201|OSN|4552-6|LNC|hemoglobin A|hemoglobin A
C0366869|T201|LN|4636-7|LNC|Hemoglobin|Hemoglobin
C0366869|T201|MTH_LN|4636-7|LNC|Hemoglobin|Hemoglobin
C0366869|T201|OSN|4636-7|LNC|Hemoglobin|Hemoglobin
C0366869|T201|LC|4636-7|LNC|Hemoglobin|Hemoglobin
C0366908|T201|LN|4679-7|LNC|reticulocytes|reticulocytes
C0366908|T201|OSN|4679-7|LNC|reticulocytes|reticulocytes
C0366908|T201|LC|4679-7|LNC|reticulocytes|reticulocytes
C0366908|T201|MTH_LN|4679-7|LNC|reticulocytes|reticulocytes
C0366908|T201|LN|4679-7|LNC|reticulocyte count|reticulocyte count
C0366908|T201|OSN|4679-7|LNC|reticulocyte count|reticulocyte count
C0366908|T201|LC|4679-7|LNC|reticulocyte count|reticulocyte count
C0366908|T201|MTH_LN|4679-7|LNC|reticulocyte count|reticulocyte count
C0367382|T201|LN|5037-7|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367382|T201|MTH_LN|5037-7|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367382|T201|OSN|5037-7|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367382|T201|LC|5037-7|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367383|T201|LN|5038-5|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367383|T201|MTH_LN|5038-5|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367383|T201|OSN|5038-5|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367383|T201|LC|5038-5|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367385|T201|LN|5039-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367385|T201|MTH_LN|5039-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367385|T201|OSN|5039-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367385|T201|LC|5039-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0367570|T201|OLC|5475-9|LNC|T cell CD40 expression|T cell CD40 expression
C0367570|T201|LO|5475-9|LNC|T cell CD40 expression|T cell CD40 expression
C0367570|T201|MTH_LO|5475-9|LNC|T cell CD40 expression|T cell CD40 expression
C0367570|T201|OOSN|5475-9|LNC|T cell CD40 expression|T cell CD40 expression
C0367570|T201|OLC|5475-9|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0367570|T201|LO|5475-9|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0367570|T201|MTH_LO|5475-9|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0367570|T201|OOSN|5475-9|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0367576|T201|OLC|5481-7|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0367576|T201|LO|5481-7|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0367576|T201|MTH_LO|5481-7|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0367576|T201|OOSN|5481-7|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0367576|T201|OLC|5481-7|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0367576|T201|LO|5481-7|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0367576|T201|MTH_LO|5481-7|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0367576|T201|OOSN|5481-7|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0367576|T201|OLC|5481-7|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0367576|T201|LO|5481-7|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0367576|T201|MTH_LO|5481-7|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0367576|T201|OOSN|5481-7|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0367576|T201|OLC|5481-7|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0367576|T201|LO|5481-7|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0367576|T201|MTH_LO|5481-7|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0367576|T201|OOSN|5481-7|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0367788|T201|LN|5631-7|LNC|copper|copper
C0367788|T201|MTH_LN|5631-7|LNC|copper|copper
C0367788|T201|OSN|5631-7|LNC|copper|copper
C0367788|T201|LC|5631-7|LNC|copper|copper
C0367788|T201|LN|5631-7|LNC|copper homeostasis|copper homeostasis
C0367788|T201|MTH_LN|5631-7|LNC|copper homeostasis|copper homeostasis
C0367788|T201|OSN|5631-7|LNC|copper homeostasis|copper homeostasis
C0367788|T201|LC|5631-7|LNC|copper homeostasis|copper homeostasis
C0367790|T201|LN|5633-3|LNC|copper|copper
C0367790|T201|MTH_LN|5633-3|LNC|copper|copper
C0367790|T201|OSN|5633-3|LNC|copper|copper
C0367790|T201|LC|5633-3|LNC|copper|copper
C0367869|T201|LN|5683-8|LNC|magnesium|magnesium
C0367869|T201|MTH_LN|5683-8|LNC|magnesium|magnesium
C0367869|T201|OSN|5683-8|LNC|magnesium|magnesium
C0367869|T201|LC|5683-8|LNC|magnesium|magnesium
C0367869|T201|LN|5683-8|LNC|magnesium metabolism|magnesium metabolism
C0367869|T201|MTH_LN|5683-8|LNC|magnesium metabolism|magnesium metabolism
C0367869|T201|OSN|5683-8|LNC|magnesium metabolism|magnesium metabolism
C0367869|T201|LC|5683-8|LNC|magnesium metabolism|magnesium metabolism
C0367869|T201|LN|5683-8|LNC|magnesium homeostasis|magnesium homeostasis
C0367869|T201|MTH_LN|5683-8|LNC|magnesium homeostasis|magnesium homeostasis
C0367869|T201|OSN|5683-8|LNC|magnesium homeostasis|magnesium homeostasis
C0367869|T201|LC|5683-8|LNC|magnesium homeostasis|magnesium homeostasis
C0367978|T201|LN|5763-8|LNC|zinc|zinc
C0367978|T201|MTH_LN|5763-8|LNC|zinc|zinc
C0367978|T201|OSN|5763-8|LNC|zinc|zinc
C0367978|T201|LC|5763-8|LNC|zinc|zinc
C0367978|T201|LN|5763-8|LNC|zinc metabolism|zinc metabolism
C0367978|T201|MTH_LN|5763-8|LNC|zinc metabolism|zinc metabolism
C0367978|T201|OSN|5763-8|LNC|zinc metabolism|zinc metabolism
C0367978|T201|LC|5763-8|LNC|zinc metabolism|zinc metabolism
C0367978|T201|LN|5763-8|LNC|zinc homeostasis|zinc homeostasis
C0367978|T201|MTH_LN|5763-8|LNC|zinc homeostasis|zinc homeostasis
C0367978|T201|OSN|5763-8|LNC|zinc homeostasis|zinc homeostasis
C0367978|T201|LC|5763-8|LNC|zinc homeostasis|zinc homeostasis
C0367984|T201|LN|5769-5|LNC|bacteria|bacteria
C0367984|T201|MTH_LN|5769-5|LNC|bacteria|bacteria
C0367984|T201|OSN|5769-5|LNC|bacteria|bacteria
C0367984|T201|LC|5769-5|LNC|bacteria|bacteria
C0368002|T201|MTH_LN|5778-6|LNC|Red|Red
C0368002|T201|LC|5778-6|LNC|Red|Red
C0368002|T201|OSN|5778-6|LNC|Red|Red
C0368002|T201|LN|5778-6|LNC|Red|Red
C0368002|T201|MTH_LN|5778-6|LNC|Red-brown|Red-brown
C0368002|T201|LC|5778-6|LNC|Red-brown|Red-brown
C0368002|T201|OSN|5778-6|LNC|Red-brown|Red-brown
C0368002|T201|LN|5778-6|LNC|Red-brown|Red-brown
C0368002|T201|MTH_LN|5778-6|LNC|red brown|red brown
C0368002|T201|LC|5778-6|LNC|red brown|red brown
C0368002|T201|OSN|5778-6|LNC|red brown|red brown
C0368002|T201|LN|5778-6|LNC|red brown|red brown
C0368002|T201|MTH_LN|5778-6|LNC|Purple|Purple
C0368002|T201|LC|5778-6|LNC|Purple|Purple
C0368002|T201|OSN|5778-6|LNC|Purple|Purple
C0368002|T201|LN|5778-6|LNC|Purple|Purple
C0368002|T201|MTH_LN|5778-6|LNC|Blue|Blue
C0368002|T201|LC|5778-6|LNC|Blue|Blue
C0368002|T201|OSN|5778-6|LNC|Blue|Blue
C0368002|T201|LN|5778-6|LNC|Blue|Blue
C0368008|T201|LN|5784-4|LNC|cystine|cystine
C0368008|T201|MTH_LN|5784-4|LNC|cystine|cystine
C0368008|T201|OSN|5784-4|LNC|cystine|cystine
C0368008|T201|LC|5784-4|LNC|cystine|cystine
C0368008|T201|LN|5784-4|LNC|amino acid|amino acid
C0368008|T201|MTH_LN|5784-4|LNC|amino acid|amino acid
C0368008|T201|OSN|5784-4|LNC|amino acid|amino acid
C0368008|T201|LC|5784-4|LNC|amino acid|amino acid
C0368008|T201|LN|5784-4|LNC|animo acids|animo acids
C0368008|T201|MTH_LN|5784-4|LNC|animo acids|animo acids
C0368008|T201|OSN|5784-4|LNC|animo acids|animo acids
C0368008|T201|LC|5784-4|LNC|animo acids|animo acids
C0368008|T201|LN|5784-4|LNC|amino-acid findings|amino-acid findings
C0368008|T201|MTH_LN|5784-4|LNC|amino-acid findings|amino-acid findings
C0368008|T201|OSN|5784-4|LNC|amino-acid findings|amino-acid findings
C0368008|T201|LC|5784-4|LNC|amino-acid findings|amino-acid findings
C0368018|T201|LN|5792-7|LNC|glucose|glucose
C0368018|T201|MTH_LN|5792-7|LNC|glucose|glucose
C0368018|T201|OSN|5792-7|LNC|glucose|glucose
C0368018|T201|LC|5792-7|LNC|glucose|glucose
C0368020|T201|LN|5794-3|LNC|Hemoglobin|Hemoglobin
C0368020|T201|MTH_LN|5794-3|LNC|Hemoglobin|Hemoglobin
C0368020|T201|OSN|5794-3|LNC|Hemoglobin|Hemoglobin
C0368020|T201|LC|5794-3|LNC|Hemoglobin|Hemoglobin
C0368036|T201|LN|5821-4|LNC|neutrophil count|neutrophil count
C0368036|T201|MTH_LN|5821-4|LNC|neutrophil count|neutrophil count
C0368036|T201|LC|5821-4|LNC|neutrophil count|neutrophil count
C0368036|T201|OSN|5821-4|LNC|neutrophil count|neutrophil count
C0368036|T201|LN|5821-4|LNC|cytology|cytology
C0368036|T201|MTH_LN|5821-4|LNC|cytology|cytology
C0368036|T201|LC|5821-4|LNC|cytology|cytology
C0368036|T201|OSN|5821-4|LNC|cytology|cytology
C0368042|T201|LN|5803-2|LNC|acid-base homeostasis|acid-base homeostasis
C0368042|T201|MTH_LN|5803-2|LNC|acid-base homeostasis|acid-base homeostasis
C0368042|T201|OSN|5803-2|LNC|acid-base homeostasis|acid-base homeostasis
C0368042|T201|LC|5803-2|LNC|acid-base homeostasis|acid-base homeostasis
C0368043|T201|LN|5804-0|LNC|Protein|Protein
C0368043|T201|MTH_LN|5804-0|LNC|Protein|Protein
C0368043|T201|OSN|5804-0|LNC|Protein|Protein
C0368043|T201|LC|5804-0|LNC|Protein|Protein
C0368059|T201|LN|5810-7|LNC|osmolality|osmolality
C0368059|T201|MTH_LN|5810-7|LNC|osmolality|osmolality
C0368059|T201|LC|5810-7|LNC|osmolality|osmolality
C0368059|T201|OSN|5810-7|LNC|osmolality|osmolality
C0368059|T201|LN|5810-7|LNC|homeostasis|homeostasis
C0368059|T201|MTH_LN|5810-7|LNC|homeostasis|homeostasis
C0368059|T201|LC|5810-7|LNC|homeostasis|homeostasis
C0368059|T201|OSN|5810-7|LNC|homeostasis|homeostasis
C0368061|T201|LN|5811-5|LNC|osmolality|osmolality
C0368061|T201|MTH_LN|5811-5|LNC|osmolality|osmolality
C0368061|T201|LC|5811-5|LNC|osmolality|osmolality
C0368061|T201|OSN|5811-5|LNC|osmolality|osmolality
C0368061|T201|LN|5811-5|LNC|homeostasis|homeostasis
C0368061|T201|MTH_LN|5811-5|LNC|homeostasis|homeostasis
C0368061|T201|LC|5811-5|LNC|homeostasis|homeostasis
C0368061|T201|OSN|5811-5|LNC|homeostasis|homeostasis
C0368078|T201|LN|5818-0|LNC|urobilinogen|urobilinogen
C0368078|T201|MTH_LN|5818-0|LNC|urobilinogen|urobilinogen
C0368078|T201|OSN|5818-0|LNC|urobilinogen|urobilinogen
C0368078|T201|LC|5818-0|LNC|urobilinogen|urobilinogen
C0368563|T201|LN|630-4|LNC|bacteria|bacteria
C0368563|T201|MTH_LN|630-4|LNC|bacteria|bacteria
C0368563|T201|OSN|630-4|LNC|bacteria|bacteria
C0368563|T201|LC|630-4|LNC|bacteria|bacteria
C0425373|T098|LN|2075-0|LNC|chloride|chloride
C0425373|T098|MTH_LN|2075-0|LNC|chloride|chloride
C0425373|T098|OSN|2075-0|LNC|chloride|chloride
C0425373|T098|LC|2075-0|LNC|chloride|chloride
C0425373|T098|LN|2075-0|LNC|chloride homeostasis|chloride homeostasis
C0425373|T098|MTH_LN|2075-0|LNC|chloride homeostasis|chloride homeostasis
C0425373|T098|OSN|2075-0|LNC|chloride homeostasis|chloride homeostasis
C0425373|T098|LC|2075-0|LNC|chloride homeostasis|chloride homeostasis
C0482460|T201|LN|1359-9|LNC|adrenocorticotropin|adrenocorticotropin
C0482460|T201|MTH_LN|1359-9|LNC|adrenocorticotropin|adrenocorticotropin
C0482460|T201|OSN|1359-9|LNC|adrenocorticotropin|adrenocorticotropin
C0482460|T201|LC|1359-9|LNC|adrenocorticotropin|adrenocorticotropin
C0482460|T201|LN|1359-9|LNC|ACTH|ACTH
C0482460|T201|MTH_LN|1359-9|LNC|ACTH|ACTH
C0482460|T201|OSN|1359-9|LNC|ACTH|ACTH
C0482460|T201|LC|1359-9|LNC|ACTH|ACTH
C0482461|T201|LN|1361-5|LNC|adrenocorticotropin|adrenocorticotropin
C0482461|T201|MTH_LN|1361-5|LNC|adrenocorticotropin|adrenocorticotropin
C0482461|T201|OSN|1361-5|LNC|adrenocorticotropin|adrenocorticotropin
C0482461|T201|LC|1361-5|LNC|adrenocorticotropin|adrenocorticotropin
C0482461|T201|LN|1361-5|LNC|ACTH|ACTH
C0482461|T201|MTH_LN|1361-5|LNC|ACTH|ACTH
C0482461|T201|OSN|1361-5|LNC|ACTH|ACTH
C0482461|T201|LC|1361-5|LNC|ACTH|ACTH
C0482462|T201|LN|1362-3|LNC|adrenocorticotropin|adrenocorticotropin
C0482462|T201|MTH_LN|1362-3|LNC|adrenocorticotropin|adrenocorticotropin
C0482462|T201|OSN|1362-3|LNC|adrenocorticotropin|adrenocorticotropin
C0482462|T201|LC|1362-3|LNC|adrenocorticotropin|adrenocorticotropin
C0482462|T201|LN|1362-3|LNC|ACTH|ACTH
C0482462|T201|MTH_LN|1362-3|LNC|ACTH|ACTH
C0482462|T201|OSN|1362-3|LNC|ACTH|ACTH
C0482462|T201|LC|1362-3|LNC|ACTH|ACTH
C0482463|T201|LN|1364-9|LNC|adrenocorticotropin|adrenocorticotropin
C0482463|T201|MTH_LN|1364-9|LNC|adrenocorticotropin|adrenocorticotropin
C0482463|T201|OSN|1364-9|LNC|adrenocorticotropin|adrenocorticotropin
C0482463|T201|LC|1364-9|LNC|adrenocorticotropin|adrenocorticotropin
C0482463|T201|LN|1364-9|LNC|ACTH|ACTH
C0482463|T201|MTH_LN|1364-9|LNC|ACTH|ACTH
C0482463|T201|OSN|1364-9|LNC|ACTH|ACTH
C0482463|T201|LC|1364-9|LNC|ACTH|ACTH
C0482464|T201|LN|1366-4|LNC|adrenocorticotropin|adrenocorticotropin
C0482464|T201|MTH_LN|1366-4|LNC|adrenocorticotropin|adrenocorticotropin
C0482464|T201|OSN|1366-4|LNC|adrenocorticotropin|adrenocorticotropin
C0482464|T201|LC|1366-4|LNC|adrenocorticotropin|adrenocorticotropin
C0482464|T201|LN|1366-4|LNC|ACTH|ACTH
C0482464|T201|MTH_LN|1366-4|LNC|ACTH|ACTH
C0482464|T201|OSN|1366-4|LNC|ACTH|ACTH
C0482464|T201|LC|1366-4|LNC|ACTH|ACTH
C0482465|T201|LN|1367-2|LNC|adrenocorticotropin|adrenocorticotropin
C0482465|T201|MTH_LN|1367-2|LNC|adrenocorticotropin|adrenocorticotropin
C0482465|T201|OSN|1367-2|LNC|adrenocorticotropin|adrenocorticotropin
C0482465|T201|LC|1367-2|LNC|adrenocorticotropin|adrenocorticotropin
C0482465|T201|LN|1367-2|LNC|ACTH|ACTH
C0482465|T201|MTH_LN|1367-2|LNC|ACTH|ACTH
C0482465|T201|OSN|1367-2|LNC|ACTH|ACTH
C0482465|T201|LC|1367-2|LNC|ACTH|ACTH
C0482466|T201|LN|1368-0|LNC|adrenocorticotropin|adrenocorticotropin
C0482466|T201|MTH_LN|1368-0|LNC|adrenocorticotropin|adrenocorticotropin
C0482466|T201|OSN|1368-0|LNC|adrenocorticotropin|adrenocorticotropin
C0482466|T201|LC|1368-0|LNC|adrenocorticotropin|adrenocorticotropin
C0482466|T201|LN|1368-0|LNC|ACTH|ACTH
C0482466|T201|MTH_LN|1368-0|LNC|ACTH|ACTH
C0482466|T201|OSN|1368-0|LNC|ACTH|ACTH
C0482466|T201|LC|1368-0|LNC|ACTH|ACTH
C0482477|T201|LN|1389-6|LNC|cortisol|cortisol
C0482477|T201|MTH_LN|1389-6|LNC|cortisol|cortisol
C0482477|T201|OSN|1389-6|LNC|cortisol|cortisol
C0482477|T201|LC|1389-6|LNC|cortisol|cortisol
// C0482477|T201|LN|1389-6|LNC||
// C0482477|T201|MTH_LN|1389-6|LNC||
// C0482477|T201|OSN|1389-6|LNC||
// C0482477|T201|LC|1389-6|LNC||
C0482478|T201|LN|1390-4|LNC|cortisol|cortisol
C0482478|T201|MTH_LN|1390-4|LNC|cortisol|cortisol
C0482478|T201|OSN|1390-4|LNC|cortisol|cortisol
C0482478|T201|LC|1390-4|LNC|cortisol|cortisol
// C0482478|T201|LN|1390-4|LNC||
// C0482478|T201|MTH_LN|1390-4|LNC||
// C0482478|T201|OSN|1390-4|LNC||
// C0482478|T201|LC|1390-4|LNC||
C0482480|T201|LN|1393-8|LNC|cortisol|cortisol
C0482480|T201|MTH_LN|1393-8|LNC|cortisol|cortisol
C0482480|T201|OSN|1393-8|LNC|cortisol|cortisol
C0482480|T201|LC|1393-8|LNC|cortisol|cortisol
// C0482480|T201|LN|1393-8|LNC||
// C0482480|T201|MTH_LN|1393-8|LNC||
// C0482480|T201|OSN|1393-8|LNC||
// C0482480|T201|LC|1393-8|LNC||
C0482481|T201|LN|1394-6|LNC|cortisol|cortisol
C0482481|T201|MTH_LN|1394-6|LNC|cortisol|cortisol
C0482481|T201|OSN|1394-6|LNC|cortisol|cortisol
C0482481|T201|LC|1394-6|LNC|cortisol|cortisol
// C0482481|T201|LN|1394-6|LNC||
// C0482481|T201|MTH_LN|1394-6|LNC||
// C0482481|T201|OSN|1394-6|LNC||
// C0482481|T201|LC|1394-6|LNC||
C0482485|T201|LN|1401-9|LNC|cortisol|cortisol
C0482485|T201|MTH_LN|1401-9|LNC|cortisol|cortisol
C0482485|T201|OSN|1401-9|LNC|cortisol|cortisol
C0482485|T201|LC|1401-9|LNC|cortisol|cortisol
C0482485|T201|LN|1401-9|LNC|cortisol low|cortisol low
C0482485|T201|MTH_LN|1401-9|LNC|cortisol low|cortisol low
C0482485|T201|OSN|1401-9|LNC|cortisol low|cortisol low
C0482485|T201|LC|1401-9|LNC|cortisol low|cortisol low
C0482485|T201|LN|1401-9|LNC|to undetectable cortisol|to undetectable cortisol
C0482485|T201|MTH_LN|1401-9|LNC|to undetectable cortisol|to undetectable cortisol
C0482485|T201|OSN|1401-9|LNC|to undetectable cortisol|to undetectable cortisol
C0482485|T201|LC|1401-9|LNC|to undetectable cortisol|to undetectable cortisol
C0482486|T201|LN|1402-7|LNC|cortisol|cortisol
C0482486|T201|MTH_LN|1402-7|LNC|cortisol|cortisol
C0482486|T201|OSN|1402-7|LNC|cortisol|cortisol
C0482486|T201|LC|1402-7|LNC|cortisol|cortisol
C0482486|T201|LN|1402-7|LNC|cortisol low|cortisol low
C0482486|T201|MTH_LN|1402-7|LNC|cortisol low|cortisol low
C0482486|T201|OSN|1402-7|LNC|cortisol low|cortisol low
C0482486|T201|LC|1402-7|LNC|cortisol low|cortisol low
C0482486|T201|LN|1402-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482486|T201|MTH_LN|1402-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482486|T201|OSN|1402-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482486|T201|LC|1402-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482487|T201|LN|1403-5|LNC|cortisol|cortisol
C0482487|T201|MTH_LN|1403-5|LNC|cortisol|cortisol
C0482487|T201|OSN|1403-5|LNC|cortisol|cortisol
C0482487|T201|LC|1403-5|LNC|cortisol|cortisol
C0482487|T201|LN|1403-5|LNC|cortisol low|cortisol low
C0482487|T201|MTH_LN|1403-5|LNC|cortisol low|cortisol low
C0482487|T201|OSN|1403-5|LNC|cortisol low|cortisol low
C0482487|T201|LC|1403-5|LNC|cortisol low|cortisol low
C0482487|T201|LN|1403-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482487|T201|MTH_LN|1403-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482487|T201|OSN|1403-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482487|T201|LC|1403-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482489|T201|LN|1408-4|LNC|cortisol|cortisol
C0482489|T201|MTH_LN|1408-4|LNC|cortisol|cortisol
C0482489|T201|OSN|1408-4|LNC|cortisol|cortisol
C0482489|T201|LC|1408-4|LNC|cortisol|cortisol
C0482489|T201|LN|1408-4|LNC|cortisol low|cortisol low
C0482489|T201|MTH_LN|1408-4|LNC|cortisol low|cortisol low
C0482489|T201|OSN|1408-4|LNC|cortisol low|cortisol low
C0482489|T201|LC|1408-4|LNC|cortisol low|cortisol low
C0482489|T201|LN|1408-4|LNC|to undetectable cortisol|to undetectable cortisol
C0482489|T201|MTH_LN|1408-4|LNC|to undetectable cortisol|to undetectable cortisol
C0482489|T201|OSN|1408-4|LNC|to undetectable cortisol|to undetectable cortisol
C0482489|T201|LC|1408-4|LNC|to undetectable cortisol|to undetectable cortisol
C0482490|T201|LN|1409-2|LNC|cortisol|cortisol
C0482490|T201|MTH_LN|1409-2|LNC|cortisol|cortisol
C0482490|T201|OSN|1409-2|LNC|cortisol|cortisol
C0482490|T201|LC|1409-2|LNC|cortisol|cortisol
C0482490|T201|LN|1409-2|LNC|cortisol low|cortisol low
C0482490|T201|MTH_LN|1409-2|LNC|cortisol low|cortisol low
C0482490|T201|OSN|1409-2|LNC|cortisol low|cortisol low
C0482490|T201|LC|1409-2|LNC|cortisol low|cortisol low
C0482490|T201|LN|1409-2|LNC|to undetectable cortisol|to undetectable cortisol
C0482490|T201|MTH_LN|1409-2|LNC|to undetectable cortisol|to undetectable cortisol
C0482490|T201|OSN|1409-2|LNC|to undetectable cortisol|to undetectable cortisol
C0482490|T201|LC|1409-2|LNC|to undetectable cortisol|to undetectable cortisol
C0482493|T201|LN|1413-4|LNC|cortisol|cortisol
C0482493|T201|MTH_LN|1413-4|LNC|cortisol|cortisol
C0482493|T201|OSN|1413-4|LNC|cortisol|cortisol
C0482493|T201|LC|1413-4|LNC|cortisol|cortisol
C0482493|T201|LN|1413-4|LNC|cortisol low|cortisol low
C0482493|T201|MTH_LN|1413-4|LNC|cortisol low|cortisol low
C0482493|T201|OSN|1413-4|LNC|cortisol low|cortisol low
C0482493|T201|LC|1413-4|LNC|cortisol low|cortisol low
C0482493|T201|LN|1413-4|LNC|to undetectable cortisol|to undetectable cortisol
C0482493|T201|MTH_LN|1413-4|LNC|to undetectable cortisol|to undetectable cortisol
C0482493|T201|OSN|1413-4|LNC|to undetectable cortisol|to undetectable cortisol
C0482493|T201|LC|1413-4|LNC|to undetectable cortisol|to undetectable cortisol
C0482495|T201|LN|1416-7|LNC|cortisol|cortisol
C0482495|T201|MTH_LN|1416-7|LNC|cortisol|cortisol
C0482495|T201|OSN|1416-7|LNC|cortisol|cortisol
C0482495|T201|LC|1416-7|LNC|cortisol|cortisol
C0482495|T201|LN|1416-7|LNC|cortisol low|cortisol low
C0482495|T201|MTH_LN|1416-7|LNC|cortisol low|cortisol low
C0482495|T201|OSN|1416-7|LNC|cortisol low|cortisol low
C0482495|T201|LC|1416-7|LNC|cortisol low|cortisol low
C0482495|T201|LN|1416-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482495|T201|MTH_LN|1416-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482495|T201|OSN|1416-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482495|T201|LC|1416-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482496|T201|LN|1417-5|LNC|cortisol|cortisol
C0482496|T201|MTH_LN|1417-5|LNC|cortisol|cortisol
C0482496|T201|OSN|1417-5|LNC|cortisol|cortisol
C0482496|T201|LC|1417-5|LNC|cortisol|cortisol
C0482496|T201|LN|1417-5|LNC|cortisol low|cortisol low
C0482496|T201|MTH_LN|1417-5|LNC|cortisol low|cortisol low
C0482496|T201|OSN|1417-5|LNC|cortisol low|cortisol low
C0482496|T201|LC|1417-5|LNC|cortisol low|cortisol low
C0482496|T201|LN|1417-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482496|T201|MTH_LN|1417-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482496|T201|OSN|1417-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482496|T201|LC|1417-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482497|T201|LN|1418-3|LNC|cortisol|cortisol
C0482497|T201|MTH_LN|1418-3|LNC|cortisol|cortisol
C0482497|T201|OSN|1418-3|LNC|cortisol|cortisol
C0482497|T201|LC|1418-3|LNC|cortisol|cortisol
C0482497|T201|LN|1418-3|LNC|cortisol low|cortisol low
C0482497|T201|MTH_LN|1418-3|LNC|cortisol low|cortisol low
C0482497|T201|OSN|1418-3|LNC|cortisol low|cortisol low
C0482497|T201|LC|1418-3|LNC|cortisol low|cortisol low
C0482497|T201|LN|1418-3|LNC|to undetectable cortisol|to undetectable cortisol
C0482497|T201|MTH_LN|1418-3|LNC|to undetectable cortisol|to undetectable cortisol
C0482497|T201|OSN|1418-3|LNC|to undetectable cortisol|to undetectable cortisol
C0482497|T201|LC|1418-3|LNC|to undetectable cortisol|to undetectable cortisol
C0482498|T201|LN|1421-7|LNC|cortisol|cortisol
C0482498|T201|MTH_LN|1421-7|LNC|cortisol|cortisol
C0482498|T201|OSN|1421-7|LNC|cortisol|cortisol
C0482498|T201|LC|1421-7|LNC|cortisol|cortisol
C0482498|T201|LN|1421-7|LNC|cortisol low|cortisol low
C0482498|T201|MTH_LN|1421-7|LNC|cortisol low|cortisol low
C0482498|T201|OSN|1421-7|LNC|cortisol low|cortisol low
C0482498|T201|LC|1421-7|LNC|cortisol low|cortisol low
C0482498|T201|LN|1421-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482498|T201|MTH_LN|1421-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482498|T201|OSN|1421-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482498|T201|LC|1421-7|LNC|to undetectable cortisol|to undetectable cortisol
C0482499|T201|LN|1422-5|LNC|cortisol|cortisol
C0482499|T201|MTH_LN|1422-5|LNC|cortisol|cortisol
C0482499|T201|OSN|1422-5|LNC|cortisol|cortisol
C0482499|T201|LC|1422-5|LNC|cortisol|cortisol
C0482499|T201|LN|1422-5|LNC|cortisol low|cortisol low
C0482499|T201|MTH_LN|1422-5|LNC|cortisol low|cortisol low
C0482499|T201|OSN|1422-5|LNC|cortisol low|cortisol low
C0482499|T201|LC|1422-5|LNC|cortisol low|cortisol low
C0482499|T201|LN|1422-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482499|T201|MTH_LN|1422-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482499|T201|OSN|1422-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482499|T201|LC|1422-5|LNC|to undetectable cortisol|to undetectable cortisol
C0482501|T201|LN|1426-6|LNC|cortisol|cortisol
C0482501|T201|MTH_LN|1426-6|LNC|cortisol|cortisol
C0482501|T201|OSN|1426-6|LNC|cortisol|cortisol
C0482501|T201|LC|1426-6|LNC|cortisol|cortisol
C0482501|T201|LN|1426-6|LNC|cortisol low|cortisol low
C0482501|T201|MTH_LN|1426-6|LNC|cortisol low|cortisol low
C0482501|T201|OSN|1426-6|LNC|cortisol low|cortisol low
C0482501|T201|LC|1426-6|LNC|cortisol low|cortisol low
C0482501|T201|LN|1426-6|LNC|to undetectable cortisol|to undetectable cortisol
C0482501|T201|MTH_LN|1426-6|LNC|to undetectable cortisol|to undetectable cortisol
C0482501|T201|OSN|1426-6|LNC|to undetectable cortisol|to undetectable cortisol
C0482501|T201|LC|1426-6|LNC|to undetectable cortisol|to undetectable cortisol
C0482504|T201|LN|1430-8|LNC|cortisol|cortisol
C0482504|T201|MTH_LN|1430-8|LNC|cortisol|cortisol
C0482504|T201|OSN|1430-8|LNC|cortisol|cortisol
C0482504|T201|LC|1430-8|LNC|cortisol|cortisol
C0482504|T201|LN|1430-8|LNC|cortisol low|cortisol low
C0482504|T201|MTH_LN|1430-8|LNC|cortisol low|cortisol low
C0482504|T201|OSN|1430-8|LNC|cortisol low|cortisol low
C0482504|T201|LC|1430-8|LNC|cortisol low|cortisol low
C0482504|T201|LN|1430-8|LNC|to undetectable cortisol|to undetectable cortisol
C0482504|T201|MTH_LN|1430-8|LNC|to undetectable cortisol|to undetectable cortisol
C0482504|T201|OSN|1430-8|LNC|to undetectable cortisol|to undetectable cortisol
C0482504|T201|LC|1430-8|LNC|to undetectable cortisol|to undetectable cortisol
C0482508|T201|LN|1438-1|LNC|cortisol|cortisol
C0482508|T201|MTH_LN|1438-1|LNC|cortisol|cortisol
C0482508|T201|OSN|1438-1|LNC|cortisol|cortisol
C0482508|T201|LC|1438-1|LNC|cortisol|cortisol
C0482508|T201|LN|1438-1|LNC|cortisol low|cortisol low
C0482508|T201|MTH_LN|1438-1|LNC|cortisol low|cortisol low
C0482508|T201|OSN|1438-1|LNC|cortisol low|cortisol low
C0482508|T201|LC|1438-1|LNC|cortisol low|cortisol low
C0482508|T201|LN|1438-1|LNC|to undetectable cortisol|to undetectable cortisol
C0482508|T201|MTH_LN|1438-1|LNC|to undetectable cortisol|to undetectable cortisol
C0482508|T201|OSN|1438-1|LNC|to undetectable cortisol|to undetectable cortisol
C0482508|T201|LC|1438-1|LNC|to undetectable cortisol|to undetectable cortisol
C0482513|T201|LN|1447-2|LNC|cortisol|cortisol
C0482513|T201|MTH_LN|1447-2|LNC|cortisol|cortisol
C0482513|T201|OSN|1447-2|LNC|cortisol|cortisol
C0482513|T201|LC|1447-2|LNC|cortisol|cortisol
C0482513|T201|LN|1447-2|LNC|cortisol low|cortisol low
C0482513|T201|MTH_LN|1447-2|LNC|cortisol low|cortisol low
C0482513|T201|OSN|1447-2|LNC|cortisol low|cortisol low
C0482513|T201|LC|1447-2|LNC|cortisol low|cortisol low
C0482513|T201|LN|1447-2|LNC|to undetectable cortisol|to undetectable cortisol
C0482513|T201|MTH_LN|1447-2|LNC|to undetectable cortisol|to undetectable cortisol
C0482513|T201|OSN|1447-2|LNC|to undetectable cortisol|to undetectable cortisol
C0482513|T201|LC|1447-2|LNC|to undetectable cortisol|to undetectable cortisol
C0482534|T201|LN|1496-9|LNC|glucose|glucose
C0482534|T201|OSN|1496-9|LNC|glucose|glucose
C0482534|T201|MTH_LN|1496-9|LNC|glucose|glucose
C0482534|T201|LC|1496-9|LNC|glucose|glucose
C0482535|T201|LN|1521-4|LNC|glucose|glucose
C0482535|T201|MTH_LN|1521-4|LNC|glucose|glucose
C0482535|T201|OSN|1521-4|LNC|glucose|glucose
C0482535|T201|LC|1521-4|LNC|glucose|glucose
C0482536|T201|LN|1524-8|LNC|glucose|glucose
C0482536|T201|MTH_LN|1524-8|LNC|glucose|glucose
C0482536|T201|OSN|1524-8|LNC|glucose|glucose
C0482536|T201|LC|1524-8|LNC|glucose|glucose
C0482537|T201|LN|1527-1|LNC|glucose|glucose
C0482537|T201|MTH_LN|1527-1|LNC|glucose|glucose
C0482537|T201|OSN|1527-1|LNC|glucose|glucose
C0482537|T201|LC|1527-1|LNC|glucose|glucose
C0482538|T201|LN|1548-7|LNC|glucose|glucose
C0482538|T201|MTH_LN|1548-7|LNC|glucose|glucose
C0482538|T201|OSN|1548-7|LNC|glucose|glucose
C0482538|T201|LC|1548-7|LNC|glucose|glucose
C0482539|T201|LN|1549-5|LNC|glucose|glucose
C0482539|T201|MTH_LN|1549-5|LNC|glucose|glucose
C0482539|T201|OSN|1549-5|LNC|glucose|glucose
C0482539|T201|LC|1549-5|LNC|glucose|glucose
C0482540|T201|LN|1550-3|LNC|glucose|glucose
C0482540|T201|MTH_LN|1550-3|LNC|glucose|glucose
C0482540|T201|OSN|1550-3|LNC|glucose|glucose
C0482540|T201|LC|1550-3|LNC|glucose|glucose
C0482541|T201|LN|1551-1|LNC|glucose|glucose
C0482541|T201|MTH_LN|1551-1|LNC|glucose|glucose
C0482541|T201|OSN|1551-1|LNC|glucose|glucose
C0482541|T201|LC|1551-1|LNC|glucose|glucose
C0482542|T201|LN|1552-9|LNC|glucose|glucose
C0482542|T201|MTH_LN|1552-9|LNC|glucose|glucose
C0482542|T201|OSN|1552-9|LNC|glucose|glucose
C0482542|T201|LC|1552-9|LNC|glucose|glucose
C0482543|T201|LN|1553-7|LNC|glucose|glucose
C0482543|T201|MTH_LN|1553-7|LNC|glucose|glucose
C0482543|T201|OSN|1553-7|LNC|glucose|glucose
C0482543|T201|LC|1553-7|LNC|glucose|glucose
C0482544|T201|MTH_LN|1558-6|LNC|glucose|glucose
C0482544|T201|LN|1558-6|LNC|glucose|glucose
C0482544|T201|OSN|1558-6|LNC|glucose|glucose
C0482544|T201|LC|1558-6|LNC|glucose|glucose
C0482562|T201|LN|1600-6|LNC|luteinizing|luteinizing
C0482562|T201|MTH_LN|1600-6|LNC|luteinizing|luteinizing
C0482562|T201|OSN|1600-6|LNC|luteinizing|luteinizing
C0482562|T201|LC|1600-6|LNC|luteinizing|luteinizing
C0482562|T201|LN|1600-6|LNC|LH|LH
C0482562|T201|MTH_LN|1600-6|LNC|LH|LH
C0482562|T201|OSN|1600-6|LNC|LH|LH
C0482562|T201|LC|1600-6|LNC|LH|LH
C0482562|T201|LN|1600-6|LNC|luteinising|luteinising
C0482562|T201|MTH_LN|1600-6|LNC|luteinising|luteinising
C0482562|T201|OSN|1600-6|LNC|luteinising|luteinising
C0482562|T201|LC|1600-6|LNC|luteinising|luteinising
C0482602|T201|LN|2842-3|LNC|prolactin|prolactin
C0482602|T201|MTH_LN|2842-3|LNC|prolactin|prolactin
C0482602|T201|OSN|2842-3|LNC|prolactin|prolactin
C0482602|T201|LC|2842-3|LNC|prolactin|prolactin
C0482617|T201|LN|3193-0|LNC|coagulation factor V activity|coagulation factor V activity
C0482617|T201|MTH_LN|3193-0|LNC|coagulation factor V activity|coagulation factor V activity
C0482617|T201|OSN|3193-0|LNC|coagulation factor V activity|coagulation factor V activity
C0482617|T201|LC|3193-0|LNC|coagulation factor V activity|coagulation factor V activity
C0482617|T201|LN|3193-0|LNC|factor V activity|factor V activity
C0482617|T201|MTH_LN|3193-0|LNC|factor V activity|factor V activity
C0482617|T201|OSN|3193-0|LNC|factor V activity|factor V activity
C0482617|T201|LC|3193-0|LNC|factor V activity|factor V activity
C0482617|T201|LN|3193-0|LNC|factor V|factor V
C0482617|T201|MTH_LN|3193-0|LNC|factor V|factor V
C0482617|T201|OSN|3193-0|LNC|factor V|factor V
C0482617|T201|LC|3193-0|LNC|factor V|factor V
C0482633|T201|LN|3209-4|LNC|factor VIII activity|factor VIII activity
C0482633|T201|MTH_LN|3209-4|LNC|factor VIII activity|factor VIII activity
C0482633|T201|OSN|3209-4|LNC|factor VIII activity|factor VIII activity
C0482633|T201|LC|3209-4|LNC|factor VIII activity|factor VIII activity
C0482677|T201|MTH_LN|5946-9|LNC|coagulation disorder|coagulation disorder
C0482677|T201|LC|5946-9|LNC|coagulation disorder|coagulation disorder
C0482677|T201|LN|5946-9|LNC|coagulation disorder|coagulation disorder
C0482677|T201|OSN|5946-9|LNC|coagulation disorder|coagulation disorder
C0482677|T201|MTH_LN|5946-9|LNC|partial thromboplastin time|partial thromboplastin time
C0482677|T201|LC|5946-9|LNC|partial thromboplastin time|partial thromboplastin time
C0482677|T201|LN|5946-9|LNC|partial thromboplastin time|partial thromboplastin time
C0482677|T201|OSN|5946-9|LNC|partial thromboplastin time|partial thromboplastin time
C0482677|T201|MTH_LN|5946-9|LNC|coagulation|coagulation
C0482677|T201|LC|5946-9|LNC|coagulation|coagulation
C0482677|T201|LN|5946-9|LNC|coagulation|coagulation
C0482677|T201|OSN|5946-9|LNC|coagulation|coagulation
C0482677|T201|MTH_LN|5946-9|LNC|Coagulationities|Coagulationities
C0482677|T201|LC|5946-9|LNC|Coagulationities|Coagulationities
C0482677|T201|LN|5946-9|LNC|Coagulationities|Coagulationities
C0482677|T201|OSN|5946-9|LNC|Coagulationities|Coagulationities
C0482677|T201|MTH_LN|5946-9|LNC|coagulation studies|coagulation studies
C0482677|T201|LC|5946-9|LNC|coagulation studies|coagulation studies
C0482677|T201|LN|5946-9|LNC|coagulation studies|coagulation studies
C0482677|T201|OSN|5946-9|LNC|coagulation studies|coagulation studies
C0482677|T201|MTH_LN|5946-9|LNC|clotting|clotting
C0482677|T201|LC|5946-9|LNC|clotting|clotting
C0482677|T201|LN|5946-9|LNC|clotting|clotting
C0482677|T201|OSN|5946-9|LNC|clotting|clotting
C0482705|T201|MTH_LN|3255-7|LNC|fibrinogen|fibrinogen
C0482705|T201|LN|3255-7|LNC|fibrinogen|fibrinogen
C0482705|T201|OSN|3255-7|LNC|fibrinogen|fibrinogen
C0482705|T201|LC|3255-7|LNC|fibrinogen|fibrinogen
C0482705|T201|MTH_LN|3255-7|LNC|fibrinogen activity|fibrinogen activity
C0482705|T201|LN|3255-7|LNC|fibrinogen activity|fibrinogen activity
C0482705|T201|OSN|3255-7|LNC|fibrinogen activity|fibrinogen activity
C0482705|T201|LC|3255-7|LNC|fibrinogen activity|fibrinogen activity
C0482780|T201|LN|4532-8|LNC|total hemolytic complement activity|total hemolytic complement activity
C0482780|T201|MTH_LN|4532-8|LNC|total hemolytic complement activity|total hemolytic complement activity
C0482780|T201|OSN|4532-8|LNC|total hemolytic complement activity|total hemolytic complement activity
C0482780|T201|LC|4532-8|LNC|total hemolytic complement activity|total hemolytic complement activity
C0482780|T201|LN|4532-8|LNC|CH50|CH50
C0482780|T201|MTH_LN|4532-8|LNC|CH50|CH50
C0482780|T201|OSN|4532-8|LNC|CH50|CH50
C0482780|T201|LC|4532-8|LNC|CH50|CH50
C0483101|T201|LN|5380-1|LNC|Autoimmune antibody|Autoimmune antibody
C0483101|T201|MTH_LN|5380-1|LNC|Autoimmune antibody|Autoimmune antibody
C0483101|T201|OSN|5380-1|LNC|Autoimmune antibody|Autoimmune antibody
C0483101|T201|LC|5380-1|LNC|Autoimmune antibody|Autoimmune antibody
C0483102|T201|LN|5381-9|LNC|Autoimmune antibody|Autoimmune antibody
C0483102|T201|MTH_LN|5381-9|LNC|Autoimmune antibody|Autoimmune antibody
C0483102|T201|OSN|5381-9|LNC|Autoimmune antibody|Autoimmune antibody
C0483102|T201|LC|5381-9|LNC|Autoimmune antibody|Autoimmune antibody
C0484424|T201|LN|6742-1|LNC|red|red
C0484424|T201|MTH_LN|6742-1|LNC|red|red
C0484424|T201|LC|6742-1|LNC|red|red
C0484424|T201|OSN|6742-1|LNC|red|red
C0484424|T201|LN|6742-1|LNC|erythrocytes|erythrocytes
C0484424|T201|MTH_LN|6742-1|LNC|erythrocytes|erythrocytes
C0484424|T201|LC|6742-1|LNC|erythrocytes|erythrocytes
C0484424|T201|OSN|6742-1|LNC|erythrocytes|erythrocytes
C0484424|T201|LN|6742-1|LNC|erythrocyte morphology|erythrocyte morphology
C0484424|T201|MTH_LN|6742-1|LNC|erythrocyte morphology|erythrocyte morphology
C0484424|T201|LC|6742-1|LNC|erythrocyte morphology|erythrocyte morphology
C0484424|T201|OSN|6742-1|LNC|erythrocyte morphology|erythrocyte morphology
C0484424|T201|LN|6742-1|LNC|erythroid lineage cell|erythroid lineage cell
C0484424|T201|MTH_LN|6742-1|LNC|erythroid lineage cell|erythroid lineage cell
C0484424|T201|LC|6742-1|LNC|erythroid lineage cell|erythroid lineage cell
C0484424|T201|OSN|6742-1|LNC|erythroid lineage cell|erythroid lineage cell
C0484430|T201|LN|6690-2|LNC|white count|white count
C0484430|T201|OSN|6690-2|LNC|white count|white count
C0484430|T201|MTH_LN|6690-2|LNC|white count|white count
C0484430|T201|LC|6690-2|LNC|white count|white count
C0484430|T201|LN|6690-2|LNC|leukocyte number|leukocyte number
C0484430|T201|OSN|6690-2|LNC|leukocyte number|leukocyte number
C0484430|T201|MTH_LN|6690-2|LNC|leukocyte number|leukocyte number
C0484430|T201|LC|6690-2|LNC|leukocyte number|leukocyte number
C0484430|T201|LN|6690-2|LNC|white cell count|white cell count
C0484430|T201|OSN|6690-2|LNC|white cell count|white cell count
C0484430|T201|MTH_LN|6690-2|LNC|white cell count|white cell count
C0484430|T201|LC|6690-2|LNC|white cell count|white cell count
C0484430|T201|LN|6690-2|LNC|leukocyte count|leukocyte count
C0484430|T201|OSN|6690-2|LNC|leukocyte count|leukocyte count
C0484430|T201|MTH_LN|6690-2|LNC|leukocyte count|leukocyte count
C0484430|T201|LC|6690-2|LNC|leukocyte count|leukocyte count
C0484511|T201|LN|10438-0|LNC|B cell count|B cell count
C0484511|T201|MTH_LN|10438-0|LNC|B cell count|B cell count
C0484511|T201|OSN|10438-0|LNC|B cell count|B cell count
C0484511|T201|LC|10438-0|LNC|B cell count|B cell count
C0484511|T201|LN|10438-0|LNC|B|B
C0484511|T201|MTH_LN|10438-0|LNC|B|B
C0484511|T201|OSN|10438-0|LNC|B|B
C0484511|T201|LC|10438-0|LNC|B|B
C0484511|T201|LN|10438-0|LNC|Increase in B|Increase in B
C0484511|T201|MTH_LN|10438-0|LNC|Increase in B|Increase in B
C0484511|T201|OSN|10438-0|LNC|Increase in B|Increase in B
C0484511|T201|LC|10438-0|LNC|Increase in B|Increase in B
C0484511|T201|LN|10438-0|LNC|Bs|Bs
C0484511|T201|MTH_LN|10438-0|LNC|Bs|Bs
C0484511|T201|OSN|10438-0|LNC|Bs|Bs
C0484511|T201|LC|10438-0|LNC|Bs|Bs
C0484511|T201|LN|10438-0|LNC|numbersB|numbersB
C0484511|T201|MTH_LN|10438-0|LNC|numbersB|numbersB
C0484511|T201|OSN|10438-0|LNC|numbersB|numbersB
C0484511|T201|LC|10438-0|LNC|numbersB|numbersB
C0484521|T201|LN|8101-8|LNC|CD8-positive T|CD8-positive T
C0484521|T201|LC|8101-8|LNC|CD8-positive T|CD8-positive T
C0484521|T201|MTH_LN|8101-8|LNC|CD8-positive T|CD8-positive T
C0484521|T201|OSN|8101-8|LNC|CD8-positive T|CD8-positive T
C0484521|T201|LN|8101-8|LNC|CD8+ T|CD8+ T
C0484521|T201|LC|8101-8|LNC|CD8+ T|CD8+ T
C0484521|T201|MTH_LN|8101-8|LNC|CD8+ T|CD8+ T
C0484521|T201|OSN|8101-8|LNC|CD8+ T|CD8+ T
C0484521|T201|LN|8101-8|LNC|CD8 T|CD8 T
C0484521|T201|LC|8101-8|LNC|CD8 T|CD8 T
C0484521|T201|MTH_LN|8101-8|LNC|CD8 T|CD8 T
C0484521|T201|OSN|8101-8|LNC|CD8 T|CD8 T
C0484548|T201|LN|8123-2|LNC|CD4-positive T|CD4-positive T
C0484548|T201|LC|8123-2|LNC|CD4-positive T|CD4-positive T
C0484548|T201|MTH_LN|8123-2|LNC|CD4-positive T|CD4-positive T
C0484548|T201|OSN|8123-2|LNC|CD4-positive T|CD4-positive T
C0484548|T201|LN|8123-2|LNC|CD4+ T|CD4+ T
C0484548|T201|LC|8123-2|LNC|CD4+ T|CD4+ T
C0484548|T201|MTH_LN|8123-2|LNC|CD4+ T|CD4+ T
C0484548|T201|OSN|8123-2|LNC|CD4+ T|CD4+ T
C0484548|T201|LN|8123-2|LNC|CD4 T|CD4 T
C0484548|T201|LC|8123-2|LNC|CD4 T|CD4 T
C0484548|T201|MTH_LN|8123-2|LNC|CD4 T|CD4 T
C0484548|T201|OSN|8123-2|LNC|CD4 T|CD4 T
C0484571|T201|LN|9612-3|LNC|cortisol|cortisol
C0484571|T201|MTH_LN|9612-3|LNC|cortisol|cortisol
C0484571|T201|OSN|9612-3|LNC|cortisol|cortisol
C0484571|T201|LC|9612-3|LNC|cortisol|cortisol
C0484571|T201|LN|9612-3|LNC|cortisol low|cortisol low
C0484571|T201|MTH_LN|9612-3|LNC|cortisol low|cortisol low
C0484571|T201|OSN|9612-3|LNC|cortisol low|cortisol low
C0484571|T201|LC|9612-3|LNC|cortisol low|cortisol low
C0484571|T201|LN|9612-3|LNC|to undetectable cortisol|to undetectable cortisol
C0484571|T201|MTH_LN|9612-3|LNC|to undetectable cortisol|to undetectable cortisol
C0484571|T201|OSN|9612-3|LNC|to undetectable cortisol|to undetectable cortisol
C0484571|T201|LC|9612-3|LNC|to undetectable cortisol|to undetectable cortisol
C0484572|T201|LN|9613-1|LNC|cortisol|cortisol
C0484572|T201|MTH_LN|9613-1|LNC|cortisol|cortisol
C0484572|T201|OSN|9613-1|LNC|cortisol|cortisol
C0484572|T201|LC|9613-1|LNC|cortisol|cortisol
C0484572|T201|LN|9613-1|LNC|cortisol low|cortisol low
C0484572|T201|MTH_LN|9613-1|LNC|cortisol low|cortisol low
C0484572|T201|OSN|9613-1|LNC|cortisol low|cortisol low
C0484572|T201|LC|9613-1|LNC|cortisol low|cortisol low
C0484572|T201|LN|9613-1|LNC|to undetectable cortisol|to undetectable cortisol
C0484572|T201|MTH_LN|9613-1|LNC|to undetectable cortisol|to undetectable cortisol
C0484572|T201|OSN|9613-1|LNC|to undetectable cortisol|to undetectable cortisol
C0484572|T201|LC|9613-1|LNC|to undetectable cortisol|to undetectable cortisol
C0484573|T201|LN|9614-9|LNC|cortisol|cortisol
C0484573|T201|MTH_LN|9614-9|LNC|cortisol|cortisol
C0484573|T201|OSN|9614-9|LNC|cortisol|cortisol
C0484573|T201|LC|9614-9|LNC|cortisol|cortisol
C0484573|T201|LN|9614-9|LNC|cortisol low|cortisol low
C0484573|T201|MTH_LN|9614-9|LNC|cortisol low|cortisol low
C0484573|T201|OSN|9614-9|LNC|cortisol low|cortisol low
C0484573|T201|LC|9614-9|LNC|cortisol low|cortisol low
C0484573|T201|LN|9614-9|LNC|to undetectable cortisol|to undetectable cortisol
C0484573|T201|MTH_LN|9614-9|LNC|to undetectable cortisol|to undetectable cortisol
C0484573|T201|OSN|9614-9|LNC|to undetectable cortisol|to undetectable cortisol
C0484573|T201|LC|9614-9|LNC|to undetectable cortisol|to undetectable cortisol
C0484574|T201|LN|9615-6|LNC|cortisol|cortisol
C0484574|T201|OSN|9615-6|LNC|cortisol|cortisol
C0484574|T201|MTH_LN|9615-6|LNC|cortisol|cortisol
C0484574|T201|LC|9615-6|LNC|cortisol|cortisol
C0484574|T201|LN|9615-6|LNC|cortisol low|cortisol low
C0484574|T201|OSN|9615-6|LNC|cortisol low|cortisol low
C0484574|T201|MTH_LN|9615-6|LNC|cortisol low|cortisol low
C0484574|T201|LC|9615-6|LNC|cortisol low|cortisol low
C0484574|T201|LN|9615-6|LNC|to undetectable cortisol|to undetectable cortisol
C0484574|T201|OSN|9615-6|LNC|to undetectable cortisol|to undetectable cortisol
C0484574|T201|MTH_LN|9615-6|LNC|to undetectable cortisol|to undetectable cortisol
C0484574|T201|LC|9615-6|LNC|to undetectable cortisol|to undetectable cortisol
C0484575|T201|LN|10332-5|LNC|cortisol|cortisol
C0484575|T201|MTH_LN|10332-5|LNC|cortisol|cortisol
C0484575|T201|OSN|10332-5|LNC|cortisol|cortisol
C0484575|T201|LC|10332-5|LNC|cortisol|cortisol
C0484575|T201|LN|10332-5|LNC|cortisol low|cortisol low
C0484575|T201|MTH_LN|10332-5|LNC|cortisol low|cortisol low
C0484575|T201|OSN|10332-5|LNC|cortisol low|cortisol low
C0484575|T201|LC|10332-5|LNC|cortisol low|cortisol low
C0484575|T201|LN|10332-5|LNC|to undetectable cortisol|to undetectable cortisol
C0484575|T201|MTH_LN|10332-5|LNC|to undetectable cortisol|to undetectable cortisol
C0484575|T201|OSN|10332-5|LNC|to undetectable cortisol|to undetectable cortisol
C0484575|T201|LC|10332-5|LNC|to undetectable cortisol|to undetectable cortisol
C0484581|T201|LN|10449-7|LNC|glucose|glucose
C0484581|T201|MTH_LN|10449-7|LNC|glucose|glucose
C0484581|T201|OSN|10449-7|LNC|glucose|glucose
C0484581|T201|LC|10449-7|LNC|glucose|glucose
C0484599|T201|LN|10450-5|LNC|glucose|glucose
C0484599|T201|MTH_LN|10450-5|LNC|glucose|glucose
C0484599|T201|OSN|10450-5|LNC|glucose|glucose
C0484599|T201|LC|10450-5|LNC|glucose|glucose
C0484638|T201|MTH_LN|6768-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0484638|T201|LN|6768-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0484638|T201|OSN|6768-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0484638|T201|LC|6768-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0484638|T201|MTH_LN|6768-6|LNC|Greatly alkaline phosphatase|Greatly alkaline phosphatase
C0484638|T201|LN|6768-6|LNC|Greatly alkaline phosphatase|Greatly alkaline phosphatase
C0484638|T201|OSN|6768-6|LNC|Greatly alkaline phosphatase|Greatly alkaline phosphatase
C0484638|T201|LC|6768-6|LNC|Greatly alkaline phosphatase|Greatly alkaline phosphatase
C0484638|T201|MTH_LN|6768-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0484638|T201|LN|6768-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0484638|T201|OSN|6768-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0484638|T201|LC|6768-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0484673|T201|LN|6874-2|LNC|calcium|calcium
C0484673|T201|MTH_LN|6874-2|LNC|calcium|calcium
C0484673|T201|OSN|6874-2|LNC|calcium|calcium
C0484673|T201|LC|6874-2|LNC|calcium|calcium
C0484692|T201|LN|6687-8|LNC|citrate|citrate
C0484692|T201|MTH_LN|6687-8|LNC|citrate|citrate
C0484692|T201|OSN|6687-8|LNC|citrate|citrate
C0484692|T201|LC|6687-8|LNC|citrate|citrate
C0484702|T201|LN|6879-1|LNC|ACTH|ACTH
C0484702|T201|MTH_LN|6879-1|LNC|ACTH|ACTH
C0484702|T201|OSN|6879-1|LNC|ACTH|ACTH
C0484702|T201|LC|6879-1|LNC|ACTH|ACTH
C0484702|T201|LN|6879-1|LNC|corticotropin|corticotropin
C0484702|T201|MTH_LN|6879-1|LNC|corticotropin|corticotropin
C0484702|T201|OSN|6879-1|LNC|corticotropin|corticotropin
C0484702|T201|LC|6879-1|LNC|corticotropin|corticotropin
C0484702|T201|LN|6879-1|LNC|adrenocorticotropin|adrenocorticotropin
C0484702|T201|MTH_LN|6879-1|LNC|adrenocorticotropin|adrenocorticotropin
C0484702|T201|OSN|6879-1|LNC|adrenocorticotropin|adrenocorticotropin
C0484702|T201|LC|6879-1|LNC|adrenocorticotropin|adrenocorticotropin
C0484705|T201|LC|9813-7|LNC|cortisol|cortisol
C0484705|T201|OSN|9813-7|LNC|cortisol|cortisol
C0484705|T201|MTH_LN|9813-7|LNC|cortisol|cortisol
C0484705|T201|LN|9813-7|LNC|cortisol|cortisol
C0484705|T201|LC|9813-7|LNC|cortisol low|cortisol low
C0484705|T201|OSN|9813-7|LNC|cortisol low|cortisol low
C0484705|T201|MTH_LN|9813-7|LNC|cortisol low|cortisol low
C0484705|T201|LN|9813-7|LNC|cortisol low|cortisol low
C0484705|T201|LC|9813-7|LNC|to undetectable cortisol|to undetectable cortisol
C0484705|T201|OSN|9813-7|LNC|to undetectable cortisol|to undetectable cortisol
C0484705|T201|MTH_LN|9813-7|LNC|to undetectable cortisol|to undetectable cortisol
C0484705|T201|LN|9813-7|LNC|to undetectable cortisol|to undetectable cortisol
C0484731|T201|MTH_LN|2345-7|LNC|glucose|glucose
C0484731|T201|LN|2345-7|LNC|glucose|glucose
C0484731|T201|OSN|2345-7|LNC|glucose|glucose
C0484731|T201|LC|2345-7|LNC|glucose|glucose
C0484734|T201|LN|10336-6|LNC|gonadotropin|gonadotropin
C0484734|T201|MTH_LN|10336-6|LNC|gonadotropin|gonadotropin
C0484734|T201|OSN|10336-6|LNC|gonadotropin|gonadotropin
C0484734|T201|LC|10336-6|LNC|gonadotropin|gonadotropin
C0484796|T201|LN|10501-5|LNC|luteinizing|luteinizing
C0484796|T201|MTH_LN|10501-5|LNC|luteinizing|luteinizing
C0484796|T201|OSN|10501-5|LNC|luteinizing|luteinizing
C0484796|T201|LC|10501-5|LNC|luteinizing|luteinizing
C0484796|T201|LN|10501-5|LNC|LH|LH
C0484796|T201|MTH_LN|10501-5|LNC|LH|LH
C0484796|T201|OSN|10501-5|LNC|LH|LH
C0484796|T201|LC|10501-5|LNC|LH|LH
C0484796|T201|LN|10501-5|LNC|luteinising|luteinising
C0484796|T201|MTH_LN|10501-5|LNC|luteinising|luteinising
C0484796|T201|OSN|10501-5|LNC|luteinising|luteinising
C0484796|T201|LC|10501-5|LNC|luteinising|luteinising
C0484841|T201|LN|9324-5|LNC|taurine|taurine
C0484841|T201|MTH_LN|9324-5|LNC|taurine|taurine
C0484841|T201|OSN|9324-5|LNC|taurine|taurine
C0484841|T201|LC|9324-5|LNC|taurine|taurine
C0484848|T201|LN|6892-4|LNC|thyroxine|thyroxine
C0484848|T201|MTH_LN|6892-4|LNC|thyroxine|thyroxine
C0484848|T201|OSN|6892-4|LNC|thyroxine|thyroxine
C0484848|T201|LC|6892-4|LNC|thyroxine|thyroxine
C0484848|T201|LN|6892-4|LNC|T4|T4
C0484848|T201|MTH_LN|6892-4|LNC|T4|T4
C0484848|T201|OSN|6892-4|LNC|T4|T4
C0484848|T201|LC|6892-4|LNC|T4|T4
C0484850|T201|LN|6597-9|LNC|troponin T|troponin T
C0484850|T201|MTH_LN|6597-9|LNC|troponin T|troponin T
C0484850|T201|OSN|6597-9|LNC|troponin T|troponin T
C0484850|T201|LC|6597-9|LNC|troponin T|troponin T
C0484851|T201|LN|6598-7|LNC|troponin T|troponin T
C0484851|T201|MTH_LN|6598-7|LNC|troponin T|troponin T
C0484851|T201|OSN|6598-7|LNC|troponin T|troponin T
C0484851|T201|LC|6598-7|LNC|troponin T|troponin T
C0484958|T201|LN|10340-8|LNC|xenobiotic|xenobiotic
C0484958|T201|MTH_LN|10340-8|LNC|xenobiotic|xenobiotic
C0484958|T201|OSN|10340-8|LNC|xenobiotic|xenobiotic
C0484958|T201|LC|10340-8|LNC|xenobiotic|xenobiotic
C0484970|T201|LN|10341-6|LNC|xenobiotic|xenobiotic
C0484970|T201|MTH_LN|10341-6|LNC|xenobiotic|xenobiotic
C0484970|T201|OSN|10341-6|LNC|xenobiotic|xenobiotic
C0484970|T201|LC|10341-6|LNC|xenobiotic|xenobiotic
C0485074|T201|LN|10611-2|LNC|sperm motility|sperm motility
C0485074|T201|MTH_LN|10611-2|LNC|sperm motility|sperm motility
C0485074|T201|LC|10611-2|LNC|sperm motility|sperm motility
C0485074|T201|OSN|10611-2|LNC|sperm motility|sperm motility
C0485076|T201|LN|10613-8|LNC|sperm count|sperm count
C0485076|T201|MTH_LN|10613-8|LNC|sperm count|sperm count
C0485076|T201|LC|10613-8|LNC|sperm count|sperm count
C0485076|T201|OSN|10613-8|LNC|sperm count|sperm count
C0485076|T201|LN|10613-8|LNC|spermatogenesis|spermatogenesis
C0485076|T201|MTH_LN|10613-8|LNC|spermatogenesis|spermatogenesis
C0485076|T201|LC|10613-8|LNC|spermatogenesis|spermatogenesis
C0485076|T201|OSN|10613-8|LNC|spermatogenesis|spermatogenesis
C0485076|T201|LN|10613-8|LNC|sperm development|sperm development
C0485076|T201|MTH_LN|10613-8|LNC|sperm development|sperm development
C0485076|T201|LC|10613-8|LNC|sperm development|sperm development
C0485076|T201|OSN|10613-8|LNC|sperm development|sperm development
C0485828|T201|LN|8058-0|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0485828|T201|MTH_LN|8058-0|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0485828|T201|OSN|8058-0|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0485828|T201|LC|8058-0|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0485832|T201|LN|8061-4|LNC|Antinuclear antibody|Antinuclear antibody
C0485832|T201|MTH_LN|8061-4|LNC|Antinuclear antibody|Antinuclear antibody
C0485832|T201|OSN|8061-4|LNC|Antinuclear antibody|Antinuclear antibody
C0485832|T201|LC|8061-4|LNC|Antinuclear antibody|Antinuclear antibody
C0485856|T201|LN|6925-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0485856|T201|MTH_LN|6925-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0485856|T201|OSN|6925-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0485856|T201|LC|6925-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0485857|T201|LN|6926-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0485857|T201|MTH_LN|6926-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0485857|T201|LC|6926-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0485857|T201|OSN|6926-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0485899|T201|LN|8098-6|LNC|Autoimmune antibody|Autoimmune antibody
C0485899|T201|OSN|8098-6|LNC|Autoimmune antibody|Autoimmune antibody
C0485899|T201|MTH_LN|8098-6|LNC|Autoimmune antibody|Autoimmune antibody
C0485899|T201|LC|8098-6|LNC|Autoimmune antibody|Autoimmune antibody
C0486102|T201|LN|10365-5|LNC|xenobiotic|xenobiotic
C0486102|T201|MTH_LN|10365-5|LNC|xenobiotic|xenobiotic
C0486102|T201|OSN|10365-5|LNC|xenobiotic|xenobiotic
C0486102|T201|LC|10365-5|LNC|xenobiotic|xenobiotic
C0486103|T201|LN|10366-3|LNC|cotinine|cotinine
C0486103|T201|MTH_LN|10366-3|LNC|cotinine|cotinine
C0486103|T201|OSN|10366-3|LNC|cotinine|cotinine
C0486103|T201|LC|10366-3|LNC|cotinine|cotinine
C0486210|T201|LN|8247-9|LNC|homeostasis|homeostasis
C0486210|T201|MTH_LN|8247-9|LNC|homeostasis|homeostasis
C0486210|T201|OSN|8247-9|LNC|homeostasis|homeostasis
C0486210|T201|LC|8247-9|LNC|homeostasis|homeostasis
C0487973|T201|LN|8287-5|LNC|head circumference|head circumference
C0487973|T201|MTH_LN|8287-5|LNC|head circumference|head circumference
C0487973|T201|OSN|8287-5|LNC|head circumference|head circumference
C0487973|T201|LC|8287-5|LNC|head circumference|head circumference
C0487973|T201|LN|8287-5|LNC|skull size|skull size
C0487973|T201|MTH_LN|8287-5|LNC|skull size|skull size
C0487973|T201|OSN|8287-5|LNC|skull size|skull size
C0487973|T201|LC|8287-5|LNC|skull size|skull size
C0487973|T201|LN|8287-5|LNC|head size|head size
C0487973|T201|MTH_LN|8287-5|LNC|head size|head size
C0487973|T201|OSN|8287-5|LNC|head size|head size
C0487973|T201|LC|8287-5|LNC|head size|head size
C0487973|T201|LN|8287-5|LNC|cranium size|cranium size
C0487973|T201|MTH_LN|8287-5|LNC|cranium size|cranium size
C0487973|T201|OSN|8287-5|LNC|cranium size|cranium size
C0487973|T201|LC|8287-5|LNC|cranium size|cranium size
C0487995|T201|MTH_LN|8310-5|LNC|ly low body temperature|ly low body temperature
C0487995|T201|LC|8310-5|LNC|ly low body temperature|ly low body temperature
C0487995|T201|OSN|8310-5|LNC|ly low body temperature|ly low body temperature
C0487995|T201|LN|8310-5|LNC|ly low body temperature|ly low body temperature
C0487995|T201|MTH_LN|8310-5|LNC|temperature regulation|temperature regulation
C0487995|T201|LC|8310-5|LNC|temperature regulation|temperature regulation
C0487995|T201|OSN|8310-5|LNC|temperature regulation|temperature regulation
C0487995|T201|LN|8310-5|LNC|temperature regulation|temperature regulation
C0488052|T201|MTH_LN|8462-4|LNC|diastolic pressure|diastolic pressure
C0488052|T201|LN|8462-4|LNC|diastolic pressure|diastolic pressure
C0488052|T201|LC|8462-4|LNC|diastolic pressure|diastolic pressure
C0488052|T201|OSN|8462-4|LNC|diastolic pressure|diastolic pressure
C0488052|T201|MTH_LN|8462-4|LNC|systemic pressure|systemic pressure
C0488052|T201|LN|8462-4|LNC|systemic pressure|systemic pressure
C0488052|T201|LC|8462-4|LNC|systemic pressure|systemic pressure
C0488052|T201|OSN|8462-4|LNC|systemic pressure|systemic pressure
C0488055|T201|MTH_LN|8480-6|LNC|systolic pressure|systolic pressure
C0488055|T201|LN|8480-6|LNC|systolic pressure|systolic pressure
C0488055|T201|LC|8480-6|LNC|systolic pressure|systolic pressure
C0488055|T201|OSN|8480-6|LNC|systolic pressure|systolic pressure
C0488055|T201|MTH_LN|8480-6|LNC|systemic pressure|systemic pressure
C0488055|T201|LN|8480-6|LNC|systemic pressure|systemic pressure
C0488055|T201|LC|8480-6|LNC|systemic pressure|systemic pressure
C0488055|T201|OSN|8480-6|LNC|systemic pressure|systemic pressure
C0488223|T201|LN|8453-3|LNC|diastolic pressure|diastolic pressure
C0488223|T201|MTH_LN|8453-3|LNC|diastolic pressure|diastolic pressure
C0488223|T201|LC|8453-3|LNC|diastolic pressure|diastolic pressure
C0488223|T201|OSN|8453-3|LNC|diastolic pressure|diastolic pressure
C0488223|T201|LN|8453-3|LNC|systemic pressure|systemic pressure
C0488223|T201|MTH_LN|8453-3|LNC|systemic pressure|systemic pressure
C0488223|T201|LC|8453-3|LNC|systemic pressure|systemic pressure
C0488223|T201|OSN|8453-3|LNC|systemic pressure|systemic pressure
C0488224|T201|LN|8454-1|LNC|diastolic pressure|diastolic pressure
C0488224|T201|MTH_LN|8454-1|LNC|diastolic pressure|diastolic pressure
C0488224|T201|LC|8454-1|LNC|diastolic pressure|diastolic pressure
C0488224|T201|OSN|8454-1|LNC|diastolic pressure|diastolic pressure
C0488224|T201|LN|8454-1|LNC|systemic pressure|systemic pressure
C0488224|T201|MTH_LN|8454-1|LNC|systemic pressure|systemic pressure
C0488224|T201|LC|8454-1|LNC|systemic pressure|systemic pressure
C0488224|T201|OSN|8454-1|LNC|systemic pressure|systemic pressure
C0488225|T201|LN|8455-8|LNC|diastolic pressure|diastolic pressure
C0488225|T201|MTH_LN|8455-8|LNC|diastolic pressure|diastolic pressure
C0488225|T201|OSN|8455-8|LNC|diastolic pressure|diastolic pressure
C0488225|T201|LC|8455-8|LNC|diastolic pressure|diastolic pressure
C0488225|T201|LN|8455-8|LNC|systemic pressure|systemic pressure
C0488225|T201|MTH_LN|8455-8|LNC|systemic pressure|systemic pressure
C0488225|T201|OSN|8455-8|LNC|systemic pressure|systemic pressure
C0488225|T201|LC|8455-8|LNC|systemic pressure|systemic pressure
C0488229|T201|LN|8459-0|LNC|systemic pressure|systemic pressure
C0488229|T201|MTH_LN|8459-0|LNC|systemic pressure|systemic pressure
C0488229|T201|LC|8459-0|LNC|systemic pressure|systemic pressure
C0488229|T201|OSN|8459-0|LNC|systemic pressure|systemic pressure
C0488230|T201|LN|8460-8|LNC|systemic pressure|systemic pressure
C0488230|T201|MTH_LN|8460-8|LNC|systemic pressure|systemic pressure
C0488230|T201|LC|8460-8|LNC|systemic pressure|systemic pressure
C0488230|T201|OSN|8460-8|LNC|systemic pressure|systemic pressure
C0488231|T201|LN|8461-6|LNC|systemic pressure|systemic pressure
C0488231|T201|MTH_LN|8461-6|LNC|systemic pressure|systemic pressure
C0488231|T201|OSN|8461-6|LNC|systemic pressure|systemic pressure
C0488231|T201|LC|8461-6|LNC|systemic pressure|systemic pressure
C0488794|T201|LC|8867-4|LNC|heart rate|heart rate
C0488794|T201|OSN|8867-4|LNC|heart rate|heart rate
C0488794|T201|MTH_LN|8867-4|LNC|heart rate|heart rate
C0488794|T201|LN|8867-4|LNC|heart rate|heart rate
C0488794|T201|LC|8867-4|LNC|cardiac conduction|cardiac conduction
C0488794|T201|OSN|8867-4|LNC|cardiac conduction|cardiac conduction
C0488794|T201|MTH_LN|8867-4|LNC|cardiac conduction|cardiac conduction
C0488794|T201|LN|8867-4|LNC|cardiac conduction|cardiac conduction
C0488794|T201|LC|8867-4|LNC|Cardiac conductionities|Cardiac conductionities
C0488794|T201|OSN|8867-4|LNC|Cardiac conductionities|Cardiac conductionities
C0488794|T201|MTH_LN|8867-4|LNC|Cardiac conductionities|Cardiac conductionities
C0488794|T201|LN|8867-4|LNC|Cardiac conductionities|Cardiac conductionities
C0489258|T201|MTH_LN|9279-1|LNC|respiratory rate or depthbreathing|respiratory rate or depthbreathing
C0489258|T201|LC|9279-1|LNC|respiratory rate or depthbreathing|respiratory rate or depthbreathing
C0489258|T201|LN|9279-1|LNC|respiratory rate or depthbreathing|respiratory rate or depthbreathing
C0489258|T201|OSN|9279-1|LNC|respiratory rate or depthbreathing|respiratory rate or depthbreathing
C0489258|T201|MTH_LN|9279-1|LNC|patternrespiration|patternrespiration
C0489258|T201|LC|9279-1|LNC|patternrespiration|patternrespiration
C0489258|T201|LN|9279-1|LNC|patternrespiration|patternrespiration
C0489258|T201|OSN|9279-1|LNC|patternrespiration|patternrespiration
C0489258|T201|MTH_LN|9279-1|LNC|respiratory patterns|respiratory patterns
C0489258|T201|LC|9279-1|LNC|respiratory patterns|respiratory patterns
C0489258|T201|LN|9279-1|LNC|respiratory patterns|respiratory patterns
C0489258|T201|OSN|9279-1|LNC|respiratory patterns|respiratory patterns
C0549842|T201|LN|11125-2|LNC|platelet morphology|platelet morphology
C0549842|T201|MTH_LN|11125-2|LNC|platelet morphology|platelet morphology
C0549842|T201|OSN|11125-2|LNC|platelet morphology|platelet morphology
C0549842|T201|LC|11125-2|LNC|platelet morphology|platelet morphology
C0549842|T201|LN|11125-2|LNC|shapeplatelets|shapeplatelets
C0549842|T201|MTH_LN|11125-2|LNC|shapeplatelets|shapeplatelets
C0549842|T201|OSN|11125-2|LNC|shapeplatelets|shapeplatelets
C0549842|T201|LC|11125-2|LNC|shapeplatelets|shapeplatelets
C0549854|T201|LN|12250-7|LNC|reticulocytes|reticulocytes
C0549854|T201|OSN|12250-7|LNC|reticulocytes|reticulocytes
C0549854|T201|LC|12250-7|LNC|reticulocytes|reticulocytes
C0549854|T201|MTH_LN|12250-7|LNC|reticulocytes|reticulocytes
C0549854|T201|LN|12250-7|LNC|reticulocyte count|reticulocyte count
C0549854|T201|OSN|12250-7|LNC|reticulocyte count|reticulocyte count
C0549854|T201|LC|12250-7|LNC|reticulocyte count|reticulocyte count
C0549854|T201|MTH_LN|12250-7|LNC|reticulocyte count|reticulocyte count
C0549872|T201|MTH_LN|13336-3|LNC|naive T|naive T
C0549872|T201|LN|13336-3|LNC|naive T|naive T
C0549872|T201|LC|13336-3|LNC|naive T|naive T
C0549872|T201|OSN|13336-3|LNC|naive T|naive T
C0549872|T201|MTH_LN|13336-3|LNC|naive T cell|naive T cell
C0549872|T201|LN|13336-3|LNC|naive T cell|naive T cell
C0549872|T201|LC|13336-3|LNC|naive T cell|naive T cell
C0549872|T201|OSN|13336-3|LNC|naive T cell|naive T cell
C0549888|T201|LN|13040-1|LNC|C-peptide|C-peptide
C0549888|T201|OSN|13040-1|LNC|C-peptide|C-peptide
C0549888|T201|MTH_LN|13040-1|LNC|C-peptide|C-peptide
C0549888|T201|LC|13040-1|LNC|C-peptide|C-peptide
C0549888|T201|LN|13040-1|LNC|C peptide|C peptide
C0549888|T201|OSN|13040-1|LNC|C peptide|C peptide
C0549888|T201|MTH_LN|13040-1|LNC|C peptide|C peptide
C0549888|T201|LC|13040-1|LNC|C peptide|C peptide
C0549889|T201|LN|13039-3|LNC|C-peptide|C-peptide
C0549889|T201|MTH_LN|13039-3|LNC|C-peptide|C-peptide
C0549889|T201|OSN|13039-3|LNC|C-peptide|C-peptide
C0549889|T201|LC|13039-3|LNC|C-peptide|C-peptide
C0549889|T201|LN|13039-3|LNC|C peptide|C peptide
C0549889|T201|MTH_LN|13039-3|LNC|C peptide|C peptide
C0549889|T201|OSN|13039-3|LNC|C peptide|C peptide
C0549889|T201|LC|13039-3|LNC|C peptide|C peptide
C0549890|T201|LN|13042-7|LNC|C-peptide|C-peptide
C0549890|T201|OSN|13042-7|LNC|C-peptide|C-peptide
C0549890|T201|MTH_LN|13042-7|LNC|C-peptide|C-peptide
C0549890|T201|LC|13042-7|LNC|C-peptide|C-peptide
C0549890|T201|LN|13042-7|LNC|C peptide|C peptide
C0549890|T201|OSN|13042-7|LNC|C peptide|C peptide
C0549890|T201|MTH_LN|13042-7|LNC|C peptide|C peptide
C0549890|T201|LC|13042-7|LNC|C peptide|C peptide
C0549891|T201|LN|13041-9|LNC|C-peptide|C-peptide
C0549891|T201|MTH_LN|13041-9|LNC|C-peptide|C-peptide
C0549891|T201|OSN|13041-9|LNC|C-peptide|C-peptide
C0549891|T201|LC|13041-9|LNC|C-peptide|C-peptide
C0549891|T201|LN|13041-9|LNC|C peptide|C peptide
C0549891|T201|MTH_LN|13041-9|LNC|C peptide|C peptide
C0549891|T201|OSN|13041-9|LNC|C peptide|C peptide
C0549891|T201|LC|13041-9|LNC|C peptide|C peptide
C0549892|T201|LN|13032-8|LNC|C-peptide|C-peptide
C0549892|T201|MTH_LN|13032-8|LNC|C-peptide|C-peptide
C0549892|T201|OSN|13032-8|LNC|C-peptide|C-peptide
C0549892|T201|LC|13032-8|LNC|C-peptide|C-peptide
C0549892|T201|LN|13032-8|LNC|C peptide|C peptide
C0549892|T201|MTH_LN|13032-8|LNC|C peptide|C peptide
C0549892|T201|OSN|13032-8|LNC|C peptide|C peptide
C0549892|T201|LC|13032-8|LNC|C peptide|C peptide
C0549893|T201|LN|13038-5|LNC|C-peptide|C-peptide
C0549893|T201|MTH_LN|13038-5|LNC|C-peptide|C-peptide
C0549893|T201|OSN|13038-5|LNC|C-peptide|C-peptide
C0549893|T201|LC|13038-5|LNC|C-peptide|C-peptide
C0549893|T201|LN|13038-5|LNC|C peptide|C peptide
C0549893|T201|MTH_LN|13038-5|LNC|C peptide|C peptide
C0549893|T201|OSN|13038-5|LNC|C peptide|C peptide
C0549893|T201|LC|13038-5|LNC|C peptide|C peptide
C0549894|T201|LN|13043-5|LNC|C-peptide|C-peptide
C0549894|T201|MTH_LN|13043-5|LNC|C-peptide|C-peptide
C0549894|T201|OSN|13043-5|LNC|C-peptide|C-peptide
C0549894|T201|LC|13043-5|LNC|C-peptide|C-peptide
C0549894|T201|LN|13043-5|LNC|C peptide|C peptide
C0549894|T201|MTH_LN|13043-5|LNC|C peptide|C peptide
C0549894|T201|OSN|13043-5|LNC|C peptide|C peptide
C0549894|T201|LC|13043-5|LNC|C peptide|C peptide
C0549895|T201|LN|13033-6|LNC|C-peptide|C-peptide
C0549895|T201|MTH_LN|13033-6|LNC|C-peptide|C-peptide
C0549895|T201|OSN|13033-6|LNC|C-peptide|C-peptide
C0549895|T201|LC|13033-6|LNC|C-peptide|C-peptide
C0549895|T201|LN|13033-6|LNC|C peptide|C peptide
C0549895|T201|MTH_LN|13033-6|LNC|C peptide|C peptide
C0549895|T201|OSN|13033-6|LNC|C peptide|C peptide
C0549895|T201|LC|13033-6|LNC|C peptide|C peptide
C0549896|T201|LN|13034-4|LNC|C-peptide|C-peptide
C0549896|T201|MTH_LN|13034-4|LNC|C-peptide|C-peptide
C0549896|T201|OSN|13034-4|LNC|C-peptide|C-peptide
C0549896|T201|LC|13034-4|LNC|C-peptide|C-peptide
C0549896|T201|LN|13034-4|LNC|C peptide|C peptide
C0549896|T201|MTH_LN|13034-4|LNC|C peptide|C peptide
C0549896|T201|OSN|13034-4|LNC|C peptide|C peptide
C0549896|T201|LC|13034-4|LNC|C peptide|C peptide
C0549897|T201|LN|13044-3|LNC|C-peptide|C-peptide
C0549897|T201|MTH_LN|13044-3|LNC|C-peptide|C-peptide
C0549897|T201|OSN|13044-3|LNC|C-peptide|C-peptide
C0549897|T201|LC|13044-3|LNC|C-peptide|C-peptide
C0549897|T201|LN|13044-3|LNC|C peptide|C peptide
C0549897|T201|MTH_LN|13044-3|LNC|C peptide|C peptide
C0549897|T201|OSN|13044-3|LNC|C peptide|C peptide
C0549897|T201|LC|13044-3|LNC|C peptide|C peptide
C0549898|T201|LN|13035-1|LNC|C-peptide|C-peptide
C0549898|T201|MTH_LN|13035-1|LNC|C-peptide|C-peptide
C0549898|T201|OSN|13035-1|LNC|C-peptide|C-peptide
C0549898|T201|LC|13035-1|LNC|C-peptide|C-peptide
C0549898|T201|LN|13035-1|LNC|C peptide|C peptide
C0549898|T201|MTH_LN|13035-1|LNC|C peptide|C peptide
C0549898|T201|OSN|13035-1|LNC|C peptide|C peptide
C0549898|T201|LC|13035-1|LNC|C peptide|C peptide
C0549899|T201|LN|13045-0|LNC|C-peptide|C-peptide
C0549899|T201|MTH_LN|13045-0|LNC|C-peptide|C-peptide
C0549899|T201|OSN|13045-0|LNC|C-peptide|C-peptide
C0549899|T201|LC|13045-0|LNC|C-peptide|C-peptide
C0549899|T201|LN|13045-0|LNC|C peptide|C peptide
C0549899|T201|MTH_LN|13045-0|LNC|C peptide|C peptide
C0549899|T201|OSN|13045-0|LNC|C peptide|C peptide
C0549899|T201|LC|13045-0|LNC|C peptide|C peptide
C0549900|T201|LN|13036-9|LNC|C-peptide|C-peptide
C0549900|T201|MTH_LN|13036-9|LNC|C-peptide|C-peptide
C0549900|T201|OSN|13036-9|LNC|C-peptide|C-peptide
C0549900|T201|LC|13036-9|LNC|C-peptide|C-peptide
C0549900|T201|LN|13036-9|LNC|C peptide|C peptide
C0549900|T201|MTH_LN|13036-9|LNC|C peptide|C peptide
C0549900|T201|OSN|13036-9|LNC|C peptide|C peptide
C0549900|T201|LC|13036-9|LNC|C peptide|C peptide
C0549901|T201|LN|13037-7|LNC|C-peptide|C-peptide
C0549901|T201|MTH_LN|13037-7|LNC|C-peptide|C-peptide
C0549901|T201|OSN|13037-7|LNC|C-peptide|C-peptide
C0549901|T201|LC|13037-7|LNC|C-peptide|C-peptide
C0549901|T201|LN|13037-7|LNC|C peptide|C peptide
C0549901|T201|MTH_LN|13037-7|LNC|C peptide|C peptide
C0549901|T201|OSN|13037-7|LNC|C peptide|C peptide
C0549901|T201|LC|13037-7|LNC|C peptide|C peptide
C0549916|T201|LN|12458-6|LNC|adrenocorticotropin|adrenocorticotropin
C0549916|T201|MTH_LN|12458-6|LNC|adrenocorticotropin|adrenocorticotropin
C0549916|T201|OSN|12458-6|LNC|adrenocorticotropin|adrenocorticotropin
C0549916|T201|LC|12458-6|LNC|adrenocorticotropin|adrenocorticotropin
C0549916|T201|LN|12458-6|LNC|ACTH|ACTH
C0549916|T201|MTH_LN|12458-6|LNC|ACTH|ACTH
C0549916|T201|OSN|12458-6|LNC|ACTH|ACTH
C0549916|T201|LC|12458-6|LNC|ACTH|ACTH
C0549917|T201|LN|12459-4|LNC|adrenocorticotropin|adrenocorticotropin
C0549917|T201|MTH_LN|12459-4|LNC|adrenocorticotropin|adrenocorticotropin
C0549917|T201|OSN|12459-4|LNC|adrenocorticotropin|adrenocorticotropin
C0549917|T201|LC|12459-4|LNC|adrenocorticotropin|adrenocorticotropin
C0549917|T201|LN|12459-4|LNC|ACTH|ACTH
C0549917|T201|MTH_LN|12459-4|LNC|ACTH|ACTH
C0549917|T201|OSN|12459-4|LNC|ACTH|ACTH
C0549917|T201|LC|12459-4|LNC|ACTH|ACTH
C0549918|T201|LN|12460-2|LNC|adrenocorticotropin|adrenocorticotropin
C0549918|T201|MTH_LN|12460-2|LNC|adrenocorticotropin|adrenocorticotropin
C0549918|T201|OSN|12460-2|LNC|adrenocorticotropin|adrenocorticotropin
C0549918|T201|LC|12460-2|LNC|adrenocorticotropin|adrenocorticotropin
C0549918|T201|LN|12460-2|LNC|ACTH|ACTH
C0549918|T201|MTH_LN|12460-2|LNC|ACTH|ACTH
C0549918|T201|OSN|12460-2|LNC|ACTH|ACTH
C0549918|T201|LC|12460-2|LNC|ACTH|ACTH
C0549919|T201|LN|12461-0|LNC|adrenocorticotropin|adrenocorticotropin
C0549919|T201|MTH_LN|12461-0|LNC|adrenocorticotropin|adrenocorticotropin
C0549919|T201|OSN|12461-0|LNC|adrenocorticotropin|adrenocorticotropin
C0549919|T201|LC|12461-0|LNC|adrenocorticotropin|adrenocorticotropin
C0549919|T201|LN|12461-0|LNC|ACTH|ACTH
C0549919|T201|MTH_LN|12461-0|LNC|ACTH|ACTH
C0549919|T201|OSN|12461-0|LNC|ACTH|ACTH
C0549919|T201|LC|12461-0|LNC|ACTH|ACTH
C0549920|T201|LN|12462-8|LNC|adrenocorticotropin|adrenocorticotropin
C0549920|T201|MTH_LN|12462-8|LNC|adrenocorticotropin|adrenocorticotropin
C0549920|T201|OSN|12462-8|LNC|adrenocorticotropin|adrenocorticotropin
C0549920|T201|LC|12462-8|LNC|adrenocorticotropin|adrenocorticotropin
C0549920|T201|LN|12462-8|LNC|ACTH|ACTH
C0549920|T201|MTH_LN|12462-8|LNC|ACTH|ACTH
C0549920|T201|OSN|12462-8|LNC|ACTH|ACTH
C0549920|T201|LC|12462-8|LNC|ACTH|ACTH
C0549921|T201|LN|12463-6|LNC|adrenocorticotropin|adrenocorticotropin
C0549921|T201|MTH_LN|12463-6|LNC|adrenocorticotropin|adrenocorticotropin
C0549921|T201|OSN|12463-6|LNC|adrenocorticotropin|adrenocorticotropin
C0549921|T201|LC|12463-6|LNC|adrenocorticotropin|adrenocorticotropin
C0549921|T201|LN|12463-6|LNC|ACTH|ACTH
C0549921|T201|MTH_LN|12463-6|LNC|ACTH|ACTH
C0549921|T201|OSN|12463-6|LNC|ACTH|ACTH
C0549921|T201|LC|12463-6|LNC|ACTH|ACTH
C0549922|T201|LN|12464-4|LNC|adrenocorticotropin|adrenocorticotropin
C0549922|T201|MTH_LN|12464-4|LNC|adrenocorticotropin|adrenocorticotropin
C0549922|T201|OSN|12464-4|LNC|adrenocorticotropin|adrenocorticotropin
C0549922|T201|LC|12464-4|LNC|adrenocorticotropin|adrenocorticotropin
C0549922|T201|LN|12464-4|LNC|ACTH|ACTH
C0549922|T201|MTH_LN|12464-4|LNC|ACTH|ACTH
C0549922|T201|OSN|12464-4|LNC|ACTH|ACTH
C0549922|T201|LC|12464-4|LNC|ACTH|ACTH
C0549964|T201|LN|12645-8|LNC|glucose|glucose
C0549964|T201|MTH_LN|12645-8|LNC|glucose|glucose
C0549964|T201|OSN|12645-8|LNC|glucose|glucose
C0549964|T201|LC|12645-8|LNC|glucose|glucose
C0549965|T201|LN|12654-0|LNC|glucose|glucose
C0549965|T201|MTH_LN|12654-0|LNC|glucose|glucose
C0549965|T201|OSN|12654-0|LNC|glucose|glucose
C0549965|T201|LC|12654-0|LNC|glucose|glucose
C0549966|T201|LN|12651-6|LNC|glucose|glucose
C0549966|T201|MTH_LN|12651-6|LNC|glucose|glucose
C0549966|T201|OSN|12651-6|LNC|glucose|glucose
C0549966|T201|LC|12651-6|LNC|glucose|glucose
C0549967|T201|LN|12622-7|LNC|glucose|glucose
C0549967|T201|MTH_LN|12622-7|LNC|glucose|glucose
C0549967|T201|OSN|12622-7|LNC|glucose|glucose
C0549967|T201|LC|12622-7|LNC|glucose|glucose
C0549968|T201|LN|12623-5|LNC|glucose|glucose
C0549968|T201|MTH_LN|12623-5|LNC|glucose|glucose
C0549968|T201|OSN|12623-5|LNC|glucose|glucose
C0549968|T201|LC|12623-5|LNC|glucose|glucose
C0549969|T201|LN|12647-4|LNC|glucose|glucose
C0549969|T201|MTH_LN|12647-4|LNC|glucose|glucose
C0549969|T201|OSN|12647-4|LNC|glucose|glucose
C0549969|T201|LC|12647-4|LNC|glucose|glucose
C0549970|T201|LN|12624-3|LNC|glucose|glucose
C0549970|T201|MTH_LN|12624-3|LNC|glucose|glucose
C0549970|T201|OSN|12624-3|LNC|glucose|glucose
C0549970|T201|LC|12624-3|LNC|glucose|glucose
C0549971|T201|LN|12625-0|LNC|glucose|glucose
C0549971|T201|MTH_LN|12625-0|LNC|glucose|glucose
C0549971|T201|OSN|12625-0|LNC|glucose|glucose
C0549971|T201|LC|12625-0|LNC|glucose|glucose
C0549972|T201|LN|12626-8|LNC|glucose|glucose
C0549972|T201|MTH_LN|12626-8|LNC|glucose|glucose
C0549972|T201|OSN|12626-8|LNC|glucose|glucose
C0549972|T201|LC|12626-8|LNC|glucose|glucose
C0549973|T201|LN|10832-4|LNC|glucose|glucose
C0549973|T201|MTH_LN|10832-4|LNC|glucose|glucose
C0549973|T201|OSN|10832-4|LNC|glucose|glucose
C0549973|T201|LC|10832-4|LNC|glucose|glucose
C0549974|T201|LN|12639-1|LNC|glucose|glucose
C0549974|T201|MTH_LN|12639-1|LNC|glucose|glucose
C0549974|T201|OSN|12639-1|LNC|glucose|glucose
C0549974|T201|LC|12639-1|LNC|glucose|glucose
C0549975|T201|LN|12648-2|LNC|glucose|glucose
C0549975|T201|MTH_LN|12648-2|LNC|glucose|glucose
C0549975|T201|OSN|12648-2|LNC|glucose|glucose
C0549975|T201|LC|12648-2|LNC|glucose|glucose
C0549976|T201|LN|12627-6|LNC|glucose|glucose
C0549976|T201|MTH_LN|12627-6|LNC|glucose|glucose
C0549976|T201|OSN|12627-6|LNC|glucose|glucose
C0549976|T201|LC|12627-6|LNC|glucose|glucose
C0549977|T201|LN|12646-6|LNC|glucose|glucose
C0549977|T201|MTH_LN|12646-6|LNC|glucose|glucose
C0549977|T201|OSN|12646-6|LNC|glucose|glucose
C0549977|T201|LC|12646-6|LNC|glucose|glucose
C0549978|T201|LN|12615-1|LNC|glucose|glucose
C0549978|T201|MTH_LN|12615-1|LNC|glucose|glucose
C0549978|T201|OSN|12615-1|LNC|glucose|glucose
C0549978|T201|LC|12615-1|LNC|glucose|glucose
C0549980|T201|LN|12655-7|LNC|glucose|glucose
C0549980|T201|MTH_LN|12655-7|LNC|glucose|glucose
C0549980|T201|OSN|12655-7|LNC|glucose|glucose
C0549980|T201|LC|12655-7|LNC|glucose|glucose
C0549981|T201|LN|12610-2|LNC|glucose|glucose
C0549981|T201|MTH_LN|12610-2|LNC|glucose|glucose
C0549981|T201|OSN|12610-2|LNC|glucose|glucose
C0549981|T201|LC|12610-2|LNC|glucose|glucose
C0549982|T201|LN|12652-4|LNC|glucose|glucose
C0549982|T201|MTH_LN|12652-4|LNC|glucose|glucose
C0549982|T201|OSN|12652-4|LNC|glucose|glucose
C0549982|T201|LC|12652-4|LNC|glucose|glucose
C0549983|T201|LN|12616-9|LNC|glucose|glucose
C0549983|T201|MTH_LN|12616-9|LNC|glucose|glucose
C0549983|T201|OSN|12616-9|LNC|glucose|glucose
C0549983|T201|LC|12616-9|LNC|glucose|glucose
C0549985|T201|LN|12650-8|LNC|glucose|glucose
C0549985|T201|MTH_LN|12650-8|LNC|glucose|glucose
C0549985|T201|OSN|12650-8|LNC|glucose|glucose
C0549985|T201|LC|12650-8|LNC|glucose|glucose
C0549986|T201|LN|12617-7|LNC|glucose|glucose
C0549986|T201|MTH_LN|12617-7|LNC|glucose|glucose
C0549986|T201|OSN|12617-7|LNC|glucose|glucose
C0549986|T201|LC|12617-7|LNC|glucose|glucose
C0549988|T201|LN|12657-3|LNC|glucose|glucose
C0549988|T201|MTH_LN|12657-3|LNC|glucose|glucose
C0549988|T201|OSN|12657-3|LNC|glucose|glucose
C0549988|T201|LC|12657-3|LNC|glucose|glucose
C0549989|T201|LN|11032-0|LNC|glucose|glucose
C0549989|T201|MTH_LN|11032-0|LNC|glucose|glucose
C0549989|T201|OSN|11032-0|LNC|glucose|glucose
C0549989|T201|LC|11032-0|LNC|glucose|glucose
C0549990|T201|LN|12656-5|LNC|glucose|glucose
C0549990|T201|MTH_LN|12656-5|LNC|glucose|glucose
C0549990|T201|OSN|12656-5|LNC|glucose|glucose
C0549990|T201|LC|12656-5|LNC|glucose|glucose
C0549991|T201|LN|12618-5|LNC|glucose|glucose
C0549991|T201|MTH_LN|12618-5|LNC|glucose|glucose
C0549991|T201|OSN|12618-5|LNC|glucose|glucose
C0549991|T201|LC|12618-5|LNC|glucose|glucose
C0549992|T201|LN|12658-1|LNC|glucose|glucose
C0549992|T201|MTH_LN|12658-1|LNC|glucose|glucose
C0549992|T201|OSN|12658-1|LNC|glucose|glucose
C0549992|T201|LC|12658-1|LNC|glucose|glucose
C0549993|T201|LN|12619-3|LNC|glucose|glucose
C0549993|T201|MTH_LN|12619-3|LNC|glucose|glucose
C0549993|T201|OSN|12619-3|LNC|glucose|glucose
C0549993|T201|LC|12619-3|LNC|glucose|glucose
C0549994|T201|LN|12640-9|LNC|glucose|glucose
C0549994|T201|MTH_LN|12640-9|LNC|glucose|glucose
C0549994|T201|OSN|12640-9|LNC|glucose|glucose
C0549994|T201|LC|12640-9|LNC|glucose|glucose
C0549995|T201|LN|12620-1|LNC|glucose|glucose
C0549995|T201|MTH_LN|12620-1|LNC|glucose|glucose
C0549995|T201|OSN|12620-1|LNC|glucose|glucose
C0549995|T201|LC|12620-1|LNC|glucose|glucose
C0549996|T201|LN|12649-0|LNC|glucose|glucose
C0549996|T201|MTH_LN|12649-0|LNC|glucose|glucose
C0549996|T201|OSN|12649-0|LNC|glucose|glucose
C0549996|T201|LC|12649-0|LNC|glucose|glucose
C0549997|T201|LN|12642-5|LNC|glucose|glucose
C0549997|T201|MTH_LN|12642-5|LNC|glucose|glucose
C0549997|T201|OSN|12642-5|LNC|glucose|glucose
C0549997|T201|LC|12642-5|LNC|glucose|glucose
C0549998|T201|LN|12659-9|LNC|glucose|glucose
C0549998|T201|MTH_LN|12659-9|LNC|glucose|glucose
C0549998|T201|OSN|12659-9|LNC|glucose|glucose
C0549998|T201|LC|12659-9|LNC|glucose|glucose
C0549999|T201|LN|12641-7|LNC|glucose|glucose
C0549999|T201|MTH_LN|12641-7|LNC|glucose|glucose
C0549999|T201|OSN|12641-7|LNC|glucose|glucose
C0549999|T201|LC|12641-7|LNC|glucose|glucose
C0550000|T201|LN|12614-4|LNC|glucose|glucose
C0550000|T201|MTH_LN|12614-4|LNC|glucose|glucose
C0550000|T201|OSN|12614-4|LNC|glucose|glucose
C0550000|T201|LC|12614-4|LNC|glucose|glucose
C0550001|T201|LN|12643-3|LNC|glucose|glucose
C0550001|T201|MTH_LN|12643-3|LNC|glucose|glucose
C0550001|T201|OSN|12643-3|LNC|glucose|glucose
C0550001|T201|LC|12643-3|LNC|glucose|glucose
C0550002|T201|LN|12653-2|LNC|glucose|glucose
C0550002|T201|MTH_LN|12653-2|LNC|glucose|glucose
C0550002|T201|OSN|12653-2|LNC|glucose|glucose
C0550002|T201|LC|12653-2|LNC|glucose|glucose
C0550004|T201|LN|12644-1|LNC|glucose|glucose
C0550004|T201|MTH_LN|12644-1|LNC|glucose|glucose
C0550004|T201|OSN|12644-1|LNC|glucose|glucose
C0550004|T201|LC|12644-1|LNC|glucose|glucose
C0550005|T201|LN|12621-9|LNC|glucose|glucose
C0550005|T201|MTH_LN|12621-9|LNC|glucose|glucose
C0550005|T201|OSN|12621-9|LNC|glucose|glucose
C0550005|T201|LC|12621-9|LNC|glucose|glucose
C0550006|T201|LN|12638-3|LNC|glucose|glucose
C0550006|T201|MTH_LN|12638-3|LNC|glucose|glucose
C0550006|T201|OSN|12638-3|LNC|glucose|glucose
C0550006|T201|LC|12638-3|LNC|glucose|glucose
C0550041|T201|LN|10833-2|LNC|insulin|insulin
C0550041|T201|MTH_LN|10833-2|LNC|insulin|insulin
C0550041|T201|OSN|10833-2|LNC|insulin|insulin
C0550041|T201|LC|10833-2|LNC|insulin|insulin
C0550046|T201|LN|12672-2|LNC|luteinizing|luteinizing
C0550046|T201|MTH_LN|12672-2|LNC|luteinizing|luteinizing
C0550046|T201|OSN|12672-2|LNC|luteinizing|luteinizing
C0550046|T201|LC|12672-2|LNC|luteinizing|luteinizing
C0550046|T201|LN|12672-2|LNC|LH|LH
C0550046|T201|MTH_LN|12672-2|LNC|LH|LH
C0550046|T201|OSN|12672-2|LNC|LH|LH
C0550046|T201|LC|12672-2|LNC|LH|LH
C0550046|T201|LN|12672-2|LNC|luteinising|luteinising
C0550046|T201|MTH_LN|12672-2|LNC|luteinising|luteinising
C0550046|T201|OSN|12672-2|LNC|luteinising|luteinising
C0550046|T201|LC|12672-2|LNC|luteinising|luteinising
C0550047|T201|LN|12674-8|LNC|luteinizing|luteinizing
C0550047|T201|MTH_LN|12674-8|LNC|luteinizing|luteinizing
C0550047|T201|OSN|12674-8|LNC|luteinizing|luteinizing
C0550047|T201|LC|12674-8|LNC|luteinizing|luteinizing
C0550047|T201|LN|12674-8|LNC|LH|LH
C0550047|T201|MTH_LN|12674-8|LNC|LH|LH
C0550047|T201|OSN|12674-8|LNC|LH|LH
C0550047|T201|LC|12674-8|LNC|LH|LH
C0550047|T201|LN|12674-8|LNC|luteinising|luteinising
C0550047|T201|MTH_LN|12674-8|LNC|luteinising|luteinising
C0550047|T201|OSN|12674-8|LNC|luteinising|luteinising
C0550047|T201|LC|12674-8|LNC|luteinising|luteinising
C0550048|T201|LN|12675-5|LNC|luteinizing|luteinizing
C0550048|T201|MTH_LN|12675-5|LNC|luteinizing|luteinizing
C0550048|T201|OSN|12675-5|LNC|luteinizing|luteinizing
C0550048|T201|LC|12675-5|LNC|luteinizing|luteinizing
C0550048|T201|LN|12675-5|LNC|LH|LH
C0550048|T201|MTH_LN|12675-5|LNC|LH|LH
C0550048|T201|OSN|12675-5|LNC|LH|LH
C0550048|T201|LC|12675-5|LNC|LH|LH
C0550048|T201|LN|12675-5|LNC|luteinising|luteinising
C0550048|T201|MTH_LN|12675-5|LNC|luteinising|luteinising
C0550048|T201|OSN|12675-5|LNC|luteinising|luteinising
C0550048|T201|LC|12675-5|LNC|luteinising|luteinising
C0550049|T201|LN|12677-1|LNC|luteinizing|luteinizing
C0550049|T201|MTH_LN|12677-1|LNC|luteinizing|luteinizing
C0550049|T201|OSN|12677-1|LNC|luteinizing|luteinizing
C0550049|T201|LC|12677-1|LNC|luteinizing|luteinizing
C0550049|T201|LN|12677-1|LNC|LH|LH
C0550049|T201|MTH_LN|12677-1|LNC|LH|LH
C0550049|T201|OSN|12677-1|LNC|LH|LH
C0550049|T201|LC|12677-1|LNC|LH|LH
C0550049|T201|LN|12677-1|LNC|luteinising|luteinising
C0550049|T201|MTH_LN|12677-1|LNC|luteinising|luteinising
C0550049|T201|OSN|12677-1|LNC|luteinising|luteinising
C0550049|T201|LC|12677-1|LNC|luteinising|luteinising
C0550050|T201|LN|12673-0|LNC|luteinizing|luteinizing
C0550050|T201|MTH_LN|12673-0|LNC|luteinizing|luteinizing
C0550050|T201|OSN|12673-0|LNC|luteinizing|luteinizing
C0550050|T201|LC|12673-0|LNC|luteinizing|luteinizing
C0550050|T201|LN|12673-0|LNC|LH|LH
C0550050|T201|MTH_LN|12673-0|LNC|LH|LH
C0550050|T201|OSN|12673-0|LNC|LH|LH
C0550050|T201|LC|12673-0|LNC|LH|LH
C0550050|T201|LN|12673-0|LNC|luteinising|luteinising
C0550050|T201|MTH_LN|12673-0|LNC|luteinising|luteinising
C0550050|T201|OSN|12673-0|LNC|luteinising|luteinising
C0550050|T201|LC|12673-0|LNC|luteinising|luteinising
C0550051|T201|LN|12678-9|LNC|luteinizing|luteinizing
C0550051|T201|MTH_LN|12678-9|LNC|luteinizing|luteinizing
C0550051|T201|OSN|12678-9|LNC|luteinizing|luteinizing
C0550051|T201|LC|12678-9|LNC|luteinizing|luteinizing
C0550051|T201|LN|12678-9|LNC|LH|LH
C0550051|T201|MTH_LN|12678-9|LNC|LH|LH
C0550051|T201|OSN|12678-9|LNC|LH|LH
C0550051|T201|LC|12678-9|LNC|LH|LH
C0550051|T201|LN|12678-9|LNC|luteinising|luteinising
C0550051|T201|MTH_LN|12678-9|LNC|luteinising|luteinising
C0550051|T201|OSN|12678-9|LNC|luteinising|luteinising
C0550051|T201|LC|12678-9|LNC|luteinising|luteinising
C0550052|T201|LN|12676-3|LNC|luteinizing|luteinizing
C0550052|T201|MTH_LN|12676-3|LNC|luteinizing|luteinizing
C0550052|T201|OSN|12676-3|LNC|luteinizing|luteinizing
C0550052|T201|LC|12676-3|LNC|luteinizing|luteinizing
C0550052|T201|LN|12676-3|LNC|LH|LH
C0550052|T201|MTH_LN|12676-3|LNC|LH|LH
C0550052|T201|OSN|12676-3|LNC|LH|LH
C0550052|T201|LC|12676-3|LNC|LH|LH
C0550052|T201|LN|12676-3|LNC|luteinising|luteinising
C0550052|T201|MTH_LN|12676-3|LNC|luteinising|luteinising
C0550052|T201|OSN|12676-3|LNC|luteinising|luteinising
C0550052|T201|LC|12676-3|LNC|luteinising|luteinising
C0550053|T201|LN|12679-7|LNC|luteinizing|luteinizing
C0550053|T201|MTH_LN|12679-7|LNC|luteinizing|luteinizing
C0550053|T201|OSN|12679-7|LNC|luteinizing|luteinizing
C0550053|T201|LC|12679-7|LNC|luteinizing|luteinizing
C0550053|T201|LN|12679-7|LNC|LH|LH
C0550053|T201|MTH_LN|12679-7|LNC|LH|LH
C0550053|T201|OSN|12679-7|LNC|LH|LH
C0550053|T201|LC|12679-7|LNC|LH|LH
C0550053|T201|LN|12679-7|LNC|luteinising|luteinising
C0550053|T201|MTH_LN|12679-7|LNC|luteinising|luteinising
C0550053|T201|OSN|12679-7|LNC|luteinising|luteinising
C0550053|T201|LC|12679-7|LNC|luteinising|luteinising
C0550054|T201|LN|12680-5|LNC|luteinizing|luteinizing
C0550054|T201|MTH_LN|12680-5|LNC|luteinizing|luteinizing
C0550054|T201|OSN|12680-5|LNC|luteinizing|luteinizing
C0550054|T201|LC|12680-5|LNC|luteinizing|luteinizing
C0550054|T201|LN|12680-5|LNC|LH|LH
C0550054|T201|MTH_LN|12680-5|LNC|LH|LH
C0550054|T201|OSN|12680-5|LNC|LH|LH
C0550054|T201|LC|12680-5|LNC|LH|LH
C0550054|T201|LN|12680-5|LNC|luteinising|luteinising
C0550054|T201|MTH_LN|12680-5|LNC|luteinising|luteinising
C0550054|T201|OSN|12680-5|LNC|luteinising|luteinising
C0550054|T201|LC|12680-5|LNC|luteinising|luteinising
C0550055|T201|LN|12681-3|LNC|luteinizing|luteinizing
C0550055|T201|MTH_LN|12681-3|LNC|luteinizing|luteinizing
C0550055|T201|OSN|12681-3|LNC|luteinizing|luteinizing
C0550055|T201|LC|12681-3|LNC|luteinizing|luteinizing
C0550055|T201|LN|12681-3|LNC|LH|LH
C0550055|T201|MTH_LN|12681-3|LNC|LH|LH
C0550055|T201|OSN|12681-3|LNC|LH|LH
C0550055|T201|LC|12681-3|LNC|LH|LH
C0550055|T201|LN|12681-3|LNC|luteinising|luteinising
C0550055|T201|MTH_LN|12681-3|LNC|luteinising|luteinising
C0550055|T201|OSN|12681-3|LNC|luteinising|luteinising
C0550055|T201|LC|12681-3|LNC|luteinising|luteinising
C0550056|T201|LN|12682-1|LNC|luteinizing|luteinizing
C0550056|T201|MTH_LN|12682-1|LNC|luteinizing|luteinizing
C0550056|T201|OSN|12682-1|LNC|luteinizing|luteinizing
C0550056|T201|LC|12682-1|LNC|luteinizing|luteinizing
C0550056|T201|LN|12682-1|LNC|LH|LH
C0550056|T201|MTH_LN|12682-1|LNC|LH|LH
C0550056|T201|OSN|12682-1|LNC|LH|LH
C0550056|T201|LC|12682-1|LNC|LH|LH
C0550056|T201|LN|12682-1|LNC|luteinising|luteinising
C0550056|T201|MTH_LN|12682-1|LNC|luteinising|luteinising
C0550056|T201|OSN|12682-1|LNC|luteinising|luteinising
C0550056|T201|LC|12682-1|LNC|luteinising|luteinising
C0550057|T201|LN|12683-9|LNC|luteinizing|luteinizing
C0550057|T201|MTH_LN|12683-9|LNC|luteinizing|luteinizing
C0550057|T201|OSN|12683-9|LNC|luteinizing|luteinizing
C0550057|T201|LC|12683-9|LNC|luteinizing|luteinizing
C0550057|T201|LN|12683-9|LNC|LH|LH
C0550057|T201|MTH_LN|12683-9|LNC|LH|LH
C0550057|T201|OSN|12683-9|LNC|LH|LH
C0550057|T201|LC|12683-9|LNC|LH|LH
C0550057|T201|LN|12683-9|LNC|luteinising|luteinising
C0550057|T201|MTH_LN|12683-9|LNC|luteinising|luteinising
C0550057|T201|OSN|12683-9|LNC|luteinising|luteinising
C0550057|T201|LC|12683-9|LNC|luteinising|luteinising
C0550058|T201|LN|12684-7|LNC|luteinizing|luteinizing
C0550058|T201|MTH_LN|12684-7|LNC|luteinizing|luteinizing
C0550058|T201|OSN|12684-7|LNC|luteinizing|luteinizing
C0550058|T201|LC|12684-7|LNC|luteinizing|luteinizing
C0550058|T201|LN|12684-7|LNC|LH|LH
C0550058|T201|MTH_LN|12684-7|LNC|LH|LH
C0550058|T201|OSN|12684-7|LNC|LH|LH
C0550058|T201|LC|12684-7|LNC|LH|LH
C0550058|T201|LN|12684-7|LNC|luteinising|luteinising
C0550058|T201|MTH_LN|12684-7|LNC|luteinising|luteinising
C0550058|T201|OSN|12684-7|LNC|luteinising|luteinising
C0550058|T201|LC|12684-7|LNC|luteinising|luteinising
C0550178|T201|LN|11034-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0550178|T201|MTH_LN|11034-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0550178|T201|OSN|11034-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0550178|T201|LC|11034-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0550196|T201|MTH_LN|12960-1|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0550196|T201|LC|12960-1|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0550196|T201|OSN|12960-1|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0550196|T201|LN|12960-1|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0550202|T201|LN|12467-7|LNC|amino acid|amino acid
C0550202|T201|MTH_LN|12467-7|LNC|amino acid|amino acid
C0550202|T201|OSN|12467-7|LNC|amino acid|amino acid
C0550202|T201|LC|12467-7|LNC|amino acid|amino acid
C0550202|T201|LN|12467-7|LNC|animo acids|animo acids
C0550202|T201|MTH_LN|12467-7|LNC|animo acids|animo acids
C0550202|T201|OSN|12467-7|LNC|animo acids|animo acids
C0550202|T201|LC|12467-7|LNC|animo acids|animo acids
C0550202|T201|LN|12467-7|LNC|amino-acid findings|amino-acid findings
C0550202|T201|MTH_LN|12467-7|LNC|amino-acid findings|amino-acid findings
C0550202|T201|OSN|12467-7|LNC|amino-acid findings|amino-acid findings
C0550202|T201|LC|12467-7|LNC|amino-acid findings|amino-acid findings
C0550203|T201|LN|12177-2|LNC|amino acid|amino acid
C0550203|T201|MTH_LN|12177-2|LNC|amino acid|amino acid
C0550203|T201|OSN|12177-2|LNC|amino acid|amino acid
C0550203|T201|LC|12177-2|LNC|amino acid|amino acid
C0550203|T201|LN|12177-2|LNC|animo acids|animo acids
C0550203|T201|MTH_LN|12177-2|LNC|animo acids|animo acids
C0550203|T201|OSN|12177-2|LNC|animo acids|animo acids
C0550203|T201|LC|12177-2|LNC|animo acids|animo acids
C0550203|T201|LN|12177-2|LNC|amino-acid findings|amino-acid findings
C0550203|T201|MTH_LN|12177-2|LNC|amino-acid findings|amino-acid findings
C0550203|T201|OSN|12177-2|LNC|amino-acid findings|amino-acid findings
C0550203|T201|LC|12177-2|LNC|amino-acid findings|amino-acid findings
C0550239|T201|LN|12180-6|LNC|calcium|calcium
C0550239|T201|MTH_LN|12180-6|LNC|calcium|calcium
C0550239|T201|OSN|12180-6|LNC|calcium|calcium
C0550239|T201|LC|12180-6|LNC|calcium|calcium
C0550239|T201|LN|12180-6|LNC|calcium homeostasis|calcium homeostasis
C0550239|T201|MTH_LN|12180-6|LNC|calcium homeostasis|calcium homeostasis
C0550239|T201|OSN|12180-6|LNC|calcium homeostasis|calcium homeostasis
C0550239|T201|LC|12180-6|LNC|calcium homeostasis|calcium homeostasis
C0550242|T201|LN|13444-5|LNC|calcium|calcium
C0550242|T201|OSN|13444-5|LNC|calcium|calcium
C0550242|T201|MTH_LN|13444-5|LNC|calcium|calcium
C0550242|T201|LC|13444-5|LNC|calcium|calcium
C0550242|T201|LN|13444-5|LNC|calcium homeostasis|calcium homeostasis
C0550242|T201|OSN|13444-5|LNC|calcium homeostasis|calcium homeostasis
C0550242|T201|MTH_LN|13444-5|LNC|calcium homeostasis|calcium homeostasis
C0550242|T201|LC|13444-5|LNC|calcium homeostasis|calcium homeostasis
C0550246|T201|LN|11557-6|LNC|carbon dioxide|carbon dioxide
C0550246|T201|LC|11557-6|LNC|carbon dioxide|carbon dioxide
C0550246|T201|MTH_LN|11557-6|LNC|carbon dioxide|carbon dioxide
C0550246|T201|OSN|11557-6|LNC|carbon dioxide|carbon dioxide
C0550259|T201|LN|12772-0|LNC|HDL cholesterol|HDL cholesterol
C0550259|T201|MTH_LN|12772-0|LNC|HDL cholesterol|HDL cholesterol
C0550259|T201|OSN|12772-0|LNC|HDL cholesterol|HDL cholesterol
C0550259|T201|LC|12772-0|LNC|HDL cholesterol|HDL cholesterol
C0550259|T201|LN|12772-0|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0550259|T201|MTH_LN|12772-0|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0550259|T201|OSN|12772-0|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0550259|T201|LC|12772-0|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0550259|T201|LN|12772-0|LNC|HDL-cholesterol|HDL-cholesterol
C0550259|T201|MTH_LN|12772-0|LNC|HDL-cholesterol|HDL-cholesterol
C0550259|T201|OSN|12772-0|LNC|HDL-cholesterol|HDL-cholesterol
C0550259|T201|LC|12772-0|LNC|HDL-cholesterol|HDL-cholesterol
C0550259|T201|LN|12772-0|LNC|high-density lipoprotein|high-density lipoprotein
C0550259|T201|MTH_LN|12772-0|LNC|high-density lipoprotein|high-density lipoprotein
C0550259|T201|OSN|12772-0|LNC|high-density lipoprotein|high-density lipoprotein
C0550259|T201|LC|12772-0|LNC|high-density lipoprotein|high-density lipoprotein
C0550259|T201|LN|12772-0|LNC|HDL|HDL
C0550259|T201|MTH_LN|12772-0|LNC|HDL|HDL
C0550259|T201|OSN|12772-0|LNC|HDL|HDL
C0550259|T201|LC|12772-0|LNC|HDL|HDL
C0550261|T201|LN|12773-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0550261|T201|MTH_LN|12773-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0550261|T201|OSN|12773-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0550261|T201|LC|12773-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0550261|T201|LN|12773-8|LNC|LDL|LDL
C0550261|T201|MTH_LN|12773-8|LNC|LDL|LDL
C0550261|T201|OSN|12773-8|LNC|LDL|LDL
C0550261|T201|LC|12773-8|LNC|LDL|LDL
C0550261|T201|LN|12773-8|LNC|LDL cholesterol|LDL cholesterol
C0550261|T201|MTH_LN|12773-8|LNC|LDL cholesterol|LDL cholesterol
C0550261|T201|OSN|12773-8|LNC|LDL cholesterol|LDL cholesterol
C0550261|T201|LC|12773-8|LNC|LDL cholesterol|LDL cholesterol
C0550261|T201|LN|12773-8|LNC|low-density lipoprotein|low-density lipoprotein
C0550261|T201|MTH_LN|12773-8|LNC|low-density lipoprotein|low-density lipoprotein
C0550261|T201|OSN|12773-8|LNC|low-density lipoprotein|low-density lipoprotein
C0550261|T201|LC|12773-8|LNC|low-density lipoprotein|low-density lipoprotein
C0550261|T201|LN|12773-8|LNC|beta-lipoproteins|beta-lipoproteins
C0550261|T201|MTH_LN|12773-8|LNC|beta-lipoproteins|beta-lipoproteins
C0550261|T201|OSN|12773-8|LNC|beta-lipoproteins|beta-lipoproteins
C0550261|T201|LC|12773-8|LNC|beta-lipoproteins|beta-lipoproteins
C0550261|T201|LN|12773-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0550261|T201|MTH_LN|12773-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0550261|T201|OSN|12773-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0550261|T201|LC|12773-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0550261|T201|LN|12773-8|LNC|LDL-C|LDL-C
C0550261|T201|MTH_LN|12773-8|LNC|LDL-C|LDL-C
C0550261|T201|OSN|12773-8|LNC|LDL-C|LDL-C
C0550261|T201|LC|12773-8|LNC|LDL-C|LDL-C
C0550262|T201|LN|13459-3|LNC|VLDL cholesterol|VLDL cholesterol
C0550262|T201|OSN|13459-3|LNC|VLDL cholesterol|VLDL cholesterol
C0550262|T201|MTH_LN|13459-3|LNC|VLDL cholesterol|VLDL cholesterol
C0550262|T201|LC|13459-3|LNC|VLDL cholesterol|VLDL cholesterol
C0550262|T201|LN|13459-3|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0550262|T201|OSN|13459-3|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0550262|T201|MTH_LN|13459-3|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0550262|T201|LC|13459-3|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0550262|T201|LN|13459-3|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0550262|T201|OSN|13459-3|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0550262|T201|MTH_LN|13459-3|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0550262|T201|LC|13459-3|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0550264|T201|LN|13457-7|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0550264|T201|MTH_LN|13457-7|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0550264|T201|OSN|13457-7|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0550264|T201|LC|13457-7|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0550264|T201|LN|13457-7|LNC|LDL|LDL
C0550264|T201|MTH_LN|13457-7|LNC|LDL|LDL
C0550264|T201|OSN|13457-7|LNC|LDL|LDL
C0550264|T201|LC|13457-7|LNC|LDL|LDL
C0550264|T201|LN|13457-7|LNC|LDL cholesterol|LDL cholesterol
C0550264|T201|MTH_LN|13457-7|LNC|LDL cholesterol|LDL cholesterol
C0550264|T201|OSN|13457-7|LNC|LDL cholesterol|LDL cholesterol
C0550264|T201|LC|13457-7|LNC|LDL cholesterol|LDL cholesterol
C0550264|T201|LN|13457-7|LNC|low-density lipoprotein|low-density lipoprotein
C0550264|T201|MTH_LN|13457-7|LNC|low-density lipoprotein|low-density lipoprotein
C0550264|T201|OSN|13457-7|LNC|low-density lipoprotein|low-density lipoprotein
C0550264|T201|LC|13457-7|LNC|low-density lipoprotein|low-density lipoprotein
C0550264|T201|LN|13457-7|LNC|beta-lipoproteins|beta-lipoproteins
C0550264|T201|MTH_LN|13457-7|LNC|beta-lipoproteins|beta-lipoproteins
C0550264|T201|OSN|13457-7|LNC|beta-lipoproteins|beta-lipoproteins
C0550264|T201|LC|13457-7|LNC|beta-lipoproteins|beta-lipoproteins
C0550264|T201|LN|13457-7|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0550264|T201|MTH_LN|13457-7|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0550264|T201|OSN|13457-7|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0550264|T201|LC|13457-7|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0550264|T201|LN|13457-7|LNC|LDL-C|LDL-C
C0550264|T201|MTH_LN|13457-7|LNC|LDL-C|LDL-C
C0550264|T201|OSN|13457-7|LNC|LDL-C|LDL-C
C0550264|T201|LC|13457-7|LNC|LDL-C|LDL-C
C0550265|T201|LN|13458-5|LNC|VLDL cholesterol|VLDL cholesterol
C0550265|T201|MTH_LN|13458-5|LNC|VLDL cholesterol|VLDL cholesterol
C0550265|T201|OSN|13458-5|LNC|VLDL cholesterol|VLDL cholesterol
C0550265|T201|LC|13458-5|LNC|VLDL cholesterol|VLDL cholesterol
C0550265|T201|LN|13458-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0550265|T201|MTH_LN|13458-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0550265|T201|OSN|13458-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0550265|T201|LC|13458-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0550265|T201|LN|13458-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0550265|T201|MTH_LN|13458-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0550265|T201|OSN|13458-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0550265|T201|LC|13458-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0550276|T201|LN|11155-9|LNC|cortisol|cortisol
C0550276|T201|OSN|11155-9|LNC|cortisol|cortisol
C0550276|T201|MTH_LN|11155-9|LNC|cortisol|cortisol
C0550276|T201|LC|11155-9|LNC|cortisol|cortisol
C0550279|T201|LN|12187-1|LNC|creatine phosphokinase|creatine phosphokinase
C0550279|T201|MTH_LN|12187-1|LNC|creatine phosphokinase|creatine phosphokinase
C0550279|T201|LC|12187-1|LNC|creatine phosphokinase|creatine phosphokinase
C0550279|T201|OSN|12187-1|LNC|creatine phosphokinase|creatine phosphokinase
C0550279|T201|LN|12187-1|LNC|CPK|CPK
C0550279|T201|MTH_LN|12187-1|LNC|CPK|CPK
C0550279|T201|LC|12187-1|LNC|CPK|CPK
C0550279|T201|OSN|12187-1|LNC|CPK|CPK
C0550279|T201|LN|12187-1|LNC|creatine kinase|creatine kinase
C0550279|T201|MTH_LN|12187-1|LNC|creatine kinase|creatine kinase
C0550279|T201|LC|12187-1|LNC|creatine kinase|creatine kinase
C0550279|T201|OSN|12187-1|LNC|creatine kinase|creatine kinase
C0550279|T201|LN|12187-1|LNC|CK|CK
C0550279|T201|MTH_LN|12187-1|LNC|CK|CK
C0550279|T201|LC|12187-1|LNC|CK|CK
C0550279|T201|OSN|12187-1|LNC|CK|CK
C0550349|T201|LN|10834-0|LNC|antibody|antibody
C0550349|T201|MTH_LN|10834-0|LNC|antibody|antibody
C0550349|T201|OSN|10834-0|LNC|antibody|antibody
C0550349|T201|LC|10834-0|LNC|antibody|antibody
C0550349|T201|LN|10834-0|LNC|gamma globulin|gamma globulin
C0550349|T201|MTH_LN|10834-0|LNC|gamma globulin|gamma globulin
C0550349|T201|OSN|10834-0|LNC|gamma globulin|gamma globulin
C0550349|T201|LC|10834-0|LNC|gamma globulin|gamma globulin
C0550349|T201|LN|10834-0|LNC|immunoglobulin|immunoglobulin
C0550349|T201|MTH_LN|10834-0|LNC|immunoglobulin|immunoglobulin
C0550349|T201|OSN|10834-0|LNC|immunoglobulin|immunoglobulin
C0550349|T201|LC|10834-0|LNC|immunoglobulin|immunoglobulin
C0550349|T201|LN|10834-0|LNC|Raised immunoglobulin|Raised immunoglobulin
C0550349|T201|MTH_LN|10834-0|LNC|Raised immunoglobulin|Raised immunoglobulin
C0550349|T201|OSN|10834-0|LNC|Raised immunoglobulin|Raised immunoglobulin
C0550349|T201|LC|10834-0|LNC|Raised immunoglobulin|Raised immunoglobulin
C0550357|T201|LN|11142-7|LNC|glucose|glucose
C0550357|T201|MTH_LN|11142-7|LNC|glucose|glucose
C0550357|T201|OSN|11142-7|LNC|glucose|glucose
C0550357|T201|LC|11142-7|LNC|glucose|glucose
C0550363|T201|LN|11143-5|LNC|glucose|glucose
C0550363|T201|MTH_LN|11143-5|LNC|glucose|glucose
C0550363|T201|OSN|11143-5|LNC|glucose|glucose
C0550363|T201|LC|11143-5|LNC|glucose|glucose
C0550366|T201|LN|12611-0|LNC|glucose|glucose
C0550366|T201|MTH_LN|12611-0|LNC|glucose|glucose
C0550366|T201|OSN|12611-0|LNC|glucose|glucose
C0550366|T201|LC|12611-0|LNC|glucose|glucose
C0550439|T201|LN|13483-3|LNC|oxalate|oxalate
C0550439|T201|OSN|13483-3|LNC|oxalate|oxalate
C0550439|T201|MTH_LN|13483-3|LNC|oxalate|oxalate
C0550439|T201|LC|13483-3|LNC|oxalate|oxalate
C0550440|T201|LN|11556-8|LNC|oxygen|oxygen
C0550440|T201|LC|11556-8|LNC|oxygen|oxygen
C0550440|T201|MTH_LN|11556-8|LNC|oxygen|oxygen
C0550440|T201|OSN|11556-8|LNC|oxygen|oxygen
C0550447|T201|LN|11558-4|LNC|acid-base homeostasis|acid-base homeostasis
C0550447|T201|LC|11558-4|LNC|acid-base homeostasis|acid-base homeostasis
C0550447|T201|MTH_LN|11558-4|LNC|acid-base homeostasis|acid-base homeostasis
C0550447|T201|OSN|11558-4|LNC|acid-base homeostasis|acid-base homeostasis
C0550473|T201|LN|11148-4|LNC|potassium|potassium
C0550473|T201|OSN|11148-4|LNC|potassium|potassium
C0550473|T201|MTH_LN|11148-4|LNC|potassium|potassium
C0550473|T201|LC|11148-4|LNC|potassium|potassium
C0550513|T201|LN|11149-2|LNC|sodium|sodium
C0550513|T201|MTH_LN|11149-2|LNC|sodium|sodium
C0550513|T201|OSN|11149-2|LNC|sodium|sodium
C0550513|T201|LC|11149-2|LNC|sodium|sodium
C0550543|T201|LN|10839-9|LNC|troponin I|troponin I
C0550543|T201|MTH_LN|10839-9|LNC|troponin I|troponin I
C0550543|T201|OSN|10839-9|LNC|troponin I|troponin I
C0550543|T201|LC|10839-9|LNC|troponin I|troponin I
C0550551|T201|LN|12962-7|LNC|BUN|BUN
C0550551|T201|MTH_LN|12962-7|LNC|BUN|BUN
C0550551|T201|OSN|12962-7|LNC|BUN|BUN
C0550551|T201|LC|12962-7|LNC|BUN|BUN
C0550551|T201|LN|12962-7|LNC|urea nitrogen|urea nitrogen
C0550551|T201|MTH_LN|12962-7|LNC|urea nitrogen|urea nitrogen
C0550551|T201|OSN|12962-7|LNC|urea nitrogen|urea nitrogen
C0550551|T201|LC|12962-7|LNC|urea nitrogen|urea nitrogen
C0550576|T201|LN|12269-7|LNC|urobilinogen|urobilinogen
C0550576|T201|MTH_LN|12269-7|LNC|urobilinogen|urobilinogen
C0550576|T201|OSN|12269-7|LNC|urobilinogen|urobilinogen
C0550576|T201|LC|12269-7|LNC|urobilinogen|urobilinogen
C0550834|T201|LN|11151-8|LNC|reticulocytes|reticulocytes
C0550834|T201|MTH_LN|11151-8|LNC|reticulocytes|reticulocytes
C0550834|T201|LC|11151-8|LNC|reticulocytes|reticulocytes
C0550834|T201|OSN|11151-8|LNC|reticulocytes|reticulocytes
C0550834|T201|LN|11151-8|LNC|reticulocyte count|reticulocyte count
C0550834|T201|MTH_LN|11151-8|LNC|reticulocyte count|reticulocyte count
C0550834|T201|LC|11151-8|LNC|reticulocyte count|reticulocyte count
C0550834|T201|OSN|11151-8|LNC|reticulocyte count|reticulocyte count
C0550835|T201|LN|11271-4|LNC|reticulocytes|reticulocytes
C0550835|T201|MTH_LN|11271-4|LNC|reticulocytes|reticulocytes
C0550835|T201|LC|11271-4|LNC|reticulocytes|reticulocytes
C0550835|T201|OSN|11271-4|LNC|reticulocytes|reticulocytes
C0550835|T201|LN|11271-4|LNC|reticulocyte count|reticulocyte count
C0550835|T201|MTH_LN|11271-4|LNC|reticulocyte count|reticulocyte count
C0550835|T201|LC|11271-4|LNC|reticulocyte count|reticulocyte count
C0550835|T201|OSN|11271-4|LNC|reticulocyte count|reticulocyte count
C0550836|T201|LN|11153-4|LNC|reticulocytes|reticulocytes
C0550836|T201|MTH_LN|11153-4|LNC|reticulocytes|reticulocytes
C0550836|T201|LC|11153-4|LNC|reticulocytes|reticulocytes
C0550836|T201|OSN|11153-4|LNC|reticulocytes|reticulocytes
C0550836|T201|LN|11153-4|LNC|reticulocyte count|reticulocyte count
C0550836|T201|MTH_LN|11153-4|LNC|reticulocyte count|reticulocyte count
C0550836|T201|LC|11153-4|LNC|reticulocyte count|reticulocyte count
C0550836|T201|OSN|11153-4|LNC|reticulocyte count|reticulocyte count
C0550846|T201|LN|12227-5|LNC|white count|white count
C0550846|T201|OSN|12227-5|LNC|white count|white count
C0550846|T201|MTH_LN|12227-5|LNC|white count|white count
C0550846|T201|LC|12227-5|LNC|white count|white count
C0550846|T201|LN|12227-5|LNC|leukocyte number|leukocyte number
C0550846|T201|OSN|12227-5|LNC|leukocyte number|leukocyte number
C0550846|T201|MTH_LN|12227-5|LNC|leukocyte number|leukocyte number
C0550846|T201|LC|12227-5|LNC|leukocyte number|leukocyte number
C0550846|T201|LN|12227-5|LNC|white cell count|white cell count
C0550846|T201|OSN|12227-5|LNC|white cell count|white cell count
C0550846|T201|MTH_LN|12227-5|LNC|white cell count|white cell count
C0550846|T201|LC|12227-5|LNC|white cell count|white cell count
C0550846|T201|LN|12227-5|LNC|leukocyte count|leukocyte count
C0550846|T201|OSN|12227-5|LNC|leukocyte count|leukocyte count
C0550846|T201|MTH_LN|12227-5|LNC|leukocyte count|leukocyte count
C0550846|T201|LC|12227-5|LNC|leukocyte count|leukocyte count
C0551273|T201|LN|11560-0|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551273|T201|MTH_LN|11560-0|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551273|T201|OSN|11560-0|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551273|T201|LC|11560-0|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551274|T201|LN|11561-8|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551274|T201|MTH_LN|11561-8|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551274|T201|OSN|11561-8|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551274|T201|LC|11561-8|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551275|T201|LN|11562-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551275|T201|MTH_LN|11562-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551275|T201|OSN|11562-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551275|T201|LC|11562-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0551356|T201|LN|11572-5|LNC|Autoimmune antibody|Autoimmune antibody
C0551356|T201|LC|11572-5|LNC|Autoimmune antibody|Autoimmune antibody
C0551356|T201|OSN|11572-5|LNC|Autoimmune antibody|Autoimmune antibody
C0551356|T201|MTH_LN|11572-5|LNC|Autoimmune antibody|Autoimmune antibody
C0551405|T201|LN|12293-7|LNC|cotinine|cotinine
C0551405|T201|MTH_LN|12293-7|LNC|cotinine|cotinine
C0551405|T201|OSN|12293-7|LNC|cotinine|cotinine
C0551405|T201|LC|12293-7|LNC|cotinine|cotinine
C0551476|T201|LN|12552-6|LNC|propylene glycol|propylene glycol
C0551476|T201|MTH_LN|12552-6|LNC|propylene glycol|propylene glycol
C0551476|T201|OSN|12552-6|LNC|propylene glycol|propylene glycol
C0551476|T201|LC|12552-6|LNC|propylene glycol|propylene glycol
C0551476|T201|LN|12552-6|LNC|propane-1,2-diol|propane-1,2-diol
C0551476|T201|MTH_LN|12552-6|LNC|propane-1,2-diol|propane-1,2-diol
C0551476|T201|OSN|12552-6|LNC|propane-1,2-diol|propane-1,2-diol
C0551476|T201|LC|12552-6|LNC|propane-1,2-diol|propane-1,2-diol
C0682110|T098|LN|1516-4|LNC|glucose|glucose
C0682110|T098|MTH_LN|1516-4|LNC|glucose|glucose
C0682110|T098|OSN|1516-4|LNC|glucose|glucose
C0682110|T098|LC|1516-4|LNC|glucose|glucose
C0682111|T098|LN|1493-6|LNC|glucose|glucose
C0682111|T098|OSN|1493-6|LNC|glucose|glucose
C0682111|T098|MTH_LN|1493-6|LNC|glucose|glucose
C0682111|T098|LC|1493-6|LNC|glucose|glucose
C0682113|T098|LN|1416-7|LNC|cortisol|cortisol
C0682113|T098|MTH_LN|1416-7|LNC|cortisol|cortisol
C0682113|T098|OSN|1416-7|LNC|cortisol|cortisol
C0682113|T098|LC|1416-7|LNC|cortisol|cortisol
C0682113|T098|LN|1416-7|LNC|cortisol low|cortisol low
C0682113|T098|MTH_LN|1416-7|LNC|cortisol low|cortisol low
C0682113|T098|OSN|1416-7|LNC|cortisol low|cortisol low
C0682113|T098|LC|1416-7|LNC|cortisol low|cortisol low
C0682113|T098|LN|1416-7|LNC|to undetectable cortisol|to undetectable cortisol
C0682113|T098|MTH_LN|1416-7|LNC|to undetectable cortisol|to undetectable cortisol
C0682113|T098|OSN|1416-7|LNC|to undetectable cortisol|to undetectable cortisol
C0682113|T098|LC|1416-7|LNC|to undetectable cortisol|to undetectable cortisol
C0700436|T201|LN|1544-6|LNC|glucose|glucose
C0700436|T201|MTH_LN|1544-6|LNC|glucose|glucose
C0700436|T201|OSN|1544-6|LNC|glucose|glucose
C0700436|T201|LC|1544-6|LNC|glucose|glucose
C0796702|T201|LN|13508-7|LNC|reticulocytes|reticulocytes
C0796702|T201|MTH_LN|13508-7|LNC|reticulocytes|reticulocytes
C0796702|T201|LC|13508-7|LNC|reticulocytes|reticulocytes
C0796702|T201|OSN|13508-7|LNC|reticulocytes|reticulocytes
C0796702|T201|LN|13508-7|LNC|reticulocyte count|reticulocyte count
C0796702|T201|MTH_LN|13508-7|LNC|reticulocyte count|reticulocyte count
C0796702|T201|LC|13508-7|LNC|reticulocyte count|reticulocyte count
C0796702|T201|OSN|13508-7|LNC|reticulocyte count|reticulocyte count
C0796797|T201|LN|13606-9|LNC|glucose|glucose
C0796797|T201|MTH_LN|13606-9|LNC|glucose|glucose
C0796797|T201|OSN|13606-9|LNC|glucose|glucose
C0796797|T201|LC|13606-9|LNC|glucose|glucose
C0796798|T201|LN|13607-7|LNC|glucose|glucose
C0796798|T201|MTH_LN|13607-7|LNC|glucose|glucose
C0796798|T201|OSN|13607-7|LNC|glucose|glucose
C0796798|T201|LC|13607-7|LNC|glucose|glucose
C0796799|T201|LN|13608-5|LNC|insulin|insulin
C0796799|T201|OSN|13608-5|LNC|insulin|insulin
C0796799|T201|MTH_LN|13608-5|LNC|insulin|insulin
C0796799|T201|LC|13608-5|LNC|insulin|insulin
C0796800|T201|LN|13609-3|LNC|insulin|insulin
C0796800|T201|OSN|13609-3|LNC|insulin|insulin
C0796800|T201|MTH_LN|13609-3|LNC|insulin|insulin
C0796800|T201|LC|13609-3|LNC|insulin|insulin
C0796849|T201|LN|13658-0|LNC|urobilinogen|urobilinogen
C0796849|T201|MTH_LN|13658-0|LNC|urobilinogen|urobilinogen
C0796849|T201|OSN|13658-0|LNC|urobilinogen|urobilinogen
C0796849|T201|LC|13658-0|LNC|urobilinogen|urobilinogen
C0796899|T201|LN|13708-3|LNC|arginine|arginine
C0796899|T201|MTH_LN|13708-3|LNC|arginine|arginine
C0796899|T201|OSN|13708-3|LNC|arginine|arginine
C0796899|T201|LC|13708-3|LNC|arginine|arginine
C0796934|T201|LN|13744-8|LNC|galactose|galactose
C0796934|T201|OSN|13744-8|LNC|galactose|galactose
C0796934|T201|MTH_LN|13744-8|LNC|galactose|galactose
C0796934|T201|LC|13744-8|LNC|galactose|galactose
C0796977|T201|LN|13787-7|LNC|orotic acid|orotic acid
C0796977|T201|OSN|13787-7|LNC|orotic acid|orotic acid
C0796977|T201|MTH_LN|13787-7|LNC|orotic acid|orotic acid
C0796977|T201|LC|13787-7|LNC|orotic acid|orotic acid
C0797004|T201|LN|13814-9|LNC|taurine|taurine
C0797004|T201|OSN|13814-9|LNC|taurine|taurine
C0797004|T201|MTH_LN|13814-9|LNC|taurine|taurine
C0797004|T201|LC|13814-9|LNC|taurine|taurine
C0797024|T201|LN|13834-7|LNC|IgE|IgE
C0797024|T201|MTH_LN|13834-7|LNC|IgE|IgE
C0797024|T201|OSN|13834-7|LNC|IgE|IgE
C0797024|T201|LC|13834-7|LNC|IgE|IgE
C0797024|T201|LN|13834-7|LNC|immunoglobulin E|immunoglobulin E
C0797024|T201|MTH_LN|13834-7|LNC|immunoglobulin E|immunoglobulin E
C0797024|T201|OSN|13834-7|LNC|immunoglobulin E|immunoglobulin E
C0797024|T201|LC|13834-7|LNC|immunoglobulin E|immunoglobulin E
C0797041|T201|LN|13852-9|LNC|aldosterone|aldosterone
C0797041|T201|MTH_LN|13852-9|LNC|aldosterone|aldosterone
C0797041|T201|OSN|13852-9|LNC|aldosterone|aldosterone
C0797041|T201|LC|13852-9|LNC|aldosterone|aldosterone
C0797044|T201|LN|13855-2|LNC|aldosterone|aldosterone
C0797044|T201|MTH_LN|13855-2|LNC|aldosterone|aldosterone
C0797044|T201|OSN|13855-2|LNC|aldosterone|aldosterone
C0797044|T201|LC|13855-2|LNC|aldosterone|aldosterone
C0797045|T201|LN|13856-0|LNC|androstenedione|androstenedione
C0797045|T201|MTH_LN|13856-0|LNC|androstenedione|androstenedione
C0797045|T201|OSN|13856-0|LNC|androstenedione|androstenedione
C0797045|T201|LC|13856-0|LNC|androstenedione|androstenedione
C0797046|T201|LN|13857-8|LNC|androstenedione|androstenedione
C0797046|T201|MTH_LN|13857-8|LNC|androstenedione|androstenedione
C0797046|T201|OSN|13857-8|LNC|androstenedione|androstenedione
C0797046|T201|LC|13857-8|LNC|androstenedione|androstenedione
C0797047|T201|LN|13858-6|LNC|androstenedione|androstenedione
C0797047|T201|MTH_LN|13858-6|LNC|androstenedione|androstenedione
C0797047|T201|OSN|13858-6|LNC|androstenedione|androstenedione
C0797047|T201|LC|13858-6|LNC|androstenedione|androstenedione
C0797048|T201|LN|13859-4|LNC|C-peptide|C-peptide
C0797048|T201|MTH_LN|13859-4|LNC|C-peptide|C-peptide
C0797048|T201|OSN|13859-4|LNC|C-peptide|C-peptide
C0797048|T201|LC|13859-4|LNC|C-peptide|C-peptide
C0797048|T201|LN|13859-4|LNC|C peptide|C peptide
C0797048|T201|MTH_LN|13859-4|LNC|C peptide|C peptide
C0797048|T201|OSN|13859-4|LNC|C peptide|C peptide
C0797048|T201|LC|13859-4|LNC|C peptide|C peptide
C0797049|T201|LN|13860-2|LNC|C-peptide|C-peptide
C0797049|T201|MTH_LN|13860-2|LNC|C-peptide|C-peptide
C0797049|T201|OSN|13860-2|LNC|C-peptide|C-peptide
C0797049|T201|LC|13860-2|LNC|C-peptide|C-peptide
C0797049|T201|LN|13860-2|LNC|C peptide|C peptide
C0797049|T201|MTH_LN|13860-2|LNC|C peptide|C peptide
C0797049|T201|OSN|13860-2|LNC|C peptide|C peptide
C0797049|T201|LC|13860-2|LNC|C peptide|C peptide
C0797050|T201|LN|13861-0|LNC|C-peptide|C-peptide
C0797050|T201|MTH_LN|13861-0|LNC|C-peptide|C-peptide
C0797050|T201|OSN|13861-0|LNC|C-peptide|C-peptide
C0797050|T201|LC|13861-0|LNC|C-peptide|C-peptide
C0797050|T201|LN|13861-0|LNC|C peptide|C peptide
C0797050|T201|MTH_LN|13861-0|LNC|C peptide|C peptide
C0797050|T201|OSN|13861-0|LNC|C peptide|C peptide
C0797050|T201|LC|13861-0|LNC|C peptide|C peptide
C0797054|T201|LN|13865-1|LNC|glucose|glucose
C0797054|T201|OSN|13865-1|LNC|glucose|glucose
C0797054|T201|MTH_LN|13865-1|LNC|glucose|glucose
C0797054|T201|LC|13865-1|LNC|glucose|glucose
C0797055|T201|LN|13866-9|LNC|glucose|glucose
C0797055|T201|MTH_LN|13866-9|LNC|glucose|glucose
C0797055|T201|OSN|13866-9|LNC|glucose|glucose
C0797055|T201|LC|13866-9|LNC|glucose|glucose
C0797063|T201|LN|13874-3|LNC|Alkaline phosphatase|Alkaline phosphatase
C0797063|T201|MTH_LN|13874-3|LNC|Alkaline phosphatase|Alkaline phosphatase
C0797063|T201|OSN|13874-3|LNC|Alkaline phosphatase|Alkaline phosphatase
C0797063|T201|LC|13874-3|LNC|Alkaline phosphatase|Alkaline phosphatase
C0797063|T201|LN|13874-3|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0797063|T201|MTH_LN|13874-3|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0797063|T201|OSN|13874-3|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0797063|T201|LC|13874-3|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0797063|T201|LN|13874-3|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0797063|T201|MTH_LN|13874-3|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0797063|T201|OSN|13874-3|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0797063|T201|LC|13874-3|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0797064|T201|LN|13875-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0797064|T201|MTH_LN|13875-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0797064|T201|OSN|13875-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0797064|T201|LC|13875-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C0797064|T201|LN|13875-0|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0797064|T201|MTH_LN|13875-0|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0797064|T201|OSN|13875-0|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0797064|T201|LC|13875-0|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0797064|T201|LN|13875-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0797064|T201|MTH_LN|13875-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0797064|T201|OSN|13875-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0797064|T201|LC|13875-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0797129|T201|OSN|13941-0|LNC|lymphocyte count|lymphocyte count
C0797129|T201|LN|13941-0|LNC|lymphocyte count|lymphocyte count
C0797129|T201|MTH_LN|13941-0|LNC|lymphocyte count|lymphocyte count
C0797129|T201|LC|13941-0|LNC|lymphocyte count|lymphocyte count
C0797129|T201|OSN|13941-0|LNC|lymphocyte number|lymphocyte number
C0797129|T201|LN|13941-0|LNC|lymphocyte number|lymphocyte number
C0797129|T201|MTH_LN|13941-0|LNC|lymphocyte number|lymphocyte number
C0797129|T201|LC|13941-0|LNC|lymphocyte number|lymphocyte number
C0797129|T201|OSN|13941-0|LNC|lymphocyte counts|lymphocyte counts
C0797129|T201|LN|13941-0|LNC|lymphocyte counts|lymphocyte counts
C0797129|T201|MTH_LN|13941-0|LNC|lymphocyte counts|lymphocyte counts
C0797129|T201|LC|13941-0|LNC|lymphocyte counts|lymphocyte counts
C0797129|T201|OSN|13941-0|LNC|lymphocytes|lymphocytes
C0797129|T201|LN|13941-0|LNC|lymphocytes|lymphocytes
C0797129|T201|MTH_LN|13941-0|LNC|lymphocytes|lymphocytes
C0797129|T201|LC|13941-0|LNC|lymphocytes|lymphocytes
C0797129|T201|OSN|13941-0|LNC|numberslymphocytes|numberslymphocytes
C0797129|T201|LN|13941-0|LNC|numberslymphocytes|numberslymphocytes
C0797129|T201|MTH_LN|13941-0|LNC|numberslymphocytes|numberslymphocytes
C0797129|T201|LC|13941-0|LNC|numberslymphocytes|numberslymphocytes
C0797147|T201|LN|13959-2|LNC|calcium|calcium
C0797147|T201|MTH_LN|13959-2|LNC|calcium|calcium
C0797147|T201|OSN|13959-2|LNC|calcium|calcium
C0797147|T201|LC|13959-2|LNC|calcium|calcium
C0797147|T201|LN|13959-2|LNC|calcium homeostasis|calcium homeostasis
C0797147|T201|MTH_LN|13959-2|LNC|calcium homeostasis|calcium homeostasis
C0797147|T201|OSN|13959-2|LNC|calcium homeostasis|calcium homeostasis
C0797147|T201|LC|13959-2|LNC|calcium homeostasis|calcium homeostasis
C0797153|T201|LN|13965-9|LNC|homocystine|homocystine
C0797153|T201|OSN|13965-9|LNC|homocystine|homocystine
C0797153|T201|MTH_LN|13965-9|LNC|homocystine|homocystine
C0797153|T201|LC|13965-9|LNC|homocystine|homocystine
C0797153|T201|LN|13965-9|LNC|homocysteine metabolism|homocysteine metabolism
C0797153|T201|OSN|13965-9|LNC|homocysteine metabolism|homocysteine metabolism
C0797153|T201|MTH_LN|13965-9|LNC|homocysteine metabolism|homocysteine metabolism
C0797153|T201|LC|13965-9|LNC|homocysteine metabolism|homocysteine metabolism
C0797154|T201|LN|13966-7|LNC|cystine|cystine
C0797154|T201|MTH_LN|13966-7|LNC|cystine|cystine
C0797154|T201|OSN|13966-7|LNC|cystine|cystine
C0797154|T201|LC|13966-7|LNC|cystine|cystine
C0797157|T201|LN|13969-1|LNC|creatine kinase|creatine kinase
C0797157|T201|MTH_LN|13969-1|LNC|creatine kinase|creatine kinase
C0797157|T201|OSN|13969-1|LNC|creatine kinase|creatine kinase
C0797157|T201|LC|13969-1|LNC|creatine kinase|creatine kinase
C0797233|T201|LN|14045-9|LNC|lactate|lactate
C0797233|T201|MTH_LN|14045-9|LNC|lactate|lactate
C0797233|T201|OSN|14045-9|LNC|lactate|lactate
C0797233|T201|LC|14045-9|LNC|lactate|lactate
C0797304|T201|LC|14118-4|LNC|lactate|lactate
C0797304|T201|MTH_LN|14118-4|LNC|lactate|lactate
C0797304|T201|LN|14118-4|LNC|lactate|lactate
C0797304|T201|OSN|14118-4|LNC|lactate|lactate
C0797321|T201|LN|14135-8|LNC|CD8-positive T|CD8-positive T
C0797321|T201|LC|14135-8|LNC|CD8-positive T|CD8-positive T
C0797321|T201|OSN|14135-8|LNC|CD8-positive T|CD8-positive T
C0797321|T201|MTH_LN|14135-8|LNC|CD8-positive T|CD8-positive T
C0797321|T201|LN|14135-8|LNC|CD8+ T|CD8+ T
C0797321|T201|LC|14135-8|LNC|CD8+ T|CD8+ T
C0797321|T201|OSN|14135-8|LNC|CD8+ T|CD8+ T
C0797321|T201|MTH_LN|14135-8|LNC|CD8+ T|CD8+ T
C0797321|T201|LN|14135-8|LNC|CD8 T|CD8 T
C0797321|T201|LC|14135-8|LNC|CD8 T|CD8 T
C0797321|T201|OSN|14135-8|LNC|CD8 T|CD8 T
C0797321|T201|MTH_LN|14135-8|LNC|CD8 T|CD8 T
C0797323|T201|LN|14137-4|LNC|glucose|glucose
C0797323|T201|MTH_LN|14137-4|LNC|glucose|glucose
C0797323|T201|OSN|14137-4|LNC|glucose|glucose
C0797323|T201|LC|14137-4|LNC|glucose|glucose
C0797340|T201|LN|14155-6|LNC|VLDL cholesterol|VLDL cholesterol
C0797340|T201|MTH_LN|14155-6|LNC|VLDL cholesterol|VLDL cholesterol
C0797340|T201|OSN|14155-6|LNC|VLDL cholesterol|VLDL cholesterol
C0797340|T201|LC|14155-6|LNC|VLDL cholesterol|VLDL cholesterol
C0797340|T201|LN|14155-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0797340|T201|MTH_LN|14155-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0797340|T201|OSN|14155-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0797340|T201|LC|14155-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0797340|T201|LN|14155-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0797340|T201|MTH_LN|14155-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0797340|T201|OSN|14155-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0797340|T201|LC|14155-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0797381|T201|LN|14196-0|LNC|reticulocytes|reticulocytes
C0797381|T201|OSN|14196-0|LNC|reticulocytes|reticulocytes
C0797381|T201|MTH_LN|14196-0|LNC|reticulocytes|reticulocytes
C0797381|T201|LC|14196-0|LNC|reticulocytes|reticulocytes
C0797381|T201|LN|14196-0|LNC|reticulocyte count|reticulocyte count
C0797381|T201|OSN|14196-0|LNC|reticulocyte count|reticulocyte count
C0797381|T201|MTH_LN|14196-0|LNC|reticulocyte count|reticulocyte count
C0797381|T201|LC|14196-0|LNC|reticulocyte count|reticulocyte count
C0797464|T201|LN|14282-8|LNC|acylcarnitine|acylcarnitine
C0797464|T201|OSN|14282-8|LNC|acylcarnitine|acylcarnitine
C0797464|T201|MTH_LN|14282-8|LNC|acylcarnitine|acylcarnitine
C0797464|T201|LC|14282-8|LNC|acylcarnitine|acylcarnitine
C0797468|T201|LN|14286-9|LNC|Carnitine|Carnitine
C0797468|T201|OSN|14286-9|LNC|Carnitine|Carnitine
C0797468|T201|MTH_LN|14286-9|LNC|Carnitine|Carnitine
C0797468|T201|LC|14286-9|LNC|Carnitine|Carnitine
C0797468|T201|LN|14286-9|LNC|carnitine metabolism|carnitine metabolism
C0797468|T201|OSN|14286-9|LNC|carnitine metabolism|carnitine metabolism
C0797468|T201|MTH_LN|14286-9|LNC|carnitine metabolism|carnitine metabolism
C0797468|T201|LC|14286-9|LNC|carnitine metabolism|carnitine metabolism
C0797468|T201|LN|14286-9|LNC|total carnitine|total carnitine
C0797468|T201|OSN|14286-9|LNC|total carnitine|total carnitine
C0797468|T201|MTH_LN|14286-9|LNC|total carnitine|total carnitine
C0797468|T201|LC|14286-9|LNC|total carnitine|total carnitine
C0797470|T201|LN|14288-5|LNC|Carnitine|Carnitine
C0797470|T201|MTH_LN|14288-5|LNC|Carnitine|Carnitine
C0797470|T201|OSN|14288-5|LNC|Carnitine|Carnitine
C0797470|T201|LC|14288-5|LNC|Carnitine|Carnitine
C0797470|T201|LN|14288-5|LNC|carnitine metabolism|carnitine metabolism
C0797470|T201|MTH_LN|14288-5|LNC|carnitine metabolism|carnitine metabolism
C0797470|T201|OSN|14288-5|LNC|carnitine metabolism|carnitine metabolism
C0797470|T201|LC|14288-5|LNC|carnitine metabolism|carnitine metabolism
C0797470|T201|LN|14288-5|LNC|total carnitine|total carnitine
C0797470|T201|MTH_LN|14288-5|LNC|total carnitine|total carnitine
C0797470|T201|OSN|14288-5|LNC|total carnitine|total carnitine
C0797470|T201|LC|14288-5|LNC|total carnitine|total carnitine
// C0797471|T201|OLC|14290-1|LNC||
// C0797471|T201|MTH_LO|14290-1|LNC||
// C0797471|T201|LO|14290-1|LNC||
// C0797471|T201|OOSN|14290-1|LNC||
C0797471|T201|OLC|14290-1|LNC|occult|occult
C0797471|T201|MTH_LO|14290-1|LNC|occult|occult
C0797471|T201|LO|14290-1|LNC|occult|occult
C0797471|T201|OOSN|14290-1|LNC|occult|occult
C0797519|T201|LN|14338-8|LNC|Serum protein|Serum protein
C0797519|T201|MTH_LN|14338-8|LNC|Serum protein|Serum protein
C0797519|T201|OSN|14338-8|LNC|Serum protein|Serum protein
C0797519|T201|LC|14338-8|LNC|Serum protein|Serum protein
C0797519|T201|LN|14338-8|LNC|protein disease|protein disease
C0797519|T201|MTH_LN|14338-8|LNC|protein disease|protein disease
C0797519|T201|OSN|14338-8|LNC|protein disease|protein disease
C0797519|T201|LC|14338-8|LNC|protein disease|protein disease
C0797519|T201|LN|14338-8|LNC|protein|protein
C0797519|T201|MTH_LN|14338-8|LNC|protein|protein
C0797519|T201|OSN|14338-8|LNC|protein|protein
C0797519|T201|LC|14338-8|LNC|protein|protein
C0797519|T201|LN|14338-8|LNC|prealbumin|prealbumin
C0797519|T201|MTH_LN|14338-8|LNC|prealbumin|prealbumin
C0797519|T201|OSN|14338-8|LNC|prealbumin|prealbumin
C0797519|T201|LC|14338-8|LNC|prealbumin|prealbumin
C0797757|T201|LN|14581-3|LNC|xenobiotic|xenobiotic
C0797757|T201|OSN|14581-3|LNC|xenobiotic|xenobiotic
C0797757|T201|MTH_LN|14581-3|LNC|xenobiotic|xenobiotic
C0797757|T201|LC|14581-3|LNC|xenobiotic|xenobiotic
C0797803|T201|LN|14628-2|LNC|bile acid|bile acid
C0797803|T201|MTH_LN|14628-2|LNC|bile acid|bile acid
C0797803|T201|OSN|14628-2|LNC|bile acid|bile acid
C0797803|T201|LC|14628-2|LNC|bile acid|bile acid
C0797803|T201|LN|14628-2|LNC|bile|bile
C0797803|T201|MTH_LN|14628-2|LNC|bile|bile
C0797803|T201|OSN|14628-2|LNC|bile|bile
C0797803|T201|LC|14628-2|LNC|bile|bile
C0797808|T201|LN|14633-2|LNC|C-peptide|C-peptide
C0797808|T201|MTH_LN|14633-2|LNC|C-peptide|C-peptide
C0797808|T201|OSN|14633-2|LNC|C-peptide|C-peptide
C0797808|T201|LC|14633-2|LNC|C-peptide|C-peptide
C0797808|T201|LN|14633-2|LNC|C peptide|C peptide
C0797808|T201|MTH_LN|14633-2|LNC|C peptide|C peptide
C0797808|T201|OSN|14633-2|LNC|C peptide|C peptide
C0797808|T201|LC|14633-2|LNC|C peptide|C peptide
C0797821|T201|LN|14646-4|LNC|HDL cholesterol|HDL cholesterol
C0797821|T201|MTH_LN|14646-4|LNC|HDL cholesterol|HDL cholesterol
C0797821|T201|OSN|14646-4|LNC|HDL cholesterol|HDL cholesterol
C0797821|T201|LC|14646-4|LNC|HDL cholesterol|HDL cholesterol
C0797821|T201|LN|14646-4|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0797821|T201|MTH_LN|14646-4|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0797821|T201|OSN|14646-4|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0797821|T201|LC|14646-4|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0797821|T201|LN|14646-4|LNC|HDL-cholesterol|HDL-cholesterol
C0797821|T201|MTH_LN|14646-4|LNC|HDL-cholesterol|HDL-cholesterol
C0797821|T201|OSN|14646-4|LNC|HDL-cholesterol|HDL-cholesterol
C0797821|T201|LC|14646-4|LNC|HDL-cholesterol|HDL-cholesterol
C0797821|T201|LN|14646-4|LNC|high-density lipoprotein|high-density lipoprotein
C0797821|T201|MTH_LN|14646-4|LNC|high-density lipoprotein|high-density lipoprotein
C0797821|T201|OSN|14646-4|LNC|high-density lipoprotein|high-density lipoprotein
C0797821|T201|LC|14646-4|LNC|high-density lipoprotein|high-density lipoprotein
C0797821|T201|LN|14646-4|LNC|HDL|HDL
C0797821|T201|MTH_LN|14646-4|LNC|HDL|HDL
C0797821|T201|OSN|14646-4|LNC|HDL|HDL
C0797821|T201|LC|14646-4|LNC|HDL|HDL
C0797848|T201|LN|14674-6|LNC|ACTH|ACTH
C0797848|T201|MTH_LN|14674-6|LNC|ACTH|ACTH
C0797848|T201|OSN|14674-6|LNC|ACTH|ACTH
C0797848|T201|LC|14674-6|LNC|ACTH|ACTH
C0797848|T201|LN|14674-6|LNC|corticotropin|corticotropin
C0797848|T201|MTH_LN|14674-6|LNC|corticotropin|corticotropin
C0797848|T201|OSN|14674-6|LNC|corticotropin|corticotropin
C0797848|T201|LC|14674-6|LNC|corticotropin|corticotropin
C0797848|T201|LN|14674-6|LNC|adrenocorticotropin|adrenocorticotropin
C0797848|T201|MTH_LN|14674-6|LNC|adrenocorticotropin|adrenocorticotropin
C0797848|T201|OSN|14674-6|LNC|adrenocorticotropin|adrenocorticotropin
C0797848|T201|LC|14674-6|LNC|adrenocorticotropin|adrenocorticotropin
C0797906|T201|LN|14732-2|LNC|folate|folate
C0797906|T201|OSN|14732-2|LNC|folate|folate
C0797906|T201|MTH_LN|14732-2|LNC|folate|folate
C0797906|T201|LC|14732-2|LNC|folate|folate
C0797917|T201|LN|14743-9|LNC|glucose|glucose
C0797917|T201|MTH_LN|14743-9|LNC|glucose|glucose
C0797917|T201|OSN|14743-9|LNC|glucose|glucose
C0797917|T201|LC|14743-9|LNC|glucose|glucose
C0797918|T201|LN|14744-7|LNC|CSF glucose|CSF glucose
C0797918|T201|MTH_LN|14744-7|LNC|CSF glucose|CSF glucose
C0797918|T201|OSN|14744-7|LNC|CSF glucose|CSF glucose
C0797918|T201|LC|14744-7|LNC|CSF glucose|CSF glucose
C0797918|T201|LN|14744-7|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C0797918|T201|MTH_LN|14744-7|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C0797918|T201|OSN|14744-7|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C0797918|T201|LC|14744-7|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C0797923|T201|LN|14749-6|LNC|glucose|glucose
C0797923|T201|MTH_LN|14749-6|LNC|glucose|glucose
C0797923|T201|OSN|14749-6|LNC|glucose|glucose
C0797923|T201|LC|14749-6|LNC|glucose|glucose
C0797925|T201|LN|14751-2|LNC|glucose|glucose
C0797925|T201|OSN|14751-2|LNC|glucose|glucose
C0797925|T201|MTH_LN|14751-2|LNC|glucose|glucose
C0797925|T201|LC|14751-2|LNC|glucose|glucose
C0797926|T201|LN|14752-0|LNC|glucose|glucose
C0797926|T201|OSN|14752-0|LNC|glucose|glucose
C0797926|T201|MTH_LN|14752-0|LNC|glucose|glucose
C0797926|T201|LC|14752-0|LNC|glucose|glucose
C0797927|T201|LN|14753-8|LNC|glucose|glucose
C0797927|T201|MTH_LN|14753-8|LNC|glucose|glucose
C0797927|T201|OSN|14753-8|LNC|glucose|glucose
C0797927|T201|LC|14753-8|LNC|glucose|glucose
C0797928|T201|LN|14754-6|LNC|glucose|glucose
C0797928|T201|MTH_LN|14754-6|LNC|glucose|glucose
C0797928|T201|OSN|14754-6|LNC|glucose|glucose
C0797928|T201|LC|14754-6|LNC|glucose|glucose
C0797929|T201|LN|14755-3|LNC|glucose|glucose
C0797929|T201|MTH_LN|14755-3|LNC|glucose|glucose
C0797929|T201|OSN|14755-3|LNC|glucose|glucose
C0797929|T201|LC|14755-3|LNC|glucose|glucose
C0797930|T201|LN|14756-1|LNC|glucose|glucose
C0797930|T201|MTH_LN|14756-1|LNC|glucose|glucose
C0797930|T201|OSN|14756-1|LNC|glucose|glucose
C0797930|T201|LC|14756-1|LNC|glucose|glucose
C0797931|T201|LN|14757-9|LNC|glucose|glucose
C0797931|T201|MTH_LN|14757-9|LNC|glucose|glucose
C0797931|T201|OSN|14757-9|LNC|glucose|glucose
C0797931|T201|LC|14757-9|LNC|glucose|glucose
C0797932|T201|LN|14758-7|LNC|glucose|glucose
C0797932|T201|MTH_LN|14758-7|LNC|glucose|glucose
C0797932|T201|OSN|14758-7|LNC|glucose|glucose
C0797932|T201|LC|14758-7|LNC|glucose|glucose
C0797933|T201|LN|14759-5|LNC|glucose|glucose
C0797933|T201|MTH_LN|14759-5|LNC|glucose|glucose
C0797933|T201|OSN|14759-5|LNC|glucose|glucose
C0797933|T201|LC|14759-5|LNC|glucose|glucose
C0797934|T201|LN|14760-3|LNC|glucose|glucose
C0797934|T201|MTH_LN|14760-3|LNC|glucose|glucose
C0797934|T201|OSN|14760-3|LNC|glucose|glucose
C0797934|T201|LC|14760-3|LNC|glucose|glucose
C0797935|T201|LN|14761-1|LNC|glucose|glucose
C0797935|T201|MTH_LN|14761-1|LNC|glucose|glucose
C0797935|T201|OSN|14761-1|LNC|glucose|glucose
C0797935|T201|LC|14761-1|LNC|glucose|glucose
C0797936|T201|LN|14762-9|LNC|glucose|glucose
C0797936|T201|MTH_LN|14762-9|LNC|glucose|glucose
C0797936|T201|OSN|14762-9|LNC|glucose|glucose
C0797936|T201|LC|14762-9|LNC|glucose|glucose
C0797937|T201|LN|14763-7|LNC|glucose|glucose
C0797937|T201|MTH_LN|14763-7|LNC|glucose|glucose
C0797937|T201|OSN|14763-7|LNC|glucose|glucose
C0797937|T201|LC|14763-7|LNC|glucose|glucose
C0797938|T201|LN|14764-5|LNC|glucose|glucose
C0797938|T201|MTH_LN|14764-5|LNC|glucose|glucose
C0797938|T201|OSN|14764-5|LNC|glucose|glucose
C0797938|T201|LC|14764-5|LNC|glucose|glucose
C0797939|T201|LN|14765-2|LNC|glucose|glucose
C0797939|T201|MTH_LN|14765-2|LNC|glucose|glucose
C0797939|T201|OSN|14765-2|LNC|glucose|glucose
C0797939|T201|LC|14765-2|LNC|glucose|glucose
C0797940|T201|LN|14766-0|LNC|glucose|glucose
C0797940|T201|MTH_LN|14766-0|LNC|glucose|glucose
C0797940|T201|OSN|14766-0|LNC|glucose|glucose
C0797940|T201|LC|14766-0|LNC|glucose|glucose
C0797941|T201|LN|14767-8|LNC|glucose|glucose
C0797941|T201|MTH_LN|14767-8|LNC|glucose|glucose
C0797941|T201|OSN|14767-8|LNC|glucose|glucose
C0797941|T201|LC|14767-8|LNC|glucose|glucose
C0797942|T201|LN|14768-6|LNC|glucose|glucose
C0797942|T201|MTH_LN|14768-6|LNC|glucose|glucose
C0797942|T201|OSN|14768-6|LNC|glucose|glucose
C0797942|T201|LC|14768-6|LNC|glucose|glucose
C0797943|T201|LN|14769-4|LNC|glucose|glucose
C0797943|T201|MTH_LN|14769-4|LNC|glucose|glucose
C0797943|T201|OSN|14769-4|LNC|glucose|glucose
C0797943|T201|LC|14769-4|LNC|glucose|glucose
C0797944|T201|LN|14770-2|LNC|glucose|glucose
C0797944|T201|MTH_LN|14770-2|LNC|glucose|glucose
C0797944|T201|OSN|14770-2|LNC|glucose|glucose
C0797944|T201|LC|14770-2|LNC|glucose|glucose
C0797945|T201|LN|14771-0|LNC|glucose|glucose
C0797945|T201|MTH_LN|14771-0|LNC|glucose|glucose
C0797945|T201|OSN|14771-0|LNC|glucose|glucose
C0797945|T201|LC|14771-0|LNC|glucose|glucose
C0797979|T201|LN|14805-6|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0797979|T201|MTH_LN|14805-6|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0797979|T201|OSN|14805-6|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0797979|T201|LC|14805-6|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C0798036|T201|LN|14862-7|LNC|oxalate|oxalate
C0798036|T201|MTH_LN|14862-7|LNC|oxalate|oxalate
C0798036|T201|OSN|14862-7|LNC|oxalate|oxalate
C0798036|T201|LC|14862-7|LNC|oxalate|oxalate
C0798049|T201|MTH_LN|14875-9|LNC|phenylalanine metabolism|phenylalanine metabolism
C0798049|T201|LN|14875-9|LNC|phenylalanine metabolism|phenylalanine metabolism
C0798049|T201|OSN|14875-9|LNC|phenylalanine metabolism|phenylalanine metabolism
C0798049|T201|LC|14875-9|LNC|phenylalanine metabolism|phenylalanine metabolism
C0798076|T201|LN|14903-9|LNC|folate|folate
C0798076|T201|MTH_LN|14903-9|LNC|folate|folate
C0798076|T201|OSN|14903-9|LNC|folate|folate
C0798076|T201|LC|14903-9|LNC|folate|folate
C0798106|T201|LN|14933-6|LNC|uric acid|uric acid
C0798106|T201|MTH_LN|14933-6|LNC|uric acid|uric acid
C0798106|T201|OSN|14933-6|LNC|uric acid|uric acid
C0798106|T201|LC|14933-6|LNC|uric acid|uric acid
C0798106|T201|LN|14933-6|LNC|purine metabolism|purine metabolism
C0798106|T201|MTH_LN|14933-6|LNC|purine metabolism|purine metabolism
C0798106|T201|OSN|14933-6|LNC|purine metabolism|purine metabolism
C0798106|T201|LC|14933-6|LNC|purine metabolism|purine metabolism
C0798107|T201|LN|14934-4|LNC|urate|urate
C0798107|T201|MTH_LN|14934-4|LNC|urate|urate
C0798107|T201|OSN|14934-4|LNC|urate|urate
C0798107|T201|LC|14934-4|LNC|urate|urate
C0798107|T201|LN|14934-4|LNC|uric acid|uric acid
C0798107|T201|MTH_LN|14934-4|LNC|uric acid|uric acid
C0798107|T201|OSN|14934-4|LNC|uric acid|uric acid
C0798107|T201|LC|14934-4|LNC|uric acid|uric acid
C0798108|T201|LN|14935-1|LNC|urate|urate
C0798108|T201|MTH_LN|14935-1|LNC|urate|urate
C0798108|T201|OSN|14935-1|LNC|urate|urate
C0798108|T201|LC|14935-1|LNC|urate|urate
C0798108|T201|LN|14935-1|LNC|uric acid|uric acid
C0798108|T201|MTH_LN|14935-1|LNC|uric acid|uric acid
C0798108|T201|OSN|14935-1|LNC|uric acid|uric acid
C0798108|T201|LC|14935-1|LNC|uric acid|uric acid
C0798130|T201|LN|14957-5|LNC|albumin|albumin
C0798130|T201|MTH_LN|14957-5|LNC|albumin|albumin
C0798130|T201|OSN|14957-5|LNC|albumin|albumin
C0798130|T201|LC|14957-5|LNC|albumin|albumin
C0798132|T201|LN|14959-1|LNC|albumin|albumin
C0798132|T201|MTH_LN|14959-1|LNC|albumin|albumin
C0798132|T201|OSN|14959-1|LNC|albumin|albumin
C0798132|T201|LC|14959-1|LNC|albumin|albumin
C0798152|T201|LN|14979-9|LNC|coagulation disorder|coagulation disorder
C0798152|T201|LC|14979-9|LNC|coagulation disorder|coagulation disorder
C0798152|T201|MTH_LN|14979-9|LNC|coagulation disorder|coagulation disorder
C0798152|T201|OSN|14979-9|LNC|coagulation disorder|coagulation disorder
C0798152|T201|LN|14979-9|LNC|partial thromboplastin time|partial thromboplastin time
C0798152|T201|LC|14979-9|LNC|partial thromboplastin time|partial thromboplastin time
C0798152|T201|MTH_LN|14979-9|LNC|partial thromboplastin time|partial thromboplastin time
C0798152|T201|OSN|14979-9|LNC|partial thromboplastin time|partial thromboplastin time
C0798152|T201|LN|14979-9|LNC|coagulation|coagulation
C0798152|T201|LC|14979-9|LNC|coagulation|coagulation
C0798152|T201|MTH_LN|14979-9|LNC|coagulation|coagulation
C0798152|T201|OSN|14979-9|LNC|coagulation|coagulation
C0798152|T201|LN|14979-9|LNC|Coagulationities|Coagulationities
C0798152|T201|LC|14979-9|LNC|Coagulationities|Coagulationities
C0798152|T201|MTH_LN|14979-9|LNC|Coagulationities|Coagulationities
C0798152|T201|OSN|14979-9|LNC|Coagulationities|Coagulationities
C0798152|T201|LN|14979-9|LNC|coagulation studies|coagulation studies
C0798152|T201|LC|14979-9|LNC|coagulation studies|coagulation studies
C0798152|T201|MTH_LN|14979-9|LNC|coagulation studies|coagulation studies
C0798152|T201|OSN|14979-9|LNC|coagulation studies|coagulation studies
C0798152|T201|LN|14979-9|LNC|clotting|clotting
C0798152|T201|LC|14979-9|LNC|clotting|clotting
C0798152|T201|MTH_LN|14979-9|LNC|clotting|clotting
C0798152|T201|OSN|14979-9|LNC|clotting|clotting
C0798168|T201|LN|14995-5|LNC|glucose|glucose
C0798168|T201|MTH_LN|14995-5|LNC|glucose|glucose
C0798168|T201|OSN|14995-5|LNC|glucose|glucose
C0798168|T201|LC|14995-5|LNC|glucose|glucose
C0798169|T201|LN|14996-3|LNC|glucose|glucose
C0798169|T201|MTH_LN|14996-3|LNC|glucose|glucose
C0798169|T201|OSN|14996-3|LNC|glucose|glucose
C0798169|T201|LC|14996-3|LNC|glucose|glucose
C0798186|T201|LN|15013-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798186|T201|MTH_LN|15013-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798186|T201|LC|15013-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798186|T201|OSN|15013-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798186|T201|LN|15013-6|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C0798186|T201|MTH_LN|15013-6|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C0798186|T201|LC|15013-6|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C0798186|T201|OSN|15013-6|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C0798186|T201|LN|15013-6|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C0798186|T201|MTH_LN|15013-6|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C0798186|T201|LC|15013-6|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C0798186|T201|OSN|15013-6|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C0798186|T201|LN|15013-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798186|T201|MTH_LN|15013-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798186|T201|LC|15013-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798186|T201|OSN|15013-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798187|T201|LN|15014-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798187|T201|MTH_LN|15014-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798187|T201|LC|15014-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798187|T201|OSN|15014-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798187|T201|LN|15014-4|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C0798187|T201|MTH_LN|15014-4|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C0798187|T201|LC|15014-4|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C0798187|T201|OSN|15014-4|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C0798187|T201|LN|15014-4|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798187|T201|MTH_LN|15014-4|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798187|T201|LC|15014-4|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798187|T201|OSN|15014-4|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798188|T201|LN|15015-1|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798188|T201|MTH_LN|15015-1|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798188|T201|LC|15015-1|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798188|T201|OSN|15015-1|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798188|T201|LN|15015-1|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798188|T201|MTH_LN|15015-1|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798188|T201|LC|15015-1|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798188|T201|OSN|15015-1|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798188|T201|LN|15015-1|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798188|T201|MTH_LN|15015-1|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798188|T201|LC|15015-1|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798188|T201|OSN|15015-1|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798215|T201|LN|15042-5|LNC|ACTH|ACTH
C0798215|T201|MTH_LN|15042-5|LNC|ACTH|ACTH
C0798215|T201|OSN|15042-5|LNC|ACTH|ACTH
C0798215|T201|LC|15042-5|LNC|ACTH|ACTH
C0798215|T201|LN|15042-5|LNC|corticotropin|corticotropin
C0798215|T201|MTH_LN|15042-5|LNC|corticotropin|corticotropin
C0798215|T201|OSN|15042-5|LNC|corticotropin|corticotropin
C0798215|T201|LC|15042-5|LNC|corticotropin|corticotropin
C0798215|T201|LN|15042-5|LNC|adrenocorticotropin|adrenocorticotropin
C0798215|T201|MTH_LN|15042-5|LNC|adrenocorticotropin|adrenocorticotropin
C0798215|T201|OSN|15042-5|LNC|adrenocorticotropin|adrenocorticotropin
C0798215|T201|LC|15042-5|LNC|adrenocorticotropin|adrenocorticotropin
C0798239|T201|LN|15067-2|LNC|follicle stimulating|follicle stimulating
C0798239|T201|MTH_LN|15067-2|LNC|follicle stimulating|follicle stimulating
C0798239|T201|OSN|15067-2|LNC|follicle stimulating|follicle stimulating
C0798239|T201|LC|15067-2|LNC|follicle stimulating|follicle stimulating
C0798239|T201|LN|15067-2|LNC|follicle-stimulating|follicle-stimulating
C0798239|T201|MTH_LN|15067-2|LNC|follicle-stimulating|follicle-stimulating
C0798239|T201|OSN|15067-2|LNC|follicle-stimulating|follicle-stimulating
C0798239|T201|LC|15067-2|LNC|follicle-stimulating|follicle-stimulating
C0798239|T201|LN|15067-2|LNC|FSH|FSH
C0798239|T201|MTH_LN|15067-2|LNC|FSH|FSH
C0798239|T201|OSN|15067-2|LNC|FSH|FSH
C0798239|T201|LC|15067-2|LNC|FSH|FSH
C0798243|T201|LN|15071-4|LNC|galactose|galactose
C0798243|T201|MTH_LN|15071-4|LNC|galactose|galactose
C0798243|T201|OSN|15071-4|LNC|galactose|galactose
C0798243|T201|LC|15071-4|LNC|galactose|galactose
C0798246|T201|LN|15074-8|LNC|glucose|glucose
C0798246|T201|MTH_LN|15074-8|LNC|glucose|glucose
C0798246|T201|OSN|15074-8|LNC|glucose|glucose
C0798246|T201|LC|15074-8|LNC|glucose|glucose
C0798248|T201|LN|15076-3|LNC|glucose|glucose
C0798248|T201|MTH_LN|15076-3|LNC|glucose|glucose
C0798248|T201|OSN|15076-3|LNC|glucose|glucose
C0798248|T201|LC|15076-3|LNC|glucose|glucose
C0798249|T201|LN|15077-1|LNC|glucose|glucose
C0798249|T201|MTH_LN|15077-1|LNC|glucose|glucose
C0798249|T201|OSN|15077-1|LNC|glucose|glucose
C0798249|T201|LC|15077-1|LNC|glucose|glucose
C0798381|T201|LN|15210-8|LNC|Autoimmune antibody|Autoimmune antibody
C0798381|T201|MTH_LN|15210-8|LNC|Autoimmune antibody|Autoimmune antibody
C0798381|T201|OSN|15210-8|LNC|Autoimmune antibody|Autoimmune antibody
C0798381|T201|LC|15210-8|LNC|Autoimmune antibody|Autoimmune antibody
C0798517|T201|LN|15348-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798517|T201|MTH_LN|15348-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798517|T201|LC|15348-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798517|T201|OSN|15348-6|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798517|T201|LN|15348-6|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798517|T201|MTH_LN|15348-6|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798517|T201|LC|15348-6|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798517|T201|OSN|15348-6|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798517|T201|LN|15348-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798517|T201|MTH_LN|15348-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798517|T201|LC|15348-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798517|T201|OSN|15348-6|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798518|T201|LN|15349-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798518|T201|MTH_LN|15349-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798518|T201|LC|15349-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798518|T201|OSN|15349-4|LNC|Alkaline phosphatase|Alkaline phosphatase
C0798518|T201|LN|15349-4|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798518|T201|MTH_LN|15349-4|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798518|T201|LC|15349-4|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798518|T201|OSN|15349-4|LNC|alkaline phosphatasehepatic origin|alkaline phosphatasehepatic origin
C0798518|T201|LN|15349-4|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798518|T201|MTH_LN|15349-4|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798518|T201|LC|15349-4|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0798518|T201|OSN|15349-4|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C0799330|T201|LN|16165-3|LNC|glucose|glucose
C0799330|T201|MTH_LN|16165-3|LNC|glucose|glucose
C0799330|T201|OSN|16165-3|LNC|glucose|glucose
C0799330|T201|LC|16165-3|LNC|glucose|glucose
C0799331|T201|LN|16166-1|LNC|glucose|glucose
C0799331|T201|MTH_LN|16166-1|LNC|glucose|glucose
C0799331|T201|OSN|16166-1|LNC|glucose|glucose
C0799331|T201|LC|16166-1|LNC|glucose|glucose
C0799332|T201|LN|16167-9|LNC|glucose|glucose
C0799332|T201|MTH_LN|16167-9|LNC|glucose|glucose
C0799332|T201|OSN|16167-9|LNC|glucose|glucose
C0799332|T201|LC|16167-9|LNC|glucose|glucose
C0799333|T201|LN|16168-7|LNC|glucose|glucose
C0799333|T201|MTH_LN|16168-7|LNC|glucose|glucose
C0799333|T201|OSN|16168-7|LNC|glucose|glucose
C0799333|T201|LC|16168-7|LNC|glucose|glucose
C0799334|T201|LN|16169-5|LNC|glucose|glucose
C0799334|T201|MTH_LN|16169-5|LNC|glucose|glucose
C0799334|T201|OSN|16169-5|LNC|glucose|glucose
C0799334|T201|LC|16169-5|LNC|glucose|glucose
C0799335|T201|LN|16170-3|LNC|glucose|glucose
C0799335|T201|MTH_LN|16170-3|LNC|glucose|glucose
C0799335|T201|OSN|16170-3|LNC|glucose|glucose
C0799335|T201|LC|16170-3|LNC|glucose|glucose
C0799364|T201|LN|16199-2|LNC|methadone test|methadone test
C0799364|T201|LC|16199-2|LNC|methadone test|methadone test
C0799364|T201|MTH_LN|16199-2|LNC|methadone test|methadone test
C0799364|T201|OSN|16199-2|LNC|methadone test|methadone test
C0799411|T201|LN|16246-1|LNC|methadone test|methadone test
C0799411|T201|LC|16246-1|LNC|methadone test|methadone test
C0799411|T201|MTH_LN|16246-1|LNC|methadone test|methadone test
C0799411|T201|OSN|16246-1|LNC|methadone test|methadone test
C0799420|T201|LN|16255-2|LNC|troponin I|troponin I
C0799420|T201|MTH_LN|16255-2|LNC|troponin I|troponin I
C0799420|T201|OSN|16255-2|LNC|troponin I|troponin I
C0799420|T201|LC|16255-2|LNC|troponin I|troponin I
C0799525|T201|LN|16362-6|LNC|ammonia|ammonia
C0799525|T201|MTH_LN|16362-6|LNC|ammonia|ammonia
C0799525|T201|OSN|16362-6|LNC|ammonia|ammonia
C0799525|T201|LC|16362-6|LNC|ammonia|ammonia
C0799554|T201|LN|16401-2|LNC|arginine|arginine
C0799554|T201|MTH_LN|16401-2|LNC|arginine|arginine
C0799554|T201|OSN|16401-2|LNC|arginine|arginine
C0799554|T201|LC|16401-2|LNC|arginine|arginine
C0799652|T201|LN|16501-9|LNC|C-peptide|C-peptide
C0799652|T201|MTH_LN|16501-9|LNC|C-peptide|C-peptide
C0799652|T201|OSN|16501-9|LNC|C-peptide|C-peptide
C0799652|T201|LC|16501-9|LNC|C-peptide|C-peptide
C0799652|T201|LN|16501-9|LNC|C peptide|C peptide
C0799652|T201|MTH_LN|16501-9|LNC|C peptide|C peptide
C0799652|T201|OSN|16501-9|LNC|C peptide|C peptide
C0799652|T201|LC|16501-9|LNC|C peptide|C peptide
C0799653|T201|LN|16502-7|LNC|C-peptide|C-peptide
C0799653|T201|MTH_LN|16502-7|LNC|C-peptide|C-peptide
C0799653|T201|OSN|16502-7|LNC|C-peptide|C-peptide
C0799653|T201|LC|16502-7|LNC|C-peptide|C-peptide
C0799653|T201|LN|16502-7|LNC|C peptide|C peptide
C0799653|T201|MTH_LN|16502-7|LNC|C peptide|C peptide
C0799653|T201|OSN|16502-7|LNC|C peptide|C peptide
C0799653|T201|LC|16502-7|LNC|C peptide|C peptide
C0799677|T201|LN|16526-6|LNC|calcium|calcium
C0799677|T201|MTH_LN|16526-6|LNC|calcium|calcium
C0799677|T201|OSN|16526-6|LNC|calcium|calcium
C0799677|T201|LC|16526-6|LNC|calcium|calcium
C0799677|T201|LN|16526-6|LNC|calcium homeostasis|calcium homeostasis
C0799677|T201|MTH_LN|16526-6|LNC|calcium homeostasis|calcium homeostasis
C0799677|T201|OSN|16526-6|LNC|calcium homeostasis|calcium homeostasis
C0799677|T201|LC|16526-6|LNC|calcium homeostasis|calcium homeostasis
C0799700|T201|LN|16551-4|LNC|carbon dioxide|carbon dioxide
C0799700|T201|MTH_LN|16551-4|LNC|carbon dioxide|carbon dioxide
C0799700|T201|OSN|16551-4|LNC|carbon dioxide|carbon dioxide
C0799700|T201|LC|16551-4|LNC|carbon dioxide|carbon dioxide
C0799762|T201|LN|16615-7|LNC|VLDL cholesterol|VLDL cholesterol
C0799762|T201|OSN|16615-7|LNC|VLDL cholesterol|VLDL cholesterol
C0799762|T201|MTH_LN|16615-7|LNC|VLDL cholesterol|VLDL cholesterol
C0799762|T201|LC|16615-7|LNC|VLDL cholesterol|VLDL cholesterol
C0799762|T201|LN|16615-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0799762|T201|OSN|16615-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0799762|T201|MTH_LN|16615-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0799762|T201|LC|16615-7|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0799762|T201|LN|16615-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0799762|T201|OSN|16615-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0799762|T201|MTH_LN|16615-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0799762|T201|LC|16615-7|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0799763|T201|LN|16616-5|LNC|HDL cholesterol|HDL cholesterol
C0799763|T201|OSN|16616-5|LNC|HDL cholesterol|HDL cholesterol
C0799763|T201|MTH_LN|16616-5|LNC|HDL cholesterol|HDL cholesterol
C0799763|T201|LC|16616-5|LNC|HDL cholesterol|HDL cholesterol
C0799763|T201|LN|16616-5|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0799763|T201|OSN|16616-5|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0799763|T201|MTH_LN|16616-5|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0799763|T201|LC|16616-5|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0799763|T201|LN|16616-5|LNC|HDL-cholesterol|HDL-cholesterol
C0799763|T201|OSN|16616-5|LNC|HDL-cholesterol|HDL-cholesterol
C0799763|T201|MTH_LN|16616-5|LNC|HDL-cholesterol|HDL-cholesterol
C0799763|T201|LC|16616-5|LNC|HDL-cholesterol|HDL-cholesterol
C0799763|T201|LN|16616-5|LNC|high-density lipoprotein|high-density lipoprotein
C0799763|T201|OSN|16616-5|LNC|high-density lipoprotein|high-density lipoprotein
C0799763|T201|MTH_LN|16616-5|LNC|high-density lipoprotein|high-density lipoprotein
C0799763|T201|LC|16616-5|LNC|high-density lipoprotein|high-density lipoprotein
C0799763|T201|LN|16616-5|LNC|HDL|HDL
C0799763|T201|OSN|16616-5|LNC|HDL|HDL
C0799763|T201|MTH_LN|16616-5|LNC|HDL|HDL
C0799763|T201|LC|16616-5|LNC|HDL|HDL
C0799800|T201|LN|16654-6|LNC|ACTH|ACTH
C0799800|T201|OSN|16654-6|LNC|ACTH|ACTH
C0799800|T201|MTH_LN|16654-6|LNC|ACTH|ACTH
C0799800|T201|LC|16654-6|LNC|ACTH|ACTH
C0799800|T201|LN|16654-6|LNC|corticotropin|corticotropin
C0799800|T201|OSN|16654-6|LNC|corticotropin|corticotropin
C0799800|T201|MTH_LN|16654-6|LNC|corticotropin|corticotropin
C0799800|T201|LC|16654-6|LNC|corticotropin|corticotropin
C0799800|T201|LN|16654-6|LNC|adrenocorticotropin|adrenocorticotropin
C0799800|T201|OSN|16654-6|LNC|adrenocorticotropin|adrenocorticotropin
C0799800|T201|MTH_LN|16654-6|LNC|adrenocorticotropin|adrenocorticotropin
C0799800|T201|LC|16654-6|LNC|adrenocorticotropin|adrenocorticotropin
C0799801|T201|LN|16655-3|LNC|ACTH|ACTH
C0799801|T201|MTH_LN|16655-3|LNC|ACTH|ACTH
C0799801|T201|OSN|16655-3|LNC|ACTH|ACTH
C0799801|T201|LC|16655-3|LNC|ACTH|ACTH
C0799801|T201|LN|16655-3|LNC|corticotropin|corticotropin
C0799801|T201|MTH_LN|16655-3|LNC|corticotropin|corticotropin
C0799801|T201|OSN|16655-3|LNC|corticotropin|corticotropin
C0799801|T201|LC|16655-3|LNC|corticotropin|corticotropin
C0799801|T201|LN|16655-3|LNC|adrenocorticotropin|adrenocorticotropin
C0799801|T201|MTH_LN|16655-3|LNC|adrenocorticotropin|adrenocorticotropin
C0799801|T201|OSN|16655-3|LNC|adrenocorticotropin|adrenocorticotropin
C0799801|T201|LC|16655-3|LNC|adrenocorticotropin|adrenocorticotropin
C0799802|T201|LN|16656-1|LNC|ACTH|ACTH
C0799802|T201|MTH_LN|16656-1|LNC|ACTH|ACTH
C0799802|T201|OSN|16656-1|LNC|ACTH|ACTH
C0799802|T201|LC|16656-1|LNC|ACTH|ACTH
C0799802|T201|LN|16656-1|LNC|corticotropin|corticotropin
C0799802|T201|MTH_LN|16656-1|LNC|corticotropin|corticotropin
C0799802|T201|OSN|16656-1|LNC|corticotropin|corticotropin
C0799802|T201|LC|16656-1|LNC|corticotropin|corticotropin
C0799802|T201|LN|16656-1|LNC|adrenocorticotropin|adrenocorticotropin
C0799802|T201|MTH_LN|16656-1|LNC|adrenocorticotropin|adrenocorticotropin
C0799802|T201|OSN|16656-1|LNC|adrenocorticotropin|adrenocorticotropin
C0799802|T201|LC|16656-1|LNC|adrenocorticotropin|adrenocorticotropin
C0799803|T201|LN|16657-9|LNC|ACTH|ACTH
C0799803|T201|MTH_LN|16657-9|LNC|ACTH|ACTH
C0799803|T201|OSN|16657-9|LNC|ACTH|ACTH
C0799803|T201|LC|16657-9|LNC|ACTH|ACTH
C0799803|T201|LN|16657-9|LNC|corticotropin|corticotropin
C0799803|T201|MTH_LN|16657-9|LNC|corticotropin|corticotropin
C0799803|T201|OSN|16657-9|LNC|corticotropin|corticotropin
C0799803|T201|LC|16657-9|LNC|corticotropin|corticotropin
C0799803|T201|LN|16657-9|LNC|adrenocorticotropin|adrenocorticotropin
C0799803|T201|MTH_LN|16657-9|LNC|adrenocorticotropin|adrenocorticotropin
C0799803|T201|OSN|16657-9|LNC|adrenocorticotropin|adrenocorticotropin
C0799803|T201|LC|16657-9|LNC|adrenocorticotropin|adrenocorticotropin
C0799804|T201|LN|16658-7|LNC|ACTH|ACTH
C0799804|T201|MTH_LN|16658-7|LNC|ACTH|ACTH
C0799804|T201|OSN|16658-7|LNC|ACTH|ACTH
C0799804|T201|LC|16658-7|LNC|ACTH|ACTH
C0799804|T201|LN|16658-7|LNC|corticotropin|corticotropin
C0799804|T201|MTH_LN|16658-7|LNC|corticotropin|corticotropin
C0799804|T201|OSN|16658-7|LNC|corticotropin|corticotropin
C0799804|T201|LC|16658-7|LNC|corticotropin|corticotropin
C0799804|T201|LN|16658-7|LNC|adrenocorticotropin|adrenocorticotropin
C0799804|T201|MTH_LN|16658-7|LNC|adrenocorticotropin|adrenocorticotropin
C0799804|T201|OSN|16658-7|LNC|adrenocorticotropin|adrenocorticotropin
C0799804|T201|LC|16658-7|LNC|adrenocorticotropin|adrenocorticotropin
C0799805|T201|LN|16659-5|LNC|ACTH|ACTH
C0799805|T201|OSN|16659-5|LNC|ACTH|ACTH
C0799805|T201|MTH_LN|16659-5|LNC|ACTH|ACTH
C0799805|T201|LC|16659-5|LNC|ACTH|ACTH
C0799805|T201|LN|16659-5|LNC|corticotropin|corticotropin
C0799805|T201|OSN|16659-5|LNC|corticotropin|corticotropin
C0799805|T201|MTH_LN|16659-5|LNC|corticotropin|corticotropin
C0799805|T201|LC|16659-5|LNC|corticotropin|corticotropin
C0799805|T201|LN|16659-5|LNC|adrenocorticotropin|adrenocorticotropin
C0799805|T201|OSN|16659-5|LNC|adrenocorticotropin|adrenocorticotropin
C0799805|T201|MTH_LN|16659-5|LNC|adrenocorticotropin|adrenocorticotropin
C0799805|T201|LC|16659-5|LNC|adrenocorticotropin|adrenocorticotropin
C0799806|T201|LN|16660-3|LNC|ACTH|ACTH
C0799806|T201|MTH_LN|16660-3|LNC|ACTH|ACTH
C0799806|T201|OSN|16660-3|LNC|ACTH|ACTH
C0799806|T201|LC|16660-3|LNC|ACTH|ACTH
C0799806|T201|LN|16660-3|LNC|corticotropin|corticotropin
C0799806|T201|MTH_LN|16660-3|LNC|corticotropin|corticotropin
C0799806|T201|OSN|16660-3|LNC|corticotropin|corticotropin
C0799806|T201|LC|16660-3|LNC|corticotropin|corticotropin
C0799806|T201|LN|16660-3|LNC|adrenocorticotropin|adrenocorticotropin
C0799806|T201|MTH_LN|16660-3|LNC|adrenocorticotropin|adrenocorticotropin
C0799806|T201|OSN|16660-3|LNC|adrenocorticotropin|adrenocorticotropin
C0799806|T201|LC|16660-3|LNC|adrenocorticotropin|adrenocorticotropin
C0799807|T201|LN|16661-1|LNC|ACTH|ACTH
C0799807|T201|MTH_LN|16661-1|LNC|ACTH|ACTH
C0799807|T201|OSN|16661-1|LNC|ACTH|ACTH
C0799807|T201|LC|16661-1|LNC|ACTH|ACTH
C0799807|T201|LN|16661-1|LNC|corticotropin|corticotropin
C0799807|T201|MTH_LN|16661-1|LNC|corticotropin|corticotropin
C0799807|T201|OSN|16661-1|LNC|corticotropin|corticotropin
C0799807|T201|LC|16661-1|LNC|corticotropin|corticotropin
C0799807|T201|LN|16661-1|LNC|adrenocorticotropin|adrenocorticotropin
C0799807|T201|MTH_LN|16661-1|LNC|adrenocorticotropin|adrenocorticotropin
C0799807|T201|OSN|16661-1|LNC|adrenocorticotropin|adrenocorticotropin
C0799807|T201|LC|16661-1|LNC|adrenocorticotropin|adrenocorticotropin
C0799808|T201|LN|16662-9|LNC|ACTH|ACTH
C0799808|T201|MTH_LN|16662-9|LNC|ACTH|ACTH
C0799808|T201|OSN|16662-9|LNC|ACTH|ACTH
C0799808|T201|LC|16662-9|LNC|ACTH|ACTH
C0799808|T201|LN|16662-9|LNC|corticotropin|corticotropin
C0799808|T201|MTH_LN|16662-9|LNC|corticotropin|corticotropin
C0799808|T201|OSN|16662-9|LNC|corticotropin|corticotropin
C0799808|T201|LC|16662-9|LNC|corticotropin|corticotropin
C0799808|T201|LN|16662-9|LNC|adrenocorticotropin|adrenocorticotropin
C0799808|T201|MTH_LN|16662-9|LNC|adrenocorticotropin|adrenocorticotropin
C0799808|T201|OSN|16662-9|LNC|adrenocorticotropin|adrenocorticotropin
C0799808|T201|LC|16662-9|LNC|adrenocorticotropin|adrenocorticotropin
C0799809|T201|LN|16663-7|LNC|ACTH|ACTH
C0799809|T201|MTH_LN|16663-7|LNC|ACTH|ACTH
C0799809|T201|OSN|16663-7|LNC|ACTH|ACTH
C0799809|T201|LC|16663-7|LNC|ACTH|ACTH
C0799809|T201|LN|16663-7|LNC|corticotropin|corticotropin
C0799809|T201|MTH_LN|16663-7|LNC|corticotropin|corticotropin
C0799809|T201|OSN|16663-7|LNC|corticotropin|corticotropin
C0799809|T201|LC|16663-7|LNC|corticotropin|corticotropin
C0799809|T201|LN|16663-7|LNC|adrenocorticotropin|adrenocorticotropin
C0799809|T201|MTH_LN|16663-7|LNC|adrenocorticotropin|adrenocorticotropin
C0799809|T201|OSN|16663-7|LNC|adrenocorticotropin|adrenocorticotropin
C0799809|T201|LC|16663-7|LNC|adrenocorticotropin|adrenocorticotropin
C0799810|T201|LN|16664-5|LNC|ACTH|ACTH
C0799810|T201|MTH_LN|16664-5|LNC|ACTH|ACTH
C0799810|T201|OSN|16664-5|LNC|ACTH|ACTH
C0799810|T201|LC|16664-5|LNC|ACTH|ACTH
C0799810|T201|LN|16664-5|LNC|corticotropin|corticotropin
C0799810|T201|MTH_LN|16664-5|LNC|corticotropin|corticotropin
C0799810|T201|OSN|16664-5|LNC|corticotropin|corticotropin
C0799810|T201|LC|16664-5|LNC|corticotropin|corticotropin
C0799810|T201|LN|16664-5|LNC|adrenocorticotropin|adrenocorticotropin
C0799810|T201|MTH_LN|16664-5|LNC|adrenocorticotropin|adrenocorticotropin
C0799810|T201|OSN|16664-5|LNC|adrenocorticotropin|adrenocorticotropin
C0799810|T201|LC|16664-5|LNC|adrenocorticotropin|adrenocorticotropin
C0799811|T201|LN|16665-2|LNC|ACTH|ACTH
C0799811|T201|MTH_LN|16665-2|LNC|ACTH|ACTH
C0799811|T201|OSN|16665-2|LNC|ACTH|ACTH
C0799811|T201|LC|16665-2|LNC|ACTH|ACTH
C0799811|T201|LN|16665-2|LNC|corticotropin|corticotropin
C0799811|T201|MTH_LN|16665-2|LNC|corticotropin|corticotropin
C0799811|T201|OSN|16665-2|LNC|corticotropin|corticotropin
C0799811|T201|LC|16665-2|LNC|corticotropin|corticotropin
C0799811|T201|LN|16665-2|LNC|adrenocorticotropin|adrenocorticotropin
C0799811|T201|MTH_LN|16665-2|LNC|adrenocorticotropin|adrenocorticotropin
C0799811|T201|OSN|16665-2|LNC|adrenocorticotropin|adrenocorticotropin
C0799811|T201|LC|16665-2|LNC|adrenocorticotropin|adrenocorticotropin
C0799812|T201|LN|16666-0|LNC|ACTH|ACTH
C0799812|T201|MTH_LN|16666-0|LNC|ACTH|ACTH
C0799812|T201|OSN|16666-0|LNC|ACTH|ACTH
C0799812|T201|LC|16666-0|LNC|ACTH|ACTH
C0799812|T201|LN|16666-0|LNC|corticotropin|corticotropin
C0799812|T201|MTH_LN|16666-0|LNC|corticotropin|corticotropin
C0799812|T201|OSN|16666-0|LNC|corticotropin|corticotropin
C0799812|T201|LC|16666-0|LNC|corticotropin|corticotropin
C0799812|T201|LN|16666-0|LNC|adrenocorticotropin|adrenocorticotropin
C0799812|T201|MTH_LN|16666-0|LNC|adrenocorticotropin|adrenocorticotropin
C0799812|T201|OSN|16666-0|LNC|adrenocorticotropin|adrenocorticotropin
C0799812|T201|LC|16666-0|LNC|adrenocorticotropin|adrenocorticotropin
C0800048|T201|LN|16914-4|LNC|glucose|glucose
C0800048|T201|MTH_LN|16914-4|LNC|glucose|glucose
C0800048|T201|OSN|16914-4|LNC|glucose|glucose
C0800048|T201|LC|16914-4|LNC|glucose|glucose
C0800049|T201|LN|16915-1|LNC|glucose|glucose
C0800049|T201|MTH_LN|16915-1|LNC|glucose|glucose
C0800049|T201|OSN|16915-1|LNC|glucose|glucose
C0800049|T201|LC|16915-1|LNC|glucose|glucose
C0800065|T201|LN|16931-8|LNC|hematocrit|hematocrit
C0800065|T201|MTH_LN|16931-8|LNC|hematocrit|hematocrit
C0800065|T201|OSN|16931-8|LNC|hematocrit|hematocrit
C0800065|T201|LC|16931-8|LNC|hematocrit|hematocrit
C0800222|T201|LN|17094-4|LNC|luteinizing|luteinizing
C0800222|T201|MTH_LN|17094-4|LNC|luteinizing|luteinizing
C0800222|T201|OSN|17094-4|LNC|luteinizing|luteinizing
C0800222|T201|LC|17094-4|LNC|luteinizing|luteinizing
C0800222|T201|LN|17094-4|LNC|LH|LH
C0800222|T201|MTH_LN|17094-4|LNC|LH|LH
C0800222|T201|OSN|17094-4|LNC|LH|LH
C0800222|T201|LC|17094-4|LNC|LH|LH
C0800222|T201|LN|17094-4|LNC|luteinising|luteinising
C0800222|T201|MTH_LN|17094-4|LNC|luteinising|luteinising
C0800222|T201|OSN|17094-4|LNC|luteinising|luteinising
C0800222|T201|LC|17094-4|LNC|luteinising|luteinising
C0800223|T201|LN|17095-1|LNC|luteinizing|luteinizing
C0800223|T201|MTH_LN|17095-1|LNC|luteinizing|luteinizing
C0800223|T201|OSN|17095-1|LNC|luteinizing|luteinizing
C0800223|T201|LC|17095-1|LNC|luteinizing|luteinizing
C0800223|T201|LN|17095-1|LNC|LH|LH
C0800223|T201|MTH_LN|17095-1|LNC|LH|LH
C0800223|T201|OSN|17095-1|LNC|LH|LH
C0800223|T201|LC|17095-1|LNC|LH|LH
C0800223|T201|LN|17095-1|LNC|luteinising|luteinising
C0800223|T201|MTH_LN|17095-1|LNC|luteinising|luteinising
C0800223|T201|OSN|17095-1|LNC|luteinising|luteinising
C0800223|T201|LC|17095-1|LNC|luteinising|luteinising
C0800274|T201|LN|17147-0|LNC|T cell CD40 expression|T cell CD40 expression
C0800274|T201|MTH_LN|17147-0|LNC|T cell CD40 expression|T cell CD40 expression
C0800274|T201|LC|17147-0|LNC|T cell CD40 expression|T cell CD40 expression
C0800274|T201|OSN|17147-0|LNC|T cell CD40 expression|T cell CD40 expression
C0800274|T201|LN|17147-0|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0800274|T201|MTH_LN|17147-0|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0800274|T201|LC|17147-0|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0800274|T201|OSN|17147-0|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C0800280|T201|LN|17153-8|LNC|naive T|naive T
C0800280|T201|MTH_LN|17153-8|LNC|naive T|naive T
C0800280|T201|LC|17153-8|LNC|naive T|naive T
C0800280|T201|OSN|17153-8|LNC|naive T|naive T
C0800280|T201|LN|17153-8|LNC|naive T cell|naive T cell
C0800280|T201|MTH_LN|17153-8|LNC|naive T cell|naive T cell
C0800280|T201|LC|17153-8|LNC|naive T cell|naive T cell
C0800280|T201|OSN|17153-8|LNC|naive T cell|naive T cell
C0800281|T201|LN|17154-6|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0800281|T201|MTH_LN|17154-6|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0800281|T201|LC|17154-6|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0800281|T201|OSN|17154-6|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0800281|T201|LN|17154-6|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0800281|T201|MTH_LN|17154-6|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0800281|T201|LC|17154-6|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0800281|T201|OSN|17154-6|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0800281|T201|LN|17154-6|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0800281|T201|MTH_LN|17154-6|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0800281|T201|LC|17154-6|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0800281|T201|OSN|17154-6|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0800281|T201|LN|17154-6|LNC|T cell subset distribution|T cell subset distribution
C0800281|T201|MTH_LN|17154-6|LNC|T cell subset distribution|T cell subset distribution
C0800281|T201|LC|17154-6|LNC|T cell subset distribution|T cell subset distribution
C0800281|T201|OSN|17154-6|LNC|T cell subset distribution|T cell subset distribution
C0800497|T201|LN|17376-5|LNC|xenobiotic|xenobiotic
C0800497|T201|LC|17376-5|LNC|xenobiotic|xenobiotic
C0800497|T201|MTH_LN|17376-5|LNC|xenobiotic|xenobiotic
C0800497|T201|OSN|17376-5|LNC|xenobiotic|xenobiotic
C0800498|T201|LN|17377-3|LNC|xenobiotic|xenobiotic
C0800498|T201|LC|17377-3|LNC|xenobiotic|xenobiotic
C0800498|T201|MTH_LN|17377-3|LNC|xenobiotic|xenobiotic
C0800498|T201|OSN|17377-3|LNC|xenobiotic|xenobiotic
C0800792|T201|LN|17678-4|LNC|taurine|taurine
C0800792|T201|MTH_LN|17678-4|LNC|taurine|taurine
C0800792|T201|OSN|17678-4|LNC|taurine|taurine
C0800792|T201|LC|17678-4|LNC|taurine|taurine
C0800816|T201|LN|17705-5|LNC|Autoimmune antibody|Autoimmune antibody
C0800816|T201|MTH_LN|17705-5|LNC|Autoimmune antibody|Autoimmune antibody
C0800816|T201|OSN|17705-5|LNC|Autoimmune antibody|Autoimmune antibody
C0800816|T201|LC|17705-5|LNC|Autoimmune antibody|Autoimmune antibody
C0800863|T201|LN|17755-0|LNC|urate|urate
C0800863|T201|MTH_LN|17755-0|LNC|urate|urate
C0800863|T201|OSN|17755-0|LNC|urate|urate
C0800863|T201|LC|17755-0|LNC|urate|urate
C0800863|T201|LN|17755-0|LNC|uric acid|uric acid
C0800863|T201|MTH_LN|17755-0|LNC|uric acid|uric acid
C0800863|T201|OSN|17755-0|LNC|uric acid|uric acid
C0800863|T201|LC|17755-0|LNC|uric acid|uric acid
C0800864|T201|LN|17756-8|LNC|urate|urate
C0800864|T201|MTH_LN|17756-8|LNC|urate|urate
C0800864|T201|OSN|17756-8|LNC|urate|urate
C0800864|T201|LC|17756-8|LNC|urate|urate
C0800864|T201|LN|17756-8|LNC|uric acid|uric acid
C0800864|T201|MTH_LN|17756-8|LNC|uric acid|uric acid
C0800864|T201|OSN|17756-8|LNC|uric acid|uric acid
C0800864|T201|LC|17756-8|LNC|uric acid|uric acid
C0800916|T201|LN|17809-5|LNC|hematocrit|hematocrit
C0800916|T201|MTH_LN|17809-5|LNC|hematocrit|hematocrit
C0800916|T201|LC|17809-5|LNC|hematocrit|hematocrit
C0800916|T201|OSN|17809-5|LNC|hematocrit|hematocrit
C0800955|T201|LN|17848-3|LNC|reticulocytes|reticulocytes
C0800955|T201|OSN|17848-3|LNC|reticulocytes|reticulocytes
C0800955|T201|LC|17848-3|LNC|reticulocytes|reticulocytes
C0800955|T201|MTH_LN|17848-3|LNC|reticulocytes|reticulocytes
C0800955|T201|LN|17848-3|LNC|reticulocyte count|reticulocyte count
C0800955|T201|OSN|17848-3|LNC|reticulocyte count|reticulocyte count
C0800955|T201|LC|17848-3|LNC|reticulocyte count|reticulocyte count
C0800955|T201|MTH_LN|17848-3|LNC|reticulocyte count|reticulocyte count
C0800956|T201|LN|17849-1|LNC|reticulocytes|reticulocytes
C0800956|T201|MTH_LN|17849-1|LNC|reticulocytes|reticulocytes
C0800956|T201|OSN|17849-1|LNC|reticulocytes|reticulocytes
C0800956|T201|LC|17849-1|LNC|reticulocytes|reticulocytes
C0800956|T201|LN|17849-1|LNC|reticulocyte count|reticulocyte count
C0800956|T201|MTH_LN|17849-1|LNC|reticulocyte count|reticulocyte count
C0800956|T201|OSN|17849-1|LNC|reticulocyte count|reticulocyte count
C0800956|T201|LC|17849-1|LNC|reticulocyte count|reticulocyte count
C0800961|T201|LN|17854-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0800961|T201|MTH_LN|17854-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0800961|T201|OSN|17854-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0800961|T201|LC|17854-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C0800963|T201|LN|17856-6|LNC|hemoglobin|hemoglobin
C0800963|T201|MTH_LN|17856-6|LNC|hemoglobin|hemoglobin
C0800963|T201|OSN|17856-6|LNC|hemoglobin|hemoglobin
C0800963|T201|LC|17856-6|LNC|hemoglobin|hemoglobin
C0800963|T201|LN|17856-6|LNC|hemoglobin A1c|hemoglobin A1c
C0800963|T201|MTH_LN|17856-6|LNC|hemoglobin A1c|hemoglobin A1c
C0800963|T201|OSN|17856-6|LNC|hemoglobin A1c|hemoglobin A1c
C0800963|T201|LC|17856-6|LNC|hemoglobin A1c|hemoglobin A1c
C0800963|T201|LN|17856-6|LNC|glycosylated hemoglobin|glycosylated hemoglobin
C0800963|T201|MTH_LN|17856-6|LNC|glycosylated hemoglobin|glycosylated hemoglobin
C0800963|T201|OSN|17856-6|LNC|glycosylated hemoglobin|glycosylated hemoglobin
C0800963|T201|LC|17856-6|LNC|glycosylated hemoglobin|glycosylated hemoglobin
C0800963|T201|LN|17856-6|LNC|HbA1c|HbA1c
C0800963|T201|MTH_LN|17856-6|LNC|HbA1c|HbA1c
C0800963|T201|OSN|17856-6|LNC|HbA1c|HbA1c
C0800963|T201|LC|17856-6|LNC|HbA1c|HbA1c
C0800963|T201|LN|17856-6|LNC|glycated hemoglobin|glycated hemoglobin
C0800963|T201|MTH_LN|17856-6|LNC|glycated hemoglobin|glycated hemoglobin
C0800963|T201|OSN|17856-6|LNC|glycated hemoglobin|glycated hemoglobin
C0800963|T201|LC|17856-6|LNC|glycated hemoglobin|glycated hemoglobin
C0800968|T201|LN|17861-6|LNC|calcium|calcium
C0800968|T201|MTH_LN|17861-6|LNC|calcium|calcium
C0800968|T201|OSN|17861-6|LNC|calcium|calcium
C0800968|T201|LC|17861-6|LNC|calcium|calcium
C0800968|T201|LN|17861-6|LNC|calcium homeostasis|calcium homeostasis
C0800968|T201|MTH_LN|17861-6|LNC|calcium homeostasis|calcium homeostasis
C0800968|T201|OSN|17861-6|LNC|calcium homeostasis|calcium homeostasis
C0800968|T201|LC|17861-6|LNC|calcium homeostasis|calcium homeostasis
C0800969|T201|LN|17862-4|LNC|calcium|calcium
C0800969|T201|MTH_LN|17862-4|LNC|calcium|calcium
C0800969|T201|OSN|17862-4|LNC|calcium|calcium
C0800969|T201|LC|17862-4|LNC|calcium|calcium
C0800970|T201|LN|17863-2|LNC|calcium|calcium
C0800970|T201|MTH_LN|17863-2|LNC|calcium|calcium
C0800970|T201|OSN|17863-2|LNC|calcium|calcium
C0800970|T201|LC|17863-2|LNC|calcium|calcium
C0800970|T201|LN|17863-2|LNC|calcium homeostasis|calcium homeostasis
C0800970|T201|MTH_LN|17863-2|LNC|calcium homeostasis|calcium homeostasis
C0800970|T201|OSN|17863-2|LNC|calcium homeostasis|calcium homeostasis
C0800970|T201|LC|17863-2|LNC|calcium homeostasis|calcium homeostasis
C0800970|T201|MTH_LN|42567-8|LNC|calcium|calcium
C0800970|T201|OSN|42567-8|LNC|calcium|calcium
C0800970|T201|LN|42567-8|LNC|calcium|calcium
C0800970|T201|LC|42567-8|LNC|calcium|calcium
C0800970|T201|MTH_LN|42567-8|LNC|calcium homeostasis|calcium homeostasis
C0800970|T201|OSN|42567-8|LNC|calcium homeostasis|calcium homeostasis
C0800970|T201|LN|42567-8|LNC|calcium homeostasis|calcium homeostasis
C0800970|T201|LC|42567-8|LNC|calcium homeostasis|calcium homeostasis
C0800971|T201|LN|17864-0|LNC|calcium|calcium
C0800971|T201|MTH_LN|17864-0|LNC|calcium|calcium
C0800971|T201|OSN|17864-0|LNC|calcium|calcium
C0800971|T201|LC|17864-0|LNC|calcium|calcium
C0800971|T201|LN|17864-0|LNC|calcium homeostasis|calcium homeostasis
C0800971|T201|MTH_LN|17864-0|LNC|calcium homeostasis|calcium homeostasis
C0800971|T201|OSN|17864-0|LNC|calcium homeostasis|calcium homeostasis
C0800971|T201|LC|17864-0|LNC|calcium homeostasis|calcium homeostasis
C0800972|T201|LN|17865-7|LNC|glucose|glucose
C0800972|T201|MTH_LN|17865-7|LNC|glucose|glucose
C0800972|T201|OSN|17865-7|LNC|glucose|glucose
C0800972|T201|LC|17865-7|LNC|glucose|glucose
C0801239|T201|LN|18191-7|LNC|amino acid|amino acid
C0801239|T201|MTH_LN|18191-7|LNC|amino acid|amino acid
C0801239|T201|OSN|18191-7|LNC|amino acid|amino acid
C0801239|T201|LC|18191-7|LNC|amino acid|amino acid
C0801239|T201|LN|18191-7|LNC|animo acids|animo acids
C0801239|T201|MTH_LN|18191-7|LNC|animo acids|animo acids
C0801239|T201|OSN|18191-7|LNC|animo acids|animo acids
C0801239|T201|LC|18191-7|LNC|animo acids|animo acids
C0801239|T201|LN|18191-7|LNC|amino-acid findings|amino-acid findings
C0801239|T201|MTH_LN|18191-7|LNC|amino-acid findings|amino-acid findings
C0801239|T201|OSN|18191-7|LNC|amino-acid findings|amino-acid findings
C0801239|T201|LC|18191-7|LNC|amino-acid findings|amino-acid findings
C0801273|T201|LN|18227-9|LNC|glucose|glucose
C0801273|T201|MTH_LN|18227-9|LNC|glucose|glucose
C0801273|T201|OSN|18227-9|LNC|glucose|glucose
C0801273|T201|LC|18227-9|LNC|glucose|glucose
C0801274|T201|LN|18228-7|LNC|glucose-6-phosphate dehydrogenase in tissue|glucose-6-phosphate dehydrogenase in tissue
C0801274|T201|LC|18228-7|LNC|glucose-6-phosphate dehydrogenase in tissue|glucose-6-phosphate dehydrogenase in tissue
C0801274|T201|MTH_LN|18228-7|LNC|glucose-6-phosphate dehydrogenase in tissue|glucose-6-phosphate dehydrogenase in tissue
C0801274|T201|OSN|18228-7|LNC|glucose-6-phosphate dehydrogenase in tissue|glucose-6-phosphate dehydrogenase in tissue
C0801274|T201|LN|18228-7|LNC|G6PD in tissue|G6PD in tissue
C0801274|T201|LC|18228-7|LNC|G6PD in tissue|G6PD in tissue
C0801274|T201|MTH_LN|18228-7|LNC|G6PD in tissue|G6PD in tissue
C0801274|T201|OSN|18228-7|LNC|G6PD in tissue|G6PD in tissue
C0801307|T201|LN|18261-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0801307|T201|MTH_LN|18261-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0801307|T201|OSN|18261-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0801307|T201|LC|18261-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0801307|T201|LN|18261-8|LNC|LDL|LDL
C0801307|T201|MTH_LN|18261-8|LNC|LDL|LDL
C0801307|T201|OSN|18261-8|LNC|LDL|LDL
C0801307|T201|LC|18261-8|LNC|LDL|LDL
C0801307|T201|LN|18261-8|LNC|LDL cholesterol|LDL cholesterol
C0801307|T201|MTH_LN|18261-8|LNC|LDL cholesterol|LDL cholesterol
C0801307|T201|OSN|18261-8|LNC|LDL cholesterol|LDL cholesterol
C0801307|T201|LC|18261-8|LNC|LDL cholesterol|LDL cholesterol
C0801307|T201|LN|18261-8|LNC|low-density lipoprotein|low-density lipoprotein
C0801307|T201|MTH_LN|18261-8|LNC|low-density lipoprotein|low-density lipoprotein
C0801307|T201|OSN|18261-8|LNC|low-density lipoprotein|low-density lipoprotein
C0801307|T201|LC|18261-8|LNC|low-density lipoprotein|low-density lipoprotein
C0801307|T201|LN|18261-8|LNC|beta-lipoproteins|beta-lipoproteins
C0801307|T201|MTH_LN|18261-8|LNC|beta-lipoproteins|beta-lipoproteins
C0801307|T201|OSN|18261-8|LNC|beta-lipoproteins|beta-lipoproteins
C0801307|T201|LC|18261-8|LNC|beta-lipoproteins|beta-lipoproteins
C0801307|T201|LN|18261-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0801307|T201|MTH_LN|18261-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0801307|T201|OSN|18261-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0801307|T201|LC|18261-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0801307|T201|LN|18261-8|LNC|LDL-C|LDL-C
C0801307|T201|MTH_LN|18261-8|LNC|LDL-C|LDL-C
C0801307|T201|OSN|18261-8|LNC|LDL-C|LDL-C
C0801307|T201|LC|18261-8|LNC|LDL-C|LDL-C
C0801308|T201|LN|18262-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0801308|T201|MTH_LN|18262-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0801308|T201|OSN|18262-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0801308|T201|LC|18262-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0801308|T201|LN|18262-6|LNC|LDL|LDL
C0801308|T201|MTH_LN|18262-6|LNC|LDL|LDL
C0801308|T201|OSN|18262-6|LNC|LDL|LDL
C0801308|T201|LC|18262-6|LNC|LDL|LDL
C0801308|T201|LN|18262-6|LNC|LDL cholesterol|LDL cholesterol
C0801308|T201|MTH_LN|18262-6|LNC|LDL cholesterol|LDL cholesterol
C0801308|T201|OSN|18262-6|LNC|LDL cholesterol|LDL cholesterol
C0801308|T201|LC|18262-6|LNC|LDL cholesterol|LDL cholesterol
C0801308|T201|LN|18262-6|LNC|low-density lipoprotein|low-density lipoprotein
C0801308|T201|MTH_LN|18262-6|LNC|low-density lipoprotein|low-density lipoprotein
C0801308|T201|OSN|18262-6|LNC|low-density lipoprotein|low-density lipoprotein
C0801308|T201|LC|18262-6|LNC|low-density lipoprotein|low-density lipoprotein
C0801308|T201|LN|18262-6|LNC|beta-lipoproteins|beta-lipoproteins
C0801308|T201|MTH_LN|18262-6|LNC|beta-lipoproteins|beta-lipoproteins
C0801308|T201|OSN|18262-6|LNC|beta-lipoproteins|beta-lipoproteins
C0801308|T201|LC|18262-6|LNC|beta-lipoproteins|beta-lipoproteins
C0801308|T201|LN|18262-6|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0801308|T201|MTH_LN|18262-6|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0801308|T201|OSN|18262-6|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0801308|T201|LC|18262-6|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0801308|T201|LN|18262-6|LNC|LDL-C|LDL-C
C0801308|T201|MTH_LN|18262-6|LNC|LDL-C|LDL-C
C0801308|T201|OSN|18262-6|LNC|LDL-C|LDL-C
C0801308|T201|LC|18262-6|LNC|LDL-C|LDL-C
C0801309|T201|LN|18263-4|LNC|HDL cholesterol|HDL cholesterol
C0801309|T201|MTH_LN|18263-4|LNC|HDL cholesterol|HDL cholesterol
C0801309|T201|OSN|18263-4|LNC|HDL cholesterol|HDL cholesterol
C0801309|T201|LC|18263-4|LNC|HDL cholesterol|HDL cholesterol
C0801309|T201|LN|18263-4|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0801309|T201|MTH_LN|18263-4|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0801309|T201|OSN|18263-4|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0801309|T201|LC|18263-4|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C0801309|T201|LN|18263-4|LNC|HDL-cholesterol|HDL-cholesterol
C0801309|T201|MTH_LN|18263-4|LNC|HDL-cholesterol|HDL-cholesterol
C0801309|T201|OSN|18263-4|LNC|HDL-cholesterol|HDL-cholesterol
C0801309|T201|LC|18263-4|LNC|HDL-cholesterol|HDL-cholesterol
C0801309|T201|LN|18263-4|LNC|high-density lipoprotein|high-density lipoprotein
C0801309|T201|MTH_LN|18263-4|LNC|high-density lipoprotein|high-density lipoprotein
C0801309|T201|OSN|18263-4|LNC|high-density lipoprotein|high-density lipoprotein
C0801309|T201|LC|18263-4|LNC|high-density lipoprotein|high-density lipoprotein
C0801309|T201|LN|18263-4|LNC|HDL|HDL
C0801309|T201|MTH_LN|18263-4|LNC|HDL|HDL
C0801309|T201|OSN|18263-4|LNC|HDL|HDL
C0801309|T201|LC|18263-4|LNC|HDL|HDL
C0801317|T201|LN|18271-7|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0801317|T201|OSN|18271-7|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0801317|T201|MTH_LN|18271-7|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0801317|T201|LC|18271-7|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0801327|T201|LN|18281-6|LNC|calcium|calcium
C0801327|T201|MTH_LN|18281-6|LNC|calcium|calcium
C0801327|T201|OSN|18281-6|LNC|calcium|calcium
C0801327|T201|LC|18281-6|LNC|calcium|calcium
C0801327|T201|LN|18281-6|LNC|calcium homeostasis|calcium homeostasis
C0801327|T201|MTH_LN|18281-6|LNC|calcium homeostasis|calcium homeostasis
C0801327|T201|OSN|18281-6|LNC|calcium homeostasis|calcium homeostasis
C0801327|T201|LC|18281-6|LNC|calcium homeostasis|calcium homeostasis
C0801384|T201|LN|18342-6|LNC|glucose|glucose
C0801384|T201|MTH_LN|18342-6|LNC|glucose|glucose
C0801384|T201|OSN|18342-6|LNC|glucose|glucose
C0801384|T201|LC|18342-6|LNC|glucose|glucose
C0801395|T201|LN|18353-3|LNC|glucose|glucose
C0801395|T201|MTH_LN|18353-3|LNC|glucose|glucose
C0801395|T201|OSN|18353-3|LNC|glucose|glucose
C0801395|T201|LC|18353-3|LNC|glucose|glucose
C0801396|T201|LN|18354-1|LNC|glucose|glucose
C0801396|T201|MTH_LN|18354-1|LNC|glucose|glucose
C0801396|T201|OSN|18354-1|LNC|glucose|glucose
C0801396|T201|LC|18354-1|LNC|glucose|glucose
C0801421|T201|LN|18379-8|LNC|urate|urate
C0801421|T201|MTH_LN|18379-8|LNC|urate|urate
C0801421|T201|OSN|18379-8|LNC|urate|urate
C0801421|T201|LC|18379-8|LNC|urate|urate
C0801421|T201|LN|18379-8|LNC|uric acid|uric acid
C0801421|T201|MTH_LN|18379-8|LNC|uric acid|uric acid
C0801421|T201|OSN|18379-8|LNC|uric acid|uric acid
C0801421|T201|LC|18379-8|LNC|uric acid|uric acid
C0801449|T201|LN|18407-7|LNC|neutrophil count|neutrophil count
C0801449|T201|OSN|18407-7|LNC|neutrophil count|neutrophil count
C0801449|T201|MTH_LN|18407-7|LNC|neutrophil count|neutrophil count
C0801449|T201|LC|18407-7|LNC|neutrophil count|neutrophil count
C0801449|T201|LN|18407-7|LNC|cytology|cytology
C0801449|T201|OSN|18407-7|LNC|cytology|cytology
C0801449|T201|MTH_LN|18407-7|LNC|cytology|cytology
C0801449|T201|LC|18407-7|LNC|cytology|cytology
C0801478|T201|LN|18436-6|LNC|acylcarnitine|acylcarnitine
C0801478|T201|OSN|18436-6|LNC|acylcarnitine|acylcarnitine
C0801478|T201|MTH_LN|18436-6|LNC|acylcarnitine|acylcarnitine
C0801478|T201|LC|18436-6|LNC|acylcarnitine|acylcarnitine
C0801529|T201|LN|18488-7|LNC|calcium|calcium
C0801529|T201|MTH_LN|18488-7|LNC|calcium|calcium
C0801529|T201|OSN|18488-7|LNC|calcium|calcium
C0801529|T201|LC|18488-7|LNC|calcium|calcium
C0802027|T201|LN|19079-3|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0802027|T201|MTH_LN|19079-3|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0802027|T201|LC|19079-3|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0802027|T201|OSN|19079-3|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C0802027|T201|LN|19079-3|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0802027|T201|MTH_LN|19079-3|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0802027|T201|LC|19079-3|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0802027|T201|OSN|19079-3|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C0802027|T201|LN|19079-3|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0802027|T201|MTH_LN|19079-3|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0802027|T201|LC|19079-3|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0802027|T201|OSN|19079-3|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C0802027|T201|LN|19079-3|LNC|T cell subset distribution|T cell subset distribution
C0802027|T201|MTH_LN|19079-3|LNC|T cell subset distribution|T cell subset distribution
C0802027|T201|LC|19079-3|LNC|T cell subset distribution|T cell subset distribution
C0802027|T201|OSN|19079-3|LNC|T cell subset distribution|T cell subset distribution
C0802050|T201|LN|19113-0|LNC|IgE|IgE
C0802050|T201|LC|19113-0|LNC|IgE|IgE
C0802050|T201|OSN|19113-0|LNC|IgE|IgE
C0802050|T201|MTH_LN|19113-0|LNC|IgE|IgE
C0802050|T201|LN|19113-0|LNC|immunoglobulin E|immunoglobulin E
C0802050|T201|LC|19113-0|LNC|immunoglobulin E|immunoglobulin E
C0802050|T201|OSN|19113-0|LNC|immunoglobulin E|immunoglobulin E
C0802050|T201|MTH_LN|19113-0|LNC|immunoglobulin E|immunoglobulin E
C0802053|T201|LC|19123-9|LNC|magnesium|magnesium
C0802053|T201|MTH_LN|19123-9|LNC|magnesium|magnesium
C0802053|T201|LN|19123-9|LNC|magnesium|magnesium
C0802053|T201|OSN|19123-9|LNC|magnesium|magnesium
C0802053|T201|LC|19123-9|LNC|magnesium metabolism|magnesium metabolism
C0802053|T201|MTH_LN|19123-9|LNC|magnesium metabolism|magnesium metabolism
C0802053|T201|LN|19123-9|LNC|magnesium metabolism|magnesium metabolism
C0802053|T201|OSN|19123-9|LNC|magnesium metabolism|magnesium metabolism
C0802053|T201|LC|19123-9|LNC|magnesium homeostasis|magnesium homeostasis
C0802053|T201|MTH_LN|19123-9|LNC|magnesium homeostasis|magnesium homeostasis
C0802053|T201|LN|19123-9|LNC|magnesium homeostasis|magnesium homeostasis
C0802053|T201|OSN|19123-9|LNC|magnesium homeostasis|magnesium homeostasis
C0802054|T201|LC|19124-7|LNC|magnesium|magnesium
C0802054|T201|MTH_LN|19124-7|LNC|magnesium|magnesium
C0802054|T201|OSN|19124-7|LNC|magnesium|magnesium
C0802054|T201|LN|19124-7|LNC|magnesium|magnesium
C0802082|T201|LN|19161-9|LNC|urobilinogen|urobilinogen
C0802082|T201|MTH_LN|19161-9|LNC|urobilinogen|urobilinogen
C0802082|T201|OSN|19161-9|LNC|urobilinogen|urobilinogen
C0802082|T201|LC|19161-9|LNC|urobilinogen|urobilinogen
C0802097|T201|LN|19176-7|LNC|alpha-fetoprotein|alpha-fetoprotein
C0802097|T201|MTH_LN|19176-7|LNC|alpha-fetoprotein|alpha-fetoprotein
C0802097|T201|OSN|19176-7|LNC|alpha-fetoprotein|alpha-fetoprotein
C0802097|T201|LC|19176-7|LNC|alpha-fetoprotein|alpha-fetoprotein
C0802097|T201|LN|19176-7|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0802097|T201|MTH_LN|19176-7|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0802097|T201|OSN|19176-7|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0802097|T201|LC|19176-7|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0802097|T201|LN|19176-7|LNC|alpha fetoprotein|alpha fetoprotein
C0802097|T201|MTH_LN|19176-7|LNC|alpha fetoprotein|alpha fetoprotein
C0802097|T201|OSN|19176-7|LNC|alpha fetoprotein|alpha fetoprotein
C0802097|T201|LC|19176-7|LNC|alpha fetoprotein|alpha fetoprotein
C0802098|T201|LN|19177-5|LNC|alpha-fetoprotein|alpha-fetoprotein
C0802098|T201|OSN|19177-5|LNC|alpha-fetoprotein|alpha-fetoprotein
C0802098|T201|MTH_LN|19177-5|LNC|alpha-fetoprotein|alpha-fetoprotein
C0802098|T201|LC|19177-5|LNC|alpha-fetoprotein|alpha-fetoprotein
C0802098|T201|LN|19177-5|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0802098|T201|OSN|19177-5|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0802098|T201|MTH_LN|19177-5|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0802098|T201|LC|19177-5|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C0802098|T201|LN|19177-5|LNC|alpha fetoprotein|alpha fetoprotein
C0802098|T201|OSN|19177-5|LNC|alpha fetoprotein|alpha fetoprotein
C0802098|T201|MTH_LN|19177-5|LNC|alpha fetoprotein|alpha fetoprotein
C0802098|T201|LC|19177-5|LNC|alpha fetoprotein|alpha fetoprotein
C0802144|T201|LN|19239-3|LNC|lactate|lactate
C0802144|T201|MTH_LN|19239-3|LNC|lactate|lactate
C0802144|T201|OSN|19239-3|LNC|lactate|lactate
C0802144|T201|LC|19239-3|LNC|lactate|lactate
C0802145|T201|LN|19240-1|LNC|lactate|lactate
C0802145|T201|MTH_LN|19240-1|LNC|lactate|lactate
C0802145|T201|OSN|19240-1|LNC|lactate|lactate
C0802145|T201|LC|19240-1|LNC|lactate|lactate
C0802146|T201|LN|19242-7|LNC|ACTH|ACTH
C0802146|T201|MTH_LN|19242-7|LNC|ACTH|ACTH
C0802146|T201|OSN|19242-7|LNC|ACTH|ACTH
C0802146|T201|LC|19242-7|LNC|ACTH|ACTH
C0802146|T201|LN|19242-7|LNC|corticotropin|corticotropin
C0802146|T201|MTH_LN|19242-7|LNC|corticotropin|corticotropin
C0802146|T201|OSN|19242-7|LNC|corticotropin|corticotropin
C0802146|T201|LC|19242-7|LNC|corticotropin|corticotropin
C0802146|T201|LN|19242-7|LNC|adrenocorticotropin|adrenocorticotropin
C0802146|T201|MTH_LN|19242-7|LNC|adrenocorticotropin|adrenocorticotropin
C0802146|T201|OSN|19242-7|LNC|adrenocorticotropin|adrenocorticotropin
C0802146|T201|LC|19242-7|LNC|adrenocorticotropin|adrenocorticotropin
C0802425|T201|LN|19550-3|LNC|methadone test|methadone test
C0802425|T201|MTH_LN|19550-3|LNC|methadone test|methadone test
C0802425|T201|OSN|19550-3|LNC|methadone test|methadone test
C0802425|T201|LC|19550-3|LNC|methadone test|methadone test
C0802426|T201|LN|19552-9|LNC|methadone test|methadone test
C0802426|T201|MTH_LN|19552-9|LNC|methadone test|methadone test
C0802426|T201|OSN|19552-9|LNC|methadone test|methadone test
C0802426|T201|LC|19552-9|LNC|methadone test|methadone test
C0802427|T201|LN|19553-7|LNC|methadone test|methadone test
C0802427|T201|LC|19553-7|LNC|methadone test|methadone test
C0802427|T201|MTH_LN|19553-7|LNC|methadone test|methadone test
C0802427|T201|OSN|19553-7|LNC|methadone test|methadone test
C0803220|T201|LN|20405-7|LNC|urobilinogen|urobilinogen
C0803220|T201|MTH_LN|20405-7|LNC|urobilinogen|urobilinogen
C0803220|T201|OSN|20405-7|LNC|urobilinogen|urobilinogen
C0803220|T201|LC|20405-7|LNC|urobilinogen|urobilinogen
C0803223|T201|LN|20408-1|LNC|neutrophil count|neutrophil count
C0803223|T201|OSN|20408-1|LNC|neutrophil count|neutrophil count
C0803223|T201|MTH_LN|20408-1|LNC|neutrophil count|neutrophil count
C0803223|T201|LC|20408-1|LNC|neutrophil count|neutrophil count
C0803223|T201|LN|20408-1|LNC|cytology|cytology
C0803223|T201|OSN|20408-1|LNC|cytology|cytology
C0803223|T201|MTH_LN|20408-1|LNC|cytology|cytology
C0803223|T201|LC|20408-1|LNC|cytology|cytology
// C0803224|T201|LN|20409-9|LNC||
// C0803224|T201|OSN|20409-9|LNC||
// C0803224|T201|MTH_LN|20409-9|LNC||
// C0803224|T201|LC|20409-9|LNC||
C0803224|T201|LN|20409-9|LNC|occult|occult
C0803224|T201|OSN|20409-9|LNC|occult|occult
C0803224|T201|MTH_LN|20409-9|LNC|occult|occult
C0803224|T201|LC|20409-9|LNC|occult|occult
C0803234|T201|LN|20419-8|LNC|luteinizing|luteinizing
C0803234|T201|MTH_LN|20419-8|LNC|luteinizing|luteinizing
C0803234|T201|OSN|20419-8|LNC|luteinizing|luteinizing
C0803234|T201|LC|20419-8|LNC|luteinizing|luteinizing
C0803234|T201|LN|20419-8|LNC|LH|LH
C0803234|T201|MTH_LN|20419-8|LNC|LH|LH
C0803234|T201|OSN|20419-8|LNC|LH|LH
C0803234|T201|LC|20419-8|LNC|LH|LH
C0803234|T201|LN|20419-8|LNC|luteinising|luteinising
C0803234|T201|MTH_LN|20419-8|LNC|luteinising|luteinising
C0803234|T201|OSN|20419-8|LNC|luteinising|luteinising
C0803234|T201|LC|20419-8|LNC|luteinising|luteinising
C0803242|T201|LN|20427-1|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0803242|T201|MTH_LN|20427-1|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0803242|T201|OSN|20427-1|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0803242|T201|LC|20427-1|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C0803251|T201|LN|20436-2|LNC|glucose|glucose
C0803251|T201|MTH_LN|20436-2|LNC|glucose|glucose
C0803251|T201|OSN|20436-2|LNC|glucose|glucose
C0803251|T201|LC|20436-2|LNC|glucose|glucose
C0803252|T201|LN|20437-0|LNC|glucose|glucose
C0803252|T201|MTH_LN|20437-0|LNC|glucose|glucose
C0803252|T201|OSN|20437-0|LNC|glucose|glucose
C0803252|T201|LC|20437-0|LNC|glucose|glucose
C0803253|T201|LN|20438-8|LNC|glucose|glucose
C0803253|T201|MTH_LN|20438-8|LNC|glucose|glucose
C0803253|T201|OSN|20438-8|LNC|glucose|glucose
C0803253|T201|LC|20438-8|LNC|glucose|glucose
C0803254|T201|LN|20439-6|LNC|glucose|glucose
C0803254|T201|MTH_LN|20439-6|LNC|glucose|glucose
C0803254|T201|OSN|20439-6|LNC|glucose|glucose
C0803254|T201|LC|20439-6|LNC|glucose|glucose
C0803255|T201|LN|20440-4|LNC|glucose|glucose
C0803255|T201|OSN|20440-4|LNC|glucose|glucose
C0803255|T201|MTH_LN|20440-4|LNC|glucose|glucose
C0803255|T201|LC|20440-4|LNC|glucose|glucose
C0803256|T201|LN|20441-2|LNC|glucose|glucose
C0803256|T201|MTH_LN|20441-2|LNC|glucose|glucose
C0803256|T201|OSN|20441-2|LNC|glucose|glucose
C0803256|T201|LC|20441-2|LNC|glucose|glucose
C0803262|T201|LN|20448-7|LNC|insulin|insulin
C0803262|T201|MTH_LN|20448-7|LNC|insulin|insulin
C0803262|T201|OSN|20448-7|LNC|insulin|insulin
C0803262|T201|LC|20448-7|LNC|insulin|insulin
C0803268|T201|LN|20454-5|LNC|Protein|Protein
C0803268|T201|MTH_LN|20454-5|LNC|Protein|Protein
C0803268|T201|OSN|20454-5|LNC|Protein|Protein
C0803268|T201|LC|20454-5|LNC|Protein|Protein
C0803269|T201|LN|20455-2|LNC|neutrophil count|neutrophil count
C0803269|T201|MTH_LN|20455-2|LNC|neutrophil count|neutrophil count
C0803269|T201|OSN|20455-2|LNC|neutrophil count|neutrophil count
C0803269|T201|LC|20455-2|LNC|neutrophil count|neutrophil count
C0803269|T201|LN|20455-2|LNC|cytology|cytology
C0803269|T201|MTH_LN|20455-2|LNC|cytology|cytology
C0803269|T201|OSN|20455-2|LNC|cytology|cytology
C0803269|T201|LC|20455-2|LNC|cytology|cytology
C0803374|T201|LN|20565-8|LNC|carbon dioxide|carbon dioxide
C0803374|T201|MTH_LN|20565-8|LNC|carbon dioxide|carbon dioxide
C0803374|T201|OSN|20565-8|LNC|carbon dioxide|carbon dioxide
C0803374|T201|LC|20565-8|LNC|carbon dioxide|carbon dioxide
C0803376|T201|LN|20567-4|LNC|ferritin|ferritin
C0803376|T201|OSN|20567-4|LNC|ferritin|ferritin
C0803376|T201|MTH_LN|20567-4|LNC|ferritin|ferritin
C0803376|T201|LC|20567-4|LNC|ferritin|ferritin
C0803378|T201|LN|20569-0|LNC|creatine phosphokinase|creatine phosphokinase
C0803378|T201|MTH_LN|20569-0|LNC|creatine phosphokinase|creatine phosphokinase
C0803378|T201|LC|20569-0|LNC|creatine phosphokinase|creatine phosphokinase
C0803378|T201|OSN|20569-0|LNC|creatine phosphokinase|creatine phosphokinase
C0803378|T201|LN|20569-0|LNC|CPK|CPK
C0803378|T201|MTH_LN|20569-0|LNC|CPK|CPK
C0803378|T201|LC|20569-0|LNC|CPK|CPK
C0803378|T201|OSN|20569-0|LNC|CPK|CPK
C0803378|T201|LN|20569-0|LNC|creatine kinase|creatine kinase
C0803378|T201|MTH_LN|20569-0|LNC|creatine kinase|creatine kinase
C0803378|T201|LC|20569-0|LNC|creatine kinase|creatine kinase
C0803378|T201|OSN|20569-0|LNC|creatine kinase|creatine kinase
C0803378|T201|LN|20569-0|LNC|CK|CK
C0803378|T201|MTH_LN|20569-0|LNC|CK|CK
C0803378|T201|LC|20569-0|LNC|CK|CK
C0803378|T201|OSN|20569-0|LNC|CK|CK
C0803379|T201|LN|20570-8|LNC|hematocrit|hematocrit
C0803379|T201|MTH_LN|20570-8|LNC|hematocrit|hematocrit
C0803379|T201|LC|20570-8|LNC|hematocrit|hematocrit
C0803379|T201|OSN|20570-8|LNC|hematocrit|hematocrit
C0803381|T201|LN|20572-4|LNC|hemoglobin|hemoglobin
C0803381|T201|MTH_LN|20572-4|LNC|hemoglobin|hemoglobin
C0803381|T201|LC|20572-4|LNC|hemoglobin|hemoglobin
C0803381|T201|OSN|20572-4|LNC|hemoglobin|hemoglobin
C0803381|T201|LN|20572-4|LNC|hemoglobin A|hemoglobin A
C0803381|T201|MTH_LN|20572-4|LNC|hemoglobin A|hemoglobin A
C0803381|T201|LC|20572-4|LNC|hemoglobin A|hemoglobin A
C0803381|T201|OSN|20572-4|LNC|hemoglobin A|hemoglobin A
C0803437|T201|LN|20633-4|LNC|histidine metabolism|histidine metabolism
C0803437|T201|MTH_LN|20633-4|LNC|histidine metabolism|histidine metabolism
C0803437|T201|OSN|20633-4|LNC|histidine metabolism|histidine metabolism
C0803437|T201|LC|20633-4|LNC|histidine metabolism|histidine metabolism
C0803439|T201|LN|20635-9|LNC|histidine metabolism|histidine metabolism
C0803439|T201|MTH_LN|20635-9|LNC|histidine metabolism|histidine metabolism
C0803439|T201|OSN|20635-9|LNC|histidine metabolism|histidine metabolism
C0803439|T201|LC|20635-9|LNC|histidine metabolism|histidine metabolism
C0803440|T201|LN|20636-7|LNC|alanine|alanine
C0803440|T201|MTH_LN|20636-7|LNC|alanine|alanine
C0803440|T201|OSN|20636-7|LNC|alanine|alanine
C0803440|T201|LC|20636-7|LNC|alanine|alanine
C0803440|T201|LN|20636-7|LNC|alanine metabolism|alanine metabolism
C0803440|T201|MTH_LN|20636-7|LNC|alanine metabolism|alanine metabolism
C0803440|T201|OSN|20636-7|LNC|alanine metabolism|alanine metabolism
C0803440|T201|LC|20636-7|LNC|alanine metabolism|alanine metabolism
C0803441|T201|LN|20637-5|LNC|arginine metabolism|arginine metabolism
C0803441|T201|MTH_LN|20637-5|LNC|arginine metabolism|arginine metabolism
C0803441|T201|OSN|20637-5|LNC|arginine metabolism|arginine metabolism
C0803441|T201|LC|20637-5|LNC|arginine metabolism|arginine metabolism
C0803441|T201|LN|20637-5|LNC|arginine|arginine
C0803441|T201|MTH_LN|20637-5|LNC|arginine|arginine
C0803441|T201|OSN|20637-5|LNC|arginine|arginine
C0803441|T201|LC|20637-5|LNC|arginine|arginine
C0803444|T201|LN|20640-9|LNC|citrulline|citrulline
C0803444|T201|MTH_LN|20640-9|LNC|citrulline|citrulline
C0803444|T201|OSN|20640-9|LNC|citrulline|citrulline
C0803444|T201|LC|20640-9|LNC|citrulline|citrulline
C0803444|T201|LN|20640-9|LNC|citrulline metabolism|citrulline metabolism
C0803444|T201|MTH_LN|20640-9|LNC|citrulline metabolism|citrulline metabolism
C0803444|T201|OSN|20640-9|LNC|citrulline metabolism|citrulline metabolism
C0803444|T201|LC|20640-9|LNC|citrulline metabolism|citrulline metabolism
C0803447|T201|LN|20643-3|LNC|glutamine|glutamine
C0803447|T201|MTH_LN|20643-3|LNC|glutamine|glutamine
C0803447|T201|OSN|20643-3|LNC|glutamine|glutamine
C0803447|T201|LC|20643-3|LNC|glutamine|glutamine
C0803447|T201|LN|20643-3|LNC|glutamine metabolism|glutamine metabolism
C0803447|T201|MTH_LN|20643-3|LNC|glutamine metabolism|glutamine metabolism
C0803447|T201|OSN|20643-3|LNC|glutamine metabolism|glutamine metabolism
C0803447|T201|LC|20643-3|LNC|glutamine metabolism|glutamine metabolism
C0803448|T201|LN|20644-1|LNC|glycine|glycine
C0803448|T201|MTH_LN|20644-1|LNC|glycine|glycine
C0803448|T201|OSN|20644-1|LNC|glycine|glycine
C0803448|T201|LC|20644-1|LNC|glycine|glycine
C0803448|T201|LN|20644-1|LNC|glycine metabolism|glycine metabolism
C0803448|T201|MTH_LN|20644-1|LNC|glycine metabolism|glycine metabolism
C0803448|T201|OSN|20644-1|LNC|glycine metabolism|glycine metabolism
C0803448|T201|LC|20644-1|LNC|glycine metabolism|glycine metabolism
C0803449|T201|LN|20645-8|LNC|histidine|histidine
C0803449|T201|MTH_LN|20645-8|LNC|histidine|histidine
C0803449|T201|OSN|20645-8|LNC|histidine|histidine
C0803449|T201|LC|20645-8|LNC|histidine|histidine
C0803449|T201|LN|20645-8|LNC|histidine metabolism|histidine metabolism
C0803449|T201|MTH_LN|20645-8|LNC|histidine metabolism|histidine metabolism
C0803449|T201|OSN|20645-8|LNC|histidine metabolism|histidine metabolism
C0803449|T201|LC|20645-8|LNC|histidine metabolism|histidine metabolism
C0803451|T201|LN|20647-4|LNC|hydroxyproline|hydroxyproline
C0803451|T201|MTH_LN|20647-4|LNC|hydroxyproline|hydroxyproline
C0803451|T201|OSN|20647-4|LNC|hydroxyproline|hydroxyproline
C0803451|T201|LC|20647-4|LNC|hydroxyproline|hydroxyproline
C0803451|T201|LN|20647-4|LNC|proline metabolism|proline metabolism
C0803451|T201|MTH_LN|20647-4|LNC|proline metabolism|proline metabolism
C0803451|T201|OSN|20647-4|LNC|proline metabolism|proline metabolism
C0803451|T201|LC|20647-4|LNC|proline metabolism|proline metabolism
C0803452|T201|LN|20648-2|LNC|isoleucine|isoleucine
C0803452|T201|MTH_LN|20648-2|LNC|isoleucine|isoleucine
C0803452|T201|OSN|20648-2|LNC|isoleucine|isoleucine
C0803452|T201|LC|20648-2|LNC|isoleucine|isoleucine
C0803452|T201|LN|20648-2|LNC|isoleucine metabolism|isoleucine metabolism
C0803452|T201|MTH_LN|20648-2|LNC|isoleucine metabolism|isoleucine metabolism
C0803452|T201|OSN|20648-2|LNC|isoleucine metabolism|isoleucine metabolism
C0803452|T201|LC|20648-2|LNC|isoleucine metabolism|isoleucine metabolism
C0803453|T201|LN|20649-0|LNC|leucine|leucine
C0803453|T201|MTH_LN|20649-0|LNC|leucine|leucine
C0803453|T201|OSN|20649-0|LNC|leucine|leucine
C0803453|T201|LC|20649-0|LNC|leucine|leucine
C0803453|T201|LN|20649-0|LNC|leucine metabolism|leucine metabolism
C0803453|T201|MTH_LN|20649-0|LNC|leucine metabolism|leucine metabolism
C0803453|T201|OSN|20649-0|LNC|leucine metabolism|leucine metabolism
C0803453|T201|LC|20649-0|LNC|leucine metabolism|leucine metabolism
C0803454|T201|LN|20650-8|LNC|lysine|lysine
C0803454|T201|MTH_LN|20650-8|LNC|lysine|lysine
C0803454|T201|OSN|20650-8|LNC|lysine|lysine
C0803454|T201|LC|20650-8|LNC|lysine|lysine
C0803454|T201|LN|20650-8|LNC|lysine metabolism|lysine metabolism
C0803454|T201|MTH_LN|20650-8|LNC|lysine metabolism|lysine metabolism
C0803454|T201|OSN|20650-8|LNC|lysine metabolism|lysine metabolism
C0803454|T201|LC|20650-8|LNC|lysine metabolism|lysine metabolism
C0803455|T201|LN|20651-6|LNC|methionine|methionine
C0803455|T201|MTH_LN|20651-6|LNC|methionine|methionine
C0803455|T201|OSN|20651-6|LNC|methionine|methionine
C0803455|T201|LC|20651-6|LNC|methionine|methionine
C0803455|T201|LN|20651-6|LNC|methionine metabolism|methionine metabolism
C0803455|T201|MTH_LN|20651-6|LNC|methionine metabolism|methionine metabolism
C0803455|T201|OSN|20651-6|LNC|methionine metabolism|methionine metabolism
C0803455|T201|LC|20651-6|LNC|methionine metabolism|methionine metabolism
C0803456|T201|LN|20652-4|LNC|ornithine|ornithine
C0803456|T201|MTH_LN|20652-4|LNC|ornithine|ornithine
C0803456|T201|OSN|20652-4|LNC|ornithine|ornithine
C0803456|T201|LC|20652-4|LNC|ornithine|ornithine
C0803456|T201|LN|20652-4|LNC|ornithine metabolism|ornithine metabolism
C0803456|T201|MTH_LN|20652-4|LNC|ornithine metabolism|ornithine metabolism
C0803456|T201|OSN|20652-4|LNC|ornithine metabolism|ornithine metabolism
C0803456|T201|LC|20652-4|LNC|ornithine metabolism|ornithine metabolism
C0803458|T201|LN|20655-7|LNC|proline metabolism|proline metabolism
C0803458|T201|MTH_LN|20655-7|LNC|proline metabolism|proline metabolism
C0803458|T201|OSN|20655-7|LNC|proline metabolism|proline metabolism
C0803458|T201|LC|20655-7|LNC|proline metabolism|proline metabolism
C0803459|T201|LN|20656-5|LNC|serine|serine
C0803459|T201|MTH_LN|20656-5|LNC|serine|serine
C0803459|T201|OSN|20656-5|LNC|serine|serine
C0803459|T201|LC|20656-5|LNC|serine|serine
C0803459|T201|LN|20656-5|LNC|serine metabolism|serine metabolism
C0803459|T201|MTH_LN|20656-5|LNC|serine metabolism|serine metabolism
C0803459|T201|OSN|20656-5|LNC|serine metabolism|serine metabolism
C0803459|T201|LC|20656-5|LNC|serine metabolism|serine metabolism
C0803461|T201|LN|20658-1|LNC|threonine|threonine
C0803461|T201|MTH_LN|20658-1|LNC|threonine|threonine
C0803461|T201|OSN|20658-1|LNC|threonine|threonine
C0803461|T201|LC|20658-1|LNC|threonine|threonine
C0803461|T201|LN|20658-1|LNC|threonine metabolism|threonine metabolism
C0803461|T201|MTH_LN|20658-1|LNC|threonine metabolism|threonine metabolism
C0803461|T201|OSN|20658-1|LNC|threonine metabolism|threonine metabolism
C0803461|T201|LC|20658-1|LNC|threonine metabolism|threonine metabolism
C0803463|T201|LN|20660-7|LNC|tyrosine|tyrosine
C0803463|T201|MTH_LN|20660-7|LNC|tyrosine|tyrosine
C0803463|T201|OSN|20660-7|LNC|tyrosine|tyrosine
C0803463|T201|LC|20660-7|LNC|tyrosine|tyrosine
C0803463|T201|LN|20660-7|LNC|tyrosine metabolism|tyrosine metabolism
C0803463|T201|MTH_LN|20660-7|LNC|tyrosine metabolism|tyrosine metabolism
C0803463|T201|OSN|20660-7|LNC|tyrosine metabolism|tyrosine metabolism
C0803463|T201|LC|20660-7|LNC|tyrosine metabolism|tyrosine metabolism
C0803464|T201|LN|20661-5|LNC|valine|valine
C0803464|T201|MTH_LN|20661-5|LNC|valine|valine
C0803464|T201|OSN|20661-5|LNC|valine|valine
C0803464|T201|LC|20661-5|LNC|valine|valine
C0803464|T201|LN|20661-5|LNC|valine metabolism|valine metabolism
C0803464|T201|MTH_LN|20661-5|LNC|valine metabolism|valine metabolism
C0803464|T201|OSN|20661-5|LNC|valine metabolism|valine metabolism
C0803464|T201|LC|20661-5|LNC|valine metabolism|valine metabolism
C0803484|T201|LN|20684-7|LNC|ammonia|ammonia
C0803484|T201|MTH_LN|20684-7|LNC|ammonia|ammonia
C0803484|T201|OSN|20684-7|LNC|ammonia|ammonia
C0803484|T201|LC|20684-7|LNC|ammonia|ammonia
C0803797|T201|LN|21000-5|LNC|red|red
C0803797|T201|MTH_LN|21000-5|LNC|red|red
C0803797|T201|OSN|21000-5|LNC|red|red
C0803797|T201|LC|21000-5|LNC|red|red
C0803797|T201|LN|21000-5|LNC|erythrocytes|erythrocytes
C0803797|T201|MTH_LN|21000-5|LNC|erythrocytes|erythrocytes
C0803797|T201|OSN|21000-5|LNC|erythrocytes|erythrocytes
C0803797|T201|LC|21000-5|LNC|erythrocytes|erythrocytes
C0803797|T201|LN|21000-5|LNC|erythrocyte morphology|erythrocyte morphology
C0803797|T201|MTH_LN|21000-5|LNC|erythrocyte morphology|erythrocyte morphology
C0803797|T201|OSN|21000-5|LNC|erythrocyte morphology|erythrocyte morphology
C0803797|T201|LC|21000-5|LNC|erythrocyte morphology|erythrocyte morphology
C0803797|T201|LN|21000-5|LNC|erythroid lineage cell|erythroid lineage cell
C0803797|T201|MTH_LN|21000-5|LNC|erythroid lineage cell|erythroid lineage cell
C0803797|T201|OSN|21000-5|LNC|erythroid lineage cell|erythroid lineage cell
C0803797|T201|LC|21000-5|LNC|erythroid lineage cell|erythroid lineage cell
C0803801|T201|MTH_LN|21004-7|LNC|glucose tolerance|glucose tolerance
C0803801|T201|LN|21004-7|LNC|glucose tolerance|glucose tolerance
C0803801|T201|OSN|21004-7|LNC|glucose tolerance|glucose tolerance
C0803801|T201|LC|21004-7|LNC|glucose tolerance|glucose tolerance
C0804013|T201|LN|21219-1|LNC|copper|copper
C0804013|T201|MTH_LN|21219-1|LNC|copper|copper
C0804013|T201|OSN|21219-1|LNC|copper|copper
C0804013|T201|LC|21219-1|LNC|copper|copper
C0804058|T201|LN|21264-7|LNC|estriol|estriol
C0804058|T201|LC|21264-7|LNC|estriol|estriol
C0804058|T201|MTH_LN|21264-7|LNC|estriol|estriol
C0804058|T201|OSN|21264-7|LNC|estriol|estriol
C0804099|T201|LN|21305-8|LNC|glucose|glucose
C0804099|T201|MTH_LN|21305-8|LNC|glucose|glucose
C0804099|T201|OSN|21305-8|LNC|glucose|glucose
C0804099|T201|LC|21305-8|LNC|glucose|glucose
C0804100|T201|LN|21306-6|LNC|glucose|glucose
C0804100|T201|MTH_LN|21306-6|LNC|glucose|glucose
C0804100|T201|OSN|21306-6|LNC|glucose|glucose
C0804100|T201|LC|21306-6|LNC|glucose|glucose
C0804101|T201|LN|21307-4|LNC|glucose|glucose
C0804101|T201|MTH_LN|21307-4|LNC|glucose|glucose
C0804101|T201|OSN|21307-4|LNC|glucose|glucose
C0804101|T201|LC|21307-4|LNC|glucose|glucose
C0804102|T201|LN|21308-2|LNC|glucose|glucose
C0804102|T201|MTH_LN|21308-2|LNC|glucose|glucose
C0804102|T201|OSN|21308-2|LNC|glucose|glucose
C0804102|T201|LC|21308-2|LNC|glucose|glucose
C0804103|T201|LN|21309-0|LNC|glucose|glucose
C0804103|T201|MTH_LN|21309-0|LNC|glucose|glucose
C0804103|T201|OSN|21309-0|LNC|glucose|glucose
C0804103|T201|LC|21309-0|LNC|glucose|glucose
C0804104|T201|LN|21310-8|LNC|glucose|glucose
C0804104|T201|MTH_LN|21310-8|LNC|glucose|glucose
C0804104|T201|OSN|21310-8|LNC|glucose|glucose
C0804104|T201|LC|21310-8|LNC|glucose|glucose
C0804319|T201|LN|21525-1|LNC|sodium|sodium
C0804319|T201|MTH_LN|21525-1|LNC|sodium|sodium
C0804319|T201|OSN|21525-1|LNC|sodium|sodium
C0804319|T201|LC|21525-1|LNC|sodium|sodium
C0804376|T201|LN|21582-2|LNC|mast cell beta-tryptase|mast cell beta-tryptase
C0804376|T201|MTH_LN|21582-2|LNC|mast cell beta-tryptase|mast cell beta-tryptase
C0804376|T201|OSN|21582-2|LNC|mast cell beta-tryptase|mast cell beta-tryptase
C0804376|T201|LC|21582-2|LNC|mast cell beta-tryptase|mast cell beta-tryptase
C0804381|T201|LC|21587-1|LNC|urate|urate
C0804381|T201|MTH_LN|21587-1|LNC|urate|urate
C0804381|T201|OSN|21587-1|LNC|urate|urate
C0804381|T201|LN|21587-1|LNC|urate|urate
C0804381|T201|LC|21587-1|LNC|uric acid|uric acid
C0804381|T201|MTH_LN|21587-1|LNC|uric acid|uric acid
C0804381|T201|OSN|21587-1|LNC|uric acid|uric acid
C0804381|T201|LN|21587-1|LNC|uric acid|uric acid
C0812462|T201|LN|19072-8|LNC|calcium|calcium
C0812462|T201|MTH_LN|19072-8|LNC|calcium|calcium
C0812462|T201|OSN|19072-8|LNC|calcium|calcium
C0812462|T201|LC|19072-8|LNC|calcium|calcium
C0812462|T201|LN|19072-8|LNC|calcium homeostasis|calcium homeostasis
C0812462|T201|MTH_LN|19072-8|LNC|calcium homeostasis|calcium homeostasis
C0812462|T201|OSN|19072-8|LNC|calcium homeostasis|calcium homeostasis
C0812462|T201|LC|19072-8|LNC|calcium homeostasis|calcium homeostasis
C0880188|T201|LN|22670-4|LNC|isoleucine|isoleucine
C0880188|T201|MTH_LN|22670-4|LNC|isoleucine|isoleucine
C0880188|T201|OSN|22670-4|LNC|isoleucine|isoleucine
C0880188|T201|LC|22670-4|LNC|isoleucine|isoleucine
C0880188|T201|LN|22670-4|LNC|isoleucine metabolism|isoleucine metabolism
C0880188|T201|MTH_LN|22670-4|LNC|isoleucine metabolism|isoleucine metabolism
C0880188|T201|OSN|22670-4|LNC|isoleucine metabolism|isoleucine metabolism
C0880188|T201|LC|22670-4|LNC|isoleucine metabolism|isoleucine metabolism
C0880189|T201|LN|22671-2|LNC|phytanic acid|phytanic acid
C0880189|T201|MTH_LN|22671-2|LNC|phytanic acid|phytanic acid
C0880189|T201|OSN|22671-2|LNC|phytanic acid|phytanic acid
C0880189|T201|LC|22671-2|LNC|phytanic acid|phytanic acid
C0880190|T201|LN|22672-0|LNC|cysteine metabolism|cysteine metabolism
C0880190|T201|MTH_LN|22672-0|LNC|cysteine metabolism|cysteine metabolism
C0880190|T201|OSN|22672-0|LNC|cysteine metabolism|cysteine metabolism
C0880190|T201|LC|22672-0|LNC|cysteine metabolism|cysteine metabolism
C0880191|T201|MTH_LN|20646-6|LNC|homocystine|homocystine
C0880191|T201|OSN|20646-6|LNC|homocystine|homocystine
C0880191|T201|LN|20646-6|LNC|homocystine|homocystine
C0880191|T201|LC|20646-6|LNC|homocystine|homocystine
C0880191|T201|MTH_LN|20646-6|LNC|homocysteine metabolism|homocysteine metabolism
C0880191|T201|OSN|20646-6|LNC|homocysteine metabolism|homocysteine metabolism
C0880191|T201|LN|20646-6|LNC|homocysteine metabolism|homocysteine metabolism
C0880191|T201|LC|20646-6|LNC|homocysteine metabolism|homocysteine metabolism
C0880214|T201|LN|22705-8|LNC|glucose|glucose
C0880214|T201|MTH_LN|22705-8|LNC|glucose|glucose
C0880214|T201|OSN|22705-8|LNC|glucose|glucose
C0880214|T201|LC|22705-8|LNC|glucose|glucose
C0880253|T201|LN|22748-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0880253|T201|MTH_LN|22748-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0880253|T201|OSN|22748-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0880253|T201|LC|22748-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C0880253|T201|LN|22748-8|LNC|LDL|LDL
C0880253|T201|MTH_LN|22748-8|LNC|LDL|LDL
C0880253|T201|OSN|22748-8|LNC|LDL|LDL
C0880253|T201|LC|22748-8|LNC|LDL|LDL
C0880253|T201|LN|22748-8|LNC|LDL cholesterol|LDL cholesterol
C0880253|T201|MTH_LN|22748-8|LNC|LDL cholesterol|LDL cholesterol
C0880253|T201|OSN|22748-8|LNC|LDL cholesterol|LDL cholesterol
C0880253|T201|LC|22748-8|LNC|LDL cholesterol|LDL cholesterol
C0880253|T201|LN|22748-8|LNC|low-density lipoprotein|low-density lipoprotein
C0880253|T201|MTH_LN|22748-8|LNC|low-density lipoprotein|low-density lipoprotein
C0880253|T201|OSN|22748-8|LNC|low-density lipoprotein|low-density lipoprotein
C0880253|T201|LC|22748-8|LNC|low-density lipoprotein|low-density lipoprotein
C0880253|T201|LN|22748-8|LNC|beta-lipoproteins|beta-lipoproteins
C0880253|T201|MTH_LN|22748-8|LNC|beta-lipoproteins|beta-lipoproteins
C0880253|T201|OSN|22748-8|LNC|beta-lipoproteins|beta-lipoproteins
C0880253|T201|LC|22748-8|LNC|beta-lipoproteins|beta-lipoproteins
C0880253|T201|LN|22748-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0880253|T201|MTH_LN|22748-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0880253|T201|OSN|22748-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0880253|T201|LC|22748-8|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C0880253|T201|LN|22748-8|LNC|LDL-C|LDL-C
C0880253|T201|MTH_LN|22748-8|LNC|LDL-C|LDL-C
C0880253|T201|OSN|22748-8|LNC|LDL-C|LDL-C
C0880253|T201|LC|22748-8|LNC|LDL-C|LDL-C
C0880263|T201|LN|22763-7|LNC|ammonia|ammonia
C0880263|T201|MTH_LN|22763-7|LNC|ammonia|ammonia
C0880263|T201|OSN|22763-7|LNC|ammonia|ammonia
C0880263|T201|LC|22763-7|LNC|ammonia|ammonia
C0880263|T201|MTH_LN|35254-2|LNC|ammonia|ammonia
C0880263|T201|OSN|35254-2|LNC|ammonia|ammonia
C0880263|T201|LN|35254-2|LNC|ammonia|ammonia
C0880263|T201|LC|35254-2|LNC|ammonia|ammonia
C0881213|T201|LN|23860-0|LNC|erythrocyte volume|erythrocyte volume
C0881213|T201|OSN|23860-0|LNC|erythrocyte volume|erythrocyte volume
C0881213|T201|MTH_LN|23860-0|LNC|erythrocyte volume|erythrocyte volume
C0881213|T201|LC|23860-0|LNC|erythrocyte volume|erythrocyte volume
C0881213|T201|LN|23860-0|LNC|mean corpuscular volume|mean corpuscular volume
C0881213|T201|OSN|23860-0|LNC|mean corpuscular volume|mean corpuscular volume
C0881213|T201|MTH_LN|23860-0|LNC|mean corpuscular volume|mean corpuscular volume
C0881213|T201|LC|23860-0|LNC|mean corpuscular volume|mean corpuscular volume
C0881630|T201|LN|24360-0|LNC|hematocrit|hematocrit
C0881630|T201|MTH_LN|24360-0|LNC|hematocrit|hematocrit
C0881630|T201|OSN|24360-0|LNC|hematocrit|hematocrit
C0881630|T201|LC|24360-0|LNC|hematocrit|hematocrit
C0881654|T201|LN|24389-9|LNC|cortisol|cortisol
C0881654|T201|MTH_LN|24389-9|LNC|cortisol|cortisol
C0881654|T201|OSN|24389-9|LNC|cortisol|cortisol
C0881654|T201|LC|24389-9|LNC|cortisol|cortisol
C0881654|T201|LN|24389-9|LNC|cortisol low|cortisol low
C0881654|T201|MTH_LN|24389-9|LNC|cortisol low|cortisol low
C0881654|T201|OSN|24389-9|LNC|cortisol low|cortisol low
C0881654|T201|LC|24389-9|LNC|cortisol low|cortisol low
C0881654|T201|LN|24389-9|LNC|to undetectable cortisol|to undetectable cortisol
C0881654|T201|MTH_LN|24389-9|LNC|to undetectable cortisol|to undetectable cortisol
C0881654|T201|OSN|24389-9|LNC|to undetectable cortisol|to undetectable cortisol
C0881654|T201|LC|24389-9|LNC|to undetectable cortisol|to undetectable cortisol
C0881655|T201|LN|24390-7|LNC|cortisol|cortisol
C0881655|T201|MTH_LN|24390-7|LNC|cortisol|cortisol
C0881655|T201|OSN|24390-7|LNC|cortisol|cortisol
C0881655|T201|LC|24390-7|LNC|cortisol|cortisol
C0881655|T201|LN|24390-7|LNC|cortisol low|cortisol low
C0881655|T201|MTH_LN|24390-7|LNC|cortisol low|cortisol low
C0881655|T201|OSN|24390-7|LNC|cortisol low|cortisol low
C0881655|T201|LC|24390-7|LNC|cortisol low|cortisol low
C0881655|T201|LN|24390-7|LNC|to undetectable cortisol|to undetectable cortisol
C0881655|T201|MTH_LN|24390-7|LNC|to undetectable cortisol|to undetectable cortisol
C0881655|T201|OSN|24390-7|LNC|to undetectable cortisol|to undetectable cortisol
C0881655|T201|LC|24390-7|LNC|to undetectable cortisol|to undetectable cortisol
C0881656|T201|LN|24391-5|LNC|cortisol|cortisol
C0881656|T201|MTH_LN|24391-5|LNC|cortisol|cortisol
C0881656|T201|OSN|24391-5|LNC|cortisol|cortisol
C0881656|T201|LC|24391-5|LNC|cortisol|cortisol
C0881656|T201|LN|24391-5|LNC|cortisol low|cortisol low
C0881656|T201|MTH_LN|24391-5|LNC|cortisol low|cortisol low
C0881656|T201|OSN|24391-5|LNC|cortisol low|cortisol low
C0881656|T201|LC|24391-5|LNC|cortisol low|cortisol low
C0881656|T201|LN|24391-5|LNC|to undetectable cortisol|to undetectable cortisol
C0881656|T201|MTH_LN|24391-5|LNC|to undetectable cortisol|to undetectable cortisol
C0881656|T201|OSN|24391-5|LNC|to undetectable cortisol|to undetectable cortisol
C0881656|T201|LC|24391-5|LNC|to undetectable cortisol|to undetectable cortisol
C0881709|T201|MTH_LN|20659-9|LNC|tryptophan metabolism|tryptophan metabolism
C0881709|T201|LN|20659-9|LNC|tryptophan metabolism|tryptophan metabolism
C0881709|T201|OSN|20659-9|LNC|tryptophan metabolism|tryptophan metabolism
C0881709|T201|LC|20659-9|LNC|tryptophan metabolism|tryptophan metabolism
C0881712|T201|LN|24461-6|LNC|free fatty acid|free fatty acid
C0881712|T201|MTH_LN|24461-6|LNC|free fatty acid|free fatty acid
C0881712|T201|OSN|24461-6|LNC|free fatty acid|free fatty acid
C0881712|T201|LC|24461-6|LNC|free fatty acid|free fatty acid
C0881712|T201|LN|24461-6|LNC|fatty acids|fatty acids
C0881712|T201|MTH_LN|24461-6|LNC|fatty acids|fatty acids
C0881712|T201|OSN|24461-6|LNC|fatty acids|fatty acids
C0881712|T201|LC|24461-6|LNC|fatty acids|fatty acids
C0881717|T201|MTH_LN|24467-3|LNC|CD4-positive T|CD4-positive T
C0881717|T201|LC|24467-3|LNC|CD4-positive T|CD4-positive T
C0881717|T201|LN|24467-3|LNC|CD4-positive T|CD4-positive T
C0881717|T201|OSN|24467-3|LNC|CD4-positive T|CD4-positive T
C0881717|T201|MTH_LN|24467-3|LNC|CD4+ T|CD4+ T
C0881717|T201|LC|24467-3|LNC|CD4+ T|CD4+ T
C0881717|T201|LN|24467-3|LNC|CD4+ T|CD4+ T
C0881717|T201|OSN|24467-3|LNC|CD4+ T|CD4+ T
C0881717|T201|MTH_LN|24467-3|LNC|CD4 T|CD4 T
C0881717|T201|LC|24467-3|LNC|CD4 T|CD4 T
C0881717|T201|LN|24467-3|LNC|CD4 T|CD4 T
C0881717|T201|OSN|24467-3|LNC|CD4 T|CD4 T
C0882311|T201|LN|22697-7|LNC|arginine|arginine
C0882311|T201|OSN|22697-7|LNC|arginine|arginine
C0882311|T201|LC|22697-7|LNC|arginine|arginine
C0882311|T201|MTH_LN|22697-7|LNC|arginine|arginine
C0941310|T201|LN|25102-5|LNC|galactose|galactose
C0941310|T201|OSN|25102-5|LNC|galactose|galactose
C0941310|T201|LC|25102-5|LNC|galactose|galactose
C0941310|T201|MTH_LN|25102-5|LNC|galactose|galactose
C0941338|T201|LN|25138-9|LNC|taurine|taurine
C0941338|T201|OSN|25138-9|LNC|taurine|taurine
C0941338|T201|LC|25138-9|LNC|taurine|taurine
C0941338|T201|MTH_LN|25138-9|LNC|taurine|taurine
C0941344|T201|LN|25145-4|LNC|bacteria|bacteria
C0941344|T201|MTH_LN|25145-4|LNC|bacteria|bacteria
C0941344|T201|OSN|25145-4|LNC|bacteria|bacteria
C0941344|T201|LC|25145-4|LNC|bacteria|bacteria
C0941475|T201|LN|25303-9|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0941475|T201|MTH_LN|25303-9|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0941475|T201|OSN|25303-9|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0941475|T201|LC|25303-9|LNC|stool alpha1-antitrypsin|stool alpha1-antitrypsin
C0941489|T201|LN|25322-9|LNC|arginine|arginine
C0941489|T201|MTH_LN|25322-9|LNC|arginine|arginine
C0941489|T201|OSN|25322-9|LNC|arginine|arginine
C0941489|T201|LC|25322-9|LNC|arginine|arginine
C0941525|T201|LN|25371-6|LNC|VLDL cholesterol|VLDL cholesterol
C0941525|T201|MTH_LN|25371-6|LNC|VLDL cholesterol|VLDL cholesterol
C0941525|T201|OSN|25371-6|LNC|VLDL cholesterol|VLDL cholesterol
C0941525|T201|LC|25371-6|LNC|VLDL cholesterol|VLDL cholesterol
C0941525|T201|LN|25371-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0941525|T201|MTH_LN|25371-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0941525|T201|OSN|25371-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0941525|T201|LC|25371-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C0941525|T201|LN|25371-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0941525|T201|MTH_LN|25371-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0941525|T201|OSN|25371-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0941525|T201|LC|25371-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C0941525|T201|LN|25371-6|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0941525|T201|MTH_LN|25371-6|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0941525|T201|OSN|25371-6|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0941525|T201|LC|25371-6|LNC|lipoprotein cholesterol|lipoprotein cholesterol
C0941562|T201|LN|25415-1|LNC|folate metabolism|folate metabolism
C0941562|T201|MTH_LN|25415-1|LNC|folate metabolism|folate metabolism
C0941562|T201|OSN|25415-1|LNC|folate metabolism|folate metabolism
C0941562|T201|LC|25415-1|LNC|folate metabolism|folate metabolism
C0941601|T201|LN|25464-9|LNC|lysine|lysine
C0941601|T201|MTH_LN|25464-9|LNC|lysine|lysine
C0941601|T201|OSN|25464-9|LNC|lysine|lysine
C0941601|T201|LC|25464-9|LNC|lysine|lysine
C0941652|T201|LN|25533-1|LNC|taurine|taurine
C0941652|T201|MTH_LN|25533-1|LNC|taurine|taurine
C0941652|T201|OSN|25533-1|LNC|taurine|taurine
C0941652|T201|LC|25533-1|LNC|taurine|taurine
C0941683|T201|LN|25568-7|LNC|C-peptide|C-peptide
C0941683|T201|MTH_LN|25568-7|LNC|C-peptide|C-peptide
C0941683|T201|OSN|25568-7|LNC|C-peptide|C-peptide
C0941683|T201|LC|25568-7|LNC|C-peptide|C-peptide
C0941683|T201|LN|25568-7|LNC|C peptide|C peptide
C0941683|T201|MTH_LN|25568-7|LNC|C peptide|C peptide
C0941683|T201|OSN|25568-7|LNC|C peptide|C peptide
C0941683|T201|LC|25568-7|LNC|C peptide|C peptide
C0941684|T201|LN|25569-5|LNC|C-peptide|C-peptide
C0941684|T201|MTH_LN|25569-5|LNC|C-peptide|C-peptide
C0941684|T201|OSN|25569-5|LNC|C-peptide|C-peptide
C0941684|T201|LC|25569-5|LNC|C-peptide|C-peptide
C0941684|T201|LN|25569-5|LNC|C peptide|C peptide
C0941684|T201|MTH_LN|25569-5|LNC|C peptide|C peptide
C0941684|T201|OSN|25569-5|LNC|C peptide|C peptide
C0941684|T201|LC|25569-5|LNC|C peptide|C peptide
C0941685|T201|LN|25570-3|LNC|C-peptide|C-peptide
C0941685|T201|MTH_LN|25570-3|LNC|C-peptide|C-peptide
C0941685|T201|OSN|25570-3|LNC|C-peptide|C-peptide
C0941685|T201|LC|25570-3|LNC|C-peptide|C-peptide
C0941685|T201|LN|25570-3|LNC|C peptide|C peptide
C0941685|T201|MTH_LN|25570-3|LNC|C peptide|C peptide
C0941685|T201|OSN|25570-3|LNC|C peptide|C peptide
C0941685|T201|LC|25570-3|LNC|C peptide|C peptide
C0941686|T201|LN|25571-1|LNC|C-peptide|C-peptide
C0941686|T201|MTH_LN|25571-1|LNC|C-peptide|C-peptide
C0941686|T201|OSN|25571-1|LNC|C-peptide|C-peptide
C0941686|T201|LC|25571-1|LNC|C-peptide|C-peptide
C0941686|T201|LN|25571-1|LNC|C peptide|C peptide
C0941686|T201|MTH_LN|25571-1|LNC|C peptide|C peptide
C0941686|T201|OSN|25571-1|LNC|C peptide|C peptide
C0941686|T201|LC|25571-1|LNC|C peptide|C peptide
C0941687|T201|LN|25572-9|LNC|C-peptide|C-peptide
C0941687|T201|MTH_LN|25572-9|LNC|C-peptide|C-peptide
C0941687|T201|OSN|25572-9|LNC|C-peptide|C-peptide
C0941687|T201|LC|25572-9|LNC|C-peptide|C-peptide
C0941687|T201|LN|25572-9|LNC|C peptide|C peptide
C0941687|T201|MTH_LN|25572-9|LNC|C peptide|C peptide
C0941687|T201|OSN|25572-9|LNC|C peptide|C peptide
C0941687|T201|LC|25572-9|LNC|C peptide|C peptide
C0941688|T201|LN|25575-2|LNC|C-peptide|C-peptide
C0941688|T201|MTH_LN|25575-2|LNC|C-peptide|C-peptide
C0941688|T201|OSN|25575-2|LNC|C-peptide|C-peptide
C0941688|T201|LC|25575-2|LNC|C-peptide|C-peptide
C0941688|T201|LN|25575-2|LNC|C peptide|C peptide
C0941688|T201|MTH_LN|25575-2|LNC|C peptide|C peptide
C0941688|T201|OSN|25575-2|LNC|C peptide|C peptide
C0941688|T201|LC|25575-2|LNC|C peptide|C peptide
C0941689|T201|LN|25576-0|LNC|C-peptide|C-peptide
C0941689|T201|MTH_LN|25576-0|LNC|C-peptide|C-peptide
C0941689|T201|OSN|25576-0|LNC|C-peptide|C-peptide
C0941689|T201|LC|25576-0|LNC|C-peptide|C-peptide
C0941689|T201|LN|25576-0|LNC|C peptide|C peptide
C0941689|T201|MTH_LN|25576-0|LNC|C peptide|C peptide
C0941689|T201|OSN|25576-0|LNC|C peptide|C peptide
C0941689|T201|LC|25576-0|LNC|C peptide|C peptide
C0941690|T201|LN|25577-8|LNC|C-peptide|C-peptide
C0941690|T201|MTH_LN|25577-8|LNC|C-peptide|C-peptide
C0941690|T201|OSN|25577-8|LNC|C-peptide|C-peptide
C0941690|T201|LC|25577-8|LNC|C-peptide|C-peptide
C0941690|T201|LN|25577-8|LNC|C peptide|C peptide
C0941690|T201|MTH_LN|25577-8|LNC|C peptide|C peptide
C0941690|T201|OSN|25577-8|LNC|C peptide|C peptide
C0941690|T201|LC|25577-8|LNC|C peptide|C peptide
C0941691|T201|LN|25578-6|LNC|C-peptide|C-peptide
C0941691|T201|MTH_LN|25578-6|LNC|C-peptide|C-peptide
C0941691|T201|OSN|25578-6|LNC|C-peptide|C-peptide
C0941691|T201|LC|25578-6|LNC|C-peptide|C-peptide
C0941691|T201|LN|25578-6|LNC|C peptide|C peptide
C0941691|T201|MTH_LN|25578-6|LNC|C peptide|C peptide
C0941691|T201|OSN|25578-6|LNC|C peptide|C peptide
C0941691|T201|LC|25578-6|LNC|C peptide|C peptide
C0941692|T201|LN|25579-4|LNC|C-peptide|C-peptide
C0941692|T201|MTH_LN|25579-4|LNC|C-peptide|C-peptide
C0941692|T201|OSN|25579-4|LNC|C-peptide|C-peptide
C0941692|T201|LC|25579-4|LNC|C-peptide|C-peptide
C0941692|T201|LN|25579-4|LNC|C peptide|C peptide
C0941692|T201|MTH_LN|25579-4|LNC|C peptide|C peptide
C0941692|T201|OSN|25579-4|LNC|C peptide|C peptide
C0941692|T201|LC|25579-4|LNC|C peptide|C peptide
C0941693|T201|LN|25580-2|LNC|C-peptide|C-peptide
C0941693|T201|MTH_LN|25580-2|LNC|C-peptide|C-peptide
C0941693|T201|OSN|25580-2|LNC|C-peptide|C-peptide
C0941693|T201|LC|25580-2|LNC|C-peptide|C-peptide
C0941693|T201|LN|25580-2|LNC|C peptide|C peptide
C0941693|T201|MTH_LN|25580-2|LNC|C peptide|C peptide
C0941693|T201|OSN|25580-2|LNC|C peptide|C peptide
C0941693|T201|LC|25580-2|LNC|C peptide|C peptide
C0941694|T201|LN|25581-0|LNC|C-peptide|C-peptide
C0941694|T201|MTH_LN|25581-0|LNC|C-peptide|C-peptide
C0941694|T201|OSN|25581-0|LNC|C-peptide|C-peptide
C0941694|T201|LC|25581-0|LNC|C-peptide|C-peptide
C0941694|T201|LN|25581-0|LNC|C peptide|C peptide
C0941694|T201|MTH_LN|25581-0|LNC|C peptide|C peptide
C0941694|T201|OSN|25581-0|LNC|C peptide|C peptide
C0941694|T201|LC|25581-0|LNC|C peptide|C peptide
C0941695|T201|LN|25582-8|LNC|C-peptide|C-peptide
C0941695|T201|MTH_LN|25582-8|LNC|C-peptide|C-peptide
C0941695|T201|OSN|25582-8|LNC|C-peptide|C-peptide
C0941695|T201|LC|25582-8|LNC|C-peptide|C-peptide
C0941695|T201|LN|25582-8|LNC|C peptide|C peptide
C0941695|T201|MTH_LN|25582-8|LNC|C peptide|C peptide
C0941695|T201|OSN|25582-8|LNC|C peptide|C peptide
C0941695|T201|LC|25582-8|LNC|C peptide|C peptide
C0941756|T201|LN|25663-6|LNC|glucose|glucose
C0941756|T201|MTH_LN|25663-6|LNC|glucose|glucose
C0941756|T201|OSN|25663-6|LNC|glucose|glucose
C0941756|T201|LC|25663-6|LNC|glucose|glucose
C0941758|T201|LN|25665-1|LNC|glucose|glucose
C0941758|T201|MTH_LN|25665-1|LNC|glucose|glucose
C0941758|T201|OSN|25665-1|LNC|glucose|glucose
C0941758|T201|LC|25665-1|LNC|glucose|glucose
C0941760|T201|LN|25668-5|LNC|glucose|glucose
C0941760|T201|MTH_LN|25668-5|LNC|glucose|glucose
C0941760|T201|OSN|25668-5|LNC|glucose|glucose
C0941760|T201|LC|25668-5|LNC|glucose|glucose
C0941761|T201|LN|25669-3|LNC|glucose|glucose
C0941761|T201|MTH_LN|25669-3|LNC|glucose|glucose
C0941761|T201|OSN|25669-3|LNC|glucose|glucose
C0941761|T201|LC|25669-3|LNC|glucose|glucose
C0941763|T201|LN|25671-9|LNC|glucose|glucose
C0941763|T201|MTH_LN|25671-9|LNC|glucose|glucose
C0941763|T201|OSN|25671-9|LNC|glucose|glucose
C0941763|T201|LC|25671-9|LNC|glucose|glucose
C0941764|T201|LN|25672-7|LNC|glucose|glucose
C0941764|T201|MTH_LN|25672-7|LNC|glucose|glucose
C0941764|T201|OSN|25672-7|LNC|glucose|glucose
C0941764|T201|LC|25672-7|LNC|glucose|glucose
C0941765|T201|LN|25673-5|LNC|glucose|glucose
C0941765|T201|MTH_LN|25673-5|LNC|glucose|glucose
C0941765|T201|OSN|25673-5|LNC|glucose|glucose
C0941765|T201|LC|25673-5|LNC|glucose|glucose
C0941766|T201|LN|25674-3|LNC|glucose|glucose
C0941766|T201|MTH_LN|25674-3|LNC|glucose|glucose
C0941766|T201|OSN|25674-3|LNC|glucose|glucose
C0941766|T201|LC|25674-3|LNC|glucose|glucose
C0941768|T201|LN|25676-8|LNC|glucose|glucose
C0941768|T201|MTH_LN|25676-8|LNC|glucose|glucose
C0941768|T201|OSN|25676-8|LNC|glucose|glucose
C0941768|T201|LC|25676-8|LNC|glucose|glucose
C0941769|T201|LN|25677-6|LNC|glucose|glucose
C0941769|T201|MTH_LN|25677-6|LNC|glucose|glucose
C0941769|T201|OSN|25677-6|LNC|glucose|glucose
C0941769|T201|LC|25677-6|LNC|glucose|glucose
C0941770|T201|LN|25679-2|LNC|glucose|glucose
C0941770|T201|OSN|25679-2|LNC|glucose|glucose
C0941770|T201|MTH_LN|25679-2|LNC|glucose|glucose
C0941770|T201|LC|25679-2|LNC|glucose|glucose
C0941771|T201|LN|25680-0|LNC|glucose|glucose
C0941771|T201|MTH_LN|25680-0|LNC|glucose|glucose
C0941771|T201|OSN|25680-0|LNC|glucose|glucose
C0941771|T201|LC|25680-0|LNC|glucose|glucose
C0941802|T201|LN|25717-0|LNC|luteinizing|luteinizing
C0941802|T201|OSN|25717-0|LNC|luteinizing|luteinizing
C0941802|T201|MTH_LN|25717-0|LNC|luteinizing|luteinizing
C0941802|T201|LC|25717-0|LNC|luteinizing|luteinizing
C0941802|T201|LN|25717-0|LNC|LH|LH
C0941802|T201|OSN|25717-0|LNC|LH|LH
C0941802|T201|MTH_LN|25717-0|LNC|LH|LH
C0941802|T201|LC|25717-0|LNC|LH|LH
C0941802|T201|LN|25717-0|LNC|luteinising|luteinising
C0941802|T201|OSN|25717-0|LNC|luteinising|luteinising
C0941802|T201|MTH_LN|25717-0|LNC|luteinising|luteinising
C0941802|T201|LC|25717-0|LNC|luteinising|luteinising
C0941803|T201|LN|25718-8|LNC|luteinizing|luteinizing
C0941803|T201|MTH_LN|25718-8|LNC|luteinizing|luteinizing
C0941803|T201|OSN|25718-8|LNC|luteinizing|luteinizing
C0941803|T201|LC|25718-8|LNC|luteinizing|luteinizing
C0941803|T201|LN|25718-8|LNC|LH|LH
C0941803|T201|MTH_LN|25718-8|LNC|LH|LH
C0941803|T201|OSN|25718-8|LNC|LH|LH
C0941803|T201|LC|25718-8|LNC|LH|LH
C0941803|T201|LN|25718-8|LNC|luteinising|luteinising
C0941803|T201|MTH_LN|25718-8|LNC|luteinising|luteinising
C0941803|T201|OSN|25718-8|LNC|luteinising|luteinising
C0941803|T201|LC|25718-8|LNC|luteinising|luteinising
C0941804|T201|LN|25719-6|LNC|luteinizing|luteinizing
C0941804|T201|MTH_LN|25719-6|LNC|luteinizing|luteinizing
C0941804|T201|OSN|25719-6|LNC|luteinizing|luteinizing
C0941804|T201|LC|25719-6|LNC|luteinizing|luteinizing
C0941804|T201|LN|25719-6|LNC|LH|LH
C0941804|T201|MTH_LN|25719-6|LNC|LH|LH
C0941804|T201|OSN|25719-6|LNC|LH|LH
C0941804|T201|LC|25719-6|LNC|LH|LH
C0941804|T201|LN|25719-6|LNC|luteinising|luteinising
C0941804|T201|MTH_LN|25719-6|LNC|luteinising|luteinising
C0941804|T201|OSN|25719-6|LNC|luteinising|luteinising
C0941804|T201|LC|25719-6|LNC|luteinising|luteinising
C0941805|T201|LN|25720-4|LNC|luteinizing|luteinizing
C0941805|T201|MTH_LN|25720-4|LNC|luteinizing|luteinizing
C0941805|T201|OSN|25720-4|LNC|luteinizing|luteinizing
C0941805|T201|LC|25720-4|LNC|luteinizing|luteinizing
C0941805|T201|LN|25720-4|LNC|LH|LH
C0941805|T201|MTH_LN|25720-4|LNC|LH|LH
C0941805|T201|OSN|25720-4|LNC|LH|LH
C0941805|T201|LC|25720-4|LNC|LH|LH
C0941805|T201|LN|25720-4|LNC|luteinising|luteinising
C0941805|T201|MTH_LN|25720-4|LNC|luteinising|luteinising
C0941805|T201|OSN|25720-4|LNC|luteinising|luteinising
C0941805|T201|LC|25720-4|LNC|luteinising|luteinising
C0941920|T201|LN|25860-8|LNC|arginine|arginine
C0941920|T201|MTH_LN|25860-8|LNC|arginine|arginine
C0941920|T201|OSN|25860-8|LNC|arginine|arginine
C0941920|T201|LC|25860-8|LNC|arginine|arginine
C0941921|T201|LN|25861-6|LNC|arginine|arginine
C0941921|T201|OSN|25861-6|LNC|arginine|arginine
C0941921|T201|LC|25861-6|LNC|arginine|arginine
C0941921|T201|MTH_LN|25861-6|LNC|arginine|arginine
C0941950|T201|LN|25899-6|LNC|lactate|lactate
C0941950|T201|OSN|25899-6|LNC|lactate|lactate
C0941950|T201|MTH_LN|25899-6|LNC|lactate|lactate
C0941950|T201|LC|25899-6|LNC|lactate|lactate
C0941951|T201|LN|25901-0|LNC|lactate|lactate
C0941951|T201|OSN|25901-0|LNC|lactate|lactate
C0941951|T201|MTH_LN|25901-0|LNC|lactate|lactate
C0941951|T201|LC|25901-0|LNC|lactate|lactate
C0941952|T201|LN|25902-8|LNC|lactate|lactate
C0941952|T201|OSN|25902-8|LNC|lactate|lactate
C0941952|T201|MTH_LN|25902-8|LNC|lactate|lactate
C0941952|T201|LC|25902-8|LNC|lactate|lactate
C0941953|T201|LN|25904-4|LNC|lactate|lactate
C0941953|T201|OSN|25904-4|LNC|lactate|lactate
C0941953|T201|MTH_LN|25904-4|LNC|lactate|lactate
C0941953|T201|LC|25904-4|LNC|lactate|lactate
C0941954|T201|LN|25905-1|LNC|lactate|lactate
C0941954|T201|OSN|25905-1|LNC|lactate|lactate
C0941954|T201|MTH_LN|25905-1|LNC|lactate|lactate
C0941954|T201|LC|25905-1|LNC|lactate|lactate
C0941985|T201|LN|25943-2|LNC|luteinizing|luteinizing
C0941985|T201|MTH_LN|25943-2|LNC|luteinizing|luteinizing
C0941985|T201|OSN|25943-2|LNC|luteinizing|luteinizing
C0941985|T201|LC|25943-2|LNC|luteinizing|luteinizing
C0941985|T201|LN|25943-2|LNC|LH|LH
C0941985|T201|MTH_LN|25943-2|LNC|LH|LH
C0941985|T201|OSN|25943-2|LNC|LH|LH
C0941985|T201|LC|25943-2|LNC|LH|LH
C0941985|T201|LN|25943-2|LNC|luteinising|luteinising
C0941985|T201|MTH_LN|25943-2|LNC|luteinising|luteinising
C0941985|T201|OSN|25943-2|LNC|luteinising|luteinising
C0941985|T201|LC|25943-2|LNC|luteinising|luteinising
C0941986|T201|LN|25944-0|LNC|luteinizing|luteinizing
C0941986|T201|MTH_LN|25944-0|LNC|luteinizing|luteinizing
C0941986|T201|OSN|25944-0|LNC|luteinizing|luteinizing
C0941986|T201|LC|25944-0|LNC|luteinizing|luteinizing
C0941986|T201|LN|25944-0|LNC|LH|LH
C0941986|T201|MTH_LN|25944-0|LNC|LH|LH
C0941986|T201|OSN|25944-0|LNC|LH|LH
C0941986|T201|LC|25944-0|LNC|LH|LH
C0941986|T201|LN|25944-0|LNC|luteinising|luteinising
C0941986|T201|MTH_LN|25944-0|LNC|luteinising|luteinising
C0941986|T201|OSN|25944-0|LNC|luteinising|luteinising
C0941986|T201|LC|25944-0|LNC|luteinising|luteinising
C0941987|T201|LN|25945-7|LNC|luteinizing|luteinizing
C0941987|T201|MTH_LN|25945-7|LNC|luteinizing|luteinizing
C0941987|T201|OSN|25945-7|LNC|luteinizing|luteinizing
C0941987|T201|LC|25945-7|LNC|luteinizing|luteinizing
C0941987|T201|LN|25945-7|LNC|LH|LH
C0941987|T201|MTH_LN|25945-7|LNC|LH|LH
C0941987|T201|OSN|25945-7|LNC|LH|LH
C0941987|T201|LC|25945-7|LNC|LH|LH
C0941987|T201|LN|25945-7|LNC|luteinising|luteinising
C0941987|T201|MTH_LN|25945-7|LNC|luteinising|luteinising
C0941987|T201|OSN|25945-7|LNC|luteinising|luteinising
C0941987|T201|LC|25945-7|LNC|luteinising|luteinising
C0941988|T201|LN|25947-3|LNC|luteinizing|luteinizing
C0941988|T201|MTH_LN|25947-3|LNC|luteinizing|luteinizing
C0941988|T201|OSN|25947-3|LNC|luteinizing|luteinizing
C0941988|T201|LC|25947-3|LNC|luteinizing|luteinizing
C0941988|T201|LN|25947-3|LNC|LH|LH
C0941988|T201|MTH_LN|25947-3|LNC|LH|LH
C0941988|T201|OSN|25947-3|LNC|LH|LH
C0941988|T201|LC|25947-3|LNC|LH|LH
C0941988|T201|LN|25947-3|LNC|luteinising|luteinising
C0941988|T201|MTH_LN|25947-3|LNC|luteinising|luteinising
C0941988|T201|OSN|25947-3|LNC|luteinising|luteinising
C0941988|T201|LC|25947-3|LNC|luteinising|luteinising
C0941989|T201|LN|25948-1|LNC|luteinizing|luteinizing
C0941989|T201|MTH_LN|25948-1|LNC|luteinizing|luteinizing
C0941989|T201|OSN|25948-1|LNC|luteinizing|luteinizing
C0941989|T201|LC|25948-1|LNC|luteinizing|luteinizing
C0941989|T201|LN|25948-1|LNC|LH|LH
C0941989|T201|MTH_LN|25948-1|LNC|LH|LH
C0941989|T201|OSN|25948-1|LNC|LH|LH
C0941989|T201|LC|25948-1|LNC|LH|LH
C0941989|T201|LN|25948-1|LNC|luteinising|luteinising
C0941989|T201|MTH_LN|25948-1|LNC|luteinising|luteinising
C0941989|T201|OSN|25948-1|LNC|luteinising|luteinising
C0941989|T201|LC|25948-1|LNC|luteinising|luteinising
C0941990|T201|LN|25949-9|LNC|luteinizing|luteinizing
C0941990|T201|MTH_LN|25949-9|LNC|luteinizing|luteinizing
C0941990|T201|OSN|25949-9|LNC|luteinizing|luteinizing
C0941990|T201|LC|25949-9|LNC|luteinizing|luteinizing
C0941990|T201|LN|25949-9|LNC|LH|LH
C0941990|T201|MTH_LN|25949-9|LNC|LH|LH
C0941990|T201|OSN|25949-9|LNC|LH|LH
C0941990|T201|LC|25949-9|LNC|LH|LH
C0941990|T201|LN|25949-9|LNC|luteinising|luteinising
C0941990|T201|MTH_LN|25949-9|LNC|luteinising|luteinising
C0941990|T201|OSN|25949-9|LNC|luteinising|luteinising
C0941990|T201|LC|25949-9|LNC|luteinising|luteinising
C0941991|T201|LN|25950-7|LNC|luteinizing|luteinizing
C0941991|T201|MTH_LN|25950-7|LNC|luteinizing|luteinizing
C0941991|T201|OSN|25950-7|LNC|luteinizing|luteinizing
C0941991|T201|LC|25950-7|LNC|luteinizing|luteinizing
C0941991|T201|LN|25950-7|LNC|LH|LH
C0941991|T201|MTH_LN|25950-7|LNC|LH|LH
C0941991|T201|OSN|25950-7|LNC|LH|LH
C0941991|T201|LC|25950-7|LNC|LH|LH
C0941991|T201|LN|25950-7|LNC|luteinising|luteinising
C0941991|T201|MTH_LN|25950-7|LNC|luteinising|luteinising
C0941991|T201|OSN|25950-7|LNC|luteinising|luteinising
C0941991|T201|LC|25950-7|LNC|luteinising|luteinising
C0941992|T201|LN|25951-5|LNC|luteinizing|luteinizing
C0941992|T201|MTH_LN|25951-5|LNC|luteinizing|luteinizing
C0941992|T201|OSN|25951-5|LNC|luteinizing|luteinizing
C0941992|T201|LC|25951-5|LNC|luteinizing|luteinizing
C0941992|T201|LN|25951-5|LNC|LH|LH
C0941992|T201|MTH_LN|25951-5|LNC|LH|LH
C0941992|T201|OSN|25951-5|LNC|LH|LH
C0941992|T201|LC|25951-5|LNC|LH|LH
C0941992|T201|LN|25951-5|LNC|luteinising|luteinising
C0941992|T201|MTH_LN|25951-5|LNC|luteinising|luteinising
C0941992|T201|OSN|25951-5|LNC|luteinising|luteinising
C0941992|T201|LC|25951-5|LNC|luteinising|luteinising
C0942023|T201|LN|25985-3|LNC|taurine|taurine
C0942023|T201|OSN|25985-3|LNC|taurine|taurine
C0942023|T201|LC|25985-3|LNC|taurine|taurine
C0942023|T201|MTH_LN|25985-3|LNC|taurine|taurine
C0942032|T201|LN|25997-8|LNC|urate|urate
C0942032|T201|MTH_LN|25997-8|LNC|urate|urate
C0942032|T201|OSN|25997-8|LNC|urate|urate
C0942032|T201|LC|25997-8|LNC|urate|urate
C0942032|T201|LN|25997-8|LNC|uric acid|uric acid
C0942032|T201|MTH_LN|25997-8|LNC|uric acid|uric acid
C0942032|T201|OSN|25997-8|LNC|uric acid|uric acid
C0942032|T201|LC|25997-8|LNC|uric acid|uric acid
C0942080|T201|LN|26054-7|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C0942080|T201|MTH_LN|26054-7|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C0942080|T201|OSN|26054-7|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C0942080|T201|LC|26054-7|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C0942414|T201|LN|26444-0|LNC|basophil count|basophil count
C0942414|T201|OSN|26444-0|LNC|basophil count|basophil count
C0942414|T201|MTH_LN|26444-0|LNC|basophil count|basophil count
C0942414|T201|LC|26444-0|LNC|basophil count|basophil count
C0942419|T201|LN|26449-9|LNC|eosinophil count|eosinophil count
C0942419|T201|OSN|26449-9|LNC|eosinophil count|eosinophil count
C0942419|T201|MTH_LN|26449-9|LNC|eosinophil count|eosinophil count
C0942419|T201|LC|26449-9|LNC|eosinophil count|eosinophil count
C0942437|T201|LN|26474-7|LNC|lymphocyte count|lymphocyte count
C0942437|T201|OSN|26474-7|LNC|lymphocyte count|lymphocyte count
C0942437|T201|MTH_LN|26474-7|LNC|lymphocyte count|lymphocyte count
C0942437|T201|LC|26474-7|LNC|lymphocyte count|lymphocyte count
C0942437|T201|LN|26474-7|LNC|lymphocyte number|lymphocyte number
C0942437|T201|OSN|26474-7|LNC|lymphocyte number|lymphocyte number
C0942437|T201|MTH_LN|26474-7|LNC|lymphocyte number|lymphocyte number
C0942437|T201|LC|26474-7|LNC|lymphocyte number|lymphocyte number
C0942437|T201|LN|26474-7|LNC|lymphocyte counts|lymphocyte counts
C0942437|T201|OSN|26474-7|LNC|lymphocyte counts|lymphocyte counts
C0942437|T201|MTH_LN|26474-7|LNC|lymphocyte counts|lymphocyte counts
C0942437|T201|LC|26474-7|LNC|lymphocyte counts|lymphocyte counts
C0942437|T201|LN|26474-7|LNC|lymphocytes|lymphocytes
C0942437|T201|OSN|26474-7|LNC|lymphocytes|lymphocytes
C0942437|T201|MTH_LN|26474-7|LNC|lymphocytes|lymphocytes
C0942437|T201|LC|26474-7|LNC|lymphocytes|lymphocytes
C0942437|T201|LN|26474-7|LNC|numberslymphocytes|numberslymphocytes
C0942437|T201|OSN|26474-7|LNC|numberslymphocytes|numberslymphocytes
C0942437|T201|MTH_LN|26474-7|LNC|numberslymphocytes|numberslymphocytes
C0942437|T201|LC|26474-7|LNC|numberslymphocytes|numberslymphocytes
C0942440|T201|LN|26478-8|LNC|lymphocyte count|lymphocyte count
C0942440|T201|OSN|26478-8|LNC|lymphocyte count|lymphocyte count
C0942440|T201|MTH_LN|26478-8|LNC|lymphocyte count|lymphocyte count
C0942440|T201|LC|26478-8|LNC|lymphocyte count|lymphocyte count
C0942440|T201|LN|26478-8|LNC|lymphocyte number|lymphocyte number
C0942440|T201|OSN|26478-8|LNC|lymphocyte number|lymphocyte number
C0942440|T201|MTH_LN|26478-8|LNC|lymphocyte number|lymphocyte number
C0942440|T201|LC|26478-8|LNC|lymphocyte number|lymphocyte number
C0942440|T201|LN|26478-8|LNC|lymphocyte counts|lymphocyte counts
C0942440|T201|OSN|26478-8|LNC|lymphocyte counts|lymphocyte counts
C0942440|T201|MTH_LN|26478-8|LNC|lymphocyte counts|lymphocyte counts
C0942440|T201|LC|26478-8|LNC|lymphocyte counts|lymphocyte counts
C0942440|T201|LN|26478-8|LNC|lymphocytes|lymphocytes
C0942440|T201|OSN|26478-8|LNC|lymphocytes|lymphocytes
C0942440|T201|MTH_LN|26478-8|LNC|lymphocytes|lymphocytes
C0942440|T201|LC|26478-8|LNC|lymphocytes|lymphocytes
C0942440|T201|LN|26478-8|LNC|numberslymphocytes|numberslymphocytes
C0942440|T201|OSN|26478-8|LNC|numberslymphocytes|numberslymphocytes
C0942440|T201|MTH_LN|26478-8|LNC|numberslymphocytes|numberslymphocytes
C0942440|T201|LC|26478-8|LNC|numberslymphocytes|numberslymphocytes
C0942441|T201|LN|26479-6|LNC|cerebrospinal fluid|cerebrospinal fluid
C0942441|T201|OSN|26479-6|LNC|cerebrospinal fluid|cerebrospinal fluid
C0942441|T201|MTH_LN|26479-6|LNC|cerebrospinal fluid|cerebrospinal fluid
C0942441|T201|LC|26479-6|LNC|cerebrospinal fluid|cerebrospinal fluid
C0942441|T201|LN|26479-6|LNC|CSF findings|CSF findings
C0942441|T201|OSN|26479-6|LNC|CSF findings|CSF findings
C0942441|T201|MTH_LN|26479-6|LNC|CSF findings|CSF findings
C0942441|T201|LC|26479-6|LNC|CSF findings|CSF findings
C0942441|T201|LN|26479-6|LNC|CSF|CSF
C0942441|T201|OSN|26479-6|LNC|CSF|CSF
C0942441|T201|MTH_LN|26479-6|LNC|CSF|CSF
C0942441|T201|LC|26479-6|LNC|CSF|CSF
C0942446|T201|LN|26484-6|LNC|monocyte number|monocyte number
C0942446|T201|OSN|26484-6|LNC|monocyte number|monocyte number
C0942446|T201|MTH_LN|26484-6|LNC|monocyte number|monocyte number
C0942446|T201|LC|26484-6|LNC|monocyte number|monocyte number
C0942446|T201|LN|26484-6|LNC|monocyte count|monocyte count
C0942446|T201|OSN|26484-6|LNC|monocyte count|monocyte count
C0942446|T201|MTH_LN|26484-6|LNC|monocyte count|monocyte count
C0942446|T201|LC|26484-6|LNC|monocyte count|monocyte count
C0942447|T201|LN|26485-3|LNC|monocyte number|monocyte number
C0942447|T201|OSN|26485-3|LNC|monocyte number|monocyte number
C0942447|T201|MTH_LN|26485-3|LNC|monocyte number|monocyte number
C0942447|T201|LC|26485-3|LNC|monocyte number|monocyte number
C0942447|T201|LN|26485-3|LNC|monocyte count|monocyte count
C0942447|T201|OSN|26485-3|LNC|monocyte count|monocyte count
C0942447|T201|MTH_LN|26485-3|LNC|monocyte count|monocyte count
C0942447|T201|LC|26485-3|LNC|monocyte count|monocyte count
C0942449|T201|LN|26487-9|LNC|monocyte number|monocyte number
C0942449|T201|OSN|26487-9|LNC|monocyte number|monocyte number
C0942449|T201|MTH_LN|26487-9|LNC|monocyte number|monocyte number
C0942449|T201|LC|26487-9|LNC|monocyte number|monocyte number
C0942449|T201|LN|26487-9|LNC|monocyte count|monocyte count
C0942449|T201|OSN|26487-9|LNC|monocyte count|monocyte count
C0942449|T201|MTH_LN|26487-9|LNC|monocyte count|monocyte count
C0942449|T201|LC|26487-9|LNC|monocyte count|monocyte count
C0942460|T201|LN|26498-6|LNC|myeloid leukocytes|myeloid leukocytes
C0942460|T201|OSN|26498-6|LNC|myeloid leukocytes|myeloid leukocytes
C0942460|T201|MTH_LN|26498-6|LNC|myeloid leukocytes|myeloid leukocytes
C0942460|T201|LC|26498-6|LNC|myeloid leukocytes|myeloid leukocytes
C0942461|T201|LN|26499-4|LNC|neutrophil counts|neutrophil counts
C0942461|T201|OSN|26499-4|LNC|neutrophil counts|neutrophil counts
C0942461|T201|MTH_LN|26499-4|LNC|neutrophil counts|neutrophil counts
C0942461|T201|LC|26499-4|LNC|neutrophil counts|neutrophil counts
C0942461|T201|LN|26499-4|LNC|neutrophil count|neutrophil count
C0942461|T201|OSN|26499-4|LNC|neutrophil count|neutrophil count
C0942461|T201|MTH_LN|26499-4|LNC|neutrophil count|neutrophil count
C0942461|T201|LC|26499-4|LNC|neutrophil count|neutrophil count
C0942461|T201|LN|26499-4|LNC|neutrophil|neutrophil
C0942461|T201|OSN|26499-4|LNC|neutrophil|neutrophil
C0942461|T201|MTH_LN|26499-4|LNC|neutrophil|neutrophil
C0942461|T201|LC|26499-4|LNC|neutrophil|neutrophil
C0942465|T201|LN|26503-3|LNC|neutrophil counts|neutrophil counts
C0942465|T201|OSN|26503-3|LNC|neutrophil counts|neutrophil counts
C0942465|T201|MTH_LN|26503-3|LNC|neutrophil counts|neutrophil counts
C0942465|T201|LC|26503-3|LNC|neutrophil counts|neutrophil counts
C0942465|T201|LN|26503-3|LNC|neutrophil count|neutrophil count
C0942465|T201|OSN|26503-3|LNC|neutrophil count|neutrophil count
C0942465|T201|MTH_LN|26503-3|LNC|neutrophil count|neutrophil count
C0942465|T201|LC|26503-3|LNC|neutrophil count|neutrophil count
C0942465|T201|LN|26503-3|LNC|neutrophil|neutrophil
C0942465|T201|OSN|26503-3|LNC|neutrophil|neutrophil
C0942465|T201|MTH_LN|26503-3|LNC|neutrophil|neutrophil
C0942465|T201|LC|26503-3|LNC|neutrophil|neutrophil
C0942468|T201|LN|26508-2|LNC|granulocyte precursors|granulocyte precursors
C0942468|T201|OSN|26508-2|LNC|granulocyte precursors|granulocyte precursors
C0942468|T201|MTH_LN|26508-2|LNC|granulocyte precursors|granulocyte precursors
C0942468|T201|LC|26508-2|LNC|granulocyte precursors|granulocyte precursors
C0942471|T201|LN|26511-6|LNC|neutrophil counts|neutrophil counts
C0942471|T201|OSN|26511-6|LNC|neutrophil counts|neutrophil counts
C0942471|T201|MTH_LN|26511-6|LNC|neutrophil counts|neutrophil counts
C0942471|T201|LC|26511-6|LNC|neutrophil counts|neutrophil counts
C0942471|T201|LN|26511-6|LNC|neutrophil count|neutrophil count
C0942471|T201|OSN|26511-6|LNC|neutrophil count|neutrophil count
C0942471|T201|MTH_LN|26511-6|LNC|neutrophil count|neutrophil count
C0942471|T201|LC|26511-6|LNC|neutrophil count|neutrophil count
C0942471|T201|LN|26511-6|LNC|neutrophil|neutrophil
C0942471|T201|OSN|26511-6|LNC|neutrophil|neutrophil
C0942471|T201|MTH_LN|26511-6|LNC|neutrophil|neutrophil
C0942471|T201|LC|26511-6|LNC|neutrophil|neutrophil
C0942474|T201|LN|26515-7|LNC|platelet count|platelet count
C0942474|T201|OSN|26515-7|LNC|platelet count|platelet count
C0942474|T201|MTH_LN|26515-7|LNC|platelet count|platelet count
C0942474|T201|LC|26515-7|LNC|platelet count|platelet count
C0942484|T201|LN|26528-0|LNC|cortisol|cortisol
C0942484|T201|MTH_LN|26528-0|LNC|cortisol|cortisol
C0942484|T201|OSN|26528-0|LNC|cortisol|cortisol
C0942484|T201|LC|26528-0|LNC|cortisol|cortisol
C0942484|T201|LN|26528-0|LNC|cortisol low|cortisol low
C0942484|T201|MTH_LN|26528-0|LNC|cortisol low|cortisol low
C0942484|T201|OSN|26528-0|LNC|cortisol low|cortisol low
C0942484|T201|LC|26528-0|LNC|cortisol low|cortisol low
C0942484|T201|LN|26528-0|LNC|to undetectable cortisol|to undetectable cortisol
C0942484|T201|MTH_LN|26528-0|LNC|to undetectable cortisol|to undetectable cortisol
C0942484|T201|OSN|26528-0|LNC|to undetectable cortisol|to undetectable cortisol
C0942484|T201|LC|26528-0|LNC|to undetectable cortisol|to undetectable cortisol
C0942485|T201|LN|26529-8|LNC|cortisol|cortisol
C0942485|T201|MTH_LN|26529-8|LNC|cortisol|cortisol
C0942485|T201|OSN|26529-8|LNC|cortisol|cortisol
C0942485|T201|LC|26529-8|LNC|cortisol|cortisol
C0942485|T201|LN|26529-8|LNC|cortisol low|cortisol low
C0942485|T201|MTH_LN|26529-8|LNC|cortisol low|cortisol low
C0942485|T201|OSN|26529-8|LNC|cortisol low|cortisol low
C0942485|T201|LC|26529-8|LNC|cortisol low|cortisol low
C0942485|T201|LN|26529-8|LNC|to undetectable cortisol|to undetectable cortisol
C0942485|T201|MTH_LN|26529-8|LNC|to undetectable cortisol|to undetectable cortisol
C0942485|T201|OSN|26529-8|LNC|to undetectable cortisol|to undetectable cortisol
C0942485|T201|LC|26529-8|LNC|to undetectable cortisol|to undetectable cortisol
C0942486|T201|LN|26530-6|LNC|cortisol|cortisol
C0942486|T201|MTH_LN|26530-6|LNC|cortisol|cortisol
C0942486|T201|OSN|26530-6|LNC|cortisol|cortisol
C0942486|T201|LC|26530-6|LNC|cortisol|cortisol
C0942486|T201|LN|26530-6|LNC|cortisol low|cortisol low
C0942486|T201|MTH_LN|26530-6|LNC|cortisol low|cortisol low
C0942486|T201|OSN|26530-6|LNC|cortisol low|cortisol low
C0942486|T201|LC|26530-6|LNC|cortisol low|cortisol low
C0942486|T201|LN|26530-6|LNC|to undetectable cortisol|to undetectable cortisol
C0942486|T201|MTH_LN|26530-6|LNC|to undetectable cortisol|to undetectable cortisol
C0942486|T201|OSN|26530-6|LNC|to undetectable cortisol|to undetectable cortisol
C0942486|T201|LC|26530-6|LNC|to undetectable cortisol|to undetectable cortisol
C0942487|T201|LN|26531-4|LNC|cortisol|cortisol
C0942487|T201|MTH_LN|26531-4|LNC|cortisol|cortisol
C0942487|T201|OSN|26531-4|LNC|cortisol|cortisol
C0942487|T201|LC|26531-4|LNC|cortisol|cortisol
C0942487|T201|LN|26531-4|LNC|cortisol low|cortisol low
C0942487|T201|MTH_LN|26531-4|LNC|cortisol low|cortisol low
C0942487|T201|OSN|26531-4|LNC|cortisol low|cortisol low
C0942487|T201|LC|26531-4|LNC|cortisol low|cortisol low
C0942487|T201|LN|26531-4|LNC|to undetectable cortisol|to undetectable cortisol
C0942487|T201|MTH_LN|26531-4|LNC|to undetectable cortisol|to undetectable cortisol
C0942487|T201|OSN|26531-4|LNC|to undetectable cortisol|to undetectable cortisol
C0942487|T201|LC|26531-4|LNC|to undetectable cortisol|to undetectable cortisol
C0942488|T201|LN|26534-8|LNC|cortisol|cortisol
C0942488|T201|MTH_LN|26534-8|LNC|cortisol|cortisol
C0942488|T201|OSN|26534-8|LNC|cortisol|cortisol
C0942488|T201|LC|26534-8|LNC|cortisol|cortisol
C0942488|T201|LN|26534-8|LNC|cortisol low|cortisol low
C0942488|T201|MTH_LN|26534-8|LNC|cortisol low|cortisol low
C0942488|T201|OSN|26534-8|LNC|cortisol low|cortisol low
C0942488|T201|LC|26534-8|LNC|cortisol low|cortisol low
C0942488|T201|LN|26534-8|LNC|to undetectable cortisol|to undetectable cortisol
C0942488|T201|MTH_LN|26534-8|LNC|to undetectable cortisol|to undetectable cortisol
C0942488|T201|OSN|26534-8|LNC|to undetectable cortisol|to undetectable cortisol
C0942488|T201|LC|26534-8|LNC|to undetectable cortisol|to undetectable cortisol
C0942489|T201|LN|26535-5|LNC|cortisol|cortisol
C0942489|T201|MTH_LN|26535-5|LNC|cortisol|cortisol
C0942489|T201|OSN|26535-5|LNC|cortisol|cortisol
C0942489|T201|LC|26535-5|LNC|cortisol|cortisol
C0942489|T201|LN|26535-5|LNC|cortisol low|cortisol low
C0942489|T201|MTH_LN|26535-5|LNC|cortisol low|cortisol low
C0942489|T201|OSN|26535-5|LNC|cortisol low|cortisol low
C0942489|T201|LC|26535-5|LNC|cortisol low|cortisol low
C0942489|T201|LN|26535-5|LNC|to undetectable cortisol|to undetectable cortisol
C0942489|T201|MTH_LN|26535-5|LNC|to undetectable cortisol|to undetectable cortisol
C0942489|T201|OSN|26535-5|LNC|to undetectable cortisol|to undetectable cortisol
C0942489|T201|LC|26535-5|LNC|to undetectable cortisol|to undetectable cortisol
C0942490|T201|LN|26536-3|LNC|cortisol|cortisol
C0942490|T201|MTH_LN|26536-3|LNC|cortisol|cortisol
C0942490|T201|OSN|26536-3|LNC|cortisol|cortisol
C0942490|T201|LC|26536-3|LNC|cortisol|cortisol
C0942490|T201|LN|26536-3|LNC|cortisol low|cortisol low
C0942490|T201|MTH_LN|26536-3|LNC|cortisol low|cortisol low
C0942490|T201|OSN|26536-3|LNC|cortisol low|cortisol low
C0942490|T201|LC|26536-3|LNC|cortisol low|cortisol low
C0942490|T201|LN|26536-3|LNC|to undetectable cortisol|to undetectable cortisol
C0942490|T201|MTH_LN|26536-3|LNC|to undetectable cortisol|to undetectable cortisol
C0942490|T201|OSN|26536-3|LNC|to undetectable cortisol|to undetectable cortisol
C0942490|T201|LC|26536-3|LNC|to undetectable cortisol|to undetectable cortisol
C0942492|T201|LN|26539-7|LNC|glucose|glucose
C0942492|T201|MTH_LN|26539-7|LNC|glucose|glucose
C0942492|T201|OSN|26539-7|LNC|glucose|glucose
C0942492|T201|LC|26539-7|LNC|glucose|glucose
C0942494|T201|LN|26541-3|LNC|glucose|glucose
C0942494|T201|MTH_LN|26541-3|LNC|glucose|glucose
C0942494|T201|OSN|26541-3|LNC|glucose|glucose
C0942494|T201|LC|26541-3|LNC|glucose|glucose
C0942496|T201|LN|26543-9|LNC|glucose|glucose
C0942496|T201|MTH_LN|26543-9|LNC|glucose|glucose
C0942496|T201|OSN|26543-9|LNC|glucose|glucose
C0942496|T201|LC|26543-9|LNC|glucose|glucose
C0942497|T201|LN|26544-7|LNC|glucose|glucose
C0942497|T201|MTH_LN|26544-7|LNC|glucose|glucose
C0942497|T201|OSN|26544-7|LNC|glucose|glucose
C0942497|T201|LC|26544-7|LNC|glucose|glucose
C0942506|T201|LN|26554-6|LNC|glucose|glucose
C0942506|T201|OSN|26554-6|LNC|glucose|glucose
C0942506|T201|MTH_LN|26554-6|LNC|glucose|glucose
C0942506|T201|LC|26554-6|LNC|glucose|glucose
C0942507|T201|LN|26555-3|LNC|glucose|glucose
C0942507|T201|MTH_LN|26555-3|LNC|glucose|glucose
C0942507|T201|OSN|26555-3|LNC|glucose|glucose
C0942507|T201|LC|26555-3|LNC|glucose|glucose
C0942546|T201|LN|26604-9|LNC|beta-alanine|beta-alanine
C0942546|T201|MTH_LN|26604-9|LNC|beta-alanine|beta-alanine
C0942546|T201|OSN|26604-9|LNC|beta-alanine|beta-alanine
C0942546|T201|LC|26604-9|LNC|beta-alanine|beta-alanine
C0942549|T201|LN|26607-2|LNC|cystathionine|cystathionine
C0942549|T201|MTH_LN|26607-2|LNC|cystathionine|cystathionine
C0942549|T201|OSN|26607-2|LNC|cystathionine|cystathionine
C0942549|T201|LC|26607-2|LNC|cystathionine|cystathionine
C0942549|T201|LN|26607-2|LNC|sulfur amino acid metabolism|sulfur amino acid metabolism
C0942549|T201|MTH_LN|26607-2|LNC|sulfur amino acid metabolism|sulfur amino acid metabolism
C0942549|T201|OSN|26607-2|LNC|sulfur amino acid metabolism|sulfur amino acid metabolism
C0942549|T201|LC|26607-2|LNC|sulfur amino acid metabolism|sulfur amino acid metabolism
C0942549|T201|LN|26607-2|LNC|sulfur-containing amino acids|sulfur-containing amino acids
C0942549|T201|MTH_LN|26607-2|LNC|sulfur-containing amino acids|sulfur-containing amino acids
C0942549|T201|OSN|26607-2|LNC|sulfur-containing amino acids|sulfur-containing amino acids
C0942549|T201|LC|26607-2|LNC|sulfur-containing amino acids|sulfur-containing amino acids
C0942624|T201|LN|26695-7|LNC|glucose|glucose
C0942624|T201|MTH_LN|26695-7|LNC|glucose|glucose
C0942624|T201|OSN|26695-7|LNC|glucose|glucose
C0942624|T201|LC|26695-7|LNC|glucose|glucose
C0942660|T201|LN|26740-1|LNC|hydroxyproline|hydroxyproline
C0942660|T201|MTH_LN|26740-1|LNC|hydroxyproline|hydroxyproline
C0942660|T201|OSN|26740-1|LNC|hydroxyproline|hydroxyproline
C0942660|T201|LC|26740-1|LNC|hydroxyproline|hydroxyproline
C0942678|T201|LN|26759-1|LNC|naive T|naive T
C0942678|T201|OSN|26759-1|LNC|naive T|naive T
C0942678|T201|MTH_LN|26759-1|LNC|naive T|naive T
C0942678|T201|LC|26759-1|LNC|naive T|naive T
C0942678|T201|LN|26759-1|LNC|naive T cell|naive T cell
C0942678|T201|OSN|26759-1|LNC|naive T cell|naive T cell
C0942678|T201|MTH_LN|26759-1|LNC|naive T cell|naive T cell
C0942678|T201|LC|26759-1|LNC|naive T cell|naive T cell
C0942692|T201|LN|26778-1|LNC|glucose|glucose
C0942692|T201|MTH_LN|26778-1|LNC|glucose|glucose
C0942692|T201|OSN|26778-1|LNC|glucose|glucose
C0942692|T201|LC|26778-1|LNC|glucose|glucose
C0942693|T201|LN|26780-7|LNC|glucose|glucose
C0942693|T201|MTH_LN|26780-7|LNC|glucose|glucose
C0942693|T201|OSN|26780-7|LNC|glucose|glucose
C0942693|T201|LC|26780-7|LNC|glucose|glucose
C0942694|T201|LN|26783-1|LNC|glucose|glucose
C0942694|T201|MTH_LN|26783-1|LNC|glucose|glucose
C0942694|T201|OSN|26783-1|LNC|glucose|glucose
C0942694|T201|LC|26783-1|LNC|glucose|glucose
C0942723|T201|LN|26817-7|LNC|glucose|glucose
C0942723|T201|MTH_LN|26817-7|LNC|glucose|glucose
C0942723|T201|OSN|26817-7|LNC|glucose|glucose
C0942723|T201|LC|26817-7|LNC|glucose|glucose
C0942729|T201|LN|26823-5|LNC|luteinizing|luteinizing
C0942729|T201|OSN|26823-5|LNC|luteinizing|luteinizing
C0942729|T201|MTH_LN|26823-5|LNC|luteinizing|luteinizing
C0942729|T201|LC|26823-5|LNC|luteinizing|luteinizing
C0942729|T201|LN|26823-5|LNC|LH|LH
C0942729|T201|OSN|26823-5|LNC|LH|LH
C0942729|T201|MTH_LN|26823-5|LNC|LH|LH
C0942729|T201|LC|26823-5|LNC|LH|LH
C0942729|T201|LN|26823-5|LNC|luteinising|luteinising
C0942729|T201|OSN|26823-5|LNC|luteinising|luteinising
C0942729|T201|MTH_LN|26823-5|LNC|luteinising|luteinising
C0942729|T201|LC|26823-5|LNC|luteinising|luteinising
C0942745|T201|LN|26843-3|LNC|cystine|cystine
C0942745|T201|MTH_LN|26843-3|LNC|cystine|cystine
C0942745|T201|OSN|26843-3|LNC|cystine|cystine
C0942745|T201|LC|26843-3|LNC|cystine|cystine
C0942751|T201|LN|26853-2|LNC|glucose|glucose
C0942751|T201|MTH_LN|26853-2|LNC|glucose|glucose
C0942751|T201|OSN|26853-2|LNC|glucose|glucose
C0942751|T201|LC|26853-2|LNC|glucose|glucose
C0942752|T201|LN|26854-0|LNC|glucose|glucose
C0942752|T201|MTH_LN|26854-0|LNC|glucose|glucose
C0942752|T201|OSN|26854-0|LNC|glucose|glucose
C0942752|T201|LC|26854-0|LNC|glucose|glucose
C0942783|T201|LN|26888-8|LNC|sulfate|sulfate
C0942783|T201|MTH_LN|26888-8|LNC|sulfate|sulfate
C0942783|T201|OSN|26888-8|LNC|sulfate|sulfate
C0942783|T201|LC|26888-8|LNC|sulfate|sulfate
C0942784|T201|LN|26889-6|LNC|sulfate|sulfate
C0942784|T201|MTH_LN|26889-6|LNC|sulfate|sulfate
C0942784|T201|OSN|26889-6|LNC|sulfate|sulfate
C0942784|T201|LC|26889-6|LNC|sulfate|sulfate
C0942947|T201|LN|27088-4|LNC|folate metabolism|folate metabolism
C0942947|T201|MTH_LN|27088-4|LNC|folate metabolism|folate metabolism
C0942947|T201|OSN|27088-4|LNC|folate metabolism|folate metabolism
C0942947|T201|LC|27088-4|LNC|folate metabolism|folate metabolism
C0943117|T201|LN|27296-3|LNC|arginine|arginine
C0943117|T201|MTH_LN|27296-3|LNC|arginine|arginine
C0943117|T201|OSN|27296-3|LNC|arginine|arginine
C0943117|T201|LC|27296-3|LNC|arginine|arginine
C0943118|T201|LN|27298-9|LNC|Protein|Protein
C0943118|T201|MTH_LN|27298-9|LNC|Protein|Protein
C0943118|T201|OSN|27298-9|LNC|Protein|Protein
C0943118|T201|LC|27298-9|LNC|Protein|Protein
C0943152|T201|LN|27340-9|LNC|HDL cholesterol|HDL cholesterol
C0943152|T201|MTH_LN|27340-9|LNC|HDL cholesterol|HDL cholesterol
C0943152|T201|OSN|27340-9|LNC|HDL cholesterol|HDL cholesterol
C0943152|T201|LC|27340-9|LNC|HDL cholesterol|HDL cholesterol
C0943152|T201|LN|27340-9|LNC|HDL|HDL
C0943152|T201|MTH_LN|27340-9|LNC|HDL|HDL
C0943152|T201|OSN|27340-9|LNC|HDL|HDL
C0943152|T201|LC|27340-9|LNC|HDL|HDL
C0943152|T201|LN|27340-9|LNC|high-density lipoprotein|high-density lipoprotein
C0943152|T201|MTH_LN|27340-9|LNC|high-density lipoprotein|high-density lipoprotein
C0943152|T201|OSN|27340-9|LNC|high-density lipoprotein|high-density lipoprotein
C0943152|T201|LC|27340-9|LNC|high-density lipoprotein|high-density lipoprotein
C0943208|T201|LN|27408-4|LNC|C-peptide|C-peptide
C0943208|T201|MTH_LN|27408-4|LNC|C-peptide|C-peptide
C0943208|T201|OSN|27408-4|LNC|C-peptide|C-peptide
C0943208|T201|LC|27408-4|LNC|C-peptide|C-peptide
C0943208|T201|LN|27408-4|LNC|C peptide|C peptide
C0943208|T201|MTH_LN|27408-4|LNC|C peptide|C peptide
C0943208|T201|OSN|27408-4|LNC|C peptide|C peptide
C0943208|T201|LC|27408-4|LNC|C peptide|C peptide
C0943219|T201|LN|27421-7|LNC|C-peptide|C-peptide
C0943219|T201|MTH_LN|27421-7|LNC|C-peptide|C-peptide
C0943219|T201|OSN|27421-7|LNC|C-peptide|C-peptide
C0943219|T201|LC|27421-7|LNC|C-peptide|C-peptide
C0943219|T201|LN|27421-7|LNC|C peptide|C peptide
C0943219|T201|MTH_LN|27421-7|LNC|C peptide|C peptide
C0943219|T201|OSN|27421-7|LNC|C peptide|C peptide
C0943219|T201|LC|27421-7|LNC|C peptide|C peptide
C0943506|T201|LN|27811-9|LNC|antithrombin III|antithrombin III
C0943506|T201|OSN|27811-9|LNC|antithrombin III|antithrombin III
C0943506|T201|MTH_LN|27811-9|LNC|antithrombin III|antithrombin III
C0943506|T201|LC|27811-9|LNC|antithrombin III|antithrombin III
C0943506|T201|LN|27811-9|LNC|antithrombin III activity|antithrombin III activity
C0943506|T201|OSN|27811-9|LNC|antithrombin III activity|antithrombin III activity
C0943506|T201|MTH_LN|27811-9|LNC|antithrombin III activity|antithrombin III activity
C0943506|T201|LC|27811-9|LNC|antithrombin III activity|antithrombin III activity
C0943529|T201|LN|27839-0|LNC|C-peptide|C-peptide
C0943529|T201|MTH_LN|27839-0|LNC|C-peptide|C-peptide
C0943529|T201|OSN|27839-0|LNC|C-peptide|C-peptide
C0943529|T201|LC|27839-0|LNC|C-peptide|C-peptide
C0943529|T201|LN|27839-0|LNC|C peptide|C peptide
C0943529|T201|MTH_LN|27839-0|LNC|C peptide|C peptide
C0943529|T201|OSN|27839-0|LNC|C peptide|C peptide
C0943529|T201|LC|27839-0|LNC|C peptide|C peptide
C0943537|T201|LN|27848-1|LNC|luteinizing|luteinizing
C0943537|T201|MTH_LN|27848-1|LNC|luteinizing|luteinizing
C0943537|T201|OSN|27848-1|LNC|luteinizing|luteinizing
C0943537|T201|LC|27848-1|LNC|luteinizing|luteinizing
C0943537|T201|LN|27848-1|LNC|LH|LH
C0943537|T201|MTH_LN|27848-1|LNC|LH|LH
C0943537|T201|OSN|27848-1|LNC|LH|LH
C0943537|T201|LC|27848-1|LNC|LH|LH
C0943537|T201|LN|27848-1|LNC|luteinising|luteinising
C0943537|T201|MTH_LN|27848-1|LNC|luteinising|luteinising
C0943537|T201|OSN|27848-1|LNC|luteinising|luteinising
C0943537|T201|LC|27848-1|LNC|luteinising|luteinising
C0943540|T201|LN|27851-5|LNC|luteinizing|luteinizing
C0943540|T201|MTH_LN|27851-5|LNC|luteinizing|luteinizing
C0943540|T201|OSN|27851-5|LNC|luteinizing|luteinizing
C0943540|T201|LC|27851-5|LNC|luteinizing|luteinizing
C0943540|T201|LN|27851-5|LNC|LH|LH
C0943540|T201|MTH_LN|27851-5|LNC|LH|LH
C0943540|T201|OSN|27851-5|LNC|LH|LH
C0943540|T201|LC|27851-5|LNC|LH|LH
C0943540|T201|LN|27851-5|LNC|luteinising|luteinising
C0943540|T201|MTH_LN|27851-5|LNC|luteinising|luteinising
C0943540|T201|OSN|27851-5|LNC|luteinising|luteinising
C0943540|T201|LC|27851-5|LNC|luteinising|luteinising
C0943542|T201|LN|27853-1|LNC|luteinizing|luteinizing
C0943542|T201|MTH_LN|27853-1|LNC|luteinizing|luteinizing
C0943542|T201|OSN|27853-1|LNC|luteinizing|luteinizing
C0943542|T201|LC|27853-1|LNC|luteinizing|luteinizing
C0943542|T201|LN|27853-1|LNC|LH|LH
C0943542|T201|MTH_LN|27853-1|LNC|LH|LH
C0943542|T201|OSN|27853-1|LNC|LH|LH
C0943542|T201|LC|27853-1|LNC|LH|LH
C0943542|T201|LN|27853-1|LNC|luteinising|luteinising
C0943542|T201|MTH_LN|27853-1|LNC|luteinising|luteinising
C0943542|T201|OSN|27853-1|LNC|luteinising|luteinising
C0943542|T201|LC|27853-1|LNC|luteinising|luteinising
C0943543|T201|LN|27854-9|LNC|luteinizing|luteinizing
C0943543|T201|MTH_LN|27854-9|LNC|luteinizing|luteinizing
C0943543|T201|OSN|27854-9|LNC|luteinizing|luteinizing
C0943543|T201|LC|27854-9|LNC|luteinizing|luteinizing
C0943543|T201|LN|27854-9|LNC|LH|LH
C0943543|T201|MTH_LN|27854-9|LNC|LH|LH
C0943543|T201|OSN|27854-9|LNC|LH|LH
C0943543|T201|LC|27854-9|LNC|LH|LH
C0943543|T201|LN|27854-9|LNC|luteinising|luteinising
C0943543|T201|MTH_LN|27854-9|LNC|luteinising|luteinising
C0943543|T201|OSN|27854-9|LNC|luteinising|luteinising
C0943543|T201|LC|27854-9|LNC|luteinising|luteinising
C0943544|T201|LN|27855-6|LNC|luteinizing|luteinizing
C0943544|T201|MTH_LN|27855-6|LNC|luteinizing|luteinizing
C0943544|T201|OSN|27855-6|LNC|luteinizing|luteinizing
C0943544|T201|LC|27855-6|LNC|luteinizing|luteinizing
C0943544|T201|LN|27855-6|LNC|LH|LH
C0943544|T201|MTH_LN|27855-6|LNC|LH|LH
C0943544|T201|OSN|27855-6|LNC|LH|LH
C0943544|T201|LC|27855-6|LNC|LH|LH
C0943544|T201|LN|27855-6|LNC|luteinising|luteinising
C0943544|T201|MTH_LN|27855-6|LNC|luteinising|luteinising
C0943544|T201|OSN|27855-6|LNC|luteinising|luteinising
C0943544|T201|LC|27855-6|LNC|luteinising|luteinising
C0943547|T201|LN|27858-0|LNC|luteinizing|luteinizing
C0943547|T201|MTH_LN|27858-0|LNC|luteinizing|luteinizing
C0943547|T201|OSN|27858-0|LNC|luteinizing|luteinizing
C0943547|T201|LC|27858-0|LNC|luteinizing|luteinizing
C0943547|T201|LN|27858-0|LNC|LH|LH
C0943547|T201|MTH_LN|27858-0|LNC|LH|LH
C0943547|T201|OSN|27858-0|LNC|LH|LH
C0943547|T201|LC|27858-0|LNC|LH|LH
C0943547|T201|LN|27858-0|LNC|luteinising|luteinising
C0943547|T201|MTH_LN|27858-0|LNC|luteinising|luteinising
C0943547|T201|OSN|27858-0|LNC|luteinising|luteinising
C0943547|T201|LC|27858-0|LNC|luteinising|luteinising
C0943569|T201|LN|27883-8|LNC|luteinizing|luteinizing
C0943569|T201|MTH_LN|27883-8|LNC|luteinizing|luteinizing
C0943569|T201|OSN|27883-8|LNC|luteinizing|luteinizing
C0943569|T201|LC|27883-8|LNC|luteinizing|luteinizing
C0943569|T201|LN|27883-8|LNC|LH|LH
C0943569|T201|MTH_LN|27883-8|LNC|LH|LH
C0943569|T201|OSN|27883-8|LNC|LH|LH
C0943569|T201|LC|27883-8|LNC|LH|LH
C0943569|T201|LN|27883-8|LNC|luteinising|luteinising
C0943569|T201|MTH_LN|27883-8|LNC|luteinising|luteinising
C0943569|T201|OSN|27883-8|LNC|luteinising|luteinising
C0943569|T201|LC|27883-8|LNC|luteinising|luteinising
C0943617|T201|LN|27941-4|LNC|CSF lactate|CSF lactate
C0943617|T201|MTH_LN|27941-4|LNC|CSF lactate|CSF lactate
C0943617|T201|OSN|27941-4|LNC|CSF lactate|CSF lactate
C0943617|T201|LC|27941-4|LNC|CSF lactate|CSF lactate
C0943617|T201|LN|27941-4|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C0943617|T201|MTH_LN|27941-4|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C0943617|T201|OSN|27941-4|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C0943617|T201|LC|27941-4|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C0943617|T201|LN|27941-4|LNC|CSF lactic acid|CSF lactic acid
C0943617|T201|MTH_LN|27941-4|LNC|CSF lactic acid|CSF lactic acid
C0943617|T201|OSN|27941-4|LNC|CSF lactic acid|CSF lactic acid
C0943617|T201|LC|27941-4|LNC|CSF lactic acid|CSF lactic acid
C0943623|T201|LN|27949-7|LNC|lactate|lactate
C0943623|T201|MTH_LN|27949-7|LNC|lactate|lactate
C0943623|T201|OSN|27949-7|LNC|lactate|lactate
C0943623|T201|LC|27949-7|LNC|lactate|lactate
C0943628|T201|LN|27955-4|LNC|lactate|lactate
C0943628|T201|MTH_LN|27955-4|LNC|lactate|lactate
C0943628|T201|OSN|27955-4|LNC|lactate|lactate
C0943628|T201|LC|27955-4|LNC|lactate|lactate
C0943634|T201|LN|27961-2|LNC|lactate|lactate
C0943634|T201|MTH_LN|27961-2|LNC|lactate|lactate
C0943634|T201|OSN|27961-2|LNC|lactate|lactate
C0943634|T201|LC|27961-2|LNC|lactate|lactate
C0943649|T201|LN|27976-0|LNC|lactate|lactate
C0943649|T201|MTH_LN|27976-0|LNC|lactate|lactate
C0943649|T201|OSN|27976-0|LNC|lactate|lactate
C0943649|T201|LC|27976-0|LNC|lactate|lactate
C0944138|T201|LN|28545-2|LNC|homeostasis|homeostasis
C0944138|T201|MTH_LN|28545-2|LNC|homeostasis|homeostasis
C0944138|T201|OSN|28545-2|LNC|homeostasis|homeostasis
C0944138|T201|LC|28545-2|LNC|homeostasis|homeostasis
C0944182|T201|LN|28595-7|LNC|taurine|taurine
C0944182|T201|MTH_LN|28595-7|LNC|taurine|taurine
C0944182|T201|OSN|28595-7|LNC|taurine|taurine
C0944182|T201|LC|28595-7|LNC|taurine|taurine
C0944184|T201|LN|28597-3|LNC|carnosine|carnosine
C0944184|T201|MTH_LN|28597-3|LNC|carnosine|carnosine
C0944184|T201|OSN|28597-3|LNC|carnosine|carnosine
C0944184|T201|LC|28597-3|LNC|carnosine|carnosine
C0944185|T201|LN|28599-9|LNC|cystathionine|cystathionine
C0944185|T201|MTH_LN|28599-9|LNC|cystathionine|cystathionine
C0944185|T201|OSN|28599-9|LNC|cystathionine|cystathionine
C0944185|T201|LC|28599-9|LNC|cystathionine|cystathionine
C0944189|T201|LN|28604-7|LNC|phosphoethanolamine|phosphoethanolamine
C0944189|T201|MTH_LN|28604-7|LNC|phosphoethanolamine|phosphoethanolamine
C0944189|T201|OSN|28604-7|LNC|phosphoethanolamine|phosphoethanolamine
C0944189|T201|LC|28604-7|LNC|phosphoethanolamine|phosphoethanolamine
C0944192|T201|LN|28608-8|LNC|tryptophan|tryptophan
C0944192|T201|MTH_LN|28608-8|LNC|tryptophan|tryptophan
C0944192|T201|OSN|28608-8|LNC|tryptophan|tryptophan
C0944192|T201|LC|28608-8|LNC|tryptophan|tryptophan
C0944223|T201|LN|28642-7|LNC|oxygen|oxygen
C0944223|T201|LC|28642-7|LNC|oxygen|oxygen
C0944223|T201|MTH_LN|28642-7|LNC|oxygen|oxygen
C0944223|T201|OSN|28642-7|LNC|oxygen|oxygen
C0944742|T201|LN|29261-5|LNC|lymphocyte count|lymphocyte count
C0944742|T201|OSN|29261-5|LNC|lymphocyte count|lymphocyte count
C0944742|T201|MTH_LN|29261-5|LNC|lymphocyte count|lymphocyte count
C0944742|T201|LC|29261-5|LNC|lymphocyte count|lymphocyte count
C0944742|T201|LN|29261-5|LNC|lymphocyte number|lymphocyte number
C0944742|T201|OSN|29261-5|LNC|lymphocyte number|lymphocyte number
C0944742|T201|MTH_LN|29261-5|LNC|lymphocyte number|lymphocyte number
C0944742|T201|LC|29261-5|LNC|lymphocyte number|lymphocyte number
C0944742|T201|LN|29261-5|LNC|lymphocyte counts|lymphocyte counts
C0944742|T201|OSN|29261-5|LNC|lymphocyte counts|lymphocyte counts
C0944742|T201|MTH_LN|29261-5|LNC|lymphocyte counts|lymphocyte counts
C0944742|T201|LC|29261-5|LNC|lymphocyte counts|lymphocyte counts
C0944742|T201|LN|29261-5|LNC|lymphocytes|lymphocytes
C0944742|T201|OSN|29261-5|LNC|lymphocytes|lymphocytes
C0944742|T201|MTH_LN|29261-5|LNC|lymphocytes|lymphocytes
C0944742|T201|LC|29261-5|LNC|lymphocytes|lymphocytes
C0944742|T201|LN|29261-5|LNC|numberslymphocytes|numberslymphocytes
C0944742|T201|OSN|29261-5|LNC|numberslymphocytes|numberslymphocytes
C0944742|T201|MTH_LN|29261-5|LNC|numberslymphocytes|numberslymphocytes
C0944742|T201|LC|29261-5|LNC|numberslymphocytes|numberslymphocytes
C0944746|T201|LN|29265-6|LNC|calcium|calcium
C0944746|T201|MTH_LN|29265-6|LNC|calcium|calcium
C0944746|T201|OSN|29265-6|LNC|calcium|calcium
C0944746|T201|LC|29265-6|LNC|calcium|calcium
C0944746|T201|LN|29265-6|LNC|calcium homeostasis|calcium homeostasis
C0944746|T201|MTH_LN|29265-6|LNC|calcium homeostasis|calcium homeostasis
C0944746|T201|OSN|29265-6|LNC|calcium homeostasis|calcium homeostasis
C0944746|T201|LC|29265-6|LNC|calcium homeostasis|calcium homeostasis
C0944796|T201|LN|29330-8|LNC|glucose|glucose
C0944796|T201|MTH_LN|29330-8|LNC|glucose|glucose
C0944796|T201|OSN|29330-8|LNC|glucose|glucose
C0944796|T201|LC|29330-8|LNC|glucose|glucose
C0944797|T201|LN|29331-6|LNC|glucose|glucose
C0944797|T201|MTH_LN|29331-6|LNC|glucose|glucose
C0944797|T201|OSN|29331-6|LNC|glucose|glucose
C0944797|T201|LC|29331-6|LNC|glucose|glucose
C0944798|T201|LN|29332-4|LNC|glucose|glucose
C0944798|T201|OSN|29332-4|LNC|glucose|glucose
C0944798|T201|MTH_LN|29332-4|LNC|glucose|glucose
C0944798|T201|LC|29332-4|LNC|glucose|glucose
C0945006|T201|LN|29572-5|LNC|phenylalanine metabolism|phenylalanine metabolism
C0945006|T201|LC|29572-5|LNC|phenylalanine metabolism|phenylalanine metabolism
C0945006|T201|MTH_LN|29572-5|LNC|phenylalanine metabolism|phenylalanine metabolism
C0945006|T201|OSN|29572-5|LNC|phenylalanine metabolism|phenylalanine metabolism
C0945007|T201|LN|29573-3|LNC|phenylalanine metabolism|phenylalanine metabolism
C0945007|T201|LC|29573-3|LNC|phenylalanine metabolism|phenylalanine metabolism
C0945007|T201|MTH_LN|29573-3|LNC|phenylalanine metabolism|phenylalanine metabolism
C0945007|T201|OSN|29573-3|LNC|phenylalanine metabolism|phenylalanine metabolism
C0945240|T201|LN|25573-7|LNC|C-peptide|C-peptide
C0945240|T201|MTH_LN|25573-7|LNC|C-peptide|C-peptide
C0945240|T201|OSN|25573-7|LNC|C-peptide|C-peptide
C0945240|T201|LC|25573-7|LNC|C-peptide|C-peptide
C0945240|T201|LN|25573-7|LNC|C peptide|C peptide
C0945240|T201|MTH_LN|25573-7|LNC|C peptide|C peptide
C0945240|T201|OSN|25573-7|LNC|C peptide|C peptide
C0945240|T201|LC|25573-7|LNC|C peptide|C peptide
C0945241|T201|LN|25574-5|LNC|C-peptide|C-peptide
C0945241|T201|MTH_LN|25574-5|LNC|C-peptide|C-peptide
C0945241|T201|OSN|25574-5|LNC|C-peptide|C-peptide
C0945241|T201|LC|25574-5|LNC|C-peptide|C-peptide
C0945241|T201|LN|25574-5|LNC|C peptide|C peptide
C0945241|T201|MTH_LN|25574-5|LNC|C peptide|C peptide
C0945241|T201|OSN|25574-5|LNC|C peptide|C peptide
C0945241|T201|LC|25574-5|LNC|C peptide|C peptide
C0945252|T201|LN|25666-9|LNC|glucose|glucose
C0945252|T201|OSN|25666-9|LNC|glucose|glucose
C0945252|T201|MTH_LN|25666-9|LNC|glucose|glucose
C0945252|T201|LC|25666-9|LNC|glucose|glucose
C0945281|T201|LN|25900-2|LNC|lactate|lactate
C0945281|T201|OSN|25900-2|LNC|lactate|lactate
C0945281|T201|MTH_LN|25900-2|LNC|lactate|lactate
C0945281|T201|LC|25900-2|LNC|lactate|lactate
C0945282|T201|LN|25903-6|LNC|lactate|lactate
C0945282|T201|OSN|25903-6|LNC|lactate|lactate
C0945282|T201|MTH_LN|25903-6|LNC|lactate|lactate
C0945282|T201|LC|25903-6|LNC|lactate|lactate
C0945289|T201|LN|25946-5|LNC|luteinizing|luteinizing
C0945289|T201|MTH_LN|25946-5|LNC|luteinizing|luteinizing
C0945289|T201|OSN|25946-5|LNC|luteinizing|luteinizing
C0945289|T201|LC|25946-5|LNC|luteinizing|luteinizing
C0945289|T201|LN|25946-5|LNC|LH|LH
C0945289|T201|MTH_LN|25946-5|LNC|LH|LH
C0945289|T201|OSN|25946-5|LNC|LH|LH
C0945289|T201|LC|25946-5|LNC|LH|LH
C0945289|T201|LN|25946-5|LNC|luteinising|luteinising
C0945289|T201|MTH_LN|25946-5|LNC|luteinising|luteinising
C0945289|T201|OSN|25946-5|LNC|luteinising|luteinising
C0945289|T201|LC|25946-5|LNC|luteinising|luteinising
C0945354|T201|LN|26450-7|LNC|eosinophil count|eosinophil count
C0945354|T201|OSN|26450-7|LNC|eosinophil count|eosinophil count
C0945354|T201|MTH_LN|26450-7|LNC|eosinophil count|eosinophil count
C0945354|T201|LC|26450-7|LNC|eosinophil count|eosinophil count
C0945354|T201|LN|26450-7|LNC|eosinophil morphology|eosinophil morphology
C0945354|T201|OSN|26450-7|LNC|eosinophil morphology|eosinophil morphology
C0945354|T201|MTH_LN|26450-7|LNC|eosinophil morphology|eosinophil morphology
C0945354|T201|LC|26450-7|LNC|eosinophil morphology|eosinophil morphology
C0945354|T201|LN|26450-7|LNC|eosinophils|eosinophils
C0945354|T201|OSN|26450-7|LNC|eosinophils|eosinophils
C0945354|T201|MTH_LN|26450-7|LNC|eosinophils|eosinophils
C0945354|T201|LC|26450-7|LNC|eosinophils|eosinophils
C0945357|T201|LN|26464-8|LNC|white count|white count
C0945357|T201|OSN|26464-8|LNC|white count|white count
C0945357|T201|MTH_LN|26464-8|LNC|white count|white count
C0945357|T201|LC|26464-8|LNC|white count|white count
C0945357|T201|LN|26464-8|LNC|leukocyte number|leukocyte number
C0945357|T201|OSN|26464-8|LNC|leukocyte number|leukocyte number
C0945357|T201|MTH_LN|26464-8|LNC|leukocyte number|leukocyte number
C0945357|T201|LC|26464-8|LNC|leukocyte number|leukocyte number
C0945357|T201|LN|26464-8|LNC|white cell count|white cell count
C0945357|T201|OSN|26464-8|LNC|white cell count|white cell count
C0945357|T201|MTH_LN|26464-8|LNC|white cell count|white cell count
C0945357|T201|LC|26464-8|LNC|white cell count|white cell count
C0945357|T201|LN|26464-8|LNC|leukocyte count|leukocyte count
C0945357|T201|OSN|26464-8|LNC|leukocyte count|leukocyte count
C0945357|T201|MTH_LN|26464-8|LNC|leukocyte count|leukocyte count
C0945357|T201|LC|26464-8|LNC|leukocyte count|leukocyte count
C0945362|T201|LN|26507-4|LNC|granulocyte precursors|granulocyte precursors
C0945362|T201|OSN|26507-4|LNC|granulocyte precursors|granulocyte precursors
C0945362|T201|MTH_LN|26507-4|LNC|granulocyte precursors|granulocyte precursors
C0945362|T201|LC|26507-4|LNC|granulocyte precursors|granulocyte precursors
C0945367|T201|LN|26533-0|LNC|cortisol|cortisol
C0945367|T201|MTH_LN|26533-0|LNC|cortisol|cortisol
C0945367|T201|OSN|26533-0|LNC|cortisol|cortisol
C0945367|T201|LC|26533-0|LNC|cortisol|cortisol
C0945367|T201|LN|26533-0|LNC|cortisol low|cortisol low
C0945367|T201|MTH_LN|26533-0|LNC|cortisol low|cortisol low
C0945367|T201|OSN|26533-0|LNC|cortisol low|cortisol low
C0945367|T201|LC|26533-0|LNC|cortisol low|cortisol low
C0945367|T201|LN|26533-0|LNC|to undetectable cortisol|to undetectable cortisol
C0945367|T201|MTH_LN|26533-0|LNC|to undetectable cortisol|to undetectable cortisol
C0945367|T201|OSN|26533-0|LNC|to undetectable cortisol|to undetectable cortisol
C0945367|T201|LC|26533-0|LNC|to undetectable cortisol|to undetectable cortisol
C0945403|T201|LN|26779-9|LNC|glucose|glucose
C0945403|T201|OSN|26779-9|LNC|glucose|glucose
C0945403|T201|MTH_LN|26779-9|LNC|glucose|glucose
C0945403|T201|LC|26779-9|LNC|glucose|glucose
C0945403|T201|LN|26779-9|LNC|glucose homeostasis|glucose homeostasis
C0945403|T201|OSN|26779-9|LNC|glucose homeostasis|glucose homeostasis
C0945403|T201|MTH_LN|26779-9|LNC|glucose homeostasis|glucose homeostasis
C0945403|T201|LC|26779-9|LNC|glucose homeostasis|glucose homeostasis
C0945404|T201|LN|26782-3|LNC|glucose|glucose
C0945404|T201|MTH_LN|26782-3|LNC|glucose|glucose
C0945404|T201|OSN|26782-3|LNC|glucose|glucose
C0945404|T201|LC|26782-3|LNC|glucose|glucose
C0945434|T201|LN|26971-2|LNC|Smooth muscle antibody|Smooth muscle antibody
C0945434|T201|MTH_LN|26971-2|LNC|Smooth muscle antibody|Smooth muscle antibody
C0945434|T201|OSN|26971-2|LNC|Smooth muscle antibody|Smooth muscle antibody
C0945434|T201|LC|26971-2|LNC|Smooth muscle antibody|Smooth muscle antibody
C0945434|T201|LN|26971-2|LNC|Anti-smooth muscle antibody|Anti-smooth muscle antibody
C0945434|T201|MTH_LN|26971-2|LNC|Anti-smooth muscle antibody|Anti-smooth muscle antibody
C0945434|T201|OSN|26971-2|LNC|Anti-smooth muscle antibody|Anti-smooth muscle antibody
C0945434|T201|LC|26971-2|LNC|Anti-smooth muscle antibody|Anti-smooth muscle antibody
C0945506|T201|LN|27432-4|LNC|glucose|glucose
C0945506|T201|MTH_LN|27432-4|LNC|glucose|glucose
C0945506|T201|OSN|27432-4|LNC|glucose|glucose
C0945506|T201|LC|27432-4|LNC|glucose|glucose
C0945549|T201|LN|27884-6|LNC|luteinizing|luteinizing
C0945549|T201|MTH_LN|27884-6|LNC|luteinizing|luteinizing
C0945549|T201|OSN|27884-6|LNC|luteinizing|luteinizing
C0945549|T201|LC|27884-6|LNC|luteinizing|luteinizing
C0945549|T201|LN|27884-6|LNC|LH|LH
C0945549|T201|MTH_LN|27884-6|LNC|LH|LH
C0945549|T201|OSN|27884-6|LNC|LH|LH
C0945549|T201|LC|27884-6|LNC|LH|LH
C0945549|T201|LN|27884-6|LNC|luteinising|luteinising
C0945549|T201|MTH_LN|27884-6|LNC|luteinising|luteinising
C0945549|T201|OSN|27884-6|LNC|luteinising|luteinising
C0945549|T201|LC|27884-6|LNC|luteinising|luteinising
C0945557|T201|LN|27946-3|LNC|lactate|lactate
C0945557|T201|MTH_LN|27946-3|LNC|lactate|lactate
C0945557|T201|OSN|27946-3|LNC|lactate|lactate
C0945557|T201|LC|27946-3|LNC|lactate|lactate
C0945564|T201|LN|28007-3|LNC|urobilinogen|urobilinogen
C0945564|T201|MTH_LN|28007-3|LNC|urobilinogen|urobilinogen
C0945564|T201|OSN|28007-3|LNC|urobilinogen|urobilinogen
C0945564|T201|LC|28007-3|LNC|urobilinogen|urobilinogen
C0945632|T201|LN|28601-3|LNC|hydroxyproline|hydroxyproline
C0945632|T201|MTH_LN|28601-3|LNC|hydroxyproline|hydroxyproline
C0945632|T201|OSN|28601-3|LNC|hydroxyproline|hydroxyproline
C0945632|T201|LC|28601-3|LNC|hydroxyproline|hydroxyproline
C0945746|T201|LN|29412-4|LNC|glucose|glucose
C0945746|T201|MTH_LN|29412-4|LNC|glucose|glucose
C0945746|T201|OSN|29412-4|LNC|glucose|glucose
C0945746|T201|LC|29412-4|LNC|glucose|glucose
C0947220|T201|LN|26532-2|LNC|cortisol|cortisol
C0947220|T201|MTH_LN|26532-2|LNC|cortisol|cortisol
C0947220|T201|OSN|26532-2|LNC|cortisol|cortisol
C0947220|T201|LC|26532-2|LNC|cortisol|cortisol
C0947220|T201|LN|26532-2|LNC|cortisol low|cortisol low
C0947220|T201|MTH_LN|26532-2|LNC|cortisol low|cortisol low
C0947220|T201|OSN|26532-2|LNC|cortisol low|cortisol low
C0947220|T201|LC|26532-2|LNC|cortisol low|cortisol low
C0947220|T201|LN|26532-2|LNC|to undetectable cortisol|to undetectable cortisol
C0947220|T201|MTH_LN|26532-2|LNC|to undetectable cortisol|to undetectable cortisol
C0947220|T201|OSN|26532-2|LNC|to undetectable cortisol|to undetectable cortisol
C0947220|T201|LC|26532-2|LNC|to undetectable cortisol|to undetectable cortisol
C0947224|T201|LN|26777-3|LNC|glucose|glucose
C0947224|T201|MTH_LN|26777-3|LNC|glucose|glucose
C0947224|T201|OSN|26777-3|LNC|glucose|glucose
C0947224|T201|LC|26777-3|LNC|glucose|glucose
C0947225|T201|LN|26781-5|LNC|glucose|glucose
C0947225|T201|MTH_LN|26781-5|LNC|glucose|glucose
C0947225|T201|OSN|26781-5|LNC|glucose|glucose
C0947225|T201|LC|26781-5|LNC|glucose|glucose
C0947235|T201|LN|27885-3|LNC|luteinizing|luteinizing
C0947235|T201|OSN|27885-3|LNC|luteinizing|luteinizing
C0947235|T201|MTH_LN|27885-3|LNC|luteinizing|luteinizing
C0947235|T201|LC|27885-3|LNC|luteinizing|luteinizing
C0947235|T201|LN|27885-3|LNC|LH|LH
C0947235|T201|OSN|27885-3|LNC|LH|LH
C0947235|T201|MTH_LN|27885-3|LNC|LH|LH
C0947235|T201|LC|27885-3|LNC|LH|LH
C0947235|T201|LN|27885-3|LNC|luteinising|luteinising
C0947235|T201|OSN|27885-3|LNC|luteinising|luteinising
C0947235|T201|MTH_LN|27885-3|LNC|luteinising|luteinising
C0947235|T201|LC|27885-3|LNC|luteinising|luteinising
C0947266|T201|LN|29329-0|LNC|glucose|glucose
C0947266|T201|MTH_LN|29329-0|LNC|glucose|glucose
C0947266|T201|OSN|29329-0|LNC|glucose|glucose
C0947266|T201|LC|29329-0|LNC|glucose|glucose
C0947495|T201|MTH_LN|14251-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C0947495|T201|LN|14251-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C0947495|T201|OSN|14251-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C0947495|T201|LC|14251-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C1113877|T201|LN|29960-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1113877|T201|OSN|29960-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1113877|T201|LC|29960-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1113877|T201|MTH_LN|29960-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1113951|T201|LN|30047-5|LNC|histidine|histidine
C1113951|T201|MTH_LN|30047-5|LNC|histidine|histidine
C1113951|T201|OSN|30047-5|LNC|histidine|histidine
C1113951|T201|LC|30047-5|LNC|histidine|histidine
C1113957|T201|LN|30057-4|LNC|threonine|threonine
C1113957|T201|MTH_LN|30057-4|LNC|threonine|threonine
C1113957|T201|OSN|30057-4|LNC|threonine|threonine
C1113957|T201|LC|30057-4|LNC|threonine|threonine
C1113962|T201|LN|30062-4|LNC|arginine|arginine
C1113962|T201|MTH_LN|30062-4|LNC|arginine|arginine
C1113962|T201|OSN|30062-4|LNC|arginine|arginine
C1113962|T201|LC|30062-4|LNC|arginine|arginine
C1113965|T201|LN|30065-7|LNC|cystine|cystine
C1113965|T201|MTH_LN|30065-7|LNC|cystine|cystine
C1113965|T201|OSN|30065-7|LNC|cystine|cystine
C1113965|T201|LC|30065-7|LNC|cystine|cystine
C1113966|T201|LN|30066-5|LNC|glycine|glycine
C1113966|T201|MTH_LN|30066-5|LNC|glycine|glycine
C1113966|T201|OSN|30066-5|LNC|glycine|glycine
C1113966|T201|LC|30066-5|LNC|glycine|glycine
C1114053|T201|LN|30166-3|LNC|thyroid stimulating|thyroid stimulating
C1114053|T201|MTH_LN|30166-3|LNC|thyroid stimulating|thyroid stimulating
C1114053|T201|OSN|30166-3|LNC|thyroid stimulating|thyroid stimulating
C1114053|T201|LC|30166-3|LNC|thyroid stimulating|thyroid stimulating
C1114053|T201|LN|30166-3|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C1114053|T201|MTH_LN|30166-3|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C1114053|T201|OSN|30166-3|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C1114053|T201|LC|30166-3|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C1114053|T201|LN|30166-3|LNC|TSH|TSH
C1114053|T201|MTH_LN|30166-3|LNC|TSH|TSH
C1114053|T201|OSN|30166-3|LNC|TSH|TSH
C1114053|T201|LC|30166-3|LNC|TSH|TSH
C1114053|T201|LN|30166-3|LNC|thyroid-stimulating|thyroid-stimulating
C1114053|T201|MTH_LN|30166-3|LNC|thyroid-stimulating|thyroid-stimulating
C1114053|T201|OSN|30166-3|LNC|thyroid-stimulating|thyroid-stimulating
C1114053|T201|LC|30166-3|LNC|thyroid-stimulating|thyroid-stimulating
C1114065|T201|LN|30180-4|LNC|basophil count|basophil count
C1114065|T201|OSN|30180-4|LNC|basophil count|basophil count
C1114065|T201|MTH_LN|30180-4|LNC|basophil count|basophil count
C1114065|T201|LC|30180-4|LNC|basophil count|basophil count
C1114076|T201|LN|30191-1|LNC|acylcarnitine|acylcarnitine
C1114076|T201|OSN|30191-1|LNC|acylcarnitine|acylcarnitine
C1114076|T201|MTH_LN|30191-1|LNC|acylcarnitine|acylcarnitine
C1114076|T201|LC|30191-1|LNC|acylcarnitine|acylcarnitine
C1114077|T201|LN|30192-9|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1114077|T201|MTH_LN|30192-9|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1114077|T201|LC|30192-9|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1114077|T201|OSN|30192-9|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1114078|T201|LN|30193-7|LNC|acylcarnitine|acylcarnitine
C1114078|T201|OSN|30193-7|LNC|acylcarnitine|acylcarnitine
C1114078|T201|LC|30193-7|LNC|acylcarnitine|acylcarnitine
C1114078|T201|MTH_LN|30193-7|LNC|acylcarnitine|acylcarnitine
C1114119|T201|LN|30241-4|LNC|lactate|lactate
C1114119|T201|MTH_LN|30241-4|LNC|lactate|lactate
C1114119|T201|OSN|30241-4|LNC|lactate|lactate
C1114119|T201|LC|30241-4|LNC|lactate|lactate
C1114120|T201|LN|30242-2|LNC|lactate|lactate
C1114120|T201|MTH_LN|30242-2|LNC|lactate|lactate
C1114120|T201|OSN|30242-2|LNC|lactate|lactate
C1114120|T201|LC|30242-2|LNC|lactate|lactate
C1114129|T201|LN|30251-3|LNC|glucose|glucose
C1114129|T201|MTH_LN|30251-3|LNC|glucose|glucose
C1114129|T201|OSN|30251-3|LNC|glucose|glucose
C1114129|T201|LC|30251-3|LNC|glucose|glucose
C1114130|T201|LN|30252-1|LNC|glucose|glucose
C1114130|T201|MTH_LN|30252-1|LNC|glucose|glucose
C1114130|T201|OSN|30252-1|LNC|glucose|glucose
C1114130|T201|LC|30252-1|LNC|glucose|glucose
C1114131|T201|LN|30253-9|LNC|glucose|glucose
C1114131|T201|MTH_LN|30253-9|LNC|glucose|glucose
C1114131|T201|OSN|30253-9|LNC|glucose|glucose
C1114131|T201|LC|30253-9|LNC|glucose|glucose
C1114140|T201|LN|30263-8|LNC|glucose|glucose
C1114140|T201|MTH_LN|30263-8|LNC|glucose|glucose
C1114140|T201|OSN|30263-8|LNC|glucose|glucose
C1114140|T201|LC|30263-8|LNC|glucose|glucose
C1114141|T201|LN|30265-3|LNC|glucose|glucose
C1114141|T201|MTH_LN|30265-3|LNC|glucose|glucose
C1114141|T201|OSN|30265-3|LNC|glucose|glucose
C1114141|T201|LC|30265-3|LNC|glucose|glucose
C1114142|T201|LN|30267-9|LNC|glucose|glucose
C1114142|T201|MTH_LN|30267-9|LNC|glucose|glucose
C1114142|T201|OSN|30267-9|LNC|glucose|glucose
C1114142|T201|LC|30267-9|LNC|glucose|glucose
C1114184|T201|LN|30313-1|LNC|hemoglobin|hemoglobin
C1114184|T201|MTH_LN|30313-1|LNC|hemoglobin|hemoglobin
C1114184|T201|OSN|30313-1|LNC|hemoglobin|hemoglobin
C1114184|T201|LC|30313-1|LNC|hemoglobin|hemoglobin
C1114209|T201|LN|30344-6|LNC|glucose|glucose
C1114209|T201|MTH_LN|30344-6|LNC|glucose|glucose
C1114209|T201|OSN|30344-6|LNC|glucose|glucose
C1114209|T201|LC|30344-6|LNC|glucose|glucose
C1114210|T201|LN|30345-3|LNC|glucose|glucose
C1114210|T201|MTH_LN|30345-3|LNC|glucose|glucose
C1114210|T201|OSN|30345-3|LNC|glucose|glucose
C1114210|T201|LC|30345-3|LNC|glucose|glucose
C1114247|T201|LN|30386-7|LNC|erythrocyte volume|erythrocyte volume
C1114247|T201|OSN|30386-7|LNC|erythrocyte volume|erythrocyte volume
C1114247|T201|MTH_LN|30386-7|LNC|erythrocyte volume|erythrocyte volume
C1114247|T201|LC|30386-7|LNC|erythrocyte volume|erythrocyte volume
C1114247|T201|LN|30386-7|LNC|mean corpuscular volume|mean corpuscular volume
C1114247|T201|OSN|30386-7|LNC|mean corpuscular volume|mean corpuscular volume
C1114247|T201|MTH_LN|30386-7|LNC|mean corpuscular volume|mean corpuscular volume
C1114247|T201|LC|30386-7|LNC|mean corpuscular volume|mean corpuscular volume
// C1114250|T201|LN|30391-7|LNC||
// C1114250|T201|OSN|30391-7|LNC||
// C1114250|T201|MTH_LN|30391-7|LNC||
// C1114250|T201|LC|30391-7|LNC||
C1114250|T201|LN|30391-7|LNC|occult|occult
C1114250|T201|OSN|30391-7|LNC|occult|occult
C1114250|T201|MTH_LN|30391-7|LNC|occult|occult
C1114250|T201|LC|30391-7|LNC|occult|occult
C1114256|T201|LN|30398-2|LNC|hematocrit|hematocrit
C1114256|T201|MTH_LN|30398-2|LNC|hematocrit|hematocrit
C1114256|T201|LC|30398-2|LNC|hematocrit|hematocrit
C1114256|T201|OSN|30398-2|LNC|hematocrit|hematocrit
C1114261|T201|LN|30405-5|LNC|neutrophil count|neutrophil count
C1114261|T201|OSN|30405-5|LNC|neutrophil count|neutrophil count
C1114261|T201|MTH_LN|30405-5|LNC|neutrophil count|neutrophil count
C1114261|T201|LC|30405-5|LNC|neutrophil count|neutrophil count
C1114261|T201|LN|30405-5|LNC|cytology|cytology
C1114261|T201|OSN|30405-5|LNC|cytology|cytology
C1114261|T201|MTH_LN|30405-5|LNC|cytology|cytology
C1114261|T201|LC|30405-5|LNC|cytology|cytology
C1114281|T201|LN|30428-7|LNC|erythrocyte volume|erythrocyte volume
C1114281|T201|OSN|30428-7|LNC|erythrocyte volume|erythrocyte volume
C1114281|T201|LC|30428-7|LNC|erythrocyte volume|erythrocyte volume
C1114281|T201|MTH_LN|30428-7|LNC|erythrocyte volume|erythrocyte volume
C1114281|T201|LN|30428-7|LNC|mean corpuscular volume|mean corpuscular volume
C1114281|T201|OSN|30428-7|LNC|mean corpuscular volume|mean corpuscular volume
C1114281|T201|LC|30428-7|LNC|mean corpuscular volume|mean corpuscular volume
C1114281|T201|MTH_LN|30428-7|LNC|mean corpuscular volume|mean corpuscular volume
C1114302|T201|LN|30451-9|LNC|neutrophil morphology|neutrophil morphology
C1114302|T201|OSN|30451-9|LNC|neutrophil morphology|neutrophil morphology
C1114302|T201|MTH_LN|30451-9|LNC|neutrophil morphology|neutrophil morphology
C1114302|T201|LC|30451-9|LNC|neutrophil morphology|neutrophil morphology
C1114363|T201|LN|30522-7|LNC|CRP|CRP
C1114363|T201|MTH_LN|30522-7|LNC|CRP|CRP
C1114363|T201|LC|30522-7|LNC|CRP|CRP
C1114363|T201|OSN|30522-7|LNC|CRP|CRP
C1114363|T201|LN|30522-7|LNC|Serum protein|Serum protein
C1114363|T201|MTH_LN|30522-7|LNC|Serum protein|Serum protein
C1114363|T201|LC|30522-7|LNC|Serum protein|Serum protein
C1114363|T201|OSN|30522-7|LNC|Serum protein|Serum protein
C1114363|T201|LN|30522-7|LNC|protein disease|protein disease
C1114363|T201|MTH_LN|30522-7|LNC|protein disease|protein disease
C1114363|T201|LC|30522-7|LNC|protein disease|protein disease
C1114363|T201|OSN|30522-7|LNC|protein disease|protein disease
C1114363|T201|LN|30522-7|LNC|C-reactive protein|C-reactive protein
C1114363|T201|MTH_LN|30522-7|LNC|C-reactive protein|C-reactive protein
C1114363|T201|LC|30522-7|LNC|C-reactive protein|C-reactive protein
C1114363|T201|OSN|30522-7|LNC|C-reactive protein|C-reactive protein
C1114363|T201|LN|30522-7|LNC|protein|protein
C1114363|T201|MTH_LN|30522-7|LNC|protein|protein
C1114363|T201|LC|30522-7|LNC|protein|protein
C1114363|T201|OSN|30522-7|LNC|protein|protein
C1114363|T201|LN|30522-7|LNC|C-peptide|C-peptide
C1114363|T201|MTH_LN|30522-7|LNC|C-peptide|C-peptide
C1114363|T201|LC|30522-7|LNC|C-peptide|C-peptide
C1114363|T201|OSN|30522-7|LNC|C-peptide|C-peptide
C1114363|T201|LN|30522-7|LNC|C peptide|C peptide
C1114363|T201|MTH_LN|30522-7|LNC|C peptide|C peptide
C1114363|T201|LC|30522-7|LNC|C peptide|C peptide
C1114363|T201|OSN|30522-7|LNC|C peptide|C peptide
C1114387|T201|LN|30552-4|LNC|vitamin b6|vitamin b6
C1114387|T201|MTH_LN|30552-4|LNC|vitamin b6|vitamin b6
C1114387|T201|OSN|30552-4|LNC|vitamin b6|vitamin b6
C1114387|T201|LC|30552-4|LNC|vitamin b6|vitamin b6
C1114387|T201|LN|30552-4|LNC|vitamin B metabolism|vitamin B metabolism
C1114387|T201|MTH_LN|30552-4|LNC|vitamin B metabolism|vitamin B metabolism
C1114387|T201|OSN|30552-4|LNC|vitamin B metabolism|vitamin B metabolism
C1114387|T201|LC|30552-4|LNC|vitamin B metabolism|vitamin B metabolism
C1114387|T201|LN|30552-4|LNC|B-vitamin metabolism|B-vitamin metabolism
C1114387|T201|MTH_LN|30552-4|LNC|B-vitamin metabolism|B-vitamin metabolism
C1114387|T201|OSN|30552-4|LNC|B-vitamin metabolism|B-vitamin metabolism
C1114387|T201|LC|30552-4|LNC|B-vitamin metabolism|B-vitamin metabolism
C1114398|T201|LN|30563-1|LNC|taurine|taurine
C1114398|T201|MTH_LN|30563-1|LNC|taurine|taurine
C1114398|T201|OSN|30563-1|LNC|taurine|taurine
C1114398|T201|LC|30563-1|LNC|taurine|taurine
C1114402|T201|LN|30567-2|LNC|thyroid stimulating|thyroid stimulating
C1114402|T201|MTH_LN|30567-2|LNC|thyroid stimulating|thyroid stimulating
C1114402|T201|OSN|30567-2|LNC|thyroid stimulating|thyroid stimulating
C1114402|T201|LC|30567-2|LNC|thyroid stimulating|thyroid stimulating
C1114402|T201|LN|30567-2|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C1114402|T201|MTH_LN|30567-2|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C1114402|T201|OSN|30567-2|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C1114402|T201|LC|30567-2|LNC|Thyroid-stimulating excess|Thyroid-stimulating excess
C1114402|T201|LN|30567-2|LNC|TSH|TSH
C1114402|T201|MTH_LN|30567-2|LNC|TSH|TSH
C1114402|T201|OSN|30567-2|LNC|TSH|TSH
C1114402|T201|LC|30567-2|LNC|TSH|TSH
C1114402|T201|LN|30567-2|LNC|thyroid-stimulating|thyroid-stimulating
C1114402|T201|MTH_LN|30567-2|LNC|thyroid-stimulating|thyroid-stimulating
C1114402|T201|OSN|30567-2|LNC|thyroid-stimulating|thyroid-stimulating
C1114402|T201|LC|30567-2|LNC|thyroid-stimulating|thyroid-stimulating
C1114721|T201|LC|30934-4|LNC|B-type natriuretic peptide|B-type natriuretic peptide
C1114721|T201|MTH_LN|30934-4|LNC|B-type natriuretic peptide|B-type natriuretic peptide
C1114721|T201|LN|30934-4|LNC|B-type natriuretic peptide|B-type natriuretic peptide
C1114721|T201|OSN|30934-4|LNC|B-type natriuretic peptide|B-type natriuretic peptide
C1114721|T201|LC|30934-4|LNC|NT-proBNP|NT-proBNP
C1114721|T201|MTH_LN|30934-4|LNC|NT-proBNP|NT-proBNP
C1114721|T201|LN|30934-4|LNC|NT-proBNP|NT-proBNP
C1114721|T201|OSN|30934-4|LNC|NT-proBNP|NT-proBNP
C1114799|T201|LN|31017-7|LNC|immunoglobulin|immunoglobulin
C1114799|T201|MTH_LN|31017-7|LNC|immunoglobulin|immunoglobulin
C1114799|T201|OSN|31017-7|LNC|immunoglobulin|immunoglobulin
C1114799|T201|LC|31017-7|LNC|immunoglobulin|immunoglobulin
C1114843|T201|LN|29953-7|LNC|Antinuclear antibody|Antinuclear antibody
C1114843|T201|MTH_LN|29953-7|LNC|Antinuclear antibody|Antinuclear antibody
C1114843|T201|OSN|29953-7|LNC|Antinuclear antibody|Antinuclear antibody
C1114843|T201|LC|29953-7|LNC|Antinuclear antibody|Antinuclear antibody
C1114856|T201|LN|30048-3|LNC|lysine|lysine
C1114856|T201|MTH_LN|30048-3|LNC|lysine|lysine
C1114856|T201|OSN|30048-3|LNC|lysine|lysine
C1114856|T201|LC|30048-3|LNC|lysine|lysine
C1114857|T201|LN|30051-7|LNC|homocystine|homocystine
C1114857|T201|OSN|30051-7|LNC|homocystine|homocystine
C1114857|T201|MTH_LN|30051-7|LNC|homocystine|homocystine
C1114857|T201|LC|30051-7|LNC|homocystine|homocystine
C1114881|T201|LN|30264-6|LNC|glucose|glucose
C1114881|T201|MTH_LN|30264-6|LNC|glucose|glucose
C1114881|T201|OSN|30264-6|LNC|glucose|glucose
C1114881|T201|LC|30264-6|LNC|glucose|glucose
C1114882|T201|LN|30266-1|LNC|glucose|glucose
C1114882|T201|MTH_LN|30266-1|LNC|glucose|glucose
C1114882|T201|OSN|30266-1|LNC|glucose|glucose
C1114882|T201|LC|30266-1|LNC|glucose|glucose
C1114891|T201|MTH_LN|30341-2|LNC|erythrocyte|erythrocyte
C1114891|T201|LC|30341-2|LNC|erythrocyte|erythrocyte
C1114891|T201|LN|30341-2|LNC|erythrocyte|erythrocyte
C1114891|T201|OSN|30341-2|LNC|erythrocyte|erythrocyte
C1114891|T201|MTH_LN|30341-2|LNC|ESR|ESR
C1114891|T201|LC|30341-2|LNC|ESR|ESR
C1114891|T201|LN|30341-2|LNC|ESR|ESR
C1114891|T201|OSN|30341-2|LNC|ESR|ESR
// C1114891|T201|MTH_LN|30341-2|LNC||
// C1114891|T201|LC|30341-2|LNC||
// C1114891|T201|LN|30341-2|LNC||
// C1114891|T201|OSN|30341-2|LNC||
C1114891|T201|MTH_LN|30341-2|LNC|Raised erythrocyte|Raised erythrocyte
C1114891|T201|LC|30341-2|LNC|Raised erythrocyte|Raised erythrocyte
C1114891|T201|LN|30341-2|LNC|Raised erythrocyte|Raised erythrocyte
C1114891|T201|OSN|30341-2|LNC|Raised erythrocyte|Raised erythrocyte
C1114891|T201|MTH_LN|30341-2|LNC|Westergren|Westergren
C1114891|T201|LC|30341-2|LNC|Westergren|Westergren
C1114891|T201|LN|30341-2|LNC|Westergren|Westergren
C1114891|T201|OSN|30341-2|LNC|Westergren|Westergren
C1114892|T201|LN|30346-1|LNC|glucose|glucose
C1114892|T201|MTH_LN|30346-1|LNC|glucose|glucose
C1114892|T201|OSN|30346-1|LNC|glucose|glucose
C1114892|T201|LC|30346-1|LNC|glucose|glucose
C1145645|T201|LN|2703-7|LNC|oxygen|oxygen
C1145645|T201|MTH_LN|2703-7|LNC|oxygen|oxygen
C1145645|T201|LC|2703-7|LNC|oxygen|oxygen
C1145645|T201|OSN|2703-7|LNC|oxygen|oxygen
C1145646|T201|LN|2704-5|LNC|oxygen|oxygen
C1145646|T201|MTH_LN|2704-5|LNC|oxygen|oxygen
C1145646|T201|LC|2704-5|LNC|oxygen|oxygen
C1145646|T201|OSN|2704-5|LNC|oxygen|oxygen
C1145647|T201|LN|2705-2|LNC|oxygen|oxygen
C1145647|T201|MTH_LN|2705-2|LNC|oxygen|oxygen
C1145647|T201|LC|2705-2|LNC|oxygen|oxygen
C1145647|T201|OSN|2705-2|LNC|oxygen|oxygen
C1146785|T201|LN|31100-1|LNC|hematocrit|hematocrit
C1146785|T201|MTH_LN|31100-1|LNC|hematocrit|hematocrit
C1146785|T201|LC|31100-1|LNC|hematocrit|hematocrit
C1146785|T201|OSN|31100-1|LNC|hematocrit|hematocrit
C1146797|T201|LN|31112-6|LNC|reticulocytes|reticulocytes
C1146797|T201|MTH_LN|31112-6|LNC|reticulocytes|reticulocytes
C1146797|T201|OSN|31112-6|LNC|reticulocytes|reticulocytes
C1146797|T201|LC|31112-6|LNC|reticulocytes|reticulocytes
C1146797|T201|LN|31112-6|LNC|reticulocyte count|reticulocyte count
C1146797|T201|MTH_LN|31112-6|LNC|reticulocyte count|reticulocyte count
C1146797|T201|OSN|31112-6|LNC|reticulocyte count|reticulocyte count
C1146797|T201|LC|31112-6|LNC|reticulocyte count|reticulocyte count
C1147090|T201|LN|31405-4|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147090|T201|OSN|31405-4|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147090|T201|MTH_LN|31405-4|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147090|T201|LC|31405-4|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147180|T201|LN|31496-3|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147180|T201|OSN|31496-3|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147180|T201|MTH_LN|31496-3|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147180|T201|LC|31496-3|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147181|T201|LN|31497-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147181|T201|MTH_LN|31497-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147181|T201|LC|31497-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147181|T201|OSN|31497-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147182|T201|LN|31498-9|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147182|T201|LC|31498-9|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147182|T201|OSN|31498-9|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147182|T201|MTH_LN|31498-9|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147183|T201|LN|31499-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147183|T201|LC|31499-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147183|T201|OSN|31499-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147183|T201|MTH_LN|31499-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147184|T201|LN|31500-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147184|T201|MTH_LN|31500-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147184|T201|LC|31500-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147184|T201|OSN|31500-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147185|T201|LN|31501-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147185|T201|MTH_LN|31501-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147185|T201|OSN|31501-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147185|T201|LC|31501-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147186|T201|LN|31502-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147186|T201|MTH_LN|31502-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147186|T201|OSN|31502-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147186|T201|LC|31502-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1147707|T201|LN|32023-4|LNC|insulin-like growth factor 1|insulin-like growth factor 1
C1147707|T201|OSN|32023-4|LNC|insulin-like growth factor 1|insulin-like growth factor 1
C1147707|T201|MTH_LN|32023-4|LNC|insulin-like growth factor 1|insulin-like growth factor 1
C1147707|T201|LC|32023-4|LNC|insulin-like growth factor 1|insulin-like growth factor 1
C1147707|T201|LN|32023-4|LNC|IGF1|IGF1
C1147707|T201|OSN|32023-4|LNC|IGF1|IGF1
C1147707|T201|MTH_LN|32023-4|LNC|IGF1|IGF1
C1147707|T201|LC|32023-4|LNC|IGF1|IGF1
C1147816|T201|LN|32132-3|LNC|lactate|lactate
C1147816|T201|MTH_LN|32132-3|LNC|lactate|lactate
C1147816|T201|OSN|32132-3|LNC|lactate|lactate
C1147816|T201|LC|32132-3|LNC|lactate|lactate
C1147817|T201|LN|32133-1|LNC|lactate|lactate
C1147817|T201|MTH_LN|32133-1|LNC|lactate|lactate
C1147817|T201|OSN|32133-1|LNC|lactate|lactate
C1147817|T201|LC|32133-1|LNC|lactate|lactate
C1147851|T201|LN|32167-9|LNC|color|color
C1147851|T201|LC|32167-9|LNC|color|color
C1147851|T201|MTH_LN|32167-9|LNC|color|color
C1147851|T201|OSN|32167-9|LNC|color|color
C1147851|T201|LN|32167-9|LNC|colour|colour
C1147851|T201|LC|32167-9|LNC|colour|colour
C1147851|T201|MTH_LN|32167-9|LNC|colour|colour
C1147851|T201|OSN|32167-9|LNC|colour|colour
C1147899|T201|LN|32215-6|LNC|thyroxine|thyroxine
C1147899|T201|OSN|32215-6|LNC|thyroxine|thyroxine
C1147899|T201|MTH_LN|32215-6|LNC|thyroxine|thyroxine
C1147899|T201|LC|32215-6|LNC|thyroxine|thyroxine
C1147899|T201|LN|32215-6|LNC|T4|T4
C1147899|T201|OSN|32215-6|LNC|T4|T4
C1147899|T201|MTH_LN|32215-6|LNC|T4|T4
C1147899|T201|LC|32215-6|LNC|T4|T4
C1148003|T201|LN|32319-6|LNC|glucose|glucose
C1148003|T201|MTH_LN|32319-6|LNC|glucose|glucose
C1148003|T201|OSN|32319-6|LNC|glucose|glucose
C1148003|T201|LC|32319-6|LNC|glucose|glucose
C1148004|T201|LN|32320-4|LNC|glucose|glucose
C1148004|T201|MTH_LN|32320-4|LNC|glucose|glucose
C1148004|T201|OSN|32320-4|LNC|glucose|glucose
C1148004|T201|LC|32320-4|LNC|glucose|glucose
C1148005|T201|LN|32321-2|LNC|glucose|glucose
C1148005|T201|MTH_LN|32321-2|LNC|glucose|glucose
C1148005|T201|OSN|32321-2|LNC|glucose|glucose
C1148005|T201|LC|32321-2|LNC|glucose|glucose
C1148006|T201|LN|32322-0|LNC|glucose|glucose
C1148006|T201|MTH_LN|32322-0|LNC|glucose|glucose
C1148006|T201|OSN|32322-0|LNC|glucose|glucose
C1148006|T201|LC|32322-0|LNC|glucose|glucose
C1148010|T201|LN|32326-1|LNC|luteinizing|luteinizing
C1148010|T201|MTH_LN|32326-1|LNC|luteinizing|luteinizing
C1148010|T201|OSN|32326-1|LNC|luteinizing|luteinizing
C1148010|T201|LC|32326-1|LNC|luteinizing|luteinizing
C1148010|T201|LN|32326-1|LNC|LH|LH
C1148010|T201|MTH_LN|32326-1|LNC|LH|LH
C1148010|T201|OSN|32326-1|LNC|LH|LH
C1148010|T201|LC|32326-1|LNC|LH|LH
C1148010|T201|LN|32326-1|LNC|luteinising|luteinising
C1148010|T201|MTH_LN|32326-1|LNC|luteinising|luteinising
C1148010|T201|OSN|32326-1|LNC|luteinising|luteinising
C1148010|T201|LC|32326-1|LNC|luteinising|luteinising
C1148011|T201|LN|32327-9|LNC|luteinizing|luteinizing
C1148011|T201|MTH_LN|32327-9|LNC|luteinizing|luteinizing
C1148011|T201|OSN|32327-9|LNC|luteinizing|luteinizing
C1148011|T201|LC|32327-9|LNC|luteinizing|luteinizing
C1148011|T201|LN|32327-9|LNC|LH|LH
C1148011|T201|MTH_LN|32327-9|LNC|LH|LH
C1148011|T201|OSN|32327-9|LNC|LH|LH
C1148011|T201|LC|32327-9|LNC|LH|LH
C1148011|T201|LN|32327-9|LNC|luteinising|luteinising
C1148011|T201|MTH_LN|32327-9|LNC|luteinising|luteinising
C1148011|T201|OSN|32327-9|LNC|luteinising|luteinising
C1148011|T201|LC|32327-9|LNC|luteinising|luteinising
C1148012|T201|LN|32328-7|LNC|luteinizing|luteinizing
C1148012|T201|MTH_LN|32328-7|LNC|luteinizing|luteinizing
C1148012|T201|OSN|32328-7|LNC|luteinizing|luteinizing
C1148012|T201|LC|32328-7|LNC|luteinizing|luteinizing
C1148012|T201|LN|32328-7|LNC|LH|LH
C1148012|T201|MTH_LN|32328-7|LNC|LH|LH
C1148012|T201|OSN|32328-7|LNC|LH|LH
C1148012|T201|LC|32328-7|LNC|LH|LH
C1148012|T201|LN|32328-7|LNC|luteinising|luteinising
C1148012|T201|MTH_LN|32328-7|LNC|luteinising|luteinising
C1148012|T201|OSN|32328-7|LNC|luteinising|luteinising
C1148012|T201|LC|32328-7|LNC|luteinising|luteinising
C1148038|T201|LN|32354-3|LNC|hematocrit|hematocrit
C1148038|T201|MTH_LN|32354-3|LNC|hematocrit|hematocrit
C1148038|T201|LC|32354-3|LNC|hematocrit|hematocrit
C1148038|T201|OSN|32354-3|LNC|hematocrit|hematocrit
C1148043|T201|LN|32359-2|LNC|glucose|glucose
C1148043|T201|MTH_LN|32359-2|LNC|glucose|glucose
C1148043|T201|OSN|32359-2|LNC|glucose|glucose
C1148043|T201|LC|32359-2|LNC|glucose|glucose
C1148230|T201|LN|32546-4|LNC|glucose-6-phosphate dehydrogenase in red|glucose-6-phosphate dehydrogenase in red
C1148230|T201|MTH_LN|32546-4|LNC|glucose-6-phosphate dehydrogenase in red|glucose-6-phosphate dehydrogenase in red
C1148230|T201|OSN|32546-4|LNC|glucose-6-phosphate dehydrogenase in red|glucose-6-phosphate dehydrogenase in red
C1148230|T201|LC|32546-4|LNC|glucose-6-phosphate dehydrogenase in red|glucose-6-phosphate dehydrogenase in red
C1148230|T201|LN|32546-4|LNC|G6PD in red|G6PD in red
C1148230|T201|MTH_LN|32546-4|LNC|G6PD in red|G6PD in red
C1148230|T201|OSN|32546-4|LNC|G6PD in red|G6PD in red
C1148230|T201|LC|32546-4|LNC|G6PD in red|G6PD in red
C1148231|T201|LN|32547-2|LNC|ketone bodies|ketone bodies
C1148231|T201|MTH_LN|32547-2|LNC|ketone bodies|ketone bodies
C1148231|T201|OSN|32547-2|LNC|ketone bodies|ketone bodies
C1148231|T201|LC|32547-2|LNC|ketone bodies|ketone bodies
C1148236|T201|LN|32552-2|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C1148236|T201|MTH_LN|32552-2|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C1148236|T201|OSN|32552-2|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C1148236|T201|LC|32552-2|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C1148236|T201|LN|32552-2|LNC|red cell pyruvate kinase activity|red cell pyruvate kinase activity
C1148236|T201|MTH_LN|32552-2|LNC|red cell pyruvate kinase activity|red cell pyruvate kinase activity
C1148236|T201|OSN|32552-2|LNC|red cell pyruvate kinase activity|red cell pyruvate kinase activity
C1148236|T201|LC|32552-2|LNC|red cell pyruvate kinase activity|red cell pyruvate kinase activity
C1148236|T201|LN|32552-2|LNC|erythrocyte pyruvate kinase activity|erythrocyte pyruvate kinase activity
C1148236|T201|MTH_LN|32552-2|LNC|erythrocyte pyruvate kinase activity|erythrocyte pyruvate kinase activity
C1148236|T201|OSN|32552-2|LNC|erythrocyte pyruvate kinase activity|erythrocyte pyruvate kinase activity
C1148236|T201|LC|32552-2|LNC|erythrocyte pyruvate kinase activity|erythrocyte pyruvate kinase activity
C1148239|T201|LN|32555-5|LNC|urate|urate
C1148239|T201|LC|32555-5|LNC|urate|urate
C1148239|T201|MTH_LN|32555-5|LNC|urate|urate
C1148239|T201|OSN|32555-5|LNC|urate|urate
C1148239|T201|LN|32555-5|LNC|uric acid|uric acid
C1148239|T201|LC|32555-5|LNC|uric acid|uric acid
C1148239|T201|MTH_LN|32555-5|LNC|uric acid|uric acid
C1148239|T201|OSN|32555-5|LNC|uric acid|uric acid
C1148283|T201|LN|32599-3|LNC|luteinizing|luteinizing
C1148283|T201|MTH_LN|32599-3|LNC|luteinizing|luteinizing
C1148283|T201|OSN|32599-3|LNC|luteinizing|luteinizing
C1148283|T201|LC|32599-3|LNC|luteinizing|luteinizing
C1148283|T201|LN|32599-3|LNC|LH|LH
C1148283|T201|MTH_LN|32599-3|LNC|LH|LH
C1148283|T201|OSN|32599-3|LNC|LH|LH
C1148283|T201|LC|32599-3|LNC|LH|LH
C1148283|T201|LN|32599-3|LNC|luteinising|luteinising
C1148283|T201|MTH_LN|32599-3|LNC|luteinising|luteinising
C1148283|T201|OSN|32599-3|LNC|luteinising|luteinising
C1148283|T201|LC|32599-3|LNC|luteinising|luteinising
C1148290|T201|LN|32606-6|LNC|luteinizing|luteinizing
C1148290|T201|MTH_LN|32606-6|LNC|luteinizing|luteinizing
C1148290|T201|OSN|32606-6|LNC|luteinizing|luteinizing
C1148290|T201|LC|32606-6|LNC|luteinizing|luteinizing
C1148290|T201|LN|32606-6|LNC|LH|LH
C1148290|T201|MTH_LN|32606-6|LNC|LH|LH
C1148290|T201|OSN|32606-6|LNC|LH|LH
C1148290|T201|LC|32606-6|LNC|LH|LH
C1148290|T201|LN|32606-6|LNC|luteinising|luteinising
C1148290|T201|MTH_LN|32606-6|LNC|luteinising|luteinising
C1148290|T201|OSN|32606-6|LNC|luteinising|luteinising
C1148290|T201|LC|32606-6|LNC|luteinising|luteinising
C1153749|T201|LN|19214-6|LNC|oxygen|oxygen
C1153749|T201|MTH_LN|19214-6|LNC|oxygen|oxygen
C1153749|T201|OSN|19214-6|LNC|oxygen|oxygen
C1153749|T201|LC|19214-6|LNC|oxygen|oxygen
C1171343|T098|LN|2157-6|LNC|creatine phosphokinase|creatine phosphokinase
C1171343|T098|MTH_LN|2157-6|LNC|creatine phosphokinase|creatine phosphokinase
C1171343|T098|OSN|2157-6|LNC|creatine phosphokinase|creatine phosphokinase
C1171343|T098|LC|2157-6|LNC|creatine phosphokinase|creatine phosphokinase
C1171343|T098|LN|2157-6|LNC|CPK|CPK
C1171343|T098|MTH_LN|2157-6|LNC|CPK|CPK
C1171343|T098|OSN|2157-6|LNC|CPK|CPK
C1171343|T098|LC|2157-6|LNC|CPK|CPK
C1171343|T098|LN|2157-6|LNC|creatine kinase|creatine kinase
C1171343|T098|MTH_LN|2157-6|LNC|creatine kinase|creatine kinase
C1171343|T098|OSN|2157-6|LNC|creatine kinase|creatine kinase
C1171343|T098|LC|2157-6|LNC|creatine kinase|creatine kinase
C1171343|T098|LN|2157-6|LNC|CK|CK
C1171343|T098|MTH_LN|2157-6|LNC|CK|CK
C1171343|T098|OSN|2157-6|LNC|CK|CK
C1171343|T098|LC|2157-6|LNC|CK|CK
C1171359|T098|LC|2160-0|LNC|creatinine|creatinine
C1171359|T098|LN|2160-0|LNC|creatinine|creatinine
C1171359|T098|MTH_LN|2160-0|LNC|creatinine|creatinine
C1171359|T098|OSN|2160-0|LNC|creatinine|creatinine
C1171364|T098|LN|2161-8|LNC|creatinine|creatinine
C1171364|T098|MTH_LN|2161-8|LNC|creatinine|creatinine
C1171364|T098|OSN|2161-8|LNC|creatinine|creatinine
C1171364|T098|LC|2161-8|LNC|creatinine|creatinine
C1171364|T098|LN|2161-8|LNC|metabolism/homeostasis|metabolism/homeostasis
C1171364|T098|MTH_LN|2161-8|LNC|metabolism/homeostasis|metabolism/homeostasis
C1171364|T098|OSN|2161-8|LNC|metabolism/homeostasis|metabolism/homeostasis
C1171364|T098|LC|2161-8|LNC|metabolism/homeostasis|metabolism/homeostasis
C1171364|T098|LN|2161-8|LNC|Metabolism|Metabolism
C1171364|T098|MTH_LN|2161-8|LNC|Metabolism|Metabolism
C1171364|T098|OSN|2161-8|LNC|Metabolism|Metabolism
C1171364|T098|LC|2161-8|LNC|Metabolism|Metabolism
C1171364|T098|LN|2161-8|LNC|Laboratory|Laboratory
C1171364|T098|MTH_LN|2161-8|LNC|Laboratory|Laboratory
C1171364|T098|OSN|2161-8|LNC|Laboratory|Laboratory
C1171364|T098|LC|2161-8|LNC|Laboratory|Laboratory
C1315089|T201|LN|32615-7|LNC|homocystine|homocystine
C1315089|T201|MTH_LN|32615-7|LNC|homocystine|homocystine
C1315089|T201|OSN|32615-7|LNC|homocystine|homocystine
C1315089|T201|LC|32615-7|LNC|homocystine|homocystine
C1315089|T201|LN|32615-7|LNC|homocysteine metabolism|homocysteine metabolism
C1315089|T201|MTH_LN|32615-7|LNC|homocysteine metabolism|homocysteine metabolism
C1315089|T201|OSN|32615-7|LNC|homocysteine metabolism|homocysteine metabolism
C1315089|T201|LC|32615-7|LNC|homocysteine metabolism|homocysteine metabolism
C1315138|T201|LN|32664-5|LNC|ammonia|ammonia
C1315138|T201|OSN|32664-5|LNC|ammonia|ammonia
C1315138|T201|MTH_LN|32664-5|LNC|ammonia|ammonia
C1315138|T201|LC|32664-5|LNC|ammonia|ammonia
C1315156|T201|LN|32682-7|LNC|hemoglobin F|hemoglobin F
C1315156|T201|MTH_LN|32682-7|LNC|hemoglobin F|hemoglobin F
C1315156|T201|LC|32682-7|LNC|hemoglobin F|hemoglobin F
C1315156|T201|OSN|32682-7|LNC|hemoglobin F|hemoglobin F
C1315156|T201|LN|32682-7|LNC|hemoglobin|hemoglobin
C1315156|T201|MTH_LN|32682-7|LNC|hemoglobin|hemoglobin
C1315156|T201|LC|32682-7|LNC|hemoglobin|hemoglobin
C1315156|T201|OSN|32682-7|LNC|hemoglobin|hemoglobin
C1315157|T201|LN|32683-5|LNC|alpha-fetoprotein|alpha-fetoprotein
C1315157|T201|MTH_LN|32683-5|LNC|alpha-fetoprotein|alpha-fetoprotein
C1315157|T201|LC|32683-5|LNC|alpha-fetoprotein|alpha-fetoprotein
C1315157|T201|OSN|32683-5|LNC|alpha-fetoprotein|alpha-fetoprotein
C1315166|T201|LN|32693-4|LNC|lactate|lactate
C1315166|T201|OSN|32693-4|LNC|lactate|lactate
C1315166|T201|MTH_LN|32693-4|LNC|lactate|lactate
C1315166|T201|LC|32693-4|LNC|lactate|lactate
C1315182|T201|MTH_LN|32623-1|LNC|mean platelet volume|mean platelet volume
C1315182|T201|LN|32623-1|LNC|mean platelet volume|mean platelet volume
C1315182|T201|LC|32623-1|LNC|mean platelet volume|mean platelet volume
C1315182|T201|OSN|32623-1|LNC|mean platelet volume|mean platelet volume
C1315182|T201|MTH_LN|32623-1|LNC|platelet volume|platelet volume
C1315182|T201|LN|32623-1|LNC|platelet volume|platelet volume
C1315182|T201|LC|32623-1|LNC|platelet volume|platelet volume
C1315182|T201|OSN|32623-1|LNC|platelet volume|platelet volume
C1315188|T201|LN|32717-1|LNC|sodium|sodium
C1315188|T201|MTH_LN|32717-1|LNC|sodium|sodium
C1315188|T201|OSN|32717-1|LNC|sodium|sodium
C1315188|T201|LC|32717-1|LNC|sodium|sodium
C1315188|T201|LN|32717-1|LNC|sodium homeostasis|sodium homeostasis
C1315188|T201|MTH_LN|32717-1|LNC|sodium homeostasis|sodium homeostasis
C1315188|T201|OSN|32717-1|LNC|sodium homeostasis|sodium homeostasis
C1315188|T201|LC|32717-1|LNC|sodium homeostasis|sodium homeostasis
C1315198|T201|LN|32727-0|LNC|urobilinogen|urobilinogen
C1315198|T201|OSN|32727-0|LNC|urobilinogen|urobilinogen
C1315198|T201|MTH_LN|32727-0|LNC|urobilinogen|urobilinogen
C1315198|T201|LC|32727-0|LNC|urobilinogen|urobilinogen
C1315242|T201|LN|32771-8|LNC|carbon dioxide|carbon dioxide
C1315242|T201|MTH_LN|32771-8|LNC|carbon dioxide|carbon dioxide
C1315242|T201|LC|32771-8|LNC|carbon dioxide|carbon dioxide
C1315242|T201|OSN|32771-8|LNC|carbon dioxide|carbon dioxide
C1315291|T201|LN|32820-3|LNC|glucose|glucose
C1315291|T201|MTH_LN|32820-3|LNC|glucose|glucose
C1315291|T201|OSN|32820-3|LNC|glucose|glucose
C1315291|T201|LC|32820-3|LNC|glucose|glucose
C1315325|T201|LN|32854-2|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C1315325|T201|MTH_LN|32854-2|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C1315325|T201|LC|32854-2|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C1315325|T201|OSN|32854-2|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C1315325|T201|LN|32854-2|LNC|17-OHP|17-OHP
C1315325|T201|MTH_LN|32854-2|LNC|17-OHP|17-OHP
C1315325|T201|LC|32854-2|LNC|17-OHP|17-OHP
C1315325|T201|OSN|32854-2|LNC|17-OHP|17-OHP
C1315466|T201|LN|32995-3|LNC|luteinizing|luteinizing
C1315466|T201|MTH_LN|32995-3|LNC|luteinizing|luteinizing
C1315466|T201|OSN|32995-3|LNC|luteinizing|luteinizing
C1315466|T201|LC|32995-3|LNC|luteinizing|luteinizing
C1315466|T201|LN|32995-3|LNC|LH|LH
C1315466|T201|MTH_LN|32995-3|LNC|LH|LH
C1315466|T201|OSN|32995-3|LNC|LH|LH
C1315466|T201|LC|32995-3|LNC|LH|LH
C1315466|T201|LN|32995-3|LNC|luteinising|luteinising
C1315466|T201|MTH_LN|32995-3|LNC|luteinising|luteinising
C1315466|T201|OSN|32995-3|LNC|luteinising|luteinising
C1315466|T201|LC|32995-3|LNC|luteinising|luteinising
C1315469|T201|LN|32998-7|LNC|immunoglobulin|immunoglobulin
C1315469|T201|OSN|32998-7|LNC|immunoglobulin|immunoglobulin
C1315469|T201|MTH_LN|32998-7|LNC|immunoglobulin|immunoglobulin
C1315469|T201|LC|32998-7|LNC|immunoglobulin|immunoglobulin
C1315495|T201|LN|33024-1|LNC|glucose|glucose
C1315495|T201|MTH_LN|33024-1|LNC|glucose|glucose
C1315495|T201|OSN|33024-1|LNC|glucose|glucose
C1315495|T201|LC|33024-1|LNC|glucose|glucose
// C1315522|T201|LN|33051-4|LNC||
// C1315522|T201|MTH_LN|33051-4|LNC||
// C1315522|T201|OSN|33051-4|LNC||
// C1315522|T201|LC|33051-4|LNC||
C1315522|T201|LN|33051-4|LNC|occult|occult
C1315522|T201|MTH_LN|33051-4|LNC|occult|occult
C1315522|T201|OSN|33051-4|LNC|occult|occult
C1315522|T201|LC|33051-4|LNC|occult|occult
C1315523|T201|LN|33052-2|LNC|neutrophil count|neutrophil count
C1315523|T201|MTH_LN|33052-2|LNC|neutrophil count|neutrophil count
C1315523|T201|OSN|33052-2|LNC|neutrophil count|neutrophil count
C1315523|T201|LC|33052-2|LNC|neutrophil count|neutrophil count
C1315523|T201|LN|33052-2|LNC|cytology|cytology
C1315523|T201|MTH_LN|33052-2|LNC|cytology|cytology
C1315523|T201|OSN|33052-2|LNC|cytology|cytology
C1315523|T201|LC|33052-2|LNC|cytology|cytology
C1315529|T201|LN|33058-9|LNC|ketone bodies|ketone bodies
C1315529|T201|MTH_LN|33058-9|LNC|ketone bodies|ketone bodies
C1315529|T201|OSN|33058-9|LNC|ketone bodies|ketone bodies
C1315529|T201|LC|33058-9|LNC|ketone bodies|ketone bodies
C1315540|T201|LN|33069-6|LNC|nuchal translucency|nuchal translucency
C1315540|T201|MTH_LN|33069-6|LNC|nuchal translucency|nuchal translucency
C1315540|T201|LC|33069-6|LNC|nuchal translucency|nuchal translucency
C1315540|T201|OSN|33069-6|LNC|nuchal translucency|nuchal translucency
C1315675|T201|LN|33204-9|LNC|troponin T|troponin T
C1315675|T201|MTH_LN|33204-9|LNC|troponin T|troponin T
C1315675|T201|OSN|33204-9|LNC|troponin T|troponin T
C1315675|T201|LC|33204-9|LNC|troponin T|troponin T
C1315725|T201|LN|33256-9|LNC|white count|white count
C1315725|T201|OSN|33256-9|LNC|white count|white count
C1315725|T201|MTH_LN|33256-9|LNC|white count|white count
C1315725|T201|LC|33256-9|LNC|white count|white count
C1315725|T201|LN|33256-9|LNC|leukocyte number|leukocyte number
C1315725|T201|OSN|33256-9|LNC|leukocyte number|leukocyte number
C1315725|T201|MTH_LN|33256-9|LNC|leukocyte number|leukocyte number
C1315725|T201|LC|33256-9|LNC|leukocyte number|leukocyte number
C1315725|T201|LN|33256-9|LNC|white cell count|white cell count
C1315725|T201|OSN|33256-9|LNC|white cell count|white cell count
C1315725|T201|MTH_LN|33256-9|LNC|white cell count|white cell count
C1315725|T201|LC|33256-9|LNC|white cell count|white cell count
C1315725|T201|LN|33256-9|LNC|leukocyte count|leukocyte count
C1315725|T201|OSN|33256-9|LNC|leukocyte count|leukocyte count
C1315725|T201|MTH_LN|33256-9|LNC|leukocyte count|leukocyte count
C1315725|T201|LC|33256-9|LNC|leukocyte count|leukocyte count
C1315743|T201|LN|33274-2|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1315743|T201|MTH_LN|33274-2|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1315743|T201|OSN|33274-2|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1315743|T201|LC|33274-2|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1315743|T201|LN|33274-2|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1315743|T201|MTH_LN|33274-2|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1315743|T201|OSN|33274-2|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1315743|T201|LC|33274-2|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1315743|T201|LN|33274-2|LNC|folate metabolism|folate metabolism
C1315743|T201|MTH_LN|33274-2|LNC|folate metabolism|folate metabolism
C1315743|T201|OSN|33274-2|LNC|folate metabolism|folate metabolism
C1315743|T201|LC|33274-2|LNC|folate metabolism|folate metabolism
C1315744|T201|LN|33275-9|LNC|7-dehydrocholesterol|7-dehydrocholesterol
C1315744|T201|OSN|33275-9|LNC|7-dehydrocholesterol|7-dehydrocholesterol
C1315744|T201|MTH_LN|33275-9|LNC|7-dehydrocholesterol|7-dehydrocholesterol
C1315744|T201|LC|33275-9|LNC|7-dehydrocholesterol|7-dehydrocholesterol
C1315744|T201|LN|33275-9|LNC|cholesta-5,7-dien-3beta-ol|cholesta-5,7-dien-3beta-ol
C1315744|T201|OSN|33275-9|LNC|cholesta-5,7-dien-3beta-ol|cholesta-5,7-dien-3beta-ol
C1315744|T201|MTH_LN|33275-9|LNC|cholesta-5,7-dien-3beta-ol|cholesta-5,7-dien-3beta-ol
C1315744|T201|LC|33275-9|LNC|cholesta-5,7-dien-3beta-ol|cholesta-5,7-dien-3beta-ol
C1315747|T201|LN|33278-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1315747|T201|OSN|33278-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1315747|T201|MTH_LN|33278-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1315747|T201|LC|33278-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1315748|T201|LN|33279-1|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1315748|T201|OSN|33279-1|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1315748|T201|MTH_LN|33279-1|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1315748|T201|LC|33279-1|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1315756|T201|LN|33287-4|LNC|glucose-6-phosphate dehydrogenase in dried spot|glucose-6-phosphate dehydrogenase in dried spot
C1315756|T201|MTH_LN|33287-4|LNC|glucose-6-phosphate dehydrogenase in dried spot|glucose-6-phosphate dehydrogenase in dried spot
C1315756|T201|LC|33287-4|LNC|glucose-6-phosphate dehydrogenase in dried spot|glucose-6-phosphate dehydrogenase in dried spot
C1315756|T201|OSN|33287-4|LNC|glucose-6-phosphate dehydrogenase in dried spot|glucose-6-phosphate dehydrogenase in dried spot
C1315756|T201|LN|33287-4|LNC|glucose-6-phosphate dehydrogenase in DBS|glucose-6-phosphate dehydrogenase in DBS
C1315756|T201|MTH_LN|33287-4|LNC|glucose-6-phosphate dehydrogenase in DBS|glucose-6-phosphate dehydrogenase in DBS
C1315756|T201|LC|33287-4|LNC|glucose-6-phosphate dehydrogenase in DBS|glucose-6-phosphate dehydrogenase in DBS
C1315756|T201|OSN|33287-4|LNC|glucose-6-phosphate dehydrogenase in DBS|glucose-6-phosphate dehydrogenase in DBS
C1315756|T201|LN|33287-4|LNC|G6PD in dried spot|G6PD in dried spot
C1315756|T201|MTH_LN|33287-4|LNC|G6PD in dried spot|G6PD in dried spot
C1315756|T201|LC|33287-4|LNC|G6PD in dried spot|G6PD in dried spot
C1315756|T201|OSN|33287-4|LNC|G6PD in dried spot|G6PD in dried spot
C1315880|T201|LN|33411-0|LNC|Hemoglobin|Hemoglobin
C1315880|T201|MTH_LN|33411-0|LNC|Hemoglobin|Hemoglobin
C1315880|T201|OSN|33411-0|LNC|Hemoglobin|Hemoglobin
C1315880|T201|LC|33411-0|LNC|Hemoglobin|Hemoglobin
C1315996|T201|LN|33527-3|LNC|methadone test|methadone test
C1315996|T201|MTH_LN|33527-3|LNC|methadone test|methadone test
C1315996|T201|OSN|33527-3|LNC|methadone test|methadone test
C1315996|T201|LC|33527-3|LNC|methadone test|methadone test
C1316226|T201|LN|33762-6|LNC|B-type natriuretic peptide|B-type natriuretic peptide
C1316226|T201|OSN|33762-6|LNC|B-type natriuretic peptide|B-type natriuretic peptide
C1316226|T201|MTH_LN|33762-6|LNC|B-type natriuretic peptide|B-type natriuretic peptide
C1316226|T201|LC|33762-6|LNC|B-type natriuretic peptide|B-type natriuretic peptide
C1316226|T201|LN|33762-6|LNC|NT-proBNP|NT-proBNP
C1316226|T201|OSN|33762-6|LNC|NT-proBNP|NT-proBNP
C1316226|T201|MTH_LN|33762-6|LNC|NT-proBNP|NT-proBNP
C1316226|T201|LC|33762-6|LNC|NT-proBNP|NT-proBNP
C1316260|T201|LN|33796-4|LNC|cotinine|cotinine
C1316260|T201|MTH_LN|33796-4|LNC|cotinine|cotinine
C1316260|T201|OSN|33796-4|LNC|cotinine|cotinine
C1316260|T201|LC|33796-4|LNC|cotinine|cotinine
C1316290|T201|LN|33826-9|LNC|luteinizing|luteinizing
C1316290|T201|MTH_LN|33826-9|LNC|luteinizing|luteinizing
C1316290|T201|OSN|33826-9|LNC|luteinizing|luteinizing
C1316290|T201|LC|33826-9|LNC|luteinizing|luteinizing
C1316290|T201|LN|33826-9|LNC|LH|LH
C1316290|T201|MTH_LN|33826-9|LNC|LH|LH
C1316290|T201|OSN|33826-9|LNC|LH|LH
C1316290|T201|LC|33826-9|LNC|LH|LH
C1316290|T201|LN|33826-9|LNC|luteinising|luteinising
C1316290|T201|MTH_LN|33826-9|LNC|luteinising|luteinising
C1316290|T201|OSN|33826-9|LNC|luteinising|luteinising
C1316290|T201|LC|33826-9|LNC|luteinising|luteinising
C1316291|T201|LN|33827-7|LNC|luteinizing|luteinizing
C1316291|T201|MTH_LN|33827-7|LNC|luteinizing|luteinizing
C1316291|T201|OSN|33827-7|LNC|luteinizing|luteinizing
C1316291|T201|LC|33827-7|LNC|luteinizing|luteinizing
C1316291|T201|LN|33827-7|LNC|LH|LH
C1316291|T201|MTH_LN|33827-7|LNC|LH|LH
C1316291|T201|OSN|33827-7|LNC|LH|LH
C1316291|T201|LC|33827-7|LNC|LH|LH
C1316291|T201|LN|33827-7|LNC|luteinising|luteinising
C1316291|T201|MTH_LN|33827-7|LNC|luteinising|luteinising
C1316291|T201|OSN|33827-7|LNC|luteinising|luteinising
C1316291|T201|LC|33827-7|LNC|luteinising|luteinising
C1316292|T201|LN|33828-5|LNC|luteinizing|luteinizing
C1316292|T201|MTH_LN|33828-5|LNC|luteinizing|luteinizing
C1316292|T201|OSN|33828-5|LNC|luteinizing|luteinizing
C1316292|T201|LC|33828-5|LNC|luteinizing|luteinizing
C1316292|T201|LN|33828-5|LNC|LH|LH
C1316292|T201|MTH_LN|33828-5|LNC|LH|LH
C1316292|T201|OSN|33828-5|LNC|LH|LH
C1316292|T201|LC|33828-5|LNC|LH|LH
C1316292|T201|LN|33828-5|LNC|luteinising|luteinising
C1316292|T201|MTH_LN|33828-5|LNC|luteinising|luteinising
C1316292|T201|OSN|33828-5|LNC|luteinising|luteinising
C1316292|T201|LC|33828-5|LNC|luteinising|luteinising
C1316293|T201|LN|33829-3|LNC|luteinizing|luteinizing
C1316293|T201|MTH_LN|33829-3|LNC|luteinizing|luteinizing
C1316293|T201|OSN|33829-3|LNC|luteinizing|luteinizing
C1316293|T201|LC|33829-3|LNC|luteinizing|luteinizing
C1316293|T201|LN|33829-3|LNC|LH|LH
C1316293|T201|MTH_LN|33829-3|LNC|LH|LH
C1316293|T201|OSN|33829-3|LNC|LH|LH
C1316293|T201|LC|33829-3|LNC|LH|LH
C1316293|T201|LN|33829-3|LNC|luteinising|luteinising
C1316293|T201|MTH_LN|33829-3|LNC|luteinising|luteinising
C1316293|T201|OSN|33829-3|LNC|luteinising|luteinising
C1316293|T201|LC|33829-3|LNC|luteinising|luteinising
C1316361|T201|LN|33898-8|LNC|bilirubin|bilirubin
C1316361|T201|OSN|33898-8|LNC|bilirubin|bilirubin
C1316361|T201|MTH_LN|33898-8|LNC|bilirubin|bilirubin
C1316361|T201|LC|33898-8|LNC|bilirubin|bilirubin
C1316361|T201|LN|33898-8|LNC|total bilirubin|total bilirubin
C1316361|T201|OSN|33898-8|LNC|total bilirubin|total bilirubin
C1316361|T201|MTH_LN|33898-8|LNC|total bilirubin|total bilirubin
C1316361|T201|LC|33898-8|LNC|total bilirubin|total bilirubin
C1316361|T201|LN|33898-8|LNC|bili total|bili total
C1316361|T201|OSN|33898-8|LNC|bili total|bili total
C1316361|T201|MTH_LN|33898-8|LNC|bili total|bili total
C1316361|T201|LC|33898-8|LNC|bili total|bili total
C1316377|T201|LN|33914-3|LNC|glomerular filtration rate|glomerular filtration rate
C1316377|T201|MTH_LN|33914-3|LNC|glomerular filtration rate|glomerular filtration rate
C1316377|T201|LC|33914-3|LNC|glomerular filtration rate|glomerular filtration rate
C1316377|T201|OSN|33914-3|LNC|glomerular filtration rate|glomerular filtration rate
C1316377|T201|LN|33914-3|LNC|creatinine clearance|creatinine clearance
C1316377|T201|MTH_LN|33914-3|LNC|creatinine clearance|creatinine clearance
C1316377|T201|LC|33914-3|LNC|creatinine clearance|creatinine clearance
C1316377|T201|OSN|33914-3|LNC|creatinine clearance|creatinine clearance
C1316518|T201|LN|34055-4|LNC|luteinizing|luteinizing
C1316518|T201|MTH_LN|34055-4|LNC|luteinizing|luteinizing
C1316518|T201|LC|34055-4|LNC|luteinizing|luteinizing
C1316518|T201|OSN|34055-4|LNC|luteinizing|luteinizing
C1316518|T201|LN|34055-4|LNC|LH|LH
C1316518|T201|MTH_LN|34055-4|LNC|LH|LH
C1316518|T201|LC|34055-4|LNC|LH|LH
C1316518|T201|OSN|34055-4|LNC|LH|LH
C1316518|T201|LN|34055-4|LNC|luteinising|luteinising
C1316518|T201|MTH_LN|34055-4|LNC|luteinising|luteinising
C1316518|T201|LC|34055-4|LNC|luteinising|luteinising
C1316518|T201|OSN|34055-4|LNC|luteinising|luteinising
C1316528|T201|LN|34065-3|LNC|cortisol|cortisol
C1316528|T201|MTH_LN|34065-3|LNC|cortisol|cortisol
C1316528|T201|LC|34065-3|LNC|cortisol|cortisol
C1316528|T201|OSN|34065-3|LNC|cortisol|cortisol
C1316528|T201|LN|34065-3|LNC|cortisol low|cortisol low
C1316528|T201|MTH_LN|34065-3|LNC|cortisol low|cortisol low
C1316528|T201|LC|34065-3|LNC|cortisol low|cortisol low
C1316528|T201|OSN|34065-3|LNC|cortisol low|cortisol low
C1316528|T201|LN|34065-3|LNC|to undetectable cortisol|to undetectable cortisol
C1316528|T201|MTH_LN|34065-3|LNC|to undetectable cortisol|to undetectable cortisol
C1316528|T201|LC|34065-3|LNC|to undetectable cortisol|to undetectable cortisol
C1316528|T201|OSN|34065-3|LNC|to undetectable cortisol|to undetectable cortisol
C1316637|T201|LN|34174-3|LNC|Hemoglobin|Hemoglobin
C1316637|T201|MTH_LN|34174-3|LNC|Hemoglobin|Hemoglobin
C1316637|T201|OSN|34174-3|LNC|Hemoglobin|Hemoglobin
C1316637|T201|LC|34174-3|LNC|Hemoglobin|Hemoglobin
C1316747|T201|LN|34284-0|LNC|delta-aminolevulinic acid|delta-aminolevulinic acid
C1316747|T201|OSN|34284-0|LNC|delta-aminolevulinic acid|delta-aminolevulinic acid
C1316747|T201|MTH_LN|34284-0|LNC|delta-aminolevulinic acid|delta-aminolevulinic acid
C1316747|T201|LC|34284-0|LNC|delta-aminolevulinic acid|delta-aminolevulinic acid
C1316773|T201|LN|34310-3|LNC|galactose|galactose
C1316773|T201|MTH_LN|34310-3|LNC|galactose|galactose
C1316773|T201|OSN|34310-3|LNC|galactose|galactose
C1316773|T201|LC|34310-3|LNC|galactose|galactose
C1316774|T201|LN|34311-1|LNC|galactose|galactose
C1316774|T201|MTH_LN|34311-1|LNC|galactose|galactose
C1316774|T201|OSN|34311-1|LNC|galactose|galactose
C1316774|T201|LC|34311-1|LNC|galactose|galactose
C1316828|T201|LN|34366-5|LNC|Protein|Protein
C1316828|T201|LC|34366-5|LNC|Protein|Protein
C1316828|T201|OSN|34366-5|LNC|Protein|Protein
C1316828|T201|MTH_LN|34366-5|LNC|Protein|Protein
C1316847|T201|LN|34385-5|LNC|urate|urate
C1316847|T201|OSN|34385-5|LNC|urate|urate
C1316847|T201|LC|34385-5|LNC|urate|urate
C1316847|T201|MTH_LN|34385-5|LNC|urate|urate
C1316847|T201|LN|34385-5|LNC|uric acid|uric acid
C1316847|T201|OSN|34385-5|LNC|uric acid|uric acid
C1316847|T201|LC|34385-5|LNC|uric acid|uric acid
C1316847|T201|MTH_LN|34385-5|LNC|uric acid|uric acid
C1316896|T201|LN|34434-1|LNC|luteinizing|luteinizing
C1316896|T201|MTH_LN|34434-1|LNC|luteinizing|luteinizing
C1316896|T201|OSN|34434-1|LNC|luteinizing|luteinizing
C1316896|T201|LC|34434-1|LNC|luteinizing|luteinizing
C1316896|T201|LN|34434-1|LNC|LH|LH
C1316896|T201|MTH_LN|34434-1|LNC|LH|LH
C1316896|T201|OSN|34434-1|LNC|LH|LH
C1316896|T201|LC|34434-1|LNC|LH|LH
C1316896|T201|LN|34434-1|LNC|luteinising|luteinising
C1316896|T201|MTH_LN|34434-1|LNC|luteinising|luteinising
C1316896|T201|OSN|34434-1|LNC|luteinising|luteinising
C1316896|T201|LC|34434-1|LNC|luteinising|luteinising
C1316938|T201|LN|34476-2|LNC|cortisol|cortisol
C1316938|T201|MTH_LN|34476-2|LNC|cortisol|cortisol
C1316938|T201|OSN|34476-2|LNC|cortisol|cortisol
C1316938|T201|LC|34476-2|LNC|cortisol|cortisol
C1316938|T201|LN|34476-2|LNC|cortisol low|cortisol low
C1316938|T201|MTH_LN|34476-2|LNC|cortisol low|cortisol low
C1316938|T201|OSN|34476-2|LNC|cortisol low|cortisol low
C1316938|T201|LC|34476-2|LNC|cortisol low|cortisol low
C1316938|T201|LN|34476-2|LNC|to undetectable cortisol|to undetectable cortisol
C1316938|T201|MTH_LN|34476-2|LNC|to undetectable cortisol|to undetectable cortisol
C1316938|T201|OSN|34476-2|LNC|to undetectable cortisol|to undetectable cortisol
C1316938|T201|LC|34476-2|LNC|to undetectable cortisol|to undetectable cortisol
C1328872|T098|LN|2069-3|LNC|chloride|chloride
C1328872|T098|MTH_LN|2069-3|LNC|chloride|chloride
C1328872|T098|OSN|2069-3|LNC|chloride|chloride
C1328872|T098|LC|2069-3|LNC|chloride|chloride
C1328872|T098|LN|2069-3|LNC|chloride homeostasis|chloride homeostasis
C1328872|T098|MTH_LN|2069-3|LNC|chloride homeostasis|chloride homeostasis
C1328872|T098|OSN|2069-3|LNC|chloride homeostasis|chloride homeostasis
C1328872|T098|LC|2069-3|LNC|chloride homeostasis|chloride homeostasis
C1369505|T201|LN|34637-9|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1369505|T201|MTH_LN|34637-9|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1369505|T201|OSN|34637-9|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1369505|T201|LC|34637-9|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1369505|T201|LN|34637-9|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1369505|T201|MTH_LN|34637-9|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1369505|T201|OSN|34637-9|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1369505|T201|LC|34637-9|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1369505|T201|LN|34637-9|LNC|folate metabolism|folate metabolism
C1369505|T201|MTH_LN|34637-9|LNC|folate metabolism|folate metabolism
C1369505|T201|OSN|34637-9|LNC|folate metabolism|folate metabolism
C1369505|T201|LC|34637-9|LNC|folate metabolism|folate metabolism
C1369580|T201|LN|34714-6|LNC|platelet aggregation|platelet aggregation
C1369580|T201|MTH_LN|34714-6|LNC|platelet aggregation|platelet aggregation
C1369580|T201|LC|34714-6|LNC|platelet aggregation|platelet aggregation
C1369580|T201|OSN|34714-6|LNC|platelet aggregation|platelet aggregation
C1369580|T201|LN|34714-6|LNC|RIPA|RIPA
C1369580|T201|MTH_LN|34714-6|LNC|RIPA|RIPA
C1369580|T201|LC|34714-6|LNC|RIPA|RIPA
C1369580|T201|OSN|34714-6|LNC|RIPA|RIPA
C1369594|T201|LN|34728-6|LNC|carbon dioxide|carbon dioxide
C1369594|T201|OSN|34728-6|LNC|carbon dioxide|carbon dioxide
C1369594|T201|MTH_LN|34728-6|LNC|carbon dioxide|carbon dioxide
C1369594|T201|LC|34728-6|LNC|carbon dioxide|carbon dioxide
C1369792|T201|LN|34927-4|LNC|urobilinogen|urobilinogen
C1369792|T201|MTH_LN|34927-4|LNC|urobilinogen|urobilinogen
C1369792|T201|OSN|34927-4|LNC|urobilinogen|urobilinogen
C1369792|T201|LC|34927-4|LNC|urobilinogen|urobilinogen
C1369793|T201|LN|34928-2|LNC|urobilinogen|urobilinogen
C1369793|T201|MTH_LN|34928-2|LNC|urobilinogen|urobilinogen
C1369793|T201|OSN|34928-2|LNC|urobilinogen|urobilinogen
C1369793|T201|LC|34928-2|LNC|urobilinogen|urobilinogen
C1369797|T201|LN|34932-4|LNC|naive T|naive T
C1369797|T201|MTH_LN|34932-4|LNC|naive T|naive T
C1369797|T201|LC|34932-4|LNC|naive T|naive T
C1369797|T201|OSN|34932-4|LNC|naive T|naive T
C1369797|T201|LN|34932-4|LNC|naive T cell|naive T cell
C1369797|T201|MTH_LN|34932-4|LNC|naive T cell|naive T cell
C1369797|T201|LC|34932-4|LNC|naive T cell|naive T cell
C1369797|T201|OSN|34932-4|LNC|naive T cell|naive T cell
C1369798|T201|LN|34933-2|LNC|naive T|naive T
C1369798|T201|MTH_LN|34933-2|LNC|naive T|naive T
C1369798|T201|LC|34933-2|LNC|naive T|naive T
C1369798|T201|OSN|34933-2|LNC|naive T|naive T
C1369798|T201|LN|34933-2|LNC|naive T cell|naive T cell
C1369798|T201|MTH_LN|34933-2|LNC|naive T cell|naive T cell
C1369798|T201|LC|34933-2|LNC|naive T cell|naive T cell
C1369798|T201|OSN|34933-2|LNC|naive T cell|naive T cell
C1369801|T201|LN|34936-5|LNC|naive T|naive T
C1369801|T201|MTH_LN|34936-5|LNC|naive T|naive T
C1369801|T201|LC|34936-5|LNC|naive T|naive T
C1369801|T201|OSN|34936-5|LNC|naive T|naive T
C1369801|T201|LN|34936-5|LNC|naive T cell|naive T cell
C1369801|T201|MTH_LN|34936-5|LNC|naive T cell|naive T cell
C1369801|T201|LC|34936-5|LNC|naive T cell|naive T cell
C1369801|T201|OSN|34936-5|LNC|naive T cell|naive T cell
C1369886|T201|MTH_LN|35094-2|LNC|pressure|pressure
C1369886|T201|LN|35094-2|LNC|pressure|pressure
C1369886|T201|LC|35094-2|LNC|pressure|pressure
C1369886|T201|OSN|35094-2|LNC|pressure|pressure
C1369886|T201|MTH_LN|35094-2|LNC|systemic pressure|systemic pressure
C1369886|T201|LN|35094-2|LNC|systemic pressure|systemic pressure
C1369886|T201|LC|35094-2|LNC|systemic pressure|systemic pressure
C1369886|T201|OSN|35094-2|LNC|systemic pressure|systemic pressure
C1369946|T201|LN|35157-7|LNC|myristic acid|myristic acid
C1369946|T201|MTH_LN|35157-7|LNC|myristic acid|myristic acid
C1369946|T201|OSN|35157-7|LNC|myristic acid|myristic acid
C1369946|T201|LC|35157-7|LNC|myristic acid|myristic acid
C1369946|T201|LN|35157-7|LNC|tetradecanoic acid|tetradecanoic acid
C1369946|T201|MTH_LN|35157-7|LNC|tetradecanoic acid|tetradecanoic acid
C1369946|T201|OSN|35157-7|LNC|tetradecanoic acid|tetradecanoic acid
C1369946|T201|LC|35157-7|LNC|tetradecanoic acid|tetradecanoic acid
C1370010|T201|MTH_LN|2777-1|LNC|phosphate|phosphate
C1370010|T201|LN|2777-1|LNC|phosphate|phosphate
C1370010|T201|OSN|2777-1|LNC|phosphate|phosphate
C1370010|T201|LC|2777-1|LNC|phosphate|phosphate
C1370010|T201|MTH_LN|2777-1|LNC|phosphate homeostasis|phosphate homeostasis
C1370010|T201|LN|2777-1|LNC|phosphate homeostasis|phosphate homeostasis
C1370010|T201|OSN|2777-1|LNC|phosphate homeostasis|phosphate homeostasis
C1370010|T201|LC|2777-1|LNC|phosphate homeostasis|phosphate homeostasis
C1507518|T201|LN|35384-7|LNC|estradiol|estradiol
C1507518|T201|LC|35384-7|LNC|estradiol|estradiol
C1507518|T201|MTH_LN|35384-7|LNC|estradiol|estradiol
C1507518|T201|OSN|35384-7|LNC|estradiol|estradiol
C1507518|T201|LN|35384-7|LNC|oestradiol|oestradiol
C1507518|T201|LC|35384-7|LNC|oestradiol|oestradiol
C1507518|T201|MTH_LN|35384-7|LNC|oestradiol|oestradiol
C1507518|T201|OSN|35384-7|LNC|oestradiol|oestradiol
C1507674|T201|LN|38230-9|LNC|calcium|calcium
C1507674|T201|OSN|38230-9|LNC|calcium|calcium
C1507674|T201|MTH_LN|38230-9|LNC|calcium|calcium
C1507674|T201|LC|38230-9|LNC|calcium|calcium
C1507674|T201|LN|38230-9|LNC|calcium homeostasis|calcium homeostasis
C1507674|T201|OSN|38230-9|LNC|calcium homeostasis|calcium homeostasis
C1507674|T201|MTH_LN|38230-9|LNC|calcium homeostasis|calcium homeostasis
C1507674|T201|LC|38230-9|LNC|calcium homeostasis|calcium homeostasis
C1507693|T201|LN|38249-9|LNC|C-peptide|C-peptide
C1507693|T201|MTH_LN|38249-9|LNC|C-peptide|C-peptide
C1507693|T201|OSN|38249-9|LNC|C-peptide|C-peptide
C1507693|T201|LC|38249-9|LNC|C-peptide|C-peptide
C1507693|T201|LN|38249-9|LNC|C peptide|C peptide
C1507693|T201|MTH_LN|38249-9|LNC|C peptide|C peptide
C1507693|T201|OSN|38249-9|LNC|C peptide|C peptide
C1507693|T201|LC|38249-9|LNC|C peptide|C peptide
C1507755|T201|LN|35595-8|LNC|xenobiotic|xenobiotic
C1507755|T201|OSN|35595-8|LNC|xenobiotic|xenobiotic
C1507755|T201|MTH_LN|35595-8|LNC|xenobiotic|xenobiotic
C1507755|T201|LC|35595-8|LNC|xenobiotic|xenobiotic
C1507778|T201|LN|35626-1|LNC|xenobiotic|xenobiotic
C1507778|T201|MTH_LN|35626-1|LNC|xenobiotic|xenobiotic
C1507778|T201|OSN|35626-1|LNC|xenobiotic|xenobiotic
C1507778|T201|LC|35626-1|LNC|xenobiotic|xenobiotic
C1507794|T201|LN|35642-8|LNC|cotinine|cotinine
C1507794|T201|LC|35642-8|LNC|cotinine|cotinine
C1507794|T201|MTH_LN|35642-8|LNC|cotinine|cotinine
C1507794|T201|OSN|35642-8|LNC|cotinine|cotinine
C1507814|T201|LN|35663-4|LNC|Protein|Protein
C1507814|T201|LC|35663-4|LNC|Protein|Protein
C1507814|T201|MTH_LN|35663-4|LNC|Protein|Protein
C1507814|T201|OSN|35663-4|LNC|Protein|Protein
C1507826|T201|LN|35675-8|LNC|calcium homeostasis|calcium homeostasis
C1507826|T201|LC|35675-8|LNC|calcium homeostasis|calcium homeostasis
C1507826|T201|MTH_LN|35675-8|LNC|calcium homeostasis|calcium homeostasis
C1507826|T201|OSN|35675-8|LNC|calcium homeostasis|calcium homeostasis
C1526422|T201|LN|38421-4|LNC|C-peptide|C-peptide
C1526422|T201|MTH_LN|38421-4|LNC|C-peptide|C-peptide
C1526422|T201|OSN|38421-4|LNC|C-peptide|C-peptide
C1526422|T201|LC|38421-4|LNC|C-peptide|C-peptide
C1526422|T201|LN|38421-4|LNC|C peptide|C peptide
C1526422|T201|MTH_LN|38421-4|LNC|C peptide|C peptide
C1526422|T201|OSN|38421-4|LNC|C peptide|C peptide
C1526422|T201|LC|38421-4|LNC|C peptide|C peptide
C1526423|T201|LN|38422-2|LNC|C-peptide|C-peptide
C1526423|T201|MTH_LN|38422-2|LNC|C-peptide|C-peptide
C1526423|T201|OSN|38422-2|LNC|C-peptide|C-peptide
C1526423|T201|LC|38422-2|LNC|C-peptide|C-peptide
C1526423|T201|LN|38422-2|LNC|C peptide|C peptide
C1526423|T201|MTH_LN|38422-2|LNC|C peptide|C peptide
C1526423|T201|OSN|38422-2|LNC|C peptide|C peptide
C1526423|T201|LC|38422-2|LNC|C peptide|C peptide
C1526424|T201|LN|38423-0|LNC|C-peptide|C-peptide
C1526424|T201|OSN|38423-0|LNC|C-peptide|C-peptide
C1526424|T201|MTH_LN|38423-0|LNC|C-peptide|C-peptide
C1526424|T201|LC|38423-0|LNC|C-peptide|C-peptide
C1526424|T201|LN|38423-0|LNC|C peptide|C peptide
C1526424|T201|OSN|38423-0|LNC|C peptide|C peptide
C1526424|T201|MTH_LN|38423-0|LNC|C peptide|C peptide
C1526424|T201|LC|38423-0|LNC|C peptide|C peptide
C1526425|T201|LN|38424-8|LNC|C-peptide|C-peptide
C1526425|T201|MTH_LN|38424-8|LNC|C-peptide|C-peptide
C1526425|T201|OSN|38424-8|LNC|C-peptide|C-peptide
C1526425|T201|LC|38424-8|LNC|C-peptide|C-peptide
C1526425|T201|LN|38424-8|LNC|C peptide|C peptide
C1526425|T201|MTH_LN|38424-8|LNC|C peptide|C peptide
C1526425|T201|OSN|38424-8|LNC|C peptide|C peptide
C1526425|T201|LC|38424-8|LNC|C peptide|C peptide
C1526426|T201|LN|38425-5|LNC|C-peptide|C-peptide
C1526426|T201|OSN|38425-5|LNC|C-peptide|C-peptide
C1526426|T201|MTH_LN|38425-5|LNC|C-peptide|C-peptide
C1526426|T201|LC|38425-5|LNC|C-peptide|C-peptide
C1526426|T201|LN|38425-5|LNC|C peptide|C peptide
C1526426|T201|OSN|38425-5|LNC|C peptide|C peptide
C1526426|T201|MTH_LN|38425-5|LNC|C peptide|C peptide
C1526426|T201|LC|38425-5|LNC|C peptide|C peptide
C1526427|T201|LN|38426-3|LNC|C-peptide|C-peptide
C1526427|T201|MTH_LN|38426-3|LNC|C-peptide|C-peptide
C1526427|T201|OSN|38426-3|LNC|C-peptide|C-peptide
C1526427|T201|LC|38426-3|LNC|C-peptide|C-peptide
C1526427|T201|LN|38426-3|LNC|C peptide|C peptide
C1526427|T201|MTH_LN|38426-3|LNC|C peptide|C peptide
C1526427|T201|OSN|38426-3|LNC|C peptide|C peptide
C1526427|T201|LC|38426-3|LNC|C peptide|C peptide
C1526475|T201|LN|38474-3|LNC|acylcarnitine|acylcarnitine
C1526475|T201|LC|38474-3|LNC|acylcarnitine|acylcarnitine
C1526475|T201|MTH_LN|38474-3|LNC|acylcarnitine|acylcarnitine
C1526475|T201|OSN|38474-3|LNC|acylcarnitine|acylcarnitine
C1526477|T201|LN|38476-8|LNC|antimullerian|antimullerian
C1526477|T201|MTH_LN|38476-8|LNC|antimullerian|antimullerian
C1526477|T201|OSN|38476-8|LNC|antimullerian|antimullerian
C1526477|T201|LC|38476-8|LNC|antimullerian|antimullerian
C1526477|T201|LN|38476-8|LNC|AMH|AMH
C1526477|T201|MTH_LN|38476-8|LNC|AMH|AMH
C1526477|T201|OSN|38476-8|LNC|AMH|AMH
C1526477|T201|LC|38476-8|LNC|AMH|AMH
C1526484|T201|LN|38483-4|LNC|creatinine|creatinine
C1526484|T201|OSN|38483-4|LNC|creatinine|creatinine
C1526484|T201|MTH_LN|38483-4|LNC|creatinine|creatinine
C1526484|T201|LC|38483-4|LNC|creatinine|creatinine
C1526494|T201|LN|38493-3|LNC|ketone bodies|ketone bodies
C1526494|T201|MTH_LN|38493-3|LNC|ketone bodies|ketone bodies
C1526494|T201|OSN|38493-3|LNC|ketone bodies|ketone bodies
C1526494|T201|LC|38493-3|LNC|ketone bodies|ketone bodies
C1526505|T201|LN|38504-7|LNC|Autoimmune antibody|Autoimmune antibody
C1526505|T201|OSN|38504-7|LNC|Autoimmune antibody|Autoimmune antibody
C1526505|T201|MTH_LN|38504-7|LNC|Autoimmune antibody|Autoimmune antibody
C1526505|T201|LC|38504-7|LNC|Autoimmune antibody|Autoimmune antibody
C1526553|T201|LN|38552-6|LNC|acylcarnitine|acylcarnitine
C1526553|T201|MTH_LN|38552-6|LNC|acylcarnitine|acylcarnitine
C1526553|T201|OSN|38552-6|LNC|acylcarnitine|acylcarnitine
C1526553|T201|LC|38552-6|LNC|acylcarnitine|acylcarnitine
C1543545|T201|LN|39469-2|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1543545|T201|OSN|39469-2|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1543545|T201|MTH_LN|39469-2|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1543545|T201|LC|39469-2|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1543545|T201|LN|39469-2|LNC|LDL|LDL
C1543545|T201|OSN|39469-2|LNC|LDL|LDL
C1543545|T201|MTH_LN|39469-2|LNC|LDL|LDL
C1543545|T201|LC|39469-2|LNC|LDL|LDL
C1543545|T201|LN|39469-2|LNC|LDL cholesterol|LDL cholesterol
C1543545|T201|OSN|39469-2|LNC|LDL cholesterol|LDL cholesterol
C1543545|T201|MTH_LN|39469-2|LNC|LDL cholesterol|LDL cholesterol
C1543545|T201|LC|39469-2|LNC|LDL cholesterol|LDL cholesterol
C1543545|T201|LN|39469-2|LNC|low-density lipoprotein|low-density lipoprotein
C1543545|T201|OSN|39469-2|LNC|low-density lipoprotein|low-density lipoprotein
C1543545|T201|MTH_LN|39469-2|LNC|low-density lipoprotein|low-density lipoprotein
C1543545|T201|LC|39469-2|LNC|low-density lipoprotein|low-density lipoprotein
C1543545|T201|LN|39469-2|LNC|beta-lipoproteins|beta-lipoproteins
C1543545|T201|OSN|39469-2|LNC|beta-lipoproteins|beta-lipoproteins
C1543545|T201|MTH_LN|39469-2|LNC|beta-lipoproteins|beta-lipoproteins
C1543545|T201|LC|39469-2|LNC|beta-lipoproteins|beta-lipoproteins
C1543545|T201|LN|39469-2|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1543545|T201|OSN|39469-2|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1543545|T201|MTH_LN|39469-2|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1543545|T201|LC|39469-2|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1543545|T201|LN|39469-2|LNC|LDL-C|LDL-C
C1543545|T201|OSN|39469-2|LNC|LDL-C|LDL-C
C1543545|T201|MTH_LN|39469-2|LNC|LDL-C|LDL-C
C1543545|T201|LC|39469-2|LNC|LDL-C|LDL-C
C1543636|T201|LN|39561-6|LNC|glucose|glucose
C1543636|T201|MTH_LN|39561-6|LNC|glucose|glucose
C1543636|T201|OSN|39561-6|LNC|glucose|glucose
C1543636|T201|LC|39561-6|LNC|glucose|glucose
C1543637|T201|LN|39562-4|LNC|glucose|glucose
C1543637|T201|MTH_LN|39562-4|LNC|glucose|glucose
C1543637|T201|OSN|39562-4|LNC|glucose|glucose
C1543637|T201|LC|39562-4|LNC|glucose|glucose
C1543638|T201|LN|39563-2|LNC|glucose|glucose
C1543638|T201|MTH_LN|39563-2|LNC|glucose|glucose
C1543638|T201|OSN|39563-2|LNC|glucose|glucose
C1543638|T201|LC|39563-2|LNC|glucose|glucose
C1543831|T201|LN|39789-3|LNC|potassium|potassium
C1543831|T201|OSN|39789-3|LNC|potassium|potassium
C1543831|T201|MTH_LN|39789-3|LNC|potassium|potassium
C1543831|T201|LC|39789-3|LNC|potassium|potassium
C1543831|T201|LN|39789-3|LNC|potassium homeostasis|potassium homeostasis
C1543831|T201|OSN|39789-3|LNC|potassium homeostasis|potassium homeostasis
C1543831|T201|MTH_LN|39789-3|LNC|potassium homeostasis|potassium homeostasis
C1543831|T201|LC|39789-3|LNC|potassium homeostasis|potassium homeostasis
C1544348|T201|LN|40373-3|LNC|luteinizing|luteinizing
C1544348|T201|MTH_LN|40373-3|LNC|luteinizing|luteinizing
C1544348|T201|OSN|40373-3|LNC|luteinizing|luteinizing
C1544348|T201|LC|40373-3|LNC|luteinizing|luteinizing
C1544348|T201|LN|40373-3|LNC|LH|LH
C1544348|T201|MTH_LN|40373-3|LNC|LH|LH
C1544348|T201|OSN|40373-3|LNC|LH|LH
C1544348|T201|LC|40373-3|LNC|LH|LH
C1544348|T201|LN|40373-3|LNC|luteinising|luteinising
C1544348|T201|MTH_LN|40373-3|LNC|luteinising|luteinising
C1544348|T201|OSN|40373-3|LNC|luteinising|luteinising
C1544348|T201|LC|40373-3|LNC|luteinising|luteinising
C1544349|T201|LN|40374-1|LNC|luteinizing|luteinizing
C1544349|T201|MTH_LN|40374-1|LNC|luteinizing|luteinizing
C1544349|T201|OSN|40374-1|LNC|luteinizing|luteinizing
C1544349|T201|LC|40374-1|LNC|luteinizing|luteinizing
C1544349|T201|LN|40374-1|LNC|LH|LH
C1544349|T201|MTH_LN|40374-1|LNC|LH|LH
C1544349|T201|OSN|40374-1|LNC|LH|LH
C1544349|T201|LC|40374-1|LNC|LH|LH
C1544349|T201|LN|40374-1|LNC|luteinising|luteinising
C1544349|T201|MTH_LN|40374-1|LNC|luteinising|luteinising
C1544349|T201|OSN|40374-1|LNC|luteinising|luteinising
C1544349|T201|LC|40374-1|LNC|luteinising|luteinising
C1544350|T201|LN|40375-8|LNC|luteinizing|luteinizing
C1544350|T201|MTH_LN|40375-8|LNC|luteinizing|luteinizing
C1544350|T201|OSN|40375-8|LNC|luteinizing|luteinizing
C1544350|T201|LC|40375-8|LNC|luteinizing|luteinizing
C1544350|T201|LN|40375-8|LNC|LH|LH
C1544350|T201|MTH_LN|40375-8|LNC|LH|LH
C1544350|T201|OSN|40375-8|LNC|LH|LH
C1544350|T201|LC|40375-8|LNC|LH|LH
C1544350|T201|LN|40375-8|LNC|luteinising|luteinising
C1544350|T201|MTH_LN|40375-8|LNC|luteinising|luteinising
C1544350|T201|OSN|40375-8|LNC|luteinising|luteinising
C1544350|T201|LC|40375-8|LNC|luteinising|luteinising
C1544351|T201|LN|40376-6|LNC|luteinizing|luteinizing
C1544351|T201|MTH_LN|40376-6|LNC|luteinizing|luteinizing
C1544351|T201|OSN|40376-6|LNC|luteinizing|luteinizing
C1544351|T201|LC|40376-6|LNC|luteinizing|luteinizing
C1544351|T201|LN|40376-6|LNC|LH|LH
C1544351|T201|MTH_LN|40376-6|LNC|LH|LH
C1544351|T201|OSN|40376-6|LNC|LH|LH
C1544351|T201|LC|40376-6|LNC|LH|LH
C1544351|T201|LN|40376-6|LNC|luteinising|luteinising
C1544351|T201|MTH_LN|40376-6|LNC|luteinising|luteinising
C1544351|T201|OSN|40376-6|LNC|luteinising|luteinising
C1544351|T201|LC|40376-6|LNC|luteinising|luteinising
C1544352|T201|LN|40377-4|LNC|luteinizing|luteinizing
C1544352|T201|MTH_LN|40377-4|LNC|luteinizing|luteinizing
C1544352|T201|OSN|40377-4|LNC|luteinizing|luteinizing
C1544352|T201|LC|40377-4|LNC|luteinizing|luteinizing
C1544352|T201|LN|40377-4|LNC|LH|LH
C1544352|T201|MTH_LN|40377-4|LNC|LH|LH
C1544352|T201|OSN|40377-4|LNC|LH|LH
C1544352|T201|LC|40377-4|LNC|LH|LH
C1544352|T201|LN|40377-4|LNC|luteinising|luteinising
C1544352|T201|MTH_LN|40377-4|LNC|luteinising|luteinising
C1544352|T201|OSN|40377-4|LNC|luteinising|luteinising
C1544352|T201|LC|40377-4|LNC|luteinising|luteinising
C1544353|T201|LN|40378-2|LNC|luteinizing|luteinizing
C1544353|T201|MTH_LN|40378-2|LNC|luteinizing|luteinizing
C1544353|T201|OSN|40378-2|LNC|luteinizing|luteinizing
C1544353|T201|LC|40378-2|LNC|luteinizing|luteinizing
C1544353|T201|LN|40378-2|LNC|LH|LH
C1544353|T201|MTH_LN|40378-2|LNC|LH|LH
C1544353|T201|OSN|40378-2|LNC|LH|LH
C1544353|T201|LC|40378-2|LNC|LH|LH
C1544353|T201|LN|40378-2|LNC|luteinising|luteinising
C1544353|T201|MTH_LN|40378-2|LNC|luteinising|luteinising
C1544353|T201|OSN|40378-2|LNC|luteinising|luteinising
C1544353|T201|LC|40378-2|LNC|luteinising|luteinising
C1544620|T201|LN|40665-2|LNC|reticulocytes|reticulocytes
C1544620|T201|OSN|40665-2|LNC|reticulocytes|reticulocytes
C1544620|T201|MTH_LN|40665-2|LNC|reticulocytes|reticulocytes
C1544620|T201|LC|40665-2|LNC|reticulocytes|reticulocytes
C1544620|T201|LN|40665-2|LNC|reticulocyte count|reticulocyte count
C1544620|T201|OSN|40665-2|LNC|reticulocyte count|reticulocyte count
C1544620|T201|MTH_LN|40665-2|LNC|reticulocyte count|reticulocyte count
C1544620|T201|LC|40665-2|LNC|reticulocyte count|reticulocyte count
C1544784|T201|LN|40829-4|LNC|ornithine|ornithine
C1544784|T201|MTH_LN|40829-4|LNC|ornithine|ornithine
C1544784|T201|OSN|40829-4|LNC|ornithine|ornithine
C1544784|T201|LC|40829-4|LNC|ornithine|ornithine
C1544784|T201|LN|40829-4|LNC|ornithine metabolism|ornithine metabolism
C1544784|T201|MTH_LN|40829-4|LNC|ornithine metabolism|ornithine metabolism
C1544784|T201|OSN|40829-4|LNC|ornithine metabolism|ornithine metabolism
C1544784|T201|LC|40829-4|LNC|ornithine metabolism|ornithine metabolism
C1544987|T201|LN|41040-7|LNC|acylcarnitine|acylcarnitine
C1544987|T201|OSN|41040-7|LNC|acylcarnitine|acylcarnitine
C1544987|T201|MTH_LN|41040-7|LNC|acylcarnitine|acylcarnitine
C1544987|T201|LC|41040-7|LNC|acylcarnitine|acylcarnitine
C1551421|T098|LN|1358-1|LNC|adrenocorticotropin|adrenocorticotropin
C1551421|T098|OSN|1358-1|LNC|adrenocorticotropin|adrenocorticotropin
C1551421|T098|MTH_LN|1358-1|LNC|adrenocorticotropin|adrenocorticotropin
C1551421|T098|LC|1358-1|LNC|adrenocorticotropin|adrenocorticotropin
C1551421|T098|LN|1358-1|LNC|ACTH|ACTH
C1551421|T098|OSN|1358-1|LNC|ACTH|ACTH
C1551421|T098|MTH_LN|1358-1|LNC|ACTH|ACTH
C1551421|T098|LC|1358-1|LNC|ACTH|ACTH
C1551422|T098|LN|1359-9|LNC|adrenocorticotropin|adrenocorticotropin
C1551422|T098|MTH_LN|1359-9|LNC|adrenocorticotropin|adrenocorticotropin
C1551422|T098|OSN|1359-9|LNC|adrenocorticotropin|adrenocorticotropin
C1551422|T098|LC|1359-9|LNC|adrenocorticotropin|adrenocorticotropin
C1551422|T098|LN|1359-9|LNC|ACTH|ACTH
C1551422|T098|MTH_LN|1359-9|LNC|ACTH|ACTH
C1551422|T098|OSN|1359-9|LNC|ACTH|ACTH
C1551422|T098|LC|1359-9|LNC|ACTH|ACTH
C1551423|T098|LN|1360-7|LNC|adrenocorticotropin|adrenocorticotropin
C1551423|T098|MTH_LN|1360-7|LNC|adrenocorticotropin|adrenocorticotropin
C1551423|T098|OSN|1360-7|LNC|adrenocorticotropin|adrenocorticotropin
C1551423|T098|LC|1360-7|LNC|adrenocorticotropin|adrenocorticotropin
C1551423|T098|LN|1360-7|LNC|ACTH|ACTH
C1551423|T098|MTH_LN|1360-7|LNC|ACTH|ACTH
C1551423|T098|OSN|1360-7|LNC|ACTH|ACTH
C1551423|T098|LC|1360-7|LNC|ACTH|ACTH
C1551424|T098|LN|1361-5|LNC|adrenocorticotropin|adrenocorticotropin
C1551424|T098|MTH_LN|1361-5|LNC|adrenocorticotropin|adrenocorticotropin
C1551424|T098|OSN|1361-5|LNC|adrenocorticotropin|adrenocorticotropin
C1551424|T098|LC|1361-5|LNC|adrenocorticotropin|adrenocorticotropin
C1551424|T098|LN|1361-5|LNC|ACTH|ACTH
C1551424|T098|MTH_LN|1361-5|LNC|ACTH|ACTH
C1551424|T098|OSN|1361-5|LNC|ACTH|ACTH
C1551424|T098|LC|1361-5|LNC|ACTH|ACTH
C1551425|T098|LN|1363-1|LNC|adrenocorticotropin|adrenocorticotropin
C1551425|T098|MTH_LN|1363-1|LNC|adrenocorticotropin|adrenocorticotropin
C1551425|T098|OSN|1363-1|LNC|adrenocorticotropin|adrenocorticotropin
C1551425|T098|LC|1363-1|LNC|adrenocorticotropin|adrenocorticotropin
C1551425|T098|LN|1363-1|LNC|ACTH|ACTH
C1551425|T098|MTH_LN|1363-1|LNC|ACTH|ACTH
C1551425|T098|OSN|1363-1|LNC|ACTH|ACTH
C1551425|T098|LC|1363-1|LNC|ACTH|ACTH
C1551426|T098|LN|1365-6|LNC|adrenocorticotropin|adrenocorticotropin
C1551426|T098|MTH_LN|1365-6|LNC|adrenocorticotropin|adrenocorticotropin
C1551426|T098|OSN|1365-6|LNC|adrenocorticotropin|adrenocorticotropin
C1551426|T098|LC|1365-6|LNC|adrenocorticotropin|adrenocorticotropin
C1551426|T098|LN|1365-6|LNC|ACTH|ACTH
C1551426|T098|MTH_LN|1365-6|LNC|ACTH|ACTH
C1551426|T098|OSN|1365-6|LNC|ACTH|ACTH
C1551426|T098|LC|1365-6|LNC|ACTH|ACTH
C1551427|T098|LN|1366-4|LNC|adrenocorticotropin|adrenocorticotropin
C1551427|T098|MTH_LN|1366-4|LNC|adrenocorticotropin|adrenocorticotropin
C1551427|T098|OSN|1366-4|LNC|adrenocorticotropin|adrenocorticotropin
C1551427|T098|LC|1366-4|LNC|adrenocorticotropin|adrenocorticotropin
C1551427|T098|LN|1366-4|LNC|ACTH|ACTH
C1551427|T098|MTH_LN|1366-4|LNC|ACTH|ACTH
C1551427|T098|OSN|1366-4|LNC|ACTH|ACTH
C1551427|T098|LC|1366-4|LNC|ACTH|ACTH
C1551428|T098|LN|1368-0|LNC|adrenocorticotropin|adrenocorticotropin
C1551428|T098|MTH_LN|1368-0|LNC|adrenocorticotropin|adrenocorticotropin
C1551428|T098|OSN|1368-0|LNC|adrenocorticotropin|adrenocorticotropin
C1551428|T098|LC|1368-0|LNC|adrenocorticotropin|adrenocorticotropin
C1551428|T098|LN|1368-0|LNC|ACTH|ACTH
C1551428|T098|MTH_LN|1368-0|LNC|ACTH|ACTH
C1551428|T098|OSN|1368-0|LNC|ACTH|ACTH
C1551428|T098|LC|1368-0|LNC|ACTH|ACTH
C1551438|T098|LN|1389-6|LNC|cortisol|cortisol
C1551438|T098|MTH_LN|1389-6|LNC|cortisol|cortisol
C1551438|T098|OSN|1389-6|LNC|cortisol|cortisol
C1551438|T098|LC|1389-6|LNC|cortisol|cortisol
// C1551438|T098|LN|1389-6|LNC||
// C1551438|T098|MTH_LN|1389-6|LNC||
// C1551438|T098|OSN|1389-6|LNC||
// C1551438|T098|LC|1389-6|LNC||
C1551441|T098|LN|1393-8|LNC|cortisol|cortisol
C1551441|T098|MTH_LN|1393-8|LNC|cortisol|cortisol
C1551441|T098|OSN|1393-8|LNC|cortisol|cortisol
C1551441|T098|LC|1393-8|LNC|cortisol|cortisol
// C1551441|T098|LN|1393-8|LNC||
// C1551441|T098|MTH_LN|1393-8|LNC||
// C1551441|T098|OSN|1393-8|LNC||
// C1551441|T098|LC|1393-8|LNC||
C1551442|T098|LN|1394-6|LNC|cortisol|cortisol
C1551442|T098|MTH_LN|1394-6|LNC|cortisol|cortisol
C1551442|T098|OSN|1394-6|LNC|cortisol|cortisol
C1551442|T098|LC|1394-6|LNC|cortisol|cortisol
// C1551442|T098|LN|1394-6|LNC||
// C1551442|T098|MTH_LN|1394-6|LNC||
// C1551442|T098|OSN|1394-6|LNC||
// C1551442|T098|LC|1394-6|LNC||
C1551449|T098|LN|1401-9|LNC|cortisol|cortisol
C1551449|T098|MTH_LN|1401-9|LNC|cortisol|cortisol
C1551449|T098|OSN|1401-9|LNC|cortisol|cortisol
C1551449|T098|LC|1401-9|LNC|cortisol|cortisol
C1551449|T098|LN|1401-9|LNC|cortisol low|cortisol low
C1551449|T098|MTH_LN|1401-9|LNC|cortisol low|cortisol low
C1551449|T098|OSN|1401-9|LNC|cortisol low|cortisol low
C1551449|T098|LC|1401-9|LNC|cortisol low|cortisol low
C1551449|T098|LN|1401-9|LNC|to undetectable cortisol|to undetectable cortisol
C1551449|T098|MTH_LN|1401-9|LNC|to undetectable cortisol|to undetectable cortisol
C1551449|T098|OSN|1401-9|LNC|to undetectable cortisol|to undetectable cortisol
C1551449|T098|LC|1401-9|LNC|to undetectable cortisol|to undetectable cortisol
C1551450|T098|LN|1403-5|LNC|cortisol|cortisol
C1551450|T098|MTH_LN|1403-5|LNC|cortisol|cortisol
C1551450|T098|OSN|1403-5|LNC|cortisol|cortisol
C1551450|T098|LC|1403-5|LNC|cortisol|cortisol
C1551450|T098|LN|1403-5|LNC|cortisol low|cortisol low
C1551450|T098|MTH_LN|1403-5|LNC|cortisol low|cortisol low
C1551450|T098|OSN|1403-5|LNC|cortisol low|cortisol low
C1551450|T098|LC|1403-5|LNC|cortisol low|cortisol low
C1551450|T098|LN|1403-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551450|T098|MTH_LN|1403-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551450|T098|OSN|1403-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551450|T098|LC|1403-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551453|T098|LN|1409-2|LNC|cortisol|cortisol
C1551453|T098|MTH_LN|1409-2|LNC|cortisol|cortisol
C1551453|T098|OSN|1409-2|LNC|cortisol|cortisol
C1551453|T098|LC|1409-2|LNC|cortisol|cortisol
C1551453|T098|LN|1409-2|LNC|cortisol low|cortisol low
C1551453|T098|MTH_LN|1409-2|LNC|cortisol low|cortisol low
C1551453|T098|OSN|1409-2|LNC|cortisol low|cortisol low
C1551453|T098|LC|1409-2|LNC|cortisol low|cortisol low
C1551453|T098|LN|1409-2|LNC|to undetectable cortisol|to undetectable cortisol
C1551453|T098|MTH_LN|1409-2|LNC|to undetectable cortisol|to undetectable cortisol
C1551453|T098|OSN|1409-2|LNC|to undetectable cortisol|to undetectable cortisol
C1551453|T098|LC|1409-2|LNC|to undetectable cortisol|to undetectable cortisol
C1551456|T098|LN|1413-4|LNC|cortisol|cortisol
C1551456|T098|MTH_LN|1413-4|LNC|cortisol|cortisol
C1551456|T098|OSN|1413-4|LNC|cortisol|cortisol
C1551456|T098|LC|1413-4|LNC|cortisol|cortisol
C1551456|T098|LN|1413-4|LNC|cortisol low|cortisol low
C1551456|T098|MTH_LN|1413-4|LNC|cortisol low|cortisol low
C1551456|T098|OSN|1413-4|LNC|cortisol low|cortisol low
C1551456|T098|LC|1413-4|LNC|cortisol low|cortisol low
C1551456|T098|LN|1413-4|LNC|to undetectable cortisol|to undetectable cortisol
C1551456|T098|MTH_LN|1413-4|LNC|to undetectable cortisol|to undetectable cortisol
C1551456|T098|OSN|1413-4|LNC|to undetectable cortisol|to undetectable cortisol
C1551456|T098|LC|1413-4|LNC|to undetectable cortisol|to undetectable cortisol
C1551458|T098|LN|1417-5|LNC|cortisol|cortisol
C1551458|T098|MTH_LN|1417-5|LNC|cortisol|cortisol
C1551458|T098|OSN|1417-5|LNC|cortisol|cortisol
C1551458|T098|LC|1417-5|LNC|cortisol|cortisol
C1551458|T098|LN|1417-5|LNC|cortisol low|cortisol low
C1551458|T098|MTH_LN|1417-5|LNC|cortisol low|cortisol low
C1551458|T098|OSN|1417-5|LNC|cortisol low|cortisol low
C1551458|T098|LC|1417-5|LNC|cortisol low|cortisol low
C1551458|T098|LN|1417-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551458|T098|MTH_LN|1417-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551458|T098|OSN|1417-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551458|T098|LC|1417-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551459|T098|LN|1418-3|LNC|cortisol|cortisol
C1551459|T098|MTH_LN|1418-3|LNC|cortisol|cortisol
C1551459|T098|OSN|1418-3|LNC|cortisol|cortisol
C1551459|T098|LC|1418-3|LNC|cortisol|cortisol
C1551459|T098|LN|1418-3|LNC|cortisol low|cortisol low
C1551459|T098|MTH_LN|1418-3|LNC|cortisol low|cortisol low
C1551459|T098|OSN|1418-3|LNC|cortisol low|cortisol low
C1551459|T098|LC|1418-3|LNC|cortisol low|cortisol low
C1551459|T098|LN|1418-3|LNC|to undetectable cortisol|to undetectable cortisol
C1551459|T098|MTH_LN|1418-3|LNC|to undetectable cortisol|to undetectable cortisol
C1551459|T098|OSN|1418-3|LNC|to undetectable cortisol|to undetectable cortisol
C1551459|T098|LC|1418-3|LNC|to undetectable cortisol|to undetectable cortisol
C1551462|T098|LN|1421-7|LNC|cortisol|cortisol
C1551462|T098|MTH_LN|1421-7|LNC|cortisol|cortisol
C1551462|T098|OSN|1421-7|LNC|cortisol|cortisol
C1551462|T098|LC|1421-7|LNC|cortisol|cortisol
C1551462|T098|LN|1421-7|LNC|cortisol low|cortisol low
C1551462|T098|MTH_LN|1421-7|LNC|cortisol low|cortisol low
C1551462|T098|OSN|1421-7|LNC|cortisol low|cortisol low
C1551462|T098|LC|1421-7|LNC|cortisol low|cortisol low
C1551462|T098|LN|1421-7|LNC|to undetectable cortisol|to undetectable cortisol
C1551462|T098|MTH_LN|1421-7|LNC|to undetectable cortisol|to undetectable cortisol
C1551462|T098|OSN|1421-7|LNC|to undetectable cortisol|to undetectable cortisol
C1551462|T098|LC|1421-7|LNC|to undetectable cortisol|to undetectable cortisol
C1551463|T098|LN|1422-5|LNC|cortisol|cortisol
C1551463|T098|MTH_LN|1422-5|LNC|cortisol|cortisol
C1551463|T098|OSN|1422-5|LNC|cortisol|cortisol
C1551463|T098|LC|1422-5|LNC|cortisol|cortisol
C1551463|T098|LN|1422-5|LNC|cortisol low|cortisol low
C1551463|T098|MTH_LN|1422-5|LNC|cortisol low|cortisol low
C1551463|T098|OSN|1422-5|LNC|cortisol low|cortisol low
C1551463|T098|LC|1422-5|LNC|cortisol low|cortisol low
C1551463|T098|LN|1422-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551463|T098|MTH_LN|1422-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551463|T098|OSN|1422-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551463|T098|LC|1422-5|LNC|to undetectable cortisol|to undetectable cortisol
C1551467|T098|LN|1426-6|LNC|cortisol|cortisol
C1551467|T098|MTH_LN|1426-6|LNC|cortisol|cortisol
C1551467|T098|OSN|1426-6|LNC|cortisol|cortisol
C1551467|T098|LC|1426-6|LNC|cortisol|cortisol
C1551467|T098|LN|1426-6|LNC|cortisol low|cortisol low
C1551467|T098|MTH_LN|1426-6|LNC|cortisol low|cortisol low
C1551467|T098|OSN|1426-6|LNC|cortisol low|cortisol low
C1551467|T098|LC|1426-6|LNC|cortisol low|cortisol low
C1551467|T098|LN|1426-6|LNC|to undetectable cortisol|to undetectable cortisol
C1551467|T098|MTH_LN|1426-6|LNC|to undetectable cortisol|to undetectable cortisol
C1551467|T098|OSN|1426-6|LNC|to undetectable cortisol|to undetectable cortisol
C1551467|T098|LC|1426-6|LNC|to undetectable cortisol|to undetectable cortisol
C1551471|T098|LN|1430-8|LNC|cortisol|cortisol
C1551471|T098|MTH_LN|1430-8|LNC|cortisol|cortisol
C1551471|T098|OSN|1430-8|LNC|cortisol|cortisol
C1551471|T098|LC|1430-8|LNC|cortisol|cortisol
C1551471|T098|LN|1430-8|LNC|cortisol low|cortisol low
C1551471|T098|MTH_LN|1430-8|LNC|cortisol low|cortisol low
C1551471|T098|OSN|1430-8|LNC|cortisol low|cortisol low
C1551471|T098|LC|1430-8|LNC|cortisol low|cortisol low
C1551471|T098|LN|1430-8|LNC|to undetectable cortisol|to undetectable cortisol
C1551471|T098|MTH_LN|1430-8|LNC|to undetectable cortisol|to undetectable cortisol
C1551471|T098|OSN|1430-8|LNC|to undetectable cortisol|to undetectable cortisol
C1551471|T098|LC|1430-8|LNC|to undetectable cortisol|to undetectable cortisol
C1551510|T098|LN|1483-7|LNC|galactose|galactose
C1551510|T098|MTH_LN|1483-7|LNC|galactose|galactose
C1551510|T098|OSN|1483-7|LNC|galactose|galactose
C1551510|T098|LC|1483-7|LNC|galactose|galactose
C1551515|T098|LN|1491-0|LNC|glucose|glucose
C1551515|T098|MTH_LN|1491-0|LNC|glucose|glucose
C1551515|T098|OSN|1491-0|LNC|glucose|glucose
C1551515|T098|LC|1491-0|LNC|glucose|glucose
C1551516|T098|LN|1492-8|LNC|glucose|glucose
C1551516|T098|OSN|1492-8|LNC|glucose|glucose
C1551516|T098|MTH_LN|1492-8|LNC|glucose|glucose
C1551516|T098|LC|1492-8|LNC|glucose|glucose
C1551517|T098|LN|1494-4|LNC|glucose|glucose
C1551517|T098|OSN|1494-4|LNC|glucose|glucose
C1551517|T098|MTH_LN|1494-4|LNC|glucose|glucose
C1551517|T098|LC|1494-4|LNC|glucose|glucose
C1551518|T098|LN|1495-1|LNC|glucose|glucose
C1551518|T098|OSN|1495-1|LNC|glucose|glucose
C1551518|T098|MTH_LN|1495-1|LNC|glucose|glucose
C1551518|T098|LC|1495-1|LNC|glucose|glucose
C1551519|T098|LN|1496-9|LNC|glucose|glucose
C1551519|T098|OSN|1496-9|LNC|glucose|glucose
C1551519|T098|MTH_LN|1496-9|LNC|glucose|glucose
C1551519|T098|LC|1496-9|LNC|glucose|glucose
C1551520|T098|LN|1497-7|LNC|glucose|glucose
C1551520|T098|OSN|1497-7|LNC|glucose|glucose
C1551520|T098|MTH_LN|1497-7|LNC|glucose|glucose
C1551520|T098|LC|1497-7|LNC|glucose|glucose
C1551521|T098|LN|1498-5|LNC|glucose|glucose
C1551521|T098|MTH_LN|1498-5|LNC|glucose|glucose
C1551521|T098|OSN|1498-5|LNC|glucose|glucose
C1551521|T098|LC|1498-5|LNC|glucose|glucose
C1551522|T098|LN|1499-3|LNC|glucose|glucose
C1551522|T098|MTH_LN|1499-3|LNC|glucose|glucose
C1551522|T098|OSN|1499-3|LNC|glucose|glucose
C1551522|T098|LC|1499-3|LNC|glucose|glucose
C1551523|T098|LN|1500-8|LNC|glucose|glucose
C1551523|T098|MTH_LN|1500-8|LNC|glucose|glucose
C1551523|T098|OSN|1500-8|LNC|glucose|glucose
C1551523|T098|LC|1500-8|LNC|glucose|glucose
C1551524|T098|LN|1501-6|LNC|glucose|glucose
C1551524|T098|MTH_LN|1501-6|LNC|glucose|glucose
C1551524|T098|OSN|1501-6|LNC|glucose|glucose
C1551524|T098|LC|1501-6|LNC|glucose|glucose
C1551526|T098|LN|1503-2|LNC|glucose|glucose
C1551526|T098|MTH_LN|1503-2|LNC|glucose|glucose
C1551526|T098|OSN|1503-2|LNC|glucose|glucose
C1551526|T098|LC|1503-2|LNC|glucose|glucose
C1551527|T098|LN|1504-0|LNC|glucose|glucose
C1551527|T098|MTH_LN|1504-0|LNC|glucose|glucose
C1551527|T098|OSN|1504-0|LNC|glucose|glucose
C1551527|T098|LC|1504-0|LNC|glucose|glucose
C1551528|T098|LN|1505-7|LNC|glucose|glucose
C1551528|T098|MTH_LN|1505-7|LNC|glucose|glucose
C1551528|T098|OSN|1505-7|LNC|glucose|glucose
C1551528|T098|LC|1505-7|LNC|glucose|glucose
C1551529|T098|LN|1506-5|LNC|glucose|glucose
C1551529|T098|MTH_LN|1506-5|LNC|glucose|glucose
C1551529|T098|OSN|1506-5|LNC|glucose|glucose
C1551529|T098|LC|1506-5|LNC|glucose|glucose
C1551530|T098|LN|1507-3|LNC|glucose|glucose
C1551530|T098|MTH_LN|1507-3|LNC|glucose|glucose
C1551530|T098|OSN|1507-3|LNC|glucose|glucose
C1551530|T098|LC|1507-3|LNC|glucose|glucose
C1551532|T098|LN|1509-9|LNC|glucose|glucose
C1551532|T098|MTH_LN|1509-9|LNC|glucose|glucose
C1551532|T098|OSN|1509-9|LNC|glucose|glucose
C1551532|T098|LC|1509-9|LNC|glucose|glucose
C1551533|T098|MTH_LN|1510-7|LNC|glucose|glucose
C1551533|T098|LN|1510-7|LNC|glucose|glucose
C1551533|T098|OSN|1510-7|LNC|glucose|glucose
C1551533|T098|LC|1510-7|LNC|glucose|glucose
C1551535|T098|LN|1512-3|LNC|glucose|glucose
C1551535|T098|MTH_LN|1512-3|LNC|glucose|glucose
C1551535|T098|OSN|1512-3|LNC|glucose|glucose
C1551535|T098|LC|1512-3|LNC|glucose|glucose
C1551536|T098|LN|1513-1|LNC|glucose|glucose
C1551536|T098|MTH_LN|1513-1|LNC|glucose|glucose
C1551536|T098|OSN|1513-1|LNC|glucose|glucose
C1551536|T098|LC|1513-1|LNC|glucose|glucose
C1551537|T098|LN|1514-9|LNC|glucose|glucose
C1551537|T098|MTH_LN|1514-9|LNC|glucose|glucose
C1551537|T098|OSN|1514-9|LNC|glucose|glucose
C1551537|T098|LC|1514-9|LNC|glucose|glucose
C1551539|T098|LN|1518-0|LNC|glucose|glucose
C1551539|T098|MTH_LN|1518-0|LNC|glucose|glucose
C1551539|T098|OSN|1518-0|LNC|glucose|glucose
C1551539|T098|LC|1518-0|LNC|glucose|glucose
C1551541|T098|LN|1520-6|LNC|glucose|glucose
C1551541|T098|MTH_LN|1520-6|LNC|glucose|glucose
C1551541|T098|OSN|1520-6|LNC|glucose|glucose
C1551541|T098|LC|1520-6|LNC|glucose|glucose
C1551542|T098|LN|1521-4|LNC|glucose|glucose
C1551542|T098|MTH_LN|1521-4|LNC|glucose|glucose
C1551542|T098|OSN|1521-4|LNC|glucose|glucose
C1551542|T098|LC|1521-4|LNC|glucose|glucose
C1551543|T098|LN|1522-2|LNC|glucose|glucose
C1551543|T098|MTH_LN|1522-2|LNC|glucose|glucose
C1551543|T098|OSN|1522-2|LNC|glucose|glucose
C1551543|T098|LC|1522-2|LNC|glucose|glucose
C1551544|T098|LN|1523-0|LNC|glucose|glucose
C1551544|T098|MTH_LN|1523-0|LNC|glucose|glucose
C1551544|T098|OSN|1523-0|LNC|glucose|glucose
C1551544|T098|LC|1523-0|LNC|glucose|glucose
C1551545|T098|LN|1524-8|LNC|glucose|glucose
C1551545|T098|MTH_LN|1524-8|LNC|glucose|glucose
C1551545|T098|OSN|1524-8|LNC|glucose|glucose
C1551545|T098|LC|1524-8|LNC|glucose|glucose
C1551546|T098|LN|1525-5|LNC|glucose|glucose
C1551546|T098|MTH_LN|1525-5|LNC|glucose|glucose
C1551546|T098|OSN|1525-5|LNC|glucose|glucose
C1551546|T098|LC|1525-5|LNC|glucose|glucose
C1551547|T098|LN|1526-3|LNC|glucose|glucose
C1551547|T098|MTH_LN|1526-3|LNC|glucose|glucose
C1551547|T098|OSN|1526-3|LNC|glucose|glucose
C1551547|T098|LC|1526-3|LNC|glucose|glucose
C1551548|T098|LN|1527-1|LNC|glucose|glucose
C1551548|T098|MTH_LN|1527-1|LNC|glucose|glucose
C1551548|T098|OSN|1527-1|LNC|glucose|glucose
C1551548|T098|LC|1527-1|LNC|glucose|glucose
C1551549|T098|MTH_LN|1528-9|LNC|glucose|glucose
C1551549|T098|LN|1528-9|LNC|glucose|glucose
C1551549|T098|OSN|1528-9|LNC|glucose|glucose
C1551549|T098|LC|1528-9|LNC|glucose|glucose
C1551551|T098|LN|1530-5|LNC|glucose|glucose
C1551551|T098|MTH_LN|1530-5|LNC|glucose|glucose
C1551551|T098|OSN|1530-5|LNC|glucose|glucose
C1551551|T098|LC|1530-5|LNC|glucose|glucose
C1551554|T098|LN|1533-9|LNC|glucose|glucose
C1551554|T098|MTH_LN|1533-9|LNC|glucose|glucose
C1551554|T098|OSN|1533-9|LNC|glucose|glucose
C1551554|T098|LC|1533-9|LNC|glucose|glucose
C1551555|T098|LN|1534-7|LNC|glucose|glucose
C1551555|T098|MTH_LN|1534-7|LNC|glucose|glucose
C1551555|T098|OSN|1534-7|LNC|glucose|glucose
C1551555|T098|LC|1534-7|LNC|glucose|glucose
C1551556|T098|LN|1535-4|LNC|glucose|glucose
C1551556|T098|MTH_LN|1535-4|LNC|glucose|glucose
C1551556|T098|OSN|1535-4|LNC|glucose|glucose
C1551556|T098|LC|1535-4|LNC|glucose|glucose
C1551557|T098|LN|1536-2|LNC|glucose|glucose
C1551557|T098|MTH_LN|1536-2|LNC|glucose|glucose
C1551557|T098|OSN|1536-2|LNC|glucose|glucose
C1551557|T098|LC|1536-2|LNC|glucose|glucose
C1551558|T098|LN|1537-0|LNC|glucose|glucose
C1551558|T098|MTH_LN|1537-0|LNC|glucose|glucose
C1551558|T098|OSN|1537-0|LNC|glucose|glucose
C1551558|T098|LC|1537-0|LNC|glucose|glucose
C1551560|T098|LN|1539-6|LNC|glucose|glucose
C1551560|T098|MTH_LN|1539-6|LNC|glucose|glucose
C1551560|T098|OSN|1539-6|LNC|glucose|glucose
C1551560|T098|LC|1539-6|LNC|glucose|glucose
C1551562|T098|LN|1543-8|LNC|glucose|glucose
C1551562|T098|MTH_LN|1543-8|LNC|glucose|glucose
C1551562|T098|OSN|1543-8|LNC|glucose|glucose
C1551562|T098|LC|1543-8|LNC|glucose|glucose
C1551564|T098|LN|1547-9|LNC|glucose|glucose
C1551564|T098|MTH_LN|1547-9|LNC|glucose|glucose
C1551564|T098|OSN|1547-9|LNC|glucose|glucose
C1551564|T098|LC|1547-9|LNC|glucose|glucose
C1551565|T098|LN|1549-5|LNC|glucose|glucose
C1551565|T098|MTH_LN|1549-5|LNC|glucose|glucose
C1551565|T098|OSN|1549-5|LNC|glucose|glucose
C1551565|T098|LC|1549-5|LNC|glucose|glucose
C1551566|T098|LN|1551-1|LNC|glucose|glucose
C1551566|T098|MTH_LN|1551-1|LNC|glucose|glucose
C1551566|T098|OSN|1551-1|LNC|glucose|glucose
C1551566|T098|LC|1551-1|LNC|glucose|glucose
C1551567|T098|LN|1552-9|LNC|glucose|glucose
C1551567|T098|MTH_LN|1552-9|LNC|glucose|glucose
C1551567|T098|OSN|1552-9|LNC|glucose|glucose
C1551567|T098|LC|1552-9|LNC|glucose|glucose
C1551568|T098|LN|1553-7|LNC|glucose|glucose
C1551568|T098|MTH_LN|1553-7|LNC|glucose|glucose
C1551568|T098|OSN|1553-7|LNC|glucose|glucose
C1551568|T098|LC|1553-7|LNC|glucose|glucose
C1551569|T098|LN|1554-5|LNC|glucose|glucose
C1551569|T098|MTH_LN|1554-5|LNC|glucose|glucose
C1551569|T098|OSN|1554-5|LNC|glucose|glucose
C1551569|T098|LC|1554-5|LNC|glucose|glucose
C1551571|T098|MTH_LN|1558-6|LNC|glucose|glucose
C1551571|T098|LN|1558-6|LNC|glucose|glucose
C1551571|T098|OSN|1558-6|LNC|glucose|glucose
C1551571|T098|LC|1558-6|LNC|glucose|glucose
C1551589|T098|LN|1588-3|LNC|luteinizing|luteinizing
C1551589|T098|OSN|1588-3|LNC|luteinizing|luteinizing
C1551589|T098|MTH_LN|1588-3|LNC|luteinizing|luteinizing
C1551589|T098|LC|1588-3|LNC|luteinizing|luteinizing
C1551589|T098|LN|1588-3|LNC|LH|LH
C1551589|T098|OSN|1588-3|LNC|LH|LH
C1551589|T098|MTH_LN|1588-3|LNC|LH|LH
C1551589|T098|LC|1588-3|LNC|LH|LH
C1551589|T098|LN|1588-3|LNC|luteinising|luteinising
C1551589|T098|OSN|1588-3|LNC|luteinising|luteinising
C1551589|T098|MTH_LN|1588-3|LNC|luteinising|luteinising
C1551589|T098|LC|1588-3|LNC|luteinising|luteinising
C1551593|T098|LN|1592-5|LNC|luteinizing|luteinizing
C1551593|T098|MTH_LN|1592-5|LNC|luteinizing|luteinizing
C1551593|T098|OSN|1592-5|LNC|luteinizing|luteinizing
C1551593|T098|LC|1592-5|LNC|luteinizing|luteinizing
C1551593|T098|LN|1592-5|LNC|LH|LH
C1551593|T098|MTH_LN|1592-5|LNC|LH|LH
C1551593|T098|OSN|1592-5|LNC|LH|LH
C1551593|T098|LC|1592-5|LNC|LH|LH
C1551593|T098|LN|1592-5|LNC|luteinising|luteinising
C1551593|T098|MTH_LN|1592-5|LNC|luteinising|luteinising
C1551593|T098|OSN|1592-5|LNC|luteinising|luteinising
C1551593|T098|LC|1592-5|LNC|luteinising|luteinising
C1551595|T098|LN|1594-1|LNC|luteinizing|luteinizing
C1551595|T098|MTH_LN|1594-1|LNC|luteinizing|luteinizing
C1551595|T098|OSN|1594-1|LNC|luteinizing|luteinizing
C1551595|T098|LC|1594-1|LNC|luteinizing|luteinizing
C1551595|T098|LN|1594-1|LNC|LH|LH
C1551595|T098|MTH_LN|1594-1|LNC|LH|LH
C1551595|T098|OSN|1594-1|LNC|LH|LH
C1551595|T098|LC|1594-1|LNC|LH|LH
C1551595|T098|LN|1594-1|LNC|luteinising|luteinising
C1551595|T098|MTH_LN|1594-1|LNC|luteinising|luteinising
C1551595|T098|OSN|1594-1|LNC|luteinising|luteinising
C1551595|T098|LC|1594-1|LNC|luteinising|luteinising
C1551597|T098|LN|1596-6|LNC|luteinizing|luteinizing
C1551597|T098|MTH_LN|1596-6|LNC|luteinizing|luteinizing
C1551597|T098|OSN|1596-6|LNC|luteinizing|luteinizing
C1551597|T098|LC|1596-6|LNC|luteinizing|luteinizing
C1551597|T098|LN|1596-6|LNC|LH|LH
C1551597|T098|MTH_LN|1596-6|LNC|LH|LH
C1551597|T098|OSN|1596-6|LNC|LH|LH
C1551597|T098|LC|1596-6|LNC|LH|LH
C1551597|T098|LN|1596-6|LNC|luteinising|luteinising
C1551597|T098|MTH_LN|1596-6|LNC|luteinising|luteinising
C1551597|T098|OSN|1596-6|LNC|luteinising|luteinising
C1551597|T098|LC|1596-6|LNC|luteinising|luteinising
C1551600|T098|LN|1599-0|LNC|luteinizing|luteinizing
C1551600|T098|MTH_LN|1599-0|LNC|luteinizing|luteinizing
C1551600|T098|OSN|1599-0|LNC|luteinizing|luteinizing
C1551600|T098|LC|1599-0|LNC|luteinizing|luteinizing
C1551600|T098|LN|1599-0|LNC|LH|LH
C1551600|T098|MTH_LN|1599-0|LNC|LH|LH
C1551600|T098|OSN|1599-0|LNC|LH|LH
C1551600|T098|LC|1599-0|LNC|LH|LH
C1551600|T098|LN|1599-0|LNC|luteinising|luteinising
C1551600|T098|MTH_LN|1599-0|LNC|luteinising|luteinising
C1551600|T098|OSN|1599-0|LNC|luteinising|luteinising
C1551600|T098|LC|1599-0|LNC|luteinising|luteinising
C1551601|T098|LN|1600-6|LNC|luteinizing|luteinizing
C1551601|T098|MTH_LN|1600-6|LNC|luteinizing|luteinizing
C1551601|T098|OSN|1600-6|LNC|luteinizing|luteinizing
C1551601|T098|LC|1600-6|LNC|luteinizing|luteinizing
C1551601|T098|LN|1600-6|LNC|LH|LH
C1551601|T098|MTH_LN|1600-6|LNC|LH|LH
C1551601|T098|OSN|1600-6|LNC|LH|LH
C1551601|T098|LC|1600-6|LNC|LH|LH
C1551601|T098|LN|1600-6|LNC|luteinising|luteinising
C1551601|T098|MTH_LN|1600-6|LNC|luteinising|luteinising
C1551601|T098|OSN|1600-6|LNC|luteinising|luteinising
C1551601|T098|LC|1600-6|LNC|luteinising|luteinising
C1551642|T098|LN|1649-3|LNC|calcium|calcium
C1551642|T098|MTH_LN|1649-3|LNC|calcium|calcium
C1551642|T098|LC|1649-3|LNC|calcium|calcium
C1551642|T098|OSN|1649-3|LNC|calcium|calcium
C1551654|T098|LN|1668-3|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C1551654|T098|MTH_LN|1668-3|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C1551654|T098|OSN|1668-3|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C1551654|T098|LC|1668-3|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C1551654|T098|LN|1668-3|LNC|17-OHP|17-OHP
C1551654|T098|MTH_LN|1668-3|LNC|17-OHP|17-OHP
C1551654|T098|OSN|1668-3|LNC|17-OHP|17-OHP
C1551654|T098|LC|1668-3|LNC|17-OHP|17-OHP
C1551660|T098|LN|1679-0|LNC|vitamin D metabolism|vitamin D metabolism
C1551660|T098|MTH_LN|1679-0|LNC|vitamin D metabolism|vitamin D metabolism
C1551660|T098|OSN|1679-0|LNC|vitamin D metabolism|vitamin D metabolism
C1551660|T098|LC|1679-0|LNC|vitamin D metabolism|vitamin D metabolism
C1551660|T098|LN|1679-0|LNC|calcifediol|calcifediol
C1551660|T098|MTH_LN|1679-0|LNC|calcifediol|calcifediol
C1551660|T098|OSN|1679-0|LNC|calcifediol|calcifediol
C1551660|T098|LC|1679-0|LNC|calcifediol|calcifediol
C1551660|T098|LN|1679-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1551660|T098|MTH_LN|1679-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1551660|T098|OSN|1679-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1551660|T098|LC|1679-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1551660|T098|LN|1679-0|LNC|calcidiol|calcidiol
C1551660|T098|MTH_LN|1679-0|LNC|calcidiol|calcidiol
C1551660|T098|OSN|1679-0|LNC|calcidiol|calcidiol
C1551660|T098|LC|1679-0|LNC|calcidiol|calcidiol
C1551660|T098|LN|1679-0|LNC|calcitriol|calcitriol
C1551660|T098|MTH_LN|1679-0|LNC|calcitriol|calcitriol
C1551660|T098|OSN|1679-0|LNC|calcitriol|calcitriol
C1551660|T098|LC|1679-0|LNC|calcitriol|calcitriol
C1551660|T098|LN|1679-0|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C1551660|T098|MTH_LN|1679-0|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C1551660|T098|OSN|1679-0|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C1551660|T098|LC|1679-0|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C1551660|T098|LN|1679-0|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C1551660|T098|MTH_LN|1679-0|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C1551660|T098|OSN|1679-0|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C1551660|T098|LC|1679-0|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C1551666|T098|LN|1688-1|LNC|vitamin b6|vitamin b6
C1551666|T098|MTH_LN|1688-1|LNC|vitamin b6|vitamin b6
C1551666|T098|OSN|1688-1|LNC|vitamin b6|vitamin b6
C1551666|T098|LC|1688-1|LNC|vitamin b6|vitamin b6
C1551666|T098|LN|1688-1|LNC|vitamin B metabolism|vitamin B metabolism
C1551666|T098|MTH_LN|1688-1|LNC|vitamin B metabolism|vitamin B metabolism
C1551666|T098|OSN|1688-1|LNC|vitamin B metabolism|vitamin B metabolism
C1551666|T098|LC|1688-1|LNC|vitamin B metabolism|vitamin B metabolism
C1551666|T098|LN|1688-1|LNC|B-vitamin metabolism|B-vitamin metabolism
C1551666|T098|MTH_LN|1688-1|LNC|B-vitamin metabolism|B-vitamin metabolism
C1551666|T098|OSN|1688-1|LNC|B-vitamin metabolism|B-vitamin metabolism
C1551666|T098|LC|1688-1|LNC|B-vitamin metabolism|B-vitamin metabolism
C1551684|T098|LN|1717-8|LNC|acylcarnitine|acylcarnitine
C1551684|T098|LC|1717-8|LNC|acylcarnitine|acylcarnitine
C1551684|T098|MTH_LN|1717-8|LNC|acylcarnitine|acylcarnitine
C1551684|T098|OSN|1717-8|LNC|acylcarnitine|acylcarnitine
C1551688|T098|LN|1722-8|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C1551688|T098|MTH_LN|1722-8|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C1551688|T098|OSN|1722-8|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C1551688|T098|LC|1722-8|LNC|erythrocyte enzyme activity|erythrocyte enzyme activity
C1551688|T098|LN|1722-8|LNC|red cell adenosine deaminase activity|red cell adenosine deaminase activity
C1551688|T098|MTH_LN|1722-8|LNC|red cell adenosine deaminase activity|red cell adenosine deaminase activity
C1551688|T098|OSN|1722-8|LNC|red cell adenosine deaminase activity|red cell adenosine deaminase activity
C1551688|T098|LC|1722-8|LNC|red cell adenosine deaminase activity|red cell adenosine deaminase activity
C1551706|T098|LN|1746-7|LNC|CSF albumin|CSF albumin
C1551706|T098|MTH_LN|1746-7|LNC|CSF albumin|CSF albumin
C1551706|T098|OSN|1746-7|LNC|CSF albumin|CSF albumin
C1551706|T098|LC|1746-7|LNC|CSF albumin|CSF albumin
C1551706|T098|LN|1746-7|LNC|CSF albumin is belowlower limitnormal.|CSF albumin is belowlower limitnormal.
C1551706|T098|MTH_LN|1746-7|LNC|CSF albumin is belowlower limitnormal.|CSF albumin is belowlower limitnormal.
C1551706|T098|OSN|1746-7|LNC|CSF albumin is belowlower limitnormal.|CSF albumin is belowlower limitnormal.
C1551706|T098|LC|1746-7|LNC|CSF albumin is belowlower limitnormal.|CSF albumin is belowlower limitnormal.
C1551706|T098|LN|1746-7|LNC|CSF protein|CSF protein
C1551706|T098|MTH_LN|1746-7|LNC|CSF protein|CSF protein
C1551706|T098|OSN|1746-7|LNC|CSF protein|CSF protein
C1551706|T098|LC|1746-7|LNC|CSF protein|CSF protein
C1551711|T098|LN|1751-7|LNC|albumin|albumin
C1551711|T098|MTH_LN|1751-7|LNC|albumin|albumin
C1551711|T098|OSN|1751-7|LNC|albumin|albumin
C1551711|T098|LC|1751-7|LNC|albumin|albumin
C1551719|T098|LN|1759-0|LNC|albumin|albumin
C1551719|T098|OSN|1759-0|LNC|albumin|albumin
C1551719|T098|MTH_LN|1759-0|LNC|albumin|albumin
C1551719|T098|LC|1759-0|LNC|albumin|albumin
C1551721|T098|LN|1761-6|LNC|aldolase|aldolase
C1551721|T098|MTH_LN|1761-6|LNC|aldolase|aldolase
C1551721|T098|OSN|1761-6|LNC|aldolase|aldolase
C1551721|T098|LC|1761-6|LNC|aldolase|aldolase
C1551723|T098|LN|1763-2|LNC|aldosterone|aldosterone
C1551723|T098|MTH_LN|1763-2|LNC|aldosterone|aldosterone
C1551723|T098|OSN|1763-2|LNC|aldosterone|aldosterone
C1551723|T098|LC|1763-2|LNC|aldosterone|aldosterone
C1551737|T098|LN|1777-2|LNC|Alkaline phosphatase|Alkaline phosphatase
C1551737|T098|MTH_LN|1777-2|LNC|Alkaline phosphatase|Alkaline phosphatase
C1551737|T098|OSN|1777-2|LNC|Alkaline phosphatase|Alkaline phosphatase
C1551737|T098|LC|1777-2|LNC|Alkaline phosphatase|Alkaline phosphatase
C1551737|T098|LN|1777-2|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C1551737|T098|MTH_LN|1777-2|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C1551737|T098|OSN|1777-2|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C1551737|T098|LC|1777-2|LNC|alkaline phosphatasebone origin|alkaline phosphatasebone origin
C1551737|T098|LN|1777-2|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C1551737|T098|MTH_LN|1777-2|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C1551737|T098|OSN|1777-2|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C1551737|T098|LC|1777-2|LNC|bone-specific alkaline phosphatase|bone-specific alkaline phosphatase
C1551737|T098|LN|1777-2|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C1551737|T098|MTH_LN|1777-2|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C1551737|T098|OSN|1777-2|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C1551737|T098|LC|1777-2|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C1551738|T098|LN|1778-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C1551738|T098|MTH_LN|1778-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C1551738|T098|OSN|1778-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C1551738|T098|LC|1778-0|LNC|Alkaline phosphatase|Alkaline phosphatase
C1551738|T098|LN|1778-0|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C1551738|T098|MTH_LN|1778-0|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C1551738|T098|OSN|1778-0|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C1551738|T098|LC|1778-0|LNC|intestinal alkaline phosphatase|intestinal alkaline phosphatase
C1551738|T098|LN|1778-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C1551738|T098|MTH_LN|1778-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C1551738|T098|OSN|1778-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C1551738|T098|LC|1778-0|LNC|alkaline phosphatase activity|alkaline phosphatase activity
C1551790|T098|LN|1834-1|LNC|alpha-fetoprotein|alpha-fetoprotein
C1551790|T098|OSN|1834-1|LNC|alpha-fetoprotein|alpha-fetoprotein
C1551790|T098|MTH_LN|1834-1|LNC|alpha-fetoprotein|alpha-fetoprotein
C1551790|T098|LC|1834-1|LNC|alpha-fetoprotein|alpha-fetoprotein
C1551790|T098|LN|1834-1|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C1551790|T098|OSN|1834-1|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C1551790|T098|MTH_LN|1834-1|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C1551790|T098|LC|1834-1|LNC|Serum alpha-fetoprotein|Serum alpha-fetoprotein
C1551790|T098|LN|1834-1|LNC|alpha fetoprotein|alpha fetoprotein
C1551790|T098|OSN|1834-1|LNC|alpha fetoprotein|alpha fetoprotein
C1551790|T098|MTH_LN|1834-1|LNC|alpha fetoprotein|alpha fetoprotein
C1551790|T098|LC|1834-1|LNC|alpha fetoprotein|alpha fetoprotein
C1551799|T098|LN|1848-1|LNC|testosterone|testosterone
C1551799|T098|MTH_LN|1848-1|LNC|testosterone|testosterone
C1551799|T098|OSN|1848-1|LNC|testosterone|testosterone
C1551799|T098|LC|1848-1|LNC|testosterone|testosterone
C1551799|T098|LN|1848-1|LNC|androgen|androgen
C1551799|T098|MTH_LN|1848-1|LNC|androgen|androgen
C1551799|T098|OSN|1848-1|LNC|androgen|androgen
C1551799|T098|LC|1848-1|LNC|androgen|androgen
C1551805|T098|LN|1854-9|LNC|androstenedione|androstenedione
C1551805|T098|MTH_LN|1854-9|LNC|androstenedione|androstenedione
C1551805|T098|OSN|1854-9|LNC|androstenedione|androstenedione
C1551805|T098|LC|1854-9|LNC|androstenedione|androstenedione
C1551805|T098|LN|1854-9|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C1551805|T098|MTH_LN|1854-9|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C1551805|T098|OSN|1854-9|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C1551805|T098|LC|1854-9|LNC|dehydroepiandrosterone|dehydroepiandrosterone
C1551805|T098|LN|1854-9|LNC|androstenolone|androstenolone
C1551805|T098|MTH_LN|1854-9|LNC|androstenolone|androstenolone
C1551805|T098|OSN|1854-9|LNC|androstenolone|androstenolone
C1551805|T098|LC|1854-9|LNC|androstenolone|androstenolone
C1551805|T098|LN|1854-9|LNC|DHEA|DHEA
C1551805|T098|MTH_LN|1854-9|LNC|DHEA|DHEA
C1551805|T098|OSN|1854-9|LNC|DHEA|DHEA
C1551805|T098|LC|1854-9|LNC|DHEA|DHEA
C1551835|T098|MTH_LN|1884-6|LNC|apolipoprotein|apolipoprotein
C1551835|T098|LN|1884-6|LNC|apolipoprotein|apolipoprotein
C1551835|T098|OSN|1884-6|LNC|apolipoprotein|apolipoprotein
C1551835|T098|LC|1884-6|LNC|apolipoprotein|apolipoprotein
C1551835|T098|MTH_LN|1884-6|LNC|apolipoprotein B|apolipoprotein B
C1551835|T098|LN|1884-6|LNC|apolipoprotein B|apolipoprotein B
C1551835|T098|OSN|1884-6|LNC|apolipoprotein B|apolipoprotein B
C1551835|T098|LC|1884-6|LNC|apolipoprotein B|apolipoprotein B
C1551835|T098|MTH_LN|1884-6|LNC|ApoB|ApoB
C1551835|T098|LN|1884-6|LNC|ApoB|ApoB
C1551835|T098|OSN|1884-6|LNC|ApoB|ApoB
C1551835|T098|LC|1884-6|LNC|ApoB|ApoB
C1551843|T098|LN|1893-7|LNC|arginine metabolism|arginine metabolism
C1551843|T098|MTH_LN|1893-7|LNC|arginine metabolism|arginine metabolism
C1551843|T098|OSN|1893-7|LNC|arginine metabolism|arginine metabolism
C1551843|T098|LC|1893-7|LNC|arginine metabolism|arginine metabolism
C1551843|T098|LN|1893-7|LNC|arginine|arginine
C1551843|T098|MTH_LN|1893-7|LNC|arginine|arginine
C1551843|T098|OSN|1893-7|LNC|arginine|arginine
C1551843|T098|LC|1893-7|LNC|arginine|arginine
C1551844|T098|LN|1894-5|LNC|arginine|arginine
C1551844|T098|MTH_LN|1894-5|LNC|arginine|arginine
C1551844|T098|OSN|1894-5|LNC|arginine|arginine
C1551844|T098|LC|1894-5|LNC|arginine|arginine
C1553258|T098|LN|1952-1|LNC|beta-2-microglobulin|beta-2-microglobulin
C1553258|T098|OSN|1952-1|LNC|beta-2-microglobulin|beta-2-microglobulin
C1553258|T098|LC|1952-1|LNC|beta-2-microglobulin|beta-2-microglobulin
C1553258|T098|MTH_LN|1952-1|LNC|beta-2-microglobulin|beta-2-microglobulin
C1553258|T098|LN|1952-1|LNC|B2M|B2M
C1553258|T098|OSN|1952-1|LNC|B2M|B2M
C1553258|T098|LC|1952-1|LNC|B2M|B2M
C1553258|T098|MTH_LN|1952-1|LNC|B2M|B2M
C1553258|T098|LN|1952-1|LNC|beta2m|beta2m
C1553258|T098|OSN|1952-1|LNC|beta2m|beta2m
C1553258|T098|LC|1952-1|LNC|beta2m|beta2m
C1553258|T098|MTH_LN|1952-1|LNC|beta2m|beta2m
C1553258|T098|LN|1952-1|LNC|beta2 microglobulin|beta2 microglobulin
C1553258|T098|OSN|1952-1|LNC|beta2 microglobulin|beta2 microglobulin
C1553258|T098|LC|1952-1|LNC|beta2 microglobulin|beta2 microglobulin
C1553258|T098|MTH_LN|1952-1|LNC|beta2 microglobulin|beta2 microglobulin
C1553258|T098|LN|1952-1|LNC|beta2-m|beta2-m
C1553258|T098|OSN|1952-1|LNC|beta2-m|beta2-m
C1553258|T098|LC|1952-1|LNC|beta2-m|beta2-m
C1553258|T098|MTH_LN|1952-1|LNC|beta2-m|beta2-m
C1553270|T098|LN|1964-6|LNC|bicarbonate|bicarbonate
C1553270|T098|MTH_LN|1964-6|LNC|bicarbonate|bicarbonate
C1553270|T098|OSN|1964-6|LNC|bicarbonate|bicarbonate
C1553270|T098|LC|1964-6|LNC|bicarbonate|bicarbonate
C1553271|T098|LN|1968-7|LNC|bilirubin|bilirubin
C1553271|T098|MTH_LN|1968-7|LNC|bilirubin|bilirubin
C1553271|T098|OSN|1968-7|LNC|bilirubin|bilirubin
C1553271|T098|LC|1968-7|LNC|bilirubin|bilirubin
C1553271|T098|LN|1968-7|LNC|metabolism/homeostasis|metabolism/homeostasis
C1553271|T098|MTH_LN|1968-7|LNC|metabolism/homeostasis|metabolism/homeostasis
C1553271|T098|OSN|1968-7|LNC|metabolism/homeostasis|metabolism/homeostasis
C1553271|T098|LC|1968-7|LNC|metabolism/homeostasis|metabolism/homeostasis
C1553271|T098|LN|1968-7|LNC|Metabolism|Metabolism
C1553271|T098|MTH_LN|1968-7|LNC|Metabolism|Metabolism
C1553271|T098|OSN|1968-7|LNC|Metabolism|Metabolism
C1553271|T098|LC|1968-7|LNC|Metabolism|Metabolism
C1553271|T098|LN|1968-7|LNC|Laboratory|Laboratory
C1553271|T098|MTH_LN|1968-7|LNC|Laboratory|Laboratory
C1553271|T098|OSN|1968-7|LNC|Laboratory|Laboratory
C1553271|T098|LC|1968-7|LNC|Laboratory|Laboratory
C1553276|T098|LN|1975-2|LNC|bilirubin|bilirubin
C1553276|T098|MTH_LN|1975-2|LNC|bilirubin|bilirubin
C1553276|T098|OSN|1975-2|LNC|bilirubin|bilirubin
C1553276|T098|LC|1975-2|LNC|bilirubin|bilirubin
C1553276|T098|LN|1975-2|LNC|total bilirubin|total bilirubin
C1553276|T098|MTH_LN|1975-2|LNC|total bilirubin|total bilirubin
C1553276|T098|OSN|1975-2|LNC|total bilirubin|total bilirubin
C1553276|T098|LC|1975-2|LNC|total bilirubin|total bilirubin
C1553276|T098|LN|1975-2|LNC|bili total|bili total
C1553276|T098|MTH_LN|1975-2|LNC|bili total|bili total
C1553276|T098|OSN|1975-2|LNC|bili total|bili total
C1553276|T098|LC|1975-2|LNC|bili total|bili total
C1553286|T098|MTH_LN|1986-9|LNC|C-peptide|C-peptide
C1553286|T098|LN|1986-9|LNC|C-peptide|C-peptide
C1553286|T098|OSN|1986-9|LNC|C-peptide|C-peptide
C1553286|T098|LC|1986-9|LNC|C-peptide|C-peptide
C1553286|T098|MTH_LN|1986-9|LNC|C peptide|C peptide
C1553286|T098|LN|1986-9|LNC|C peptide|C peptide
C1553286|T098|OSN|1986-9|LNC|C peptide|C peptide
C1553286|T098|LC|1986-9|LNC|C peptide|C peptide
C1553288|T098|LN|1988-5|LNC|CRP|CRP
C1553288|T098|MTH_LN|1988-5|LNC|CRP|CRP
C1553288|T098|OSN|1988-5|LNC|CRP|CRP
C1553288|T098|LC|1988-5|LNC|CRP|CRP
C1553288|T098|LN|1988-5|LNC|C-reactive protein|C-reactive protein
C1553288|T098|MTH_LN|1988-5|LNC|C-reactive protein|C-reactive protein
C1553288|T098|OSN|1988-5|LNC|C-reactive protein|C-reactive protein
C1553288|T098|LC|1988-5|LNC|C-reactive protein|C-reactive protein
C1553288|T098|LN|1988-5|LNC|C-peptide|C-peptide
C1553288|T098|MTH_LN|1988-5|LNC|C-peptide|C-peptide
C1553288|T098|OSN|1988-5|LNC|C-peptide|C-peptide
C1553288|T098|LC|1988-5|LNC|C-peptide|C-peptide
C1553288|T098|LN|1988-5|LNC|C peptide|C peptide
C1553288|T098|MTH_LN|1988-5|LNC|C peptide|C peptide
C1553288|T098|OSN|1988-5|LNC|C peptide|C peptide
C1553288|T098|LC|1988-5|LNC|C peptide|C peptide
C1553292|T098|LN|1994-3|LNC|calcium|calcium
C1553292|T098|MTH_LN|1994-3|LNC|calcium|calcium
C1553292|T098|OSN|1994-3|LNC|calcium|calcium
C1553292|T098|LC|1994-3|LNC|calcium|calcium
C1553292|T098|LN|1994-3|LNC|calcium homeostasis|calcium homeostasis
C1553292|T098|MTH_LN|1994-3|LNC|calcium homeostasis|calcium homeostasis
C1553292|T098|OSN|1994-3|LNC|calcium homeostasis|calcium homeostasis
C1553292|T098|LC|1994-3|LNC|calcium homeostasis|calcium homeostasis
C1553293|T098|LN|1995-0|LNC|calcium|calcium
C1553293|T098|MTH_LN|1995-0|LNC|calcium|calcium
C1553293|T098|OSN|1995-0|LNC|calcium|calcium
C1553293|T098|LC|1995-0|LNC|calcium|calcium
C1553293|T098|LN|1995-0|LNC|calcium homeostasis|calcium homeostasis
C1553293|T098|MTH_LN|1995-0|LNC|calcium homeostasis|calcium homeostasis
C1553293|T098|OSN|1995-0|LNC|calcium homeostasis|calcium homeostasis
C1553293|T098|LC|1995-0|LNC|calcium homeostasis|calcium homeostasis
C1553294|T098|LN|1996-8|LNC|calcium|calcium
C1553294|T098|MTH_LN|1996-8|LNC|calcium|calcium
C1553294|T098|OSN|1996-8|LNC|calcium|calcium
C1553294|T098|LC|1996-8|LNC|calcium|calcium
C1553294|T098|LN|1996-8|LNC|calcium homeostasis|calcium homeostasis
C1553294|T098|MTH_LN|1996-8|LNC|calcium homeostasis|calcium homeostasis
C1553294|T098|OSN|1996-8|LNC|calcium homeostasis|calcium homeostasis
C1553294|T098|LC|1996-8|LNC|calcium homeostasis|calcium homeostasis
C1553298|T098|LN|2000-8|LNC|calcium|calcium
C1553298|T098|MTH_LN|2000-8|LNC|calcium|calcium
C1553298|T098|OSN|2000-8|LNC|calcium|calcium
C1553298|T098|LC|2000-8|LNC|calcium|calcium
C1553298|T098|LN|2000-8|LNC|calcium homeostasis|calcium homeostasis
C1553298|T098|MTH_LN|2000-8|LNC|calcium homeostasis|calcium homeostasis
C1553298|T098|OSN|2000-8|LNC|calcium homeostasis|calcium homeostasis
C1553298|T098|LC|2000-8|LNC|calcium homeostasis|calcium homeostasis
C1553314|T098|LN|2019-8|LNC|carbon dioxide|carbon dioxide
C1553314|T098|MTH_LN|2019-8|LNC|carbon dioxide|carbon dioxide
C1553314|T098|LC|2019-8|LNC|carbon dioxide|carbon dioxide
C1553314|T098|OSN|2019-8|LNC|carbon dioxide|carbon dioxide
C1553315|T098|LN|2020-6|LNC|carbon dioxide|carbon dioxide
C1553315|T098|MTH_LN|2020-6|LNC|carbon dioxide|carbon dioxide
C1553315|T098|LC|2020-6|LNC|carbon dioxide|carbon dioxide
C1553315|T098|OSN|2020-6|LNC|carbon dioxide|carbon dioxide
C1553316|T098|LN|2021-4|LNC|carbon dioxide|carbon dioxide
C1553316|T098|MTH_LN|2021-4|LNC|carbon dioxide|carbon dioxide
C1553316|T098|OSN|2021-4|LNC|carbon dioxide|carbon dioxide
C1553316|T098|LC|2021-4|LNC|carbon dioxide|carbon dioxide
C1553338|T098|LN|2069-3|LNC|chloride|chloride
C1553338|T098|MTH_LN|2069-3|LNC|chloride|chloride
C1553338|T098|OSN|2069-3|LNC|chloride|chloride
C1553338|T098|LC|2069-3|LNC|chloride|chloride
C1553338|T098|LN|2069-3|LNC|chloride homeostasis|chloride homeostasis
C1553338|T098|MTH_LN|2069-3|LNC|chloride homeostasis|chloride homeostasis
C1553338|T098|OSN|2069-3|LNC|chloride homeostasis|chloride homeostasis
C1553338|T098|LC|2069-3|LNC|chloride homeostasis|chloride homeostasis
C1553342|T098|OLC|2086-7|LNC|HDL cholesterol|HDL cholesterol
C1553342|T098|MTH_LO|2086-7|LNC|HDL cholesterol|HDL cholesterol
C1553342|T098|LO|2086-7|LNC|HDL cholesterol|HDL cholesterol
C1553342|T098|OOSN|2086-7|LNC|HDL cholesterol|HDL cholesterol
C1553342|T098|OLC|2086-7|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1553342|T098|MTH_LO|2086-7|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1553342|T098|LO|2086-7|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1553342|T098|OOSN|2086-7|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1553342|T098|OLC|2086-7|LNC|HDL-cholesterol|HDL-cholesterol
C1553342|T098|MTH_LO|2086-7|LNC|HDL-cholesterol|HDL-cholesterol
C1553342|T098|LO|2086-7|LNC|HDL-cholesterol|HDL-cholesterol
C1553342|T098|OOSN|2086-7|LNC|HDL-cholesterol|HDL-cholesterol
C1553342|T098|OLC|2086-7|LNC|high-density lipoprotein|high-density lipoprotein
C1553342|T098|MTH_LO|2086-7|LNC|high-density lipoprotein|high-density lipoprotein
C1553342|T098|LO|2086-7|LNC|high-density lipoprotein|high-density lipoprotein
C1553342|T098|OOSN|2086-7|LNC|high-density lipoprotein|high-density lipoprotein
C1553342|T098|OLC|2086-7|LNC|HDL|HDL
C1553342|T098|MTH_LO|2086-7|LNC|HDL|HDL
C1553342|T098|LO|2086-7|LNC|HDL|HDL
C1553342|T098|OOSN|2086-7|LNC|HDL|HDL
C1553344|T098|MTH_LN|2089-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1553344|T098|LN|2089-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1553344|T098|OSN|2089-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1553344|T098|LC|2089-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1553344|T098|MTH_LN|2089-1|LNC|LDL|LDL
C1553344|T098|LN|2089-1|LNC|LDL|LDL
C1553344|T098|OSN|2089-1|LNC|LDL|LDL
C1553344|T098|LC|2089-1|LNC|LDL|LDL
C1553344|T098|MTH_LN|2089-1|LNC|LDL cholesterol|LDL cholesterol
C1553344|T098|LN|2089-1|LNC|LDL cholesterol|LDL cholesterol
C1553344|T098|OSN|2089-1|LNC|LDL cholesterol|LDL cholesterol
C1553344|T098|LC|2089-1|LNC|LDL cholesterol|LDL cholesterol
C1553344|T098|MTH_LN|2089-1|LNC|low-density lipoprotein|low-density lipoprotein
C1553344|T098|LN|2089-1|LNC|low-density lipoprotein|low-density lipoprotein
C1553344|T098|OSN|2089-1|LNC|low-density lipoprotein|low-density lipoprotein
C1553344|T098|LC|2089-1|LNC|low-density lipoprotein|low-density lipoprotein
C1553344|T098|MTH_LN|2089-1|LNC|beta-lipoproteins|beta-lipoproteins
C1553344|T098|LN|2089-1|LNC|beta-lipoproteins|beta-lipoproteins
C1553344|T098|OSN|2089-1|LNC|beta-lipoproteins|beta-lipoproteins
C1553344|T098|LC|2089-1|LNC|beta-lipoproteins|beta-lipoproteins
C1553344|T098|MTH_LN|2089-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1553344|T098|LN|2089-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1553344|T098|OSN|2089-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1553344|T098|LC|2089-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1553344|T098|MTH_LN|2089-1|LNC|LDL-C|LDL-C
C1553344|T098|LN|2089-1|LNC|LDL-C|LDL-C
C1553344|T098|OSN|2089-1|LNC|LDL-C|LDL-C
C1553344|T098|LC|2089-1|LNC|LDL-C|LDL-C
C1553346|T098|MTH_LN|2093-3|LNC|cholesterol|cholesterol
C1553346|T098|LN|2093-3|LNC|cholesterol|cholesterol
C1553346|T098|OSN|2093-3|LNC|cholesterol|cholesterol
C1553346|T098|LC|2093-3|LNC|cholesterol|cholesterol
C1553346|T098|MTH_LN|2093-3|LNC|total cholesterol|total cholesterol
C1553346|T098|LN|2093-3|LNC|total cholesterol|total cholesterol
C1553346|T098|OSN|2093-3|LNC|total cholesterol|total cholesterol
C1553346|T098|LC|2093-3|LNC|total cholesterol|total cholesterol
C1553346|T098|MTH_LN|2093-3|LNC|cholesterol metabolism|cholesterol metabolism
C1553346|T098|LN|2093-3|LNC|cholesterol metabolism|cholesterol metabolism
C1553346|T098|OSN|2093-3|LNC|cholesterol metabolism|cholesterol metabolism
C1553346|T098|LC|2093-3|LNC|cholesterol metabolism|cholesterol metabolism
C1553351|T098|LC|2500-7|LNC|total iron binding capacity|total iron binding capacity
C1553351|T098|MTH_LN|2500-7|LNC|total iron binding capacity|total iron binding capacity
C1553351|T098|LN|2500-7|LNC|total iron binding capacity|total iron binding capacity
C1553351|T098|OSN|2500-7|LNC|total iron binding capacity|total iron binding capacity
C1553351|T098|LC|2500-7|LNC|iron homeostasis|iron homeostasis
C1553351|T098|MTH_LN|2500-7|LNC|iron homeostasis|iron homeostasis
C1553351|T098|LN|2500-7|LNC|iron homeostasis|iron homeostasis
C1553351|T098|OSN|2500-7|LNC|iron homeostasis|iron homeostasis
C1553353|T098|LN|2118-8|LNC|maternal chorionic gonadotropin|maternal chorionic gonadotropin
C1553353|T098|MTH_LN|2118-8|LNC|maternal chorionic gonadotropin|maternal chorionic gonadotropin
C1553353|T098|LC|2118-8|LNC|maternal chorionic gonadotropin|maternal chorionic gonadotropin
C1553353|T098|OSN|2118-8|LNC|maternal chorionic gonadotropin|maternal chorionic gonadotropin
C1553353|T098|LN|2118-8|LNC|maternal hCG|maternal hCG
C1553353|T098|MTH_LN|2118-8|LNC|maternal hCG|maternal hCG
C1553353|T098|LC|2118-8|LNC|maternal hCG|maternal hCG
C1553353|T098|OSN|2118-8|LNC|maternal hCG|maternal hCG
C1553353|T098|LN|2118-8|LNC|maternal screening|maternal screening
C1553353|T098|MTH_LN|2118-8|LNC|maternal screening|maternal screening
C1553353|T098|LC|2118-8|LNC|maternal screening|maternal screening
C1553353|T098|OSN|2118-8|LNC|maternal screening|maternal screening
C1553360|T098|LN|2139-4|LNC|corticosterone|corticosterone
C1553360|T098|MTH_LN|2139-4|LNC|corticosterone|corticosterone
C1553360|T098|LC|2139-4|LNC|corticosterone|corticosterone
C1553360|T098|OSN|2139-4|LNC|corticosterone|corticosterone
C1553362|T098|LC|2141-0|LNC|ACTH|ACTH
C1553362|T098|MTH_LN|2141-0|LNC|ACTH|ACTH
C1553362|T098|LN|2141-0|LNC|ACTH|ACTH
C1553362|T098|OSN|2141-0|LNC|ACTH|ACTH
C1553362|T098|LC|2141-0|LNC|corticotropin|corticotropin
C1553362|T098|MTH_LN|2141-0|LNC|corticotropin|corticotropin
C1553362|T098|LN|2141-0|LNC|corticotropin|corticotropin
C1553362|T098|OSN|2141-0|LNC|corticotropin|corticotropin
C1553362|T098|LC|2141-0|LNC|adrenocorticotropin|adrenocorticotropin
C1553362|T098|MTH_LN|2141-0|LNC|adrenocorticotropin|adrenocorticotropin
C1553362|T098|LN|2141-0|LNC|adrenocorticotropin|adrenocorticotropin
C1553362|T098|OSN|2141-0|LNC|adrenocorticotropin|adrenocorticotropin
C1553364|T098|LN|2143-6|LNC|cortisol|cortisol
C1553364|T098|MTH_LN|2143-6|LNC|cortisol|cortisol
C1553364|T098|OSN|2143-6|LNC|cortisol|cortisol
C1553364|T098|LC|2143-6|LNC|cortisol|cortisol
C1553364|T098|LN|2143-6|LNC|cortisol low|cortisol low
C1553364|T098|MTH_LN|2143-6|LNC|cortisol low|cortisol low
C1553364|T098|OSN|2143-6|LNC|cortisol low|cortisol low
C1553364|T098|LC|2143-6|LNC|cortisol low|cortisol low
C1553364|T098|LN|2143-6|LNC|to undetectable cortisol|to undetectable cortisol
C1553364|T098|MTH_LN|2143-6|LNC|to undetectable cortisol|to undetectable cortisol
C1553364|T098|OSN|2143-6|LNC|to undetectable cortisol|to undetectable cortisol
C1553364|T098|LC|2143-6|LNC|to undetectable cortisol|to undetectable cortisol
C1556094|T098|LN|2039-6|LNC|carcinoembryonic antigen|carcinoembryonic antigen
C1556094|T098|MTH_LN|2039-6|LNC|carcinoembryonic antigen|carcinoembryonic antigen
C1556094|T098|OSN|2039-6|LNC|carcinoembryonic antigen|carcinoembryonic antigen
C1556094|T098|LC|2039-6|LNC|carcinoembryonic antigen|carcinoembryonic antigen
C1556094|T098|LN|2039-6|LNC|CEA|CEA
C1556094|T098|MTH_LN|2039-6|LNC|CEA|CEA
C1556094|T098|OSN|2039-6|LNC|CEA|CEA
C1556094|T098|LC|2039-6|LNC|CEA|CEA
C1556099|T098|LC|2085-9|LNC|HDL cholesterol|HDL cholesterol
C1556099|T098|MTH_LN|2085-9|LNC|HDL cholesterol|HDL cholesterol
C1556099|T098|LN|2085-9|LNC|HDL cholesterol|HDL cholesterol
C1556099|T098|OSN|2085-9|LNC|HDL cholesterol|HDL cholesterol
C1556099|T098|LC|2085-9|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1556099|T098|MTH_LN|2085-9|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1556099|T098|LN|2085-9|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1556099|T098|OSN|2085-9|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1556099|T098|LC|2085-9|LNC|HDL-cholesterol|HDL-cholesterol
C1556099|T098|MTH_LN|2085-9|LNC|HDL-cholesterol|HDL-cholesterol
C1556099|T098|LN|2085-9|LNC|HDL-cholesterol|HDL-cholesterol
C1556099|T098|OSN|2085-9|LNC|HDL-cholesterol|HDL-cholesterol
C1556099|T098|LC|2085-9|LNC|high-density lipoprotein|high-density lipoprotein
C1556099|T098|MTH_LN|2085-9|LNC|high-density lipoprotein|high-density lipoprotein
C1556099|T098|LN|2085-9|LNC|high-density lipoprotein|high-density lipoprotein
C1556099|T098|OSN|2085-9|LNC|high-density lipoprotein|high-density lipoprotein
C1556099|T098|LC|2085-9|LNC|HDL|HDL
C1556099|T098|MTH_LN|2085-9|LNC|HDL|HDL
C1556099|T098|LN|2085-9|LNC|HDL|HDL
C1556099|T098|OSN|2085-9|LNC|HDL|HDL
C1556108|T098|LN|2082-6|LNC|cholesterol|cholesterol
C1556108|T098|MTH_LN|2082-6|LNC|cholesterol|cholesterol
C1556108|T098|OSN|2082-6|LNC|cholesterol|cholesterol
C1556108|T098|LC|2082-6|LNC|cholesterol|cholesterol
C1556108|T098|LN|2082-6|LNC|total cholesterol|total cholesterol
C1556108|T098|MTH_LN|2082-6|LNC|total cholesterol|total cholesterol
C1556108|T098|OSN|2082-6|LNC|total cholesterol|total cholesterol
C1556108|T098|LC|2082-6|LNC|total cholesterol|total cholesterol
C1556108|T098|LN|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C1556108|T098|MTH_LN|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C1556108|T098|OSN|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C1556108|T098|LC|2082-6|LNC|cholesterol metabolism|cholesterol metabolism
C1624127|T201|LN|42678-3|LNC|urate|urate
C1624127|T201|MTH_LN|42678-3|LNC|urate|urate
C1624127|T201|OSN|42678-3|LNC|urate|urate
C1624127|T201|LC|42678-3|LNC|urate|urate
C1624127|T201|LN|42678-3|LNC|uric acid|uric acid
C1624127|T201|MTH_LN|42678-3|LNC|uric acid|uric acid
C1624127|T201|OSN|42678-3|LNC|uric acid|uric acid
C1624127|T201|LC|42678-3|LNC|uric acid|uric acid
C1624714|T201|LN|42758-3|LNC|reticulocytes|reticulocytes
C1624714|T201|OSN|42758-3|LNC|reticulocytes|reticulocytes
C1624714|T201|MTH_LN|42758-3|LNC|reticulocytes|reticulocytes
C1624714|T201|LC|42758-3|LNC|reticulocytes|reticulocytes
C1624714|T201|LN|42758-3|LNC|reticulocyte count|reticulocyte count
C1624714|T201|OSN|42758-3|LNC|reticulocyte count|reticulocyte count
C1624714|T201|MTH_LN|42758-3|LNC|reticulocyte count|reticulocyte count
C1624714|T201|LC|42758-3|LNC|reticulocyte count|reticulocyte count
C1626179|T201|LN|42180-0|LNC|C-peptide|C-peptide
C1626179|T201|MTH_LN|42180-0|LNC|C-peptide|C-peptide
C1626179|T201|OSN|42180-0|LNC|C-peptide|C-peptide
C1626179|T201|LC|42180-0|LNC|C-peptide|C-peptide
C1626179|T201|LN|42180-0|LNC|C peptide|C peptide
C1626179|T201|MTH_LN|42180-0|LNC|C peptide|C peptide
C1626179|T201|OSN|42180-0|LNC|C peptide|C peptide
C1626179|T201|LC|42180-0|LNC|C peptide|C peptide
C1627306|T201|LN|42203-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1627306|T201|OSN|42203-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1627306|T201|MTH_LN|42203-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1627306|T201|LC|42203-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1627910|T201|LN|42908-4|LNC|hematocrit|hematocrit
C1627910|T201|MTH_LN|42908-4|LNC|hematocrit|hematocrit
C1627910|T201|LC|42908-4|LNC|hematocrit|hematocrit
C1627910|T201|OSN|42908-4|LNC|hematocrit|hematocrit
C1632378|T201|LN|41654-5|LNC|hematocrit|hematocrit
C1632378|T201|MTH_LN|41654-5|LNC|hematocrit|hematocrit
C1632378|T201|LC|41654-5|LNC|hematocrit|hematocrit
C1632378|T201|OSN|41654-5|LNC|hematocrit|hematocrit
C1633476|T201|LN|42857-3|LNC|calcium|calcium
C1633476|T201|OSN|42857-3|LNC|calcium|calcium
C1633476|T201|MTH_LN|42857-3|LNC|calcium|calcium
C1633476|T201|LC|42857-3|LNC|calcium|calcium
C1633476|T201|LN|42857-3|LNC|calcium homeostasis|calcium homeostasis
C1633476|T201|OSN|42857-3|LNC|calcium homeostasis|calcium homeostasis
C1633476|T201|MTH_LN|42857-3|LNC|calcium homeostasis|calcium homeostasis
C1633476|T201|LC|42857-3|LNC|calcium homeostasis|calcium homeostasis
C1638459|T201|LN|42937-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1638459|T201|MTH_LN|42937-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1638459|T201|LC|42937-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1638459|T201|OSN|42937-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1639938|T201|LN|42593-4|LNC|calcium|calcium
C1639938|T201|OSN|42593-4|LNC|calcium|calcium
C1639938|T201|MTH_LN|42593-4|LNC|calcium|calcium
C1639938|T201|LC|42593-4|LNC|calcium|calcium
C1639938|T201|LN|42593-4|LNC|calcium homeostasis|calcium homeostasis
C1639938|T201|OSN|42593-4|LNC|calcium homeostasis|calcium homeostasis
C1639938|T201|MTH_LN|42593-4|LNC|calcium homeostasis|calcium homeostasis
C1639938|T201|LC|42593-4|LNC|calcium homeostasis|calcium homeostasis
C1641514|T201|LN|41646-1|LNC|calcium|calcium
C1641514|T201|OSN|41646-1|LNC|calcium|calcium
C1641514|T201|MTH_LN|41646-1|LNC|calcium|calcium
C1641514|T201|LC|41646-1|LNC|calcium|calcium
C1641514|T201|LN|41646-1|LNC|calcium homeostasis|calcium homeostasis
C1641514|T201|OSN|41646-1|LNC|calcium homeostasis|calcium homeostasis
C1641514|T201|MTH_LN|41646-1|LNC|calcium homeostasis|calcium homeostasis
C1641514|T201|LC|41646-1|LNC|calcium homeostasis|calcium homeostasis
C1641515|T201|LN|41647-9|LNC|carbon dioxide|carbon dioxide
C1641515|T201|MTH_LN|41647-9|LNC|carbon dioxide|carbon dioxide
C1641515|T201|OSN|41647-9|LNC|carbon dioxide|carbon dioxide
C1641515|T201|LC|41647-9|LNC|carbon dioxide|carbon dioxide
C1642078|T201|LN|41655-2|LNC|hematocrit|hematocrit
C1642078|T201|MTH_LN|41655-2|LNC|hematocrit|hematocrit
C1642078|T201|LC|41655-2|LNC|hematocrit|hematocrit
C1642078|T201|OSN|41655-2|LNC|hematocrit|hematocrit
C1642581|T201|LN|41644-6|LNC|calcium|calcium
C1642581|T201|OSN|41644-6|LNC|calcium|calcium
C1642581|T201|MTH_LN|41644-6|LNC|calcium|calcium
C1642581|T201|LC|41644-6|LNC|calcium|calcium
C1642581|T201|LN|41644-6|LNC|calcium homeostasis|calcium homeostasis
C1642581|T201|OSN|41644-6|LNC|calcium homeostasis|calcium homeostasis
C1642581|T201|MTH_LN|41644-6|LNC|calcium homeostasis|calcium homeostasis
C1642581|T201|LC|41644-6|LNC|calcium homeostasis|calcium homeostasis
C1645723|T201|LN|41653-7|LNC|glucose|glucose
C1645723|T201|OSN|41653-7|LNC|glucose|glucose
C1645723|T201|MTH_LN|41653-7|LNC|glucose|glucose
C1645723|T201|LC|41653-7|LNC|glucose|glucose
C1646772|T201|LN|42757-5|LNC|troponin I|troponin I
C1646772|T201|OSN|42757-5|LNC|troponin I|troponin I
C1646772|T201|MTH_LN|42757-5|LNC|troponin I|troponin I
C1646772|T201|LC|42757-5|LNC|troponin I|troponin I
C1649478|T201|LN|41407-8|LNC|cortisol|cortisol
C1649478|T201|OSN|41407-8|LNC|cortisol|cortisol
C1649478|T201|MTH_LN|41407-8|LNC|cortisol|cortisol
C1649478|T201|LC|41407-8|LNC|cortisol|cortisol
C1649478|T201|LN|41407-8|LNC|cortisol low|cortisol low
C1649478|T201|OSN|41407-8|LNC|cortisol low|cortisol low
C1649478|T201|MTH_LN|41407-8|LNC|cortisol low|cortisol low
C1649478|T201|LC|41407-8|LNC|cortisol low|cortisol low
C1649478|T201|LN|41407-8|LNC|to undetectable cortisol|to undetectable cortisol
C1649478|T201|OSN|41407-8|LNC|to undetectable cortisol|to undetectable cortisol
C1649478|T201|MTH_LN|41407-8|LNC|to undetectable cortisol|to undetectable cortisol
C1649478|T201|LC|41407-8|LNC|to undetectable cortisol|to undetectable cortisol
C1651491|T201|LN|41645-3|LNC|calcium|calcium
C1651491|T201|OSN|41645-3|LNC|calcium|calcium
C1651491|T201|MTH_LN|41645-3|LNC|calcium|calcium
C1651491|T201|LC|41645-3|LNC|calcium|calcium
C1651491|T201|LN|41645-3|LNC|calcium homeostasis|calcium homeostasis
C1651491|T201|OSN|41645-3|LNC|calcium homeostasis|calcium homeostasis
C1651491|T201|MTH_LN|41645-3|LNC|calcium homeostasis|calcium homeostasis
C1651491|T201|LC|41645-3|LNC|calcium homeostasis|calcium homeostasis
C1652145|T201|LN|42251-9|LNC|methadone test|methadone test
C1652145|T201|MTH_LN|42251-9|LNC|methadone test|methadone test
C1652145|T201|OSN|42251-9|LNC|methadone test|methadone test
C1652145|T201|LC|42251-9|LNC|methadone test|methadone test
C1654330|T201|LN|42932-4|LNC|T cell CD40 expression|T cell CD40 expression
C1654330|T201|MTH_LN|42932-4|LNC|T cell CD40 expression|T cell CD40 expression
C1654330|T201|LC|42932-4|LNC|T cell CD40 expression|T cell CD40 expression
C1654330|T201|OSN|42932-4|LNC|T cell CD40 expression|T cell CD40 expression
C1654330|T201|LN|42932-4|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C1654330|T201|MTH_LN|42932-4|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C1654330|T201|LC|42932-4|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C1654330|T201|OSN|42932-4|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C1714488|T201|LN|43576-8|LNC|acylcarnitine|acylcarnitine
C1714488|T201|MTH_LN|43576-8|LNC|acylcarnitine|acylcarnitine
C1714488|T201|OSN|43576-8|LNC|acylcarnitine|acylcarnitine
C1714488|T201|LC|43576-8|LNC|acylcarnitine|acylcarnitine
C1714568|T201|LN|43196-5|LNC|xenobiotic|xenobiotic
C1714568|T201|LC|43196-5|LNC|xenobiotic|xenobiotic
C1714568|T201|OSN|43196-5|LNC|xenobiotic|xenobiotic
C1714568|T201|MTH_LN|43196-5|LNC|xenobiotic|xenobiotic
C1714607|T201|LN|43240-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1714607|T201|OSN|43240-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1714607|T201|MTH_LN|43240-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1714607|T201|LC|43240-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1714608|T201|LN|43241-9|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1714608|T201|OSN|43241-9|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1714608|T201|MTH_LN|43241-9|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1714608|T201|LC|43241-9|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1714736|T201|LN|43392-0|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714736|T201|OSN|43392-0|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714736|T201|LC|43392-0|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714736|T201|MTH_LN|43392-0|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714736|T201|LN|43392-0|LNC|LDL|LDL
C1714736|T201|OSN|43392-0|LNC|LDL|LDL
C1714736|T201|LC|43392-0|LNC|LDL|LDL
C1714736|T201|MTH_LN|43392-0|LNC|LDL|LDL
C1714736|T201|LN|43392-0|LNC|LDL cholesterol|LDL cholesterol
C1714736|T201|OSN|43392-0|LNC|LDL cholesterol|LDL cholesterol
C1714736|T201|LC|43392-0|LNC|LDL cholesterol|LDL cholesterol
C1714736|T201|MTH_LN|43392-0|LNC|LDL cholesterol|LDL cholesterol
C1714736|T201|LN|43392-0|LNC|low-density lipoprotein|low-density lipoprotein
C1714736|T201|OSN|43392-0|LNC|low-density lipoprotein|low-density lipoprotein
C1714736|T201|LC|43392-0|LNC|low-density lipoprotein|low-density lipoprotein
C1714736|T201|MTH_LN|43392-0|LNC|low-density lipoprotein|low-density lipoprotein
C1714736|T201|LN|43392-0|LNC|beta-lipoproteins|beta-lipoproteins
C1714736|T201|OSN|43392-0|LNC|beta-lipoproteins|beta-lipoproteins
C1714736|T201|LC|43392-0|LNC|beta-lipoproteins|beta-lipoproteins
C1714736|T201|MTH_LN|43392-0|LNC|beta-lipoproteins|beta-lipoproteins
C1714736|T201|LN|43392-0|LNC|LDL-C|LDL-C
C1714736|T201|OSN|43392-0|LNC|LDL-C|LDL-C
C1714736|T201|LC|43392-0|LNC|LDL-C|LDL-C
C1714736|T201|MTH_LN|43392-0|LNC|LDL-C|LDL-C
C1714737|T201|LN|43393-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714737|T201|LC|43393-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714737|T201|MTH_LN|43393-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714737|T201|OSN|43393-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714737|T201|LN|43393-8|LNC|LDL|LDL
C1714737|T201|LC|43393-8|LNC|LDL|LDL
C1714737|T201|MTH_LN|43393-8|LNC|LDL|LDL
C1714737|T201|OSN|43393-8|LNC|LDL|LDL
C1714737|T201|LN|43393-8|LNC|LDL cholesterol|LDL cholesterol
C1714737|T201|LC|43393-8|LNC|LDL cholesterol|LDL cholesterol
C1714737|T201|MTH_LN|43393-8|LNC|LDL cholesterol|LDL cholesterol
C1714737|T201|OSN|43393-8|LNC|LDL cholesterol|LDL cholesterol
C1714737|T201|LN|43393-8|LNC|low-density lipoprotein|low-density lipoprotein
C1714737|T201|LC|43393-8|LNC|low-density lipoprotein|low-density lipoprotein
C1714737|T201|MTH_LN|43393-8|LNC|low-density lipoprotein|low-density lipoprotein
C1714737|T201|OSN|43393-8|LNC|low-density lipoprotein|low-density lipoprotein
C1714737|T201|LN|43393-8|LNC|beta-lipoproteins|beta-lipoproteins
C1714737|T201|LC|43393-8|LNC|beta-lipoproteins|beta-lipoproteins
C1714737|T201|MTH_LN|43393-8|LNC|beta-lipoproteins|beta-lipoproteins
C1714737|T201|OSN|43393-8|LNC|beta-lipoproteins|beta-lipoproteins
C1714737|T201|LN|43393-8|LNC|LDL-C|LDL-C
C1714737|T201|LC|43393-8|LNC|LDL-C|LDL-C
C1714737|T201|MTH_LN|43393-8|LNC|LDL-C|LDL-C
C1714737|T201|OSN|43393-8|LNC|LDL-C|LDL-C
C1714738|T201|LN|43394-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714738|T201|OSN|43394-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714738|T201|MTH_LN|43394-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714738|T201|LC|43394-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1714738|T201|LN|43394-6|LNC|LDL|LDL
C1714738|T201|OSN|43394-6|LNC|LDL|LDL
C1714738|T201|MTH_LN|43394-6|LNC|LDL|LDL
C1714738|T201|LC|43394-6|LNC|LDL|LDL
C1714738|T201|LN|43394-6|LNC|LDL cholesterol|LDL cholesterol
C1714738|T201|OSN|43394-6|LNC|LDL cholesterol|LDL cholesterol
C1714738|T201|MTH_LN|43394-6|LNC|LDL cholesterol|LDL cholesterol
C1714738|T201|LC|43394-6|LNC|LDL cholesterol|LDL cholesterol
C1714738|T201|LN|43394-6|LNC|low-density lipoprotein|low-density lipoprotein
C1714738|T201|OSN|43394-6|LNC|low-density lipoprotein|low-density lipoprotein
C1714738|T201|MTH_LN|43394-6|LNC|low-density lipoprotein|low-density lipoprotein
C1714738|T201|LC|43394-6|LNC|low-density lipoprotein|low-density lipoprotein
C1714738|T201|LN|43394-6|LNC|beta-lipoproteins|beta-lipoproteins
C1714738|T201|OSN|43394-6|LNC|beta-lipoproteins|beta-lipoproteins
C1714738|T201|MTH_LN|43394-6|LNC|beta-lipoproteins|beta-lipoproteins
C1714738|T201|LC|43394-6|LNC|beta-lipoproteins|beta-lipoproteins
C1714738|T201|LN|43394-6|LNC|LDL-C|LDL-C
C1714738|T201|OSN|43394-6|LNC|LDL-C|LDL-C
C1714738|T201|MTH_LN|43394-6|LNC|LDL-C|LDL-C
C1714738|T201|LC|43394-6|LNC|LDL-C|LDL-C
C1714757|T201|LN|43416-7|LNC|hematocrit|hematocrit
C1714757|T201|MTH_LN|43416-7|LNC|hematocrit|hematocrit
C1714757|T201|LC|43416-7|LNC|hematocrit|hematocrit
C1714757|T201|OSN|43416-7|LNC|hematocrit|hematocrit
C1714998|T201|LN|43623-8|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1714998|T201|MTH_LN|43623-8|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1714998|T201|OSN|43623-8|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1714998|T201|LC|43623-8|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1714999|T201|LN|43624-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1714999|T201|MTH_LN|43624-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1714999|T201|OSN|43624-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1714999|T201|LC|43624-6|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1715000|T201|LN|43625-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1715000|T201|MTH_LN|43625-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1715000|T201|OSN|43625-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1715000|T201|LC|43625-3|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C1715064|T201|LN|43715-2|LNC|acylcarnitine|acylcarnitine
C1715064|T201|MTH_LN|43715-2|LNC|acylcarnitine|acylcarnitine
C1715064|T201|OSN|43715-2|LNC|acylcarnitine|acylcarnitine
C1715064|T201|LC|43715-2|LNC|acylcarnitine|acylcarnitine
C1715066|T201|LN|43717-8|LNC|acylcarnitine|acylcarnitine
C1715066|T201|MTH_LN|43717-8|LNC|acylcarnitine|acylcarnitine
C1715066|T201|LC|43717-8|LNC|acylcarnitine|acylcarnitine
C1715066|T201|OSN|43717-8|LNC|acylcarnitine|acylcarnitine
C1715250|T201|LN|43962-0|LNC|naive T|naive T
C1715250|T201|MTH_LN|43962-0|LNC|naive T|naive T
C1715250|T201|LC|43962-0|LNC|naive T|naive T
C1715250|T201|OSN|43962-0|LNC|naive T|naive T
C1715250|T201|LN|43962-0|LNC|naive T cell|naive T cell
C1715250|T201|MTH_LN|43962-0|LNC|naive T cell|naive T cell
C1715250|T201|LC|43962-0|LNC|naive T cell|naive T cell
C1715250|T201|OSN|43962-0|LNC|naive T cell|naive T cell
C1715251|T201|LN|43963-8|LNC|naive T|naive T
C1715251|T201|MTH_LN|43963-8|LNC|naive T|naive T
C1715251|T201|LC|43963-8|LNC|naive T|naive T
C1715251|T201|OSN|43963-8|LNC|naive T|naive T
C1715251|T201|LN|43963-8|LNC|naive T cell|naive T cell
C1715251|T201|MTH_LN|43963-8|LNC|naive T cell|naive T cell
C1715251|T201|LC|43963-8|LNC|naive T cell|naive T cell
C1715251|T201|OSN|43963-8|LNC|naive T cell|naive T cell
C1715252|T201|LN|43964-6|LNC|naive T|naive T
C1715252|T201|MTH_LN|43964-6|LNC|naive T|naive T
C1715252|T201|LC|43964-6|LNC|naive T|naive T
C1715252|T201|OSN|43964-6|LNC|naive T|naive T
C1715252|T201|LN|43964-6|LNC|naive T cell|naive T cell
C1715252|T201|MTH_LN|43964-6|LNC|naive T cell|naive T cell
C1715252|T201|LC|43964-6|LNC|naive T cell|naive T cell
C1715252|T201|OSN|43964-6|LNC|naive T cell|naive T cell
C1715253|T201|LN|43965-3|LNC|naive T|naive T
C1715253|T201|MTH_LN|43965-3|LNC|naive T|naive T
C1715253|T201|LC|43965-3|LNC|naive T|naive T
C1715253|T201|OSN|43965-3|LNC|naive T|naive T
C1715253|T201|LN|43965-3|LNC|naive T cell|naive T cell
C1715253|T201|MTH_LN|43965-3|LNC|naive T cell|naive T cell
C1715253|T201|LC|43965-3|LNC|naive T cell|naive T cell
C1715253|T201|OSN|43965-3|LNC|naive T cell|naive T cell
C1715553|T201|LN|44299-6|LNC|arginine|arginine
C1715553|T201|MTH_LN|44299-6|LNC|arginine|arginine
C1715553|T201|OSN|44299-6|LNC|arginine|arginine
C1715553|T201|LC|44299-6|LNC|arginine|arginine
C1715640|T201|LN|44411-7|LNC|taurine|taurine
C1715640|T201|MTH_LN|44411-7|LNC|taurine|taurine
C1715640|T201|OSN|44411-7|LNC|taurine|taurine
C1715640|T201|LC|44411-7|LNC|taurine|taurine
C1715977|T201|LN|44750-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1715977|T201|MTH_LN|44750-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1715977|T201|LC|44750-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1715977|T201|OSN|44750-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1716121|T201|LN|44915-7|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1716121|T201|OSN|44915-7|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1716121|T201|LC|44915-7|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1716121|T201|MTH_LN|44915-7|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1716121|T201|LN|44915-7|LNC|LDL|LDL
C1716121|T201|OSN|44915-7|LNC|LDL|LDL
C1716121|T201|LC|44915-7|LNC|LDL|LDL
C1716121|T201|MTH_LN|44915-7|LNC|LDL|LDL
C1716121|T201|LN|44915-7|LNC|LDL cholesterol|LDL cholesterol
C1716121|T201|OSN|44915-7|LNC|LDL cholesterol|LDL cholesterol
C1716121|T201|LC|44915-7|LNC|LDL cholesterol|LDL cholesterol
C1716121|T201|MTH_LN|44915-7|LNC|LDL cholesterol|LDL cholesterol
C1716121|T201|LN|44915-7|LNC|low-density lipoprotein|low-density lipoprotein
C1716121|T201|OSN|44915-7|LNC|low-density lipoprotein|low-density lipoprotein
C1716121|T201|LC|44915-7|LNC|low-density lipoprotein|low-density lipoprotein
C1716121|T201|MTH_LN|44915-7|LNC|low-density lipoprotein|low-density lipoprotein
C1716121|T201|LN|44915-7|LNC|beta-lipoproteins|beta-lipoproteins
C1716121|T201|OSN|44915-7|LNC|beta-lipoproteins|beta-lipoproteins
C1716121|T201|LC|44915-7|LNC|beta-lipoproteins|beta-lipoproteins
C1716121|T201|MTH_LN|44915-7|LNC|beta-lipoproteins|beta-lipoproteins
C1716121|T201|LN|44915-7|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1716121|T201|OSN|44915-7|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1716121|T201|LC|44915-7|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1716121|T201|MTH_LN|44915-7|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1716121|T201|LN|44915-7|LNC|LDL-C|LDL-C
C1716121|T201|OSN|44915-7|LNC|LDL-C|LDL-C
C1716121|T201|LC|44915-7|LNC|LDL-C|LDL-C
C1716121|T201|MTH_LN|44915-7|LNC|LDL-C|LDL-C
C1716137|T201|LN|44933-0|LNC|osmolality|osmolality
C1716137|T201|MTH_LN|44933-0|LNC|osmolality|osmolality
C1716137|T201|OSN|44933-0|LNC|osmolality|osmolality
C1716137|T201|LC|44933-0|LNC|osmolality|osmolality
C1716137|T201|LN|44933-0|LNC|homeostasis|homeostasis
C1716137|T201|MTH_LN|44933-0|LNC|homeostasis|homeostasis
C1716137|T201|OSN|44933-0|LNC|homeostasis|homeostasis
C1716137|T201|LC|44933-0|LNC|homeostasis|homeostasis
C1716316|T201|LN|45169-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1716316|T201|MTH_LN|45169-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1716316|T201|OSN|45169-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1716316|T201|LC|45169-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1716495|T201|LN|45383-7|LNC|neutrophil count|neutrophil count
C1716495|T201|MTH_LN|45383-7|LNC|neutrophil count|neutrophil count
C1716495|T201|OSN|45383-7|LNC|neutrophil count|neutrophil count
C1716495|T201|LC|45383-7|LNC|neutrophil count|neutrophil count
C1716495|T201|LN|45383-7|LNC|cytology|cytology
C1716495|T201|MTH_LN|45383-7|LNC|cytology|cytology
C1716495|T201|OSN|45383-7|LNC|cytology|cytology
C1716495|T201|LC|45383-7|LNC|cytology|cytology
C1717133|T201|LN|46099-8|LNC|calcium|calcium
C1717133|T201|OSN|46099-8|LNC|calcium|calcium
C1717133|T201|MTH_LN|46099-8|LNC|calcium|calcium
C1717133|T201|LC|46099-8|LNC|calcium|calcium
C1717133|T201|LN|46099-8|LNC|calcium homeostasis|calcium homeostasis
C1717133|T201|OSN|46099-8|LNC|calcium homeostasis|calcium homeostasis
C1717133|T201|MTH_LN|46099-8|LNC|calcium homeostasis|calcium homeostasis
C1717133|T201|LC|46099-8|LNC|calcium homeostasis|calcium homeostasis
C1717305|T201|LN|44050-3|LNC|glucosephosphate isomerase activity|glucosephosphate isomerase activity
C1717305|T201|OSN|44050-3|LNC|glucosephosphate isomerase activity|glucosephosphate isomerase activity
C1717305|T201|MTH_LN|44050-3|LNC|glucosephosphate isomerase activity|glucosephosphate isomerase activity
C1717305|T201|LC|44050-3|LNC|glucosephosphate isomerase activity|glucosephosphate isomerase activity
C1717305|T201|LN|44050-3|LNC|glucose phosphate isomerase activity|glucose phosphate isomerase activity
C1717305|T201|OSN|44050-3|LNC|glucose phosphate isomerase activity|glucose phosphate isomerase activity
C1717305|T201|MTH_LN|44050-3|LNC|glucose phosphate isomerase activity|glucose phosphate isomerase activity
C1717305|T201|LC|44050-3|LNC|glucose phosphate isomerase activity|glucose phosphate isomerase activity
C1744633|T201|LN|24122-4|LNC|neutrophil count|neutrophil count
C1744633|T201|OSN|24122-4|LNC|neutrophil count|neutrophil count
C1744633|T201|MTH_LN|24122-4|LNC|neutrophil count|neutrophil count
C1744633|T201|LC|24122-4|LNC|neutrophil count|neutrophil count
C1744633|T201|LN|24122-4|LNC|cytology|cytology
C1744633|T201|OSN|24122-4|LNC|cytology|cytology
C1744633|T201|MTH_LN|24122-4|LNC|cytology|cytology
C1744633|T201|LC|24122-4|LNC|cytology|cytology
C1830099|T201|LN|46269-7|LNC|vitamin D metabolism|vitamin D metabolism
C1830099|T201|MTH_LN|46269-7|LNC|vitamin D metabolism|vitamin D metabolism
C1830099|T201|LC|46269-7|LNC|vitamin D metabolism|vitamin D metabolism
C1830099|T201|OSN|46269-7|LNC|vitamin D metabolism|vitamin D metabolism
C1830099|T201|LN|46269-7|LNC|calcifediol|calcifediol
C1830099|T201|MTH_LN|46269-7|LNC|calcifediol|calcifediol
C1830099|T201|LC|46269-7|LNC|calcifediol|calcifediol
C1830099|T201|OSN|46269-7|LNC|calcifediol|calcifediol
C1830099|T201|LN|46269-7|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1830099|T201|MTH_LN|46269-7|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1830099|T201|LC|46269-7|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1830099|T201|OSN|46269-7|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1830099|T201|LN|46269-7|LNC|calcidiol|calcidiol
C1830099|T201|MTH_LN|46269-7|LNC|calcidiol|calcidiol
C1830099|T201|LC|46269-7|LNC|calcidiol|calcidiol
C1830099|T201|OSN|46269-7|LNC|calcidiol|calcidiol
C1830289|T201|LN|46400-8|LNC|ACTH|ACTH
C1830289|T201|MTH_LN|46400-8|LNC|ACTH|ACTH
C1830289|T201|OSN|46400-8|LNC|ACTH|ACTH
C1830289|T201|LC|46400-8|LNC|ACTH|ACTH
C1830289|T201|LN|46400-8|LNC|corticotropin|corticotropin
C1830289|T201|MTH_LN|46400-8|LNC|corticotropin|corticotropin
C1830289|T201|OSN|46400-8|LNC|corticotropin|corticotropin
C1830289|T201|LC|46400-8|LNC|corticotropin|corticotropin
C1830289|T201|LN|46400-8|LNC|adrenocorticotropin|adrenocorticotropin
C1830289|T201|MTH_LN|46400-8|LNC|adrenocorticotropin|adrenocorticotropin
C1830289|T201|OSN|46400-8|LNC|adrenocorticotropin|adrenocorticotropin
C1830289|T201|LC|46400-8|LNC|adrenocorticotropin|adrenocorticotropin
C1830290|T201|LN|46401-6|LNC|ACTH|ACTH
C1830290|T201|MTH_LN|46401-6|LNC|ACTH|ACTH
C1830290|T201|OSN|46401-6|LNC|ACTH|ACTH
C1830290|T201|LC|46401-6|LNC|ACTH|ACTH
C1830290|T201|LN|46401-6|LNC|corticotropin|corticotropin
C1830290|T201|MTH_LN|46401-6|LNC|corticotropin|corticotropin
C1830290|T201|OSN|46401-6|LNC|corticotropin|corticotropin
C1830290|T201|LC|46401-6|LNC|corticotropin|corticotropin
C1830290|T201|LN|46401-6|LNC|adrenocorticotropin|adrenocorticotropin
C1830290|T201|MTH_LN|46401-6|LNC|adrenocorticotropin|adrenocorticotropin
C1830290|T201|OSN|46401-6|LNC|adrenocorticotropin|adrenocorticotropin
C1830290|T201|LC|46401-6|LNC|adrenocorticotropin|adrenocorticotropin
C1830291|T201|LN|46402-4|LNC|ACTH|ACTH
C1830291|T201|OSN|46402-4|LNC|ACTH|ACTH
C1830291|T201|MTH_LN|46402-4|LNC|ACTH|ACTH
C1830291|T201|LC|46402-4|LNC|ACTH|ACTH
C1830291|T201|LN|46402-4|LNC|corticotropin|corticotropin
C1830291|T201|OSN|46402-4|LNC|corticotropin|corticotropin
C1830291|T201|MTH_LN|46402-4|LNC|corticotropin|corticotropin
C1830291|T201|LC|46402-4|LNC|corticotropin|corticotropin
C1830291|T201|LN|46402-4|LNC|adrenocorticotropin|adrenocorticotropin
C1830291|T201|OSN|46402-4|LNC|adrenocorticotropin|adrenocorticotropin
C1830291|T201|MTH_LN|46402-4|LNC|adrenocorticotropin|adrenocorticotropin
C1830291|T201|LC|46402-4|LNC|adrenocorticotropin|adrenocorticotropin
C1830303|T201|LN|46414-9|LNC|luteinizing|luteinizing
C1830303|T201|MTH_LN|46414-9|LNC|luteinizing|luteinizing
C1830303|T201|OSN|46414-9|LNC|luteinizing|luteinizing
C1830303|T201|LC|46414-9|LNC|luteinizing|luteinizing
C1830303|T201|LN|46414-9|LNC|LH|LH
C1830303|T201|MTH_LN|46414-9|LNC|LH|LH
C1830303|T201|OSN|46414-9|LNC|LH|LH
C1830303|T201|LC|46414-9|LNC|LH|LH
C1830303|T201|LN|46414-9|LNC|luteinising|luteinising
C1830303|T201|MTH_LN|46414-9|LNC|luteinising|luteinising
C1830303|T201|OSN|46414-9|LNC|luteinising|luteinising
C1830303|T201|LC|46414-9|LNC|luteinising|luteinising
C1830304|T201|LN|46415-6|LNC|luteinizing|luteinizing
C1830304|T201|OSN|46415-6|LNC|luteinizing|luteinizing
C1830304|T201|MTH_LN|46415-6|LNC|luteinizing|luteinizing
C1830304|T201|LC|46415-6|LNC|luteinizing|luteinizing
C1830304|T201|LN|46415-6|LNC|LH|LH
C1830304|T201|OSN|46415-6|LNC|LH|LH
C1830304|T201|MTH_LN|46415-6|LNC|LH|LH
C1830304|T201|LC|46415-6|LNC|LH|LH
C1830304|T201|LN|46415-6|LNC|luteinising|luteinising
C1830304|T201|OSN|46415-6|LNC|luteinising|luteinising
C1830304|T201|MTH_LN|46415-6|LNC|luteinising|luteinising
C1830304|T201|LC|46415-6|LNC|luteinising|luteinising
// C1830308|T201|LN|46419-8|LNC||
// C1830308|T201|OSN|46419-8|LNC||
// C1830308|T201|MTH_LN|46419-8|LNC||
// C1830308|T201|LC|46419-8|LNC||
C1830308|T201|LN|46419-8|LNC|occult|occult
C1830308|T201|OSN|46419-8|LNC|occult|occult
C1830308|T201|MTH_LN|46419-8|LNC|occult|occult
C1830308|T201|LC|46419-8|LNC|occult|occult
C1830310|T201|LN|46421-4|LNC|homeostasis|homeostasis
C1830310|T201|MTH_LN|46421-4|LNC|homeostasis|homeostasis
C1830310|T201|LC|46421-4|LNC|homeostasis|homeostasis
C1830310|T201|OSN|46421-4|LNC|homeostasis|homeostasis
C1830776|T201|LN|46702-7|LNC|neutrophil count|neutrophil count
C1830776|T201|MTH_LN|46702-7|LNC|neutrophil count|neutrophil count
C1830776|T201|OSN|46702-7|LNC|neutrophil count|neutrophil count
C1830776|T201|LC|46702-7|LNC|neutrophil count|neutrophil count
C1831046|T201|LN|46967-6|LNC|T cell CD40 expression|T cell CD40 expression
C1831046|T201|OSN|46967-6|LNC|T cell CD40 expression|T cell CD40 expression
C1831046|T201|MTH_LN|46967-6|LNC|T cell CD40 expression|T cell CD40 expression
C1831046|T201|LC|46967-6|LNC|T cell CD40 expression|T cell CD40 expression
C1831046|T201|LN|46967-6|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C1831046|T201|OSN|46967-6|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C1831046|T201|MTH_LN|46967-6|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C1831046|T201|LC|46967-6|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C1831079|T201|LN|46984-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1831079|T201|LC|46984-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1831079|T201|MTH_LN|46984-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1831079|T201|OSN|46984-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1831079|T201|LN|46984-1|LNC|LDL|LDL
C1831079|T201|LC|46984-1|LNC|LDL|LDL
C1831079|T201|MTH_LN|46984-1|LNC|LDL|LDL
C1831079|T201|OSN|46984-1|LNC|LDL|LDL
C1831079|T201|LN|46984-1|LNC|LDL cholesterol|LDL cholesterol
C1831079|T201|LC|46984-1|LNC|LDL cholesterol|LDL cholesterol
C1831079|T201|MTH_LN|46984-1|LNC|LDL cholesterol|LDL cholesterol
C1831079|T201|OSN|46984-1|LNC|LDL cholesterol|LDL cholesterol
C1831079|T201|LN|46984-1|LNC|low-density lipoprotein|low-density lipoprotein
C1831079|T201|LC|46984-1|LNC|low-density lipoprotein|low-density lipoprotein
C1831079|T201|MTH_LN|46984-1|LNC|low-density lipoprotein|low-density lipoprotein
C1831079|T201|OSN|46984-1|LNC|low-density lipoprotein|low-density lipoprotein
C1831079|T201|LN|46984-1|LNC|beta-lipoproteins|beta-lipoproteins
C1831079|T201|LC|46984-1|LNC|beta-lipoproteins|beta-lipoproteins
C1831079|T201|MTH_LN|46984-1|LNC|beta-lipoproteins|beta-lipoproteins
C1831079|T201|OSN|46984-1|LNC|beta-lipoproteins|beta-lipoproteins
C1831079|T201|LN|46984-1|LNC|LDL-C|LDL-C
C1831079|T201|LC|46984-1|LNC|LDL-C|LDL-C
C1831079|T201|MTH_LN|46984-1|LNC|LDL-C|LDL-C
C1831079|T201|OSN|46984-1|LNC|LDL-C|LDL-C
C1831080|T201|LN|46985-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1831080|T201|MTH_LN|46985-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1831080|T201|OSN|46985-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1831080|T201|LC|46985-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1831080|T201|LN|46985-8|LNC|LDL|LDL
C1831080|T201|MTH_LN|46985-8|LNC|LDL|LDL
C1831080|T201|OSN|46985-8|LNC|LDL|LDL
C1831080|T201|LC|46985-8|LNC|LDL|LDL
C1831080|T201|LN|46985-8|LNC|LDL cholesterol|LDL cholesterol
C1831080|T201|MTH_LN|46985-8|LNC|LDL cholesterol|LDL cholesterol
C1831080|T201|OSN|46985-8|LNC|LDL cholesterol|LDL cholesterol
C1831080|T201|LC|46985-8|LNC|LDL cholesterol|LDL cholesterol
C1831080|T201|LN|46985-8|LNC|low-density lipoprotein|low-density lipoprotein
C1831080|T201|MTH_LN|46985-8|LNC|low-density lipoprotein|low-density lipoprotein
C1831080|T201|OSN|46985-8|LNC|low-density lipoprotein|low-density lipoprotein
C1831080|T201|LC|46985-8|LNC|low-density lipoprotein|low-density lipoprotein
C1831080|T201|LN|46985-8|LNC|beta-lipoproteins|beta-lipoproteins
C1831080|T201|MTH_LN|46985-8|LNC|beta-lipoproteins|beta-lipoproteins
C1831080|T201|OSN|46985-8|LNC|beta-lipoproteins|beta-lipoproteins
C1831080|T201|LC|46985-8|LNC|beta-lipoproteins|beta-lipoproteins
C1831080|T201|LN|46985-8|LNC|LDL-C|LDL-C
C1831080|T201|MTH_LN|46985-8|LNC|LDL-C|LDL-C
C1831080|T201|OSN|46985-8|LNC|LDL-C|LDL-C
C1831080|T201|LC|46985-8|LNC|LDL-C|LDL-C
C1831081|T201|LN|46986-6|LNC|VLDL cholesterol|VLDL cholesterol
C1831081|T201|MTH_LN|46986-6|LNC|VLDL cholesterol|VLDL cholesterol
C1831081|T201|OSN|46986-6|LNC|VLDL cholesterol|VLDL cholesterol
C1831081|T201|LC|46986-6|LNC|VLDL cholesterol|VLDL cholesterol
C1831081|T201|LN|46986-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1831081|T201|MTH_LN|46986-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1831081|T201|OSN|46986-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1831081|T201|LC|46986-6|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1831081|T201|LN|46986-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1831081|T201|MTH_LN|46986-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1831081|T201|OSN|46986-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1831081|T201|LC|46986-6|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1952650|T201|LN|47843-8|LNC|ACTH|ACTH
C1952650|T201|OSN|47843-8|LNC|ACTH|ACTH
C1952650|T201|MTH_LN|47843-8|LNC|ACTH|ACTH
C1952650|T201|LC|47843-8|LNC|ACTH|ACTH
C1952650|T201|LN|47843-8|LNC|corticotropin|corticotropin
C1952650|T201|OSN|47843-8|LNC|corticotropin|corticotropin
C1952650|T201|MTH_LN|47843-8|LNC|corticotropin|corticotropin
C1952650|T201|LC|47843-8|LNC|corticotropin|corticotropin
C1952650|T201|LN|47843-8|LNC|adrenocorticotropin|adrenocorticotropin
C1952650|T201|OSN|47843-8|LNC|adrenocorticotropin|adrenocorticotropin
C1952650|T201|MTH_LN|47843-8|LNC|adrenocorticotropin|adrenocorticotropin
C1952650|T201|LC|47843-8|LNC|adrenocorticotropin|adrenocorticotropin
C1952753|T201|LN|47547-5|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1952753|T201|MTH_LN|47547-5|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1952753|T201|OSN|47547-5|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1952753|T201|LC|47547-5|LNC|cerebrospinal fluid 5-methyltetrahydrofolate|cerebrospinal fluid 5-methyltetrahydrofolate
C1952753|T201|LN|47547-5|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1952753|T201|MTH_LN|47547-5|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1952753|T201|OSN|47547-5|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1952753|T201|LC|47547-5|LNC|CSF 5-methyltetrahydrofolate|CSF 5-methyltetrahydrofolate
C1952753|T201|LN|47547-5|LNC|folate metabolism|folate metabolism
C1952753|T201|MTH_LN|47547-5|LNC|folate metabolism|folate metabolism
C1952753|T201|OSN|47547-5|LNC|folate metabolism|folate metabolism
C1952753|T201|LC|47547-5|LNC|folate metabolism|folate metabolism
C1952809|T201|LN|47579-8|LNC|bicarbonate|bicarbonate
C1952809|T201|MTH_LN|47579-8|LNC|bicarbonate|bicarbonate
C1952809|T201|OSN|47579-8|LNC|bicarbonate|bicarbonate
C1952809|T201|LC|47579-8|LNC|bicarbonate|bicarbonate
C1952810|T201|LN|47580-6|LNC|bicarbonate|bicarbonate
C1952810|T201|OSN|47580-6|LNC|bicarbonate|bicarbonate
C1952810|T201|MTH_LN|47580-6|LNC|bicarbonate|bicarbonate
C1952810|T201|LC|47580-6|LNC|bicarbonate|bicarbonate
C1952814|T201|LN|47583-0|LNC|C-peptide|C-peptide
C1952814|T201|OSN|47583-0|LNC|C-peptide|C-peptide
C1952814|T201|MTH_LN|47583-0|LNC|C-peptide|C-peptide
C1952814|T201|LC|47583-0|LNC|C-peptide|C-peptide
C1952814|T201|LN|47583-0|LNC|C peptide|C peptide
C1952814|T201|OSN|47583-0|LNC|C peptide|C peptide
C1952814|T201|MTH_LN|47583-0|LNC|C peptide|C peptide
C1952814|T201|LC|47583-0|LNC|C peptide|C peptide
C1952815|T201|LN|47584-8|LNC|C-peptide|C-peptide
C1952815|T201|MTH_LN|47584-8|LNC|C-peptide|C-peptide
C1952815|T201|OSN|47584-8|LNC|C-peptide|C-peptide
C1952815|T201|LC|47584-8|LNC|C-peptide|C-peptide
C1952815|T201|LN|47584-8|LNC|C peptide|C peptide
C1952815|T201|MTH_LN|47584-8|LNC|C peptide|C peptide
C1952815|T201|OSN|47584-8|LNC|C peptide|C peptide
C1952815|T201|LC|47584-8|LNC|C peptide|C peptide
C1952816|T201|LN|47585-5|LNC|C-peptide|C-peptide
C1952816|T201|OSN|47585-5|LNC|C-peptide|C-peptide
C1952816|T201|MTH_LN|47585-5|LNC|C-peptide|C-peptide
C1952816|T201|LC|47585-5|LNC|C-peptide|C-peptide
C1952816|T201|LN|47585-5|LNC|C peptide|C peptide
C1952816|T201|OSN|47585-5|LNC|C peptide|C peptide
C1952816|T201|MTH_LN|47585-5|LNC|C peptide|C peptide
C1952816|T201|LC|47585-5|LNC|C peptide|C peptide
C1952817|T201|LN|47586-3|LNC|C-peptide|C-peptide
C1952817|T201|OSN|47586-3|LNC|C-peptide|C-peptide
C1952817|T201|MTH_LN|47586-3|LNC|C-peptide|C-peptide
C1952817|T201|LC|47586-3|LNC|C-peptide|C-peptide
C1952817|T201|LN|47586-3|LNC|C peptide|C peptide
C1952817|T201|OSN|47586-3|LNC|C peptide|C peptide
C1952817|T201|MTH_LN|47586-3|LNC|C peptide|C peptide
C1952817|T201|LC|47586-3|LNC|C peptide|C peptide
C1952818|T201|LN|47587-1|LNC|C-peptide|C-peptide
C1952818|T201|OSN|47587-1|LNC|C-peptide|C-peptide
C1952818|T201|MTH_LN|47587-1|LNC|C-peptide|C-peptide
C1952818|T201|LC|47587-1|LNC|C-peptide|C-peptide
C1952818|T201|LN|47587-1|LNC|C peptide|C peptide
C1952818|T201|OSN|47587-1|LNC|C peptide|C peptide
C1952818|T201|MTH_LN|47587-1|LNC|C peptide|C peptide
C1952818|T201|LC|47587-1|LNC|C peptide|C peptide
C1952819|T201|LN|47588-9|LNC|C-peptide|C-peptide
C1952819|T201|MTH_LN|47588-9|LNC|C-peptide|C-peptide
C1952819|T201|OSN|47588-9|LNC|C-peptide|C-peptide
C1952819|T201|LC|47588-9|LNC|C-peptide|C-peptide
C1952819|T201|LN|47588-9|LNC|C peptide|C peptide
C1952819|T201|MTH_LN|47588-9|LNC|C peptide|C peptide
C1952819|T201|OSN|47588-9|LNC|C peptide|C peptide
C1952819|T201|LC|47588-9|LNC|C peptide|C peptide
C1952820|T201|LN|47589-7|LNC|C-peptide|C-peptide
C1952820|T201|MTH_LN|47589-7|LNC|C-peptide|C-peptide
C1952820|T201|OSN|47589-7|LNC|C-peptide|C-peptide
C1952820|T201|LC|47589-7|LNC|C-peptide|C-peptide
C1952820|T201|LN|47589-7|LNC|C peptide|C peptide
C1952820|T201|MTH_LN|47589-7|LNC|C peptide|C peptide
C1952820|T201|OSN|47589-7|LNC|C peptide|C peptide
C1952820|T201|LC|47589-7|LNC|C peptide|C peptide
C1952821|T201|LN|47590-5|LNC|C-peptide|C-peptide
C1952821|T201|OSN|47590-5|LNC|C-peptide|C-peptide
C1952821|T201|MTH_LN|47590-5|LNC|C-peptide|C-peptide
C1952821|T201|LC|47590-5|LNC|C-peptide|C-peptide
C1952821|T201|LN|47590-5|LNC|C peptide|C peptide
C1952821|T201|OSN|47590-5|LNC|C peptide|C peptide
C1952821|T201|MTH_LN|47590-5|LNC|C peptide|C peptide
C1952821|T201|LC|47590-5|LNC|C peptide|C peptide
C1952822|T201|LN|47591-3|LNC|C-peptide|C-peptide
C1952822|T201|MTH_LN|47591-3|LNC|C-peptide|C-peptide
C1952822|T201|OSN|47591-3|LNC|C-peptide|C-peptide
C1952822|T201|LC|47591-3|LNC|C-peptide|C-peptide
C1952822|T201|LN|47591-3|LNC|C peptide|C peptide
C1952822|T201|MTH_LN|47591-3|LNC|C peptide|C peptide
C1952822|T201|OSN|47591-3|LNC|C peptide|C peptide
C1952822|T201|LC|47591-3|LNC|C peptide|C peptide
C1952823|T201|LN|47592-1|LNC|C-peptide|C-peptide
C1952823|T201|MTH_LN|47592-1|LNC|C-peptide|C-peptide
C1952823|T201|OSN|47592-1|LNC|C-peptide|C-peptide
C1952823|T201|LC|47592-1|LNC|C-peptide|C-peptide
C1952823|T201|LN|47592-1|LNC|C peptide|C peptide
C1952823|T201|MTH_LN|47592-1|LNC|C peptide|C peptide
C1952823|T201|OSN|47592-1|LNC|C peptide|C peptide
C1952823|T201|LC|47592-1|LNC|C peptide|C peptide
C1952824|T201|LN|47593-9|LNC|C-peptide|C-peptide
C1952824|T201|OSN|47593-9|LNC|C-peptide|C-peptide
C1952824|T201|MTH_LN|47593-9|LNC|C-peptide|C-peptide
C1952824|T201|LC|47593-9|LNC|C-peptide|C-peptide
C1952824|T201|LN|47593-9|LNC|C peptide|C peptide
C1952824|T201|OSN|47593-9|LNC|C peptide|C peptide
C1952824|T201|MTH_LN|47593-9|LNC|C peptide|C peptide
C1952824|T201|LC|47593-9|LNC|C peptide|C peptide
C1952825|T201|LN|47594-7|LNC|C-peptide|C-peptide
C1952825|T201|MTH_LN|47594-7|LNC|C-peptide|C-peptide
C1952825|T201|OSN|47594-7|LNC|C-peptide|C-peptide
C1952825|T201|LC|47594-7|LNC|C-peptide|C-peptide
C1952825|T201|LN|47594-7|LNC|C peptide|C peptide
C1952825|T201|MTH_LN|47594-7|LNC|C peptide|C peptide
C1952825|T201|OSN|47594-7|LNC|C peptide|C peptide
C1952825|T201|LC|47594-7|LNC|C peptide|C peptide
C1952826|T201|LN|47595-4|LNC|C-peptide|C-peptide
C1952826|T201|OSN|47595-4|LNC|C-peptide|C-peptide
C1952826|T201|MTH_LN|47595-4|LNC|C-peptide|C-peptide
C1952826|T201|LC|47595-4|LNC|C-peptide|C-peptide
C1952826|T201|LN|47595-4|LNC|C peptide|C peptide
C1952826|T201|OSN|47595-4|LNC|C peptide|C peptide
C1952826|T201|MTH_LN|47595-4|LNC|C peptide|C peptide
C1952826|T201|LC|47595-4|LNC|C peptide|C peptide
C1952827|T201|LN|47596-2|LNC|calcium|calcium
C1952827|T201|OSN|47596-2|LNC|calcium|calcium
C1952827|T201|MTH_LN|47596-2|LNC|calcium|calcium
C1952827|T201|LC|47596-2|LNC|calcium|calcium
C1952827|T201|LN|47596-2|LNC|calcium homeostasis|calcium homeostasis
C1952827|T201|OSN|47596-2|LNC|calcium homeostasis|calcium homeostasis
C1952827|T201|MTH_LN|47596-2|LNC|calcium homeostasis|calcium homeostasis
C1952827|T201|LC|47596-2|LNC|calcium homeostasis|calcium homeostasis
C1952828|T201|LN|47597-0|LNC|calcium|calcium
C1952828|T201|OSN|47597-0|LNC|calcium|calcium
C1952828|T201|MTH_LN|47597-0|LNC|calcium|calcium
C1952828|T201|LC|47597-0|LNC|calcium|calcium
C1952828|T201|LN|47597-0|LNC|calcium homeostasis|calcium homeostasis
C1952828|T201|OSN|47597-0|LNC|calcium homeostasis|calcium homeostasis
C1952828|T201|MTH_LN|47597-0|LNC|calcium homeostasis|calcium homeostasis
C1952828|T201|LC|47597-0|LNC|calcium homeostasis|calcium homeostasis
C1952829|T201|LN|47598-8|LNC|calcium|calcium
C1952829|T201|OSN|47598-8|LNC|calcium|calcium
C1952829|T201|MTH_LN|47598-8|LNC|calcium|calcium
C1952829|T201|LC|47598-8|LNC|calcium|calcium
C1952829|T201|LN|47598-8|LNC|calcium homeostasis|calcium homeostasis
C1952829|T201|OSN|47598-8|LNC|calcium homeostasis|calcium homeostasis
C1952829|T201|MTH_LN|47598-8|LNC|calcium homeostasis|calcium homeostasis
C1952829|T201|LC|47598-8|LNC|calcium homeostasis|calcium homeostasis
C1952839|T201|LN|47608-5|LNC|cortisol|cortisol
C1952839|T201|OSN|47608-5|LNC|cortisol|cortisol
C1952839|T201|MTH_LN|47608-5|LNC|cortisol|cortisol
C1952839|T201|LC|47608-5|LNC|cortisol|cortisol
C1952839|T201|LN|47608-5|LNC|cortisol low|cortisol low
C1952839|T201|OSN|47608-5|LNC|cortisol low|cortisol low
C1952839|T201|MTH_LN|47608-5|LNC|cortisol low|cortisol low
C1952839|T201|LC|47608-5|LNC|cortisol low|cortisol low
C1952839|T201|LN|47608-5|LNC|to undetectable cortisol|to undetectable cortisol
C1952839|T201|OSN|47608-5|LNC|to undetectable cortisol|to undetectable cortisol
C1952839|T201|MTH_LN|47608-5|LNC|to undetectable cortisol|to undetectable cortisol
C1952839|T201|LC|47608-5|LNC|to undetectable cortisol|to undetectable cortisol
C1952877|T201|LN|47640-8|LNC|hematocrit|hematocrit
C1952877|T201|MTH_LN|47640-8|LNC|hematocrit|hematocrit
C1952877|T201|LC|47640-8|LNC|hematocrit|hematocrit
C1952877|T201|OSN|47640-8|LNC|hematocrit|hematocrit
C1952922|T201|LN|47687-9|LNC|luteinizing|luteinizing
C1952922|T201|OSN|47687-9|LNC|luteinizing|luteinizing
C1952922|T201|MTH_LN|47687-9|LNC|luteinizing|luteinizing
C1952922|T201|LC|47687-9|LNC|luteinizing|luteinizing
C1952922|T201|LN|47687-9|LNC|LH|LH
C1952922|T201|OSN|47687-9|LNC|LH|LH
C1952922|T201|MTH_LN|47687-9|LNC|LH|LH
C1952922|T201|LC|47687-9|LNC|LH|LH
C1952922|T201|LN|47687-9|LNC|luteinising|luteinising
C1952922|T201|OSN|47687-9|LNC|luteinising|luteinising
C1952922|T201|MTH_LN|47687-9|LNC|luteinising|luteinising
C1952922|T201|LC|47687-9|LNC|luteinising|luteinising
C1952923|T201|LN|47688-7|LNC|luteinizing|luteinizing
C1952923|T201|OSN|47688-7|LNC|luteinizing|luteinizing
C1952923|T201|MTH_LN|47688-7|LNC|luteinizing|luteinizing
C1952923|T201|LC|47688-7|LNC|luteinizing|luteinizing
C1952923|T201|LN|47688-7|LNC|LH|LH
C1952923|T201|OSN|47688-7|LNC|LH|LH
C1952923|T201|MTH_LN|47688-7|LNC|LH|LH
C1952923|T201|LC|47688-7|LNC|LH|LH
C1952923|T201|LN|47688-7|LNC|luteinising|luteinising
C1952923|T201|OSN|47688-7|LNC|luteinising|luteinising
C1952923|T201|MTH_LN|47688-7|LNC|luteinising|luteinising
C1952923|T201|LC|47688-7|LNC|luteinising|luteinising
C1953159|T201|LN|47832-1|LNC|C-peptide|C-peptide
C1953159|T201|MTH_LN|47832-1|LNC|C-peptide|C-peptide
C1953159|T201|OSN|47832-1|LNC|C-peptide|C-peptide
C1953159|T201|LC|47832-1|LNC|C-peptide|C-peptide
C1953159|T201|LN|47832-1|LNC|C peptide|C peptide
C1953159|T201|MTH_LN|47832-1|LNC|C peptide|C peptide
C1953159|T201|OSN|47832-1|LNC|C peptide|C peptide
C1953159|T201|LC|47832-1|LNC|C peptide|C peptide
C1953160|T201|LN|47833-9|LNC|C-peptide|C-peptide
C1953160|T201|MTH_LN|47833-9|LNC|C-peptide|C-peptide
C1953160|T201|OSN|47833-9|LNC|C-peptide|C-peptide
C1953160|T201|LC|47833-9|LNC|C-peptide|C-peptide
C1953160|T201|LN|47833-9|LNC|C peptide|C peptide
C1953160|T201|MTH_LN|47833-9|LNC|C peptide|C peptide
C1953160|T201|OSN|47833-9|LNC|C peptide|C peptide
C1953160|T201|LC|47833-9|LNC|C peptide|C peptide
C1953161|T201|LN|47834-7|LNC|C-peptide|C-peptide
C1953161|T201|OSN|47834-7|LNC|C-peptide|C-peptide
C1953161|T201|MTH_LN|47834-7|LNC|C-peptide|C-peptide
C1953161|T201|LC|47834-7|LNC|C-peptide|C-peptide
C1953161|T201|LN|47834-7|LNC|C peptide|C peptide
C1953161|T201|OSN|47834-7|LNC|C peptide|C peptide
C1953161|T201|MTH_LN|47834-7|LNC|C peptide|C peptide
C1953161|T201|LC|47834-7|LNC|C peptide|C peptide
C1953170|T201|LN|47850-3|LNC|cortisol|cortisol
C1953170|T201|MTH_LN|47850-3|LNC|cortisol|cortisol
C1953170|T201|OSN|47850-3|LNC|cortisol|cortisol
C1953170|T201|LC|47850-3|LNC|cortisol|cortisol
C1953170|T201|LN|47850-3|LNC|cortisol low|cortisol low
C1953170|T201|MTH_LN|47850-3|LNC|cortisol low|cortisol low
C1953170|T201|OSN|47850-3|LNC|cortisol low|cortisol low
C1953170|T201|LC|47850-3|LNC|cortisol low|cortisol low
C1953170|T201|LN|47850-3|LNC|to undetectable cortisol|to undetectable cortisol
C1953170|T201|MTH_LN|47850-3|LNC|to undetectable cortisol|to undetectable cortisol
C1953170|T201|OSN|47850-3|LNC|to undetectable cortisol|to undetectable cortisol
C1953170|T201|LC|47850-3|LNC|to undetectable cortisol|to undetectable cortisol
C1953186|T201|LN|47864-4|LNC|luteinizing|luteinizing
C1953186|T201|MTH_LN|47864-4|LNC|luteinizing|luteinizing
C1953186|T201|OSN|47864-4|LNC|luteinizing|luteinizing
C1953186|T201|LC|47864-4|LNC|luteinizing|luteinizing
C1953186|T201|LN|47864-4|LNC|LH|LH
C1953186|T201|MTH_LN|47864-4|LNC|LH|LH
C1953186|T201|OSN|47864-4|LNC|LH|LH
C1953186|T201|LC|47864-4|LNC|LH|LH
C1953186|T201|LN|47864-4|LNC|luteinising|luteinising
C1953186|T201|MTH_LN|47864-4|LNC|luteinising|luteinising
C1953186|T201|OSN|47864-4|LNC|luteinising|luteinising
C1953186|T201|LC|47864-4|LNC|luteinising|luteinising
C1953264|T201|LN|47941-0|LNC|androgen|androgen
C1953264|T201|OSN|47941-0|LNC|androgen|androgen
C1953264|T201|MTH_LN|47941-0|LNC|androgen|androgen
C1953264|T201|LC|47941-0|LNC|androgen|androgen
C1953269|T201|LN|47946-9|LNC|androgen|androgen
C1953269|T201|OSN|47946-9|LNC|androgen|androgen
C1953269|T201|MTH_LN|47946-9|LNC|androgen|androgen
C1953269|T201|LC|47946-9|LNC|androgen|androgen
C1953449|T201|LN|48065-7|LNC|coagulation disorder|coagulation disorder
C1953449|T201|OSN|48065-7|LNC|coagulation disorder|coagulation disorder
C1953449|T201|MTH_LN|48065-7|LNC|coagulation disorder|coagulation disorder
C1953449|T201|LC|48065-7|LNC|coagulation disorder|coagulation disorder
C1953449|T201|LN|48065-7|LNC|coagulation|coagulation
C1953449|T201|OSN|48065-7|LNC|coagulation|coagulation
C1953449|T201|MTH_LN|48065-7|LNC|coagulation|coagulation
C1953449|T201|LC|48065-7|LNC|coagulation|coagulation
C1953449|T201|LN|48065-7|LNC|Coagulationities|Coagulationities
C1953449|T201|OSN|48065-7|LNC|Coagulationities|Coagulationities
C1953449|T201|MTH_LN|48065-7|LNC|Coagulationities|Coagulationities
C1953449|T201|LC|48065-7|LNC|Coagulationities|Coagulationities
C1953449|T201|LN|48065-7|LNC|coagulation studies|coagulation studies
C1953449|T201|OSN|48065-7|LNC|coagulation studies|coagulation studies
C1953449|T201|MTH_LN|48065-7|LNC|coagulation studies|coagulation studies
C1953449|T201|LC|48065-7|LNC|coagulation studies|coagulation studies
C1953449|T201|LN|48065-7|LNC|clotting|clotting
C1953449|T201|OSN|48065-7|LNC|clotting|clotting
C1953449|T201|MTH_LN|48065-7|LNC|clotting|clotting
C1953449|T201|LC|48065-7|LNC|clotting|clotting
C1953490|T201|LN|48090-5|LNC|HDL cholesterol|HDL cholesterol
C1953490|T201|OSN|48090-5|LNC|HDL cholesterol|HDL cholesterol
C1953490|T201|MTH_LN|48090-5|LNC|HDL cholesterol|HDL cholesterol
C1953490|T201|LC|48090-5|LNC|HDL cholesterol|HDL cholesterol
C1953490|T201|LN|48090-5|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1953490|T201|OSN|48090-5|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1953490|T201|MTH_LN|48090-5|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1953490|T201|LC|48090-5|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1953490|T201|LN|48090-5|LNC|HDL-cholesterol|HDL-cholesterol
C1953490|T201|OSN|48090-5|LNC|HDL-cholesterol|HDL-cholesterol
C1953490|T201|MTH_LN|48090-5|LNC|HDL-cholesterol|HDL-cholesterol
C1953490|T201|LC|48090-5|LNC|HDL-cholesterol|HDL-cholesterol
C1953490|T201|LN|48090-5|LNC|high-density lipoprotein|high-density lipoprotein
C1953490|T201|OSN|48090-5|LNC|high-density lipoprotein|high-density lipoprotein
C1953490|T201|MTH_LN|48090-5|LNC|high-density lipoprotein|high-density lipoprotein
C1953490|T201|LC|48090-5|LNC|high-density lipoprotein|high-density lipoprotein
C1953490|T201|LN|48090-5|LNC|HDL|HDL
C1953490|T201|OSN|48090-5|LNC|HDL|HDL
C1953490|T201|MTH_LN|48090-5|LNC|HDL|HDL
C1953490|T201|LC|48090-5|LNC|HDL|HDL
C1953492|T201|LN|48091-3|LNC|ACTH|ACTH
C1953492|T201|MTH_LN|48091-3|LNC|ACTH|ACTH
C1953492|T201|OSN|48091-3|LNC|ACTH|ACTH
C1953492|T201|LC|48091-3|LNC|ACTH|ACTH
C1953492|T201|LN|48091-3|LNC|corticotropin|corticotropin
C1953492|T201|MTH_LN|48091-3|LNC|corticotropin|corticotropin
C1953492|T201|OSN|48091-3|LNC|corticotropin|corticotropin
C1953492|T201|LC|48091-3|LNC|corticotropin|corticotropin
// C1953492|T201|LN|48091-3|LNC||
// C1953492|T201|MTH_LN|48091-3|LNC||
// C1953492|T201|OSN|48091-3|LNC||
// C1953492|T201|LC|48091-3|LNC||
C1953493|T201|LN|48092-1|LNC|ACTH|ACTH
C1953493|T201|OSN|48092-1|LNC|ACTH|ACTH
C1953493|T201|MTH_LN|48092-1|LNC|ACTH|ACTH
C1953493|T201|LC|48092-1|LNC|ACTH|ACTH
C1953493|T201|LN|48092-1|LNC|corticotropin|corticotropin
C1953493|T201|OSN|48092-1|LNC|corticotropin|corticotropin
C1953493|T201|MTH_LN|48092-1|LNC|corticotropin|corticotropin
C1953493|T201|LC|48092-1|LNC|corticotropin|corticotropin
// C1953493|T201|LN|48092-1|LNC||
// C1953493|T201|OSN|48092-1|LNC||
// C1953493|T201|MTH_LN|48092-1|LNC||
// C1953493|T201|LC|48092-1|LNC||
C1953494|T201|LN|48093-9|LNC|ACTH|ACTH
C1953494|T201|MTH_LN|48093-9|LNC|ACTH|ACTH
C1953494|T201|OSN|48093-9|LNC|ACTH|ACTH
C1953494|T201|LC|48093-9|LNC|ACTH|ACTH
C1953494|T201|LN|48093-9|LNC|corticotropin|corticotropin
C1953494|T201|MTH_LN|48093-9|LNC|corticotropin|corticotropin
C1953494|T201|OSN|48093-9|LNC|corticotropin|corticotropin
C1953494|T201|LC|48093-9|LNC|corticotropin|corticotropin
// C1953494|T201|LN|48093-9|LNC||
// C1953494|T201|MTH_LN|48093-9|LNC||
// C1953494|T201|OSN|48093-9|LNC||
// C1953494|T201|LC|48093-9|LNC||
C1953495|T201|LN|48094-7|LNC|ACTH|ACTH
C1953495|T201|OSN|48094-7|LNC|ACTH|ACTH
C1953495|T201|MTH_LN|48094-7|LNC|ACTH|ACTH
C1953495|T201|LC|48094-7|LNC|ACTH|ACTH
C1953495|T201|LN|48094-7|LNC|corticotropin|corticotropin
C1953495|T201|OSN|48094-7|LNC|corticotropin|corticotropin
C1953495|T201|MTH_LN|48094-7|LNC|corticotropin|corticotropin
C1953495|T201|LC|48094-7|LNC|corticotropin|corticotropin
// C1953495|T201|LN|48094-7|LNC||
// C1953495|T201|OSN|48094-7|LNC||
// C1953495|T201|MTH_LN|48094-7|LNC||
// C1953495|T201|LC|48094-7|LNC||
C1953496|T201|LN|48095-4|LNC|ACTH|ACTH
C1953496|T201|MTH_LN|48095-4|LNC|ACTH|ACTH
C1953496|T201|OSN|48095-4|LNC|ACTH|ACTH
C1953496|T201|LC|48095-4|LNC|ACTH|ACTH
C1953496|T201|LN|48095-4|LNC|corticotropin|corticotropin
C1953496|T201|MTH_LN|48095-4|LNC|corticotropin|corticotropin
C1953496|T201|OSN|48095-4|LNC|corticotropin|corticotropin
C1953496|T201|LC|48095-4|LNC|corticotropin|corticotropin
// C1953496|T201|LN|48095-4|LNC||
// C1953496|T201|MTH_LN|48095-4|LNC||
// C1953496|T201|OSN|48095-4|LNC||
// C1953496|T201|LC|48095-4|LNC||
C1953497|T201|LN|48096-2|LNC|ACTH|ACTH
C1953497|T201|OSN|48096-2|LNC|ACTH|ACTH
C1953497|T201|MTH_LN|48096-2|LNC|ACTH|ACTH
C1953497|T201|LC|48096-2|LNC|ACTH|ACTH
C1953497|T201|LN|48096-2|LNC|corticotropin|corticotropin
C1953497|T201|OSN|48096-2|LNC|corticotropin|corticotropin
C1953497|T201|MTH_LN|48096-2|LNC|corticotropin|corticotropin
C1953497|T201|LC|48096-2|LNC|corticotropin|corticotropin
// C1953497|T201|LN|48096-2|LNC||
// C1953497|T201|OSN|48096-2|LNC||
// C1953497|T201|MTH_LN|48096-2|LNC||
// C1953497|T201|LC|48096-2|LNC||
C1953498|T201|LN|48097-0|LNC|ACTH|ACTH
C1953498|T201|MTH_LN|48097-0|LNC|ACTH|ACTH
C1953498|T201|OSN|48097-0|LNC|ACTH|ACTH
C1953498|T201|LC|48097-0|LNC|ACTH|ACTH
C1953498|T201|LN|48097-0|LNC|corticotropin|corticotropin
C1953498|T201|MTH_LN|48097-0|LNC|corticotropin|corticotropin
C1953498|T201|OSN|48097-0|LNC|corticotropin|corticotropin
C1953498|T201|LC|48097-0|LNC|corticotropin|corticotropin
// C1953498|T201|LN|48097-0|LNC||
// C1953498|T201|MTH_LN|48097-0|LNC||
// C1953498|T201|OSN|48097-0|LNC||
// C1953498|T201|LC|48097-0|LNC||
C1953526|T201|LN|48118-4|LNC|luteinizing|luteinizing
C1953526|T201|MTH_LN|48118-4|LNC|luteinizing|luteinizing
C1953526|T201|OSN|48118-4|LNC|luteinizing|luteinizing
C1953526|T201|LC|48118-4|LNC|luteinizing|luteinizing
C1953526|T201|LN|48118-4|LNC|LH|LH
C1953526|T201|MTH_LN|48118-4|LNC|LH|LH
C1953526|T201|OSN|48118-4|LNC|LH|LH
C1953526|T201|LC|48118-4|LNC|LH|LH
C1953526|T201|LN|48118-4|LNC|luteinising|luteinising
C1953526|T201|MTH_LN|48118-4|LNC|luteinising|luteinising
C1953526|T201|OSN|48118-4|LNC|luteinising|luteinising
C1953526|T201|LC|48118-4|LNC|luteinising|luteinising
C1953928|T201|LN|48425-3|LNC|troponin T|troponin T
C1953928|T201|MTH_LN|48425-3|LNC|troponin T|troponin T
C1953928|T201|OSN|48425-3|LNC|troponin T|troponin T
C1953928|T201|LC|48425-3|LNC|troponin T|troponin T
C1953929|T201|LN|48426-1|LNC|troponin T|troponin T
C1953929|T201|MTH_LN|48426-1|LNC|troponin T|troponin T
C1953929|T201|OSN|48426-1|LNC|troponin T|troponin T
C1953929|T201|LC|48426-1|LNC|troponin T|troponin T
C1954149|T201|LN|48581-3|LNC|luteinizing|luteinizing
C1954149|T201|MTH_LN|48581-3|LNC|luteinizing|luteinizing
C1954149|T201|OSN|48581-3|LNC|luteinizing|luteinizing
C1954149|T201|LC|48581-3|LNC|luteinizing|luteinizing
C1954149|T201|LN|48581-3|LNC|LH|LH
C1954149|T201|MTH_LN|48581-3|LNC|LH|LH
C1954149|T201|OSN|48581-3|LNC|LH|LH
C1954149|T201|LC|48581-3|LNC|LH|LH
C1954149|T201|LN|48581-3|LNC|luteinising|luteinising
C1954149|T201|MTH_LN|48581-3|LNC|luteinising|luteinising
C1954149|T201|OSN|48581-3|LNC|luteinising|luteinising
C1954149|T201|LC|48581-3|LNC|luteinising|luteinising
C1954150|T201|LN|48582-1|LNC|luteinizing|luteinizing
C1954150|T201|MTH_LN|48582-1|LNC|luteinizing|luteinizing
C1954150|T201|OSN|48582-1|LNC|luteinizing|luteinizing
C1954150|T201|LC|48582-1|LNC|luteinizing|luteinizing
C1954150|T201|LN|48582-1|LNC|LH|LH
C1954150|T201|MTH_LN|48582-1|LNC|LH|LH
C1954150|T201|OSN|48582-1|LNC|LH|LH
C1954150|T201|LC|48582-1|LNC|LH|LH
C1954150|T201|LN|48582-1|LNC|luteinising|luteinising
C1954150|T201|MTH_LN|48582-1|LNC|luteinising|luteinising
C1954150|T201|OSN|48582-1|LNC|luteinising|luteinising
C1954150|T201|LC|48582-1|LNC|luteinising|luteinising
C1954151|T201|LN|48583-9|LNC|luteinizing|luteinizing
C1954151|T201|MTH_LN|48583-9|LNC|luteinizing|luteinizing
C1954151|T201|OSN|48583-9|LNC|luteinizing|luteinizing
C1954151|T201|LC|48583-9|LNC|luteinizing|luteinizing
C1954151|T201|LN|48583-9|LNC|LH|LH
C1954151|T201|MTH_LN|48583-9|LNC|LH|LH
C1954151|T201|OSN|48583-9|LNC|LH|LH
C1954151|T201|LC|48583-9|LNC|LH|LH
C1954151|T201|LN|48583-9|LNC|luteinising|luteinising
C1954151|T201|MTH_LN|48583-9|LNC|luteinising|luteinising
C1954151|T201|OSN|48583-9|LNC|luteinising|luteinising
C1954151|T201|LC|48583-9|LNC|luteinising|luteinising
C1954199|T201|LN|48618-3|LNC|VLDL cholesterol|VLDL cholesterol
C1954199|T201|OSN|48618-3|LNC|VLDL cholesterol|VLDL cholesterol
C1954199|T201|MTH_LN|48618-3|LNC|VLDL cholesterol|VLDL cholesterol
C1954199|T201|LC|48618-3|LNC|VLDL cholesterol|VLDL cholesterol
C1954199|T201|LN|48618-3|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1954199|T201|OSN|48618-3|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1954199|T201|MTH_LN|48618-3|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1954199|T201|LC|48618-3|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1954199|T201|LN|48618-3|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1954199|T201|OSN|48618-3|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1954199|T201|MTH_LN|48618-3|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1954199|T201|LC|48618-3|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1954228|T201|LN|48642-3|LNC|glomerular filtration rate|glomerular filtration rate
C1954228|T201|LC|48642-3|LNC|glomerular filtration rate|glomerular filtration rate
C1954228|T201|OSN|48642-3|LNC|glomerular filtration rate|glomerular filtration rate
C1954228|T201|MTH_LN|48642-3|LNC|glomerular filtration rate|glomerular filtration rate
C1954228|T201|LN|48642-3|LNC|creatinine clearance|creatinine clearance
C1954228|T201|LC|48642-3|LNC|creatinine clearance|creatinine clearance
C1954228|T201|OSN|48642-3|LNC|creatinine clearance|creatinine clearance
C1954228|T201|MTH_LN|48642-3|LNC|creatinine clearance|creatinine clearance
C1954230|T201|LN|48643-1|LNC|glomerular filtration rate|glomerular filtration rate
C1954230|T201|MTH_LN|48643-1|LNC|glomerular filtration rate|glomerular filtration rate
C1954230|T201|LC|48643-1|LNC|glomerular filtration rate|glomerular filtration rate
C1954230|T201|OSN|48643-1|LNC|glomerular filtration rate|glomerular filtration rate
C1954230|T201|LN|48643-1|LNC|creatinine clearance|creatinine clearance
C1954230|T201|MTH_LN|48643-1|LNC|creatinine clearance|creatinine clearance
C1954230|T201|LC|48643-1|LNC|creatinine clearance|creatinine clearance
C1954230|T201|OSN|48643-1|LNC|creatinine clearance|creatinine clearance
C1954256|T201|LN|48660-5|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1954256|T201|OSN|48660-5|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1954256|T201|MTH_LN|48660-5|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1954256|T201|LC|48660-5|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1954321|T201|LN|48703-3|LNC|hematocrit|hematocrit
C1954321|T201|MTH_LN|48703-3|LNC|hematocrit|hematocrit
C1954321|T201|LC|48703-3|LNC|hematocrit|hematocrit
C1954321|T201|OSN|48703-3|LNC|hematocrit|hematocrit
C1954746|T201|LN|49026-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954746|T201|MTH_LN|49026-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954746|T201|LC|49026-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954746|T201|OSN|49026-8|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954746|T201|LN|49026-8|LNC|LDL|LDL
C1954746|T201|MTH_LN|49026-8|LNC|LDL|LDL
C1954746|T201|LC|49026-8|LNC|LDL|LDL
C1954746|T201|OSN|49026-8|LNC|LDL|LDL
C1954746|T201|LN|49026-8|LNC|LDL cholesterol|LDL cholesterol
C1954746|T201|MTH_LN|49026-8|LNC|LDL cholesterol|LDL cholesterol
C1954746|T201|LC|49026-8|LNC|LDL cholesterol|LDL cholesterol
C1954746|T201|OSN|49026-8|LNC|LDL cholesterol|LDL cholesterol
C1954746|T201|LN|49026-8|LNC|low-density lipoprotein|low-density lipoprotein
C1954746|T201|MTH_LN|49026-8|LNC|low-density lipoprotein|low-density lipoprotein
C1954746|T201|LC|49026-8|LNC|low-density lipoprotein|low-density lipoprotein
C1954746|T201|OSN|49026-8|LNC|low-density lipoprotein|low-density lipoprotein
C1954746|T201|LN|49026-8|LNC|beta-lipoproteins|beta-lipoproteins
C1954746|T201|MTH_LN|49026-8|LNC|beta-lipoproteins|beta-lipoproteins
C1954746|T201|LC|49026-8|LNC|beta-lipoproteins|beta-lipoproteins
C1954746|T201|OSN|49026-8|LNC|beta-lipoproteins|beta-lipoproteins
C1954746|T201|LN|49026-8|LNC|LDL-C|LDL-C
C1954746|T201|MTH_LN|49026-8|LNC|LDL-C|LDL-C
C1954746|T201|LC|49026-8|LNC|LDL-C|LDL-C
C1954746|T201|OSN|49026-8|LNC|LDL-C|LDL-C
C1954748|T201|LN|49027-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954748|T201|MTH_LN|49027-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954748|T201|OSN|49027-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954748|T201|LC|49027-6|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954748|T201|LN|49027-6|LNC|LDL|LDL
C1954748|T201|MTH_LN|49027-6|LNC|LDL|LDL
C1954748|T201|OSN|49027-6|LNC|LDL|LDL
C1954748|T201|LC|49027-6|LNC|LDL|LDL
C1954748|T201|LN|49027-6|LNC|LDL cholesterol|LDL cholesterol
C1954748|T201|MTH_LN|49027-6|LNC|LDL cholesterol|LDL cholesterol
C1954748|T201|OSN|49027-6|LNC|LDL cholesterol|LDL cholesterol
C1954748|T201|LC|49027-6|LNC|LDL cholesterol|LDL cholesterol
C1954748|T201|LN|49027-6|LNC|low-density lipoprotein|low-density lipoprotein
C1954748|T201|MTH_LN|49027-6|LNC|low-density lipoprotein|low-density lipoprotein
C1954748|T201|OSN|49027-6|LNC|low-density lipoprotein|low-density lipoprotein
C1954748|T201|LC|49027-6|LNC|low-density lipoprotein|low-density lipoprotein
C1954748|T201|LN|49027-6|LNC|beta-lipoproteins|beta-lipoproteins
C1954748|T201|MTH_LN|49027-6|LNC|beta-lipoproteins|beta-lipoproteins
C1954748|T201|OSN|49027-6|LNC|beta-lipoproteins|beta-lipoproteins
C1954748|T201|LC|49027-6|LNC|beta-lipoproteins|beta-lipoproteins
C1954748|T201|LN|49027-6|LNC|LDL-C|LDL-C
C1954748|T201|MTH_LN|49027-6|LNC|LDL-C|LDL-C
C1954748|T201|OSN|49027-6|LNC|LDL-C|LDL-C
C1954748|T201|LC|49027-6|LNC|LDL-C|LDL-C
C1954793|T201|LN|49054-0|LNC|vitamin D metabolism|vitamin D metabolism
C1954793|T201|MTH_LN|49054-0|LNC|vitamin D metabolism|vitamin D metabolism
C1954793|T201|LC|49054-0|LNC|vitamin D metabolism|vitamin D metabolism
C1954793|T201|OSN|49054-0|LNC|vitamin D metabolism|vitamin D metabolism
C1954793|T201|LN|49054-0|LNC|calcifediol|calcifediol
C1954793|T201|MTH_LN|49054-0|LNC|calcifediol|calcifediol
C1954793|T201|LC|49054-0|LNC|calcifediol|calcifediol
C1954793|T201|OSN|49054-0|LNC|calcifediol|calcifediol
C1954793|T201|LN|49054-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1954793|T201|MTH_LN|49054-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1954793|T201|LC|49054-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1954793|T201|OSN|49054-0|LNC|25-hydroxycholecalciferol|25-hydroxycholecalciferol
C1954793|T201|LN|49054-0|LNC|calcidiol|calcidiol
C1954793|T201|MTH_LN|49054-0|LNC|calcidiol|calcidiol
C1954793|T201|LC|49054-0|LNC|calcidiol|calcidiol
C1954793|T201|OSN|49054-0|LNC|calcidiol|calcidiol
C1954893|T201|LN|49130-8|LNC|HDL cholesterol|HDL cholesterol
C1954893|T201|MTH_LN|49130-8|LNC|HDL cholesterol|HDL cholesterol
C1954893|T201|OSN|49130-8|LNC|HDL cholesterol|HDL cholesterol
C1954893|T201|LC|49130-8|LNC|HDL cholesterol|HDL cholesterol
C1954893|T201|LN|49130-8|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1954893|T201|MTH_LN|49130-8|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1954893|T201|OSN|49130-8|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1954893|T201|LC|49130-8|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C1954893|T201|LN|49130-8|LNC|HDL-cholesterol|HDL-cholesterol
C1954893|T201|MTH_LN|49130-8|LNC|HDL-cholesterol|HDL-cholesterol
C1954893|T201|OSN|49130-8|LNC|HDL-cholesterol|HDL-cholesterol
C1954893|T201|LC|49130-8|LNC|HDL-cholesterol|HDL-cholesterol
C1954893|T201|LN|49130-8|LNC|high-density lipoprotein|high-density lipoprotein
C1954893|T201|MTH_LN|49130-8|LNC|high-density lipoprotein|high-density lipoprotein
C1954893|T201|OSN|49130-8|LNC|high-density lipoprotein|high-density lipoprotein
C1954893|T201|LC|49130-8|LNC|high-density lipoprotein|high-density lipoprotein
C1954893|T201|LN|49130-8|LNC|HDL|HDL
C1954893|T201|MTH_LN|49130-8|LNC|HDL|HDL
C1954893|T201|OSN|49130-8|LNC|HDL|HDL
C1954893|T201|LC|49130-8|LNC|HDL|HDL
C1954896|T201|LN|49132-4|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954896|T201|MTH_LN|49132-4|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954896|T201|OSN|49132-4|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954896|T201|LC|49132-4|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C1954896|T201|LN|49132-4|LNC|LDL|LDL
C1954896|T201|MTH_LN|49132-4|LNC|LDL|LDL
C1954896|T201|OSN|49132-4|LNC|LDL|LDL
C1954896|T201|LC|49132-4|LNC|LDL|LDL
C1954896|T201|LN|49132-4|LNC|LDL cholesterol|LDL cholesterol
C1954896|T201|MTH_LN|49132-4|LNC|LDL cholesterol|LDL cholesterol
C1954896|T201|OSN|49132-4|LNC|LDL cholesterol|LDL cholesterol
C1954896|T201|LC|49132-4|LNC|LDL cholesterol|LDL cholesterol
C1954896|T201|LN|49132-4|LNC|low-density lipoprotein|low-density lipoprotein
C1954896|T201|MTH_LN|49132-4|LNC|low-density lipoprotein|low-density lipoprotein
C1954896|T201|OSN|49132-4|LNC|low-density lipoprotein|low-density lipoprotein
C1954896|T201|LC|49132-4|LNC|low-density lipoprotein|low-density lipoprotein
C1954896|T201|LN|49132-4|LNC|beta-lipoproteins|beta-lipoproteins
C1954896|T201|MTH_LN|49132-4|LNC|beta-lipoproteins|beta-lipoproteins
C1954896|T201|OSN|49132-4|LNC|beta-lipoproteins|beta-lipoproteins
C1954896|T201|LC|49132-4|LNC|beta-lipoproteins|beta-lipoproteins
C1954896|T201|LN|49132-4|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1954896|T201|MTH_LN|49132-4|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1954896|T201|OSN|49132-4|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1954896|T201|LC|49132-4|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C1954896|T201|LN|49132-4|LNC|LDL-C|LDL-C
C1954896|T201|MTH_LN|49132-4|LNC|LDL-C|LDL-C
C1954896|T201|OSN|49132-4|LNC|LDL-C|LDL-C
C1954896|T201|LC|49132-4|LNC|LDL-C|LDL-C
C1954897|T201|LN|49133-2|LNC|VLDL cholesterol|VLDL cholesterol
C1954897|T201|OSN|49133-2|LNC|VLDL cholesterol|VLDL cholesterol
C1954897|T201|MTH_LN|49133-2|LNC|VLDL cholesterol|VLDL cholesterol
C1954897|T201|LC|49133-2|LNC|VLDL cholesterol|VLDL cholesterol
C1954897|T201|LN|49133-2|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1954897|T201|OSN|49133-2|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1954897|T201|MTH_LN|49133-2|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1954897|T201|LC|49133-2|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1954897|T201|LN|49133-2|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1954897|T201|OSN|49133-2|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1954897|T201|MTH_LN|49133-2|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1954897|T201|LC|49133-2|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1954901|T201|LN|49137-3|LNC|Hemoglobin|Hemoglobin
C1954901|T201|MTH_LN|49137-3|LNC|Hemoglobin|Hemoglobin
C1954901|T201|OSN|49137-3|LNC|Hemoglobin|Hemoglobin
C1954901|T201|LC|49137-3|LNC|Hemoglobin|Hemoglobin
C1976903|T201|LN|50192-4|LNC|VLDL cholesterol|VLDL cholesterol
C1976903|T201|MTH_LN|50192-4|LNC|VLDL cholesterol|VLDL cholesterol
C1976903|T201|OSN|50192-4|LNC|VLDL cholesterol|VLDL cholesterol
C1976903|T201|LC|50192-4|LNC|VLDL cholesterol|VLDL cholesterol
C1976903|T201|LN|50192-4|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1976903|T201|MTH_LN|50192-4|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1976903|T201|OSN|50192-4|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1976903|T201|LC|50192-4|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1976903|T201|LN|50192-4|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1976903|T201|MTH_LN|50192-4|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1976903|T201|OSN|50192-4|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1976903|T201|LC|50192-4|LNC|very-low-density lipoprotein|very-low-density lipoprotein
// C1977255|T201|LN|49505-1|LNC||
// C1977255|T201|LC|49505-1|LNC||
// C1977255|T201|MTH_LN|49505-1|LNC||
// C1977255|T201|OSN|49505-1|LNC||
C1977255|T201|LN|49505-1|LNC|occult|occult
C1977255|T201|LC|49505-1|LNC|occult|occult
C1977255|T201|MTH_LN|49505-1|LNC|occult|occult
C1977255|T201|OSN|49505-1|LNC|occult|occult
C1977318|T201|LN|49563-0|LNC|troponin I|troponin I
C1977318|T201|MTH_LN|49563-0|LNC|troponin I|troponin I
C1977318|T201|OSN|49563-0|LNC|troponin I|troponin I
C1977318|T201|LC|49563-0|LNC|troponin I|troponin I
C1977402|T201|LN|49624-0|LNC|VLDL cholesterol|VLDL cholesterol
C1977402|T201|OSN|49624-0|LNC|VLDL cholesterol|VLDL cholesterol
C1977402|T201|MTH_LN|49624-0|LNC|VLDL cholesterol|VLDL cholesterol
C1977402|T201|LC|49624-0|LNC|VLDL cholesterol|VLDL cholesterol
C1977402|T201|LN|49624-0|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1977402|T201|OSN|49624-0|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1977402|T201|MTH_LN|49624-0|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1977402|T201|LC|49624-0|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C1977402|T201|LN|49624-0|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1977402|T201|OSN|49624-0|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1977402|T201|MTH_LN|49624-0|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1977402|T201|LC|49624-0|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C1977516|T201|LN|49765-1|LNC|calcium|calcium
C1977516|T201|MTH_LN|49765-1|LNC|calcium|calcium
C1977516|T201|OSN|49765-1|LNC|calcium|calcium
C1977516|T201|LC|49765-1|LNC|calcium|calcium
C1977516|T201|LN|49765-1|LNC|calcium homeostasis|calcium homeostasis
C1977516|T201|MTH_LN|49765-1|LNC|calcium homeostasis|calcium homeostasis
C1977516|T201|OSN|49765-1|LNC|calcium homeostasis|calcium homeostasis
C1977516|T201|LC|49765-1|LNC|calcium homeostasis|calcium homeostasis
C1977524|T201|LN|49781-8|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C1977524|T201|OSN|49781-8|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C1977524|T201|MTH_LN|49781-8|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C1977524|T201|LC|49781-8|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C1977690|T201|LN|50202-1|LNC|iron|iron
C1977690|T201|OSN|50202-1|LNC|iron|iron
C1977690|T201|MTH_LN|50202-1|LNC|iron|iron
C1977690|T201|LC|50202-1|LNC|iron|iron
C1977691|T201|LN|50203-9|LNC|iron|iron
C1977691|T201|OSN|50203-9|LNC|iron|iron
C1977691|T201|MTH_LN|50203-9|LNC|iron|iron
C1977691|T201|LC|50203-9|LNC|iron|iron
C1977692|T201|LN|50204-7|LNC|iron|iron
C1977692|T201|MTH_LN|50204-7|LNC|iron|iron
C1977692|T201|OSN|50204-7|LNC|iron|iron
C1977692|T201|LC|50204-7|LNC|iron|iron
C1977693|T201|LN|50205-4|LNC|iron|iron
C1977693|T201|MTH_LN|50205-4|LNC|iron|iron
C1977693|T201|OSN|50205-4|LNC|iron|iron
C1977693|T201|LC|50205-4|LNC|iron|iron
C1977831|T201|LN|49959-0|LNC|osmolality|osmolality
C1977831|T201|MTH_LN|49959-0|LNC|osmolality|osmolality
C1977831|T201|LC|49959-0|LNC|osmolality|osmolality
C1977831|T201|OSN|49959-0|LNC|osmolality|osmolality
C1977831|T201|LN|49959-0|LNC|homeostasis|homeostasis
C1977831|T201|MTH_LN|49959-0|LNC|homeostasis|homeostasis
C1977831|T201|LC|49959-0|LNC|homeostasis|homeostasis
C1977831|T201|OSN|49959-0|LNC|homeostasis|homeostasis
C1977844|T201|LN|49968-1|LNC|cortisol|cortisol
C1977844|T201|OSN|49968-1|LNC|cortisol|cortisol
C1977844|T201|MTH_LN|49968-1|LNC|cortisol|cortisol
C1977844|T201|LC|49968-1|LNC|cortisol|cortisol
C1977844|T201|LN|49968-1|LNC|cortisol low|cortisol low
C1977844|T201|OSN|49968-1|LNC|cortisol low|cortisol low
C1977844|T201|MTH_LN|49968-1|LNC|cortisol low|cortisol low
C1977844|T201|LC|49968-1|LNC|cortisol low|cortisol low
C1977844|T201|LN|49968-1|LNC|to undetectable cortisol|to undetectable cortisol
C1977844|T201|OSN|49968-1|LNC|to undetectable cortisol|to undetectable cortisol
C1977844|T201|MTH_LN|49968-1|LNC|to undetectable cortisol|to undetectable cortisol
C1977844|T201|LC|49968-1|LNC|to undetectable cortisol|to undetectable cortisol
C1977845|T201|LN|49969-9|LNC|cortisol|cortisol
C1977845|T201|OSN|49969-9|LNC|cortisol|cortisol
C1977845|T201|MTH_LN|49969-9|LNC|cortisol|cortisol
C1977845|T201|LC|49969-9|LNC|cortisol|cortisol
C1977845|T201|LN|49969-9|LNC|cortisol low|cortisol low
C1977845|T201|OSN|49969-9|LNC|cortisol low|cortisol low
C1977845|T201|MTH_LN|49969-9|LNC|cortisol low|cortisol low
C1977845|T201|LC|49969-9|LNC|cortisol low|cortisol low
C1977845|T201|LN|49969-9|LNC|to undetectable cortisol|to undetectable cortisol
C1977845|T201|OSN|49969-9|LNC|to undetectable cortisol|to undetectable cortisol
C1977845|T201|MTH_LN|49969-9|LNC|to undetectable cortisol|to undetectable cortisol
C1977845|T201|LC|49969-9|LNC|to undetectable cortisol|to undetectable cortisol
C1978030|T201|LN|50171-8|LNC|aldosterone|aldosterone
C1978030|T201|OSN|50171-8|LNC|aldosterone|aldosterone
C1978030|T201|MTH_LN|50171-8|LNC|aldosterone|aldosterone
C1978030|T201|LC|50171-8|LNC|aldosterone|aldosterone
C1978031|T201|LN|50172-6|LNC|aldosterone|aldosterone
C1978031|T201|OSN|50172-6|LNC|aldosterone|aldosterone
C1978031|T201|MTH_LN|50172-6|LNC|aldosterone|aldosterone
C1978031|T201|LC|50172-6|LNC|aldosterone|aldosterone
C1978032|T201|LN|50173-4|LNC|aldosterone|aldosterone
C1978032|T201|MTH_LN|50173-4|LNC|aldosterone|aldosterone
C1978032|T201|OSN|50173-4|LNC|aldosterone|aldosterone
C1978032|T201|LC|50173-4|LNC|aldosterone|aldosterone
C1978037|T201|LN|50198-1|LNC|iron|iron
C1978037|T201|OSN|50198-1|LNC|iron|iron
C1978037|T201|MTH_LN|50198-1|LNC|iron|iron
C1978037|T201|LC|50198-1|LNC|iron|iron
C1978038|T201|LN|50199-9|LNC|iron|iron
C1978038|T201|MTH_LN|50199-9|LNC|iron|iron
C1978038|T201|OSN|50199-9|LNC|iron|iron
C1978038|T201|LC|50199-9|LNC|iron|iron
C1978039|T201|LN|50200-5|LNC|iron|iron
C1978039|T201|MTH_LN|50200-5|LNC|iron|iron
C1978039|T201|OSN|50200-5|LNC|iron|iron
C1978039|T201|LC|50200-5|LNC|iron|iron
C1978040|T201|LN|50201-3|LNC|iron|iron
C1978040|T201|OSN|50201-3|LNC|iron|iron
C1978040|T201|MTH_LN|50201-3|LNC|iron|iron
C1978040|T201|LC|50201-3|LNC|iron|iron
// C1978061|T201|LN|50226-0|LNC||
// C1978061|T201|MTH_LN|50226-0|LNC||
// C1978061|T201|OSN|50226-0|LNC||
// C1978061|T201|LC|50226-0|LNC||
C1978061|T201|LN|50226-0|LNC|occult|occult
C1978061|T201|MTH_LN|50226-0|LNC|occult|occult
C1978061|T201|OSN|50226-0|LNC|occult|occult
C1978061|T201|LC|50226-0|LNC|occult|occult
C1978070|T201|LN|50235-1|LNC|homeostasis|homeostasis
C1978070|T201|MTH_LN|50235-1|LNC|homeostasis|homeostasis
C1978070|T201|OSN|50235-1|LNC|homeostasis|homeostasis
C1978070|T201|LC|50235-1|LNC|homeostasis|homeostasis
C1978283|T201|LN|50410-0|LNC|Autoimmune antibody|Autoimmune antibody
C1978283|T201|OSN|50410-0|LNC|Autoimmune antibody|Autoimmune antibody
C1978283|T201|LC|50410-0|LNC|Autoimmune antibody|Autoimmune antibody
C1978283|T201|MTH_LN|50410-0|LNC|Autoimmune antibody|Autoimmune antibody
C1978287|T201|LN|50413-4|LNC|ACTH|ACTH
C1978287|T201|MTH_LN|50413-4|LNC|ACTH|ACTH
C1978287|T201|OSN|50413-4|LNC|ACTH|ACTH
C1978287|T201|LC|50413-4|LNC|ACTH|ACTH
C1978287|T201|LN|50413-4|LNC|corticotropin|corticotropin
C1978287|T201|MTH_LN|50413-4|LNC|corticotropin|corticotropin
C1978287|T201|OSN|50413-4|LNC|corticotropin|corticotropin
C1978287|T201|LC|50413-4|LNC|corticotropin|corticotropin
C1978287|T201|LN|50413-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978287|T201|MTH_LN|50413-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978287|T201|OSN|50413-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978287|T201|LC|50413-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978288|T201|LN|50414-2|LNC|ACTH|ACTH
C1978288|T201|OSN|50414-2|LNC|ACTH|ACTH
C1978288|T201|MTH_LN|50414-2|LNC|ACTH|ACTH
C1978288|T201|LC|50414-2|LNC|ACTH|ACTH
C1978288|T201|LN|50414-2|LNC|corticotropin|corticotropin
C1978288|T201|OSN|50414-2|LNC|corticotropin|corticotropin
C1978288|T201|MTH_LN|50414-2|LNC|corticotropin|corticotropin
C1978288|T201|LC|50414-2|LNC|corticotropin|corticotropin
C1978288|T201|LN|50414-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978288|T201|OSN|50414-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978288|T201|MTH_LN|50414-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978288|T201|LC|50414-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978291|T201|LN|50417-5|LNC|ACTH|ACTH
C1978291|T201|MTH_LN|50417-5|LNC|ACTH|ACTH
C1978291|T201|OSN|50417-5|LNC|ACTH|ACTH
C1978291|T201|LC|50417-5|LNC|ACTH|ACTH
C1978291|T201|LN|50417-5|LNC|corticotropin|corticotropin
C1978291|T201|MTH_LN|50417-5|LNC|corticotropin|corticotropin
C1978291|T201|OSN|50417-5|LNC|corticotropin|corticotropin
C1978291|T201|LC|50417-5|LNC|corticotropin|corticotropin
C1978291|T201|LN|50417-5|LNC|adrenocorticotropin|adrenocorticotropin
C1978291|T201|MTH_LN|50417-5|LNC|adrenocorticotropin|adrenocorticotropin
C1978291|T201|OSN|50417-5|LNC|adrenocorticotropin|adrenocorticotropin
C1978291|T201|LC|50417-5|LNC|adrenocorticotropin|adrenocorticotropin
C1978292|T201|LN|50418-3|LNC|ACTH|ACTH
C1978292|T201|MTH_LN|50418-3|LNC|ACTH|ACTH
C1978292|T201|OSN|50418-3|LNC|ACTH|ACTH
C1978292|T201|LC|50418-3|LNC|ACTH|ACTH
C1978292|T201|LN|50418-3|LNC|corticotropin|corticotropin
C1978292|T201|MTH_LN|50418-3|LNC|corticotropin|corticotropin
C1978292|T201|OSN|50418-3|LNC|corticotropin|corticotropin
C1978292|T201|LC|50418-3|LNC|corticotropin|corticotropin
C1978292|T201|LN|50418-3|LNC|adrenocorticotropin|adrenocorticotropin
C1978292|T201|MTH_LN|50418-3|LNC|adrenocorticotropin|adrenocorticotropin
C1978292|T201|OSN|50418-3|LNC|adrenocorticotropin|adrenocorticotropin
C1978292|T201|LC|50418-3|LNC|adrenocorticotropin|adrenocorticotropin
C1978293|T201|LN|50419-1|LNC|ACTH|ACTH
C1978293|T201|MTH_LN|50419-1|LNC|ACTH|ACTH
C1978293|T201|OSN|50419-1|LNC|ACTH|ACTH
C1978293|T201|LC|50419-1|LNC|ACTH|ACTH
C1978293|T201|LN|50419-1|LNC|corticotropin|corticotropin
C1978293|T201|MTH_LN|50419-1|LNC|corticotropin|corticotropin
C1978293|T201|OSN|50419-1|LNC|corticotropin|corticotropin
C1978293|T201|LC|50419-1|LNC|corticotropin|corticotropin
C1978293|T201|LN|50419-1|LNC|adrenocorticotropin|adrenocorticotropin
C1978293|T201|MTH_LN|50419-1|LNC|adrenocorticotropin|adrenocorticotropin
C1978293|T201|OSN|50419-1|LNC|adrenocorticotropin|adrenocorticotropin
C1978293|T201|LC|50419-1|LNC|adrenocorticotropin|adrenocorticotropin
C1978294|T201|LN|50420-9|LNC|ACTH|ACTH
C1978294|T201|MTH_LN|50420-9|LNC|ACTH|ACTH
C1978294|T201|OSN|50420-9|LNC|ACTH|ACTH
C1978294|T201|LC|50420-9|LNC|ACTH|ACTH
C1978294|T201|LN|50420-9|LNC|corticotropin|corticotropin
C1978294|T201|MTH_LN|50420-9|LNC|corticotropin|corticotropin
C1978294|T201|OSN|50420-9|LNC|corticotropin|corticotropin
C1978294|T201|LC|50420-9|LNC|corticotropin|corticotropin
C1978294|T201|LN|50420-9|LNC|adrenocorticotropin|adrenocorticotropin
C1978294|T201|MTH_LN|50420-9|LNC|adrenocorticotropin|adrenocorticotropin
C1978294|T201|OSN|50420-9|LNC|adrenocorticotropin|adrenocorticotropin
C1978294|T201|LC|50420-9|LNC|adrenocorticotropin|adrenocorticotropin
C1978299|T201|LN|50425-8|LNC|ACTH|ACTH
C1978299|T201|MTH_LN|50425-8|LNC|ACTH|ACTH
C1978299|T201|OSN|50425-8|LNC|ACTH|ACTH
C1978299|T201|LC|50425-8|LNC|ACTH|ACTH
C1978299|T201|LN|50425-8|LNC|corticotropin|corticotropin
C1978299|T201|MTH_LN|50425-8|LNC|corticotropin|corticotropin
C1978299|T201|OSN|50425-8|LNC|corticotropin|corticotropin
C1978299|T201|LC|50425-8|LNC|corticotropin|corticotropin
C1978299|T201|LN|50425-8|LNC|adrenocorticotropin|adrenocorticotropin
C1978299|T201|MTH_LN|50425-8|LNC|adrenocorticotropin|adrenocorticotropin
C1978299|T201|OSN|50425-8|LNC|adrenocorticotropin|adrenocorticotropin
C1978299|T201|LC|50425-8|LNC|adrenocorticotropin|adrenocorticotropin
C1978300|T201|LN|50426-6|LNC|ACTH|ACTH
C1978300|T201|OSN|50426-6|LNC|ACTH|ACTH
C1978300|T201|MTH_LN|50426-6|LNC|ACTH|ACTH
C1978300|T201|LC|50426-6|LNC|ACTH|ACTH
C1978300|T201|LN|50426-6|LNC|corticotropin|corticotropin
C1978300|T201|OSN|50426-6|LNC|corticotropin|corticotropin
C1978300|T201|MTH_LN|50426-6|LNC|corticotropin|corticotropin
C1978300|T201|LC|50426-6|LNC|corticotropin|corticotropin
C1978300|T201|LN|50426-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978300|T201|OSN|50426-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978300|T201|MTH_LN|50426-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978300|T201|LC|50426-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978301|T201|LN|50427-4|LNC|ACTH|ACTH
C1978301|T201|MTH_LN|50427-4|LNC|ACTH|ACTH
C1978301|T201|OSN|50427-4|LNC|ACTH|ACTH
C1978301|T201|LC|50427-4|LNC|ACTH|ACTH
C1978301|T201|LN|50427-4|LNC|corticotropin|corticotropin
C1978301|T201|MTH_LN|50427-4|LNC|corticotropin|corticotropin
C1978301|T201|OSN|50427-4|LNC|corticotropin|corticotropin
C1978301|T201|LC|50427-4|LNC|corticotropin|corticotropin
C1978301|T201|LN|50427-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978301|T201|MTH_LN|50427-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978301|T201|OSN|50427-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978301|T201|LC|50427-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978302|T201|LN|50428-2|LNC|ACTH|ACTH
C1978302|T201|MTH_LN|50428-2|LNC|ACTH|ACTH
C1978302|T201|OSN|50428-2|LNC|ACTH|ACTH
C1978302|T201|LC|50428-2|LNC|ACTH|ACTH
C1978302|T201|LN|50428-2|LNC|corticotropin|corticotropin
C1978302|T201|MTH_LN|50428-2|LNC|corticotropin|corticotropin
C1978302|T201|OSN|50428-2|LNC|corticotropin|corticotropin
C1978302|T201|LC|50428-2|LNC|corticotropin|corticotropin
C1978302|T201|LN|50428-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978302|T201|MTH_LN|50428-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978302|T201|OSN|50428-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978302|T201|LC|50428-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978309|T201|LN|50435-7|LNC|ACTH|ACTH
C1978309|T201|MTH_LN|50435-7|LNC|ACTH|ACTH
C1978309|T201|OSN|50435-7|LNC|ACTH|ACTH
C1978309|T201|LC|50435-7|LNC|ACTH|ACTH
C1978309|T201|LN|50435-7|LNC|corticotropin|corticotropin
C1978309|T201|MTH_LN|50435-7|LNC|corticotropin|corticotropin
C1978309|T201|OSN|50435-7|LNC|corticotropin|corticotropin
C1978309|T201|LC|50435-7|LNC|corticotropin|corticotropin
C1978309|T201|LN|50435-7|LNC|adrenocorticotropin|adrenocorticotropin
C1978309|T201|MTH_LN|50435-7|LNC|adrenocorticotropin|adrenocorticotropin
C1978309|T201|OSN|50435-7|LNC|adrenocorticotropin|adrenocorticotropin
C1978309|T201|LC|50435-7|LNC|adrenocorticotropin|adrenocorticotropin
C1978310|T201|LN|50436-5|LNC|ACTH|ACTH
C1978310|T201|MTH_LN|50436-5|LNC|ACTH|ACTH
C1978310|T201|OSN|50436-5|LNC|ACTH|ACTH
C1978310|T201|LC|50436-5|LNC|ACTH|ACTH
C1978310|T201|LN|50436-5|LNC|corticotropin|corticotropin
C1978310|T201|MTH_LN|50436-5|LNC|corticotropin|corticotropin
C1978310|T201|OSN|50436-5|LNC|corticotropin|corticotropin
C1978310|T201|LC|50436-5|LNC|corticotropin|corticotropin
C1978310|T201|LN|50436-5|LNC|adrenocorticotropin|adrenocorticotropin
C1978310|T201|MTH_LN|50436-5|LNC|adrenocorticotropin|adrenocorticotropin
C1978310|T201|OSN|50436-5|LNC|adrenocorticotropin|adrenocorticotropin
C1978310|T201|LC|50436-5|LNC|adrenocorticotropin|adrenocorticotropin
C1978311|T201|LN|50437-3|LNC|ACTH|ACTH
C1978311|T201|OSN|50437-3|LNC|ACTH|ACTH
C1978311|T201|MTH_LN|50437-3|LNC|ACTH|ACTH
C1978311|T201|LC|50437-3|LNC|ACTH|ACTH
C1978311|T201|LN|50437-3|LNC|corticotropin|corticotropin
C1978311|T201|OSN|50437-3|LNC|corticotropin|corticotropin
C1978311|T201|MTH_LN|50437-3|LNC|corticotropin|corticotropin
C1978311|T201|LC|50437-3|LNC|corticotropin|corticotropin
C1978311|T201|LN|50437-3|LNC|adrenocorticotropin|adrenocorticotropin
C1978311|T201|OSN|50437-3|LNC|adrenocorticotropin|adrenocorticotropin
C1978311|T201|MTH_LN|50437-3|LNC|adrenocorticotropin|adrenocorticotropin
C1978311|T201|LC|50437-3|LNC|adrenocorticotropin|adrenocorticotropin
C1978312|T201|LN|50438-1|LNC|ACTH|ACTH
C1978312|T201|MTH_LN|50438-1|LNC|ACTH|ACTH
C1978312|T201|OSN|50438-1|LNC|ACTH|ACTH
C1978312|T201|LC|50438-1|LNC|ACTH|ACTH
C1978312|T201|LN|50438-1|LNC|corticotropin|corticotropin
C1978312|T201|MTH_LN|50438-1|LNC|corticotropin|corticotropin
C1978312|T201|OSN|50438-1|LNC|corticotropin|corticotropin
C1978312|T201|LC|50438-1|LNC|corticotropin|corticotropin
C1978312|T201|LN|50438-1|LNC|adrenocorticotropin|adrenocorticotropin
C1978312|T201|MTH_LN|50438-1|LNC|adrenocorticotropin|adrenocorticotropin
C1978312|T201|OSN|50438-1|LNC|adrenocorticotropin|adrenocorticotropin
C1978312|T201|LC|50438-1|LNC|adrenocorticotropin|adrenocorticotropin
C1978313|T201|LN|50439-9|LNC|ACTH|ACTH
C1978313|T201|MTH_LN|50439-9|LNC|ACTH|ACTH
C1978313|T201|OSN|50439-9|LNC|ACTH|ACTH
C1978313|T201|LC|50439-9|LNC|ACTH|ACTH
C1978313|T201|LN|50439-9|LNC|corticotropin|corticotropin
C1978313|T201|MTH_LN|50439-9|LNC|corticotropin|corticotropin
C1978313|T201|OSN|50439-9|LNC|corticotropin|corticotropin
C1978313|T201|LC|50439-9|LNC|corticotropin|corticotropin
C1978313|T201|LN|50439-9|LNC|adrenocorticotropin|adrenocorticotropin
C1978313|T201|MTH_LN|50439-9|LNC|adrenocorticotropin|adrenocorticotropin
C1978313|T201|OSN|50439-9|LNC|adrenocorticotropin|adrenocorticotropin
C1978313|T201|LC|50439-9|LNC|adrenocorticotropin|adrenocorticotropin
C1978314|T201|LN|50440-7|LNC|ACTH|ACTH
C1978314|T201|MTH_LN|50440-7|LNC|ACTH|ACTH
C1978314|T201|OSN|50440-7|LNC|ACTH|ACTH
C1978314|T201|LC|50440-7|LNC|ACTH|ACTH
C1978314|T201|LN|50440-7|LNC|corticotropin|corticotropin
C1978314|T201|MTH_LN|50440-7|LNC|corticotropin|corticotropin
C1978314|T201|OSN|50440-7|LNC|corticotropin|corticotropin
C1978314|T201|LC|50440-7|LNC|corticotropin|corticotropin
C1978314|T201|LN|50440-7|LNC|adrenocorticotropin|adrenocorticotropin
C1978314|T201|MTH_LN|50440-7|LNC|adrenocorticotropin|adrenocorticotropin
C1978314|T201|OSN|50440-7|LNC|adrenocorticotropin|adrenocorticotropin
C1978314|T201|LC|50440-7|LNC|adrenocorticotropin|adrenocorticotropin
C1978319|T201|LN|50445-6|LNC|ACTH|ACTH
C1978319|T201|MTH_LN|50445-6|LNC|ACTH|ACTH
C1978319|T201|OSN|50445-6|LNC|ACTH|ACTH
C1978319|T201|LC|50445-6|LNC|ACTH|ACTH
C1978319|T201|LN|50445-6|LNC|corticotropin|corticotropin
C1978319|T201|MTH_LN|50445-6|LNC|corticotropin|corticotropin
C1978319|T201|OSN|50445-6|LNC|corticotropin|corticotropin
C1978319|T201|LC|50445-6|LNC|corticotropin|corticotropin
C1978319|T201|LN|50445-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978319|T201|MTH_LN|50445-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978319|T201|OSN|50445-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978319|T201|LC|50445-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978320|T201|LN|50446-4|LNC|ACTH|ACTH
C1978320|T201|MTH_LN|50446-4|LNC|ACTH|ACTH
C1978320|T201|OSN|50446-4|LNC|ACTH|ACTH
C1978320|T201|LC|50446-4|LNC|ACTH|ACTH
C1978320|T201|LN|50446-4|LNC|corticotropin|corticotropin
C1978320|T201|MTH_LN|50446-4|LNC|corticotropin|corticotropin
C1978320|T201|OSN|50446-4|LNC|corticotropin|corticotropin
C1978320|T201|LC|50446-4|LNC|corticotropin|corticotropin
C1978320|T201|LN|50446-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978320|T201|MTH_LN|50446-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978320|T201|OSN|50446-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978320|T201|LC|50446-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978321|T201|LN|50447-2|LNC|ACTH|ACTH
C1978321|T201|MTH_LN|50447-2|LNC|ACTH|ACTH
C1978321|T201|OSN|50447-2|LNC|ACTH|ACTH
C1978321|T201|LC|50447-2|LNC|ACTH|ACTH
C1978321|T201|LN|50447-2|LNC|corticotropin|corticotropin
C1978321|T201|MTH_LN|50447-2|LNC|corticotropin|corticotropin
C1978321|T201|OSN|50447-2|LNC|corticotropin|corticotropin
C1978321|T201|LC|50447-2|LNC|corticotropin|corticotropin
C1978321|T201|LN|50447-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978321|T201|MTH_LN|50447-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978321|T201|OSN|50447-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978321|T201|LC|50447-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978322|T201|LN|50448-0|LNC|ACTH|ACTH
C1978322|T201|MTH_LN|50448-0|LNC|ACTH|ACTH
C1978322|T201|OSN|50448-0|LNC|ACTH|ACTH
C1978322|T201|LC|50448-0|LNC|ACTH|ACTH
C1978322|T201|LN|50448-0|LNC|corticotropin|corticotropin
C1978322|T201|MTH_LN|50448-0|LNC|corticotropin|corticotropin
C1978322|T201|OSN|50448-0|LNC|corticotropin|corticotropin
C1978322|T201|LC|50448-0|LNC|corticotropin|corticotropin
C1978322|T201|LN|50448-0|LNC|adrenocorticotropin|adrenocorticotropin
C1978322|T201|MTH_LN|50448-0|LNC|adrenocorticotropin|adrenocorticotropin
C1978322|T201|OSN|50448-0|LNC|adrenocorticotropin|adrenocorticotropin
C1978322|T201|LC|50448-0|LNC|adrenocorticotropin|adrenocorticotropin
C1978323|T201|LN|50449-8|LNC|ACTH|ACTH
C1978323|T201|OSN|50449-8|LNC|ACTH|ACTH
C1978323|T201|MTH_LN|50449-8|LNC|ACTH|ACTH
C1978323|T201|LC|50449-8|LNC|ACTH|ACTH
C1978323|T201|LN|50449-8|LNC|corticotropin|corticotropin
C1978323|T201|OSN|50449-8|LNC|corticotropin|corticotropin
C1978323|T201|MTH_LN|50449-8|LNC|corticotropin|corticotropin
C1978323|T201|LC|50449-8|LNC|corticotropin|corticotropin
C1978323|T201|LN|50449-8|LNC|adrenocorticotropin|adrenocorticotropin
C1978323|T201|OSN|50449-8|LNC|adrenocorticotropin|adrenocorticotropin
C1978323|T201|MTH_LN|50449-8|LNC|adrenocorticotropin|adrenocorticotropin
C1978323|T201|LC|50449-8|LNC|adrenocorticotropin|adrenocorticotropin
C1978324|T201|LN|50450-6|LNC|ACTH|ACTH
C1978324|T201|MTH_LN|50450-6|LNC|ACTH|ACTH
C1978324|T201|OSN|50450-6|LNC|ACTH|ACTH
C1978324|T201|LC|50450-6|LNC|ACTH|ACTH
C1978324|T201|LN|50450-6|LNC|corticotropin|corticotropin
C1978324|T201|MTH_LN|50450-6|LNC|corticotropin|corticotropin
C1978324|T201|OSN|50450-6|LNC|corticotropin|corticotropin
C1978324|T201|LC|50450-6|LNC|corticotropin|corticotropin
C1978324|T201|LN|50450-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978324|T201|MTH_LN|50450-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978324|T201|OSN|50450-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978324|T201|LC|50450-6|LNC|adrenocorticotropin|adrenocorticotropin
C1978325|T201|LN|50451-4|LNC|ACTH|ACTH
C1978325|T201|MTH_LN|50451-4|LNC|ACTH|ACTH
C1978325|T201|OSN|50451-4|LNC|ACTH|ACTH
C1978325|T201|LC|50451-4|LNC|ACTH|ACTH
C1978325|T201|LN|50451-4|LNC|corticotropin|corticotropin
C1978325|T201|MTH_LN|50451-4|LNC|corticotropin|corticotropin
C1978325|T201|OSN|50451-4|LNC|corticotropin|corticotropin
C1978325|T201|LC|50451-4|LNC|corticotropin|corticotropin
C1978325|T201|LN|50451-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978325|T201|MTH_LN|50451-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978325|T201|OSN|50451-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978325|T201|LC|50451-4|LNC|adrenocorticotropin|adrenocorticotropin
C1978326|T201|LN|50452-2|LNC|ACTH|ACTH
C1978326|T201|OSN|50452-2|LNC|ACTH|ACTH
C1978326|T201|MTH_LN|50452-2|LNC|ACTH|ACTH
C1978326|T201|LC|50452-2|LNC|ACTH|ACTH
C1978326|T201|LN|50452-2|LNC|corticotropin|corticotropin
C1978326|T201|OSN|50452-2|LNC|corticotropin|corticotropin
C1978326|T201|MTH_LN|50452-2|LNC|corticotropin|corticotropin
C1978326|T201|LC|50452-2|LNC|corticotropin|corticotropin
C1978326|T201|LN|50452-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978326|T201|OSN|50452-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978326|T201|MTH_LN|50452-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978326|T201|LC|50452-2|LNC|adrenocorticotropin|adrenocorticotropin
C1978335|T201|LN|50461-3|LNC|C-peptide|C-peptide
C1978335|T201|MTH_LN|50461-3|LNC|C-peptide|C-peptide
C1978335|T201|OSN|50461-3|LNC|C-peptide|C-peptide
C1978335|T201|LC|50461-3|LNC|C-peptide|C-peptide
C1978335|T201|LN|50461-3|LNC|C peptide|C peptide
C1978335|T201|MTH_LN|50461-3|LNC|C peptide|C peptide
C1978335|T201|OSN|50461-3|LNC|C peptide|C peptide
C1978335|T201|LC|50461-3|LNC|C peptide|C peptide
C1978336|T201|LN|50462-1|LNC|C-peptide|C-peptide
C1978336|T201|MTH_LN|50462-1|LNC|C-peptide|C-peptide
C1978336|T201|OSN|50462-1|LNC|C-peptide|C-peptide
C1978336|T201|LC|50462-1|LNC|C-peptide|C-peptide
C1978336|T201|LN|50462-1|LNC|C peptide|C peptide
C1978336|T201|MTH_LN|50462-1|LNC|C peptide|C peptide
C1978336|T201|OSN|50462-1|LNC|C peptide|C peptide
C1978336|T201|LC|50462-1|LNC|C peptide|C peptide
C1978337|T201|LN|50463-9|LNC|C-peptide|C-peptide
C1978337|T201|OSN|50463-9|LNC|C-peptide|C-peptide
C1978337|T201|MTH_LN|50463-9|LNC|C-peptide|C-peptide
C1978337|T201|LC|50463-9|LNC|C-peptide|C-peptide
C1978337|T201|LN|50463-9|LNC|C peptide|C peptide
C1978337|T201|OSN|50463-9|LNC|C peptide|C peptide
C1978337|T201|MTH_LN|50463-9|LNC|C peptide|C peptide
C1978337|T201|LC|50463-9|LNC|C peptide|C peptide
C1978338|T201|LN|50464-7|LNC|C-peptide|C-peptide
C1978338|T201|OSN|50464-7|LNC|C-peptide|C-peptide
C1978338|T201|MTH_LN|50464-7|LNC|C-peptide|C-peptide
C1978338|T201|LC|50464-7|LNC|C-peptide|C-peptide
C1978338|T201|LN|50464-7|LNC|C peptide|C peptide
C1978338|T201|OSN|50464-7|LNC|C peptide|C peptide
C1978338|T201|MTH_LN|50464-7|LNC|C peptide|C peptide
C1978338|T201|LC|50464-7|LNC|C peptide|C peptide
C1978339|T201|LN|50465-4|LNC|C-peptide|C-peptide
C1978339|T201|OSN|50465-4|LNC|C-peptide|C-peptide
C1978339|T201|MTH_LN|50465-4|LNC|C-peptide|C-peptide
C1978339|T201|LC|50465-4|LNC|C-peptide|C-peptide
C1978339|T201|LN|50465-4|LNC|C peptide|C peptide
C1978339|T201|OSN|50465-4|LNC|C peptide|C peptide
C1978339|T201|MTH_LN|50465-4|LNC|C peptide|C peptide
C1978339|T201|LC|50465-4|LNC|C peptide|C peptide
C1978340|T201|LN|50466-2|LNC|C-peptide|C-peptide
C1978340|T201|MTH_LN|50466-2|LNC|C-peptide|C-peptide
C1978340|T201|OSN|50466-2|LNC|C-peptide|C-peptide
C1978340|T201|LC|50466-2|LNC|C-peptide|C-peptide
C1978340|T201|LN|50466-2|LNC|C peptide|C peptide
C1978340|T201|MTH_LN|50466-2|LNC|C peptide|C peptide
C1978340|T201|OSN|50466-2|LNC|C peptide|C peptide
C1978340|T201|LC|50466-2|LNC|C peptide|C peptide
C1978341|T201|LN|50467-0|LNC|C-peptide|C-peptide
C1978341|T201|MTH_LN|50467-0|LNC|C-peptide|C-peptide
C1978341|T201|OSN|50467-0|LNC|C-peptide|C-peptide
C1978341|T201|LC|50467-0|LNC|C-peptide|C-peptide
C1978341|T201|LN|50467-0|LNC|C peptide|C peptide
C1978341|T201|MTH_LN|50467-0|LNC|C peptide|C peptide
C1978341|T201|OSN|50467-0|LNC|C peptide|C peptide
C1978341|T201|LC|50467-0|LNC|C peptide|C peptide
C1978342|T201|LN|50468-8|LNC|C-peptide|C-peptide
C1978342|T201|OSN|50468-8|LNC|C-peptide|C-peptide
C1978342|T201|MTH_LN|50468-8|LNC|C-peptide|C-peptide
C1978342|T201|LC|50468-8|LNC|C-peptide|C-peptide
C1978342|T201|LN|50468-8|LNC|C peptide|C peptide
C1978342|T201|OSN|50468-8|LNC|C peptide|C peptide
C1978342|T201|MTH_LN|50468-8|LNC|C peptide|C peptide
C1978342|T201|LC|50468-8|LNC|C peptide|C peptide
C1978383|T201|LN|50509-9|LNC|luteinizing|luteinizing
C1978383|T201|MTH_LN|50509-9|LNC|luteinizing|luteinizing
C1978383|T201|OSN|50509-9|LNC|luteinizing|luteinizing
C1978383|T201|LC|50509-9|LNC|luteinizing|luteinizing
C1978383|T201|LN|50509-9|LNC|LH|LH
C1978383|T201|MTH_LN|50509-9|LNC|LH|LH
C1978383|T201|OSN|50509-9|LNC|LH|LH
C1978383|T201|LC|50509-9|LNC|LH|LH
C1978383|T201|LN|50509-9|LNC|luteinising|luteinising
C1978383|T201|MTH_LN|50509-9|LNC|luteinising|luteinising
C1978383|T201|OSN|50509-9|LNC|luteinising|luteinising
C1978383|T201|LC|50509-9|LNC|luteinising|luteinising
C1978384|T201|LN|50510-7|LNC|luteinizing|luteinizing
C1978384|T201|OSN|50510-7|LNC|luteinizing|luteinizing
C1978384|T201|MTH_LN|50510-7|LNC|luteinizing|luteinizing
C1978384|T201|LC|50510-7|LNC|luteinizing|luteinizing
C1978384|T201|LN|50510-7|LNC|LH|LH
C1978384|T201|OSN|50510-7|LNC|LH|LH
C1978384|T201|MTH_LN|50510-7|LNC|LH|LH
C1978384|T201|LC|50510-7|LNC|LH|LH
C1978384|T201|LN|50510-7|LNC|luteinising|luteinising
C1978384|T201|OSN|50510-7|LNC|luteinising|luteinising
C1978384|T201|MTH_LN|50510-7|LNC|luteinising|luteinising
C1978384|T201|LC|50510-7|LNC|luteinising|luteinising
C1978385|T201|LN|50511-5|LNC|luteinizing|luteinizing
C1978385|T201|OSN|50511-5|LNC|luteinizing|luteinizing
C1978385|T201|MTH_LN|50511-5|LNC|luteinizing|luteinizing
C1978385|T201|LC|50511-5|LNC|luteinizing|luteinizing
C1978385|T201|LN|50511-5|LNC|LH|LH
C1978385|T201|OSN|50511-5|LNC|LH|LH
C1978385|T201|MTH_LN|50511-5|LNC|LH|LH
C1978385|T201|LC|50511-5|LNC|LH|LH
C1978385|T201|LN|50511-5|LNC|luteinising|luteinising
C1978385|T201|OSN|50511-5|LNC|luteinising|luteinising
C1978385|T201|MTH_LN|50511-5|LNC|luteinising|luteinising
C1978385|T201|LC|50511-5|LNC|luteinising|luteinising
C1978386|T201|LN|50512-3|LNC|luteinizing|luteinizing
C1978386|T201|OSN|50512-3|LNC|luteinizing|luteinizing
C1978386|T201|MTH_LN|50512-3|LNC|luteinizing|luteinizing
C1978386|T201|LC|50512-3|LNC|luteinizing|luteinizing
C1978386|T201|LN|50512-3|LNC|LH|LH
C1978386|T201|OSN|50512-3|LNC|LH|LH
C1978386|T201|MTH_LN|50512-3|LNC|LH|LH
C1978386|T201|LC|50512-3|LNC|LH|LH
C1978386|T201|LN|50512-3|LNC|luteinising|luteinising
C1978386|T201|OSN|50512-3|LNC|luteinising|luteinising
C1978386|T201|MTH_LN|50512-3|LNC|luteinising|luteinising
C1978386|T201|LC|50512-3|LNC|luteinising|luteinising
C1978387|T201|LN|50513-1|LNC|luteinizing|luteinizing
C1978387|T201|MTH_LN|50513-1|LNC|luteinizing|luteinizing
C1978387|T201|OSN|50513-1|LNC|luteinizing|luteinizing
C1978387|T201|LC|50513-1|LNC|luteinizing|luteinizing
C1978387|T201|LN|50513-1|LNC|LH|LH
C1978387|T201|MTH_LN|50513-1|LNC|LH|LH
C1978387|T201|OSN|50513-1|LNC|LH|LH
C1978387|T201|LC|50513-1|LNC|LH|LH
C1978387|T201|LN|50513-1|LNC|luteinising|luteinising
C1978387|T201|MTH_LN|50513-1|LNC|luteinising|luteinising
C1978387|T201|OSN|50513-1|LNC|luteinising|luteinising
C1978387|T201|LC|50513-1|LNC|luteinising|luteinising
C1978388|T201|LN|50514-9|LNC|luteinizing|luteinizing
C1978388|T201|OSN|50514-9|LNC|luteinizing|luteinizing
C1978388|T201|MTH_LN|50514-9|LNC|luteinizing|luteinizing
C1978388|T201|LC|50514-9|LNC|luteinizing|luteinizing
C1978388|T201|LN|50514-9|LNC|LH|LH
C1978388|T201|OSN|50514-9|LNC|LH|LH
C1978388|T201|MTH_LN|50514-9|LNC|LH|LH
C1978388|T201|LC|50514-9|LNC|LH|LH
C1978388|T201|LN|50514-9|LNC|luteinising|luteinising
C1978388|T201|OSN|50514-9|LNC|luteinising|luteinising
C1978388|T201|MTH_LN|50514-9|LNC|luteinising|luteinising
C1978388|T201|LC|50514-9|LNC|luteinising|luteinising
C1978389|T201|LN|50515-6|LNC|luteinizing|luteinizing
C1978389|T201|OSN|50515-6|LNC|luteinizing|luteinizing
C1978389|T201|MTH_LN|50515-6|LNC|luteinizing|luteinizing
C1978389|T201|LC|50515-6|LNC|luteinizing|luteinizing
C1978389|T201|LN|50515-6|LNC|LH|LH
C1978389|T201|OSN|50515-6|LNC|LH|LH
C1978389|T201|MTH_LN|50515-6|LNC|LH|LH
C1978389|T201|LC|50515-6|LNC|LH|LH
C1978389|T201|LN|50515-6|LNC|luteinising|luteinising
C1978389|T201|OSN|50515-6|LNC|luteinising|luteinising
C1978389|T201|MTH_LN|50515-6|LNC|luteinising|luteinising
C1978389|T201|LC|50515-6|LNC|luteinising|luteinising
C1978390|T201|LN|50516-4|LNC|luteinizing|luteinizing
C1978390|T201|OSN|50516-4|LNC|luteinizing|luteinizing
C1978390|T201|MTH_LN|50516-4|LNC|luteinizing|luteinizing
C1978390|T201|LC|50516-4|LNC|luteinizing|luteinizing
C1978390|T201|LN|50516-4|LNC|LH|LH
C1978390|T201|OSN|50516-4|LNC|LH|LH
C1978390|T201|MTH_LN|50516-4|LNC|LH|LH
C1978390|T201|LC|50516-4|LNC|LH|LH
C1978390|T201|LN|50516-4|LNC|luteinising|luteinising
C1978390|T201|OSN|50516-4|LNC|luteinising|luteinising
C1978390|T201|MTH_LN|50516-4|LNC|luteinising|luteinising
C1978390|T201|LC|50516-4|LNC|luteinising|luteinising
C1978480|T201|LN|50553-7|LNC|Red|Red
C1978480|T201|OSN|50553-7|LNC|Red|Red
C1978480|T201|MTH_LN|50553-7|LNC|Red|Red
C1978480|T201|LC|50553-7|LNC|Red|Red
C1978480|T201|LN|50553-7|LNC|Red-brown|Red-brown
C1978480|T201|OSN|50553-7|LNC|Red-brown|Red-brown
C1978480|T201|MTH_LN|50553-7|LNC|Red-brown|Red-brown
C1978480|T201|LC|50553-7|LNC|Red-brown|Red-brown
C1978480|T201|LN|50553-7|LNC|red brown|red brown
C1978480|T201|OSN|50553-7|LNC|red brown|red brown
C1978480|T201|MTH_LN|50553-7|LNC|red brown|red brown
C1978480|T201|LC|50553-7|LNC|red brown|red brown
C1978480|T201|LN|50553-7|LNC|Purple|Purple
C1978480|T201|OSN|50553-7|LNC|Purple|Purple
C1978480|T201|MTH_LN|50553-7|LNC|Purple|Purple
C1978480|T201|LC|50553-7|LNC|Purple|Purple
C1978480|T201|LN|50553-7|LNC|Blue|Blue
C1978480|T201|OSN|50553-7|LNC|Blue|Blue
C1978480|T201|MTH_LN|50553-7|LNC|Blue|Blue
C1978480|T201|LC|50553-7|LNC|Blue|Blue
C1978486|T201|LN|50559-4|LNC|Hemoglobin|Hemoglobin
C1978486|T201|OSN|50559-4|LNC|Hemoglobin|Hemoglobin
C1978486|T201|MTH_LN|50559-4|LNC|Hemoglobin|Hemoglobin
C1978486|T201|LC|50559-4|LNC|Hemoglobin|Hemoglobin
C1978489|T201|LN|50562-8|LNC|osmolality|osmolality
C1978489|T201|MTH_LN|50562-8|LNC|osmolality|osmolality
C1978489|T201|OSN|50562-8|LNC|osmolality|osmolality
C1978489|T201|LC|50562-8|LNC|osmolality|osmolality
C1978489|T201|LN|50562-8|LNC|homeostasis|homeostasis
C1978489|T201|MTH_LN|50562-8|LNC|homeostasis|homeostasis
C1978489|T201|OSN|50562-8|LNC|homeostasis|homeostasis
C1978489|T201|LC|50562-8|LNC|homeostasis|homeostasis
C1978490|T201|LN|50563-6|LNC|urobilinogen|urobilinogen
C1978490|T201|OSN|50563-6|LNC|urobilinogen|urobilinogen
C1978490|T201|MTH_LN|50563-6|LNC|urobilinogen|urobilinogen
C1978490|T201|LC|50563-6|LNC|urobilinogen|urobilinogen
C1978568|T201|LN|50609-7|LNC|nitroblue tetrazolium reduction test|nitroblue tetrazolium reduction test
C1978568|T201|OSN|50609-7|LNC|nitroblue tetrazolium reduction test|nitroblue tetrazolium reduction test
C1978568|T201|MTH_LN|50609-7|LNC|nitroblue tetrazolium reduction test|nitroblue tetrazolium reduction test
C1978568|T201|LC|50609-7|LNC|nitroblue tetrazolium reduction test|nitroblue tetrazolium reduction test
C1978568|T201|LN|50609-7|LNC|NBT reduction test|NBT reduction test
C1978568|T201|OSN|50609-7|LNC|NBT reduction test|NBT reduction test
C1978568|T201|MTH_LN|50609-7|LNC|NBT reduction test|NBT reduction test
C1978568|T201|LC|50609-7|LNC|NBT reduction test|NBT reduction test
C1978782|T201|LN|50770-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1978782|T201|OSN|50770-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1978782|T201|MTH_LN|50770-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1978782|T201|LC|50770-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C1979375|T201|LN|51329-1|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979375|T201|MTH_LN|51329-1|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979375|T201|LC|51329-1|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979375|T201|OSN|51329-1|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979375|T201|LN|51329-1|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979375|T201|MTH_LN|51329-1|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979375|T201|LC|51329-1|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979375|T201|OSN|51329-1|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979375|T201|LN|51329-1|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979375|T201|MTH_LN|51329-1|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979375|T201|LC|51329-1|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979375|T201|OSN|51329-1|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979375|T201|LN|51329-1|LNC|T cell subset distribution|T cell subset distribution
C1979375|T201|MTH_LN|51329-1|LNC|T cell subset distribution|T cell subset distribution
C1979375|T201|LC|51329-1|LNC|T cell subset distribution|T cell subset distribution
C1979375|T201|OSN|51329-1|LNC|T cell subset distribution|T cell subset distribution
C1979376|T201|LN|51330-9|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979376|T201|MTH_LN|51330-9|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979376|T201|LC|51330-9|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979376|T201|OSN|51330-9|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979376|T201|LN|51330-9|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979376|T201|MTH_LN|51330-9|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979376|T201|LC|51330-9|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979376|T201|OSN|51330-9|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979376|T201|LN|51330-9|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979376|T201|MTH_LN|51330-9|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979376|T201|LC|51330-9|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979376|T201|OSN|51330-9|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979376|T201|LN|51330-9|LNC|T cell subset distribution|T cell subset distribution
C1979376|T201|MTH_LN|51330-9|LNC|T cell subset distribution|T cell subset distribution
C1979376|T201|LC|51330-9|LNC|T cell subset distribution|T cell subset distribution
C1979376|T201|OSN|51330-9|LNC|T cell subset distribution|T cell subset distribution
C1979377|T201|LN|51331-7|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979377|T201|MTH_LN|51331-7|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979377|T201|LC|51331-7|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979377|T201|OSN|51331-7|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979377|T201|LN|51331-7|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979377|T201|MTH_LN|51331-7|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979377|T201|LC|51331-7|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979377|T201|OSN|51331-7|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979377|T201|LN|51331-7|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979377|T201|MTH_LN|51331-7|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979377|T201|LC|51331-7|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979377|T201|OSN|51331-7|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979377|T201|LN|51331-7|LNC|T cell subset distribution|T cell subset distribution
C1979377|T201|MTH_LN|51331-7|LNC|T cell subset distribution|T cell subset distribution
C1979377|T201|LC|51331-7|LNC|T cell subset distribution|T cell subset distribution
C1979377|T201|OSN|51331-7|LNC|T cell subset distribution|T cell subset distribution
C1979378|T201|LN|51332-5|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979378|T201|MTH_LN|51332-5|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979378|T201|LC|51332-5|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979378|T201|OSN|51332-5|LNC|lymphocyte surface expressionCD43|lymphocyte surface expressionCD43
C1979378|T201|LN|51332-5|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979378|T201|MTH_LN|51332-5|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979378|T201|LC|51332-5|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979378|T201|OSN|51332-5|LNC|Cd43 defectively expressed on surface of|Cd43 defectively expressed on surface of
C1979378|T201|LN|51332-5|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979378|T201|MTH_LN|51332-5|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979378|T201|LC|51332-5|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979378|T201|OSN|51332-5|LNC|lymphocyte surface expressionsialophorin|lymphocyte surface expressionsialophorin
C1979378|T201|LN|51332-5|LNC|T cell subset distribution|T cell subset distribution
C1979378|T201|MTH_LN|51332-5|LNC|T cell subset distribution|T cell subset distribution
C1979378|T201|LC|51332-5|LNC|T cell subset distribution|T cell subset distribution
C1979378|T201|OSN|51332-5|LNC|T cell subset distribution|T cell subset distribution
C1979446|T201|LN|51423-2|LNC|ACTH|ACTH
C1979446|T201|MTH_LN|51423-2|LNC|ACTH|ACTH
C1979446|T201|OSN|51423-2|LNC|ACTH|ACTH
C1979446|T201|LC|51423-2|LNC|ACTH|ACTH
C1979446|T201|LN|51423-2|LNC|corticotropin|corticotropin
C1979446|T201|MTH_LN|51423-2|LNC|corticotropin|corticotropin
C1979446|T201|OSN|51423-2|LNC|corticotropin|corticotropin
C1979446|T201|LC|51423-2|LNC|corticotropin|corticotropin
C1979446|T201|LN|51423-2|LNC|adrenocorticotropin|adrenocorticotropin
C1979446|T201|MTH_LN|51423-2|LNC|adrenocorticotropin|adrenocorticotropin
C1979446|T201|OSN|51423-2|LNC|adrenocorticotropin|adrenocorticotropin
C1979446|T201|LC|51423-2|LNC|adrenocorticotropin|adrenocorticotropin
C1979451|T201|LN|51428-1|LNC|lactate|lactate
C1979451|T201|LC|51428-1|LNC|lactate|lactate
C1979451|T201|MTH_LN|51428-1|LNC|lactate|lactate
C1979451|T201|OSN|51428-1|LNC|lactate|lactate
C1979494|T201|LN|51478-6|LNC|homeostasis|homeostasis
C1979494|T201|OSN|51478-6|LNC|homeostasis|homeostasis
C1979494|T201|MTH_LN|51478-6|LNC|homeostasis|homeostasis
C1979494|T201|LC|51478-6|LNC|homeostasis|homeostasis
C1979503|T201|LN|51487-7|LNC|neutrophil count|neutrophil count
C1979503|T201|MTH_LN|51487-7|LNC|neutrophil count|neutrophil count
C1979503|T201|OSN|51487-7|LNC|neutrophil count|neutrophil count
C1979503|T201|LC|51487-7|LNC|neutrophil count|neutrophil count
C1979503|T201|LN|51487-7|LNC|cytology|cytology
C1979503|T201|MTH_LN|51487-7|LNC|cytology|cytology
C1979503|T201|OSN|51487-7|LNC|cytology|cytology
C1979503|T201|LC|51487-7|LNC|cytology|cytology
C2360374|T201|LN|51696-3|LNC|ACTH|ACTH
C2360374|T201|LC|51696-3|LNC|ACTH|ACTH
C2360374|T201|MTH_LN|51696-3|LNC|ACTH|ACTH
C2360374|T201|OSN|51696-3|LNC|ACTH|ACTH
C2360374|T201|LN|51696-3|LNC|corticotropin|corticotropin
C2360374|T201|LC|51696-3|LNC|corticotropin|corticotropin
C2360374|T201|MTH_LN|51696-3|LNC|corticotropin|corticotropin
C2360374|T201|OSN|51696-3|LNC|corticotropin|corticotropin
C2360374|T201|LN|51696-3|LNC|adrenocorticotropin|adrenocorticotropin
C2360374|T201|LC|51696-3|LNC|adrenocorticotropin|adrenocorticotropin
C2360374|T201|MTH_LN|51696-3|LNC|adrenocorticotropin|adrenocorticotropin
C2360374|T201|OSN|51696-3|LNC|adrenocorticotropin|adrenocorticotropin
C2360383|T201|LN|51703-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C2360383|T201|OSN|51703-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C2360383|T201|MTH_LN|51703-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C2360383|T201|LC|51703-7|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C2360395|T201|LN|51715-1|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2360395|T201|OSN|51715-1|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2360395|T201|MTH_LN|51715-1|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2360395|T201|LC|51715-1|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2360412|T201|LN|51729-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C2360412|T201|OSN|51729-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C2360412|T201|MTH_LN|51729-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C2360412|T201|LC|51729-2|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C2360416|T201|LN|51733-4|LNC|oxygen|oxygen
C2360416|T201|MTH_LN|51733-4|LNC|oxygen|oxygen
C2360416|T201|LC|51733-4|LNC|oxygen|oxygen
C2360416|T201|OSN|51733-4|LNC|oxygen|oxygen
C2360498|T201|LN|51794-6|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2360498|T201|MTH_LN|51794-6|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2360498|T201|OSN|51794-6|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2360498|T201|LC|51794-6|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2360520|T201|LN|51829-0|LNC|lactate|lactate
C2360520|T201|OSN|51829-0|LNC|lactate|lactate
C2360520|T201|MTH_LN|51829-0|LNC|lactate|lactate
C2360520|T201|LC|51829-0|LNC|lactate|lactate
C2361322|T201|LN|53316-6|LNC|neutrophil count|neutrophil count
C2361322|T201|MTH_LN|53316-6|LNC|neutrophil count|neutrophil count
C2361322|T201|OSN|53316-6|LNC|neutrophil count|neutrophil count
C2361322|T201|LC|53316-6|LNC|neutrophil count|neutrophil count
C2361322|T201|LN|53316-6|LNC|cytology|cytology
C2361322|T201|MTH_LN|53316-6|LNC|cytology|cytology
C2361322|T201|OSN|53316-6|LNC|cytology|cytology
C2361322|T201|LC|53316-6|LNC|cytology|cytology
C2361327|T201|LN|53321-6|LNC|homeostasis|homeostasis
C2361327|T201|MTH_LN|53321-6|LNC|homeostasis|homeostasis
C2361327|T201|OSN|53321-6|LNC|homeostasis|homeostasis
C2361327|T201|LC|53321-6|LNC|homeostasis|homeostasis
C2361444|T201|LN|52958-6|LNC|methadone test|methadone test
C2361444|T201|MTH_LN|52958-6|LNC|methadone test|methadone test
C2361444|T201|OSN|52958-6|LNC|methadone test|methadone test
C2361444|T201|LC|52958-6|LNC|methadone test|methadone test
C2361549|T201|LN|53061-8|LNC|ketone bodies|ketone bodies
C2361549|T201|OSN|53061-8|LNC|ketone bodies|ketone bodies
C2361549|T201|MTH_LN|53061-8|LNC|ketone bodies|ketone bodies
C2361549|T201|LC|53061-8|LNC|ketone bodies|ketone bodies
C2361616|T201|LN|53133-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2361616|T201|MTH_LN|53133-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2361616|T201|OSN|53133-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2361616|T201|LC|53133-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2361616|T201|LN|53133-5|LNC|LDL|LDL
C2361616|T201|MTH_LN|53133-5|LNC|LDL|LDL
C2361616|T201|OSN|53133-5|LNC|LDL|LDL
C2361616|T201|LC|53133-5|LNC|LDL|LDL
C2361616|T201|LN|53133-5|LNC|LDL cholesterol|LDL cholesterol
C2361616|T201|MTH_LN|53133-5|LNC|LDL cholesterol|LDL cholesterol
C2361616|T201|OSN|53133-5|LNC|LDL cholesterol|LDL cholesterol
C2361616|T201|LC|53133-5|LNC|LDL cholesterol|LDL cholesterol
C2361616|T201|LN|53133-5|LNC|low-density lipoprotein|low-density lipoprotein
C2361616|T201|MTH_LN|53133-5|LNC|low-density lipoprotein|low-density lipoprotein
C2361616|T201|OSN|53133-5|LNC|low-density lipoprotein|low-density lipoprotein
C2361616|T201|LC|53133-5|LNC|low-density lipoprotein|low-density lipoprotein
C2361616|T201|LN|53133-5|LNC|beta-lipoproteins|beta-lipoproteins
C2361616|T201|MTH_LN|53133-5|LNC|beta-lipoproteins|beta-lipoproteins
C2361616|T201|OSN|53133-5|LNC|beta-lipoproteins|beta-lipoproteins
C2361616|T201|LC|53133-5|LNC|beta-lipoproteins|beta-lipoproteins
C2361616|T201|LN|53133-5|LNC|LDL-C|LDL-C
C2361616|T201|MTH_LN|53133-5|LNC|LDL-C|LDL-C
C2361616|T201|OSN|53133-5|LNC|LDL-C|LDL-C
C2361616|T201|LC|53133-5|LNC|LDL-C|LDL-C
C2361628|T201|LN|53145-9|LNC|luteinizing|luteinizing
C2361628|T201|OSN|53145-9|LNC|luteinizing|luteinizing
C2361628|T201|MTH_LN|53145-9|LNC|luteinizing|luteinizing
C2361628|T201|LC|53145-9|LNC|luteinizing|luteinizing
C2361628|T201|LN|53145-9|LNC|LH|LH
C2361628|T201|OSN|53145-9|LNC|LH|LH
C2361628|T201|MTH_LN|53145-9|LNC|LH|LH
C2361628|T201|LC|53145-9|LNC|LH|LH
C2361628|T201|LN|53145-9|LNC|luteinising|luteinising
C2361628|T201|OSN|53145-9|LNC|luteinising|luteinising
C2361628|T201|MTH_LN|53145-9|LNC|luteinising|luteinising
C2361628|T201|LC|53145-9|LNC|luteinising|luteinising
// C2361818|T201|LN|53292-9|LNC||
// C2361818|T201|MTH_LN|53292-9|LNC||
// C2361818|T201|OSN|53292-9|LNC||
// C2361818|T201|LC|53292-9|LNC||
C2361818|T201|LN|53292-9|LNC|occult|occult
C2361818|T201|MTH_LN|53292-9|LNC|occult|occult
C2361818|T201|OSN|53292-9|LNC|occult|occult
C2361818|T201|LC|53292-9|LNC|occult|occult
C2361846|T201|LN|53326-5|LNC|osmolality|osmolality
C2361846|T201|MTH_LN|53326-5|LNC|osmolality|osmolality
C2361846|T201|OSN|53326-5|LNC|osmolality|osmolality
C2361846|T201|LC|53326-5|LNC|osmolality|osmolality
C2361846|T201|LN|53326-5|LNC|homeostasis|homeostasis
C2361846|T201|MTH_LN|53326-5|LNC|homeostasis|homeostasis
C2361846|T201|OSN|53326-5|LNC|homeostasis|homeostasis
C2361846|T201|LC|53326-5|LNC|homeostasis|homeostasis
C2361881|T201|LN|53358-8|LNC|y|y
C2361881|T201|MTH_LN|53358-8|LNC|y|y
C2361881|T201|OSN|53358-8|LNC|y|y
C2361881|T201|LC|53358-8|LNC|y|y
C2361883|T201|LN|53360-4|LNC|y|y
C2361883|T201|MTH_LN|53360-4|LNC|y|y
C2361883|T201|OSN|53360-4|LNC|y|y
C2361883|T201|LC|53360-4|LNC|y|y
C2363250|T201|MTH_LN|35214-6|LNC|iron|iron
C2363250|T201|LN|35214-6|LNC|iron|iron
C2363250|T201|OSN|35214-6|LNC|iron|iron
C2363250|T201|LC|35214-6|LNC|iron|iron
C2363268|T201|MTH_LN|35233-6|LNC|urate|urate
C2363268|T201|OSN|35233-6|LNC|urate|urate
C2363268|T201|LN|35233-6|LNC|urate|urate
C2363268|T201|LC|35233-6|LNC|urate|urate
C2363268|T201|MTH_LN|35233-6|LNC|uric acid|uric acid
C2363268|T201|OSN|35233-6|LNC|uric acid|uric acid
C2363268|T201|LN|35233-6|LNC|uric acid|uric acid
C2363268|T201|LC|35233-6|LNC|uric acid|uric acid
C2363271|T201|MTH_LN|35236-9|LNC|urobilinogen|urobilinogen
C2363271|T201|OSN|35236-9|LNC|urobilinogen|urobilinogen
C2363271|T201|LN|35236-9|LNC|urobilinogen|urobilinogen
C2363271|T201|LC|35236-9|LNC|urobilinogen|urobilinogen
C2363286|T201|MTH_LN|35232-8|LNC|uric acid|uric acid
C2363286|T201|LN|35232-8|LNC|uric acid|uric acid
C2363286|T201|OSN|35232-8|LNC|uric acid|uric acid
C2363286|T201|LC|35232-8|LNC|uric acid|uric acid
C2363286|T201|MTH_LN|35232-8|LNC|purine metabolism|purine metabolism
C2363286|T201|LN|35232-8|LNC|purine metabolism|purine metabolism
C2363286|T201|OSN|35232-8|LNC|purine metabolism|purine metabolism
C2363286|T201|LC|35232-8|LNC|purine metabolism|purine metabolism
C2363327|T201|MTH_LN|26513-2|LNC|neutrophil counts|neutrophil counts
C2363327|T201|OSN|26513-2|LNC|neutrophil counts|neutrophil counts
C2363327|T201|LN|26513-2|LNC|neutrophil counts|neutrophil counts
C2363327|T201|LC|26513-2|LNC|neutrophil counts|neutrophil counts
C2363327|T201|MTH_LN|26513-2|LNC|neutrophil count|neutrophil count
C2363327|T201|OSN|26513-2|LNC|neutrophil count|neutrophil count
C2363327|T201|LN|26513-2|LNC|neutrophil count|neutrophil count
C2363327|T201|LC|26513-2|LNC|neutrophil count|neutrophil count
C2363327|T201|MTH_LN|26513-2|LNC|neutrophil|neutrophil
C2363327|T201|OSN|26513-2|LNC|neutrophil|neutrophil
C2363327|T201|LN|26513-2|LNC|neutrophil|neutrophil
C2363327|T201|LC|26513-2|LNC|neutrophil|neutrophil
C2363361|T201|MTH_LN|35245-0|LNC|lactate|lactate
C2363361|T201|LN|35245-0|LNC|lactate|lactate
C2363361|T201|OSN|35245-0|LNC|lactate|lactate
C2363361|T201|LC|35245-0|LNC|lactate|lactate
C2363362|T201|MTH_LN|35253-4|LNC|urate|urate
C2363362|T201|OSN|35253-4|LNC|urate|urate
C2363362|T201|LN|35253-4|LNC|urate|urate
C2363362|T201|LC|35253-4|LNC|urate|urate
C2363362|T201|MTH_LN|35253-4|LNC|uric acid|uric acid
C2363362|T201|OSN|35253-4|LNC|uric acid|uric acid
C2363362|T201|LN|35253-4|LNC|uric acid|uric acid
C2363362|T201|LC|35253-4|LNC|uric acid|uric acid
C2598498|T201|LN|53964-3|LNC|neutrophil count|neutrophil count
C2598498|T201|MTH_LN|53964-3|LNC|neutrophil count|neutrophil count
C2598498|T201|LC|53964-3|LNC|neutrophil count|neutrophil count
C2598498|T201|OSN|53964-3|LNC|neutrophil count|neutrophil count
C2598498|T201|LN|53964-3|LNC|cytology|cytology
C2598498|T201|MTH_LN|53964-3|LNC|cytology|cytology
C2598498|T201|LC|53964-3|LNC|cytology|cytology
C2598498|T201|OSN|53964-3|LNC|cytology|cytology
C2598649|T201|LN|53531-0|LNC|albumin|albumin
C2598649|T201|MTH_LN|53531-0|LNC|albumin|albumin
C2598649|T201|OSN|53531-0|LNC|albumin|albumin
C2598649|T201|LC|53531-0|LNC|albumin|albumin
C2599044|T201|LN|53835-5|LNC|1,5 anhydroglucitol|1,5 anhydroglucitol
C2599044|T201|LC|53835-5|LNC|1,5 anhydroglucitol|1,5 anhydroglucitol
C2599044|T201|OSN|53835-5|LNC|1,5 anhydroglucitol|1,5 anhydroglucitol
C2599044|T201|MTH_LN|53835-5|LNC|1,5 anhydroglucitol|1,5 anhydroglucitol
C2599044|T201|LN|53835-5|LNC|1,5-anhydroglucitol|1,5-anhydroglucitol
C2599044|T201|LC|53835-5|LNC|1,5-anhydroglucitol|1,5-anhydroglucitol
C2599044|T201|OSN|53835-5|LNC|1,5-anhydroglucitol|1,5-anhydroglucitol
C2599044|T201|MTH_LN|53835-5|LNC|1,5-anhydroglucitol|1,5-anhydroglucitol
C2599044|T201|LN|53835-5|LNC|1,5-anhydro-D-glucitol|1,5-anhydro-D-glucitol
C2599044|T201|LC|53835-5|LNC|1,5-anhydro-D-glucitol|1,5-anhydro-D-glucitol
C2599044|T201|OSN|53835-5|LNC|1,5-anhydro-D-glucitol|1,5-anhydro-D-glucitol
C2599044|T201|MTH_LN|53835-5|LNC|1,5-anhydro-D-glucitol|1,5-anhydro-D-glucitol
C2599044|T201|LN|53835-5|LNC|1,5-AG|1,5-AG
C2599044|T201|LC|53835-5|LNC|1,5-AG|1,5-AG
C2599044|T201|OSN|53835-5|LNC|1,5-AG|1,5-AG
C2599044|T201|MTH_LN|53835-5|LNC|1,5-AG|1,5-AG
C2599167|T201|LN|53919-7|LNC|Autoimmune antibody|Autoimmune antibody
C2599167|T201|MTH_LN|53919-7|LNC|Autoimmune antibody|Autoimmune antibody
C2599167|T201|OSN|53919-7|LNC|Autoimmune antibody|Autoimmune antibody
C2599167|T201|LC|53919-7|LNC|Autoimmune antibody|Autoimmune antibody
C2599169|T201|LN|53921-3|LNC|Autoimmune antibody|Autoimmune antibody
C2599169|T201|MTH_LN|53921-3|LNC|Autoimmune antibody|Autoimmune antibody
C2599169|T201|LC|53921-3|LNC|Autoimmune antibody|Autoimmune antibody
C2599169|T201|OSN|53921-3|LNC|Autoimmune antibody|Autoimmune antibody
C2603387|T201|MTH_LN|35197-3|LNC|HDL cholesterol|HDL cholesterol
C2603387|T201|LN|35197-3|LNC|HDL cholesterol|HDL cholesterol
C2603387|T201|OSN|35197-3|LNC|HDL cholesterol|HDL cholesterol
C2603387|T201|LC|35197-3|LNC|HDL cholesterol|HDL cholesterol
C2603387|T201|MTH_LN|35197-3|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C2603387|T201|LN|35197-3|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C2603387|T201|OSN|35197-3|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C2603387|T201|LC|35197-3|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C2603387|T201|MTH_LN|35197-3|LNC|HDL-cholesterol|HDL-cholesterol
C2603387|T201|LN|35197-3|LNC|HDL-cholesterol|HDL-cholesterol
C2603387|T201|OSN|35197-3|LNC|HDL-cholesterol|HDL-cholesterol
C2603387|T201|LC|35197-3|LNC|HDL-cholesterol|HDL-cholesterol
C2603387|T201|MTH_LN|35197-3|LNC|high-density lipoprotein|high-density lipoprotein
C2603387|T201|LN|35197-3|LNC|high-density lipoprotein|high-density lipoprotein
C2603387|T201|OSN|35197-3|LNC|high-density lipoprotein|high-density lipoprotein
C2603387|T201|LC|35197-3|LNC|high-density lipoprotein|high-density lipoprotein
C2603387|T201|MTH_LN|35197-3|LNC|HDL|HDL
C2603387|T201|LN|35197-3|LNC|HDL|HDL
C2603387|T201|OSN|35197-3|LNC|HDL|HDL
C2603387|T201|LC|35197-3|LNC|HDL|HDL
C2603388|T201|MTH_LN|35198-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2603388|T201|LN|35198-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2603388|T201|OSN|35198-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2603388|T201|LC|35198-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2603388|T201|MTH_LN|35198-1|LNC|LDL|LDL
C2603388|T201|LN|35198-1|LNC|LDL|LDL
C2603388|T201|OSN|35198-1|LNC|LDL|LDL
C2603388|T201|LC|35198-1|LNC|LDL|LDL
C2603388|T201|MTH_LN|35198-1|LNC|LDL cholesterol|LDL cholesterol
C2603388|T201|LN|35198-1|LNC|LDL cholesterol|LDL cholesterol
C2603388|T201|OSN|35198-1|LNC|LDL cholesterol|LDL cholesterol
C2603388|T201|LC|35198-1|LNC|LDL cholesterol|LDL cholesterol
C2603388|T201|MTH_LN|35198-1|LNC|low-density lipoprotein|low-density lipoprotein
C2603388|T201|LN|35198-1|LNC|low-density lipoprotein|low-density lipoprotein
C2603388|T201|OSN|35198-1|LNC|low-density lipoprotein|low-density lipoprotein
C2603388|T201|LC|35198-1|LNC|low-density lipoprotein|low-density lipoprotein
C2603388|T201|MTH_LN|35198-1|LNC|beta-lipoproteins|beta-lipoproteins
C2603388|T201|LN|35198-1|LNC|beta-lipoproteins|beta-lipoproteins
C2603388|T201|OSN|35198-1|LNC|beta-lipoproteins|beta-lipoproteins
C2603388|T201|LC|35198-1|LNC|beta-lipoproteins|beta-lipoproteins
C2603388|T201|MTH_LN|35198-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C2603388|T201|LN|35198-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C2603388|T201|OSN|35198-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C2603388|T201|LC|35198-1|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C2603388|T201|MTH_LN|35198-1|LNC|LDL-C|LDL-C
C2603388|T201|LN|35198-1|LNC|LDL-C|LDL-C
C2603388|T201|OSN|35198-1|LNC|LDL-C|LDL-C
C2603388|T201|LC|35198-1|LNC|LDL-C|LDL-C
C2603389|T201|MTH_LN|35199-9|LNC|VLDL cholesterol|VLDL cholesterol
C2603389|T201|LN|35199-9|LNC|VLDL cholesterol|VLDL cholesterol
C2603389|T201|OSN|35199-9|LNC|VLDL cholesterol|VLDL cholesterol
C2603389|T201|LC|35199-9|LNC|VLDL cholesterol|VLDL cholesterol
C2603389|T201|MTH_LN|35199-9|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C2603389|T201|LN|35199-9|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C2603389|T201|OSN|35199-9|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C2603389|T201|LC|35199-9|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C2603389|T201|MTH_LN|35199-9|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C2603389|T201|LN|35199-9|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C2603389|T201|OSN|35199-9|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C2603389|T201|LC|35199-9|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C2607829|T201|LC|35209-6|LNC|ferritin|ferritin
C2607829|T201|MTH_LN|35209-6|LNC|ferritin|ferritin
C2607829|T201|LN|35209-6|LNC|ferritin|ferritin
C2607829|T201|OSN|35209-6|LNC|ferritin|ferritin
C2607831|T201|OSN|35210-4|LNC|folate metabolism|folate metabolism
C2607831|T201|LN|35210-4|LNC|folate metabolism|folate metabolism
C2607831|T201|MTH_LN|35210-4|LNC|folate metabolism|folate metabolism
C2607831|T201|LC|35210-4|LNC|folate metabolism|folate metabolism
C2607836|T201|MTH_LN|35211-2|LNC|glucose|glucose
C2607836|T201|LN|35211-2|LNC|glucose|glucose
C2607836|T201|OSN|35211-2|LNC|glucose|glucose
C2607836|T201|LC|35211-2|LNC|glucose|glucose
C2706775|T201|LN|54213-4|LNC|cortisol|cortisol
C2706775|T201|OSN|54213-4|LNC|cortisol|cortisol
C2706775|T201|MTH_LN|54213-4|LNC|cortisol|cortisol
C2706775|T201|LC|54213-4|LNC|cortisol|cortisol
C2706775|T201|LN|54213-4|LNC|cortisol low|cortisol low
C2706775|T201|OSN|54213-4|LNC|cortisol low|cortisol low
C2706775|T201|MTH_LN|54213-4|LNC|cortisol low|cortisol low
C2706775|T201|LC|54213-4|LNC|cortisol low|cortisol low
C2706775|T201|LN|54213-4|LNC|to undetectable cortisol|to undetectable cortisol
C2706775|T201|OSN|54213-4|LNC|to undetectable cortisol|to undetectable cortisol
C2706775|T201|MTH_LN|54213-4|LNC|to undetectable cortisol|to undetectable cortisol
C2706775|T201|LC|54213-4|LNC|to undetectable cortisol|to undetectable cortisol
C2706777|T201|LN|54215-9|LNC|cortisol|cortisol
C2706777|T201|OSN|54215-9|LNC|cortisol|cortisol
C2706777|T201|MTH_LN|54215-9|LNC|cortisol|cortisol
C2706777|T201|LC|54215-9|LNC|cortisol|cortisol
C2706777|T201|LN|54215-9|LNC|cortisol low|cortisol low
C2706777|T201|OSN|54215-9|LNC|cortisol low|cortisol low
C2706777|T201|MTH_LN|54215-9|LNC|cortisol low|cortisol low
C2706777|T201|LC|54215-9|LNC|cortisol low|cortisol low
C2706777|T201|LN|54215-9|LNC|to undetectable cortisol|to undetectable cortisol
C2706777|T201|OSN|54215-9|LNC|to undetectable cortisol|to undetectable cortisol
C2706777|T201|MTH_LN|54215-9|LNC|to undetectable cortisol|to undetectable cortisol
C2706777|T201|LC|54215-9|LNC|to undetectable cortisol|to undetectable cortisol
C2706780|T201|MTH_LN|54218-3|LNC|CD4:CD8 ratio|CD4:CD8 ratio
C2706780|T201|LC|54218-3|LNC|CD4:CD8 ratio|CD4:CD8 ratio
C2706780|T201|LN|54218-3|LNC|CD4:CD8 ratio|CD4:CD8 ratio
C2706780|T201|OSN|54218-3|LNC|CD4:CD8 ratio|CD4:CD8 ratio
C2706800|T201|LN|54237-3|LNC|ACTH|ACTH
C2706800|T201|OSN|54237-3|LNC|ACTH|ACTH
C2706800|T201|LC|54237-3|LNC|ACTH|ACTH
C2706800|T201|MTH_LN|54237-3|LNC|ACTH|ACTH
C2706800|T201|LN|54237-3|LNC|corticotropin|corticotropin
C2706800|T201|OSN|54237-3|LNC|corticotropin|corticotropin
C2706800|T201|LC|54237-3|LNC|corticotropin|corticotropin
C2706800|T201|MTH_LN|54237-3|LNC|corticotropin|corticotropin
C2706800|T201|LN|54237-3|LNC|adrenocorticotropin|adrenocorticotropin
C2706800|T201|OSN|54237-3|LNC|adrenocorticotropin|adrenocorticotropin
C2706800|T201|LC|54237-3|LNC|adrenocorticotropin|adrenocorticotropin
C2706800|T201|MTH_LN|54237-3|LNC|adrenocorticotropin|adrenocorticotropin
C2706875|T201|LN|54309-0|LNC|CSF lactate|CSF lactate
C2706875|T201|OSN|54309-0|LNC|CSF lactate|CSF lactate
C2706875|T201|LC|54309-0|LNC|CSF lactate|CSF lactate
C2706875|T201|MTH_LN|54309-0|LNC|CSF lactate|CSF lactate
C2706875|T201|LN|54309-0|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C2706875|T201|OSN|54309-0|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C2706875|T201|LC|54309-0|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C2706875|T201|MTH_LN|54309-0|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C2706875|T201|LN|54309-0|LNC|CSF lactic acid|CSF lactic acid
C2706875|T201|OSN|54309-0|LNC|CSF lactic acid|CSF lactic acid
C2706875|T201|LC|54309-0|LNC|CSF lactic acid|CSF lactic acid
C2706875|T201|MTH_LN|54309-0|LNC|CSF lactic acid|CSF lactic acid
C2708273|T201|LN|55440-2|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2708273|T201|LC|55440-2|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2708273|T201|OSN|55440-2|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2708273|T201|MTH_LN|55440-2|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2708273|T201|LN|55440-2|LNC|LDL|LDL
C2708273|T201|LC|55440-2|LNC|LDL|LDL
C2708273|T201|OSN|55440-2|LNC|LDL|LDL
C2708273|T201|MTH_LN|55440-2|LNC|LDL|LDL
C2708273|T201|LN|55440-2|LNC|LDL cholesterol|LDL cholesterol
C2708273|T201|LC|55440-2|LNC|LDL cholesterol|LDL cholesterol
C2708273|T201|OSN|55440-2|LNC|LDL cholesterol|LDL cholesterol
C2708273|T201|MTH_LN|55440-2|LNC|LDL cholesterol|LDL cholesterol
C2708273|T201|LN|55440-2|LNC|low-density lipoprotein|low-density lipoprotein
C2708273|T201|LC|55440-2|LNC|low-density lipoprotein|low-density lipoprotein
C2708273|T201|OSN|55440-2|LNC|low-density lipoprotein|low-density lipoprotein
C2708273|T201|MTH_LN|55440-2|LNC|low-density lipoprotein|low-density lipoprotein
C2708273|T201|LN|55440-2|LNC|beta-lipoproteins|beta-lipoproteins
C2708273|T201|LC|55440-2|LNC|beta-lipoproteins|beta-lipoproteins
C2708273|T201|OSN|55440-2|LNC|beta-lipoproteins|beta-lipoproteins
C2708273|T201|MTH_LN|55440-2|LNC|beta-lipoproteins|beta-lipoproteins
C2708273|T201|LN|55440-2|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C2708273|T201|LC|55440-2|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C2708273|T201|OSN|55440-2|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C2708273|T201|MTH_LN|55440-2|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C2708273|T201|LN|55440-2|LNC|LDL-C|LDL-C
C2708273|T201|LC|55440-2|LNC|LDL-C|LDL-C
C2708273|T201|OSN|55440-2|LNC|LDL-C|LDL-C
C2708273|T201|MTH_LN|55440-2|LNC|LDL-C|LDL-C
C2708749|T201|LN|55469-1|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C2708749|T201|MTH_LN|55469-1|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C2708749|T201|OSN|55469-1|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C2708749|T201|LC|55469-1|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C2708749|T201|LN|55469-1|LNC|17-OHP|17-OHP
C2708749|T201|MTH_LN|55469-1|LNC|17-OHP|17-OHP
C2708749|T201|OSN|55469-1|LNC|17-OHP|17-OHP
C2708749|T201|LC|55469-1|LNC|17-OHP|17-OHP
C2708750|T201|LN|55470-9|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C2708750|T201|MTH_LN|55470-9|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C2708750|T201|OSN|55470-9|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C2708750|T201|LC|55470-9|LNC|17-hydroxyprogesterone|17-hydroxyprogesterone
C2708750|T201|LN|55470-9|LNC|17-OHP|17-OHP
C2708750|T201|MTH_LN|55470-9|LNC|17-OHP|17-OHP
C2708750|T201|OSN|55470-9|LNC|17-OHP|17-OHP
C2708750|T201|LC|55470-9|LNC|17-OHP|17-OHP
C2708781|T201|LN|55501-1|LNC|luteinizing|luteinizing
C2708781|T201|LC|55501-1|LNC|luteinizing|luteinizing
C2708781|T201|OSN|55501-1|LNC|luteinizing|luteinizing
C2708781|T201|MTH_LN|55501-1|LNC|luteinizing|luteinizing
C2708781|T201|LN|55501-1|LNC|LH|LH
C2708781|T201|LC|55501-1|LNC|LH|LH
C2708781|T201|OSN|55501-1|LNC|LH|LH
C2708781|T201|MTH_LN|55501-1|LNC|LH|LH
C2708781|T201|LN|55501-1|LNC|luteinising|luteinising
C2708781|T201|LC|55501-1|LNC|luteinising|luteinising
C2708781|T201|OSN|55501-1|LNC|luteinising|luteinising
C2708781|T201|MTH_LN|55501-1|LNC|luteinising|luteinising
C2708824|T201|LN|55559-9|LNC|xenobiotic|xenobiotic
C2708824|T201|OSN|55559-9|LNC|xenobiotic|xenobiotic
C2708824|T201|MTH_LN|55559-9|LNC|xenobiotic|xenobiotic
C2708824|T201|LC|55559-9|LNC|xenobiotic|xenobiotic
C2713261|T201|OLC|2086-7|LNC|HDL cholesterol|HDL cholesterol
C2713261|T201|MTH_LO|2086-7|LNC|HDL cholesterol|HDL cholesterol
C2713261|T201|LO|2086-7|LNC|HDL cholesterol|HDL cholesterol
C2713261|T201|OOSN|2086-7|LNC|HDL cholesterol|HDL cholesterol
C2713261|T201|OLC|2086-7|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C2713261|T201|MTH_LO|2086-7|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C2713261|T201|LO|2086-7|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C2713261|T201|OOSN|2086-7|LNC|high-density lipoprotein cholesterol|high-density lipoprotein cholesterol
C2713261|T201|OLC|2086-7|LNC|HDL-cholesterol|HDL-cholesterol
C2713261|T201|MTH_LO|2086-7|LNC|HDL-cholesterol|HDL-cholesterol
C2713261|T201|LO|2086-7|LNC|HDL-cholesterol|HDL-cholesterol
C2713261|T201|OOSN|2086-7|LNC|HDL-cholesterol|HDL-cholesterol
C2713261|T201|OLC|2086-7|LNC|high-density lipoprotein|high-density lipoprotein
C2713261|T201|MTH_LO|2086-7|LNC|high-density lipoprotein|high-density lipoprotein
C2713261|T201|LO|2086-7|LNC|high-density lipoprotein|high-density lipoprotein
C2713261|T201|OOSN|2086-7|LNC|high-density lipoprotein|high-density lipoprotein
C2713261|T201|OLC|2086-7|LNC|HDL|HDL
C2713261|T201|MTH_LO|2086-7|LNC|HDL|HDL
C2713261|T201|LO|2086-7|LNC|HDL|HDL
C2713261|T201|OOSN|2086-7|LNC|HDL|HDL
C2733675|T201|LN|55781-9|LNC|hematocrit|hematocrit
C2733675|T201|MTH_LN|55781-9|LNC|hematocrit|hematocrit
C2733675|T201|LC|55781-9|LNC|hematocrit|hematocrit
C2733675|T201|OSN|55781-9|LNC|hematocrit|hematocrit
C2733831|T201|LN|55859-3|LNC|folate metabolism|folate metabolism
C2733831|T201|OSN|55859-3|LNC|folate metabolism|folate metabolism
C2733831|T201|LC|55859-3|LNC|folate metabolism|folate metabolism
C2733831|T201|MTH_LN|55859-3|LNC|folate metabolism|folate metabolism
C2733887|T201|LN|55918-7|LNC|C-peptide|C-peptide
C2733887|T201|OSN|55918-7|LNC|C-peptide|C-peptide
C2733887|T201|LC|55918-7|LNC|C-peptide|C-peptide
C2733887|T201|MTH_LN|55918-7|LNC|C-peptide|C-peptide
C2733887|T201|LN|55918-7|LNC|C peptide|C peptide
C2733887|T201|OSN|55918-7|LNC|C peptide|C peptide
C2733887|T201|LC|55918-7|LNC|C peptide|C peptide
C2733887|T201|MTH_LN|55918-7|LNC|C peptide|C peptide
C2733888|T201|LN|55919-5|LNC|C-peptide|C-peptide
C2733888|T201|OSN|55919-5|LNC|C-peptide|C-peptide
C2733888|T201|LC|55919-5|LNC|C-peptide|C-peptide
C2733888|T201|MTH_LN|55919-5|LNC|C-peptide|C-peptide
C2733888|T201|LN|55919-5|LNC|C peptide|C peptide
C2733888|T201|OSN|55919-5|LNC|C peptide|C peptide
C2733888|T201|LC|55919-5|LNC|C peptide|C peptide
C2733888|T201|MTH_LN|55919-5|LNC|C peptide|C peptide
C2733903|T201|LN|55932-8|LNC|lactate|lactate
C2733903|T201|LC|55932-8|LNC|lactate|lactate
C2733903|T201|OSN|55932-8|LNC|lactate|lactate
C2733903|T201|MTH_LN|55932-8|LNC|lactate|lactate
C2734094|T201|LN|56136-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734094|T201|LC|56136-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734094|T201|OSN|56136-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734094|T201|MTH_LN|56136-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734094|T201|LN|56136-5|LNC|LDL|LDL
C2734094|T201|LC|56136-5|LNC|LDL|LDL
C2734094|T201|OSN|56136-5|LNC|LDL|LDL
C2734094|T201|MTH_LN|56136-5|LNC|LDL|LDL
C2734094|T201|LN|56136-5|LNC|LDL cholesterol|LDL cholesterol
C2734094|T201|LC|56136-5|LNC|LDL cholesterol|LDL cholesterol
C2734094|T201|OSN|56136-5|LNC|LDL cholesterol|LDL cholesterol
C2734094|T201|MTH_LN|56136-5|LNC|LDL cholesterol|LDL cholesterol
C2734094|T201|LN|56136-5|LNC|low-density lipoprotein|low-density lipoprotein
C2734094|T201|LC|56136-5|LNC|low-density lipoprotein|low-density lipoprotein
C2734094|T201|OSN|56136-5|LNC|low-density lipoprotein|low-density lipoprotein
C2734094|T201|MTH_LN|56136-5|LNC|low-density lipoprotein|low-density lipoprotein
C2734094|T201|LN|56136-5|LNC|beta-lipoproteins|beta-lipoproteins
C2734094|T201|LC|56136-5|LNC|beta-lipoproteins|beta-lipoproteins
C2734094|T201|OSN|56136-5|LNC|beta-lipoproteins|beta-lipoproteins
C2734094|T201|MTH_LN|56136-5|LNC|beta-lipoproteins|beta-lipoproteins
C2734094|T201|LN|56136-5|LNC|LDL-C|LDL-C
C2734094|T201|LC|56136-5|LNC|LDL-C|LDL-C
C2734094|T201|OSN|56136-5|LNC|LDL-C|LDL-C
C2734094|T201|MTH_LN|56136-5|LNC|LDL-C|LDL-C
C2734095|T201|LN|56137-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734095|T201|OSN|56137-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734095|T201|LC|56137-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734095|T201|MTH_LN|56137-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734095|T201|LN|56137-3|LNC|LDL|LDL
C2734095|T201|OSN|56137-3|LNC|LDL|LDL
C2734095|T201|LC|56137-3|LNC|LDL|LDL
C2734095|T201|MTH_LN|56137-3|LNC|LDL|LDL
C2734095|T201|LN|56137-3|LNC|LDL cholesterol|LDL cholesterol
C2734095|T201|OSN|56137-3|LNC|LDL cholesterol|LDL cholesterol
C2734095|T201|LC|56137-3|LNC|LDL cholesterol|LDL cholesterol
C2734095|T201|MTH_LN|56137-3|LNC|LDL cholesterol|LDL cholesterol
C2734095|T201|LN|56137-3|LNC|low-density lipoprotein|low-density lipoprotein
C2734095|T201|OSN|56137-3|LNC|low-density lipoprotein|low-density lipoprotein
C2734095|T201|LC|56137-3|LNC|low-density lipoprotein|low-density lipoprotein
C2734095|T201|MTH_LN|56137-3|LNC|low-density lipoprotein|low-density lipoprotein
C2734095|T201|LN|56137-3|LNC|beta-lipoproteins|beta-lipoproteins
C2734095|T201|OSN|56137-3|LNC|beta-lipoproteins|beta-lipoproteins
C2734095|T201|LC|56137-3|LNC|beta-lipoproteins|beta-lipoproteins
C2734095|T201|MTH_LN|56137-3|LNC|beta-lipoproteins|beta-lipoproteins
C2734095|T201|LN|56137-3|LNC|LDL-C|LDL-C
C2734095|T201|OSN|56137-3|LNC|LDL-C|LDL-C
C2734095|T201|LC|56137-3|LNC|LDL-C|LDL-C
C2734095|T201|MTH_LN|56137-3|LNC|LDL-C|LDL-C
C2734096|T201|LN|56138-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734096|T201|LC|56138-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734096|T201|MTH_LN|56138-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734096|T201|OSN|56138-1|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734096|T201|LN|56138-1|LNC|LDL|LDL
C2734096|T201|LC|56138-1|LNC|LDL|LDL
C2734096|T201|MTH_LN|56138-1|LNC|LDL|LDL
C2734096|T201|OSN|56138-1|LNC|LDL|LDL
C2734096|T201|LN|56138-1|LNC|LDL cholesterol|LDL cholesterol
C2734096|T201|LC|56138-1|LNC|LDL cholesterol|LDL cholesterol
C2734096|T201|MTH_LN|56138-1|LNC|LDL cholesterol|LDL cholesterol
C2734096|T201|OSN|56138-1|LNC|LDL cholesterol|LDL cholesterol
C2734096|T201|LN|56138-1|LNC|low-density lipoprotein|low-density lipoprotein
C2734096|T201|LC|56138-1|LNC|low-density lipoprotein|low-density lipoprotein
C2734096|T201|MTH_LN|56138-1|LNC|low-density lipoprotein|low-density lipoprotein
C2734096|T201|OSN|56138-1|LNC|low-density lipoprotein|low-density lipoprotein
C2734096|T201|LN|56138-1|LNC|beta-lipoproteins|beta-lipoproteins
C2734096|T201|LC|56138-1|LNC|beta-lipoproteins|beta-lipoproteins
C2734096|T201|MTH_LN|56138-1|LNC|beta-lipoproteins|beta-lipoproteins
C2734096|T201|OSN|56138-1|LNC|beta-lipoproteins|beta-lipoproteins
C2734096|T201|LN|56138-1|LNC|LDL-C|LDL-C
C2734096|T201|LC|56138-1|LNC|LDL-C|LDL-C
C2734096|T201|MTH_LN|56138-1|LNC|LDL-C|LDL-C
C2734096|T201|OSN|56138-1|LNC|LDL-C|LDL-C
C2734097|T201|LN|56139-9|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734097|T201|LC|56139-9|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734097|T201|MTH_LN|56139-9|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734097|T201|OSN|56139-9|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2734097|T201|LN|56139-9|LNC|LDL|LDL
C2734097|T201|LC|56139-9|LNC|LDL|LDL
C2734097|T201|MTH_LN|56139-9|LNC|LDL|LDL
C2734097|T201|OSN|56139-9|LNC|LDL|LDL
C2734097|T201|LN|56139-9|LNC|LDL cholesterol|LDL cholesterol
C2734097|T201|LC|56139-9|LNC|LDL cholesterol|LDL cholesterol
C2734097|T201|MTH_LN|56139-9|LNC|LDL cholesterol|LDL cholesterol
C2734097|T201|OSN|56139-9|LNC|LDL cholesterol|LDL cholesterol
C2734097|T201|LN|56139-9|LNC|low-density lipoprotein|low-density lipoprotein
C2734097|T201|LC|56139-9|LNC|low-density lipoprotein|low-density lipoprotein
C2734097|T201|MTH_LN|56139-9|LNC|low-density lipoprotein|low-density lipoprotein
C2734097|T201|OSN|56139-9|LNC|low-density lipoprotein|low-density lipoprotein
C2734097|T201|LN|56139-9|LNC|beta-lipoproteins|beta-lipoproteins
C2734097|T201|LC|56139-9|LNC|beta-lipoproteins|beta-lipoproteins
C2734097|T201|MTH_LN|56139-9|LNC|beta-lipoproteins|beta-lipoproteins
C2734097|T201|OSN|56139-9|LNC|beta-lipoproteins|beta-lipoproteins
C2734097|T201|LN|56139-9|LNC|LDL-C|LDL-C
C2734097|T201|LC|56139-9|LNC|LDL-C|LDL-C
C2734097|T201|MTH_LN|56139-9|LNC|LDL-C|LDL-C
C2734097|T201|OSN|56139-9|LNC|LDL-C|LDL-C
C2734587|T201|LN|56493-0|LNC|luteinizing|luteinizing
C2734587|T201|LC|56493-0|LNC|luteinizing|luteinizing
C2734587|T201|MTH_LN|56493-0|LNC|luteinizing|luteinizing
C2734587|T201|OSN|56493-0|LNC|luteinizing|luteinizing
C2734587|T201|LN|56493-0|LNC|LH|LH
C2734587|T201|LC|56493-0|LNC|LH|LH
C2734587|T201|MTH_LN|56493-0|LNC|LH|LH
C2734587|T201|OSN|56493-0|LNC|LH|LH
C2734587|T201|LN|56493-0|LNC|luteinising|luteinising
C2734587|T201|LC|56493-0|LNC|luteinising|luteinising
C2734587|T201|MTH_LN|56493-0|LNC|luteinising|luteinising
C2734587|T201|OSN|56493-0|LNC|luteinising|luteinising
C2734588|T201|LN|56494-8|LNC|luteinizing|luteinizing
C2734588|T201|OSN|56494-8|LNC|luteinizing|luteinizing
C2734588|T201|MTH_LN|56494-8|LNC|luteinizing|luteinizing
C2734588|T201|LC|56494-8|LNC|luteinizing|luteinizing
C2734588|T201|LN|56494-8|LNC|LH|LH
C2734588|T201|OSN|56494-8|LNC|LH|LH
C2734588|T201|MTH_LN|56494-8|LNC|LH|LH
C2734588|T201|LC|56494-8|LNC|LH|LH
C2734588|T201|LN|56494-8|LNC|luteinising|luteinising
C2734588|T201|OSN|56494-8|LNC|luteinising|luteinising
C2734588|T201|MTH_LN|56494-8|LNC|luteinising|luteinising
C2734588|T201|LC|56494-8|LNC|luteinising|luteinising
C2734589|T201|LN|56495-5|LNC|luteinizing|luteinizing
C2734589|T201|MTH_LN|56495-5|LNC|luteinizing|luteinizing
C2734589|T201|LC|56495-5|LNC|luteinizing|luteinizing
C2734589|T201|OSN|56495-5|LNC|luteinizing|luteinizing
C2734589|T201|LN|56495-5|LNC|LH|LH
C2734589|T201|MTH_LN|56495-5|LNC|LH|LH
C2734589|T201|LC|56495-5|LNC|LH|LH
C2734589|T201|OSN|56495-5|LNC|LH|LH
C2734589|T201|LN|56495-5|LNC|luteinising|luteinising
C2734589|T201|MTH_LN|56495-5|LNC|luteinising|luteinising
C2734589|T201|LC|56495-5|LNC|luteinising|luteinising
C2734589|T201|OSN|56495-5|LNC|luteinising|luteinising
C2734598|T201|LN|56504-4|LNC|ACTH|ACTH
C2734598|T201|OSN|56504-4|LNC|ACTH|ACTH
C2734598|T201|MTH_LN|56504-4|LNC|ACTH|ACTH
C2734598|T201|LC|56504-4|LNC|ACTH|ACTH
C2734598|T201|LN|56504-4|LNC|corticotropin|corticotropin
C2734598|T201|OSN|56504-4|LNC|corticotropin|corticotropin
C2734598|T201|MTH_LN|56504-4|LNC|corticotropin|corticotropin
C2734598|T201|LC|56504-4|LNC|corticotropin|corticotropin
C2734598|T201|LN|56504-4|LNC|adrenocorticotropin|adrenocorticotropin
C2734598|T201|OSN|56504-4|LNC|adrenocorticotropin|adrenocorticotropin
C2734598|T201|MTH_LN|56504-4|LNC|adrenocorticotropin|adrenocorticotropin
C2734598|T201|LC|56504-4|LNC|adrenocorticotropin|adrenocorticotropin
C2734599|T201|LN|56505-1|LNC|ACTH|ACTH
C2734599|T201|LC|56505-1|LNC|ACTH|ACTH
C2734599|T201|OSN|56505-1|LNC|ACTH|ACTH
C2734599|T201|MTH_LN|56505-1|LNC|ACTH|ACTH
C2734599|T201|LN|56505-1|LNC|corticotropin|corticotropin
C2734599|T201|LC|56505-1|LNC|corticotropin|corticotropin
C2734599|T201|OSN|56505-1|LNC|corticotropin|corticotropin
C2734599|T201|MTH_LN|56505-1|LNC|corticotropin|corticotropin
C2734599|T201|LN|56505-1|LNC|adrenocorticotropin|adrenocorticotropin
C2734599|T201|LC|56505-1|LNC|adrenocorticotropin|adrenocorticotropin
C2734599|T201|OSN|56505-1|LNC|adrenocorticotropin|adrenocorticotropin
C2734599|T201|MTH_LN|56505-1|LNC|adrenocorticotropin|adrenocorticotropin
C2734600|T201|LN|56506-9|LNC|ACTH|ACTH
C2734600|T201|OSN|56506-9|LNC|ACTH|ACTH
C2734600|T201|MTH_LN|56506-9|LNC|ACTH|ACTH
C2734600|T201|LC|56506-9|LNC|ACTH|ACTH
C2734600|T201|LN|56506-9|LNC|corticotropin|corticotropin
C2734600|T201|OSN|56506-9|LNC|corticotropin|corticotropin
C2734600|T201|MTH_LN|56506-9|LNC|corticotropin|corticotropin
C2734600|T201|LC|56506-9|LNC|corticotropin|corticotropin
C2734600|T201|LN|56506-9|LNC|adrenocorticotropin|adrenocorticotropin
C2734600|T201|OSN|56506-9|LNC|adrenocorticotropin|adrenocorticotropin
C2734600|T201|MTH_LN|56506-9|LNC|adrenocorticotropin|adrenocorticotropin
C2734600|T201|LC|56506-9|LNC|adrenocorticotropin|adrenocorticotropin
C2734609|T201|LN|56516-8|LNC|C-peptide|C-peptide
C2734609|T201|OSN|56516-8|LNC|C-peptide|C-peptide
C2734609|T201|MTH_LN|56516-8|LNC|C-peptide|C-peptide
C2734609|T201|LC|56516-8|LNC|C-peptide|C-peptide
C2734609|T201|LN|56516-8|LNC|C peptide|C peptide
C2734609|T201|OSN|56516-8|LNC|C peptide|C peptide
C2734609|T201|MTH_LN|56516-8|LNC|C peptide|C peptide
C2734609|T201|LC|56516-8|LNC|C peptide|C peptide
C2734629|T201|LN|56536-6|LNC|Autoimmune antibody|Autoimmune antibody
C2734629|T201|LC|56536-6|LNC|Autoimmune antibody|Autoimmune antibody
C2734629|T201|MTH_LN|56536-6|LNC|Autoimmune antibody|Autoimmune antibody
C2734629|T201|OSN|56536-6|LNC|Autoimmune antibody|Autoimmune antibody
C2734748|T201|LN|56582-0|LNC|C-peptide|C-peptide
C2734748|T201|LC|56582-0|LNC|C-peptide|C-peptide
C2734748|T201|OSN|56582-0|LNC|C-peptide|C-peptide
C2734748|T201|MTH_LN|56582-0|LNC|C-peptide|C-peptide
C2734748|T201|LN|56582-0|LNC|C peptide|C peptide
C2734748|T201|LC|56582-0|LNC|C peptide|C peptide
C2734748|T201|OSN|56582-0|LNC|C peptide|C peptide
C2734748|T201|MTH_LN|56582-0|LNC|C peptide|C peptide
C2734749|T201|LN|56583-8|LNC|C-peptide|C-peptide
C2734749|T201|OSN|56583-8|LNC|C-peptide|C-peptide
C2734749|T201|MTH_LN|56583-8|LNC|C-peptide|C-peptide
C2734749|T201|LC|56583-8|LNC|C-peptide|C-peptide
C2734749|T201|LN|56583-8|LNC|C peptide|C peptide
C2734749|T201|OSN|56583-8|LNC|C peptide|C peptide
C2734749|T201|MTH_LN|56583-8|LNC|C peptide|C peptide
C2734749|T201|LC|56583-8|LNC|C peptide|C peptide
C2734750|T201|LN|56584-6|LNC|C-peptide|C-peptide
C2734750|T201|OSN|56584-6|LNC|C-peptide|C-peptide
C2734750|T201|LC|56584-6|LNC|C-peptide|C-peptide
C2734750|T201|MTH_LN|56584-6|LNC|C-peptide|C-peptide
C2734750|T201|LN|56584-6|LNC|C peptide|C peptide
C2734750|T201|OSN|56584-6|LNC|C peptide|C peptide
C2734750|T201|LC|56584-6|LNC|C peptide|C peptide
C2734750|T201|MTH_LN|56584-6|LNC|C peptide|C peptide
C2734787|T201|LN|56632-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2734787|T201|LC|56632-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2734787|T201|MTH_LN|56632-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2734787|T201|OSN|56632-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2734790|T201|LN|56635-6|LNC|Autoimmune antibody|Autoimmune antibody
C2734790|T201|OSN|56635-6|LNC|Autoimmune antibody|Autoimmune antibody
C2734790|T201|MTH_LN|56635-6|LNC|Autoimmune antibody|Autoimmune antibody
C2734790|T201|LC|56635-6|LNC|Autoimmune antibody|Autoimmune antibody
C2734826|T201|LN|56672-9|LNC|arginine|arginine
C2734826|T201|MTH_LN|56672-9|LNC|arginine|arginine
C2734826|T201|LC|56672-9|LNC|arginine|arginine
C2734826|T201|OSN|56672-9|LNC|arginine|arginine
C2734917|T201|LN|57386-5|LNC|urate|urate
C2734917|T201|LC|57386-5|LNC|urate|urate
C2734917|T201|MTH_LN|57386-5|LNC|urate|urate
C2734917|T201|OSN|57386-5|LNC|urate|urate
C2734917|T201|LN|57386-5|LNC|uric acid|uric acid
C2734917|T201|LC|57386-5|LNC|uric acid|uric acid
C2734917|T201|MTH_LN|57386-5|LNC|uric acid|uric acid
C2734917|T201|OSN|57386-5|LNC|uric acid|uric acid
C2734918|T201|LN|57387-3|LNC|urate|urate
C2734918|T201|LC|57387-3|LNC|urate|urate
C2734918|T201|OSN|57387-3|LNC|urate|urate
C2734918|T201|MTH_LN|57387-3|LNC|urate|urate
C2734918|T201|LN|57387-3|LNC|uric acid|uric acid
C2734918|T201|LC|57387-3|LNC|uric acid|uric acid
C2734918|T201|OSN|57387-3|LNC|uric acid|uric acid
C2734918|T201|MTH_LN|57387-3|LNC|uric acid|uric acid
C2734953|T201|LN|56735-4|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2734953|T201|MTH_LN|56735-4|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2734953|T201|LC|56735-4|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2734953|T201|OSN|56735-4|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C2735191|T201|LN|56913-7|LNC|ACTH|ACTH
C2735191|T201|LC|56913-7|LNC|ACTH|ACTH
C2735191|T201|MTH_LN|56913-7|LNC|ACTH|ACTH
C2735191|T201|OSN|56913-7|LNC|ACTH|ACTH
C2735191|T201|LN|56913-7|LNC|corticotropin|corticotropin
C2735191|T201|LC|56913-7|LNC|corticotropin|corticotropin
C2735191|T201|MTH_LN|56913-7|LNC|corticotropin|corticotropin
C2735191|T201|OSN|56913-7|LNC|corticotropin|corticotropin
C2735191|T201|LN|56913-7|LNC|adrenocorticotropin|adrenocorticotropin
C2735191|T201|LC|56913-7|LNC|adrenocorticotropin|adrenocorticotropin
C2735191|T201|MTH_LN|56913-7|LNC|adrenocorticotropin|adrenocorticotropin
C2735191|T201|OSN|56913-7|LNC|adrenocorticotropin|adrenocorticotropin
C2735192|T201|LN|56914-5|LNC|ACTH|ACTH
C2735192|T201|OSN|56914-5|LNC|ACTH|ACTH
C2735192|T201|MTH_LN|56914-5|LNC|ACTH|ACTH
C2735192|T201|LC|56914-5|LNC|ACTH|ACTH
C2735192|T201|LN|56914-5|LNC|corticotropin|corticotropin
C2735192|T201|OSN|56914-5|LNC|corticotropin|corticotropin
C2735192|T201|MTH_LN|56914-5|LNC|corticotropin|corticotropin
C2735192|T201|LC|56914-5|LNC|corticotropin|corticotropin
C2735192|T201|LN|56914-5|LNC|adrenocorticotropin|adrenocorticotropin
C2735192|T201|OSN|56914-5|LNC|adrenocorticotropin|adrenocorticotropin
C2735192|T201|MTH_LN|56914-5|LNC|adrenocorticotropin|adrenocorticotropin
C2735192|T201|LC|56914-5|LNC|adrenocorticotropin|adrenocorticotropin
C2735264|T201|LN|56985-5|LNC|taurine|taurine
C2735264|T201|MTH_LN|56985-5|LNC|taurine|taurine
C2735264|T201|LC|56985-5|LNC|taurine|taurine
C2735264|T201|OSN|56985-5|LNC|taurine|taurine
C2735391|T201|LN|57102-6|LNC|luteinizing|luteinizing
C2735391|T201|OSN|57102-6|LNC|luteinizing|luteinizing
C2735391|T201|LC|57102-6|LNC|luteinizing|luteinizing
C2735391|T201|MTH_LN|57102-6|LNC|luteinizing|luteinizing
C2735391|T201|LN|57102-6|LNC|LH|LH
C2735391|T201|OSN|57102-6|LNC|LH|LH
C2735391|T201|LC|57102-6|LNC|LH|LH
C2735391|T201|MTH_LN|57102-6|LNC|LH|LH
C2735391|T201|LN|57102-6|LNC|luteinising|luteinising
C2735391|T201|OSN|57102-6|LNC|luteinising|luteinising
C2735391|T201|LC|57102-6|LNC|luteinising|luteinising
C2735391|T201|MTH_LN|57102-6|LNC|luteinising|luteinising
C2735392|T201|LN|57103-4|LNC|luteinizing|luteinizing
C2735392|T201|MTH_LN|57103-4|LNC|luteinizing|luteinizing
C2735392|T201|LC|57103-4|LNC|luteinizing|luteinizing
C2735392|T201|OSN|57103-4|LNC|luteinizing|luteinizing
C2735392|T201|LN|57103-4|LNC|LH|LH
C2735392|T201|MTH_LN|57103-4|LNC|LH|LH
C2735392|T201|LC|57103-4|LNC|LH|LH
C2735392|T201|OSN|57103-4|LNC|LH|LH
C2735392|T201|LN|57103-4|LNC|luteinising|luteinising
C2735392|T201|MTH_LN|57103-4|LNC|luteinising|luteinising
C2735392|T201|LC|57103-4|LNC|luteinising|luteinising
C2735392|T201|OSN|57103-4|LNC|luteinising|luteinising
C2735393|T201|LN|57104-2|LNC|luteinizing|luteinizing
C2735393|T201|LC|57104-2|LNC|luteinizing|luteinizing
C2735393|T201|MTH_LN|57104-2|LNC|luteinizing|luteinizing
C2735393|T201|OSN|57104-2|LNC|luteinizing|luteinizing
C2735393|T201|LN|57104-2|LNC|LH|LH
C2735393|T201|LC|57104-2|LNC|LH|LH
C2735393|T201|MTH_LN|57104-2|LNC|LH|LH
C2735393|T201|OSN|57104-2|LNC|LH|LH
C2735393|T201|LN|57104-2|LNC|luteinising|luteinising
C2735393|T201|LC|57104-2|LNC|luteinising|luteinising
C2735393|T201|MTH_LN|57104-2|LNC|luteinising|luteinising
C2735393|T201|OSN|57104-2|LNC|luteinising|luteinising
C2735394|T201|LN|57105-9|LNC|luteinizing|luteinizing
C2735394|T201|LC|57105-9|LNC|luteinizing|luteinizing
C2735394|T201|MTH_LN|57105-9|LNC|luteinizing|luteinizing
C2735394|T201|OSN|57105-9|LNC|luteinizing|luteinizing
C2735394|T201|LN|57105-9|LNC|LH|LH
C2735394|T201|LC|57105-9|LNC|LH|LH
C2735394|T201|MTH_LN|57105-9|LNC|LH|LH
C2735394|T201|OSN|57105-9|LNC|LH|LH
C2735394|T201|LN|57105-9|LNC|luteinising|luteinising
C2735394|T201|LC|57105-9|LNC|luteinising|luteinising
C2735394|T201|MTH_LN|57105-9|LNC|luteinising|luteinising
C2735394|T201|OSN|57105-9|LNC|luteinising|luteinising
C2735395|T201|LN|57106-7|LNC|luteinizing|luteinizing
C2735395|T201|MTH_LN|57106-7|LNC|luteinizing|luteinizing
C2735395|T201|LC|57106-7|LNC|luteinizing|luteinizing
C2735395|T201|OSN|57106-7|LNC|luteinizing|luteinizing
C2735395|T201|LN|57106-7|LNC|LH|LH
C2735395|T201|MTH_LN|57106-7|LNC|LH|LH
C2735395|T201|LC|57106-7|LNC|LH|LH
C2735395|T201|OSN|57106-7|LNC|LH|LH
C2735395|T201|LN|57106-7|LNC|luteinising|luteinising
C2735395|T201|MTH_LN|57106-7|LNC|luteinising|luteinising
C2735395|T201|LC|57106-7|LNC|luteinising|luteinising
C2735395|T201|OSN|57106-7|LNC|luteinising|luteinising
C2735396|T201|LN|57107-5|LNC|luteinizing|luteinizing
C2735396|T201|OSN|57107-5|LNC|luteinizing|luteinizing
C2735396|T201|MTH_LN|57107-5|LNC|luteinizing|luteinizing
C2735396|T201|LC|57107-5|LNC|luteinizing|luteinizing
C2735396|T201|LN|57107-5|LNC|LH|LH
C2735396|T201|OSN|57107-5|LNC|LH|LH
C2735396|T201|MTH_LN|57107-5|LNC|LH|LH
C2735396|T201|LC|57107-5|LNC|LH|LH
C2735396|T201|LN|57107-5|LNC|luteinising|luteinising
C2735396|T201|OSN|57107-5|LNC|luteinising|luteinising
C2735396|T201|MTH_LN|57107-5|LNC|luteinising|luteinising
C2735396|T201|LC|57107-5|LNC|luteinising|luteinising
C2735471|T201|LN|57938-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2735471|T201|LC|57938-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2735471|T201|OSN|57938-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2735471|T201|MTH_LN|57938-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2735471|T201|LN|57938-3|LNC|LDL|LDL
C2735471|T201|LC|57938-3|LNC|LDL|LDL
C2735471|T201|OSN|57938-3|LNC|LDL|LDL
C2735471|T201|MTH_LN|57938-3|LNC|LDL|LDL
C2735471|T201|LN|57938-3|LNC|LDL cholesterol|LDL cholesterol
C2735471|T201|LC|57938-3|LNC|LDL cholesterol|LDL cholesterol
C2735471|T201|OSN|57938-3|LNC|LDL cholesterol|LDL cholesterol
C2735471|T201|MTH_LN|57938-3|LNC|LDL cholesterol|LDL cholesterol
C2735471|T201|LN|57938-3|LNC|low-density lipoprotein|low-density lipoprotein
C2735471|T201|LC|57938-3|LNC|low-density lipoprotein|low-density lipoprotein
C2735471|T201|OSN|57938-3|LNC|low-density lipoprotein|low-density lipoprotein
C2735471|T201|MTH_LN|57938-3|LNC|low-density lipoprotein|low-density lipoprotein
C2735471|T201|LN|57938-3|LNC|beta-lipoproteins|beta-lipoproteins
C2735471|T201|LC|57938-3|LNC|beta-lipoproteins|beta-lipoproteins
C2735471|T201|OSN|57938-3|LNC|beta-lipoproteins|beta-lipoproteins
C2735471|T201|MTH_LN|57938-3|LNC|beta-lipoproteins|beta-lipoproteins
C2735471|T201|LN|57938-3|LNC|LDL-C|LDL-C
C2735471|T201|LC|57938-3|LNC|LDL-C|LDL-C
C2735471|T201|OSN|57938-3|LNC|LDL-C|LDL-C
C2735471|T201|MTH_LN|57938-3|LNC|LDL-C|LDL-C
C2735528|T201|LN|57376-6|LNC|C-peptide|C-peptide
C2735528|T201|MTH_LN|57376-6|LNC|C-peptide|C-peptide
C2735528|T201|LC|57376-6|LNC|C-peptide|C-peptide
C2735528|T201|OSN|57376-6|LNC|C-peptide|C-peptide
C2735528|T201|LN|57376-6|LNC|C peptide|C peptide
C2735528|T201|MTH_LN|57376-6|LNC|C peptide|C peptide
C2735528|T201|LC|57376-6|LNC|C peptide|C peptide
C2735528|T201|OSN|57376-6|LNC|C peptide|C peptide
C2735755|T201|LN|57356-8|LNC|lactate|lactate
C2735755|T201|MTH_LN|57356-8|LNC|lactate|lactate
C2735755|T201|OSN|57356-8|LNC|lactate|lactate
C2735755|T201|LC|57356-8|LNC|lactate|lactate
C2735756|T201|LN|57357-6|LNC|lactate|lactate
C2735756|T201|MTH_LN|57357-6|LNC|lactate|lactate
C2735756|T201|OSN|57357-6|LNC|lactate|lactate
C2735756|T201|LC|57357-6|LNC|lactate|lactate
C2735757|T201|LN|57358-4|LNC|lactate|lactate
C2735757|T201|OSN|57358-4|LNC|lactate|lactate
C2735757|T201|LC|57358-4|LNC|lactate|lactate
C2735757|T201|MTH_LN|57358-4|LNC|lactate|lactate
C2735758|T201|LN|57359-2|LNC|lactate|lactate
C2735758|T201|OSN|57359-2|LNC|lactate|lactate
C2735758|T201|MTH_LN|57359-2|LNC|lactate|lactate
C2735758|T201|LC|57359-2|LNC|lactate|lactate
C2735759|T201|LN|57360-0|LNC|lactate|lactate
C2735759|T201|MTH_LN|57360-0|LNC|lactate|lactate
C2735759|T201|LC|57360-0|LNC|lactate|lactate
C2735759|T201|OSN|57360-0|LNC|lactate|lactate
C2735760|T201|LN|57361-8|LNC|lactate|lactate
C2735760|T201|OSN|57361-8|LNC|lactate|lactate
C2735760|T201|LC|57361-8|LNC|lactate|lactate
C2735760|T201|MTH_LN|57361-8|LNC|lactate|lactate
C2735761|T201|LN|57362-6|LNC|lactate|lactate
C2735761|T201|LC|57362-6|LNC|lactate|lactate
C2735761|T201|OSN|57362-6|LNC|lactate|lactate
C2735761|T201|MTH_LN|57362-6|LNC|lactate|lactate
C2735762|T201|LN|57363-4|LNC|lactate|lactate
C2735762|T201|MTH_LN|57363-4|LNC|lactate|lactate
C2735762|T201|OSN|57363-4|LNC|lactate|lactate
C2735762|T201|LC|57363-4|LNC|lactate|lactate
C2735763|T201|LN|57364-2|LNC|lactate|lactate
C2735763|T201|MTH_LN|57364-2|LNC|lactate|lactate
C2735763|T201|OSN|57364-2|LNC|lactate|lactate
C2735763|T201|LC|57364-2|LNC|lactate|lactate
C2735764|T201|LN|57365-9|LNC|lactate|lactate
C2735764|T201|OSN|57365-9|LNC|lactate|lactate
C2735764|T201|LC|57365-9|LNC|lactate|lactate
C2735764|T201|MTH_LN|57365-9|LNC|lactate|lactate
C2735789|T201|LN|57422-8|LNC|T cell CD40 expression|T cell CD40 expression
C2735789|T201|MTH_LN|57422-8|LNC|T cell CD40 expression|T cell CD40 expression
C2735789|T201|LC|57422-8|LNC|T cell CD40 expression|T cell CD40 expression
C2735789|T201|OSN|57422-8|LNC|T cell CD40 expression|T cell CD40 expression
C2735789|T201|LN|57422-8|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C2735789|T201|MTH_LN|57422-8|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C2735789|T201|LC|57422-8|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C2735789|T201|OSN|57422-8|LNC|lymphocyte surface marker expression|lymphocyte surface marker expression
C2736059|T201|LN|57646-2|LNC|C-peptide|C-peptide
C2736059|T201|OSN|57646-2|LNC|C-peptide|C-peptide
C2736059|T201|MTH_LN|57646-2|LNC|C-peptide|C-peptide
C2736059|T201|LC|57646-2|LNC|C-peptide|C-peptide
C2736059|T201|LN|57646-2|LNC|C peptide|C peptide
C2736059|T201|OSN|57646-2|LNC|C peptide|C peptide
C2736059|T201|MTH_LN|57646-2|LNC|C peptide|C peptide
C2736059|T201|LC|57646-2|LNC|C peptide|C peptide
C2736060|T201|LN|57647-0|LNC|C-peptide|C-peptide
C2736060|T201|OSN|57647-0|LNC|C-peptide|C-peptide
C2736060|T201|MTH_LN|57647-0|LNC|C-peptide|C-peptide
C2736060|T201|LC|57647-0|LNC|C-peptide|C-peptide
C2736060|T201|LN|57647-0|LNC|C peptide|C peptide
C2736060|T201|OSN|57647-0|LNC|C peptide|C peptide
C2736060|T201|MTH_LN|57647-0|LNC|C peptide|C peptide
C2736060|T201|LC|57647-0|LNC|C peptide|C peptide
C2736061|T201|LN|57651-2|LNC|C-peptide|C-peptide
C2736061|T201|OSN|57651-2|LNC|C-peptide|C-peptide
C2736061|T201|MTH_LN|57651-2|LNC|C-peptide|C-peptide
C2736061|T201|LC|57651-2|LNC|C-peptide|C-peptide
C2736061|T201|LN|57651-2|LNC|C peptide|C peptide
C2736061|T201|OSN|57651-2|LNC|C peptide|C peptide
C2736061|T201|MTH_LN|57651-2|LNC|C peptide|C peptide
C2736061|T201|LC|57651-2|LNC|C peptide|C peptide
C2736108|T201|LN|57698-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2736108|T201|OSN|57698-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2736108|T201|MTH_LN|57698-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2736108|T201|LC|57698-3|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C2736108|T201|LN|57698-3|LNC|LDL|LDL
C2736108|T201|OSN|57698-3|LNC|LDL|LDL
C2736108|T201|MTH_LN|57698-3|LNC|LDL|LDL
C2736108|T201|LC|57698-3|LNC|LDL|LDL
C2736108|T201|LN|57698-3|LNC|LDL cholesterol|LDL cholesterol
C2736108|T201|OSN|57698-3|LNC|LDL cholesterol|LDL cholesterol
C2736108|T201|MTH_LN|57698-3|LNC|LDL cholesterol|LDL cholesterol
C2736108|T201|LC|57698-3|LNC|LDL cholesterol|LDL cholesterol
C2736108|T201|LN|57698-3|LNC|low-density lipoprotein|low-density lipoprotein
C2736108|T201|OSN|57698-3|LNC|low-density lipoprotein|low-density lipoprotein
C2736108|T201|MTH_LN|57698-3|LNC|low-density lipoprotein|low-density lipoprotein
C2736108|T201|LC|57698-3|LNC|low-density lipoprotein|low-density lipoprotein
C2736108|T201|LN|57698-3|LNC|beta-lipoproteins|beta-lipoproteins
C2736108|T201|OSN|57698-3|LNC|beta-lipoproteins|beta-lipoproteins
C2736108|T201|MTH_LN|57698-3|LNC|beta-lipoproteins|beta-lipoproteins
C2736108|T201|LC|57698-3|LNC|beta-lipoproteins|beta-lipoproteins
C2736108|T201|LN|57698-3|LNC|LDL-C|LDL-C
C2736108|T201|OSN|57698-3|LNC|LDL-C|LDL-C
C2736108|T201|MTH_LN|57698-3|LNC|LDL-C|LDL-C
C2736108|T201|LC|57698-3|LNC|LDL-C|LDL-C
C2736136|T201|LN|57725-4|LNC|ACTH|ACTH
C2736136|T201|MTH_LN|57725-4|LNC|ACTH|ACTH
C2736136|T201|LC|57725-4|LNC|ACTH|ACTH
C2736136|T201|OSN|57725-4|LNC|ACTH|ACTH
C2736136|T201|LN|57725-4|LNC|corticotropin|corticotropin
C2736136|T201|MTH_LN|57725-4|LNC|corticotropin|corticotropin
C2736136|T201|LC|57725-4|LNC|corticotropin|corticotropin
C2736136|T201|OSN|57725-4|LNC|corticotropin|corticotropin
C2736136|T201|LN|57725-4|LNC|adrenocorticotropin|adrenocorticotropin
C2736136|T201|MTH_LN|57725-4|LNC|adrenocorticotropin|adrenocorticotropin
C2736136|T201|LC|57725-4|LNC|adrenocorticotropin|adrenocorticotropin
C2736136|T201|OSN|57725-4|LNC|adrenocorticotropin|adrenocorticotropin
C2736140|T201|LN|57728-8|LNC|lactate|lactate
C2736140|T201|MTH_LN|57728-8|LNC|lactate|lactate
C2736140|T201|LC|57728-8|LNC|lactate|lactate
C2736140|T201|OSN|57728-8|LNC|lactate|lactate
C2736141|T201|LN|57729-6|LNC|lactate|lactate
C2736141|T201|OSN|57729-6|LNC|lactate|lactate
C2736141|T201|MTH_LN|57729-6|LNC|lactate|lactate
C2736141|T201|LC|57729-6|LNC|lactate|lactate
C2736146|T201|LN|57735-3|LNC|Protein|Protein
C2736146|T201|MTH_LN|57735-3|LNC|Protein|Protein
C2736146|T201|OSN|57735-3|LNC|Protein|Protein
C2736146|T201|LC|57735-3|LNC|Protein|Protein
// C2736161|T201|LN|57747-8|LNC||
// C2736161|T201|LC|57747-8|LNC||
// C2736161|T201|MTH_LN|57747-8|LNC||
// C2736161|T201|OSN|57747-8|LNC||
C2736161|T201|LN|57747-8|LNC|occult|occult
C2736161|T201|LC|57747-8|LNC|occult|occult
C2736161|T201|MTH_LN|57747-8|LNC|occult|occult
C2736161|T201|OSN|57747-8|LNC|occult|occult
C2736165|T201|LN|57751-0|LNC|Hemoglobin|Hemoglobin
C2736165|T201|MTH_LN|57751-0|LNC|Hemoglobin|Hemoglobin
C2736165|T201|OSN|57751-0|LNC|Hemoglobin|Hemoglobin
C2736165|T201|LC|57751-0|LNC|Hemoglobin|Hemoglobin
C2736262|T201|LN|57838-5|LNC|Autoimmune antibody|Autoimmune antibody
C2736262|T201|OSN|57838-5|LNC|Autoimmune antibody|Autoimmune antibody
C2736262|T201|LC|57838-5|LNC|Autoimmune antibody|Autoimmune antibody
C2736262|T201|MTH_LN|57838-5|LNC|Autoimmune antibody|Autoimmune antibody
C2736320|T201|LN|57894-8|LNC|C-peptide|C-peptide
C2736320|T201|MTH_LN|57894-8|LNC|C-peptide|C-peptide
C2736320|T201|OSN|57894-8|LNC|C-peptide|C-peptide
C2736320|T201|LC|57894-8|LNC|C-peptide|C-peptide
C2736320|T201|LN|57894-8|LNC|C peptide|C peptide
C2736320|T201|MTH_LN|57894-8|LNC|C peptide|C peptide
C2736320|T201|OSN|57894-8|LNC|C peptide|C peptide
C2736320|T201|LC|57894-8|LNC|C peptide|C peptide
C2738971|T201|LN|57330-3|LNC|ACTH|ACTH
C2738971|T201|OSN|57330-3|LNC|ACTH|ACTH
C2738971|T201|MTH_LN|57330-3|LNC|ACTH|ACTH
C2738971|T201|LC|57330-3|LNC|ACTH|ACTH
C2738971|T201|LN|57330-3|LNC|corticotropin|corticotropin
C2738971|T201|OSN|57330-3|LNC|corticotropin|corticotropin
C2738971|T201|MTH_LN|57330-3|LNC|corticotropin|corticotropin
C2738971|T201|LC|57330-3|LNC|corticotropin|corticotropin
C2738971|T201|LN|57330-3|LNC|adrenocorticotropin|adrenocorticotropin
C2738971|T201|OSN|57330-3|LNC|adrenocorticotropin|adrenocorticotropin
C2738971|T201|MTH_LN|57330-3|LNC|adrenocorticotropin|adrenocorticotropin
C2738971|T201|LC|57330-3|LNC|adrenocorticotropin|adrenocorticotropin
C2738972|T201|LN|57332-9|LNC|urate|urate
C2738972|T201|OSN|57332-9|LNC|urate|urate
C2738972|T201|MTH_LN|57332-9|LNC|urate|urate
C2738972|T201|LC|57332-9|LNC|urate|urate
C2738972|T201|LN|57332-9|LNC|uric acid|uric acid
C2738972|T201|OSN|57332-9|LNC|uric acid|uric acid
C2738972|T201|MTH_LN|57332-9|LNC|uric acid|uric acid
C2738972|T201|LC|57332-9|LNC|uric acid|uric acid
C2923139|T201|LN|58805-3|LNC|neutrophil count|neutrophil count
C2923139|T201|MTH_LN|58805-3|LNC|neutrophil count|neutrophil count
C2923139|T201|LC|58805-3|LNC|neutrophil count|neutrophil count
C2923139|T201|OSN|58805-3|LNC|neutrophil count|neutrophil count
C2923139|T201|LN|58805-3|LNC|cytology|cytology
C2923139|T201|MTH_LN|58805-3|LNC|cytology|cytology
C2923139|T201|LC|58805-3|LNC|cytology|cytology
C2923139|T201|OSN|58805-3|LNC|cytology|cytology
C2923208|T201|LN|58896-2|LNC|C-peptide|C-peptide
C2923208|T201|MTH_LN|58896-2|LNC|C-peptide|C-peptide
C2923208|T201|LC|58896-2|LNC|C-peptide|C-peptide
C2923208|T201|OSN|58896-2|LNC|C-peptide|C-peptide
C2923208|T201|LN|58896-2|LNC|C peptide|C peptide
C2923208|T201|MTH_LN|58896-2|LNC|C peptide|C peptide
C2923208|T201|LC|58896-2|LNC|C peptide|C peptide
C2923208|T201|OSN|58896-2|LNC|C peptide|C peptide
C2923267|T201|LN|58946-5|LNC|luteinizing|luteinizing
C2923267|T201|MTH_LN|58946-5|LNC|luteinizing|luteinizing
C2923267|T201|OSN|58946-5|LNC|luteinizing|luteinizing
C2923267|T201|LC|58946-5|LNC|luteinizing|luteinizing
C2923267|T201|LN|58946-5|LNC|LH|LH
C2923267|T201|MTH_LN|58946-5|LNC|LH|LH
C2923267|T201|OSN|58946-5|LNC|LH|LH
C2923267|T201|LC|58946-5|LNC|LH|LH
C2923267|T201|LN|58946-5|LNC|luteinising|luteinising
C2923267|T201|MTH_LN|58946-5|LNC|luteinising|luteinising
C2923267|T201|OSN|58946-5|LNC|luteinising|luteinising
C2923267|T201|LC|58946-5|LNC|luteinising|luteinising
C2923319|T201|LN|58990-3|LNC|urate|urate
C2923319|T201|LC|58990-3|LNC|urate|urate
C2923319|T201|OSN|58990-3|LNC|urate|urate
C2923319|T201|MTH_LN|58990-3|LNC|urate|urate
C2923319|T201|LN|58990-3|LNC|uric acid|uric acid
C2923319|T201|LC|58990-3|LNC|uric acid|uric acid
C2923319|T201|OSN|58990-3|LNC|uric acid|uric acid
C2923319|T201|MTH_LN|58990-3|LNC|uric acid|uric acid
C2923333|T201|LN|59004-2|LNC|lactate|lactate
C2923333|T201|OSN|59004-2|LNC|lactate|lactate
C2923333|T201|LC|59004-2|LNC|lactate|lactate
C2923333|T201|MTH_LN|59004-2|LNC|lactate|lactate
C2923334|T201|LN|59005-9|LNC|lactate|lactate
C2923334|T201|OSN|59005-9|LNC|lactate|lactate
C2923334|T201|MTH_LN|59005-9|LNC|lactate|lactate
C2923334|T201|LC|59005-9|LNC|lactate|lactate
C2923335|T201|LN|59006-7|LNC|lactate|lactate
C2923335|T201|LC|59006-7|LNC|lactate|lactate
C2923335|T201|MTH_LN|59006-7|LNC|lactate|lactate
C2923335|T201|OSN|59006-7|LNC|lactate|lactate
C2923336|T201|LN|59007-5|LNC|lactate|lactate
C2923336|T201|OSN|59007-5|LNC|lactate|lactate
C2923336|T201|LC|59007-5|LNC|lactate|lactate
C2923336|T201|MTH_LN|59007-5|LNC|lactate|lactate
C2923341|T201|LN|59011-7|LNC|lactate|lactate
C2923341|T201|OSN|59011-7|LNC|lactate|lactate
C2923341|T201|MTH_LN|59011-7|LNC|lactate|lactate
C2923341|T201|LC|59011-7|LNC|lactate|lactate
C2923342|T201|LN|59012-5|LNC|lactate|lactate
C2923342|T201|LC|59012-5|LNC|lactate|lactate
C2923342|T201|MTH_LN|59012-5|LNC|lactate|lactate
C2923342|T201|OSN|59012-5|LNC|lactate|lactate
C2923343|T201|LN|59013-3|LNC|lactate|lactate
C2923343|T201|LC|59013-3|LNC|lactate|lactate
C2923343|T201|OSN|59013-3|LNC|lactate|lactate
C2923343|T201|MTH_LN|59013-3|LNC|lactate|lactate
C2923353|T201|LN|59048-9|LNC|lactate|lactate
C2923353|T201|OSN|59048-9|LNC|lactate|lactate
C2923353|T201|MTH_LN|59048-9|LNC|lactate|lactate
C2923353|T201|LC|59048-9|LNC|lactate|lactate
C2923385|T201|LN|59069-5|LNC|Antinuclear antibody|Antinuclear antibody
C2923385|T201|MTH_LN|59069-5|LNC|Antinuclear antibody|Antinuclear antibody
C2923385|T201|LC|59069-5|LNC|Antinuclear antibody|Antinuclear antibody
C2923385|T201|OSN|59069-5|LNC|Antinuclear antibody|Antinuclear antibody
C2923805|T201|LN|59408-5|LNC|oxygen|oxygen
C2923805|T201|LC|59408-5|LNC|oxygen|oxygen
C2923805|T201|MTH_LN|59408-5|LNC|oxygen|oxygen
C2923805|T201|OSN|59408-5|LNC|oxygen|oxygen
C2923932|T201|LN|59645-2|LNC|xenobiotic|xenobiotic
C2923932|T201|MTH_LN|59645-2|LNC|xenobiotic|xenobiotic
C2923932|T201|OSN|59645-2|LNC|xenobiotic|xenobiotic
C2923932|T201|LC|59645-2|LNC|xenobiotic|xenobiotic
C2923933|T201|LN|59646-0|LNC|cotinine|cotinine
C2923933|T201|MTH_LN|59646-0|LNC|cotinine|cotinine
C2923933|T201|LC|59646-0|LNC|cotinine|cotinine
C2923933|T201|OSN|59646-0|LNC|cotinine|cotinine
C2924077|T201|LN|59829-2|LNC|neutrophil count|neutrophil count
C2924077|T201|LC|59829-2|LNC|neutrophil count|neutrophil count
C2924077|T201|OSN|59829-2|LNC|neutrophil count|neutrophil count
C2924077|T201|MTH_LN|59829-2|LNC|neutrophil count|neutrophil count
C2924077|T201|LN|59829-2|LNC|cytology|cytology
C2924077|T201|LC|59829-2|LNC|cytology|cytology
C2924077|T201|OSN|59829-2|LNC|cytology|cytology
C2924077|T201|MTH_LN|59829-2|LNC|cytology|cytology
C2925635|T201|LN|57366-7|LNC|lactate|lactate
C2925635|T201|OSN|57366-7|LNC|lactate|lactate
C2925635|T201|MTH_LN|57366-7|LNC|lactate|lactate
C2925635|T201|LC|57366-7|LNC|lactate|lactate
C2925655|T201|LN|58816-0|LNC|C-peptide|C-peptide
C2925655|T201|LC|58816-0|LNC|C-peptide|C-peptide
C2925655|T201|OSN|58816-0|LNC|C-peptide|C-peptide
C2925655|T201|MTH_LN|58816-0|LNC|C-peptide|C-peptide
C2925655|T201|LN|58816-0|LNC|C peptide|C peptide
C2925655|T201|LC|58816-0|LNC|C peptide|C peptide
C2925655|T201|OSN|58816-0|LNC|C peptide|C peptide
C2925655|T201|MTH_LN|58816-0|LNC|C peptide|C peptide
C2925954|T201|LN|58494-6|LNC|C-peptide|C-peptide
C2925954|T201|OSN|58494-6|LNC|C-peptide|C-peptide
C2925954|T201|MTH_LN|58494-6|LNC|C-peptide|C-peptide
C2925954|T201|LC|58494-6|LNC|C-peptide|C-peptide
C2925954|T201|LN|58494-6|LNC|C peptide|C peptide
C2925954|T201|OSN|58494-6|LNC|C peptide|C peptide
C2925954|T201|MTH_LN|58494-6|LNC|C peptide|C peptide
C2925954|T201|LC|58494-6|LNC|C peptide|C peptide
C2925955|T201|LN|58495-3|LNC|C-peptide|C-peptide
C2925955|T201|OSN|58495-3|LNC|C-peptide|C-peptide
C2925955|T201|LC|58495-3|LNC|C-peptide|C-peptide
C2925955|T201|MTH_LN|58495-3|LNC|C-peptide|C-peptide
C2925955|T201|LN|58495-3|LNC|C peptide|C peptide
C2925955|T201|OSN|58495-3|LNC|C peptide|C peptide
C2925955|T201|LC|58495-3|LNC|C peptide|C peptide
C2925955|T201|MTH_LN|58495-3|LNC|C peptide|C peptide
C2926016|T201|LN|59032-3|LNC|lactate|lactate
C2926016|T201|LC|59032-3|LNC|lactate|lactate
C2926016|T201|MTH_LN|59032-3|LNC|lactate|lactate
C2926016|T201|OSN|59032-3|LNC|lactate|lactate
C2926027|T201|LN|58540-6|LNC|ACTH|ACTH
C2926027|T201|MTH_LN|58540-6|LNC|ACTH|ACTH
C2926027|T201|OSN|58540-6|LNC|ACTH|ACTH
C2926027|T201|LC|58540-6|LNC|ACTH|ACTH
C2926027|T201|LN|58540-6|LNC|corticotropin|corticotropin
C2926027|T201|MTH_LN|58540-6|LNC|corticotropin|corticotropin
C2926027|T201|OSN|58540-6|LNC|corticotropin|corticotropin
C2926027|T201|LC|58540-6|LNC|corticotropin|corticotropin
C2926027|T201|LN|58540-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926027|T201|MTH_LN|58540-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926027|T201|OSN|58540-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926027|T201|LC|58540-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926028|T201|LN|58541-4|LNC|ACTH|ACTH
C2926028|T201|OSN|58541-4|LNC|ACTH|ACTH
C2926028|T201|LC|58541-4|LNC|ACTH|ACTH
C2926028|T201|MTH_LN|58541-4|LNC|ACTH|ACTH
C2926028|T201|LN|58541-4|LNC|corticotropin|corticotropin
C2926028|T201|OSN|58541-4|LNC|corticotropin|corticotropin
C2926028|T201|LC|58541-4|LNC|corticotropin|corticotropin
C2926028|T201|MTH_LN|58541-4|LNC|corticotropin|corticotropin
C2926028|T201|LN|58541-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926028|T201|OSN|58541-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926028|T201|LC|58541-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926028|T201|MTH_LN|58541-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926029|T201|LN|58542-2|LNC|ACTH|ACTH
C2926029|T201|OSN|58542-2|LNC|ACTH|ACTH
C2926029|T201|MTH_LN|58542-2|LNC|ACTH|ACTH
C2926029|T201|LC|58542-2|LNC|ACTH|ACTH
C2926029|T201|LN|58542-2|LNC|corticotropin|corticotropin
C2926029|T201|OSN|58542-2|LNC|corticotropin|corticotropin
C2926029|T201|MTH_LN|58542-2|LNC|corticotropin|corticotropin
C2926029|T201|LC|58542-2|LNC|corticotropin|corticotropin
C2926029|T201|LN|58542-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926029|T201|OSN|58542-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926029|T201|MTH_LN|58542-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926029|T201|LC|58542-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926030|T201|LN|58543-0|LNC|ACTH|ACTH
C2926030|T201|LC|58543-0|LNC|ACTH|ACTH
C2926030|T201|MTH_LN|58543-0|LNC|ACTH|ACTH
C2926030|T201|OSN|58543-0|LNC|ACTH|ACTH
C2926030|T201|LN|58543-0|LNC|corticotropin|corticotropin
C2926030|T201|LC|58543-0|LNC|corticotropin|corticotropin
C2926030|T201|MTH_LN|58543-0|LNC|corticotropin|corticotropin
C2926030|T201|OSN|58543-0|LNC|corticotropin|corticotropin
C2926030|T201|LN|58543-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926030|T201|LC|58543-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926030|T201|MTH_LN|58543-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926030|T201|OSN|58543-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926031|T201|LN|58544-8|LNC|ACTH|ACTH
C2926031|T201|LC|58544-8|LNC|ACTH|ACTH
C2926031|T201|OSN|58544-8|LNC|ACTH|ACTH
C2926031|T201|MTH_LN|58544-8|LNC|ACTH|ACTH
C2926031|T201|LN|58544-8|LNC|corticotropin|corticotropin
C2926031|T201|LC|58544-8|LNC|corticotropin|corticotropin
C2926031|T201|OSN|58544-8|LNC|corticotropin|corticotropin
C2926031|T201|MTH_LN|58544-8|LNC|corticotropin|corticotropin
C2926031|T201|LN|58544-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926031|T201|LC|58544-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926031|T201|OSN|58544-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926031|T201|MTH_LN|58544-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926032|T201|LN|58545-5|LNC|ACTH|ACTH
C2926032|T201|LC|58545-5|LNC|ACTH|ACTH
C2926032|T201|OSN|58545-5|LNC|ACTH|ACTH
C2926032|T201|MTH_LN|58545-5|LNC|ACTH|ACTH
C2926032|T201|LN|58545-5|LNC|corticotropin|corticotropin
C2926032|T201|LC|58545-5|LNC|corticotropin|corticotropin
C2926032|T201|OSN|58545-5|LNC|corticotropin|corticotropin
C2926032|T201|MTH_LN|58545-5|LNC|corticotropin|corticotropin
C2926032|T201|LN|58545-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926032|T201|LC|58545-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926032|T201|OSN|58545-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926032|T201|MTH_LN|58545-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926033|T201|LN|58546-3|LNC|ACTH|ACTH
C2926033|T201|MTH_LN|58546-3|LNC|ACTH|ACTH
C2926033|T201|OSN|58546-3|LNC|ACTH|ACTH
C2926033|T201|LC|58546-3|LNC|ACTH|ACTH
C2926033|T201|LN|58546-3|LNC|corticotropin|corticotropin
C2926033|T201|MTH_LN|58546-3|LNC|corticotropin|corticotropin
C2926033|T201|OSN|58546-3|LNC|corticotropin|corticotropin
C2926033|T201|LC|58546-3|LNC|corticotropin|corticotropin
C2926033|T201|LN|58546-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926033|T201|MTH_LN|58546-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926033|T201|OSN|58546-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926033|T201|LC|58546-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926035|T201|LN|58686-7|LNC|C-peptide|C-peptide
C2926035|T201|LC|58686-7|LNC|C-peptide|C-peptide
C2926035|T201|OSN|58686-7|LNC|C-peptide|C-peptide
C2926035|T201|MTH_LN|58686-7|LNC|C-peptide|C-peptide
C2926035|T201|LN|58686-7|LNC|C peptide|C peptide
C2926035|T201|LC|58686-7|LNC|C peptide|C peptide
C2926035|T201|OSN|58686-7|LNC|C peptide|C peptide
C2926035|T201|MTH_LN|58686-7|LNC|C peptide|C peptide
C2926036|T201|LN|58687-5|LNC|ACTH|ACTH
C2926036|T201|MTH_LN|58687-5|LNC|ACTH|ACTH
C2926036|T201|OSN|58687-5|LNC|ACTH|ACTH
C2926036|T201|LC|58687-5|LNC|ACTH|ACTH
C2926036|T201|LN|58687-5|LNC|corticotropin|corticotropin
C2926036|T201|MTH_LN|58687-5|LNC|corticotropin|corticotropin
C2926036|T201|OSN|58687-5|LNC|corticotropin|corticotropin
C2926036|T201|LC|58687-5|LNC|corticotropin|corticotropin
C2926036|T201|LN|58687-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926036|T201|MTH_LN|58687-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926036|T201|OSN|58687-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926036|T201|LC|58687-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926049|T201|LN|58841-8|LNC|C-peptide|C-peptide
C2926049|T201|OSN|58841-8|LNC|C-peptide|C-peptide
C2926049|T201|LC|58841-8|LNC|C-peptide|C-peptide
C2926049|T201|MTH_LN|58841-8|LNC|C-peptide|C-peptide
C2926049|T201|LN|58841-8|LNC|C peptide|C peptide
C2926049|T201|OSN|58841-8|LNC|C peptide|C peptide
C2926049|T201|LC|58841-8|LNC|C peptide|C peptide
C2926049|T201|MTH_LN|58841-8|LNC|C peptide|C peptide
C2926219|T201|LN|58448-2|LNC|albumin|albumin
C2926219|T201|MTH_LN|58448-2|LNC|albumin|albumin
C2926219|T201|LC|58448-2|LNC|albumin|albumin
C2926219|T201|OSN|58448-2|LNC|albumin|albumin
C2926245|T201|LN|58496-1|LNC|C-peptide|C-peptide
C2926245|T201|LC|58496-1|LNC|C-peptide|C-peptide
C2926245|T201|OSN|58496-1|LNC|C-peptide|C-peptide
C2926245|T201|MTH_LN|58496-1|LNC|C-peptide|C-peptide
C2926245|T201|LN|58496-1|LNC|C peptide|C peptide
C2926245|T201|LC|58496-1|LNC|C peptide|C peptide
C2926245|T201|OSN|58496-1|LNC|C peptide|C peptide
C2926245|T201|MTH_LN|58496-1|LNC|C peptide|C peptide
C2926246|T201|LN|58497-9|LNC|C-peptide|C-peptide
C2926246|T201|MTH_LN|58497-9|LNC|C-peptide|C-peptide
C2926246|T201|LC|58497-9|LNC|C-peptide|C-peptide
C2926246|T201|OSN|58497-9|LNC|C-peptide|C-peptide
C2926246|T201|LN|58497-9|LNC|C peptide|C peptide
C2926246|T201|MTH_LN|58497-9|LNC|C peptide|C peptide
C2926246|T201|LC|58497-9|LNC|C peptide|C peptide
C2926246|T201|OSN|58497-9|LNC|C peptide|C peptide
C2926247|T201|LN|58498-7|LNC|C-peptide|C-peptide
C2926247|T201|LC|58498-7|LNC|C-peptide|C-peptide
C2926247|T201|OSN|58498-7|LNC|C-peptide|C-peptide
C2926247|T201|MTH_LN|58498-7|LNC|C-peptide|C-peptide
C2926247|T201|LN|58498-7|LNC|C peptide|C peptide
C2926247|T201|LC|58498-7|LNC|C peptide|C peptide
C2926247|T201|OSN|58498-7|LNC|C peptide|C peptide
C2926247|T201|MTH_LN|58498-7|LNC|C peptide|C peptide
C2926248|T201|LN|58499-5|LNC|C-peptide|C-peptide
C2926248|T201|OSN|58499-5|LNC|C-peptide|C-peptide
C2926248|T201|LC|58499-5|LNC|C-peptide|C-peptide
C2926248|T201|MTH_LN|58499-5|LNC|C-peptide|C-peptide
C2926248|T201|LN|58499-5|LNC|C peptide|C peptide
C2926248|T201|OSN|58499-5|LNC|C peptide|C peptide
C2926248|T201|LC|58499-5|LNC|C peptide|C peptide
C2926248|T201|MTH_LN|58499-5|LNC|C peptide|C peptide
C2926249|T201|LN|58500-0|LNC|C-peptide|C-peptide
C2926249|T201|OSN|58500-0|LNC|C-peptide|C-peptide
C2926249|T201|MTH_LN|58500-0|LNC|C-peptide|C-peptide
C2926249|T201|LC|58500-0|LNC|C-peptide|C-peptide
C2926249|T201|LN|58500-0|LNC|C peptide|C peptide
C2926249|T201|OSN|58500-0|LNC|C peptide|C peptide
C2926249|T201|MTH_LN|58500-0|LNC|C peptide|C peptide
C2926249|T201|LC|58500-0|LNC|C peptide|C peptide
C2926250|T201|LN|58501-8|LNC|C-peptide|C-peptide
C2926250|T201|MTH_LN|58501-8|LNC|C-peptide|C-peptide
C2926250|T201|OSN|58501-8|LNC|C-peptide|C-peptide
C2926250|T201|LC|58501-8|LNC|C-peptide|C-peptide
C2926250|T201|LN|58501-8|LNC|C peptide|C peptide
C2926250|T201|MTH_LN|58501-8|LNC|C peptide|C peptide
C2926250|T201|OSN|58501-8|LNC|C peptide|C peptide
C2926250|T201|LC|58501-8|LNC|C peptide|C peptide
C2926251|T201|LN|58502-6|LNC|C-peptide|C-peptide
C2926251|T201|LC|58502-6|LNC|C-peptide|C-peptide
C2926251|T201|OSN|58502-6|LNC|C-peptide|C-peptide
C2926251|T201|MTH_LN|58502-6|LNC|C-peptide|C-peptide
C2926251|T201|LN|58502-6|LNC|C peptide|C peptide
C2926251|T201|LC|58502-6|LNC|C peptide|C peptide
C2926251|T201|OSN|58502-6|LNC|C peptide|C peptide
C2926251|T201|MTH_LN|58502-6|LNC|C peptide|C peptide
C2926252|T201|LN|58503-4|LNC|C-peptide|C-peptide
C2926252|T201|MTH_LN|58503-4|LNC|C-peptide|C-peptide
C2926252|T201|LC|58503-4|LNC|C-peptide|C-peptide
C2926252|T201|OSN|58503-4|LNC|C-peptide|C-peptide
C2926252|T201|LN|58503-4|LNC|C peptide|C peptide
C2926252|T201|MTH_LN|58503-4|LNC|C peptide|C peptide
C2926252|T201|LC|58503-4|LNC|C peptide|C peptide
C2926252|T201|OSN|58503-4|LNC|C peptide|C peptide
C2926253|T201|LN|58504-2|LNC|C-peptide|C-peptide
C2926253|T201|LC|58504-2|LNC|C-peptide|C-peptide
C2926253|T201|MTH_LN|58504-2|LNC|C-peptide|C-peptide
C2926253|T201|OSN|58504-2|LNC|C-peptide|C-peptide
C2926253|T201|LN|58504-2|LNC|C peptide|C peptide
C2926253|T201|LC|58504-2|LNC|C peptide|C peptide
C2926253|T201|MTH_LN|58504-2|LNC|C peptide|C peptide
C2926253|T201|OSN|58504-2|LNC|C peptide|C peptide
C2926254|T201|LN|58505-9|LNC|C-peptide|C-peptide
C2926254|T201|OSN|58505-9|LNC|C-peptide|C-peptide
C2926254|T201|LC|58505-9|LNC|C-peptide|C-peptide
C2926254|T201|MTH_LN|58505-9|LNC|C-peptide|C-peptide
C2926254|T201|LN|58505-9|LNC|C peptide|C peptide
C2926254|T201|OSN|58505-9|LNC|C peptide|C peptide
C2926254|T201|LC|58505-9|LNC|C peptide|C peptide
C2926254|T201|MTH_LN|58505-9|LNC|C peptide|C peptide
C2926255|T201|LN|58506-7|LNC|C-peptide|C-peptide
C2926255|T201|LC|58506-7|LNC|C-peptide|C-peptide
C2926255|T201|OSN|58506-7|LNC|C-peptide|C-peptide
C2926255|T201|MTH_LN|58506-7|LNC|C-peptide|C-peptide
C2926255|T201|LN|58506-7|LNC|C peptide|C peptide
C2926255|T201|LC|58506-7|LNC|C peptide|C peptide
C2926255|T201|OSN|58506-7|LNC|C peptide|C peptide
C2926255|T201|MTH_LN|58506-7|LNC|C peptide|C peptide
C2926256|T201|LN|58507-5|LNC|C-peptide|C-peptide
C2926256|T201|OSN|58507-5|LNC|C-peptide|C-peptide
C2926256|T201|MTH_LN|58507-5|LNC|C-peptide|C-peptide
C2926256|T201|LC|58507-5|LNC|C-peptide|C-peptide
C2926256|T201|LN|58507-5|LNC|C peptide|C peptide
C2926256|T201|OSN|58507-5|LNC|C peptide|C peptide
C2926256|T201|MTH_LN|58507-5|LNC|C peptide|C peptide
C2926256|T201|LC|58507-5|LNC|C peptide|C peptide
C2926257|T201|LN|58508-3|LNC|C-peptide|C-peptide
C2926257|T201|LC|58508-3|LNC|C-peptide|C-peptide
C2926257|T201|OSN|58508-3|LNC|C-peptide|C-peptide
C2926257|T201|MTH_LN|58508-3|LNC|C-peptide|C-peptide
C2926257|T201|LN|58508-3|LNC|C peptide|C peptide
C2926257|T201|LC|58508-3|LNC|C peptide|C peptide
C2926257|T201|OSN|58508-3|LNC|C peptide|C peptide
C2926257|T201|MTH_LN|58508-3|LNC|C peptide|C peptide
C2926258|T201|LN|58509-1|LNC|C-peptide|C-peptide
C2926258|T201|LC|58509-1|LNC|C-peptide|C-peptide
C2926258|T201|MTH_LN|58509-1|LNC|C-peptide|C-peptide
C2926258|T201|OSN|58509-1|LNC|C-peptide|C-peptide
C2926258|T201|LN|58509-1|LNC|C peptide|C peptide
C2926258|T201|LC|58509-1|LNC|C peptide|C peptide
C2926258|T201|MTH_LN|58509-1|LNC|C peptide|C peptide
C2926258|T201|OSN|58509-1|LNC|C peptide|C peptide
C2926259|T201|LN|58510-9|LNC|C-peptide|C-peptide
C2926259|T201|LC|58510-9|LNC|C-peptide|C-peptide
C2926259|T201|MTH_LN|58510-9|LNC|C-peptide|C-peptide
C2926259|T201|OSN|58510-9|LNC|C-peptide|C-peptide
C2926259|T201|LN|58510-9|LNC|C peptide|C peptide
C2926259|T201|LC|58510-9|LNC|C peptide|C peptide
C2926259|T201|MTH_LN|58510-9|LNC|C peptide|C peptide
C2926259|T201|OSN|58510-9|LNC|C peptide|C peptide
C2926260|T201|LN|58511-7|LNC|C-peptide|C-peptide
C2926260|T201|OSN|58511-7|LNC|C-peptide|C-peptide
C2926260|T201|LC|58511-7|LNC|C-peptide|C-peptide
C2926260|T201|MTH_LN|58511-7|LNC|C-peptide|C-peptide
C2926260|T201|LN|58511-7|LNC|C peptide|C peptide
C2926260|T201|OSN|58511-7|LNC|C peptide|C peptide
C2926260|T201|LC|58511-7|LNC|C peptide|C peptide
C2926260|T201|MTH_LN|58511-7|LNC|C peptide|C peptide
C2926261|T201|LN|58512-5|LNC|C-peptide|C-peptide
C2926261|T201|MTH_LN|58512-5|LNC|C-peptide|C-peptide
C2926261|T201|OSN|58512-5|LNC|C-peptide|C-peptide
C2926261|T201|LC|58512-5|LNC|C-peptide|C-peptide
C2926261|T201|LN|58512-5|LNC|C peptide|C peptide
C2926261|T201|MTH_LN|58512-5|LNC|C peptide|C peptide
C2926261|T201|OSN|58512-5|LNC|C peptide|C peptide
C2926261|T201|LC|58512-5|LNC|C peptide|C peptide
C2926262|T201|LN|58513-3|LNC|C-peptide|C-peptide
C2926262|T201|MTH_LN|58513-3|LNC|C-peptide|C-peptide
C2926262|T201|OSN|58513-3|LNC|C-peptide|C-peptide
C2926262|T201|LC|58513-3|LNC|C-peptide|C-peptide
C2926262|T201|LN|58513-3|LNC|C peptide|C peptide
C2926262|T201|MTH_LN|58513-3|LNC|C peptide|C peptide
C2926262|T201|OSN|58513-3|LNC|C peptide|C peptide
C2926262|T201|LC|58513-3|LNC|C peptide|C peptide
C2926263|T201|LN|58514-1|LNC|C-peptide|C-peptide
C2926263|T201|MTH_LN|58514-1|LNC|C-peptide|C-peptide
C2926263|T201|OSN|58514-1|LNC|C-peptide|C-peptide
C2926263|T201|LC|58514-1|LNC|C-peptide|C-peptide
C2926263|T201|LN|58514-1|LNC|C peptide|C peptide
C2926263|T201|MTH_LN|58514-1|LNC|C peptide|C peptide
C2926263|T201|OSN|58514-1|LNC|C peptide|C peptide
C2926263|T201|LC|58514-1|LNC|C peptide|C peptide
C2926264|T201|LN|58515-8|LNC|C-peptide|C-peptide
C2926264|T201|OSN|58515-8|LNC|C-peptide|C-peptide
C2926264|T201|MTH_LN|58515-8|LNC|C-peptide|C-peptide
C2926264|T201|LC|58515-8|LNC|C-peptide|C-peptide
C2926264|T201|LN|58515-8|LNC|C peptide|C peptide
C2926264|T201|OSN|58515-8|LNC|C peptide|C peptide
C2926264|T201|MTH_LN|58515-8|LNC|C peptide|C peptide
C2926264|T201|LC|58515-8|LNC|C peptide|C peptide
C2926265|T201|LN|58516-6|LNC|C-peptide|C-peptide
C2926265|T201|MTH_LN|58516-6|LNC|C-peptide|C-peptide
C2926265|T201|OSN|58516-6|LNC|C-peptide|C-peptide
C2926265|T201|LC|58516-6|LNC|C-peptide|C-peptide
C2926265|T201|LN|58516-6|LNC|C peptide|C peptide
C2926265|T201|MTH_LN|58516-6|LNC|C peptide|C peptide
C2926265|T201|OSN|58516-6|LNC|C peptide|C peptide
C2926265|T201|LC|58516-6|LNC|C peptide|C peptide
C2926266|T201|LN|58517-4|LNC|C-peptide|C-peptide
C2926266|T201|LC|58517-4|LNC|C-peptide|C-peptide
C2926266|T201|OSN|58517-4|LNC|C-peptide|C-peptide
C2926266|T201|MTH_LN|58517-4|LNC|C-peptide|C-peptide
C2926266|T201|LN|58517-4|LNC|C peptide|C peptide
C2926266|T201|LC|58517-4|LNC|C peptide|C peptide
C2926266|T201|OSN|58517-4|LNC|C peptide|C peptide
C2926266|T201|MTH_LN|58517-4|LNC|C peptide|C peptide
C2926267|T201|LN|58518-2|LNC|C-peptide|C-peptide
C2926267|T201|OSN|58518-2|LNC|C-peptide|C-peptide
C2926267|T201|MTH_LN|58518-2|LNC|C-peptide|C-peptide
C2926267|T201|LC|58518-2|LNC|C-peptide|C-peptide
C2926267|T201|LN|58518-2|LNC|C peptide|C peptide
C2926267|T201|OSN|58518-2|LNC|C peptide|C peptide
C2926267|T201|MTH_LN|58518-2|LNC|C peptide|C peptide
C2926267|T201|LC|58518-2|LNC|C peptide|C peptide
C2926268|T201|LN|58519-0|LNC|C-peptide|C-peptide
C2926268|T201|LC|58519-0|LNC|C-peptide|C-peptide
C2926268|T201|OSN|58519-0|LNC|C-peptide|C-peptide
C2926268|T201|MTH_LN|58519-0|LNC|C-peptide|C-peptide
C2926268|T201|LN|58519-0|LNC|C peptide|C peptide
C2926268|T201|LC|58519-0|LNC|C peptide|C peptide
C2926268|T201|OSN|58519-0|LNC|C peptide|C peptide
C2926268|T201|MTH_LN|58519-0|LNC|C peptide|C peptide
C2926269|T201|LN|58520-8|LNC|C-peptide|C-peptide
C2926269|T201|LC|58520-8|LNC|C-peptide|C-peptide
C2926269|T201|OSN|58520-8|LNC|C-peptide|C-peptide
C2926269|T201|MTH_LN|58520-8|LNC|C-peptide|C-peptide
C2926269|T201|LN|58520-8|LNC|C peptide|C peptide
C2926269|T201|LC|58520-8|LNC|C peptide|C peptide
C2926269|T201|OSN|58520-8|LNC|C peptide|C peptide
C2926269|T201|MTH_LN|58520-8|LNC|C peptide|C peptide
C2926270|T201|LN|58521-6|LNC|C-peptide|C-peptide
C2926270|T201|LC|58521-6|LNC|C-peptide|C-peptide
C2926270|T201|MTH_LN|58521-6|LNC|C-peptide|C-peptide
C2926270|T201|OSN|58521-6|LNC|C-peptide|C-peptide
C2926270|T201|LN|58521-6|LNC|C peptide|C peptide
C2926270|T201|LC|58521-6|LNC|C peptide|C peptide
C2926270|T201|MTH_LN|58521-6|LNC|C peptide|C peptide
C2926270|T201|OSN|58521-6|LNC|C peptide|C peptide
C2926271|T201|LN|58522-4|LNC|C-peptide|C-peptide
C2926271|T201|OSN|58522-4|LNC|C-peptide|C-peptide
C2926271|T201|LC|58522-4|LNC|C-peptide|C-peptide
C2926271|T201|MTH_LN|58522-4|LNC|C-peptide|C-peptide
C2926271|T201|LN|58522-4|LNC|C peptide|C peptide
C2926271|T201|OSN|58522-4|LNC|C peptide|C peptide
C2926271|T201|LC|58522-4|LNC|C peptide|C peptide
C2926271|T201|MTH_LN|58522-4|LNC|C peptide|C peptide
C2926272|T201|LN|58523-2|LNC|ACTH|ACTH
C2926272|T201|LC|58523-2|LNC|ACTH|ACTH
C2926272|T201|MTH_LN|58523-2|LNC|ACTH|ACTH
C2926272|T201|OSN|58523-2|LNC|ACTH|ACTH
C2926272|T201|LN|58523-2|LNC|corticotropin|corticotropin
C2926272|T201|LC|58523-2|LNC|corticotropin|corticotropin
C2926272|T201|MTH_LN|58523-2|LNC|corticotropin|corticotropin
C2926272|T201|OSN|58523-2|LNC|corticotropin|corticotropin
C2926272|T201|LN|58523-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926272|T201|LC|58523-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926272|T201|MTH_LN|58523-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926272|T201|OSN|58523-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926273|T201|LN|58524-0|LNC|ACTH|ACTH
C2926273|T201|MTH_LN|58524-0|LNC|ACTH|ACTH
C2926273|T201|LC|58524-0|LNC|ACTH|ACTH
C2926273|T201|OSN|58524-0|LNC|ACTH|ACTH
C2926273|T201|LN|58524-0|LNC|corticotropin|corticotropin
C2926273|T201|MTH_LN|58524-0|LNC|corticotropin|corticotropin
C2926273|T201|LC|58524-0|LNC|corticotropin|corticotropin
C2926273|T201|OSN|58524-0|LNC|corticotropin|corticotropin
C2926273|T201|LN|58524-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926273|T201|MTH_LN|58524-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926273|T201|LC|58524-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926273|T201|OSN|58524-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926274|T201|LN|58525-7|LNC|ACTH|ACTH
C2926274|T201|LC|58525-7|LNC|ACTH|ACTH
C2926274|T201|MTH_LN|58525-7|LNC|ACTH|ACTH
C2926274|T201|OSN|58525-7|LNC|ACTH|ACTH
C2926274|T201|LN|58525-7|LNC|corticotropin|corticotropin
C2926274|T201|LC|58525-7|LNC|corticotropin|corticotropin
C2926274|T201|MTH_LN|58525-7|LNC|corticotropin|corticotropin
C2926274|T201|OSN|58525-7|LNC|corticotropin|corticotropin
C2926274|T201|LN|58525-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926274|T201|LC|58525-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926274|T201|MTH_LN|58525-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926274|T201|OSN|58525-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926275|T201|LN|58526-5|LNC|ACTH|ACTH
C2926275|T201|LC|58526-5|LNC|ACTH|ACTH
C2926275|T201|OSN|58526-5|LNC|ACTH|ACTH
C2926275|T201|MTH_LN|58526-5|LNC|ACTH|ACTH
C2926275|T201|LN|58526-5|LNC|corticotropin|corticotropin
C2926275|T201|LC|58526-5|LNC|corticotropin|corticotropin
C2926275|T201|OSN|58526-5|LNC|corticotropin|corticotropin
C2926275|T201|MTH_LN|58526-5|LNC|corticotropin|corticotropin
C2926275|T201|LN|58526-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926275|T201|LC|58526-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926275|T201|OSN|58526-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926275|T201|MTH_LN|58526-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926276|T201|LN|58527-3|LNC|ACTH|ACTH
C2926276|T201|OSN|58527-3|LNC|ACTH|ACTH
C2926276|T201|LC|58527-3|LNC|ACTH|ACTH
C2926276|T201|MTH_LN|58527-3|LNC|ACTH|ACTH
C2926276|T201|LN|58527-3|LNC|corticotropin|corticotropin
C2926276|T201|OSN|58527-3|LNC|corticotropin|corticotropin
C2926276|T201|LC|58527-3|LNC|corticotropin|corticotropin
C2926276|T201|MTH_LN|58527-3|LNC|corticotropin|corticotropin
C2926276|T201|LN|58527-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926276|T201|OSN|58527-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926276|T201|LC|58527-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926276|T201|MTH_LN|58527-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926277|T201|LN|58528-1|LNC|ACTH|ACTH
C2926277|T201|LC|58528-1|LNC|ACTH|ACTH
C2926277|T201|OSN|58528-1|LNC|ACTH|ACTH
C2926277|T201|MTH_LN|58528-1|LNC|ACTH|ACTH
C2926277|T201|LN|58528-1|LNC|corticotropin|corticotropin
C2926277|T201|LC|58528-1|LNC|corticotropin|corticotropin
C2926277|T201|OSN|58528-1|LNC|corticotropin|corticotropin
C2926277|T201|MTH_LN|58528-1|LNC|corticotropin|corticotropin
C2926277|T201|LN|58528-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926277|T201|LC|58528-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926277|T201|OSN|58528-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926277|T201|MTH_LN|58528-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926278|T201|LN|58529-9|LNC|ACTH|ACTH
C2926278|T201|OSN|58529-9|LNC|ACTH|ACTH
C2926278|T201|MTH_LN|58529-9|LNC|ACTH|ACTH
C2926278|T201|LC|58529-9|LNC|ACTH|ACTH
C2926278|T201|LN|58529-9|LNC|corticotropin|corticotropin
C2926278|T201|OSN|58529-9|LNC|corticotropin|corticotropin
C2926278|T201|MTH_LN|58529-9|LNC|corticotropin|corticotropin
C2926278|T201|LC|58529-9|LNC|corticotropin|corticotropin
C2926278|T201|LN|58529-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926278|T201|OSN|58529-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926278|T201|MTH_LN|58529-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926278|T201|LC|58529-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926279|T201|LN|58530-7|LNC|ACTH|ACTH
C2926279|T201|LC|58530-7|LNC|ACTH|ACTH
C2926279|T201|OSN|58530-7|LNC|ACTH|ACTH
C2926279|T201|MTH_LN|58530-7|LNC|ACTH|ACTH
C2926279|T201|LN|58530-7|LNC|corticotropin|corticotropin
C2926279|T201|LC|58530-7|LNC|corticotropin|corticotropin
C2926279|T201|OSN|58530-7|LNC|corticotropin|corticotropin
C2926279|T201|MTH_LN|58530-7|LNC|corticotropin|corticotropin
C2926279|T201|LN|58530-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926279|T201|LC|58530-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926279|T201|OSN|58530-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926279|T201|MTH_LN|58530-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926280|T201|LN|58531-5|LNC|ACTH|ACTH
C2926280|T201|OSN|58531-5|LNC|ACTH|ACTH
C2926280|T201|LC|58531-5|LNC|ACTH|ACTH
C2926280|T201|MTH_LN|58531-5|LNC|ACTH|ACTH
C2926280|T201|LN|58531-5|LNC|corticotropin|corticotropin
C2926280|T201|OSN|58531-5|LNC|corticotropin|corticotropin
C2926280|T201|LC|58531-5|LNC|corticotropin|corticotropin
C2926280|T201|MTH_LN|58531-5|LNC|corticotropin|corticotropin
C2926280|T201|LN|58531-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926280|T201|OSN|58531-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926280|T201|LC|58531-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926280|T201|MTH_LN|58531-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926281|T201|LN|58532-3|LNC|ACTH|ACTH
C2926281|T201|OSN|58532-3|LNC|ACTH|ACTH
C2926281|T201|LC|58532-3|LNC|ACTH|ACTH
C2926281|T201|MTH_LN|58532-3|LNC|ACTH|ACTH
C2926281|T201|LN|58532-3|LNC|corticotropin|corticotropin
C2926281|T201|OSN|58532-3|LNC|corticotropin|corticotropin
C2926281|T201|LC|58532-3|LNC|corticotropin|corticotropin
C2926281|T201|MTH_LN|58532-3|LNC|corticotropin|corticotropin
C2926281|T201|LN|58532-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926281|T201|OSN|58532-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926281|T201|LC|58532-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926281|T201|MTH_LN|58532-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926282|T201|LN|58533-1|LNC|ACTH|ACTH
C2926282|T201|OSN|58533-1|LNC|ACTH|ACTH
C2926282|T201|LC|58533-1|LNC|ACTH|ACTH
C2926282|T201|MTH_LN|58533-1|LNC|ACTH|ACTH
C2926282|T201|LN|58533-1|LNC|corticotropin|corticotropin
C2926282|T201|OSN|58533-1|LNC|corticotropin|corticotropin
C2926282|T201|LC|58533-1|LNC|corticotropin|corticotropin
C2926282|T201|MTH_LN|58533-1|LNC|corticotropin|corticotropin
C2926282|T201|LN|58533-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926282|T201|OSN|58533-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926282|T201|LC|58533-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926282|T201|MTH_LN|58533-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926283|T201|LN|58534-9|LNC|ACTH|ACTH
C2926283|T201|MTH_LN|58534-9|LNC|ACTH|ACTH
C2926283|T201|OSN|58534-9|LNC|ACTH|ACTH
C2926283|T201|LC|58534-9|LNC|ACTH|ACTH
C2926283|T201|LN|58534-9|LNC|corticotropin|corticotropin
C2926283|T201|MTH_LN|58534-9|LNC|corticotropin|corticotropin
C2926283|T201|OSN|58534-9|LNC|corticotropin|corticotropin
C2926283|T201|LC|58534-9|LNC|corticotropin|corticotropin
C2926283|T201|LN|58534-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926283|T201|MTH_LN|58534-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926283|T201|OSN|58534-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926283|T201|LC|58534-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926284|T201|LN|58535-6|LNC|ACTH|ACTH
C2926284|T201|OSN|58535-6|LNC|ACTH|ACTH
C2926284|T201|LC|58535-6|LNC|ACTH|ACTH
C2926284|T201|MTH_LN|58535-6|LNC|ACTH|ACTH
C2926284|T201|LN|58535-6|LNC|corticotropin|corticotropin
C2926284|T201|OSN|58535-6|LNC|corticotropin|corticotropin
C2926284|T201|LC|58535-6|LNC|corticotropin|corticotropin
C2926284|T201|MTH_LN|58535-6|LNC|corticotropin|corticotropin
C2926284|T201|LN|58535-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926284|T201|OSN|58535-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926284|T201|LC|58535-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926284|T201|MTH_LN|58535-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926285|T201|LN|58536-4|LNC|ACTH|ACTH
C2926285|T201|OSN|58536-4|LNC|ACTH|ACTH
C2926285|T201|LC|58536-4|LNC|ACTH|ACTH
C2926285|T201|MTH_LN|58536-4|LNC|ACTH|ACTH
C2926285|T201|LN|58536-4|LNC|corticotropin|corticotropin
C2926285|T201|OSN|58536-4|LNC|corticotropin|corticotropin
C2926285|T201|LC|58536-4|LNC|corticotropin|corticotropin
C2926285|T201|MTH_LN|58536-4|LNC|corticotropin|corticotropin
C2926285|T201|LN|58536-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926285|T201|OSN|58536-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926285|T201|LC|58536-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926285|T201|MTH_LN|58536-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926286|T201|LN|58537-2|LNC|ACTH|ACTH
C2926286|T201|MTH_LN|58537-2|LNC|ACTH|ACTH
C2926286|T201|OSN|58537-2|LNC|ACTH|ACTH
C2926286|T201|LC|58537-2|LNC|ACTH|ACTH
C2926286|T201|LN|58537-2|LNC|corticotropin|corticotropin
C2926286|T201|MTH_LN|58537-2|LNC|corticotropin|corticotropin
C2926286|T201|OSN|58537-2|LNC|corticotropin|corticotropin
C2926286|T201|LC|58537-2|LNC|corticotropin|corticotropin
C2926286|T201|LN|58537-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926286|T201|MTH_LN|58537-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926286|T201|OSN|58537-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926286|T201|LC|58537-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926287|T201|LN|58538-0|LNC|ACTH|ACTH
C2926287|T201|MTH_LN|58538-0|LNC|ACTH|ACTH
C2926287|T201|LC|58538-0|LNC|ACTH|ACTH
C2926287|T201|OSN|58538-0|LNC|ACTH|ACTH
C2926287|T201|LN|58538-0|LNC|corticotropin|corticotropin
C2926287|T201|MTH_LN|58538-0|LNC|corticotropin|corticotropin
C2926287|T201|LC|58538-0|LNC|corticotropin|corticotropin
C2926287|T201|OSN|58538-0|LNC|corticotropin|corticotropin
C2926287|T201|LN|58538-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926287|T201|MTH_LN|58538-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926287|T201|LC|58538-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926287|T201|OSN|58538-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926288|T201|LN|58539-8|LNC|ACTH|ACTH
C2926288|T201|LC|58539-8|LNC|ACTH|ACTH
C2926288|T201|OSN|58539-8|LNC|ACTH|ACTH
C2926288|T201|MTH_LN|58539-8|LNC|ACTH|ACTH
C2926288|T201|LN|58539-8|LNC|corticotropin|corticotropin
C2926288|T201|LC|58539-8|LNC|corticotropin|corticotropin
C2926288|T201|OSN|58539-8|LNC|corticotropin|corticotropin
C2926288|T201|MTH_LN|58539-8|LNC|corticotropin|corticotropin
C2926288|T201|LN|58539-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926288|T201|LC|58539-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926288|T201|OSN|58539-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926288|T201|MTH_LN|58539-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926289|T201|LN|58547-1|LNC|ACTH|ACTH
C2926289|T201|LC|58547-1|LNC|ACTH|ACTH
C2926289|T201|OSN|58547-1|LNC|ACTH|ACTH
C2926289|T201|MTH_LN|58547-1|LNC|ACTH|ACTH
C2926289|T201|LN|58547-1|LNC|corticotropin|corticotropin
C2926289|T201|LC|58547-1|LNC|corticotropin|corticotropin
C2926289|T201|OSN|58547-1|LNC|corticotropin|corticotropin
C2926289|T201|MTH_LN|58547-1|LNC|corticotropin|corticotropin
C2926289|T201|LN|58547-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926289|T201|LC|58547-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926289|T201|OSN|58547-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926289|T201|MTH_LN|58547-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926290|T201|LN|58548-9|LNC|ACTH|ACTH
C2926290|T201|LC|58548-9|LNC|ACTH|ACTH
C2926290|T201|OSN|58548-9|LNC|ACTH|ACTH
C2926290|T201|MTH_LN|58548-9|LNC|ACTH|ACTH
C2926290|T201|LN|58548-9|LNC|corticotropin|corticotropin
C2926290|T201|LC|58548-9|LNC|corticotropin|corticotropin
C2926290|T201|OSN|58548-9|LNC|corticotropin|corticotropin
C2926290|T201|MTH_LN|58548-9|LNC|corticotropin|corticotropin
C2926290|T201|LN|58548-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926290|T201|LC|58548-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926290|T201|OSN|58548-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926290|T201|MTH_LN|58548-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926291|T201|LN|58549-7|LNC|ACTH|ACTH
C2926291|T201|LC|58549-7|LNC|ACTH|ACTH
C2926291|T201|OSN|58549-7|LNC|ACTH|ACTH
C2926291|T201|MTH_LN|58549-7|LNC|ACTH|ACTH
C2926291|T201|LN|58549-7|LNC|corticotropin|corticotropin
C2926291|T201|LC|58549-7|LNC|corticotropin|corticotropin
C2926291|T201|OSN|58549-7|LNC|corticotropin|corticotropin
C2926291|T201|MTH_LN|58549-7|LNC|corticotropin|corticotropin
C2926291|T201|LN|58549-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926291|T201|LC|58549-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926291|T201|OSN|58549-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926291|T201|MTH_LN|58549-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926292|T201|LN|58550-5|LNC|ACTH|ACTH
C2926292|T201|OSN|58550-5|LNC|ACTH|ACTH
C2926292|T201|MTH_LN|58550-5|LNC|ACTH|ACTH
C2926292|T201|LC|58550-5|LNC|ACTH|ACTH
C2926292|T201|LN|58550-5|LNC|corticotropin|corticotropin
C2926292|T201|OSN|58550-5|LNC|corticotropin|corticotropin
C2926292|T201|MTH_LN|58550-5|LNC|corticotropin|corticotropin
C2926292|T201|LC|58550-5|LNC|corticotropin|corticotropin
C2926292|T201|LN|58550-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926292|T201|OSN|58550-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926292|T201|MTH_LN|58550-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926292|T201|LC|58550-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926293|T201|LN|58551-3|LNC|ACTH|ACTH
C2926293|T201|OSN|58551-3|LNC|ACTH|ACTH
C2926293|T201|LC|58551-3|LNC|ACTH|ACTH
C2926293|T201|MTH_LN|58551-3|LNC|ACTH|ACTH
C2926293|T201|LN|58551-3|LNC|corticotropin|corticotropin
C2926293|T201|OSN|58551-3|LNC|corticotropin|corticotropin
C2926293|T201|LC|58551-3|LNC|corticotropin|corticotropin
C2926293|T201|MTH_LN|58551-3|LNC|corticotropin|corticotropin
C2926293|T201|LN|58551-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926293|T201|OSN|58551-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926293|T201|LC|58551-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926293|T201|MTH_LN|58551-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926294|T201|LN|58552-1|LNC|ACTH|ACTH
C2926294|T201|OSN|58552-1|LNC|ACTH|ACTH
C2926294|T201|MTH_LN|58552-1|LNC|ACTH|ACTH
C2926294|T201|LC|58552-1|LNC|ACTH|ACTH
C2926294|T201|LN|58552-1|LNC|corticotropin|corticotropin
C2926294|T201|OSN|58552-1|LNC|corticotropin|corticotropin
C2926294|T201|MTH_LN|58552-1|LNC|corticotropin|corticotropin
C2926294|T201|LC|58552-1|LNC|corticotropin|corticotropin
C2926294|T201|LN|58552-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926294|T201|OSN|58552-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926294|T201|MTH_LN|58552-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926294|T201|LC|58552-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926295|T201|LN|58553-9|LNC|ACTH|ACTH
C2926295|T201|OSN|58553-9|LNC|ACTH|ACTH
C2926295|T201|LC|58553-9|LNC|ACTH|ACTH
C2926295|T201|MTH_LN|58553-9|LNC|ACTH|ACTH
C2926295|T201|LN|58553-9|LNC|corticotropin|corticotropin
C2926295|T201|OSN|58553-9|LNC|corticotropin|corticotropin
C2926295|T201|LC|58553-9|LNC|corticotropin|corticotropin
C2926295|T201|MTH_LN|58553-9|LNC|corticotropin|corticotropin
C2926295|T201|LN|58553-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926295|T201|OSN|58553-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926295|T201|LC|58553-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926295|T201|MTH_LN|58553-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926296|T201|LN|58554-7|LNC|ACTH|ACTH
C2926296|T201|LC|58554-7|LNC|ACTH|ACTH
C2926296|T201|OSN|58554-7|LNC|ACTH|ACTH
C2926296|T201|MTH_LN|58554-7|LNC|ACTH|ACTH
C2926296|T201|LN|58554-7|LNC|corticotropin|corticotropin
C2926296|T201|LC|58554-7|LNC|corticotropin|corticotropin
C2926296|T201|OSN|58554-7|LNC|corticotropin|corticotropin
C2926296|T201|MTH_LN|58554-7|LNC|corticotropin|corticotropin
C2926296|T201|LN|58554-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926296|T201|LC|58554-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926296|T201|OSN|58554-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926296|T201|MTH_LN|58554-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926297|T201|LN|58555-4|LNC|ACTH|ACTH
C2926297|T201|OSN|58555-4|LNC|ACTH|ACTH
C2926297|T201|MTH_LN|58555-4|LNC|ACTH|ACTH
C2926297|T201|LC|58555-4|LNC|ACTH|ACTH
C2926297|T201|LN|58555-4|LNC|corticotropin|corticotropin
C2926297|T201|OSN|58555-4|LNC|corticotropin|corticotropin
C2926297|T201|MTH_LN|58555-4|LNC|corticotropin|corticotropin
C2926297|T201|LC|58555-4|LNC|corticotropin|corticotropin
C2926297|T201|LN|58555-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926297|T201|OSN|58555-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926297|T201|MTH_LN|58555-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926297|T201|LC|58555-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926298|T201|LN|58556-2|LNC|ACTH|ACTH
C2926298|T201|MTH_LN|58556-2|LNC|ACTH|ACTH
C2926298|T201|OSN|58556-2|LNC|ACTH|ACTH
C2926298|T201|LC|58556-2|LNC|ACTH|ACTH
C2926298|T201|LN|58556-2|LNC|corticotropin|corticotropin
C2926298|T201|MTH_LN|58556-2|LNC|corticotropin|corticotropin
C2926298|T201|OSN|58556-2|LNC|corticotropin|corticotropin
C2926298|T201|LC|58556-2|LNC|corticotropin|corticotropin
C2926298|T201|LN|58556-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926298|T201|MTH_LN|58556-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926298|T201|OSN|58556-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926298|T201|LC|58556-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926299|T201|LN|58557-0|LNC|ACTH|ACTH
C2926299|T201|OSN|58557-0|LNC|ACTH|ACTH
C2926299|T201|MTH_LN|58557-0|LNC|ACTH|ACTH
C2926299|T201|LC|58557-0|LNC|ACTH|ACTH
C2926299|T201|LN|58557-0|LNC|corticotropin|corticotropin
C2926299|T201|OSN|58557-0|LNC|corticotropin|corticotropin
C2926299|T201|MTH_LN|58557-0|LNC|corticotropin|corticotropin
C2926299|T201|LC|58557-0|LNC|corticotropin|corticotropin
C2926299|T201|LN|58557-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926299|T201|OSN|58557-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926299|T201|MTH_LN|58557-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926299|T201|LC|58557-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926300|T201|LN|58558-8|LNC|ACTH|ACTH
C2926300|T201|MTH_LN|58558-8|LNC|ACTH|ACTH
C2926300|T201|LC|58558-8|LNC|ACTH|ACTH
C2926300|T201|OSN|58558-8|LNC|ACTH|ACTH
C2926300|T201|LN|58558-8|LNC|corticotropin|corticotropin
C2926300|T201|MTH_LN|58558-8|LNC|corticotropin|corticotropin
C2926300|T201|LC|58558-8|LNC|corticotropin|corticotropin
C2926300|T201|OSN|58558-8|LNC|corticotropin|corticotropin
C2926300|T201|LN|58558-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926300|T201|MTH_LN|58558-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926300|T201|LC|58558-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926300|T201|OSN|58558-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926301|T201|LN|58559-6|LNC|ACTH|ACTH
C2926301|T201|LC|58559-6|LNC|ACTH|ACTH
C2926301|T201|MTH_LN|58559-6|LNC|ACTH|ACTH
C2926301|T201|OSN|58559-6|LNC|ACTH|ACTH
C2926301|T201|LN|58559-6|LNC|corticotropin|corticotropin
C2926301|T201|LC|58559-6|LNC|corticotropin|corticotropin
C2926301|T201|MTH_LN|58559-6|LNC|corticotropin|corticotropin
C2926301|T201|OSN|58559-6|LNC|corticotropin|corticotropin
C2926301|T201|LN|58559-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926301|T201|LC|58559-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926301|T201|MTH_LN|58559-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926301|T201|OSN|58559-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926302|T201|LN|58560-4|LNC|ACTH|ACTH
C2926302|T201|OSN|58560-4|LNC|ACTH|ACTH
C2926302|T201|MTH_LN|58560-4|LNC|ACTH|ACTH
C2926302|T201|LC|58560-4|LNC|ACTH|ACTH
C2926302|T201|LN|58560-4|LNC|corticotropin|corticotropin
C2926302|T201|OSN|58560-4|LNC|corticotropin|corticotropin
C2926302|T201|MTH_LN|58560-4|LNC|corticotropin|corticotropin
C2926302|T201|LC|58560-4|LNC|corticotropin|corticotropin
C2926302|T201|LN|58560-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926302|T201|OSN|58560-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926302|T201|MTH_LN|58560-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926302|T201|LC|58560-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926303|T201|LN|58561-2|LNC|ACTH|ACTH
C2926303|T201|LC|58561-2|LNC|ACTH|ACTH
C2926303|T201|MTH_LN|58561-2|LNC|ACTH|ACTH
C2926303|T201|OSN|58561-2|LNC|ACTH|ACTH
C2926303|T201|LN|58561-2|LNC|corticotropin|corticotropin
C2926303|T201|LC|58561-2|LNC|corticotropin|corticotropin
C2926303|T201|MTH_LN|58561-2|LNC|corticotropin|corticotropin
C2926303|T201|OSN|58561-2|LNC|corticotropin|corticotropin
C2926303|T201|LN|58561-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926303|T201|LC|58561-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926303|T201|MTH_LN|58561-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926303|T201|OSN|58561-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926304|T201|LN|58562-0|LNC|ACTH|ACTH
C2926304|T201|LC|58562-0|LNC|ACTH|ACTH
C2926304|T201|MTH_LN|58562-0|LNC|ACTH|ACTH
C2926304|T201|OSN|58562-0|LNC|ACTH|ACTH
C2926304|T201|LN|58562-0|LNC|corticotropin|corticotropin
C2926304|T201|LC|58562-0|LNC|corticotropin|corticotropin
C2926304|T201|MTH_LN|58562-0|LNC|corticotropin|corticotropin
C2926304|T201|OSN|58562-0|LNC|corticotropin|corticotropin
C2926304|T201|LN|58562-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926304|T201|LC|58562-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926304|T201|MTH_LN|58562-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926304|T201|OSN|58562-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926305|T201|LN|58563-8|LNC|ACTH|ACTH
C2926305|T201|MTH_LN|58563-8|LNC|ACTH|ACTH
C2926305|T201|LC|58563-8|LNC|ACTH|ACTH
C2926305|T201|OSN|58563-8|LNC|ACTH|ACTH
C2926305|T201|LN|58563-8|LNC|corticotropin|corticotropin
C2926305|T201|MTH_LN|58563-8|LNC|corticotropin|corticotropin
C2926305|T201|LC|58563-8|LNC|corticotropin|corticotropin
C2926305|T201|OSN|58563-8|LNC|corticotropin|corticotropin
C2926305|T201|LN|58563-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926305|T201|MTH_LN|58563-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926305|T201|LC|58563-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926305|T201|OSN|58563-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926306|T201|LN|58564-6|LNC|ACTH|ACTH
C2926306|T201|LC|58564-6|LNC|ACTH|ACTH
C2926306|T201|OSN|58564-6|LNC|ACTH|ACTH
C2926306|T201|MTH_LN|58564-6|LNC|ACTH|ACTH
C2926306|T201|LN|58564-6|LNC|corticotropin|corticotropin
C2926306|T201|LC|58564-6|LNC|corticotropin|corticotropin
C2926306|T201|OSN|58564-6|LNC|corticotropin|corticotropin
C2926306|T201|MTH_LN|58564-6|LNC|corticotropin|corticotropin
C2926306|T201|LN|58564-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926306|T201|LC|58564-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926306|T201|OSN|58564-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926306|T201|MTH_LN|58564-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926307|T201|LN|58565-3|LNC|ACTH|ACTH
C2926307|T201|LC|58565-3|LNC|ACTH|ACTH
C2926307|T201|OSN|58565-3|LNC|ACTH|ACTH
C2926307|T201|MTH_LN|58565-3|LNC|ACTH|ACTH
C2926307|T201|LN|58565-3|LNC|corticotropin|corticotropin
C2926307|T201|LC|58565-3|LNC|corticotropin|corticotropin
C2926307|T201|OSN|58565-3|LNC|corticotropin|corticotropin
C2926307|T201|MTH_LN|58565-3|LNC|corticotropin|corticotropin
C2926307|T201|LN|58565-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926307|T201|LC|58565-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926307|T201|OSN|58565-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926307|T201|MTH_LN|58565-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926308|T201|LN|58566-1|LNC|ACTH|ACTH
C2926308|T201|LC|58566-1|LNC|ACTH|ACTH
C2926308|T201|OSN|58566-1|LNC|ACTH|ACTH
C2926308|T201|MTH_LN|58566-1|LNC|ACTH|ACTH
C2926308|T201|LN|58566-1|LNC|corticotropin|corticotropin
C2926308|T201|LC|58566-1|LNC|corticotropin|corticotropin
C2926308|T201|OSN|58566-1|LNC|corticotropin|corticotropin
C2926308|T201|MTH_LN|58566-1|LNC|corticotropin|corticotropin
C2926308|T201|LN|58566-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926308|T201|LC|58566-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926308|T201|OSN|58566-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926308|T201|MTH_LN|58566-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926309|T201|LN|58567-9|LNC|ACTH|ACTH
C2926309|T201|OSN|58567-9|LNC|ACTH|ACTH
C2926309|T201|MTH_LN|58567-9|LNC|ACTH|ACTH
C2926309|T201|LC|58567-9|LNC|ACTH|ACTH
C2926309|T201|LN|58567-9|LNC|corticotropin|corticotropin
C2926309|T201|OSN|58567-9|LNC|corticotropin|corticotropin
C2926309|T201|MTH_LN|58567-9|LNC|corticotropin|corticotropin
C2926309|T201|LC|58567-9|LNC|corticotropin|corticotropin
C2926309|T201|LN|58567-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926309|T201|OSN|58567-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926309|T201|MTH_LN|58567-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926309|T201|LC|58567-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926310|T201|LN|58568-7|LNC|ACTH|ACTH
C2926310|T201|MTH_LN|58568-7|LNC|ACTH|ACTH
C2926310|T201|LC|58568-7|LNC|ACTH|ACTH
C2926310|T201|OSN|58568-7|LNC|ACTH|ACTH
C2926310|T201|LN|58568-7|LNC|corticotropin|corticotropin
C2926310|T201|MTH_LN|58568-7|LNC|corticotropin|corticotropin
C2926310|T201|LC|58568-7|LNC|corticotropin|corticotropin
C2926310|T201|OSN|58568-7|LNC|corticotropin|corticotropin
C2926310|T201|LN|58568-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926310|T201|MTH_LN|58568-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926310|T201|LC|58568-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926310|T201|OSN|58568-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926311|T201|LN|58569-5|LNC|ACTH|ACTH
C2926311|T201|OSN|58569-5|LNC|ACTH|ACTH
C2926311|T201|LC|58569-5|LNC|ACTH|ACTH
C2926311|T201|MTH_LN|58569-5|LNC|ACTH|ACTH
C2926311|T201|LN|58569-5|LNC|corticotropin|corticotropin
C2926311|T201|OSN|58569-5|LNC|corticotropin|corticotropin
C2926311|T201|LC|58569-5|LNC|corticotropin|corticotropin
C2926311|T201|MTH_LN|58569-5|LNC|corticotropin|corticotropin
C2926311|T201|LN|58569-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926311|T201|OSN|58569-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926311|T201|LC|58569-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926311|T201|MTH_LN|58569-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926312|T201|LN|58570-3|LNC|ACTH|ACTH
C2926312|T201|LC|58570-3|LNC|ACTH|ACTH
C2926312|T201|OSN|58570-3|LNC|ACTH|ACTH
C2926312|T201|MTH_LN|58570-3|LNC|ACTH|ACTH
C2926312|T201|LN|58570-3|LNC|corticotropin|corticotropin
C2926312|T201|LC|58570-3|LNC|corticotropin|corticotropin
C2926312|T201|OSN|58570-3|LNC|corticotropin|corticotropin
C2926312|T201|MTH_LN|58570-3|LNC|corticotropin|corticotropin
C2926312|T201|LN|58570-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926312|T201|LC|58570-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926312|T201|OSN|58570-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926312|T201|MTH_LN|58570-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926313|T201|LN|58571-1|LNC|ACTH|ACTH
C2926313|T201|OSN|58571-1|LNC|ACTH|ACTH
C2926313|T201|LC|58571-1|LNC|ACTH|ACTH
C2926313|T201|MTH_LN|58571-1|LNC|ACTH|ACTH
C2926313|T201|LN|58571-1|LNC|corticotropin|corticotropin
C2926313|T201|OSN|58571-1|LNC|corticotropin|corticotropin
C2926313|T201|LC|58571-1|LNC|corticotropin|corticotropin
C2926313|T201|MTH_LN|58571-1|LNC|corticotropin|corticotropin
C2926313|T201|LN|58571-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926313|T201|OSN|58571-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926313|T201|LC|58571-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926313|T201|MTH_LN|58571-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926314|T201|LN|58572-9|LNC|ACTH|ACTH
C2926314|T201|LC|58572-9|LNC|ACTH|ACTH
C2926314|T201|OSN|58572-9|LNC|ACTH|ACTH
C2926314|T201|MTH_LN|58572-9|LNC|ACTH|ACTH
C2926314|T201|LN|58572-9|LNC|corticotropin|corticotropin
C2926314|T201|LC|58572-9|LNC|corticotropin|corticotropin
C2926314|T201|OSN|58572-9|LNC|corticotropin|corticotropin
C2926314|T201|MTH_LN|58572-9|LNC|corticotropin|corticotropin
C2926314|T201|LN|58572-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926314|T201|LC|58572-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926314|T201|OSN|58572-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926314|T201|MTH_LN|58572-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926315|T201|LN|58573-7|LNC|ACTH|ACTH
C2926315|T201|LC|58573-7|LNC|ACTH|ACTH
C2926315|T201|MTH_LN|58573-7|LNC|ACTH|ACTH
C2926315|T201|OSN|58573-7|LNC|ACTH|ACTH
C2926315|T201|LN|58573-7|LNC|corticotropin|corticotropin
C2926315|T201|LC|58573-7|LNC|corticotropin|corticotropin
C2926315|T201|MTH_LN|58573-7|LNC|corticotropin|corticotropin
C2926315|T201|OSN|58573-7|LNC|corticotropin|corticotropin
C2926315|T201|LN|58573-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926315|T201|LC|58573-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926315|T201|MTH_LN|58573-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926315|T201|OSN|58573-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926316|T201|LN|58574-5|LNC|ACTH|ACTH
C2926316|T201|LC|58574-5|LNC|ACTH|ACTH
C2926316|T201|OSN|58574-5|LNC|ACTH|ACTH
C2926316|T201|MTH_LN|58574-5|LNC|ACTH|ACTH
C2926316|T201|LN|58574-5|LNC|corticotropin|corticotropin
C2926316|T201|LC|58574-5|LNC|corticotropin|corticotropin
C2926316|T201|OSN|58574-5|LNC|corticotropin|corticotropin
C2926316|T201|MTH_LN|58574-5|LNC|corticotropin|corticotropin
C2926316|T201|LN|58574-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926316|T201|LC|58574-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926316|T201|OSN|58574-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926316|T201|MTH_LN|58574-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926317|T201|LN|58575-2|LNC|ACTH|ACTH
C2926317|T201|MTH_LN|58575-2|LNC|ACTH|ACTH
C2926317|T201|OSN|58575-2|LNC|ACTH|ACTH
C2926317|T201|LC|58575-2|LNC|ACTH|ACTH
C2926317|T201|LN|58575-2|LNC|corticotropin|corticotropin
C2926317|T201|MTH_LN|58575-2|LNC|corticotropin|corticotropin
C2926317|T201|OSN|58575-2|LNC|corticotropin|corticotropin
C2926317|T201|LC|58575-2|LNC|corticotropin|corticotropin
C2926317|T201|LN|58575-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926317|T201|MTH_LN|58575-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926317|T201|OSN|58575-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926317|T201|LC|58575-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926318|T201|LN|58576-0|LNC|ACTH|ACTH
C2926318|T201|OSN|58576-0|LNC|ACTH|ACTH
C2926318|T201|LC|58576-0|LNC|ACTH|ACTH
C2926318|T201|MTH_LN|58576-0|LNC|ACTH|ACTH
C2926318|T201|LN|58576-0|LNC|corticotropin|corticotropin
C2926318|T201|OSN|58576-0|LNC|corticotropin|corticotropin
C2926318|T201|LC|58576-0|LNC|corticotropin|corticotropin
C2926318|T201|MTH_LN|58576-0|LNC|corticotropin|corticotropin
C2926318|T201|LN|58576-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926318|T201|OSN|58576-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926318|T201|LC|58576-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926318|T201|MTH_LN|58576-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926319|T201|LN|58577-8|LNC|ACTH|ACTH
C2926319|T201|OSN|58577-8|LNC|ACTH|ACTH
C2926319|T201|LC|58577-8|LNC|ACTH|ACTH
C2926319|T201|MTH_LN|58577-8|LNC|ACTH|ACTH
C2926319|T201|LN|58577-8|LNC|corticotropin|corticotropin
C2926319|T201|OSN|58577-8|LNC|corticotropin|corticotropin
C2926319|T201|LC|58577-8|LNC|corticotropin|corticotropin
C2926319|T201|MTH_LN|58577-8|LNC|corticotropin|corticotropin
C2926319|T201|LN|58577-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926319|T201|OSN|58577-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926319|T201|LC|58577-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926319|T201|MTH_LN|58577-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926320|T201|LN|58578-6|LNC|ACTH|ACTH
C2926320|T201|OSN|58578-6|LNC|ACTH|ACTH
C2926320|T201|MTH_LN|58578-6|LNC|ACTH|ACTH
C2926320|T201|LC|58578-6|LNC|ACTH|ACTH
C2926320|T201|LN|58578-6|LNC|corticotropin|corticotropin
C2926320|T201|OSN|58578-6|LNC|corticotropin|corticotropin
C2926320|T201|MTH_LN|58578-6|LNC|corticotropin|corticotropin
C2926320|T201|LC|58578-6|LNC|corticotropin|corticotropin
C2926320|T201|LN|58578-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926320|T201|OSN|58578-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926320|T201|MTH_LN|58578-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926320|T201|LC|58578-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926321|T201|LN|58579-4|LNC|ACTH|ACTH
C2926321|T201|OSN|58579-4|LNC|ACTH|ACTH
C2926321|T201|LC|58579-4|LNC|ACTH|ACTH
C2926321|T201|MTH_LN|58579-4|LNC|ACTH|ACTH
C2926321|T201|LN|58579-4|LNC|corticotropin|corticotropin
C2926321|T201|OSN|58579-4|LNC|corticotropin|corticotropin
C2926321|T201|LC|58579-4|LNC|corticotropin|corticotropin
C2926321|T201|MTH_LN|58579-4|LNC|corticotropin|corticotropin
C2926321|T201|LN|58579-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926321|T201|OSN|58579-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926321|T201|LC|58579-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926321|T201|MTH_LN|58579-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926322|T201|LN|58580-2|LNC|ACTH|ACTH
C2926322|T201|OSN|58580-2|LNC|ACTH|ACTH
C2926322|T201|LC|58580-2|LNC|ACTH|ACTH
C2926322|T201|MTH_LN|58580-2|LNC|ACTH|ACTH
C2926322|T201|LN|58580-2|LNC|corticotropin|corticotropin
C2926322|T201|OSN|58580-2|LNC|corticotropin|corticotropin
C2926322|T201|LC|58580-2|LNC|corticotropin|corticotropin
C2926322|T201|MTH_LN|58580-2|LNC|corticotropin|corticotropin
C2926322|T201|LN|58580-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926322|T201|OSN|58580-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926322|T201|LC|58580-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926322|T201|MTH_LN|58580-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926323|T201|LN|58581-0|LNC|ACTH|ACTH
C2926323|T201|OSN|58581-0|LNC|ACTH|ACTH
C2926323|T201|LC|58581-0|LNC|ACTH|ACTH
C2926323|T201|MTH_LN|58581-0|LNC|ACTH|ACTH
C2926323|T201|LN|58581-0|LNC|corticotropin|corticotropin
C2926323|T201|OSN|58581-0|LNC|corticotropin|corticotropin
C2926323|T201|LC|58581-0|LNC|corticotropin|corticotropin
C2926323|T201|MTH_LN|58581-0|LNC|corticotropin|corticotropin
C2926323|T201|LN|58581-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926323|T201|OSN|58581-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926323|T201|LC|58581-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926323|T201|MTH_LN|58581-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926324|T201|LN|58582-8|LNC|ACTH|ACTH
C2926324|T201|MTH_LN|58582-8|LNC|ACTH|ACTH
C2926324|T201|OSN|58582-8|LNC|ACTH|ACTH
C2926324|T201|LC|58582-8|LNC|ACTH|ACTH
C2926324|T201|LN|58582-8|LNC|corticotropin|corticotropin
C2926324|T201|MTH_LN|58582-8|LNC|corticotropin|corticotropin
C2926324|T201|OSN|58582-8|LNC|corticotropin|corticotropin
C2926324|T201|LC|58582-8|LNC|corticotropin|corticotropin
C2926324|T201|LN|58582-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926324|T201|MTH_LN|58582-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926324|T201|OSN|58582-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926324|T201|LC|58582-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926325|T201|LN|58583-6|LNC|ACTH|ACTH
C2926325|T201|LC|58583-6|LNC|ACTH|ACTH
C2926325|T201|OSN|58583-6|LNC|ACTH|ACTH
C2926325|T201|MTH_LN|58583-6|LNC|ACTH|ACTH
C2926325|T201|LN|58583-6|LNC|corticotropin|corticotropin
C2926325|T201|LC|58583-6|LNC|corticotropin|corticotropin
C2926325|T201|OSN|58583-6|LNC|corticotropin|corticotropin
C2926325|T201|MTH_LN|58583-6|LNC|corticotropin|corticotropin
C2926325|T201|LN|58583-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926325|T201|LC|58583-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926325|T201|OSN|58583-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926325|T201|MTH_LN|58583-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926326|T201|LN|58584-4|LNC|ACTH|ACTH
C2926326|T201|LC|58584-4|LNC|ACTH|ACTH
C2926326|T201|OSN|58584-4|LNC|ACTH|ACTH
C2926326|T201|MTH_LN|58584-4|LNC|ACTH|ACTH
C2926326|T201|LN|58584-4|LNC|corticotropin|corticotropin
C2926326|T201|LC|58584-4|LNC|corticotropin|corticotropin
C2926326|T201|OSN|58584-4|LNC|corticotropin|corticotropin
C2926326|T201|MTH_LN|58584-4|LNC|corticotropin|corticotropin
C2926326|T201|LN|58584-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926326|T201|LC|58584-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926326|T201|OSN|58584-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926326|T201|MTH_LN|58584-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926327|T201|LN|58585-1|LNC|ACTH|ACTH
C2926327|T201|OSN|58585-1|LNC|ACTH|ACTH
C2926327|T201|MTH_LN|58585-1|LNC|ACTH|ACTH
C2926327|T201|LC|58585-1|LNC|ACTH|ACTH
C2926327|T201|LN|58585-1|LNC|corticotropin|corticotropin
C2926327|T201|OSN|58585-1|LNC|corticotropin|corticotropin
C2926327|T201|MTH_LN|58585-1|LNC|corticotropin|corticotropin
C2926327|T201|LC|58585-1|LNC|corticotropin|corticotropin
C2926327|T201|LN|58585-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926327|T201|OSN|58585-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926327|T201|MTH_LN|58585-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926327|T201|LC|58585-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926328|T201|LN|58586-9|LNC|ACTH|ACTH
C2926328|T201|OSN|58586-9|LNC|ACTH|ACTH
C2926328|T201|LC|58586-9|LNC|ACTH|ACTH
C2926328|T201|MTH_LN|58586-9|LNC|ACTH|ACTH
C2926328|T201|LN|58586-9|LNC|corticotropin|corticotropin
C2926328|T201|OSN|58586-9|LNC|corticotropin|corticotropin
C2926328|T201|LC|58586-9|LNC|corticotropin|corticotropin
C2926328|T201|MTH_LN|58586-9|LNC|corticotropin|corticotropin
C2926328|T201|LN|58586-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926328|T201|OSN|58586-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926328|T201|LC|58586-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926328|T201|MTH_LN|58586-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926329|T201|LN|58587-7|LNC|ACTH|ACTH
C2926329|T201|LC|58587-7|LNC|ACTH|ACTH
C2926329|T201|MTH_LN|58587-7|LNC|ACTH|ACTH
C2926329|T201|OSN|58587-7|LNC|ACTH|ACTH
C2926329|T201|LN|58587-7|LNC|corticotropin|corticotropin
C2926329|T201|LC|58587-7|LNC|corticotropin|corticotropin
C2926329|T201|MTH_LN|58587-7|LNC|corticotropin|corticotropin
C2926329|T201|OSN|58587-7|LNC|corticotropin|corticotropin
C2926329|T201|LN|58587-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926329|T201|LC|58587-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926329|T201|MTH_LN|58587-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926329|T201|OSN|58587-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926330|T201|LN|58588-5|LNC|ACTH|ACTH
C2926330|T201|MTH_LN|58588-5|LNC|ACTH|ACTH
C2926330|T201|OSN|58588-5|LNC|ACTH|ACTH
C2926330|T201|LC|58588-5|LNC|ACTH|ACTH
C2926330|T201|LN|58588-5|LNC|corticotropin|corticotropin
C2926330|T201|MTH_LN|58588-5|LNC|corticotropin|corticotropin
C2926330|T201|OSN|58588-5|LNC|corticotropin|corticotropin
C2926330|T201|LC|58588-5|LNC|corticotropin|corticotropin
C2926330|T201|LN|58588-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926330|T201|MTH_LN|58588-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926330|T201|OSN|58588-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926330|T201|LC|58588-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926331|T201|LN|58589-3|LNC|ACTH|ACTH
C2926331|T201|OSN|58589-3|LNC|ACTH|ACTH
C2926331|T201|LC|58589-3|LNC|ACTH|ACTH
C2926331|T201|MTH_LN|58589-3|LNC|ACTH|ACTH
C2926331|T201|LN|58589-3|LNC|corticotropin|corticotropin
C2926331|T201|OSN|58589-3|LNC|corticotropin|corticotropin
C2926331|T201|LC|58589-3|LNC|corticotropin|corticotropin
C2926331|T201|MTH_LN|58589-3|LNC|corticotropin|corticotropin
C2926331|T201|LN|58589-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926331|T201|OSN|58589-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926331|T201|LC|58589-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926331|T201|MTH_LN|58589-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926332|T201|LN|58590-1|LNC|ACTH|ACTH
C2926332|T201|MTH_LN|58590-1|LNC|ACTH|ACTH
C2926332|T201|LC|58590-1|LNC|ACTH|ACTH
C2926332|T201|OSN|58590-1|LNC|ACTH|ACTH
C2926332|T201|LN|58590-1|LNC|corticotropin|corticotropin
C2926332|T201|MTH_LN|58590-1|LNC|corticotropin|corticotropin
C2926332|T201|LC|58590-1|LNC|corticotropin|corticotropin
C2926332|T201|OSN|58590-1|LNC|corticotropin|corticotropin
C2926332|T201|LN|58590-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926332|T201|MTH_LN|58590-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926332|T201|LC|58590-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926332|T201|OSN|58590-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926333|T201|LN|58591-9|LNC|ACTH|ACTH
C2926333|T201|LC|58591-9|LNC|ACTH|ACTH
C2926333|T201|MTH_LN|58591-9|LNC|ACTH|ACTH
C2926333|T201|OSN|58591-9|LNC|ACTH|ACTH
C2926333|T201|LN|58591-9|LNC|corticotropin|corticotropin
C2926333|T201|LC|58591-9|LNC|corticotropin|corticotropin
C2926333|T201|MTH_LN|58591-9|LNC|corticotropin|corticotropin
C2926333|T201|OSN|58591-9|LNC|corticotropin|corticotropin
C2926333|T201|LN|58591-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926333|T201|LC|58591-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926333|T201|MTH_LN|58591-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926333|T201|OSN|58591-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926334|T201|LN|58592-7|LNC|ACTH|ACTH
C2926334|T201|MTH_LN|58592-7|LNC|ACTH|ACTH
C2926334|T201|LC|58592-7|LNC|ACTH|ACTH
C2926334|T201|OSN|58592-7|LNC|ACTH|ACTH
C2926334|T201|LN|58592-7|LNC|corticotropin|corticotropin
C2926334|T201|MTH_LN|58592-7|LNC|corticotropin|corticotropin
C2926334|T201|LC|58592-7|LNC|corticotropin|corticotropin
C2926334|T201|OSN|58592-7|LNC|corticotropin|corticotropin
C2926334|T201|LN|58592-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926334|T201|MTH_LN|58592-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926334|T201|LC|58592-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926334|T201|OSN|58592-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926335|T201|LN|58593-5|LNC|ACTH|ACTH
C2926335|T201|LC|58593-5|LNC|ACTH|ACTH
C2926335|T201|OSN|58593-5|LNC|ACTH|ACTH
C2926335|T201|MTH_LN|58593-5|LNC|ACTH|ACTH
C2926335|T201|LN|58593-5|LNC|corticotropin|corticotropin
C2926335|T201|LC|58593-5|LNC|corticotropin|corticotropin
C2926335|T201|OSN|58593-5|LNC|corticotropin|corticotropin
C2926335|T201|MTH_LN|58593-5|LNC|corticotropin|corticotropin
C2926335|T201|LN|58593-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926335|T201|LC|58593-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926335|T201|OSN|58593-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926335|T201|MTH_LN|58593-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926336|T201|LN|58594-3|LNC|ACTH|ACTH
C2926336|T201|MTH_LN|58594-3|LNC|ACTH|ACTH
C2926336|T201|OSN|58594-3|LNC|ACTH|ACTH
C2926336|T201|LC|58594-3|LNC|ACTH|ACTH
C2926336|T201|LN|58594-3|LNC|corticotropin|corticotropin
C2926336|T201|MTH_LN|58594-3|LNC|corticotropin|corticotropin
C2926336|T201|OSN|58594-3|LNC|corticotropin|corticotropin
C2926336|T201|LC|58594-3|LNC|corticotropin|corticotropin
C2926336|T201|LN|58594-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926336|T201|MTH_LN|58594-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926336|T201|OSN|58594-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926336|T201|LC|58594-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926337|T201|LN|58595-0|LNC|ACTH|ACTH
C2926337|T201|LC|58595-0|LNC|ACTH|ACTH
C2926337|T201|MTH_LN|58595-0|LNC|ACTH|ACTH
C2926337|T201|OSN|58595-0|LNC|ACTH|ACTH
C2926337|T201|LN|58595-0|LNC|corticotropin|corticotropin
C2926337|T201|LC|58595-0|LNC|corticotropin|corticotropin
C2926337|T201|MTH_LN|58595-0|LNC|corticotropin|corticotropin
C2926337|T201|OSN|58595-0|LNC|corticotropin|corticotropin
C2926337|T201|LN|58595-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926337|T201|LC|58595-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926337|T201|MTH_LN|58595-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926337|T201|OSN|58595-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926338|T201|LN|58596-8|LNC|ACTH|ACTH
C2926338|T201|MTH_LN|58596-8|LNC|ACTH|ACTH
C2926338|T201|OSN|58596-8|LNC|ACTH|ACTH
C2926338|T201|LC|58596-8|LNC|ACTH|ACTH
C2926338|T201|LN|58596-8|LNC|corticotropin|corticotropin
C2926338|T201|MTH_LN|58596-8|LNC|corticotropin|corticotropin
C2926338|T201|OSN|58596-8|LNC|corticotropin|corticotropin
C2926338|T201|LC|58596-8|LNC|corticotropin|corticotropin
C2926338|T201|LN|58596-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926338|T201|MTH_LN|58596-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926338|T201|OSN|58596-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926338|T201|LC|58596-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926339|T201|LN|58597-6|LNC|ACTH|ACTH
C2926339|T201|OSN|58597-6|LNC|ACTH|ACTH
C2926339|T201|MTH_LN|58597-6|LNC|ACTH|ACTH
C2926339|T201|LC|58597-6|LNC|ACTH|ACTH
C2926339|T201|LN|58597-6|LNC|corticotropin|corticotropin
C2926339|T201|OSN|58597-6|LNC|corticotropin|corticotropin
C2926339|T201|MTH_LN|58597-6|LNC|corticotropin|corticotropin
C2926339|T201|LC|58597-6|LNC|corticotropin|corticotropin
C2926339|T201|LN|58597-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926339|T201|OSN|58597-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926339|T201|MTH_LN|58597-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926339|T201|LC|58597-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926340|T201|LN|58598-4|LNC|ACTH|ACTH
C2926340|T201|OSN|58598-4|LNC|ACTH|ACTH
C2926340|T201|MTH_LN|58598-4|LNC|ACTH|ACTH
C2926340|T201|LC|58598-4|LNC|ACTH|ACTH
C2926340|T201|LN|58598-4|LNC|corticotropin|corticotropin
C2926340|T201|OSN|58598-4|LNC|corticotropin|corticotropin
C2926340|T201|MTH_LN|58598-4|LNC|corticotropin|corticotropin
C2926340|T201|LC|58598-4|LNC|corticotropin|corticotropin
C2926340|T201|LN|58598-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926340|T201|OSN|58598-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926340|T201|MTH_LN|58598-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926340|T201|LC|58598-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926341|T201|LN|58599-2|LNC|ACTH|ACTH
C2926341|T201|LC|58599-2|LNC|ACTH|ACTH
C2926341|T201|MTH_LN|58599-2|LNC|ACTH|ACTH
C2926341|T201|OSN|58599-2|LNC|ACTH|ACTH
C2926341|T201|LN|58599-2|LNC|corticotropin|corticotropin
C2926341|T201|LC|58599-2|LNC|corticotropin|corticotropin
C2926341|T201|MTH_LN|58599-2|LNC|corticotropin|corticotropin
C2926341|T201|OSN|58599-2|LNC|corticotropin|corticotropin
C2926341|T201|LN|58599-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926341|T201|LC|58599-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926341|T201|MTH_LN|58599-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926341|T201|OSN|58599-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926342|T201|LN|58600-8|LNC|ACTH|ACTH
C2926342|T201|MTH_LN|58600-8|LNC|ACTH|ACTH
C2926342|T201|OSN|58600-8|LNC|ACTH|ACTH
C2926342|T201|LC|58600-8|LNC|ACTH|ACTH
C2926342|T201|LN|58600-8|LNC|corticotropin|corticotropin
C2926342|T201|MTH_LN|58600-8|LNC|corticotropin|corticotropin
C2926342|T201|OSN|58600-8|LNC|corticotropin|corticotropin
C2926342|T201|LC|58600-8|LNC|corticotropin|corticotropin
C2926342|T201|LN|58600-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926342|T201|MTH_LN|58600-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926342|T201|OSN|58600-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926342|T201|LC|58600-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926343|T201|LN|58601-6|LNC|ACTH|ACTH
C2926343|T201|MTH_LN|58601-6|LNC|ACTH|ACTH
C2926343|T201|OSN|58601-6|LNC|ACTH|ACTH
C2926343|T201|LC|58601-6|LNC|ACTH|ACTH
C2926343|T201|LN|58601-6|LNC|corticotropin|corticotropin
C2926343|T201|MTH_LN|58601-6|LNC|corticotropin|corticotropin
C2926343|T201|OSN|58601-6|LNC|corticotropin|corticotropin
C2926343|T201|LC|58601-6|LNC|corticotropin|corticotropin
C2926343|T201|LN|58601-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926343|T201|MTH_LN|58601-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926343|T201|OSN|58601-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926343|T201|LC|58601-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926344|T201|LN|58602-4|LNC|ACTH|ACTH
C2926344|T201|OSN|58602-4|LNC|ACTH|ACTH
C2926344|T201|LC|58602-4|LNC|ACTH|ACTH
C2926344|T201|MTH_LN|58602-4|LNC|ACTH|ACTH
C2926344|T201|LN|58602-4|LNC|corticotropin|corticotropin
C2926344|T201|OSN|58602-4|LNC|corticotropin|corticotropin
C2926344|T201|LC|58602-4|LNC|corticotropin|corticotropin
C2926344|T201|MTH_LN|58602-4|LNC|corticotropin|corticotropin
C2926344|T201|LN|58602-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926344|T201|OSN|58602-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926344|T201|LC|58602-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926344|T201|MTH_LN|58602-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926345|T201|LN|58603-2|LNC|ACTH|ACTH
C2926345|T201|LC|58603-2|LNC|ACTH|ACTH
C2926345|T201|MTH_LN|58603-2|LNC|ACTH|ACTH
C2926345|T201|OSN|58603-2|LNC|ACTH|ACTH
C2926345|T201|LN|58603-2|LNC|corticotropin|corticotropin
C2926345|T201|LC|58603-2|LNC|corticotropin|corticotropin
C2926345|T201|MTH_LN|58603-2|LNC|corticotropin|corticotropin
C2926345|T201|OSN|58603-2|LNC|corticotropin|corticotropin
C2926345|T201|LN|58603-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926345|T201|LC|58603-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926345|T201|MTH_LN|58603-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926345|T201|OSN|58603-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926346|T201|LN|58604-0|LNC|ACTH|ACTH
C2926346|T201|LC|58604-0|LNC|ACTH|ACTH
C2926346|T201|MTH_LN|58604-0|LNC|ACTH|ACTH
C2926346|T201|OSN|58604-0|LNC|ACTH|ACTH
C2926346|T201|LN|58604-0|LNC|corticotropin|corticotropin
C2926346|T201|LC|58604-0|LNC|corticotropin|corticotropin
C2926346|T201|MTH_LN|58604-0|LNC|corticotropin|corticotropin
C2926346|T201|OSN|58604-0|LNC|corticotropin|corticotropin
C2926346|T201|LN|58604-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926346|T201|LC|58604-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926346|T201|MTH_LN|58604-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926346|T201|OSN|58604-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926347|T201|LN|58605-7|LNC|ACTH|ACTH
C2926347|T201|OSN|58605-7|LNC|ACTH|ACTH
C2926347|T201|MTH_LN|58605-7|LNC|ACTH|ACTH
C2926347|T201|LC|58605-7|LNC|ACTH|ACTH
C2926347|T201|LN|58605-7|LNC|corticotropin|corticotropin
C2926347|T201|OSN|58605-7|LNC|corticotropin|corticotropin
C2926347|T201|MTH_LN|58605-7|LNC|corticotropin|corticotropin
C2926347|T201|LC|58605-7|LNC|corticotropin|corticotropin
C2926347|T201|LN|58605-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926347|T201|OSN|58605-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926347|T201|MTH_LN|58605-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926347|T201|LC|58605-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926348|T201|LN|58606-5|LNC|ACTH|ACTH
C2926348|T201|MTH_LN|58606-5|LNC|ACTH|ACTH
C2926348|T201|OSN|58606-5|LNC|ACTH|ACTH
C2926348|T201|LC|58606-5|LNC|ACTH|ACTH
C2926348|T201|LN|58606-5|LNC|corticotropin|corticotropin
C2926348|T201|MTH_LN|58606-5|LNC|corticotropin|corticotropin
C2926348|T201|OSN|58606-5|LNC|corticotropin|corticotropin
C2926348|T201|LC|58606-5|LNC|corticotropin|corticotropin
C2926348|T201|LN|58606-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926348|T201|MTH_LN|58606-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926348|T201|OSN|58606-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926348|T201|LC|58606-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926349|T201|LN|58607-3|LNC|ACTH|ACTH
C2926349|T201|LC|58607-3|LNC|ACTH|ACTH
C2926349|T201|OSN|58607-3|LNC|ACTH|ACTH
C2926349|T201|MTH_LN|58607-3|LNC|ACTH|ACTH
C2926349|T201|LN|58607-3|LNC|corticotropin|corticotropin
C2926349|T201|LC|58607-3|LNC|corticotropin|corticotropin
C2926349|T201|OSN|58607-3|LNC|corticotropin|corticotropin
C2926349|T201|MTH_LN|58607-3|LNC|corticotropin|corticotropin
C2926349|T201|LN|58607-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926349|T201|LC|58607-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926349|T201|OSN|58607-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926349|T201|MTH_LN|58607-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926350|T201|LN|58608-1|LNC|ACTH|ACTH
C2926350|T201|MTH_LN|58608-1|LNC|ACTH|ACTH
C2926350|T201|LC|58608-1|LNC|ACTH|ACTH
C2926350|T201|OSN|58608-1|LNC|ACTH|ACTH
C2926350|T201|LN|58608-1|LNC|corticotropin|corticotropin
C2926350|T201|MTH_LN|58608-1|LNC|corticotropin|corticotropin
C2926350|T201|LC|58608-1|LNC|corticotropin|corticotropin
C2926350|T201|OSN|58608-1|LNC|corticotropin|corticotropin
C2926350|T201|LN|58608-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926350|T201|MTH_LN|58608-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926350|T201|LC|58608-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926350|T201|OSN|58608-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926351|T201|LN|58609-9|LNC|ACTH|ACTH
C2926351|T201|MTH_LN|58609-9|LNC|ACTH|ACTH
C2926351|T201|OSN|58609-9|LNC|ACTH|ACTH
C2926351|T201|LC|58609-9|LNC|ACTH|ACTH
C2926351|T201|LN|58609-9|LNC|corticotropin|corticotropin
C2926351|T201|MTH_LN|58609-9|LNC|corticotropin|corticotropin
C2926351|T201|OSN|58609-9|LNC|corticotropin|corticotropin
C2926351|T201|LC|58609-9|LNC|corticotropin|corticotropin
C2926351|T201|LN|58609-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926351|T201|MTH_LN|58609-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926351|T201|OSN|58609-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926351|T201|LC|58609-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926352|T201|LN|58610-7|LNC|ACTH|ACTH
C2926352|T201|LC|58610-7|LNC|ACTH|ACTH
C2926352|T201|MTH_LN|58610-7|LNC|ACTH|ACTH
C2926352|T201|OSN|58610-7|LNC|ACTH|ACTH
C2926352|T201|LN|58610-7|LNC|corticotropin|corticotropin
C2926352|T201|LC|58610-7|LNC|corticotropin|corticotropin
C2926352|T201|MTH_LN|58610-7|LNC|corticotropin|corticotropin
C2926352|T201|OSN|58610-7|LNC|corticotropin|corticotropin
C2926352|T201|LN|58610-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926352|T201|LC|58610-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926352|T201|MTH_LN|58610-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926352|T201|OSN|58610-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926353|T201|LN|58611-5|LNC|ACTH|ACTH
C2926353|T201|OSN|58611-5|LNC|ACTH|ACTH
C2926353|T201|LC|58611-5|LNC|ACTH|ACTH
C2926353|T201|MTH_LN|58611-5|LNC|ACTH|ACTH
C2926353|T201|LN|58611-5|LNC|corticotropin|corticotropin
C2926353|T201|OSN|58611-5|LNC|corticotropin|corticotropin
C2926353|T201|LC|58611-5|LNC|corticotropin|corticotropin
C2926353|T201|MTH_LN|58611-5|LNC|corticotropin|corticotropin
C2926353|T201|LN|58611-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926353|T201|OSN|58611-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926353|T201|LC|58611-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926353|T201|MTH_LN|58611-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926354|T201|LN|58612-3|LNC|ACTH|ACTH
C2926354|T201|OSN|58612-3|LNC|ACTH|ACTH
C2926354|T201|LC|58612-3|LNC|ACTH|ACTH
C2926354|T201|MTH_LN|58612-3|LNC|ACTH|ACTH
C2926354|T201|LN|58612-3|LNC|corticotropin|corticotropin
C2926354|T201|OSN|58612-3|LNC|corticotropin|corticotropin
C2926354|T201|LC|58612-3|LNC|corticotropin|corticotropin
C2926354|T201|MTH_LN|58612-3|LNC|corticotropin|corticotropin
C2926354|T201|LN|58612-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926354|T201|OSN|58612-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926354|T201|LC|58612-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926354|T201|MTH_LN|58612-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926355|T201|LN|58613-1|LNC|ACTH|ACTH
C2926355|T201|OSN|58613-1|LNC|ACTH|ACTH
C2926355|T201|LC|58613-1|LNC|ACTH|ACTH
C2926355|T201|MTH_LN|58613-1|LNC|ACTH|ACTH
C2926355|T201|LN|58613-1|LNC|corticotropin|corticotropin
C2926355|T201|OSN|58613-1|LNC|corticotropin|corticotropin
C2926355|T201|LC|58613-1|LNC|corticotropin|corticotropin
C2926355|T201|MTH_LN|58613-1|LNC|corticotropin|corticotropin
C2926355|T201|LN|58613-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926355|T201|OSN|58613-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926355|T201|LC|58613-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926355|T201|MTH_LN|58613-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926356|T201|LN|58614-9|LNC|ACTH|ACTH
C2926356|T201|MTH_LN|58614-9|LNC|ACTH|ACTH
C2926356|T201|OSN|58614-9|LNC|ACTH|ACTH
C2926356|T201|LC|58614-9|LNC|ACTH|ACTH
C2926356|T201|LN|58614-9|LNC|corticotropin|corticotropin
C2926356|T201|MTH_LN|58614-9|LNC|corticotropin|corticotropin
C2926356|T201|OSN|58614-9|LNC|corticotropin|corticotropin
C2926356|T201|LC|58614-9|LNC|corticotropin|corticotropin
C2926356|T201|LN|58614-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926356|T201|MTH_LN|58614-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926356|T201|OSN|58614-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926356|T201|LC|58614-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926357|T201|LN|58615-6|LNC|ACTH|ACTH
C2926357|T201|LC|58615-6|LNC|ACTH|ACTH
C2926357|T201|MTH_LN|58615-6|LNC|ACTH|ACTH
C2926357|T201|OSN|58615-6|LNC|ACTH|ACTH
C2926357|T201|LN|58615-6|LNC|corticotropin|corticotropin
C2926357|T201|LC|58615-6|LNC|corticotropin|corticotropin
C2926357|T201|MTH_LN|58615-6|LNC|corticotropin|corticotropin
C2926357|T201|OSN|58615-6|LNC|corticotropin|corticotropin
C2926357|T201|LN|58615-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926357|T201|LC|58615-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926357|T201|MTH_LN|58615-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926357|T201|OSN|58615-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926358|T201|LN|58616-4|LNC|ACTH|ACTH
C2926358|T201|MTH_LN|58616-4|LNC|ACTH|ACTH
C2926358|T201|OSN|58616-4|LNC|ACTH|ACTH
C2926358|T201|LC|58616-4|LNC|ACTH|ACTH
C2926358|T201|LN|58616-4|LNC|corticotropin|corticotropin
C2926358|T201|MTH_LN|58616-4|LNC|corticotropin|corticotropin
C2926358|T201|OSN|58616-4|LNC|corticotropin|corticotropin
C2926358|T201|LC|58616-4|LNC|corticotropin|corticotropin
C2926358|T201|LN|58616-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926358|T201|MTH_LN|58616-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926358|T201|OSN|58616-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926358|T201|LC|58616-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926359|T201|LN|58617-2|LNC|ACTH|ACTH
C2926359|T201|OSN|58617-2|LNC|ACTH|ACTH
C2926359|T201|MTH_LN|58617-2|LNC|ACTH|ACTH
C2926359|T201|LC|58617-2|LNC|ACTH|ACTH
C2926359|T201|LN|58617-2|LNC|corticotropin|corticotropin
C2926359|T201|OSN|58617-2|LNC|corticotropin|corticotropin
C2926359|T201|MTH_LN|58617-2|LNC|corticotropin|corticotropin
C2926359|T201|LC|58617-2|LNC|corticotropin|corticotropin
C2926359|T201|LN|58617-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926359|T201|OSN|58617-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926359|T201|MTH_LN|58617-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926359|T201|LC|58617-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926360|T201|LN|58618-0|LNC|ACTH|ACTH
C2926360|T201|LC|58618-0|LNC|ACTH|ACTH
C2926360|T201|MTH_LN|58618-0|LNC|ACTH|ACTH
C2926360|T201|OSN|58618-0|LNC|ACTH|ACTH
C2926360|T201|LN|58618-0|LNC|corticotropin|corticotropin
C2926360|T201|LC|58618-0|LNC|corticotropin|corticotropin
C2926360|T201|MTH_LN|58618-0|LNC|corticotropin|corticotropin
C2926360|T201|OSN|58618-0|LNC|corticotropin|corticotropin
C2926360|T201|LN|58618-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926360|T201|LC|58618-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926360|T201|MTH_LN|58618-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926360|T201|OSN|58618-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926361|T201|LN|58619-8|LNC|ACTH|ACTH
C2926361|T201|MTH_LN|58619-8|LNC|ACTH|ACTH
C2926361|T201|LC|58619-8|LNC|ACTH|ACTH
C2926361|T201|OSN|58619-8|LNC|ACTH|ACTH
C2926361|T201|LN|58619-8|LNC|corticotropin|corticotropin
C2926361|T201|MTH_LN|58619-8|LNC|corticotropin|corticotropin
C2926361|T201|LC|58619-8|LNC|corticotropin|corticotropin
C2926361|T201|OSN|58619-8|LNC|corticotropin|corticotropin
C2926361|T201|LN|58619-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926361|T201|MTH_LN|58619-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926361|T201|LC|58619-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926361|T201|OSN|58619-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926362|T201|LN|58620-6|LNC|ACTH|ACTH
C2926362|T201|OSN|58620-6|LNC|ACTH|ACTH
C2926362|T201|MTH_LN|58620-6|LNC|ACTH|ACTH
C2926362|T201|LC|58620-6|LNC|ACTH|ACTH
C2926362|T201|LN|58620-6|LNC|corticotropin|corticotropin
C2926362|T201|OSN|58620-6|LNC|corticotropin|corticotropin
C2926362|T201|MTH_LN|58620-6|LNC|corticotropin|corticotropin
C2926362|T201|LC|58620-6|LNC|corticotropin|corticotropin
C2926362|T201|LN|58620-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926362|T201|OSN|58620-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926362|T201|MTH_LN|58620-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926362|T201|LC|58620-6|LNC|adrenocorticotropin|adrenocorticotropin
C2926363|T201|LN|58621-4|LNC|ACTH|ACTH
C2926363|T201|MTH_LN|58621-4|LNC|ACTH|ACTH
C2926363|T201|OSN|58621-4|LNC|ACTH|ACTH
C2926363|T201|LC|58621-4|LNC|ACTH|ACTH
C2926363|T201|LN|58621-4|LNC|corticotropin|corticotropin
C2926363|T201|MTH_LN|58621-4|LNC|corticotropin|corticotropin
C2926363|T201|OSN|58621-4|LNC|corticotropin|corticotropin
C2926363|T201|LC|58621-4|LNC|corticotropin|corticotropin
C2926363|T201|LN|58621-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926363|T201|MTH_LN|58621-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926363|T201|OSN|58621-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926363|T201|LC|58621-4|LNC|adrenocorticotropin|adrenocorticotropin
C2926364|T201|LN|58622-2|LNC|ACTH|ACTH
C2926364|T201|OSN|58622-2|LNC|ACTH|ACTH
C2926364|T201|LC|58622-2|LNC|ACTH|ACTH
C2926364|T201|MTH_LN|58622-2|LNC|ACTH|ACTH
C2926364|T201|LN|58622-2|LNC|corticotropin|corticotropin
C2926364|T201|OSN|58622-2|LNC|corticotropin|corticotropin
C2926364|T201|LC|58622-2|LNC|corticotropin|corticotropin
C2926364|T201|MTH_LN|58622-2|LNC|corticotropin|corticotropin
C2926364|T201|LN|58622-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926364|T201|OSN|58622-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926364|T201|LC|58622-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926364|T201|MTH_LN|58622-2|LNC|adrenocorticotropin|adrenocorticotropin
C2926365|T201|LN|58623-0|LNC|ACTH|ACTH
C2926365|T201|MTH_LN|58623-0|LNC|ACTH|ACTH
C2926365|T201|LC|58623-0|LNC|ACTH|ACTH
C2926365|T201|OSN|58623-0|LNC|ACTH|ACTH
C2926365|T201|LN|58623-0|LNC|corticotropin|corticotropin
C2926365|T201|MTH_LN|58623-0|LNC|corticotropin|corticotropin
C2926365|T201|LC|58623-0|LNC|corticotropin|corticotropin
C2926365|T201|OSN|58623-0|LNC|corticotropin|corticotropin
C2926365|T201|LN|58623-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926365|T201|MTH_LN|58623-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926365|T201|LC|58623-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926365|T201|OSN|58623-0|LNC|adrenocorticotropin|adrenocorticotropin
C2926366|T201|LN|58624-8|LNC|ACTH|ACTH
C2926366|T201|OSN|58624-8|LNC|ACTH|ACTH
C2926366|T201|LC|58624-8|LNC|ACTH|ACTH
C2926366|T201|MTH_LN|58624-8|LNC|ACTH|ACTH
C2926366|T201|LN|58624-8|LNC|corticotropin|corticotropin
C2926366|T201|OSN|58624-8|LNC|corticotropin|corticotropin
C2926366|T201|LC|58624-8|LNC|corticotropin|corticotropin
C2926366|T201|MTH_LN|58624-8|LNC|corticotropin|corticotropin
C2926366|T201|LN|58624-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926366|T201|OSN|58624-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926366|T201|LC|58624-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926366|T201|MTH_LN|58624-8|LNC|adrenocorticotropin|adrenocorticotropin
C2926367|T201|LN|58625-5|LNC|ACTH|ACTH
C2926367|T201|OSN|58625-5|LNC|ACTH|ACTH
C2926367|T201|LC|58625-5|LNC|ACTH|ACTH
C2926367|T201|MTH_LN|58625-5|LNC|ACTH|ACTH
C2926367|T201|LN|58625-5|LNC|corticotropin|corticotropin
C2926367|T201|OSN|58625-5|LNC|corticotropin|corticotropin
C2926367|T201|LC|58625-5|LNC|corticotropin|corticotropin
C2926367|T201|MTH_LN|58625-5|LNC|corticotropin|corticotropin
C2926367|T201|LN|58625-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926367|T201|OSN|58625-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926367|T201|LC|58625-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926367|T201|MTH_LN|58625-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926368|T201|LN|58626-3|LNC|ACTH|ACTH
C2926368|T201|OSN|58626-3|LNC|ACTH|ACTH
C2926368|T201|LC|58626-3|LNC|ACTH|ACTH
C2926368|T201|MTH_LN|58626-3|LNC|ACTH|ACTH
C2926368|T201|LN|58626-3|LNC|corticotropin|corticotropin
C2926368|T201|OSN|58626-3|LNC|corticotropin|corticotropin
C2926368|T201|LC|58626-3|LNC|corticotropin|corticotropin
C2926368|T201|MTH_LN|58626-3|LNC|corticotropin|corticotropin
C2926368|T201|LN|58626-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926368|T201|OSN|58626-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926368|T201|LC|58626-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926368|T201|MTH_LN|58626-3|LNC|adrenocorticotropin|adrenocorticotropin
C2926369|T201|LN|58627-1|LNC|ACTH|ACTH
C2926369|T201|LC|58627-1|LNC|ACTH|ACTH
C2926369|T201|MTH_LN|58627-1|LNC|ACTH|ACTH
C2926369|T201|OSN|58627-1|LNC|ACTH|ACTH
C2926369|T201|LN|58627-1|LNC|corticotropin|corticotropin
C2926369|T201|LC|58627-1|LNC|corticotropin|corticotropin
C2926369|T201|MTH_LN|58627-1|LNC|corticotropin|corticotropin
C2926369|T201|OSN|58627-1|LNC|corticotropin|corticotropin
C2926369|T201|LN|58627-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926369|T201|LC|58627-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926369|T201|MTH_LN|58627-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926369|T201|OSN|58627-1|LNC|adrenocorticotropin|adrenocorticotropin
C2926370|T201|LN|58628-9|LNC|ACTH|ACTH
C2926370|T201|OSN|58628-9|LNC|ACTH|ACTH
C2926370|T201|LC|58628-9|LNC|ACTH|ACTH
C2926370|T201|MTH_LN|58628-9|LNC|ACTH|ACTH
C2926370|T201|LN|58628-9|LNC|corticotropin|corticotropin
C2926370|T201|OSN|58628-9|LNC|corticotropin|corticotropin
C2926370|T201|LC|58628-9|LNC|corticotropin|corticotropin
C2926370|T201|MTH_LN|58628-9|LNC|corticotropin|corticotropin
C2926370|T201|LN|58628-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926370|T201|OSN|58628-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926370|T201|LC|58628-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926370|T201|MTH_LN|58628-9|LNC|adrenocorticotropin|adrenocorticotropin
C2926371|T201|LN|58629-7|LNC|ACTH|ACTH
C2926371|T201|MTH_LN|58629-7|LNC|ACTH|ACTH
C2926371|T201|LC|58629-7|LNC|ACTH|ACTH
C2926371|T201|OSN|58629-7|LNC|ACTH|ACTH
C2926371|T201|LN|58629-7|LNC|corticotropin|corticotropin
C2926371|T201|MTH_LN|58629-7|LNC|corticotropin|corticotropin
C2926371|T201|LC|58629-7|LNC|corticotropin|corticotropin
C2926371|T201|OSN|58629-7|LNC|corticotropin|corticotropin
C2926371|T201|LN|58629-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926371|T201|MTH_LN|58629-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926371|T201|LC|58629-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926371|T201|OSN|58629-7|LNC|adrenocorticotropin|adrenocorticotropin
C2926372|T201|LN|58630-5|LNC|ACTH|ACTH
C2926372|T201|MTH_LN|58630-5|LNC|ACTH|ACTH
C2926372|T201|OSN|58630-5|LNC|ACTH|ACTH
C2926372|T201|LC|58630-5|LNC|ACTH|ACTH
C2926372|T201|LN|58630-5|LNC|corticotropin|corticotropin
C2926372|T201|MTH_LN|58630-5|LNC|corticotropin|corticotropin
C2926372|T201|OSN|58630-5|LNC|corticotropin|corticotropin
C2926372|T201|LC|58630-5|LNC|corticotropin|corticotropin
C2926372|T201|LN|58630-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926372|T201|MTH_LN|58630-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926372|T201|OSN|58630-5|LNC|adrenocorticotropin|adrenocorticotropin
C2926372|T201|LC|58630-5|LNC|adrenocorticotropin|adrenocorticotropin
C2966814|T201|LN|60014-8|LNC|ACTH|ACTH
C2966814|T201|OSN|60014-8|LNC|ACTH|ACTH
C2966814|T201|MTH_LN|60014-8|LNC|ACTH|ACTH
C2966814|T201|LC|60014-8|LNC|ACTH|ACTH
C2966814|T201|LN|60014-8|LNC|corticotropin|corticotropin
C2966814|T201|OSN|60014-8|LNC|corticotropin|corticotropin
C2966814|T201|MTH_LN|60014-8|LNC|corticotropin|corticotropin
C2966814|T201|LC|60014-8|LNC|corticotropin|corticotropin
C2966814|T201|LN|60014-8|LNC|adrenocorticotropin|adrenocorticotropin
C2966814|T201|OSN|60014-8|LNC|adrenocorticotropin|adrenocorticotropin
C2966814|T201|MTH_LN|60014-8|LNC|adrenocorticotropin|adrenocorticotropin
C2966814|T201|LC|60014-8|LNC|adrenocorticotropin|adrenocorticotropin
C2966815|T201|LN|60015-5|LNC|ACTH|ACTH
C2966815|T201|LC|60015-5|LNC|ACTH|ACTH
C2966815|T201|MTH_LN|60015-5|LNC|ACTH|ACTH
C2966815|T201|OSN|60015-5|LNC|ACTH|ACTH
C2966815|T201|LN|60015-5|LNC|corticotropin|corticotropin
C2966815|T201|LC|60015-5|LNC|corticotropin|corticotropin
C2966815|T201|MTH_LN|60015-5|LNC|corticotropin|corticotropin
C2966815|T201|OSN|60015-5|LNC|corticotropin|corticotropin
C2966815|T201|LN|60015-5|LNC|adrenocorticotropin|adrenocorticotropin
C2966815|T201|LC|60015-5|LNC|adrenocorticotropin|adrenocorticotropin
C2966815|T201|MTH_LN|60015-5|LNC|adrenocorticotropin|adrenocorticotropin
C2966815|T201|OSN|60015-5|LNC|adrenocorticotropin|adrenocorticotropin
C2966816|T201|LN|60016-3|LNC|ACTH|ACTH
C2966816|T201|LC|60016-3|LNC|ACTH|ACTH
C2966816|T201|MTH_LN|60016-3|LNC|ACTH|ACTH
C2966816|T201|OSN|60016-3|LNC|ACTH|ACTH
C2966816|T201|LN|60016-3|LNC|corticotropin|corticotropin
C2966816|T201|LC|60016-3|LNC|corticotropin|corticotropin
C2966816|T201|MTH_LN|60016-3|LNC|corticotropin|corticotropin
C2966816|T201|OSN|60016-3|LNC|corticotropin|corticotropin
C2966816|T201|LN|60016-3|LNC|adrenocorticotropin|adrenocorticotropin
C2966816|T201|LC|60016-3|LNC|adrenocorticotropin|adrenocorticotropin
C2966816|T201|MTH_LN|60016-3|LNC|adrenocorticotropin|adrenocorticotropin
C2966816|T201|OSN|60016-3|LNC|adrenocorticotropin|adrenocorticotropin
C2969748|T201|LN|59849-0|LNC|lactate|lactate
C2969748|T201|OSN|59849-0|LNC|lactate|lactate
C2969748|T201|MTH_LN|59849-0|LNC|lactate|lactate
C2969748|T201|LC|59849-0|LNC|lactate|lactate
C2969770|T201|LN|60025-4|LNC|urobilinogen|urobilinogen
C2969770|T201|MTH_LN|60025-4|LNC|urobilinogen|urobilinogen
C2969770|T201|LC|60025-4|LNC|urobilinogen|urobilinogen
C2969770|T201|OSN|60025-4|LNC|urobilinogen|urobilinogen
C2969825|T201|LN|59891-2|LNC|xenobiotic|xenobiotic
C2969825|T201|OSN|59891-2|LNC|xenobiotic|xenobiotic
C2969825|T201|LC|59891-2|LNC|xenobiotic|xenobiotic
C2969825|T201|MTH_LN|59891-2|LNC|xenobiotic|xenobiotic
C2969934|T201|LN|60017-1|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C2969934|T201|OSN|60017-1|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C2969934|T201|MTH_LN|60017-1|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C2969934|T201|LC|60017-1|LNC|lactate dehydrogenase activity|lactate dehydrogenase activity
C2969949|T201|LN|60048-6|LNC|xenobiotic|xenobiotic
C2969949|T201|OSN|60048-6|LNC|xenobiotic|xenobiotic
C2969949|T201|MTH_LN|60048-6|LNC|xenobiotic|xenobiotic
C2969949|T201|LC|60048-6|LNC|xenobiotic|xenobiotic
C2970267|T201|LN|60474-4|LNC|reticulocytes|reticulocytes
C2970267|T201|LC|60474-4|LNC|reticulocytes|reticulocytes
C2970267|T201|MTH_LN|60474-4|LNC|reticulocytes|reticulocytes
C2970267|T201|OSN|60474-4|LNC|reticulocytes|reticulocytes
C2970267|T201|LN|60474-4|LNC|reticulocyte count|reticulocyte count
C2970267|T201|LC|60474-4|LNC|reticulocyte count|reticulocyte count
C2970267|T201|MTH_LN|60474-4|LNC|reticulocyte count|reticulocyte count
C2970267|T201|OSN|60474-4|LNC|reticulocyte count|reticulocyte count
C2970588|T201|LN|61128-5|LNC|xenobiotic|xenobiotic
C2970588|T201|MTH_LN|61128-5|LNC|xenobiotic|xenobiotic
C2970588|T201|OSN|61128-5|LNC|xenobiotic|xenobiotic
C2970588|T201|LC|61128-5|LNC|xenobiotic|xenobiotic
C2973163|T201|LN|62241-5|LNC|hematocrit|hematocrit
C2973163|T201|MTH_LN|62241-5|LNC|hematocrit|hematocrit
C2973163|T201|OSN|62241-5|LNC|hematocrit|hematocrit
C2973163|T201|LC|62241-5|LNC|hematocrit|hematocrit
C2973199|T201|LN|62290-2|LNC|vitamin D metabolism|vitamin D metabolism
C2973199|T201|OSN|62290-2|LNC|vitamin D metabolism|vitamin D metabolism
C2973199|T201|LC|62290-2|LNC|vitamin D metabolism|vitamin D metabolism
C2973199|T201|MTH_LN|62290-2|LNC|vitamin D metabolism|vitamin D metabolism
C2973199|T201|LN|62290-2|LNC|calcitriol|calcitriol
C2973199|T201|OSN|62290-2|LNC|calcitriol|calcitriol
C2973199|T201|LC|62290-2|LNC|calcitriol|calcitriol
C2973199|T201|MTH_LN|62290-2|LNC|calcitriol|calcitriol
C2973199|T201|LN|62290-2|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C2973199|T201|OSN|62290-2|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C2973199|T201|LC|62290-2|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C2973199|T201|MTH_LN|62290-2|LNC|1,25-dihydroxyvitamin D3|1,25-dihydroxyvitamin D3
C2973199|T201|LN|62290-2|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C2973199|T201|OSN|62290-2|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C2973199|T201|LC|62290-2|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C2973199|T201|MTH_LN|62290-2|LNC|1,25-dihydroxycholecalciferol|1,25-dihydroxycholecalciferol
C3166946|T201|LN|57645-4|LNC|C-peptide|C-peptide
C3166946|T201|LC|57645-4|LNC|C-peptide|C-peptide
C3166946|T201|MTH_LN|57645-4|LNC|C-peptide|C-peptide
C3166946|T201|OSN|57645-4|LNC|C-peptide|C-peptide
C3166946|T201|LN|57645-4|LNC|C peptide|C peptide
C3166946|T201|LC|57645-4|LNC|C peptide|C peptide
C3166946|T201|MTH_LN|57645-4|LNC|C peptide|C peptide
C3166946|T201|OSN|57645-4|LNC|C peptide|C peptide
C3167213|T201|LN|57648-8|LNC|C-peptide|C-peptide
C3167213|T201|MTH_LN|57648-8|LNC|C-peptide|C-peptide
C3167213|T201|OSN|57648-8|LNC|C-peptide|C-peptide
C3167213|T201|LC|57648-8|LNC|C-peptide|C-peptide
C3167213|T201|LN|57648-8|LNC|C peptide|C peptide
C3167213|T201|MTH_LN|57648-8|LNC|C peptide|C peptide
C3167213|T201|OSN|57648-8|LNC|C peptide|C peptide
C3167213|T201|LC|57648-8|LNC|C peptide|C peptide
C3167214|T201|LN|57649-6|LNC|C-peptide|C-peptide
C3167214|T201|LC|57649-6|LNC|C-peptide|C-peptide
C3167214|T201|MTH_LN|57649-6|LNC|C-peptide|C-peptide
C3167214|T201|OSN|57649-6|LNC|C-peptide|C-peptide
C3167214|T201|LN|57649-6|LNC|C peptide|C peptide
C3167214|T201|LC|57649-6|LNC|C peptide|C peptide
C3167214|T201|MTH_LN|57649-6|LNC|C peptide|C peptide
C3167214|T201|OSN|57649-6|LNC|C peptide|C peptide
C3167215|T201|LN|57650-4|LNC|C-peptide|C-peptide
C3167215|T201|LC|57650-4|LNC|C-peptide|C-peptide
C3167215|T201|MTH_LN|57650-4|LNC|C-peptide|C-peptide
C3167215|T201|OSN|57650-4|LNC|C-peptide|C-peptide
C3167215|T201|LN|57650-4|LNC|C peptide|C peptide
C3167215|T201|LC|57650-4|LNC|C peptide|C peptide
C3167215|T201|MTH_LN|57650-4|LNC|C peptide|C peptide
C3167215|T201|OSN|57650-4|LNC|C peptide|C peptide
C3169574|T201|LN|62487-4|LNC|urobilinogen|urobilinogen
C3169574|T201|OSN|62487-4|LNC|urobilinogen|urobilinogen
C3169574|T201|LC|62487-4|LNC|urobilinogen|urobilinogen
C3169574|T201|MTH_LN|62487-4|LNC|urobilinogen|urobilinogen
C3172328|T201|LN|63243-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172328|T201|LC|63243-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172328|T201|OSN|63243-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172328|T201|MTH_LN|63243-0|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172329|T201|LN|63244-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172329|T201|LC|63244-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172329|T201|MTH_LN|63244-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172329|T201|OSN|63244-8|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172332|T201|LN|63247-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172332|T201|LC|63247-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172332|T201|MTH_LN|63247-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172332|T201|OSN|63247-1|LNC|Anti-ganglioside GM1 IgM antibody|Anti-ganglioside GM1 IgM antibody
C3172373|T201|LN|63283-6|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C3172373|T201|LC|63283-6|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C3172373|T201|OSN|63283-6|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C3172373|T201|MTH_LN|63283-6|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C3172428|T201|LN|63359-4|LNC|Autoimmune antibody|Autoimmune antibody
C3172428|T201|LC|63359-4|LNC|Autoimmune antibody|Autoimmune antibody
C3172428|T201|MTH_LN|63359-4|LNC|Autoimmune antibody|Autoimmune antibody
C3172428|T201|OSN|63359-4|LNC|Autoimmune antibody|Autoimmune antibody
C3172429|T201|LN|63360-2|LNC|Autoimmune antibody|Autoimmune antibody
C3172429|T201|MTH_LN|63360-2|LNC|Autoimmune antibody|Autoimmune antibody
C3172429|T201|LC|63360-2|LNC|Autoimmune antibody|Autoimmune antibody
C3172429|T201|OSN|63360-2|LNC|Autoimmune antibody|Autoimmune antibody
C3172449|T201|LN|63378-4|LNC|y|y
C3172449|T201|OSN|63378-4|LNC|y|y
C3172449|T201|LC|63378-4|LNC|y|y
C3172449|T201|MTH_LN|63378-4|LNC|y|y
C3172620|T201|LN|63554-0|LNC|neutrophil count|neutrophil count
C3172620|T201|MTH_LN|63554-0|LNC|neutrophil count|neutrophil count
C3172620|T201|OSN|63554-0|LNC|neutrophil count|neutrophil count
C3172620|T201|LC|63554-0|LNC|neutrophil count|neutrophil count
C3172620|T201|LN|63554-0|LNC|cytology|cytology
C3172620|T201|MTH_LN|63554-0|LNC|cytology|cytology
C3172620|T201|OSN|63554-0|LNC|cytology|cytology
C3172620|T201|LC|63554-0|LNC|cytology|cytology
C3258901|T201|LN|66126-4|LNC|VLDL cholesterol|VLDL cholesterol
C3258901|T201|OSN|66126-4|LNC|VLDL cholesterol|VLDL cholesterol
C3258901|T201|LC|66126-4|LNC|VLDL cholesterol|VLDL cholesterol
C3258901|T201|MTH_LN|66126-4|LNC|VLDL cholesterol|VLDL cholesterol
C3258901|T201|LN|66126-4|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3258901|T201|OSN|66126-4|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3258901|T201|LC|66126-4|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3258901|T201|MTH_LN|66126-4|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3258901|T201|LN|66126-4|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3258901|T201|OSN|66126-4|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3258901|T201|LC|66126-4|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3258901|T201|MTH_LN|66126-4|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3258971|T201|LN|66139-7|LNC|neutrophil counts|neutrophil counts
C3258971|T201|LC|66139-7|LNC|neutrophil counts|neutrophil counts
C3258971|T201|OSN|66139-7|LNC|neutrophil counts|neutrophil counts
C3258971|T201|MTH_LN|66139-7|LNC|neutrophil counts|neutrophil counts
C3258971|T201|LN|66139-7|LNC|neutrophil count|neutrophil count
C3258971|T201|LC|66139-7|LNC|neutrophil count|neutrophil count
C3258971|T201|OSN|66139-7|LNC|neutrophil count|neutrophil count
C3258971|T201|MTH_LN|66139-7|LNC|neutrophil count|neutrophil count
C3258971|T201|LN|66139-7|LNC|neutrophil|neutrophil
C3258971|T201|LC|66139-7|LNC|neutrophil|neutrophil
C3258971|T201|OSN|66139-7|LNC|neutrophil|neutrophil
C3258971|T201|MTH_LN|66139-7|LNC|neutrophil|neutrophil
C3259342|T201|LN|67151-1|LNC|troponin T|troponin T
C3259342|T201|OSN|67151-1|LNC|troponin T|troponin T
C3259342|T201|MTH_LN|67151-1|LNC|troponin T|troponin T
C3259342|T201|LC|67151-1|LNC|troponin T|troponin T
C3259432|T201|LN|66499-5|LNC|VLDL cholesterol|VLDL cholesterol
C3259432|T201|OSN|66499-5|LNC|VLDL cholesterol|VLDL cholesterol
C3259432|T201|LC|66499-5|LNC|VLDL cholesterol|VLDL cholesterol
C3259432|T201|MTH_LN|66499-5|LNC|VLDL cholesterol|VLDL cholesterol
C3259432|T201|LN|66499-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3259432|T201|OSN|66499-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3259432|T201|LC|66499-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3259432|T201|MTH_LN|66499-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3259432|T201|LN|66499-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3259432|T201|OSN|66499-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3259432|T201|LC|66499-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3259432|T201|MTH_LN|66499-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3259749|T201|LC|66732-9|LNC|ACTH|ACTH
C3259749|T201|MTH_LN|66732-9|LNC|ACTH|ACTH
C3259749|T201|OSN|66732-9|LNC|ACTH|ACTH
C3259749|T201|LN|66732-9|LNC|ACTH|ACTH
C3259749|T201|LC|66732-9|LNC|corticotropin|corticotropin
C3259749|T201|MTH_LN|66732-9|LNC|corticotropin|corticotropin
C3259749|T201|OSN|66732-9|LNC|corticotropin|corticotropin
C3259749|T201|LN|66732-9|LNC|corticotropin|corticotropin
C3259749|T201|LC|66732-9|LNC|adrenocorticotropin|adrenocorticotropin
C3259749|T201|MTH_LN|66732-9|LNC|adrenocorticotropin|adrenocorticotropin
C3259749|T201|OSN|66732-9|LNC|adrenocorticotropin|adrenocorticotropin
C3259749|T201|LN|66732-9|LNC|adrenocorticotropin|adrenocorticotropin
C3262207|T201|LN|68324-3|LNC|von Willebrand factor|von Willebrand factor
C3262207|T201|OSN|68324-3|LNC|von Willebrand factor|von Willebrand factor
C3262207|T201|MTH_LN|68324-3|LNC|von Willebrand factor|von Willebrand factor
C3262207|T201|LC|68324-3|LNC|von Willebrand factor|von Willebrand factor
C3262207|T201|LN|68324-3|LNC|von Willebrand factor activity|von Willebrand factor activity
C3262207|T201|OSN|68324-3|LNC|von Willebrand factor activity|von Willebrand factor activity
C3262207|T201|MTH_LN|68324-3|LNC|von Willebrand factor activity|von Willebrand factor activity
C3262207|T201|LC|68324-3|LNC|von Willebrand factor activity|von Willebrand factor activity
// C3262756|T201|LN|68902-6|LNC||
// C3262756|T201|OSN|68902-6|LNC||
// C3262756|T201|MTH_LN|68902-6|LNC||
// C3262756|T201|LC|68902-6|LNC||
C3262756|T201|LN|68902-6|LNC|occult|occult
C3262756|T201|OSN|68902-6|LNC|occult|occult
C3262756|T201|MTH_LN|68902-6|LNC|occult|occult
C3262756|T201|LC|68902-6|LNC|occult|occult
// C3262757|T201|LN|68903-4|LNC||
// C3262757|T201|OSN|68903-4|LNC||
// C3262757|T201|MTH_LN|68903-4|LNC||
// C3262757|T201|LC|68903-4|LNC||
C3262757|T201|LN|68903-4|LNC|occult|occult
C3262757|T201|OSN|68903-4|LNC|occult|occult
C3262757|T201|MTH_LN|68903-4|LNC|occult|occult
C3262757|T201|LC|68903-4|LNC|occult|occult
C3262759|T201|LN|68911-7|LNC|lactate|lactate
C3262759|T201|MTH_LN|68911-7|LNC|lactate|lactate
C3262759|T201|OSN|68911-7|LNC|lactate|lactate
C3262759|T201|LC|68911-7|LNC|lactate|lactate
C3262763|T201|LN|68916-6|LNC|Autoimmune antibody|Autoimmune antibody
C3262763|T201|MTH_LN|68916-6|LNC|Autoimmune antibody|Autoimmune antibody
C3262763|T201|OSN|68916-6|LNC|Autoimmune antibody|Autoimmune antibody
C3262763|T201|LC|68916-6|LNC|Autoimmune antibody|Autoimmune antibody
C3262782|T201|LN|68937-2|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C3262782|T201|LC|68937-2|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C3262782|T201|MTH_LN|68937-2|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C3262782|T201|OSN|68937-2|LNC|Acetylcholine receptor antibody|Acetylcholine receptor antibody
C3262796|T201|LN|68955-4|LNC|ketone bodies|ketone bodies
C3262796|T201|OSN|68955-4|LNC|ketone bodies|ketone bodies
C3262796|T201|LC|68955-4|LNC|ketone bodies|ketone bodies
C3262796|T201|MTH_LN|68955-4|LNC|ketone bodies|ketone bodies
C3481648|T201|LN|70198-7|LNC|xenobiotic|xenobiotic
C3481648|T201|MTH_LN|70198-7|LNC|xenobiotic|xenobiotic
C3481648|T201|LC|70198-7|LNC|xenobiotic|xenobiotic
C3481648|T201|OSN|70198-7|LNC|xenobiotic|xenobiotic
C3481653|T201|LN|70203-5|LNC|VLDL cholesterol|VLDL cholesterol
C3481653|T201|MTH_LN|70203-5|LNC|VLDL cholesterol|VLDL cholesterol
C3481653|T201|LC|70203-5|LNC|VLDL cholesterol|VLDL cholesterol
C3481653|T201|OSN|70203-5|LNC|VLDL cholesterol|VLDL cholesterol
C3481653|T201|LN|70203-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3481653|T201|MTH_LN|70203-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3481653|T201|LC|70203-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3481653|T201|OSN|70203-5|LNC|very-low-density lipoprotein cholesterol|very-low-density lipoprotein cholesterol
C3481653|T201|LN|70203-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3481653|T201|MTH_LN|70203-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3481653|T201|LC|70203-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3481653|T201|OSN|70203-5|LNC|very-low-density lipoprotein|very-low-density lipoprotein
C3481704|T201|LN|69419-0|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C3481704|T201|MTH_LN|69419-0|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C3481704|T201|OSN|69419-0|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C3481704|T201|LC|69419-0|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C3481704|T201|LN|69419-0|LNC|LDL|LDL
C3481704|T201|MTH_LN|69419-0|LNC|LDL|LDL
C3481704|T201|OSN|69419-0|LNC|LDL|LDL
C3481704|T201|LC|69419-0|LNC|LDL|LDL
C3481704|T201|LN|69419-0|LNC|LDL cholesterol|LDL cholesterol
C3481704|T201|MTH_LN|69419-0|LNC|LDL cholesterol|LDL cholesterol
C3481704|T201|OSN|69419-0|LNC|LDL cholesterol|LDL cholesterol
C3481704|T201|LC|69419-0|LNC|LDL cholesterol|LDL cholesterol
C3481704|T201|LN|69419-0|LNC|low-density lipoprotein|low-density lipoprotein
C3481704|T201|MTH_LN|69419-0|LNC|low-density lipoprotein|low-density lipoprotein
C3481704|T201|OSN|69419-0|LNC|low-density lipoprotein|low-density lipoprotein
C3481704|T201|LC|69419-0|LNC|low-density lipoprotein|low-density lipoprotein
C3481704|T201|LN|69419-0|LNC|beta-lipoproteins|beta-lipoproteins
C3481704|T201|MTH_LN|69419-0|LNC|beta-lipoproteins|beta-lipoproteins
C3481704|T201|OSN|69419-0|LNC|beta-lipoproteins|beta-lipoproteins
C3481704|T201|LC|69419-0|LNC|beta-lipoproteins|beta-lipoproteins
C3481704|T201|LN|69419-0|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C3481704|T201|MTH_LN|69419-0|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C3481704|T201|OSN|69419-0|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C3481704|T201|LC|69419-0|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C3481704|T201|LN|69419-0|LNC|LDL-C|LDL-C
C3481704|T201|MTH_LN|69419-0|LNC|LDL-C|LDL-C
C3481704|T201|OSN|69419-0|LNC|LDL-C|LDL-C
C3481704|T201|LC|69419-0|LNC|LDL-C|LDL-C
C3482218|T201|LN|70149-0|LNC|methadone test|methadone test
C3482218|T201|LC|70149-0|LNC|methadone test|methadone test
C3482218|T201|OSN|70149-0|LNC|methadone test|methadone test
C3482218|T201|MTH_LN|70149-0|LNC|methadone test|methadone test
C3482237|T201|LN|70168-0|LNC|hematocrit|hematocrit
C3482237|T201|OSN|70168-0|LNC|hematocrit|hematocrit
C3482237|T201|LC|70168-0|LNC|hematocrit|hematocrit
C3482237|T201|MTH_LN|70168-0|LNC|hematocrit|hematocrit
C3482238|T201|LN|70169-8|LNC|hematocrit|hematocrit
C3482238|T201|LC|70169-8|LNC|hematocrit|hematocrit
C3482238|T201|OSN|70169-8|LNC|hematocrit|hematocrit
C3482238|T201|MTH_LN|70169-8|LNC|hematocrit|hematocrit
C3483886|T201|LN|71847-8|LNC|oxygen|oxygen
C3483886|T201|LC|71847-8|LNC|oxygen|oxygen
C3483886|T201|MTH_LN|71847-8|LNC|oxygen|oxygen
C3483886|T201|OSN|71847-8|LNC|oxygen|oxygen
C3484058|T201|LN|71828-8|LNC|hematocrit|hematocrit
C3484058|T201|MTH_LN|71828-8|LNC|hematocrit|hematocrit
C3484058|T201|OSN|71828-8|LNC|hematocrit|hematocrit
C3484058|T201|LC|71828-8|LNC|hematocrit|hematocrit
C3484059|T201|LN|71829-6|LNC|hematocrit|hematocrit
C3484059|T201|LC|71829-6|LNC|hematocrit|hematocrit
C3484059|T201|MTH_LN|71829-6|LNC|hematocrit|hematocrit
C3484059|T201|OSN|71829-6|LNC|hematocrit|hematocrit
C3484060|T201|LN|71830-4|LNC|hematocrit|hematocrit
C3484060|T201|MTH_LN|71830-4|LNC|hematocrit|hematocrit
C3484060|T201|OSN|71830-4|LNC|hematocrit|hematocrit
C3484060|T201|LC|71830-4|LNC|hematocrit|hematocrit
C3484061|T201|LN|71831-2|LNC|hematocrit|hematocrit
C3484061|T201|MTH_LN|71831-2|LNC|hematocrit|hematocrit
C3484061|T201|OSN|71831-2|LNC|hematocrit|hematocrit
C3484061|T201|LC|71831-2|LNC|hematocrit|hematocrit
C3484062|T201|LN|71832-0|LNC|hematocrit|hematocrit
C3484062|T201|OSN|71832-0|LNC|hematocrit|hematocrit
C3484062|T201|MTH_LN|71832-0|LNC|hematocrit|hematocrit
C3484062|T201|LC|71832-0|LNC|hematocrit|hematocrit
C3484063|T201|LN|71833-8|LNC|hematocrit|hematocrit
C3484063|T201|OSN|71833-8|LNC|hematocrit|hematocrit
C3484063|T201|LC|71833-8|LNC|hematocrit|hematocrit
C3484063|T201|MTH_LN|71833-8|LNC|hematocrit|hematocrit
C3533399|T201|LN|72786-7|LNC|cotinine|cotinine
C3533399|T201|MTH_LN|72786-7|LNC|cotinine|cotinine
C3533399|T201|OSN|72786-7|LNC|cotinine|cotinine
C3533399|T201|LC|72786-7|LNC|cotinine|cotinine
C3654079|T201|LN|73978-9|LNC|von Willebrand factor|von Willebrand factor
C3654079|T201|MTH_LN|73978-9|LNC|von Willebrand factor|von Willebrand factor
C3654079|T201|LC|73978-9|LNC|von Willebrand factor|von Willebrand factor
C3654079|T201|OSN|73978-9|LNC|von Willebrand factor|von Willebrand factor
C3654079|T201|LN|73978-9|LNC|von Willebrand factor activity|von Willebrand factor activity
C3654079|T201|MTH_LN|73978-9|LNC|von Willebrand factor activity|von Willebrand factor activity
C3654079|T201|LC|73978-9|LNC|von Willebrand factor activity|von Willebrand factor activity
C3654079|T201|OSN|73978-9|LNC|von Willebrand factor activity|von Willebrand factor activity
C3654405|T201|LN|73572-0|LNC|magnesium|magnesium
C3654405|T201|LC|73572-0|LNC|magnesium|magnesium
C3654405|T201|MTH_LN|73572-0|LNC|magnesium|magnesium
C3654405|T201|OSN|73572-0|LNC|magnesium|magnesium
C3654405|T201|LN|73572-0|LNC|magnesium metabolism|magnesium metabolism
C3654405|T201|LC|73572-0|LNC|magnesium metabolism|magnesium metabolism
C3654405|T201|MTH_LN|73572-0|LNC|magnesium metabolism|magnesium metabolism
C3654405|T201|OSN|73572-0|LNC|magnesium metabolism|magnesium metabolism
C3654405|T201|LN|73572-0|LNC|magnesium homeostasis|magnesium homeostasis
C3654405|T201|LC|73572-0|LNC|magnesium homeostasis|magnesium homeostasis
C3654405|T201|MTH_LN|73572-0|LNC|magnesium homeostasis|magnesium homeostasis
C3654405|T201|OSN|73572-0|LNC|magnesium homeostasis|magnesium homeostasis
C3655182|T201|LN|70148-2|LNC|methadone test|methadone test
C3655182|T201|OSN|70148-2|LNC|methadone test|methadone test
C3655182|T201|LC|70148-2|LNC|methadone test|methadone test
C3655182|T201|MTH_LN|70148-2|LNC|methadone test|methadone test
C3655183|T201|LN|70147-4|LNC|methadone test|methadone test
C3655183|T201|LC|70147-4|LNC|methadone test|methadone test
C3655183|T201|MTH_LN|70147-4|LNC|methadone test|methadone test
C3655183|T201|OSN|70147-4|LNC|methadone test|methadone test
C3699844|T201|LN|74398-9|LNC|neutrophil counts|neutrophil counts
C3699844|T201|LC|74398-9|LNC|neutrophil counts|neutrophil counts
C3699844|T201|MTH_LN|74398-9|LNC|neutrophil counts|neutrophil counts
C3699844|T201|OSN|74398-9|LNC|neutrophil counts|neutrophil counts
C3699844|T201|LN|74398-9|LNC|neutrophil count|neutrophil count
C3699844|T201|LC|74398-9|LNC|neutrophil count|neutrophil count
C3699844|T201|MTH_LN|74398-9|LNC|neutrophil count|neutrophil count
C3699844|T201|OSN|74398-9|LNC|neutrophil count|neutrophil count
C3699844|T201|LN|74398-9|LNC|neutrophil|neutrophil
C3699844|T201|LC|74398-9|LNC|neutrophil|neutrophil
C3699844|T201|MTH_LN|74398-9|LNC|neutrophil|neutrophil
C3699844|T201|OSN|74398-9|LNC|neutrophil|neutrophil
C3699850|T201|LN|74404-5|LNC|eosinophil count|eosinophil count
C3699850|T201|MTH_LN|74404-5|LNC|eosinophil count|eosinophil count
C3699850|T201|LC|74404-5|LNC|eosinophil count|eosinophil count
C3699850|T201|OSN|74404-5|LNC|eosinophil count|eosinophil count
C3699850|T201|LN|74404-5|LNC|eosinophil morphology|eosinophil morphology
C3699850|T201|MTH_LN|74404-5|LNC|eosinophil morphology|eosinophil morphology
C3699850|T201|LC|74404-5|LNC|eosinophil morphology|eosinophil morphology
C3699850|T201|OSN|74404-5|LNC|eosinophil morphology|eosinophil morphology
C3699850|T201|LN|74404-5|LNC|eosinophils|eosinophils
C3699850|T201|MTH_LN|74404-5|LNC|eosinophils|eosinophils
C3699850|T201|LC|74404-5|LNC|eosinophils|eosinophils
C3699850|T201|OSN|74404-5|LNC|eosinophils|eosinophils
C3699851|T201|LN|74405-2|LNC|eosinophil count|eosinophil count
C3699851|T201|MTH_LN|74405-2|LNC|eosinophil count|eosinophil count
C3699851|T201|LC|74405-2|LNC|eosinophil count|eosinophil count
C3699851|T201|OSN|74405-2|LNC|eosinophil count|eosinophil count
C3699851|T201|LN|74405-2|LNC|eosinophil morphology|eosinophil morphology
C3699851|T201|MTH_LN|74405-2|LNC|eosinophil morphology|eosinophil morphology
C3699851|T201|LC|74405-2|LNC|eosinophil morphology|eosinophil morphology
C3699851|T201|OSN|74405-2|LNC|eosinophil morphology|eosinophil morphology
C3699851|T201|LN|74405-2|LNC|eosinophils|eosinophils
C3699851|T201|MTH_LN|74405-2|LNC|eosinophils|eosinophils
C3699851|T201|LC|74405-2|LNC|eosinophils|eosinophils
C3699851|T201|OSN|74405-2|LNC|eosinophils|eosinophils
C3846945|T201|LN|75040-6|LNC|CSF lactate|CSF lactate
C3846945|T201|LC|75040-6|LNC|CSF lactate|CSF lactate
C3846945|T201|OSN|75040-6|LNC|CSF lactate|CSF lactate
C3846945|T201|MTH_LN|75040-6|LNC|CSF lactate|CSF lactate
C3846945|T201|LN|75040-6|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C3846945|T201|LC|75040-6|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C3846945|T201|OSN|75040-6|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C3846945|T201|MTH_LN|75040-6|LNC|cerebrospinal fluid lactate|cerebrospinal fluid lactate
C3846945|T201|LN|75040-6|LNC|CSF lactic acid|CSF lactic acid
C3846945|T201|LC|75040-6|LNC|CSF lactic acid|CSF lactic acid
C3846945|T201|OSN|75040-6|LNC|CSF lactic acid|CSF lactic acid
C3846945|T201|MTH_LN|75040-6|LNC|CSF lactic acid|CSF lactic acid
C3847065|T201|LN|74893-9|LNC|D-mannose|D-mannose
C3847065|T201|OSN|74893-9|LNC|D-mannose|D-mannose
C3847065|T201|LC|74893-9|LNC|D-mannose|D-mannose
C3847065|T201|MTH_LN|74893-9|LNC|D-mannose|D-mannose
C3847419|T201|LN|74809-5|LNC|von Willebrand factor|von Willebrand factor
C3847419|T201|OSN|74809-5|LNC|von Willebrand factor|von Willebrand factor
C3847419|T201|MTH_LN|74809-5|LNC|von Willebrand factor|von Willebrand factor
C3847419|T201|LC|74809-5|LNC|von Willebrand factor|von Willebrand factor
C3847419|T201|LN|74809-5|LNC|von Willebrand factor activity|von Willebrand factor activity
C3847419|T201|OSN|74809-5|LNC|von Willebrand factor activity|von Willebrand factor activity
C3847419|T201|MTH_LN|74809-5|LNC|von Willebrand factor activity|von Willebrand factor activity
C3847419|T201|LC|74809-5|LNC|von Willebrand factor activity|von Willebrand factor activity
C3847420|T201|LN|74808-7|LNC|von Willebrand factor|von Willebrand factor
C3847420|T201|LC|74808-7|LNC|von Willebrand factor|von Willebrand factor
C3847420|T201|OSN|74808-7|LNC|von Willebrand factor|von Willebrand factor
C3847420|T201|MTH_LN|74808-7|LNC|von Willebrand factor|von Willebrand factor
C3847420|T201|LN|74808-7|LNC|von Willebrand factor activity|von Willebrand factor activity
C3847420|T201|LC|74808-7|LNC|von Willebrand factor activity|von Willebrand factor activity
C3847420|T201|OSN|74808-7|LNC|von Willebrand factor activity|von Willebrand factor activity
C3847420|T201|MTH_LN|74808-7|LNC|von Willebrand factor activity|von Willebrand factor activity
C3870010|T201|LN|75913-4|LNC|Autoimmune antibody|Autoimmune antibody
C3870010|T201|LC|75913-4|LNC|Autoimmune antibody|Autoimmune antibody
C3870010|T201|MTH_LN|75913-4|LNC|Autoimmune antibody|Autoimmune antibody
C3870010|T201|OSN|75913-4|LNC|Autoimmune antibody|Autoimmune antibody
C3870037|T201|LN|75883-9|LNC|Autoimmune antibody|Autoimmune antibody
C3870037|T201|OSN|75883-9|LNC|Autoimmune antibody|Autoimmune antibody
C3870037|T201|LC|75883-9|LNC|Autoimmune antibody|Autoimmune antibody
C3870037|T201|MTH_LN|75883-9|LNC|Autoimmune antibody|Autoimmune antibody
C3870342|T201|LN|75511-6|LNC|Autoimmune antibody|Autoimmune antibody
C3870342|T201|MTH_LN|75511-6|LNC|Autoimmune antibody|Autoimmune antibody
C3870342|T201|LC|75511-6|LNC|Autoimmune antibody|Autoimmune antibody
C3870342|T201|OSN|75511-6|LNC|Autoimmune antibody|Autoimmune antibody
C3870449|T201|LN|75366-5|LNC|lactate|lactate
C3870449|T201|OSN|75366-5|LNC|lactate|lactate
C3870449|T201|LC|75366-5|LNC|lactate|lactate
C3870449|T201|MTH_LN|75366-5|LNC|lactate|lactate
C4036476|T201|LN|76483-7|LNC|apolipoprotein AI|apolipoprotein AI
C4036476|T201|MTH_LN|76483-7|LNC|apolipoprotein AI|apolipoprotein AI
C4036476|T201|OSN|76483-7|LNC|apolipoprotein AI|apolipoprotein AI
C4036476|T201|LC|76483-7|LNC|apolipoprotein AI|apolipoprotein AI
C4036476|T201|LN|76483-7|LNC|apoA-I|apoA-I
C4036476|T201|MTH_LN|76483-7|LNC|apoA-I|apoA-I
C4036476|T201|OSN|76483-7|LNC|apoA-I|apoA-I
C4036476|T201|LC|76483-7|LNC|apoA-I|apoA-I
C4036476|T201|LN|76483-7|LNC|apo-AI|apo-AI
C4036476|T201|MTH_LN|76483-7|LNC|apo-AI|apo-AI
C4036476|T201|OSN|76483-7|LNC|apo-AI|apo-AI
C4036476|T201|LC|76483-7|LNC|apo-AI|apo-AI
C4036527|T201|LN|77939-7|LNC|ACTH|ACTH
C4036527|T201|MTH_LN|77939-7|LNC|ACTH|ACTH
C4036527|T201|OSN|77939-7|LNC|ACTH|ACTH
C4036527|T201|LC|77939-7|LNC|ACTH|ACTH
C4036527|T201|LN|77939-7|LNC|corticotropin|corticotropin
C4036527|T201|MTH_LN|77939-7|LNC|corticotropin|corticotropin
C4036527|T201|OSN|77939-7|LNC|corticotropin|corticotropin
C4036527|T201|LC|77939-7|LNC|corticotropin|corticotropin
C4036527|T201|LN|77939-7|LNC|adrenocorticotropin|adrenocorticotropin
C4036527|T201|MTH_LN|77939-7|LNC|adrenocorticotropin|adrenocorticotropin
C4036527|T201|OSN|77939-7|LNC|adrenocorticotropin|adrenocorticotropin
C4036527|T201|LC|77939-7|LNC|adrenocorticotropin|adrenocorticotropin
C4036769|T201|LN|77612-0|LNC|C-peptide|C-peptide
C4036769|T201|OSN|77612-0|LNC|C-peptide|C-peptide
C4036769|T201|MTH_LN|77612-0|LNC|C-peptide|C-peptide
C4036769|T201|LC|77612-0|LNC|C-peptide|C-peptide
C4036769|T201|LN|77612-0|LNC|C peptide|C peptide
C4036769|T201|OSN|77612-0|LNC|C peptide|C peptide
C4036769|T201|MTH_LN|77612-0|LNC|C peptide|C peptide
C4036769|T201|LC|77612-0|LNC|C peptide|C peptide
C4036770|T201|LN|77611-2|LNC|C-peptide|C-peptide
C4036770|T201|OSN|77611-2|LNC|C-peptide|C-peptide
C4036770|T201|LC|77611-2|LNC|C-peptide|C-peptide
C4036770|T201|MTH_LN|77611-2|LNC|C-peptide|C-peptide
C4036770|T201|LN|77611-2|LNC|C peptide|C peptide
C4036770|T201|OSN|77611-2|LNC|C peptide|C peptide
C4036770|T201|LC|77611-2|LNC|C peptide|C peptide
C4036770|T201|MTH_LN|77611-2|LNC|C peptide|C peptide
C4036771|T201|LN|77610-4|LNC|C-peptide|C-peptide
C4036771|T201|LC|77610-4|LNC|C-peptide|C-peptide
C4036771|T201|OSN|77610-4|LNC|C-peptide|C-peptide
C4036771|T201|MTH_LN|77610-4|LNC|C-peptide|C-peptide
C4036771|T201|LN|77610-4|LNC|C peptide|C peptide
C4036771|T201|LC|77610-4|LNC|C peptide|C peptide
C4036771|T201|OSN|77610-4|LNC|C peptide|C peptide
C4036771|T201|MTH_LN|77610-4|LNC|C peptide|C peptide
C4037465|T201|LN|77652-6|LNC|C-peptide|C-peptide
C4037465|T201|MTH_LN|77652-6|LNC|C-peptide|C-peptide
C4037465|T201|OSN|77652-6|LNC|C-peptide|C-peptide
C4037465|T201|LC|77652-6|LNC|C-peptide|C-peptide
C4037465|T201|LN|77652-6|LNC|C peptide|C peptide
C4037465|T201|MTH_LN|77652-6|LNC|C peptide|C peptide
C4037465|T201|OSN|77652-6|LNC|C peptide|C peptide
C4037465|T201|LC|77652-6|LNC|C peptide|C peptide
C4037466|T201|LN|77651-8|LNC|C-peptide|C-peptide
C4037466|T201|LC|77651-8|LNC|C-peptide|C-peptide
C4037466|T201|OSN|77651-8|LNC|C-peptide|C-peptide
C4037466|T201|MTH_LN|77651-8|LNC|C-peptide|C-peptide
C4037466|T201|LN|77651-8|LNC|C peptide|C peptide
C4037466|T201|LC|77651-8|LNC|C peptide|C peptide
C4037466|T201|OSN|77651-8|LNC|C peptide|C peptide
C4037466|T201|MTH_LN|77651-8|LNC|C peptide|C peptide
C4037566|T201|LN|76672-5|LNC|CSF glucose|CSF glucose
C4037566|T201|LC|76672-5|LNC|CSF glucose|CSF glucose
C4037566|T201|MTH_LN|76672-5|LNC|CSF glucose|CSF glucose
C4037566|T201|OSN|76672-5|LNC|CSF glucose|CSF glucose
C4037566|T201|LN|76672-5|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037566|T201|LC|76672-5|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037566|T201|MTH_LN|76672-5|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037566|T201|OSN|76672-5|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037567|T201|LN|76671-7|LNC|CSF glucose|CSF glucose
C4037567|T201|MTH_LN|76671-7|LNC|CSF glucose|CSF glucose
C4037567|T201|LC|76671-7|LNC|CSF glucose|CSF glucose
C4037567|T201|OSN|76671-7|LNC|CSF glucose|CSF glucose
C4037567|T201|LN|76671-7|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037567|T201|MTH_LN|76671-7|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037567|T201|LC|76671-7|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037567|T201|OSN|76671-7|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037568|T201|LN|76670-9|LNC|CSF glucose|CSF glucose
C4037568|T201|MTH_LN|76670-9|LNC|CSF glucose|CSF glucose
C4037568|T201|OSN|76670-9|LNC|CSF glucose|CSF glucose
C4037568|T201|LC|76670-9|LNC|CSF glucose|CSF glucose
C4037568|T201|LN|76670-9|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037568|T201|MTH_LN|76670-9|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037568|T201|OSN|76670-9|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037568|T201|LC|76670-9|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037569|T201|LN|76669-1|LNC|CSF glucose|CSF glucose
C4037569|T201|OSN|76669-1|LNC|CSF glucose|CSF glucose
C4037569|T201|LC|76669-1|LNC|CSF glucose|CSF glucose
C4037569|T201|MTH_LN|76669-1|LNC|CSF glucose|CSF glucose
C4037569|T201|LN|76669-1|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037569|T201|OSN|76669-1|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037569|T201|LC|76669-1|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037569|T201|MTH_LN|76669-1|LNC|glucose in cerebral spinal fluid|glucose in cerebral spinal fluid
C4037570|T201|LN|76668-3|LNC|CSF protein|CSF protein
C4037570|T201|LC|76668-3|LNC|CSF protein|CSF protein
C4037570|T201|MTH_LN|76668-3|LNC|CSF protein|CSF protein
C4037570|T201|OSN|76668-3|LNC|CSF protein|CSF protein
C4037570|T201|LN|76668-3|LNC|protein in csf|protein in csf
C4037570|T201|LC|76668-3|LNC|protein in csf|protein in csf
C4037570|T201|MTH_LN|76668-3|LNC|protein in csf|protein in csf
C4037570|T201|OSN|76668-3|LNC|protein in csf|protein in csf
C4037570|T201|LN|76668-3|LNC|Spinal fluid protein|Spinal fluid protein
C4037570|T201|LC|76668-3|LNC|Spinal fluid protein|Spinal fluid protein
C4037570|T201|MTH_LN|76668-3|LNC|Spinal fluid protein|Spinal fluid protein
C4037570|T201|OSN|76668-3|LNC|Spinal fluid protein|Spinal fluid protein
C4037570|T201|LN|76668-3|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037570|T201|LC|76668-3|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037570|T201|MTH_LN|76668-3|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037570|T201|OSN|76668-3|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037570|T201|LN|76668-3|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037570|T201|LC|76668-3|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037570|T201|MTH_LN|76668-3|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037570|T201|OSN|76668-3|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037570|T201|LN|76668-3|LNC|CSF total protein|CSF total protein
C4037570|T201|LC|76668-3|LNC|CSF total protein|CSF total protein
C4037570|T201|MTH_LN|76668-3|LNC|CSF total protein|CSF total protein
C4037570|T201|OSN|76668-3|LNC|CSF total protein|CSF total protein
C4037570|T201|LN|76668-3|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037570|T201|LC|76668-3|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037570|T201|MTH_LN|76668-3|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037570|T201|OSN|76668-3|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037676|T201|LN|76667-5|LNC|CSF protein|CSF protein
C4037676|T201|OSN|76667-5|LNC|CSF protein|CSF protein
C4037676|T201|LC|76667-5|LNC|CSF protein|CSF protein
C4037676|T201|MTH_LN|76667-5|LNC|CSF protein|CSF protein
C4037676|T201|LN|76667-5|LNC|protein in csf|protein in csf
C4037676|T201|OSN|76667-5|LNC|protein in csf|protein in csf
C4037676|T201|LC|76667-5|LNC|protein in csf|protein in csf
C4037676|T201|MTH_LN|76667-5|LNC|protein in csf|protein in csf
C4037676|T201|LN|76667-5|LNC|Spinal fluid protein|Spinal fluid protein
C4037676|T201|OSN|76667-5|LNC|Spinal fluid protein|Spinal fluid protein
C4037676|T201|LC|76667-5|LNC|Spinal fluid protein|Spinal fluid protein
C4037676|T201|MTH_LN|76667-5|LNC|Spinal fluid protein|Spinal fluid protein
C4037676|T201|LN|76667-5|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037676|T201|OSN|76667-5|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037676|T201|LC|76667-5|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037676|T201|MTH_LN|76667-5|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037676|T201|LN|76667-5|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037676|T201|OSN|76667-5|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037676|T201|LC|76667-5|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037676|T201|MTH_LN|76667-5|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037676|T201|LN|76667-5|LNC|CSF total protein|CSF total protein
C4037676|T201|OSN|76667-5|LNC|CSF total protein|CSF total protein
C4037676|T201|LC|76667-5|LNC|CSF total protein|CSF total protein
C4037676|T201|MTH_LN|76667-5|LNC|CSF total protein|CSF total protein
C4037676|T201|LN|76667-5|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037676|T201|OSN|76667-5|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037676|T201|LC|76667-5|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037676|T201|MTH_LN|76667-5|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037677|T201|LN|76666-7|LNC|CSF protein|CSF protein
C4037677|T201|OSN|76666-7|LNC|CSF protein|CSF protein
C4037677|T201|MTH_LN|76666-7|LNC|CSF protein|CSF protein
C4037677|T201|LC|76666-7|LNC|CSF protein|CSF protein
C4037677|T201|LN|76666-7|LNC|protein in csf|protein in csf
C4037677|T201|OSN|76666-7|LNC|protein in csf|protein in csf
C4037677|T201|MTH_LN|76666-7|LNC|protein in csf|protein in csf
C4037677|T201|LC|76666-7|LNC|protein in csf|protein in csf
C4037677|T201|LN|76666-7|LNC|Spinal fluid protein|Spinal fluid protein
C4037677|T201|OSN|76666-7|LNC|Spinal fluid protein|Spinal fluid protein
C4037677|T201|MTH_LN|76666-7|LNC|Spinal fluid protein|Spinal fluid protein
C4037677|T201|LC|76666-7|LNC|Spinal fluid protein|Spinal fluid protein
C4037677|T201|LN|76666-7|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037677|T201|OSN|76666-7|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037677|T201|MTH_LN|76666-7|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037677|T201|LC|76666-7|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037677|T201|LN|76666-7|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037677|T201|OSN|76666-7|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037677|T201|MTH_LN|76666-7|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037677|T201|LC|76666-7|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037677|T201|LN|76666-7|LNC|CSF total protein|CSF total protein
C4037677|T201|OSN|76666-7|LNC|CSF total protein|CSF total protein
C4037677|T201|MTH_LN|76666-7|LNC|CSF total protein|CSF total protein
C4037677|T201|LC|76666-7|LNC|CSF total protein|CSF total protein
C4037677|T201|LN|76666-7|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037677|T201|OSN|76666-7|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037677|T201|MTH_LN|76666-7|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037677|T201|LC|76666-7|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037678|T201|LN|76665-9|LNC|CSF protein|CSF protein
C4037678|T201|OSN|76665-9|LNC|CSF protein|CSF protein
C4037678|T201|MTH_LN|76665-9|LNC|CSF protein|CSF protein
C4037678|T201|LC|76665-9|LNC|CSF protein|CSF protein
C4037678|T201|LN|76665-9|LNC|protein in csf|protein in csf
C4037678|T201|OSN|76665-9|LNC|protein in csf|protein in csf
C4037678|T201|MTH_LN|76665-9|LNC|protein in csf|protein in csf
C4037678|T201|LC|76665-9|LNC|protein in csf|protein in csf
C4037678|T201|LN|76665-9|LNC|Spinal fluid protein|Spinal fluid protein
C4037678|T201|OSN|76665-9|LNC|Spinal fluid protein|Spinal fluid protein
C4037678|T201|MTH_LN|76665-9|LNC|Spinal fluid protein|Spinal fluid protein
C4037678|T201|LC|76665-9|LNC|Spinal fluid protein|Spinal fluid protein
C4037678|T201|LN|76665-9|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037678|T201|OSN|76665-9|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037678|T201|MTH_LN|76665-9|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037678|T201|LC|76665-9|LNC|Cerebrospinal fluid protein|Cerebrospinal fluid protein
C4037678|T201|LN|76665-9|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037678|T201|OSN|76665-9|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037678|T201|MTH_LN|76665-9|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037678|T201|LC|76665-9|LNC|Cerebrospinal fluid with protein|Cerebrospinal fluid with protein
C4037678|T201|LN|76665-9|LNC|CSF total protein|CSF total protein
C4037678|T201|OSN|76665-9|LNC|CSF total protein|CSF total protein
C4037678|T201|MTH_LN|76665-9|LNC|CSF total protein|CSF total protein
C4037678|T201|LC|76665-9|LNC|CSF total protein|CSF total protein
C4037678|T201|LN|76665-9|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037678|T201|OSN|76665-9|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037678|T201|MTH_LN|76665-9|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037678|T201|LC|76665-9|LNC|cerebrospinal fluid total protein|cerebrospinal fluid total protein
C4037760|T201|LN|76482-9|LNC|apolipoprotein B|apolipoprotein B
C4037760|T201|OSN|76482-9|LNC|apolipoprotein B|apolipoprotein B
C4037760|T201|LC|76482-9|LNC|apolipoprotein B|apolipoprotein B
C4037760|T201|MTH_LN|76482-9|LNC|apolipoprotein B|apolipoprotein B
C4037760|T201|LN|76482-9|LNC|ApoB|ApoB
C4037760|T201|OSN|76482-9|LNC|ApoB|ApoB
C4037760|T201|LC|76482-9|LNC|ApoB|ApoB
C4037760|T201|MTH_LN|76482-9|LNC|ApoB|ApoB
C4037792|T201|LN|76399-5|LNC|troponin I|troponin I
C4037792|T201|LC|76399-5|LNC|troponin I|troponin I
C4037792|T201|OSN|76399-5|LNC|troponin I|troponin I
C4037792|T201|MTH_LN|76399-5|LNC|troponin I|troponin I
C4070134|T201|LN|79469-3|LNC|uridine diphosphate glucose-4-epimerase activity in red|uridine diphosphate glucose-4-epimerase activity in red
C4070134|T201|OSN|79469-3|LNC|uridine diphosphate glucose-4-epimerase activity in red|uridine diphosphate glucose-4-epimerase activity in red
C4070134|T201|LC|79469-3|LNC|uridine diphosphate glucose-4-epimerase activity in red|uridine diphosphate glucose-4-epimerase activity in red
C4070134|T201|MTH_LN|79469-3|LNC|uridine diphosphate glucose-4-epimerase activity in red|uridine diphosphate glucose-4-epimerase activity in red
C4070134|T201|LN|79469-3|LNC|UDP-glucose 4-epimerase activity activity in red|UDP-glucose 4-epimerase activity activity in red
C4070134|T201|OSN|79469-3|LNC|UDP-glucose 4-epimerase activity activity in red|UDP-glucose 4-epimerase activity activity in red
C4070134|T201|LC|79469-3|LNC|UDP-glucose 4-epimerase activity activity in red|UDP-glucose 4-epimerase activity activity in red
C4070134|T201|MTH_LN|79469-3|LNC|UDP-glucose 4-epimerase activity activity in red|UDP-glucose 4-epimerase activity activity in red
C4070658|T201|LN|78857-0|LNC|methadone test|methadone test
C4070658|T201|MTH_LN|78857-0|LNC|methadone test|methadone test
C4070658|T201|OSN|78857-0|LNC|methadone test|methadone test
C4070658|T201|LC|78857-0|LNC|methadone test|methadone test
C4070824|T201|LN|78770-5|LNC|methadone test|methadone test
C4070824|T201|MTH_LN|78770-5|LNC|methadone test|methadone test
C4070824|T201|LC|78770-5|LNC|methadone test|methadone test
C4070824|T201|OSN|78770-5|LNC|methadone test|methadone test
C4265794|T201|LN|80964-0|LNC|xenobiotic|xenobiotic
C4265794|T201|LC|80964-0|LNC|xenobiotic|xenobiotic
C4265794|T201|OSN|80964-0|LNC|xenobiotic|xenobiotic
C4265794|T201|MTH_LN|80964-0|LNC|xenobiotic|xenobiotic
C4297159|T201|LN|85066-9|LNC|estradiol|estradiol
C4297159|T201|LC|85066-9|LNC|estradiol|estradiol
C4297159|T201|MTH_LN|85066-9|LNC|estradiol|estradiol
C4297159|T201|OSN|85066-9|LNC|estradiol|estradiol
C4298232|T201|LN|83103-2|LNC|luteinizing|luteinizing
C4298232|T201|LC|83103-2|LNC|luteinizing|luteinizing
C4298232|T201|MTH_LN|83103-2|LNC|luteinizing|luteinizing
C4298232|T201|OSN|83103-2|LNC|luteinizing|luteinizing
C4298232|T201|LN|83103-2|LNC|LH|LH
C4298232|T201|LC|83103-2|LNC|LH|LH
C4298232|T201|MTH_LN|83103-2|LNC|LH|LH
C4298232|T201|OSN|83103-2|LNC|LH|LH
C4298232|T201|LN|83103-2|LNC|luteinising|luteinising
C4298232|T201|LC|83103-2|LNC|luteinising|luteinising
C4298232|T201|MTH_LN|83103-2|LNC|luteinising|luteinising
C4298232|T201|OSN|83103-2|LNC|luteinising|luteinising
C4298267|T201|LN|83117-2|LNC|Autoimmune antibody|Autoimmune antibody
C4298267|T201|OSN|83117-2|LNC|Autoimmune antibody|Autoimmune antibody
C4298267|T201|LC|83117-2|LNC|Autoimmune antibody|Autoimmune antibody
C4298267|T201|MTH_LN|83117-2|LNC|Autoimmune antibody|Autoimmune antibody
C4298342|T201|LN|82928-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C4298342|T201|MTH_LN|82928-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C4298342|T201|LC|82928-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C4298342|T201|OSN|82928-3|LNC|Anti-mitochondrial M2 antibody|Anti-mitochondrial M2 antibody
C4482807|T201|LN|85369-7|LNC|neutrophil counts|neutrophil counts
C4482807|T201|MTH_LN|85369-7|LNC|neutrophil counts|neutrophil counts
C4482807|T201|OSN|85369-7|LNC|neutrophil counts|neutrophil counts
C4482807|T201|LC|85369-7|LNC|neutrophil counts|neutrophil counts
C4482807|T201|LN|85369-7|LNC|neutrophil count|neutrophil count
C4482807|T201|MTH_LN|85369-7|LNC|neutrophil count|neutrophil count
C4482807|T201|OSN|85369-7|LNC|neutrophil count|neutrophil count
C4482807|T201|LC|85369-7|LNC|neutrophil count|neutrophil count
C4482807|T201|LN|85369-7|LNC|neutrophil|neutrophil
C4482807|T201|MTH_LN|85369-7|LNC|neutrophil|neutrophil
C4482807|T201|OSN|85369-7|LNC|neutrophil|neutrophil
C4482807|T201|LC|85369-7|LNC|neutrophil|neutrophil
C4531914|T201|LN|86911-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C4531914|T201|OSN|86911-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C4531914|T201|LC|86911-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C4531914|T201|MTH_LN|86911-5|LNC|low-density lipoprotein cholesterol|low-density lipoprotein cholesterol
C4531914|T201|LN|86911-5|LNC|LDL|LDL
C4531914|T201|OSN|86911-5|LNC|LDL|LDL
C4531914|T201|LC|86911-5|LNC|LDL|LDL
C4531914|T201|MTH_LN|86911-5|LNC|LDL|LDL
C4531914|T201|LN|86911-5|LNC|LDL cholesterol|LDL cholesterol
C4531914|T201|OSN|86911-5|LNC|LDL cholesterol|LDL cholesterol
C4531914|T201|LC|86911-5|LNC|LDL cholesterol|LDL cholesterol
C4531914|T201|MTH_LN|86911-5|LNC|LDL cholesterol|LDL cholesterol
C4531914|T201|LN|86911-5|LNC|low-density lipoprotein|low-density lipoprotein
C4531914|T201|OSN|86911-5|LNC|low-density lipoprotein|low-density lipoprotein
C4531914|T201|LC|86911-5|LNC|low-density lipoprotein|low-density lipoprotein
C4531914|T201|MTH_LN|86911-5|LNC|low-density lipoprotein|low-density lipoprotein
C4531914|T201|LN|86911-5|LNC|beta-lipoproteins|beta-lipoproteins
C4531914|T201|OSN|86911-5|LNC|beta-lipoproteins|beta-lipoproteins
C4531914|T201|LC|86911-5|LNC|beta-lipoproteins|beta-lipoproteins
C4531914|T201|MTH_LN|86911-5|LNC|beta-lipoproteins|beta-lipoproteins
C4531914|T201|LN|86911-5|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C4531914|T201|OSN|86911-5|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C4531914|T201|LC|86911-5|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C4531914|T201|MTH_LN|86911-5|LNC|LDL cholesterol conncentration|LDL cholesterol conncentration
C4531914|T201|LN|86911-5|LNC|LDL-C|LDL-C
C4531914|T201|OSN|86911-5|LNC|LDL-C|LDL-C
C4531914|T201|LC|86911-5|LNC|LDL-C|LDL-C
C4531914|T201|MTH_LN|86911-5|LNC|LDL-C|LDL-C
C4533466|T201|LN|88059-1|LNC|xenobiotic|xenobiotic
C4533466|T201|OSN|88059-1|LNC|xenobiotic|xenobiotic
C4533466|T201|LC|88059-1|LNC|xenobiotic|xenobiotic
C4533466|T201|MTH_LN|88059-1|LNC|xenobiotic|xenobiotic
