C0002059|T034||LNC|ALKALINE PHOSPHATASE
C0201850|T034||LNC|ALKALINE PHOSPHATASE MEASUREMENT
C0443450|T034||LNC|ALK. PHOS. - BILE ISOENZYME
C0443450|T034||LNC|THIS IS THE MORE SPECFIC ISOENZYME OF AP THAT YOU'D ACTUALLY CARE ABOUT WHEN LOOKING AT LFTS. I'M NOT SURE IF IT'S AN INCLUDE OR EXCLUDE, I'D ASK YOUR CMO ABOUT APPROPRIATENESS
C0443450|T034||LNC|ALKALINE PHOSPHATASE BILIARY ISOENZYME 
C0301810|T034|LP18187-2|LNC|SAME AS ABOVE, MORE SPECIFIC BUT MAY WANT TO INCLUDE|ALKALINE PHOSPHATASE ISOENZYME
C0301810|T034|LP18187-2|LNC|ALKALINE PHOSPHATASE ISOENZYME|ALKALINE PHOSPHATASE ISOENZYME
C0301810|T034|LP18187-2|LNC|ALKALINE PHOSPHATASE ISOENZYME |ALKALINE PHOSPHATASE ISOENZYME
C0301810|T034|LP18187-2|LNC|ALKALINE PHOSPHATASE ISOENZYME, NOS|ALKALINE PHOSPHATASE ISOENZYME
C0312398|T034||LNC|ALKALINE PHOSPHATASE.LIVER
C0312398|T034||LNC|ALK. PHOS. - LIVER ISOENZYME
C0312398|T034||LNC|LIVER ALKALINE PHOSPHATASE
C0312398|T034||LNC|ALKALINE PHOSPHATASE ISOENZYME, LIVER FRACTION
C0312398|T034||LNC|ALKALINE PHOSPHATASE LIVER ISOENZYME
C0312398|T034||LNC|ALKALINE PHOSPHATASE ISOENZYME, LIVER FRACTION 
C0002059|T034||LNC|ALKALINE PHOSPHATASE
C0002059|T034||LNC|AP
C0002059|T034||LNC|ALKALINE PHOSPHOMONOESTERASE
C0002059|T034||LNC|APPARENTLY THIS IS AP, NEVER SEEN THIS NAME USED
C0002059|T034||LNC|ALKALINE PHOSPHATASE [CHEMICAL/INGREDIENT]
C0002059|T034||LNC|ALP - ALKALINE PHOSPHATASE
C0002059|T034||LNC|AP - ALKALINE PHOSPHATASE
C0002059|T034||LNC|ALKALINE PHOSPHATASE 
C2932888|T034||LNC|ALKALINE PHOSPHATASE, LIVER-BONE-KIDNEY, HUMAN
C2932888|T034||LNC|THIS IS THE TISSUE NON-SPECIFIC AP SO IS A SYNONYM, BUT WOULD BE SURPRISED TO SEE IT EVER LISTED THIS WAY
C2932888|T034||LNC|TNAP PHOSPHATASE, HUMAN
C2932888|T034||LNC|TISSUE-NON SPECIFIC ALKALINE PHOSPHATASE, HUMAN
C2932888|T034||LNC|LIVER/BONE/KIDNEY-TYPE ALKALINE PHOSPHATASE
C2932888|T034||LNC|ALKALINE PHOSPHATASE, TISSUE-NONSPECIFIC ISOZYME
C2932888|T034||LNC|TISSUE-NONSPECIFIC ALP
C2932888|T034||LNC|EC 3.1.3.1
C2932888|T034||LNC|ALKALINE PHOSPHOMONOESTERASE
C1318717|T034||LNC|ALKALINE PHOSPHATASE
C1980986|T034|LP45609-2|LNC|ALKALINE PHOSPHATASE &#X7C; BLD-SER-PLAS|ALKALINE PHOSPHATASE &#X7C; BLD-SER-PLAS
C2930591|T034||LNC|SYNONYM FOR AP - RARE
C1148297|T034||LNC|THIS IS THE LIVER SPECIFIC AP (BONE IS NOT HEAT STABLE?) - SAME AS SOME OTHERS, NOT SPECIFICALLY WHAT YOU'D TYPICALLY EXPECT, BUT IS VERY RELEVANT ??INCLUDE?? HTTPS://WWW.SHH.ORG/OUTPATIENT-SERVICES/LABORATORY-SERVICES/LABORATORY-TEST-PRINT.ASP?ID=55
C1148297|T034||LNC|HEAT STABLE ALKALINE PHOSPHATASE 
C1148297|T034||LNC|HEAT STABLE ALKALINE PHOSPHATASE
C0201850|T034||LNC|ALKALINE PHOSPHATASE MEASUREMENT
C0201850|T034||LNC|PHOSPHATASE, ALKALINE
C0201850|T034||LNC|ALP
C0201850|T034||LNC|TEST;ALKALINE PHOSPHATASE
C0201850|T034||LNC|MEASUREMENT OF ALKALINE PHOSPHATASE
C0201850|T034||LNC|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T034||LNC|ALKALINE PHOSPHATASE
C0201850|T034||LNC|ALK PHOSPH
C0201850|T034||LNC|ALK PHOS
C0201850|T034||LNC|ALKPHOS
C0201850|T034||LNC|ALK-PHOS
C0201850|T034||LNC|ALKALINE PHOSPHATASE MEASUREMENT 
C0201850|T034||LNC|ASSAY ALKALINE PHOSPHATASE
C0201850|T034||LNC|ALKALINE PHOSPHATASE TEST
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE MEASUREMENT
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE MEASUREMENT 
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE (& LEVEL)
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE (& LEVEL) 
C0036776|T034||LNC|ALK. PHOSPHATASE -SERUM
C0036776|T034||LNC|ALKALINE PHOSPHATASE (& LEVEL (& SERUM))
C0036776|T034||LNC|PHOSPH.- ALK. - SERUM
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE NOS
C0036776|T034||LNC|ALKALINE PHOSPHATASE (& LEVEL (& SERUM)) 
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE NOS 
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE TEST
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE LEVEL
C0036776|T034||LNC|SERUM ALKALINE PHOSPHATASE MEASUREMENT 
C0201851|T034||LNC|PHOSPHATASE, ALKALINE; ISOENZYMES
C0201851|T034||LNC|MEASUREMENT OF ALKALINE PHOSPHATASE ISOENZYMES
C0201851|T034||LNC|ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES
C0201851|T034||LNC|ALKALINE PHOSPHATASE ISOENZYMES MEASUREMENT
C0201851|T034||LNC|ALKALINE PHOSPHATASE ISOENZYMES MEASUREMENT 
C0201851|T034||LNC|ASSAY ALKALINE PHOSPHATASES
C0201855|T034||LNC|ALKALINE PHOSPHATASE, HEAT STABLE MEASUREMENT
C0201855|T034||LNC|PHOSPHATASE, ALKALINE; HEAT STABLE (TOTAL NOT INCLUDED)
C0201855|T034||LNC|MEASUREMENT OF HEAT STABLE ALKALINE PHOSPHATASE
C0201855|T034||LNC|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C0201855|T034||LNC|THERMOSTABLE ALKALINE PHOSPHATASE MEASUREMENT
C0201855|T034||LNC|ALKALINE PHOSPHATASE, HEAT STABLE MEASUREMENT 
C0201855|T034||LNC|ASSAY ALKALINE PHOSPHATASE
C3898585|T034||LNC|LIVER SPECIFIC ALKALINE PHOSPHATASE MEASUREMENT
C3898585|T034||LNC|ALPLS
C3898585|T034||LNC|LIVER SPECIFIC ALKALINE PHOSPHATASE
C3898710|T034||LNC|INTESTINAL SPECIFIC ALKALINE PHOSPHATASE
C1272113|T034||LNC|PLASMA ALKALINE PHOSPHATASE LEVEL 
C1272113|T034||LNC|PLASMA ALKALINE PHOSPHATASE LEVEL
