C1255280|T034||LNC|25-OH D VITAMIN TEST
C1255280|T034||LNC|VIT D 25-OH
C1255280|T034||LNC|VITAMIN D 25-OH
C1255280|T034||LNC|VITAMIN D 25-OH
