C0333106|T047|57052009|SNOMEDCT_US|BLEEDING VARICES|BLEEDING VARICES (MORPHOLOGIC ABNORMALITY)
C3837381|T047||SNOMEDCT_US|GASTRIC VARICEAL PROCEDURES
C4288030|T047||SNOMEDCT_US|VARICEAL BANDING
C0192331|T047|149327003|SNOMEDCT_US|LIGATION OF ESOPHAGEAL VARICES|LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192558|T047|80444007|SNOMEDCT_US|STAPLING OF GASTRIC VARICES|STAPLING OF GASTRIC VARICES (PROCEDURE)
C0852804|T047||SNOMEDCT_US|OESOPHAGEAL VARICEAL INJECTION
C1739112|T047||SNOMEDCT_US|GASTROOESOPHAGEAL VARICEAL HAEMORRHAGE PROPHYLAXIS
C2062316|T047||SNOMEDCT_US|ACUTE BLEEDING OF ESOPHAGEAL VARICES
C2065631|T047||SNOMEDCT_US|ESOPHAGOSCOPY RIGID VARICEAL SCLEROTHERAPY
C2960232|T047|446740007|SNOMEDCT_US|BANDING OF VARIX OF STOMACH|BANDING OF GASTRIC VARICES
C3837654|T047||SNOMEDCT_US|ESOPHAGUS VARICEAL SURGERY
C3888799|T047||SNOMEDCT_US|GASTRIC VARICEAL INJECTION
C3888800|T047||SNOMEDCT_US|GASTRIC VARICEAL LIGATION
C4272078|T047||SNOMEDCT_US|SUGIURA VARICEAL PROCEDURE
C3694764|T047||SNOMEDCT_US|ESOPHAGOSCOPY TRANSORAL FLEXIBLE WITH VARICEAL SCLEROTHERAPY
C0547715|T047||SNOMEDCT_US|FOLLOW PROTOCOL FOR VASOPRESSIN OR NITROGLYCERINE THERAPY OF VARICEAL HEMORRHAGE
C0333106|T047|57052009|SNOMEDCT_US|BLEEDING VARICES|BLEEDING VARICES (MORPHOLOGIC ABNORMALITY)
C0333106|T047|57052009|SNOMEDCT_US|BLEEDING VARICES (MORPHOLOGIC ABNORMALITY)|BLEEDING VARICES (MORPHOLOGIC ABNORMALITY)
C3837379|T047||SNOMEDCT_US|GASTRIC SURGERY VARICEAL STAPLING 
C3837379|T047||SNOMEDCT_US|GASTRIC SURGERY VARICEAL STAPLING
C2960232|T047|446740007|SNOMEDCT_US|BANDING OF VARIX OF STOMACH |BANDING OF GASTRIC VARICES
C2960232|T047|446740007|SNOMEDCT_US|BANDING OF GASTRIC VARICES|BANDING OF GASTRIC VARICES
C2960232|T047|446740007|SNOMEDCT_US|BANDING OF VARIX OF STOMACH|BANDING OF GASTRIC VARICES
C2960232|T047|446740007|SNOMEDCT_US|GASTRIC SURGERY VARICEAL BANDING|BANDING OF GASTRIC VARICES
C2960232|T047|446740007|SNOMEDCT_US|BANDING OF GASTRIC VARICES |BANDING OF GASTRIC VARICES
C3837380|T047||SNOMEDCT_US|GASTRIC SURGERY VARICEAL LIGATION
C3837380|T047||SNOMEDCT_US|GASTRIC SURGERY VARICEAL LIGATION 
C0192331|T047|149327003|SNOMEDCT_US|LIGATION OF ESOPHAGEAL VARICES |LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192331|T047|149327003|SNOMEDCT_US|LIGATION OF ESOPHAGEAL VARICES|LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192331|T047|149327003|SNOMEDCT_US|OESOPHAGEAL VARICEAL LIGATION|LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192331|T047|149327003|SNOMEDCT_US|LIGATION ESOPH VARIX|LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192331|T047|149327003|SNOMEDCT_US|LOCAL LIGATION OF OESOPHAGEAL VARICES |LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192331|T047|149327003|SNOMEDCT_US|LOCAL LIGATION OF ESOPHAGEAL VARICES|LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192331|T047|149327003|SNOMEDCT_US|LOCAL LIGATION OF OESOPHAGEAL VARICES|LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192331|T047|149327003|SNOMEDCT_US|LIGATION OF OESOPHAGEAL VARICES|LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192331|T047|149327003|SNOMEDCT_US|ESOPHAGEAL VARICEAL LIGATION|LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0192331|T047|149327003|SNOMEDCT_US|LIGATION OF ESOPHAGEAL VARICES |LOCAL LIGATION OF OESOPHAGEAL VARICES (PROCEDURE)
C0372009|T047||SNOMEDCT_US|LIGATION, DIRECT, ESOPHAGEAL VARICES
C0372009|T047||SNOMEDCT_US|LIGATION DIRECT ESOPHAGEAL VARICES
C0372009|T047||SNOMEDCT_US|DIRECT LIGATION OF ESOPHAGEAL VARICES
C0372009|T047||SNOMEDCT_US|LIGATE ESOPHAGUS VEINS
C0852804|T047||SNOMEDCT_US|OESOPHAGEAL VARICEAL INJECTION
C0852804|T047||SNOMEDCT_US|ESOPHAGEAL VARICEAL INJECTION
C0852804|T047||SNOMEDCT_US|INJECTION OF ESOPHAGEAL VARICES
C0852804|T047||SNOMEDCT_US|INJECTION OF OESOPHAGEAL VARICES
C1739112|T047||SNOMEDCT_US|GASTROOESOPHAGEAL VARICEAL HAEMORRHAGE PROPHYLAXIS
C1739112|T047||SNOMEDCT_US|GASTROOESOPHAGEAL VARICEAL HEMORRHAGE PROPHYLAXIS
C1739112|T047||SNOMEDCT_US|GASTROESOPHAGEAL VARICEAL HEMORRHAGE PROPHYLAXIS
C1739112|T047||SNOMEDCT_US|PROPHYLAXIS OF GASTROOESOPHAGEAL VARICEAL BLEEDING
C1739112|T047||SNOMEDCT_US|PROPHYLAXIS OF GASTROESOPHAGEAL VARICEAL BLEEDING
C0472988|T047|173660005|SNOMEDCT_US|ENDOSCOPIC INJECTION SCLEROTHERAPY TO VARICES OF ESOPHAGUS USING RIGID ESOPHAGOSCOPE|RIGID ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES (PROCEDURE)
C0472988|T047|173660005|SNOMEDCT_US|ENDOSCOPIC INJECTION SCLEROTHERAPY TO VARICES OF OESOPHAGUS USING RIGID OESOPHAGOSCOPE|RIGID ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES (PROCEDURE)
C0472988|T047|173660005|SNOMEDCT_US|RIGID ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES|RIGID ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES (PROCEDURE)
C0472988|T047|173660005|SNOMEDCT_US|RIGID OESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES|RIGID ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES (PROCEDURE)
C0472988|T047|173660005|SNOMEDCT_US|RIGID ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES |RIGID ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES (PROCEDURE)
C2959927|T047|446743009|SNOMEDCT_US|OESOPHAGOGASTRODUODENOSCOPY AND BANDING OF GASTRIC VARICES|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF STOMACH (PROCEDURE)
C2959927|T047|446743009|SNOMEDCT_US|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF STOMACH|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF STOMACH (PROCEDURE)
C2959927|T047|446743009|SNOMEDCT_US|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF GASTRIC VARICES|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF STOMACH (PROCEDURE)
C2959927|T047|446743009|SNOMEDCT_US|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF STOMACH |ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF STOMACH (PROCEDURE)
C2959927|T047|446743009|SNOMEDCT_US|ESOPHAGOGASTRODUODENOSCOPY AND BANDING OF GASTRIC VARICES|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF STOMACH (PROCEDURE)
C0472950|T047|265863006|SNOMEDCT_US|OESOPH. VARICES OPN.|VARICES - OESOPH.- OPN.
C0472950|T047|265863006|SNOMEDCT_US|OPERATION ON OESOPHAGEAL VARICES|VARICES - OESOPH.- OPN.
C0472950|T047|265863006|SNOMEDCT_US|VARICES - OESOPH.- OPN.|VARICES - OESOPH.- OPN.
C0472950|T047|265863006|SNOMEDCT_US|OPERATION ON ESOPHAGEAL VARICES|VARICES - OESOPH.- OPN.
C0472950|T047|265863006|SNOMEDCT_US|OPERATION ON ESOPHAGEAL VARICES |VARICES - OESOPH.- OPN.
C3888799|T047||SNOMEDCT_US|GASTRIC VARICEAL INJECTION
C3888800|T047||SNOMEDCT_US|GASTRIC VARICEAL LIGATION
