C0201838|T034||LNC|ALBUMIN MEASUREMENT
C0523464|T034||LNC|ALBUMIN RENAL CLEARANCE MEASUREMENT
C0523464|T034||LNC|ALBUMIN RENAL CLEARANCE MEASUREMENT 
C0523465|T034||LNC|SERUM ALBUMIN
C0523465|T034||LNC|SERUM ALBUMIN MEASUREMENT
C0523465|T034||LNC|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T034||LNC|ALBUMIN; SERUM, PLASMA OR WHOLE BLOOD
C0523465|T034||LNC|SERUM ALBUMIN MEASUREMENT 
C0523465|T034||LNC|MEASUREMENT OF ALBUMIN IN SERUM
C0523465|T034||LNC|SERUM ALBUMIN (& LEVEL) 
C0523465|T034||LNC|ALBUMIN - SERUM
C0523465|T034||LNC|SERUM ALBUMIN (& LEVEL)
C0523465|T034||LNC|SERUM ALBUMIN TEST
C0523465|T034||LNC|ALBUMIN MEASUREMENT, SERUM
C0523465|T034||LNC|SERUM ALBUMIN LEVEL
C0523465|T034||LNC|SA - SERUM ALBUMIN
C0523465|T034||LNC|ALBUMIN MEASUREMENT, SERUM 
C0523465|T034||LNC|ASSAY OF SERUM ALBUMIN
C0201838|T034||LNC|ALBUMIN MEASUREMENT
C0201838|T034||LNC|TEST;ALBUMIN
C0201838|T034||LNC|MEASUREMENT OF ALBUMIN
C0201838|T034||LNC|ALBUMIN
C0201838|T034||LNC|ALB
C0201838|T034||LNC|ALBUMIN MEASUREMENT 
C0201838|T034||LNC|ALBUMIN TEST
# C0428520|T034||LNC|I SUSPECT THIS WILL WIND UP RETURNING ALBUMIN LEVELS FROM PERITONEAL FLUID ETC. KEEP IT ON YOUR RADAR TO EXCLUDE - YOU CARE ONLY ABOUT SERUM ALBUMIN (FOR YOUR FORM)
C1272106|T034||LNC|PLASMA ALBUMIN LEVEL 
C1272106|T034||LNC|PLASMA ALBUMIN LEVEL
