C0018935|T034|LP15101-6|LNC|HCT|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT PROCEDURE|HEMATOCRIT
C0518014|T034||LNC|HEMATOCRIT
C1542366|T034||LNC|HEMATOCRIT
C1545323|T034|MTHU017408|LNC|HEMATOCRIT TEST STATUS|HEMATOCRIT TEST STATUS
C1627395|T034|MTHU018856|LNC|HEMATOCRIT TEST RESULTS|HEMATOCRIT TEST STATUS &OR RESULTS
C1627395|T034|MTHU018856|LNC|HEMATOCRIT TEST STATUS &OR RESULTS|HEMATOCRIT TEST STATUS &OR RESULTS
C1627395|T034|MTHU018856|LNC|HEMATOCRIT TEST STATUS OR RESULTS|HEMATOCRIT TEST STATUS &OR RESULTS
C1254918|T034||LNC|OPERATING ROOM MISC LABS: HCT
C0018935|T034|LP15101-6|LNC|HCT|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|ERYTHROCYTE VOLUMES, PACKED|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRITS|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PACKED ERYTHROCYTE VOLUME|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PACKED ERYTHROCYTE VOLUMES|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PACKED RED CELL VOLUME|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PACKED RED-CELL VOLUMES|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|RED-CELL VOLUME, PACKED|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|RED-CELL VOLUMES, PACKED|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|VOLUME, PACKED ERYTHROCYTE|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|VOLUME, PACKED RED-CELL|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|VOLUMES, PACKED ERYTHROCYTE|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|VOLUMES, PACKED RED-CELL|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HAEMATOCRIT|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT PROCEDURE|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT |HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT MEASUREMENT|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|BLOOD COUNT HEMATOCRIT|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|MEASUREMENT OF HEMATOCRIT (HCT)|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PACKED CELL VOLUME (OBSERVABLE ENTITY)|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HAEMATOCRIT - PCV - NOS|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PACKED CELL VOLUME|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HAEMATOCRIT (OBSERVABLE ENTITY)|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HAEMATOCRIT |HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT - PCV - NOS|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HAEMATOCRIT - PCV - NOS |HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT - PCV - NOS |HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT PACKED CELL VOLUME |HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT PACKED CELL VOLUME|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|EVF|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PCV|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|ERYTHROCYTE VOLUME FRACTION|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|BLOOD COUNT; HEMATOCRIT (HCT)|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PACKED RED-CELL VOLUME|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|ERYTHROCYTE VOLUME, PACKED|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|WHOLE BLOOD HEMATOCRIT TEST|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT DETERMINATION|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HAEMATOCRIT - PCV|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HCT - HAEMATOCRIT|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HCT - HEMATOCRIT|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT - PCV|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HAEMATOCRIT DETERMINATION|HEMATOCRIT
C0018935|T034|LP15101-6|LNC|HEMATOCRIT DETERMINATION |HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PACKED CELL VOLUME MEASUREMENT |HEMATOCRIT
C0018935|T034|LP15101-6|LNC|PACKED CELL VOLUME MEASUREMENT|HEMATOCRIT
C0373755|T034||LNC|EQUIVALENT BUT DIFFERENT THAN A CBC HCT
C0373755|T034||LNC|MICROHEMATOCRIT (SPUN) 
C0373755|T034||LNC|MICROHEMATOCRIT (SPUN)
C0373755|T034||LNC|MICROHEMATOCRIT LEVEL
C0373755|T034||LNC|BLOOD COUNT SPUN MICROHEMATOCRIT
C0373755|T034||LNC|MEASUREMENT OF SPUN MICROHEMATOCRIT
C0373755|T034||LNC|SPUN MICROHEMATOCRIT
C0518014|T034||LNC|HEMATOCRIT
C0518014|T034||LNC|HEMATOCRIT LEVEL
C0518014|T034||LNC|HEMATOCRIT (HCT)
C0518014|T034||LNC|FINDING OF HAEMATOCRIT
C0518014|T034||LNC|FINDING OF HEMATOCRIT
C0518014|T034||LNC|HEMATOCRIT FINDING
C0518014|T034||LNC|HEMATOCRIT FINDING 
C0518014|T034||LNC|HAEMATOCRIT
C0518014|T034||LNC|FINDING OF HEMATOCRIT 
C0518014|T034||LNC|HAEMATOCRIT - FINDING
C0518014|T034||LNC|HEMATOCRIT - FINDING
C1988891|T034|LP52614-2|LNC|HEMATOCRIT &#X7C; BLOOD CAPILLARY|HEMATOCRIT &#X7C; BLOOD CAPILLARY
C1988890|T034|LP50017-0|LNC|HEMATOCRIT &#X7C; BLOOD ARTERIAL|HEMATOCRIT &#X7C; BLOOD ARTERIAL
C1988893|T034|LP52291-9|LNC|HEMATOCRIT &#X7C; BLOOD MIXED VENOUS|HEMATOCRIT &#X7C; BLOOD MIXED VENOUS
C1988889|T034|LP45040-0|LNC|HEMATOCRIT &#X7C; BLD-SER-PLAS|HEMATOCRIT &#X7C; BLD-SER-PLAS
C1988894|T034|LP52290-1|LNC|HEMATOCRIT &#X7C; BLOOD VENOUS|HEMATOCRIT &#X7C; BLOOD VENOUS
C3837271|T034||LNC|HEMATOCRIT PACKED CELL VOLUME FINDING
C3837271|T034||LNC|HEMATOCRIT PACKED CELL VOLUME FINDING 
C4028949|T034||LNC|HEMATOCRIT LEVEL BY AUTOMATED COUNT
C4028949|T034||LNC|HEMATOCRIT LEVEL BY AUTOMATED COUNT 
C4028949|T034||LNC|HEMATOCRIT BY AUTOMATED COUNT
C4064964|T034||LNC|HEMATOCRIT LEVEL BY IMPEDANCE 
C4064964|T034||LNC|HEMATOCRIT BY IMPEDANCE
C4064964|T034||LNC|HEMATOCRIT LEVEL BY IMPEDANCE
C0523148|T034||LNC|HAEMATOCRIT, SPUN MICROHAEMATOCRIT METHOD
C0523148|T034||LNC|HEMATOCRIT, SPUN MICROHEMATOCRIT METHOD
C0523148|T034||LNC|HEMATOCRIT, SPUN MICROHEMATOCRIT METHOD 
C1443988|T034||LNC|SERIAL HAEMATOCRIT DETERMINATIONS
C1443988|T034||LNC|SERIAL HEMATOCRIT DETERMINATIONS 
C1443988|T034||LNC|SERIAL HEMATOCRIT DETERMINATIONS
C0580315|T034||LNC|HAEMATOCRIT - PCV ABNORMAL 
C0580315|T034||LNC|HEMATOCRIT - PCV ABNORMAL
C0580315|T034||LNC|HAEMATOCRIT - PCV ABNORMAL
C0580315|T034||LNC|HEMATOCRIT - PACKED CELL VOLUME ABNORMAL 
C0580315|T034||LNC|HEMATOCRIT - PCV ABNORMAL 
C0580315|T034||LNC|HEMATOCRIT - PACKED CELL VOLUME ABNORMAL
C0580315|T034||LNC|HAEMATOCRIT - PACKED CELL VOLUME ABNORMAL
C0474548|T034||LNC|HAEMATOCRIT - PCV - NORMAL
C0474548|T034||LNC|HAEMATOCRIT - PCV - NORMAL 
C0474548|T034||LNC|HEMATOCRIT - PCV - NORMAL
C0474548|T034||LNC|HEMATOCRIT - PACKED CELL VOLUME - NORMAL
C0474548|T034||LNC|HEMATOCRIT - PACKED CELL VOLUME - NORMAL 
C0474548|T034||LNC|HEMATOCRIT - PCV - NORMAL 
C0474548|T034||LNC|HAEMATOCRIT - PACKED CELL VOLUME - NORMAL
C0474550|T034||LNC|HAEMATOCRIT - PCV - LOW 
C0474550|T034||LNC|HAEMATOCRIT - PCV - LOW
C0474550|T034||LNC|HEMATOCRIT - PCV - LOW
C0474550|T034||LNC|PACKED CELL VOLUME DECREASED BELOW NORMAL
C0474550|T034||LNC|HEMATOCRIT DECREASED BELOW NORMAL
C0474550|T034||LNC|HCT DECREASED
C0474550|T034||LNC|PCV DECREASED BELOW NORMAL
C0474550|T034||LNC|HEMATOCRIT - PACKED CELL VOLUME - LOW
C0474550|T034||LNC|HEMATOCRIT - PCV - LOW 
C0474550|T034||LNC|HEMATOCRIT - PACKED CELL VOLUME - LOW 
C0474550|T034||LNC|HAEMATOCRIT - PACKED CELL VOLUME - LOW
C0549409|T034||LNC|HAEMATOCRIT - PCV - HIGH 
C0549409|T034||LNC|HAEMATOCRIT - PCV - HIGH
C0549409|T034||LNC|HEMATOCRIT - PCV - HIGH
C0549409|T034||LNC|PCV INCREASED
C0549409|T034||LNC|HCT INCREASED
C0549409|T034||LNC|HEMATOCRIT INCREASED ABOVE NORMAL
C0549409|T034||LNC|HEMOCONCENTRATION
C0549409|T034||LNC|PACKED CELL VOLUME INCREASED ABOVE NORMAL
C0549409|T034||LNC|HEMATOCRIT - PCV - HIGH 
C0549409|T034||LNC|HEMATOCRIT - PACKED CELL VOLUME - HIGH 
C0549409|T034||LNC|HEMATOCRIT - PACKED CELL VOLUME - HIGH
C0549409|T034||LNC|HAEMATOCRIT - PACKED CELL VOLUME - HIGH
C0549409|T034||LNC|PACKED CELL VOLUME INCREASED
C0474547|T034||LNC|HAEMATOCRIT - BORDERLINE HIGH
C0474547|T034||LNC|HAEMATOCRIT - BORDERLINE HIGH 
C0474547|T034||LNC|HEMATOCRIT - BORDERLINE HIGH
C0474547|T034||LNC|HEMATOCRIT - BORDERLINE HIGH 
C0474551|T034||LNC|HAEMATOCRIT - BORDERLINE LOW 
C0474551|T034||LNC|HAEMATOCRIT - BORDERLINE LOW
C0474551|T034||LNC|HEMATOCRIT - BORDERLINE LOW
C0474551|T034||LNC|HEMATOCRIT - BORDERLINE LOW 
C2004297|T034||LNC|FINDING OF HEMATOCRIT - PACKED CELL VOLUME LEVEL
C2004297|T034||LNC|FINDING OF HAEMATOCRIT - PACKED CELL VOLUME LEVEL
C2004297|T034||LNC|HEMATOCRIT - PCV
C2004297|T034||LNC|HEMATOCRIT - P.C.V
C2004297|T034||LNC|HAEMATOCRIT - PCV
C2004297|T034||LNC|HAEMATOCRIT - P.C.V
C2004297|T034||LNC|HAEMATOCRIT - PCV LEVEL
C2004297|T034||LNC|HEMATOCRIT - PCV LEVEL
C2004297|T034||LNC|FINDING OF HEMATOCRIT - PACKED CELL VOLUME LEVEL 
C2004297|T034||LNC|HAEMATOCRIT - PCV LEVEL - FINDING
C2004297|T034||LNC|HEMATOCRIT - PCV LEVEL - FINDING
C1443990|T034||LNC|STABLE HAEMATOCRIT
C1443990|T034||LNC|STABLE HEMATOCRIT 
C1443990|T034||LNC|STABLE HEMATOCRIT
C0878707|T034||LNC|PRECIPITOUS DROP IN HEMATOCRIT
C0878707|T034||LNC|PRECIPITOUS DROP IN HEMATOCRIT 
C0878707|T034||LNC|DROP, HEMATOCRIT, PRECIP
C0878707|T034||LNC|PRECIPITOUS DROP IN HAEMATOCRIT
C0878707|T034||LNC|PRECIPITOUS DROP IN HEMATOCRIT 
