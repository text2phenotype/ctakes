C0003289|T121||RXNORM|ANTIDEPRESSIVE AGENTS
C0003289|T121||RXNORM|ANTIDEPRESSIVE DRUGS
C0003289|T121||RXNORM|ANTIDEPRESSIVE MEDICATIONS
C0360105|T121||RXNORM|SELECTIVE SEROTONIN REUPTAKE INHIBITORS
C0360105|T121||RXNORM|SSRI
C0719199|T121|215928|RXNORM|CELEXA|CELEXA
C0162373|T121|58827|RXNORM|PROZAC|PROZAC
C0376414|T121|114228|RXNORM|PAXIL|PAXIL
C0284660|T121|82728|RXNORM|ZOLOFT|ZOLOFT
C0678176|T121|196498|RXNORM|NEURONTIN|NEURONTIN
C0657912|T121|187832|RXNORM|PREGABALIN|PREGABALIN
C1570232|T121|593441|RXNORM|LYRICA|LYRICA
C0074393|T121|36437|RXNORM|SERTRALINE|SERTRALINE
C0074393|T121|36437|RXNORM|1-NAPHTHALENAMINE,1,2,3,4-TETRAHYDRO-4-(3,4-DICHLOROPHENYL)-N-METHYL-, (1S-CIS)-|SERTRALINE
C0074393|T121|36437|RXNORM|SERTRALINE [CHEMICAL/INGREDIENT]|SERTRALINE
C0074393|T121|36437|RXNORM|SERTRALINE |SERTRALINE
C0074393|T121|36437|RXNORM|SERTRALINE |SERTRALINE
C0078569|T121|39786|RXNORM|VENLAFAXINE|VENLAFAXINE
C0078569|T121|39786|RXNORM|ANTIDEPRESSANTS VENLAFAXINE|VENLAFAXINE
C0078569|T121|39786|RXNORM|VENLAFAXINE |VENLAFAXINE
C0078569|T121|39786|RXNORM|1-(2-(DIMETHYLAMINO)-1-(4-METHOXYPHENYL)ETHYL)CYCLOHEXANOL|VENLAFAXINE
C0078569|T121|39786|RXNORM|VENLAFAXINE [CHEMICAL/INGREDIENT]|VENLAFAXINE
C0078569|T121|39786|RXNORM|VENLAFAXINE |VENLAFAXINE
C0078569|T121|39786|RXNORM|VENLAFAXINE |VENLAFAXINE
C0078569|T121|39786|RXNORM|VNF|VENLAFAXINE
C0003290|T121||RXNORM|AGENTS, TRICYCLIC ANTIDEPRESSIVE
C0003290|T121||RXNORM|ANTIDEPRESSIVE AGENTS, TRICYCLIC
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSANT
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSANTS
C0003290|T121||RXNORM|DRUGS, TRICYCLIC ANTIDEPRESSANT
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSANT DRUGS
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSANTS 
C0003290|T121||RXNORM|[CN601] TRICYCLIC ANTIDEPRESSANTS
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSIVE AGENTS
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSANT DRUG
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSANT DRUG 
C0003290|T121||RXNORM|ANTIDEPRESSANTS, TRICYCLIC
C0003290|T121||RXNORM|ANTIDEPRESSANT DRUGS, TRICYCLIC
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSANT 
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSANT 
C0003290|T121||RXNORM|TRICYCLIC ANTIDEPRESSANT, NOS
C0016365|T121|4493|RXNORM|FLUOXETINE|FLUOXETINE
C0016365|T121|4493|RXNORM|BENZENEPROPANAMINE, N-METHYL-GAMMA-(4-(TRIFLUOROMETHYL)PHENOXY)-, (+-)-|FLUOXETINE
C0016365|T121|4493|RXNORM|N-METHYL-GAMMA-(4-(TRIFLUOROMETHYL) -PHENOXY)-BENZENEPROPANAMINE|FLUOXETINE
C0016365|T121|4493|RXNORM|FLUOXETIN|FLUOXETINE
C0016365|T121|4493|RXNORM|N-METHYL-GAMMA-(4-(TRIFLUOROMETHYL)PHENOXY)BENZENEPROPANAMINE|FLUOXETINE
C0016365|T121|4493|RXNORM|FLUOXETINE [CHEMICAL/INGREDIENT]|FLUOXETINE
C0016365|T121|4493|RXNORM|FLUOXETINE |FLUOXETINE
C0016365|T121|4493|RXNORM|FLUOXETINE |FLUOXETINE
C0016365|T121|4493|RXNORM|FLUOX|FLUOXETINE
C0031392|T121|8123|RXNORM|2 PHENETHYLHYDRAZINE|PHENELZINE
C0031392|T121|8123|RXNORM|PHENELZINE|PHENELZINE
C0031392|T121|8123|RXNORM|BETA PHENYLETHYLHYDRAZINE|PHENELZINE
C0031392|T121|8123|RXNORM|HYDRAZINE, (2-PHENYLETHYL)-|PHENELZINE
C0031392|T121|8123|RXNORM|FENELZIN|PHENELZINE
C0031392|T121|8123|RXNORM|BETA-PHENYLETHYLHYDRAZINE|PHENELZINE
C0031392|T121|8123|RXNORM|PHENETHYLHYDRAZINE|PHENELZINE
C0031392|T121|8123|RXNORM|PHENELZINE [CHEMICAL/INGREDIENT]|PHENELZINE
C0031392|T121|8123|RXNORM|2-PHENETHYLHYDRAZINE|PHENELZINE
C0031392|T121|8123|RXNORM|ANTIDEPRESSANTS PHENELZINE|PHENELZINE
C0031392|T121|8123|RXNORM|PHENELZINE |PHENELZINE
C0031392|T121|8123|RXNORM|MAOI - PHENELZINE|PHENELZINE
C0031392|T121|8123|RXNORM|PHENELZINE |PHENELZINE
C0031392|T121|8123|RXNORM|PHENELZINE |PHENELZINE
C0085208|T121|42347|RXNORM|BUPROPION|BUPROPION
C0085208|T121|42347|RXNORM|1-PROPANONE, 1-(3-CHLOROPHENYL)-2-((1,1-DIMETHYLETHYL)AMINO)-|BUPROPION
C0085208|T121|42347|RXNORM|AMFEBUTAMONE|BUPROPION
C0085208|T121|42347|RXNORM|BUPROPION |BUPROPION
C0085208|T121|42347|RXNORM|(+-)-1-(3-CHLOROPHENYL)-2-((1,1-DIMETHYLETHYL)AMINO)-1-PROPANONE|BUPROPION
C0085208|T121|42347|RXNORM|BUPROPION [CHEMICAL/INGREDIENT]|BUPROPION
C0085208|T121|42347|RXNORM|AMFEBUTAMON|BUPROPION
C0085208|T121|42347|RXNORM|BUPROPION |BUPROPION
C0085208|T121|42347|RXNORM|BUPROPION |BUPROPION
C0085208|T121|42347|RXNORM|BUP|BUPROPION
C0085208|T121|42347|RXNORM|BUPROPION [DUP] |BUPROPION
C0070122|T121|32937|RXNORM|PAROXETINE|PAROXETINE
C0070122|T121|32937|RXNORM|PIPERIDINE, 3-((1,3-BENZODIOXOL-5-YLOXY)METHYL)-4-(4-FLUOROPHENYL)-, (3S-TRANS)-|PAROXETINE
C0070122|T121|32937|RXNORM|(-)-TRANS-4-(P-FLUOROPHENYL)-3-((3,4-(METHYLENEDIOXY)PHENOXY)METHYL)PIPERIDINE|PAROXETINE
C0070122|T121|32937|RXNORM|(-)-(3S,4R)-4-(P-FLUOROPHENYL)-3-((3,4-(METHYLENEDIOXY)PHENOXY)METHYL)PIPERIDINE|PAROXETINE
C0070122|T121|32937|RXNORM|PAROXETINE [CHEMICAL/INGREDIENT]|PAROXETINE
C0070122|T121|32937|RXNORM|PAROXETINE |PAROXETINE
C0070122|T121|32937|RXNORM|PAROXETINE |PAROXETINE
C0008845|T121|2556|RXNORM|CITALOPRAM|CITALOPRAM
C0008845|T121|2556|RXNORM|5-ISOBENZOFURANCARBONITRILE, 1-(3-(DIMETHYLAMINO)PROPYL)-1-(4-FLUOROPHENYL)-1,3-DIHYDRO-|CITALOPRAM
C0008845|T121|2556|RXNORM|CYTALOPRAM|CITALOPRAM
C0008845|T121|2556|RXNORM|CITALOPRAM [CHEMICAL/INGREDIENT]|CITALOPRAM
C0008845|T121|2556|RXNORM|NITALAPRAM|CITALOPRAM
C0008845|T121|2556|RXNORM|1,3-DIHYDRO-1-(3-(DIMETHYLAMINO)PROPYL)-1-(4-FLUOROPHENYL)-5-ISOBENZOFURANCARBONITRILE|CITALOPRAM
C0008845|T121|2556|RXNORM|CITALOPRAM |CITALOPRAM
C0008845|T121|2556|RXNORM|CITALOPRAM |CITALOPRAM
C0085228|T121|42355|RXNORM|FLUVOXAMINE|FLUVOXAMINE
C0085228|T121|42355|RXNORM|1-PENTANONE, 5-METHOXY-1-(4-(TRIFLUOROMETHYL)PHENYL)-, O-(2-AMINOETHYL)OXIME, (E)-|FLUVOXAMINE
C0085228|T121|42355|RXNORM|FLUVOXAMINE [CHEMICAL/INGREDIENT]|FLUVOXAMINE
C0085228|T121|42355|RXNORM|FLUVOXAMINE |FLUVOXAMINE
C0085228|T121|42355|RXNORM|FLUVOXAMINE |FLUVOXAMINE
C0085228|T121|42355|RXNORM|FLUOXAMINE|FLUVOXAMINE
C0004962|T121|1361|RXNORM|BENACTYZINE|BENACTYZINE
C0004962|T121|1361|RXNORM|BENZENEACETIC ACID, ALPHA-HYDROXY-ALPHA-PHENYL-, 2-(DIETHYLAMINO)ETHYL ESTER|BENACTYZINE
C0004962|T121|1361|RXNORM|BENACTYZINE [CHEMICAL/INGREDIENT]|BENACTYZINE
C0004962|T121|1361|RXNORM|BENACTYZINE |BENACTYZINE
C0009035|T121||RXNORM|CLORGYLINE
C0009035|T121||RXNORM|2-PROPYN-1-AMINE, N-(3-(2,4-DICHLOROPHENOXY)PROPYL)-N-METHYL-
C0009035|T121||RXNORM|CLORGILINE
C0009035|T121||RXNORM|CLORGYLINE [CHEMICAL/INGREDIENT]
C0009035|T121||RXNORM|CLORGILIN
C0009035|T121||RXNORM|CHLORGYLINE
C0011064|T121|3116|RXNORM|DEANOL|DEANOL
C0011064|T121|3116|RXNORM|ETHANOL, 2-(DIMETHYLAMINO)-|DEANOL
C0011064|T121|3116|RXNORM|N,N DIMETHYL 2 HYDROXYETHYLAMINE|DEANOL
C0011064|T121|3116|RXNORM|DIMETHYLETHANOLAMINE|DEANOL
C0011064|T121|3116|RXNORM|DIMETHYL ETHANOLAMINE|DEANOL
C0011064|T121|3116|RXNORM|PARASYMPATHOMIMETICS DEANOL|DEANOL
C0011064|T121|3116|RXNORM|DEANOL |DEANOL
C0011064|T121|3116|RXNORM|N,N-DIMETHYL-N-(2-HYDROXYETHYL)AMINE|DEANOL
C0011064|T121|3116|RXNORM|2-DIMETHYLAMINOETHANOL|DEANOL
C0011064|T121|3116|RXNORM|DIMETHYLAMINOETHANOL|DEANOL
C0011064|T121|3116|RXNORM|DEMANYL|DEANOL
C0011064|T121|3116|RXNORM|DEMANOL|DEANOL
C0011064|T121|3116|RXNORM|N,N-DIMETHYL-2-HYDROXYETHYLAMINE|DEANOL
C0011064|T121|3116|RXNORM|N,N-DIMETHYLETHANOLAMINE|DEANOL
C0011064|T121|3116|RXNORM|DEANOL [CHEMICAL/INGREDIENT]|DEANOL
C0011064|T121|3116|RXNORM|DIMETHYL ETHANOLAMINE |DEANOL
C0011064|T121|3116|RXNORM|DEANOL |DEANOL
C0011064|T121|3116|RXNORM|2 DIMETHYLAMINOETHANOL|DEANOL
C0022059|T121|5981|RXNORM|IPRONIAZID|IPRONIAZID
C0022059|T121|5981|RXNORM|4-PYRIDINECARBOXYLIC ACID, 2-(1-METHYLETHYL)HYDRAZIDE|IPRONIAZID
C0022059|T121|5981|RXNORM|IPRAZID|IPRONIAZID
C0022059|T121|5981|RXNORM|IPRONIAZID [CHEMICAL/INGREDIENT]|IPRONIAZID
C0022059|T121|5981|RXNORM|1-ISONICOTINOYL-2-ISOPROPYLHYDRAZINE|IPRONIAZID
C0022059|T121|5981|RXNORM|IPRONIAZID |IPRONIAZID
C0022059|T121|5981|RXNORM|IPRONIAZID |IPRONIAZID
C0022154|T121|6011|RXNORM|ISOCARBOXAZID|ISOCARBOXAZID
C0022154|T121|6011|RXNORM|3-ISOXAZOLECARBOXYLIC ACID, 5-METHYL-, 2-(PHENYLMETHYL)HYDRAZIDE|ISOCARBOXAZID
C0022154|T121|6011|RXNORM|RO 5-0831|ISOCARBOXAZID
C0022154|T121|6011|RXNORM|ISOCARBOXAZID |ISOCARBOXAZID
C0022154|T121|6011|RXNORM|ISOCARBOXAZID [CHEMICAL/INGREDIENT]|ISOCARBOXAZID
C0022154|T121|6011|RXNORM|MAOI - ISOCARBOXAZID|ISOCARBOXAZID
C0022154|T121|6011|RXNORM|ISOCARBOXAZID |ISOCARBOXAZID
C0022154|T121|6011|RXNORM|ISOCARBOXAZID |ISOCARBOXAZID
C0027999|T121|7394|RXNORM|NIALAMIDE|NIALAMIDE
C0027999|T121|7394|RXNORM|4-PYRIDINECARBOXYLIC ACID, 2-(3-OXO-3-((PHENYLMETHYL)AMINO)PROPYL)HYDRAZIDE|NIALAMIDE
C0027999|T121|7394|RXNORM|1-(2-(BENZYLCARBAMOYL)ETHYL)-2-ISONICOTINOYLHYDRAZINE|NIALAMIDE
C0027999|T121|7394|RXNORM|NIALAMIDE [CHEMICAL/INGREDIENT]|NIALAMIDE
C0027999|T121|7394|RXNORM|NIALAMIDE |NIALAMIDE
C0032036|T121|8373|RXNORM|PIZOTYLINE|PIZOTYLINE
C0032036|T121|8373|RXNORM|PIPERIDINE, 4-(9,10-DIHYDRO-4H-BENZO(4,5)CYCLOHEPTA(1,2-B)THIEN-4-YLIDENE)-1-METHYL-|PIZOTYLINE
C0032036|T121|8373|RXNORM|PIZOTYLINE PRODUCT|PIZOTYLINE
C0032036|T121|8373|RXNORM|PIZOTIFEN|PIZOTYLINE
C0032036|T121|8373|RXNORM|PIZOTYLINE [CHEMICAL/INGREDIENT]|PIZOTYLINE
C0032036|T121|8373|RXNORM|4-(9,10-DIHYDRO-4H-BENZO(4,5)CYCLOHEPTA(1,2-B)THIEN-4-YLIDENE)-1-METHYLPIPERIDINE|PIZOTYLINE
C0032036|T121|8373|RXNORM|PIZOTIFEN PRODUCT |PIZOTYLINE
C0032036|T121|8373|RXNORM|PIZOTIFEN PRODUCT|PIZOTYLINE
C0032036|T121|8373|RXNORM|PIZOTIFEN |PIZOTYLINE
C0032036|T121|8373|RXNORM|PIZOTIFEN |PIZOTYLINE
C0040778|T121|10734|RXNORM|TRANYLCYPROMINE|TRANYLCYPROMINE
C0040778|T121|10734|RXNORM|TRANS 2 PHENYLCYCLOPROPYLAMINE|TRANYLCYPROMINE
C0040778|T121|10734|RXNORM|CYCLOPROPANAMINE, 2-PHENYL-, TRANS-(+-)-|TRANYLCYPROMINE
C0040778|T121|10734|RXNORM|TRANYLCYPROMINE [CHEMICAL/INGREDIENT]|TRANYLCYPROMINE
C0040778|T121|10734|RXNORM|TRANS-2-PHENYLCYCLOPROPYLAMINE|TRANYLCYPROMINE
C0040778|T121|10734|RXNORM|ANTIDEPRESSANTS TRANYLCYPROMINE|TRANYLCYPROMINE
C0040778|T121|10734|RXNORM|TRANYLCYPROMINE |TRANYLCYPROMINE
C0040778|T121|10734|RXNORM|MAOI - TRANYLCYPROMINE|TRANYLCYPROMINE
C0040778|T121|10734|RXNORM|TRANYLCYPROMINE |TRANYLCYPROMINE
C0040778|T121|10734|RXNORM|TRANYLCYPROMINE |TRANYLCYPROMINE
C0206486|T121||RXNORM|LITHIUM COMPOUNDS
C0206486|T121||RXNORM|COMPOUNDS, LITHIUM
C0206486|T121||RXNORM|LITHIUM CPDS
C0206486|T121||RXNORM|LITHIUM COMPOUNDS [CHEMICAL/INGREDIENT]
C0206486|T121||RXNORM|LITHIUM COMPOUND 
C0206486|T121||RXNORM|LITHIUM COMPOUND
C0206486|T121||RXNORM|LITHIUM COMPOUND, NOS
C0073561|T121||RXNORM|ROLIPRAM
C0073561|T121||RXNORM|PYRROLIDONE, 4-(3-CYCLOPENTYLOXY-4-METHOXYPHENYL)-2-
C0073561|T121||RXNORM|ROLIPRAM [CHEMICAL/INGREDIENT]
C0073561|T121||RXNORM|(+/-)-ROLIPRAM
C0073561|T121||RXNORM|(R,S)-ROLIPRAM
C0066673|T121|30121|RXNORM|MOCLOBEMIDE|MOCLOBEMIDE
C0066673|T121|30121|RXNORM|MOCLOBEMIDE |MOCLOBEMIDE
C0066673|T121|30121|RXNORM|BENZAMIDE, 4-CHLORO-N-(2-(4-MORPHOLINYL)ETHYL)-|MOCLOBEMIDE
C0066673|T121|30121|RXNORM|MOCLOBAMIDE|MOCLOBEMIDE
C0066673|T121|30121|RXNORM|MOCLOBEMIDE [CHEMICAL/INGREDIENT]|MOCLOBEMIDE
C0066673|T121|30121|RXNORM|P-CHLORO-N-(2-MORPHOLINOETHYL)BENZAMIDE|MOCLOBEMIDE
C0066673|T121|30121|RXNORM|MOCLOBEMIDE |MOCLOBEMIDE
C0066673|T121|30121|RXNORM|MOCLOBEMIDE |MOCLOBEMIDE
C0242905|T121||RXNORM|AGENTS, SECOND-GENERATION ANTIDEPRESSIVE
C0242905|T121||RXNORM|ANTIDEPRESSIVE AGENTS, SECOND GENERATION
C0242905|T121||RXNORM|ANTIDEPRESSIVE AGENTS, SECOND-GENERATION
C0242905|T121||RXNORM|ANTIDEPRESSIVE DRUGS, SECOND GENERATION
C0242905|T121||RXNORM|DRUGS, SECOND-GENERATION ANTIDEPRESSIVE
C0242905|T121||RXNORM|SECOND GENERATION ANTIDEPRESSIVE AGENTS
C0242905|T121||RXNORM|SECOND-GENERATION ANTIDEPRESSIVE DRUGS
C0242905|T121||RXNORM|SECOND-GENERATION ANTIDEPRESSIVE AGENTS
C0242905|T121||RXNORM|ANTIDEPRESSANTS, ATYPICAL
C0242905|T121||RXNORM|ANTIDEPRESSIVE DRUGS, SECOND-GENERATION
C0242905|T121||RXNORM|ATYPICAL ANTIDEPRESSANTS
C0085217|T121|42351|RXNORM|CARBONATE, LITHIUM|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|CARBONATE, DILITHIUM|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|CARBONIC ACID, DILITHIUM SALT|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE |LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE [CHEMICAL/INGREDIENT]|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|DILITHIUM CARBONATE|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE PREPARATION|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE |LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE |LITHIUM CARBONATE
C0003289|T121||RXNORM|AGENTS, ANTIDEPRESSIVE
C0003289|T121||RXNORM|ANTIDEPRESSIVE AGENTS
C0003289|T121||RXNORM|ANTIDEPRESSANT
C0003289|T121||RXNORM|DRUGS, ANTIDEPRESSANT
C0003289|T121||RXNORM|ANTIDEPRESSANTS
C0003289|T121||RXNORM|ANTIDEPRESSANTS 
C0003289|T121||RXNORM|ANTIDEPRESSIVE
C0003289|T121||RXNORM|ANTIDEPRESSIVE AGENT [TC]
C0003289|T121||RXNORM|[CN600] ANTIDEPRESSANTS
C0003289|T121||RXNORM|ANTIDEPRESSIVE AGENT
C0003289|T121||RXNORM|ANTIDEPRESSANT DRUG
C0003289|T121||RXNORM|ANTIDEPRESSANT DRUG 
C0003289|T121||RXNORM|ANTIDEPRESSANT DRUGS
C0003289|T121||RXNORM|ANTIDEPRESSANT 
C0003289|T121||RXNORM|ANTIDEPRESSANT 
C0003289|T121||RXNORM|ANTIDEPRESSANT, NOS
C0003289|T121||RXNORM|ANTIDEPRESSANT AGENT
C1337136|T121||RXNORM|L-METHYLFOLATE
C1337136|T121||RXNORM|L-METHYLFOLATE 
C1337136|T121||RXNORM|L-METHYLFOLATE 
C1337136|T121||RXNORM|6(S)-5-METHYLTETRAHYDROFOLATE
C1337136|T121||RXNORM|L-METHYL FOLIC ACID
C1337136|T121||RXNORM|5-MTHF
C1337136|T121||RXNORM|5-METHYLTETRAHYDROFOLATE
C1337136|T121||RXNORM|L-GLUTAMIC ACID, N-(4-(((2-AMINO-1,4,5,6,7,8-HEXAHYDRO-5- METHYL-4-OXO-6-PTERIDINYL)METHYL)AMINO)BENZOYL)-
C1337136|T121||RXNORM|L-METHYLTETRAHYDROFOLATE
C1337136|T121||RXNORM|5-METHYL TERAHYDROFOLIC ACID
C2316497|T121|993548|RXNORM|BUPROPION HYDROBROMIDE |BUPROPION HYDROBROMIDE
C2316497|T121|993548|RXNORM|BUPROPION HYDROBROMIDE|BUPROPION HYDROBROMIDE
C2316497|T121|993548|RXNORM|1-PROPANONE, 1-(3-CHLOROPHENYL)-2-((1,1-DIMETHYLETHYL)AMINO)-, HYDROBROMIDE|BUPROPION HYDROBROMIDE
C2316497|T121|993548|RXNORM|BUPROPION HBR|BUPROPION HYDROBROMIDE
C2316497|T121|993548|RXNORM|BUPROPION HYDROBROMIDE |BUPROPION HYDROBROMIDE
C0215087|T121||RXNORM|N,N-DIMETHYL-ALPHA-(2-(1-NAPHTHALENYLOXY)ETHYL)BENZENEMETHANAMINE
C0215087|T121||RXNORM|DAPOXETINE
C0215087|T121||RXNORM|BENZENEMETHANAMINE, N,N-DIMETHYL-ALPHA-(2-(1-NAPHTHALENYLOXY)ETHYL)-, (+)-
C0215087|T121||RXNORM|DAPOXETINE 
C2699580|T121||RXNORM|DELFAPRAZINE
C2699584|T121||RXNORM|DELUCEMINE HYDROCHLORIDE
C0957739|T121||RXNORM|ECLANAMINE MALEATE
C0068785|T121||RXNORM|3-(2-METHOXYPHENOXY)-N-METHYL-3-PHENYLPROPYLAMINE
C0068785|T121||RXNORM|3-(O-METHOXYPHENOXY)-N-METHYL-3-PHENYLPROPYLAMINE
C0068785|T121||RXNORM|N-METHYL-GAMMA-(2-METHYLPHENOXY)PHENYLPROPANOLAMINE
C0068785|T121||RXNORM|NISOXETINE
C2698483|T121||RXNORM|NOMELIDINE
C2698505|T121||RXNORM|NOXIPTILINE
C0069709|T121||RXNORM|2-(3-TRIFLUOROMETHYLPHENYL)-4-ISOPROPYLTETRAHYDRO-1,4-OXAZINE
C0069709|T121||RXNORM|4-(1-METHYLETHYL)-2-(3-(TRIFLUOROMETHYL)PHENYL)MORPHOLINE
C0069709|T121||RXNORM|OXAFLOZANE
C2699092|T121||RXNORM|ROFELODINE
C2699289|T121||RXNORM|SEPROXETINE
C0069628|T121||RXNORM|1,2,3,4-TETRAHYDRO-2-METHYL-9H-DIBENZO(3,4-6,7)CYCLOHEPTA(1,2-C)PYRIDINE
C0069628|T121||RXNORM|13B,4A-CARBA-MIANSERIN
C0069628|T121||RXNORM|SETIPTILINE
C2699506|T121||RXNORM|SPIROXEPIN
C0144486|T121||RXNORM|TALSUPRAM
C2699901|T121||RXNORM|TEBATIZOLE
C0075496|T121||RXNORM|SUFOXAZINE
C0075496|T121||RXNORM|TENILOXAZINE
C2699942|T121||RXNORM|TIENOPRAMINE
C0607615|T121||RXNORM|TETRAHYDRO-6-(PHENOXYMETHYL)-2H-1,3-OXAZINE-2- THIONE
C0607615|T121||RXNORM|TIFEMOXONE
C0538554|T121||RXNORM|(S)-2-(((7-FLUORO-4-INDANYL)OXY)METHYL)MORPHOLINE MONOHYDROCHLORIDE
C0538554|T121||RXNORM|LUBAZODONE HYDROCHLORIDE
C0055961|T121||RXNORM|(E)-1-(4- CHLOROPHENYL)-5-METHOXY-1-PENTANONE O-(2- AMINOETHYL)OXIME, (E)-2-BUTENEDIOATE (1:1)
C0055961|T121||RXNORM|CLOVOXAMINE
C0600943|T121||RXNORM|COTRIPTYLINE
C0600943|T121||RXNORM|10,11-DIHYDRO-5H-DIBENZO(A,D)CYCLOHEPTENYLIDENE-5-3-DIMETHYLAMINO-2-PROPANONE
C0663336|T121||RXNORM|ALPHA-2-PROPENYL BENZENEETHANAMINE
C0663336|T121||RXNORM|ALETAMINE
C0663336|T121||RXNORM|ALFETADRINE
C0663336|T121||RXNORM|ALFETAMIN
C0663336|T121||RXNORM|ALFETAMINE
C0663336|T121||RXNORM|ALPHA-ALLYL-PHENETHYLAMIN
C0663336|T121||RXNORM|ALPHA-ALLYLPHENETHYLAMINE
C1702222|T121||RXNORM|BEFETUPITANT
C2698343|T121||RXNORM|BELOXEPIN
C0621294|T121||RXNORM|CLOBAMINE MESYLATE
C0621294|T121||RXNORM|CILOBAMINE MESYLATE
C2699221|T121||RXNORM|CINFENINE
C0047305|T121||RXNORM|3-CHLORO-5-(3-(4-PIPERIDINO-4- CARBAMOYLPIPERIDINO)PROPYL)-10,11-DIHYDRO-5H- DIBENZ(B,F)AZEPINE DIHYDROCHLORIDE MONOHYDRATE
C0047305|T121||RXNORM|3-CHLOROCARPIPRAMINE
C0047305|T121||RXNORM|CLOCAPRAMINE
C2699359|T121||RXNORM|CLODAZON
C2699360|T121||RXNORM|CLODAZON HYDROCHLORIDE
C0615823|T121||RXNORM|5H-DIBENXO(A,D)CYCLOHEPTEN-5-ONE O-(2-(METHYLAMINO)ETHYL)OXIME
C0615823|T121||RXNORM|DEMEXIPTILINE
C0044643|T121||RXNORM|5-(3-(DIMETHYLAMINO)PROPYL)-5H-DIBENZ- (B,F)AZEPINE
C0044643|T121||RXNORM|DEPRAMINE
C0044643|T121||RXNORM|10,11-DEHYDROIMIPRAMINE
C2699611|T121||RXNORM|DEXIMAFEN
C0131796|T121||RXNORM|(2-(2-DIMETHYLAMINO)ETHYL)-2-PHENYL-3,4-DIHYDRO-1(2H)-NAPHTHALENONE
C0131796|T121||RXNORM|(S)-NAFENODONE
C0131796|T121||RXNORM|NAFENODONE
C0131796|T121||RXNORM|DEXNAFENODONE
C0057877|T121||RXNORM|DICLOFENSINE
C0543452|T121|142133|RXNORM|HYDROCHLORIDE, DOTHIEPIN|DOTHIEPIN HYDROCHLORIDE
C0543452|T121|142133|RXNORM|DOTHIEPIN HYDROCHLORIDE |DOTHIEPIN HYDROCHLORIDE
C0543452|T121|142133|RXNORM|DOTHIEPIN HYDROCHLORIDE|DOTHIEPIN HYDROCHLORIDE
C0543452|T121|142133|RXNORM|ANTIDEPRESSANTS DOTHIEPIN HYDROCHLORIDE|DOTHIEPIN HYDROCHLORIDE
C0543452|T121|142133|RXNORM|DOTHIEPIN HYDROCHLORIDE |DOTHIEPIN HYDROCHLORIDE
C0543452|T121|142133|RXNORM|DOTHIEPIN HYDROCHLORIDE |DOTHIEPIN HYDROCHLORIDE
C0543452|T121|142133|RXNORM|DOSULEPIN HYDROCHLORIDE|DOTHIEPIN HYDROCHLORIDE
C2699861|T121||RXNORM|ELANZEPINE
C2697947|T121||RXNORM|LUBAZODONE
C1533126|T121|588250|RXNORM|CYCLOPROPANECARBOXAMIDE, 2-(AMINOMETHYL)-N,N-DIETHYL-1-PHENYL-, CIS-(+-)-|MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN|MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN |MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN |MILNACIPRAN
C1533126|T121|588250|RXNORM|MIDALCIPRAN|MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN [CHEMICAL/INGREDIENT]|MILNACIPRAN
C1533126|T121|588250|RXNORM|ANTIDEPRESSANTS SNRI MILNACIPRAN|MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN |MILNACIPRAN
C0066529|T121|30003|RXNORM|MILNACIPRAN HYDROCHLORIDE|MILNACIPRAN HYDROCHLORIDE
C0066529|T121|30003|RXNORM|MILNACIPRAN HYDROCHLORIDE |MILNACIPRAN HYDROCHLORIDE
C0066529|T121|30003|RXNORM|MILNACIPRAN HYDROCHLORIDE |MILNACIPRAN HYDROCHLORIDE
C0066529|T121|30003|RXNORM|MILNACIPRAN HYDROCHLORIDE |MILNACIPRAN HYDROCHLORIDE
C0066529|T121|30003|RXNORM|1-PHENYL-1-DIETHYLAMINOCARBONYL-2-AMINOMETHYLCYCLOPROPANE HCL|MILNACIPRAN HYDROCHLORIDE
C2698946|T121||RXNORM|RADAFAXINE HYDROCHLORIDE
C2699361|T121||RXNORM|CLODAZON HYDROCHLORIDE ANHYDROUS
C0052237|T121||RXNORM|1,3,4,14B-TETRAHYDRO-2-METHYL-10H-PYRAZINO-(1,2-A)PYRROLO(2,1-C)(1,4)BENZODIAZEPINE
C0052237|T121||RXNORM|APTAZAPINE
C0052237|T121||RXNORM|2H,10H-PARAZINO(1,2-A)PYRROLO(2,1-C)(1,4)BENZODIAZEPINE,1,3,4,14B-TETRAHYDRO-2-METHYL-
C2698177|T121||RXNORM|APTAZAPINE MALEATE
C2698177|T121||RXNORM|2H,10H-PYRAZINO(1,2-A)PYRROLO(2,1-C)(1,4)BENZODIAZEPINE, 1,3,4,14B-TETRAHYDRO-2-METHYL-, (+-)-, (Z)-2-BUTENEDIOATE (1:1)
C2698082|T121||RXNORM|2H- INDOL-2-ONE, L,3-DIHYDRO-3-METHYL-3-[3-(METHYLAMINO)-PROPYL]-L-PHENYL-
C2698082|T121||RXNORM|AMEDALIN
C2607957|T121||RXNORM|BENZAPRINOXIDE
C2607957|T121||RXNORM|1-PROPANAMINE, 3-(1-CHLORO-5H-DIBENZO(A,D)CYCLOHEPTEN-5-YLIDENE)-N,N-DIMETHYL-, N-OXIDE
C2698511|T121||RXNORM|BIPENAMOL
C0054270|T121|19895|RXNORM|10,11-DIHYDRO-N,N,BETA-TRIMETHYL-5H-DIBENZO(A,D) CYCLOHEPTANE-5-PROPYLAMINE|BUTRIPTYLINE
C0054270|T121|19895|RXNORM|BUTRIPTYLENE|BUTRIPTYLINE
C0054270|T121|19895|RXNORM|BUTRIPTYLINE|BUTRIPTYLINE
C0054270|T121|19895|RXNORM|10,11-DIHYDRO-N,N,BETA-TRIMETHYL-5H-DIBENZO(A,D)CYCLOHEPTENE-5-PROPYLAMINE|BUTRIPTYLINE
C0054270|T121|19895|RXNORM|BUTRIPTYLINE |BUTRIPTYLINE
C0054270|T121|19895|RXNORM|BUTRIPTYLINE |BUTRIPTYLINE
C1108795|T121|324004|RXNORM|BUTRIPTYLINE HYDROCHLORIDE |BUTRIPTYLINE HYDROCHLORIDE
C1108795|T121|324004|RXNORM|ANTIDEPRESSANTS BUTRIPTYLINE HYDROCHLORIDE|BUTRIPTYLINE HYDROCHLORIDE
C1108795|T121|324004|RXNORM|BUTRIPTYLINE HYDROCHLORIDE|BUTRIPTYLINE HYDROCHLORIDE
C1108795|T121|324004|RXNORM|5H-DIBENZO(A,D)CYCLOHEPTENE-5-PROPYLAMINE, 10,11-DIHYDRO-N,N,BETA-TRIMETHYL-, HYDROCHLORIDE, DL-|BUTRIPTYLINE HYDROCHLORIDE
C2699208|T121||RXNORM|CICLOPRAMINE
C2699208|T121||RXNORM|2,3,7,8-TETRAHYDRO-3-METHYLAMINO-1H-CHINO(1,8-A,B)BENZAZEPIN
C2699343|T121||RXNORM|3-(3-CHLORPHENYL)-1-(DIMETHYLAMINO)-3-PHENYL-2-PROPANOL
C2699343|T121||RXNORM|CLEMEPROL
C2699343|T121||RXNORM|M-CHLORO-ALPHA-((DIMETHYLAMINO)METHYL)-BETA-PHENYLPHENETYL ALCOHOL
C0055708|T121||RXNORM|CICLAZINDOL
C0055708|T121||RXNORM|PYRIMIDO(1,2-A)INDOL-10-OL, 10-(3-CHLOROPHENYL)-2,3,4,10-TETRAHYDRO-
C0951496|T121||RXNORM|3-(2-MORPHOLINO-ETHYLAMINO)-4-METHYL-6-PHENYL PYRIDAZINE, DIHYDROCHLORIDE
C0951496|T121||RXNORM|N-(4-METHYL-6-PHENYL-3-PYRIDAZINYL)-4-MORPHOLINEETHANAMINE DIHYDROCHLORIDE
C0951496|T121||RXNORM|MINAPRINE HYDROCHLORIDE
C0951496|T121||RXNORM|MORPHOLINE, 4-(2-((4-METHYL-6-PHENYL-3-PYRIDAZINYL)AMINO)ETHYL)-, DIHYDROCHLORIDE
C0951496|T121||RXNORM|MINAPRINE DIHYDROCHLORIDE
C0959897|T121||RXNORM|ALPHA-ALLYLPHENETHYLAMINE HYDROCHLORIDE
C0959897|T121||RXNORM|ALFETAMINE HYDROCHLORIDE
C0959897|T121||RXNORM|ALETAMINE HYDROCHLORIDE
C0959897|T121||RXNORM|BENZENEETHANAMINE, ALPHA-2-PROPENYL-, HYDROCHLORIDE
C0970823|T121||RXNORM|DAPOXETINE HYDROCHLORIDE
C0621295|T121||RXNORM|2-(3,4-DICHLOROPHENYL)-3-((1-METHYLETHYL)AMINO)BICYCLO(2.2.2)OCTAN-2-OL MONOMETHANESULFONATE
C0621295|T121||RXNORM|CILOBAMINE
C2825651|T121||RXNORM|AMEDALIN HYDROCHLORIDE
C0953067|T121|1311672|RXNORM|INDELOXAZINE HYDROCHLORIDE|INDELOXAZINE HYDROCHLORIDE
C2825652|T121||RXNORM|DILOPETINE
C0635054|T121||RXNORM|ECLANAMINE
C2825653|T121||RXNORM|NUCLOTIXENE
C2825654|T121||RXNORM|ADOPRAZINE
C2825655|T121||RXNORM|CAPROXAMINE
C0063456|T121|1311673|RXNORM|2-(7-INDENYLOXYMETHYL)MORPHOLINE|INDELOXAZINE
C0063456|T121|1311673|RXNORM|INDELOXAZINE|INDELOXAZINE
C0063456|T121|1311673|RXNORM|MORPHOLINE, 2-((1H-INDEN-7-YLOXY)METHYL)-|INDELOXAZINE
C0054826|T121|20342|RXNORM|5-(3-(4-PIPERIDINO-4-CARBAMOYLPIPERIDINO)PROPYL)- 10,11-DIHYDRO-5(H)-DIBENZ(B,F)AZEPINE|CARPIPRAMINE
C0054826|T121|20342|RXNORM|CARBADIPIMIDINE|CARPIPRAMINE
C0054826|T121|20342|RXNORM|CARPIPRAMINE|CARPIPRAMINE
C2825656|T121||RXNORM|FENMETOZOLE HYDROCHLORIDE
C0060175|T121||RXNORM|FENMETAZOLE
C0060175|T121||RXNORM|FENMETOZOLE
C0060175|T121||RXNORM|2-((3,4-DICHLOROPHENOXY)METHYL)-2-IMIDAZOLINE
C0056704|T121||RXNORM|2,3,4,9-TETRAHYDRO-N,N-DIMETHYL-1H-CARBAZOL-3- AMINE
C0056704|T121||RXNORM|2,3,4,9-TETRAHYDRO-N,N-DIMETHYL-1H-CARBAZOLE-3-AMINE
C0056704|T121||RXNORM|3-(DIMETHYLAMINO)-1,2,3,4-TETRAHYDROCARBAZOLE
C0056704|T121||RXNORM|CYCLINDOLE
C2825657|T121||RXNORM|LOSINDOLE
C0058199|T121||RXNORM|DIMETACRINE
C0058199|T121||RXNORM|DIMETHACRINE
C0058199|T121||RXNORM|ISOTONIL
C0058199|T121||RXNORM|ISTONIL
C2825658|T121||RXNORM|LOMEVACTONE
C2825659|T121||RXNORM|FENMETRAMIDE
C2826066|T121||RXNORM|MARIPTILINE
C2826066|T121||RXNORM|1A,10B-DIHYDRODIBENZO(A,E)CYCLOPROPA(C)CYCLOHEPTEN-6(1H)-ONE O-(2-AMINOETHYL)OXIME
C0886642|T121|1298842|RXNORM|PAROXETINE HYDROCHLORIDE HEMIHYDRATE|PAROXETINE HYDROCHLORIDE, HEMIHYDRATE
C0886642|T121|1298842|RXNORM|PAROXETINE HYDROCHLORIDE, HEMIHYDRATE|PAROXETINE HYDROCHLORIDE, HEMIHYDRATE
C0886642|T121|1298842|RXNORM|HEMIHYDRATE, PAROXETINE HYDROCHLORIDE|PAROXETINE HYDROCHLORIDE, HEMIHYDRATE
C0886642|T121|1298842|RXNORM|HYDROCHLORIDE HEMIHYDRATE, PAROXETINE|PAROXETINE HYDROCHLORIDE, HEMIHYDRATE
C0886642|T121|1298842|RXNORM|HYDROCHLORIDE, HEMIHYDRATE PAROXETINE|PAROXETINE HYDROCHLORIDE, HEMIHYDRATE
C0886642|T121|1298842|RXNORM|HEMIHYDRATE PAROXETINE HYDROCHLORIDE|PAROXETINE HYDROCHLORIDE, HEMIHYDRATE
C0886642|T121|1298842|RXNORM|(3S-TRANS)-3-[(1,3-BENZODIOXOL-5-YLOXY)METHYL]-4-(4-FLUOROPHENYL)PIPERIDINE HYDROCHLORIDE HEMIHYDRATE|PAROXETINE HYDROCHLORIDE, HEMIHYDRATE
C2827083|T121||RXNORM|AZEPINDOLE
C2827119|T121||RXNORM|CUTAMESINE
C2827119|T121||RXNORM|1-(2-(3,4-DIMETHOXYPHENYL)ETHYL)-4-(3-PHENYLPROPYL)PIPERAZINE
C2827129|T121||RXNORM|DAZADROL
C2827129|T121||RXNORM|2-PYRIDINEMETHANOL, ALPHA-(4-CHLOROPHENYL)-ALPHA-(4,5-DIHYDRO-1H-IMIDAZOL-2-YL)-
C2827129|T121||RXNORM|ALPHA-(P-CHLOROPHENYL)-ALPHA-2-IMIDAZOLIN-2-YL-2-PYRIDINEMETHANOL
C2827130|T121||RXNORM|DAZADROL MALEATE
C2827154|T121||RXNORM|FANTRIDONE
C0963192|T121||RXNORM|(+-)-TRANS-3-(3,4-DICHLOROPHENYL)-N-METHYL-1-INDANAMINE
C0963192|T121||RXNORM|INDATRALINE
C0611882|T121||RXNORM|5-(3-(DIMETHYLAMINO)PROPYL)-5,11-DIHYDRO-10H-DIBENZ(B,F)AZEPIN-10-ONE
C0611882|T121||RXNORM|KETIMIPRAMINE
C0611882|T121||RXNORM|KETIPRAMINE
C0611882|T121||RXNORM|1-ALPHA-4,5-ALPHA-H-TROPANIUM, 3-ALPHA-HYDROXY-8-(P-PHENYLPHENACYL)-, (-)-TROPATE
C2827221|T121||RXNORM|KETIPRAMINE FUMARATE
C0125662|T121||RXNORM|LEVOPROTILINE
C0125662|T121||RXNORM|HYDROXYMAPROTILIN, (+R)-ISOMER
C1565971|T121||RXNORM|TALOPRAM
C1565971|T121||RXNORM|1,3-DIHYDRO-N,3,3-TRIMETHYL-1-PHENYLBENZO(C)FURAN-1-PROPANAMINE
C0025912|T121|6929|RXNORM|MIANSERIN|MIANSERIN
C0025912|T121|6929|RXNORM|DIBENZO(C,F)PYRAZINO(1,2-A)AZEPINE, 1,2,3,4,10,14B-HEXAHYDRO-2-METHYL-|MIANSERIN
C0025912|T121|6929|RXNORM|MIANSERIN [CHEMICAL/INGREDIENT]|MIANSERIN
C0025912|T121|6929|RXNORM|1,2,3,4,10,14B-HEXAHYDRO-2-METHYLDIBENZO(C,F)-PYRAZINO(1,2-A)AZEPINE|MIANSERIN
C0025912|T121|6929|RXNORM|ANTIDEPRESSANTS MIANSERIN|MIANSERIN
C0025912|T121|6929|RXNORM|MIANSERIN |MIANSERIN
C0025912|T121|6929|RXNORM|MIANSERIN |MIANSERIN
C0025912|T121|6929|RXNORM|MIANSERIN |MIANSERIN
C0700456|T121|203127|RXNORM|HYDROCHLORIDE, MIANSERIN|MIANSERIN HYDROCHLORIDE
C0700456|T121|203127|RXNORM|MIANSERIN HYDROCHLORIDE |MIANSERIN HYDROCHLORIDE
C0700456|T121|203127|RXNORM|MIANSERIN HYDROCHLORIDE|MIANSERIN HYDROCHLORIDE
C0700456|T121|203127|RXNORM|ANTIDEPRESSANTS MIANSERIN HYDROCHLORIDE|MIANSERIN HYDROCHLORIDE
C0700456|T121|203127|RXNORM|DIBENZO(C,F)PYRAZINO(1,2-A)AZEPINE, 1,2,3,4,10,14B-HEXAHYDRO-2-METHYL-, MONOHYDROCHLORIDE|MIANSERIN HYDROCHLORIDE
C0700456|T121|203127|RXNORM|1,2,3,4,10,14B-HEXAHYDRO-2-METHYLDIBENZO(C,F)-PYRAZINO(1,2-A)AZEPINE MONOHYDROCHLORIDE|MIANSERIN HYDROCHLORIDE
C0700456|T121|203127|RXNORM|MONOHYDROCHLORIDE, MIANSERIN|MIANSERIN HYDROCHLORIDE
C0700456|T121|203127|RXNORM|MIANSERIN MONOHYDROCHLORIDE|MIANSERIN HYDROCHLORIDE
C0700456|T121|203127|RXNORM|MIANSERIN HYDROCHLORIDE |MIANSERIN HYDROCHLORIDE
C0700456|T121|203127|RXNORM|MIANSERIN HYDROCHLORIDE |MIANSERIN HYDROCHLORIDE
C0031974|T121||RXNORM|PIPRADROL
C0031974|T121||RXNORM|PYRIDROL
C0031974|T121||RXNORM|PIPRADOL
C0031974|T121||RXNORM|PIPRADROL 
C0020934|T121|5691|RXNORM|IMIPRAMINE|IMIPRAMINE
C0020934|T121|5691|RXNORM|5H-DIBENZ(B,F)AZEPINE-5-PROPANAMINE, 10,11-DIHYDRO-N,N-DIMETHYL-|IMIPRAMINE
C0020934|T121|5691|RXNORM|IMIDOBENZYLE|IMIPRAMINE
C0020934|T121|5691|RXNORM|IMIPRAMINE [CHEMICAL/INGREDIENT]|IMIPRAMINE
C0020934|T121|5691|RXNORM|IMIZIN|IMIPRAMINE
C0020934|T121|5691|RXNORM|NORCHLORIMIPRAMINE|IMIPRAMINE
C0020934|T121|5691|RXNORM|IMIPRAMINE |IMIPRAMINE
C0020934|T121|5691|RXNORM|IMIPRAMINE |IMIPRAMINE
C0026388|T121|7019|RXNORM|MOLINDONE|MOLINDONE
C0026388|T121|7019|RXNORM|4H-INDOL-4-ONE, 3-ETHYL-1,5,6,7-TETRAHYDRO-2-METHYL-5-(4-MORPHOLINYLMETHYL)-|MOLINDONE
C0026388|T121|7019|RXNORM|MOLINDONE [CHEMICAL/INGREDIENT]|MOLINDONE
C0026388|T121|7019|RXNORM|MOLINDONE |MOLINDONE
C0026388|T121|7019|RXNORM|MOLINDONE |MOLINDONE
C0040805|T121|10737|RXNORM|TRAZODONE|TRAZODONE
C0040805|T121|10737|RXNORM|1,2,4-TRIAZOLO(4,3-A)PYRIDIN-3(2H)-ONE, 2-(3-(4-(3-CHLOROPHENYL)-1-PIPERAZINYL)PROPYL)-|TRAZODONE
C0040805|T121|10737|RXNORM|TRADOZONE|TRAZODONE
C0040805|T121|10737|RXNORM|SEARLE BRAND OF TRAZODONE HYDROCHLORIDE|TRAZODONE
C0040805|T121|10737|RXNORM|TRAZODONE [CHEMICAL/INGREDIENT]|TRAZODONE
C0040805|T121|10737|RXNORM|TRAZODONE |TRAZODONE
C0040805|T121|10737|RXNORM|ANTIDEPRESSANTS TRAZODONE|TRAZODONE
C0040805|T121|10737|RXNORM|TRAZODONE |TRAZODONE
C0040805|T121|10737|RXNORM|TRAZODONE |TRAZODONE
C0038803|T121|10239|RXNORM|SULPIRIDE|SULPIRIDE
C0038803|T121|10239|RXNORM|BENZAMIDE, 5-(AMINOSULFONYL)-N-((1-ETHYL-2-PYRROLIDINYL)METHYL)-2-METHOXY-|SULPIRIDE
C0038803|T121|10239|RXNORM|SULPIRIDE [CHEMICAL/INGREDIENT]|SULPIRIDE
C0038803|T121|10239|RXNORM|SULPERIDE|SULPIRIDE
C0038803|T121|10239|RXNORM|N-((1-ETHYL-2-PYRROLIDINYL)METHYL)-5-SULFAMOYL-O-ANISAMIDE|SULPIRIDE
C0038803|T121|10239|RXNORM|ANTIDEPRESSANTS SULPIRIDE|SULPIRIDE
C0038803|T121|10239|RXNORM|SULPIRIDE |SULPIRIDE
C0038803|T121|10239|RXNORM|SULPIRIDE |SULPIRIDE
C0038803|T121|10239|RXNORM|SULPIRIDE |SULPIRIDE
C0043479|T121||RXNORM|ZIMELDINE
C0043479|T121||RXNORM|2-PROPEN-1-AMINE, 3-(4-BROMOPHENYL)-N,N-DIMETHYL-3-(3-PYRIDINYL)-, (Z)-
C0043479|T121||RXNORM|ZIMELDINE [CHEMICAL/INGREDIENT]
C0043479|T121||RXNORM|ZIMELIDIN
C0043479|T121||RXNORM|ZIMELIDINE
C0043479|T121||RXNORM|ZIMELDINE 
C0028420|T121|7531|RXNORM|NORTRIPTYLINE|NORTRIPTYLINE
C0028420|T121|7531|RXNORM|1-PROPANAMINE, 3-(10,11-DIHYDRO-5H-DIBENZO(A,D)CYCLOHEPTEN-5-YLIDENE)-N-METHYL-|NORTRIPTYLINE
C0028420|T121|7531|RXNORM|DESITRIPTYLINE|NORTRIPTYLINE
C0028420|T121|7531|RXNORM|NORTRIPTYLINE [CHEMICAL/INGREDIENT]|NORTRIPTYLINE
C0028420|T121|7531|RXNORM|DESMETHYLAMITRIPTYLIN|NORTRIPTYLINE
C0028420|T121|7531|RXNORM|NORTRIPTYLINE |NORTRIPTYLINE
C0028420|T121|7531|RXNORM|NORTRYPTYLINE|NORTRIPTYLINE
C0028420|T121|7531|RXNORM|NORTRIPTYLINE |NORTRIPTYLINE
C0028420|T121|7531|RXNORM|NTPL|NORTRIPTYLINE
C0025810|T121|6901|RXNORM|METHYLPHENIDATE|METHYLPHENIDATE
C0025810|T121|6901|RXNORM|2-PIPERIDINEACETIC ACID, ALPHA-PHENYL-, METHYL ESTER|METHYLPHENIDATE
C0025810|T121|6901|RXNORM|ALPHA-PHENYL-2-PIPERIDINEACETIC ACID METHYL ESTER|METHYLPHENIDATE
C0025810|T121|6901|RXNORM|METHYLPHENIDATE [CHEMICAL/INGREDIENT]|METHYLPHENIDATE
C0025810|T121|6901|RXNORM|METHYLPHENIDATE |METHYLPHENIDATE
C0025810|T121|6901|RXNORM|CNS STIMULANTS METHYLPHENIDATE|METHYLPHENIDATE
C0025810|T121|6901|RXNORM|METHYLPHENIDATE |METHYLPHENIDATE
C0025810|T121|6901|RXNORM|METHYLPHENIDATE |METHYLPHENIDATE
C0025810|T121|6901|RXNORM|D-METHYLPHENIDATE|METHYLPHENIDATE
C0031407|T121||RXNORM|BETA-PHENYLISOPROPYLHYDRAZINE
C0031407|T121||RXNORM|PHENIPRAZINE
C0031407|T121||RXNORM|HYDRAZINE, (1-METHYL-2-PHENYLETHYL)-
C0013085|T121|3638|RXNORM|DOXEPIN|DOXEPIN
C0013085|T121|3638|RXNORM|1-PROPANAMINE, 3-DIBENZ(B,E)OXEPIN-11(6H)-YLIDENE-N,N-DIMETHYL-|DOXEPIN
C0013085|T121|3638|RXNORM|DOXEPIN [CHEMICAL/INGREDIENT]|DOXEPIN
C0013085|T121|3638|RXNORM|DOXEPIN |DOXEPIN
C0013085|T121|3638|RXNORM|DOXEPIN |DOXEPIN
C0024778|T121|6646|RXNORM|MAPROTILINE|MAPROTILINE
C0024778|T121|6646|RXNORM|9,10-ETHANOANTHRACENE-9(10H)-PROPANAMINE, N-METHYL-|MAPROTILINE
C0024778|T121|6646|RXNORM|MAPROTILIN|MAPROTILINE
C0024778|T121|6646|RXNORM|N-METHYL-9,10-ETHANOANTHRACENE-9(10H)-PROPYLAMINE|MAPROTILINE
C0024778|T121|6646|RXNORM|DIBENCYCLADINE|MAPROTILINE
C0024778|T121|6646|RXNORM|MAPROTILINE [CHEMICAL/INGREDIENT]|MAPROTILINE
C0024778|T121|6646|RXNORM|MAPROTILINE |MAPROTILINE
C0024778|T121|6646|RXNORM|MAPROTILINE |MAPROTILINE
C0011685|T121|3247|RXNORM|DESIPRAMINE|DESIPRAMINE
C0011685|T121|3247|RXNORM|5H-DIBENZ(B,F)AZEPINE-5-PROPANAMINE, 10,11-DIHYDRO-N-METHYL-|DESIPRAMINE
C0011685|T121|3247|RXNORM|DESMETHYLIMIPRAMINE|DESIPRAMINE
C0011685|T121|3247|RXNORM|DEMETHYLIMIPRAMINE|DESIPRAMINE
C0011685|T121|3247|RXNORM|DESIPRAMINE [CHEMICAL/INGREDIENT]|DESIPRAMINE
C0011685|T121|3247|RXNORM|ANTIDEPRESSANTS DESIPRAMINE|DESIPRAMINE
C0011685|T121|3247|RXNORM|DESIPRAMINE |DESIPRAMINE
C0011685|T121|3247|RXNORM|DESIPRAMINE |DESIPRAMINE
C0011685|T121|3247|RXNORM|DESIPRAMINE |DESIPRAMINE
C0009010|T121|2597|RXNORM|CLOMIPRAMINE|CLOMIPRAMINE
C0009010|T121|2597|RXNORM|5H-DIBENZ(B,F)AZEPINE-5-PROPANAMINE, 3-CHLORO-10,11-DIHYDRO-N,N-DIMETHYL-|CLOMIPRAMINE
C0009010|T121|2597|RXNORM|3-CHLORO-5-(3-(DIMETHYLAMINO)PROPYL)-10,11-DIHYDRO-5H-DIBENZ(B,F)AZEPINE|CLOMIPRAMINE
C0009010|T121|2597|RXNORM|CHLOMIPRAMINE|CLOMIPRAMINE
C0009010|T121|2597|RXNORM|CLOMIPRAMINE [CHEMICAL/INGREDIENT]|CLOMIPRAMINE
C0009010|T121|2597|RXNORM|CHLORIMIPRAMINE|CLOMIPRAMINE
C0009010|T121|2597|RXNORM|CLOMIPRAMINE |CLOMIPRAMINE
C0009010|T121|2597|RXNORM|CLOMIPRAMINE |CLOMIPRAMINE
C0028277|T121|7500|RXNORM|NOMIFENSINE|NOMIFENSINE
C0028277|T121|7500|RXNORM|8-ISOQUINOLINAMINE, 1,2,3,4-TETRAHYDRO-2-METHYL-4-PHENYL-|NOMIFENSINE
C0028277|T121|7500|RXNORM|NOMIFENSIN|NOMIFENSINE
C0028277|T121|7500|RXNORM|LINAMIPHEN|NOMIFENSINE
C0028277|T121|7500|RXNORM|NOMIFENSINE [CHEMICAL/INGREDIENT]|NOMIFENSINE
C0009170|T121|2653|RXNORM|COCAINE|COCAINE
C0009170|T121|2653|RXNORM|8-AZABICYCLO(3.2.1)OCTANE-2-CARBOXYLIC ACID, 3-(BENZOYLOXY)-8-METHYL-, METHYL ESTER, (1R-(EXO,EXO))-|COCAINE
C0009170|T121|2653|RXNORM|(1R,2R,3S,5S)-2-METHOXYCARBONYLTROPAN-3-YL BENZOATE|COCAINE
C0009170|T121|2653|RXNORM|COCAINE [CHEMICAL/INGREDIENT]|COCAINE
C0009170|T121|2653|RXNORM|COCAINE (SCHEDULE I SUBSTANCE)|COCAINE
C0009170|T121|2653|RXNORM|BLOW|COCAINE
C0009170|T121|2653|RXNORM|SNOW|COCAINE
C0009170|T121|2653|RXNORM|COKE|COCAINE
C0009170|T121|2653|RXNORM|COCA|COCAINE
C0009170|T121|2653|RXNORM|COCAINE PRODUCT|COCAINE
C0009170|T121|2653|RXNORM|COCAINE |COCAINE
C0009170|T121|2653|RXNORM|COCAINE |COCAINE
C0355303|T121||RXNORM|COMPOUND ANTIDEPRESSANTS
C0355303|T121||RXNORM|COMPOUND ANTIDEPRESSANTS 
C0355303|T121||RXNORM|COMPOUND ANTIDEPRESSANTS 
C0771200|T121|235988|RXNORM|VENLAFAXINE HYDROCHLORIDE|VENLAFAXINE HYDROCHLORIDE
C0771200|T121|235988|RXNORM|VENLAFAXINE HYDROCHLORIDE |VENLAFAXINE HYDROCHLORIDE
C0771200|T121|235988|RXNORM|ANTIDEPRESSANTS VENLAFAXINE HYDROCHLORIDE|VENLAFAXINE HYDROCHLORIDE
C0771200|T121|235988|RXNORM|HYDROCHLORIDE, VENLAFAXINE|VENLAFAXINE HYDROCHLORIDE
C0771200|T121|235988|RXNORM|CYCLOHEXANOL, 1-(2-(DIMETHYLAMINO)-1-(4-METHOXYPHENYL)ETHYL)-, HYDROCHLORIDE|VENLAFAXINE HYDROCHLORIDE
C0771200|T121|235988|RXNORM|VENLAFAXINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|VENLAFAXINE HYDROCHLORIDE
C0771200|T121|235988|RXNORM|1-(2-(DIMETHYLAMINO)-1-(4-METHOXYPHENYL)ETHYL)CYCLOHEXANOL HCL|VENLAFAXINE HYDROCHLORIDE
C0771200|T121|235988|RXNORM|VENLAFAXINE HYDROCHLORIDE |VENLAFAXINE HYDROCHLORIDE
C0771200|T121|235988|RXNORM|VENLAFAXINE HYDROCHLORIDE |VENLAFAXINE HYDROCHLORIDE
C0600356|T121||RXNORM|H 102 09
C0600356|T121||RXNORM|H10209
C0600356|T121||RXNORM|H-102-09
C0002600|T121|704|RXNORM|AMITRIPTYLINE|AMITRIPTYLINE
C0002600|T121|704|RXNORM|1-PROPANAMINE, 3-(10,11-DIHYDRO-5H-DIBENZO(A,D)CYCLOHEPTEN-5-YLIDENE)-N,N-DIMETHYL-|AMITRIPTYLINE
C0002600|T121|704|RXNORM|AMITRIPTYLINE [CHEMICAL/INGREDIENT]|AMITRIPTYLINE
C0002600|T121|704|RXNORM|AMITRIPTYLINE |AMITRIPTYLINE
C0002600|T121|704|RXNORM|AMITRIPTYLINE |AMITRIPTYLINE
C0678139|T121|196471|RXNORM|SEROXAT|SEROXAT
C0591911|T121|152158|RXNORM|OPTIMAX|OPTIMAX
C0591911|T121|152158|RXNORM|MERCK BRAND OF TRYPTOPHAN|OPTIMAX
C0360105|T121||RXNORM|SELECTIVE SEROTONIN REUPTAKE INHIBITORS 
C0360105|T121||RXNORM|SEROTONIN REUPTAKE INHIBITORS
C0360105|T121||RXNORM|SELECTIVE SEROTONIN REUPTAKE INHIBITORS (SSRIS)
C0360105|T121||RXNORM|SELECTIVE SEROTONIN REUPTAKE INHIBITORS
C0360105|T121||RXNORM|SELECTIVE SEROTONIN REUPTAKE INHIBITOR
C0360105|T121||RXNORM|SSRIS
C0360105|T121||RXNORM|SSRI
C0360105|T121||RXNORM|SSRI - SELECTIVE SEROTONIN RE-UPTAKE INHIBITOR
C0360105|T121||RXNORM|SELECTIVE SEROTONIN RE-UPTAKE INHIBITOR
C0360105|T121||RXNORM|SELECTIVE SEROTONIN RE-UPTAKE INHIBITOR 
C0360105|T121||RXNORM|SELECTIVE SEROTONIN RE-UPTAKE INHIBITOR 
C0543469|T121|142143|RXNORM|VILOXAZINE HYDROCHLORIDE |VILOXAZINE HYDROCHLORIDE
C0543469|T121|142143|RXNORM|ANTIDEPRESSANTS VILOXAZINE HYDROCHLORIDE|VILOXAZINE HYDROCHLORIDE
C0543469|T121|142143|RXNORM|VILOXAZINE HYDROCHLORIDE|VILOXAZINE HYDROCHLORIDE
C0543469|T121|142143|RXNORM|VILOXAZINE HYDROCHLORIDE |VILOXAZINE HYDROCHLORIDE
C0543469|T121|142143|RXNORM|VILOXAZINE HYDROCHLORIDE |VILOXAZINE HYDROCHLORIDE
C1529955|T121||RXNORM|ANTIDEPRESSANTS DIBENZEPIN HYDROCHLORIDE
C1529955|T121||RXNORM|DIBENZEPIN HYDROCHLORIDE
C1529955|T121||RXNORM|DIBENZEPIN HYDROCHLORIDE 
C0877847|T121|262302|RXNORM|MALEATE, NOMIFENSINE|NOMIFENSINE MALEATE
C0877847|T121|262302|RXNORM|NOMIFENSINE MALEATE |NOMIFENSINE MALEATE
C0877847|T121|262302|RXNORM|NOMIFENSINE MALEATE|NOMIFENSINE MALEATE
C0877847|T121|262302|RXNORM|NOMIFENSINE MALEATE (1:1)|NOMIFENSINE MALEATE
C2079567|T121|814600|RXNORM|PERPHENAZINE + NORTRIPTYLINE |NORTRIPTYLINE / PERPHENAZINE
C2079567|T121|814600|RXNORM|PERPHENAZINE + NORTRIPTYLINE|NORTRIPTYLINE / PERPHENAZINE
C2079567|T121|814600|RXNORM|NORTRIPTYLINE / PERPHENAZINE|NORTRIPTYLINE / PERPHENAZINE
C2189302|T121|816810|RXNORM|VERALIPRIDE + BROMAZEPAM|BROMAZEPAM / VERALIPRIDE
C2189302|T121|816810|RXNORM|VERALIPRIDE + BROMAZEPAM |BROMAZEPAM / VERALIPRIDE
C2189302|T121|816810|RXNORM|BROMAZEPAM / VERALIPRIDE|BROMAZEPAM / VERALIPRIDE
C0041056|T121|10834|RXNORM|TRIMIPRAMINE|TRIMIPRAMINE
C0041056|T121|10834|RXNORM|5H-DIBENZ(B,F)AZEPINE-5-PROPANAMINE, 10,11-DIHYDRO-N,N,BETA-TRIMETHYL-|TRIMIPRAMINE
C0041056|T121|10834|RXNORM|TRIMIPRAMINE |TRIMIPRAMINE
C0041056|T121|10834|RXNORM|TRIMEPRIMINE|TRIMIPRAMINE
C0041056|T121|10834|RXNORM|10,11 DIHYDRO-N,N,BETA-TRIMETHYL-5H-DIBENZ(B,F)AZEPINE-5-PROPANAMINE|TRIMIPRAMINE
C0041056|T121|10834|RXNORM|TRIMIPRAMINE [CHEMICAL/INGREDIENT]|TRIMIPRAMINE
C0041056|T121|10834|RXNORM|TRIMIPRAMINE |TRIMIPRAMINE
C0041056|T121|10834|RXNORM|TRIMIPRAMINE |TRIMIPRAMINE
C0036579|T121|9639|RXNORM|SELEGILINE|SELEGILINE
C0036579|T121|9639|RXNORM|BENZENEETHANAMINE, N,ALPHA-DIMETHYL-N-2-PROPYNYL-, (R)-|SELEGILINE
C0036579|T121|9639|RXNORM|SELEGILINE |SELEGILINE
C0036579|T121|9639|RXNORM|(-)-DEPRENIL|SELEGILINE
C0036579|T121|9639|RXNORM|(-)-PHENYLISOPROPYLMETHYLPROPYNYLAMINE|SELEGILINE
C0036579|T121|9639|RXNORM|L-DEPRENYL|SELEGILINE
C0036579|T121|9639|RXNORM|SELEGILINE [CHEMICAL/INGREDIENT]|SELEGILINE
C0036579|T121|9639|RXNORM|SELEGYLINE|SELEGILINE
C0036579|T121|9639|RXNORM|SELEGILINE, (R)-ISOMER|SELEGILINE
C0036579|T121|9639|RXNORM|(-)-SELEGILINE|SELEGILINE
C0036579|T121|9639|RXNORM|SELEGILINE |SELEGILINE
C0036579|T121|9639|RXNORM|SELEGILINE |SELEGILINE
C1579361|T121||RXNORM|SNRI ANTIDEPRESSANTS
C1579361|T121||RXNORM|SEROTONIN AND NOREPINEPHRINE REUPTAKE INHIBITORS (SNRIS)
C1579361|T121||RXNORM|SEROTONIN AND NOREPINEPHRINE REUPTAKE INHIBITORS 
C1579361|T121||RXNORM|ANTIDEPRESSANTS SEROTONIN AND NOREPINEPHRINE REUPTAKE INHIBITORS
C1579361|T121||RXNORM|SEROTONIN AND NOREPINEPHRINE REUPTAKE INHIBITORS
C1579361|T121||RXNORM|SEROTONIN AND NORADRENALINE REUPTAKE INHIBITORS
C1579361|T121||RXNORM|NRIS AND SSRIS
C1579361|T121||RXNORM|SEROTONIN AND NOREPINEPHRINE UPTAKE INHIBITORS
C1579361|T121||RXNORM|SSRIS AND NRIS
C1579361|T121||RXNORM|SEROTONIN AND NORADRENALINE UPTAKE INHIBITORS
C1579361|T121||RXNORM|SNRIS
C2064901|T121||RXNORM|BENACTYZINE HYDROCHLORIDE + MEPROBAMATE
C2064901|T121||RXNORM|BENACTYZINE HYDROCHLORIDE + MEPROBAMATE 
C1616289|T121||RXNORM|HYDROGENATED ERGOT ALKALOIDS 
C1616289|T121||RXNORM|HYDROGENATED ERGOT ALKALOIDS
C1616289|T121||RXNORM|ERGOT ALKALOIDS, HYDROGENATED
C1616289|T121||RXNORM|HYDROGENATED ERGOT ALKALOID
C1616289|T121||RXNORM|ALKALOIDS, HYDROGENATED ERGOT
C0026457|T121||RXNORM|INHIBITOR, MONOAMINE OXIDASE
C0026457|T121||RXNORM|INHIBITORS, MONOAMINE OXIDASE
C0026457|T121||RXNORM|MONOAMINE OXIDASE INHIBITORS
C0026457|T121||RXNORM|MAO INHIBITOR
C0026457|T121||RXNORM|INHIBITORS, MAO
C0026457|T121||RXNORM|MAO INHIB
C0026457|T121||RXNORM|MONOAMINE OXIDASE INHIB
C0026457|T121||RXNORM|MONOAMINE OXIDASE INHIBITOR
C0026457|T121||RXNORM|MONOAMINE OXIDASE INHIBITORS 
C0026457|T121||RXNORM|MAO INHIBITORS
C0026457|T121||RXNORM|MONOAMINE OXIDASE INHIBITORS (MAOI)
C0026457|T121||RXNORM|MAOI
C0026457|T121||RXNORM|MONOAMINE OXIDASE--INHIBITORS
C0026457|T121||RXNORM|MAOI - MONOAMINE-OXIDASE INHIBITOR
C0026457|T121||RXNORM|MONOAMINE-OXIDASE INHIBITOR
C0026457|T121||RXNORM|MONOAMINE OXIDASE INHIBITOR 
C0026457|T121||RXNORM|MONOAMINE OXIDASE INHIBITOR 
C0026457|T121||RXNORM|MONOAMINE OXIDASE INHIBITOR, NOS
C0026457|T121||RXNORM|AMINE OXIDASE INHIBITORS
C1302097|T121||RXNORM|PERPHENAZINE + AMITRIPTYLINE HYDROCHLORIDE 
C1302097|T121||RXNORM|PERPHENAZINE + AMITRIPTYLINE HYDROCHLORIDE
C1302097|T121||RXNORM|ANTIDEPRESSANTS PERPHENAZINE + AMITRIPTYLINE HCL
C1302097|T121||RXNORM|AMITRIPTYLINE HYDROCHLORIDE + PERPHENAZINE
C1302097|T121||RXNORM|AMITRIPTYLINE HYDROCHLORIDE + PERPHENAZINE 
C0002644|T121|722|RXNORM|AMOXAPINE|AMOXAPINE
C0002644|T121|722|RXNORM|DIBENZ(B,F)(1,4)OXAZEPINE, 2-CHLORO-11-(1-PIPERAZINYL)-|AMOXAPINE
C0002644|T121|722|RXNORM|AMOXAPINE |AMOXAPINE
C0002644|T121|722|RXNORM|AMOXAPINE [CHEMICAL/INGREDIENT]|AMOXAPINE
C0002644|T121|722|RXNORM|DESMETHYLLOXAPINE|AMOXAPINE
C0002644|T121|722|RXNORM|2-CHLORO-11-(1-PIPERAZINYL)DIBENZ(B,F)(1,4)OXAZEPINE|AMOXAPINE
C0002644|T121|722|RXNORM|AMOXAPINE - CHEMICAL|AMOXAPINE
C0002644|T121|722|RXNORM|AMOXAPINE - CHEMICAL |AMOXAPINE
C0002644|T121|722|RXNORM|AMOXAPINE |AMOXAPINE
C0002644|T121|722|RXNORM|AMOXAPINE |AMOXAPINE
C0049506|T121|15996|RXNORM|6-AZAMIANSERIN|MIRTAZAPINE
C0049506|T121|15996|RXNORM|PYRAZINO(2,1-A)PYRIDO(2,3-C)(2)BENZAZEPINE, 1,2,3,4,10,14B-HEXAHYDRO-2-METHYL-|MIRTAZAPINE
C0049506|T121|15996|RXNORM|MIRTAZAPINE|MIRTAZAPINE
C0049506|T121|15996|RXNORM|MIRTAZAPINE |MIRTAZAPINE
C0049506|T121|15996|RXNORM|MIRTAZAPINE [CHEMICAL/INGREDIENT]|MIRTAZAPINE
C0049506|T121|15996|RXNORM|MIRTAZAPINE |MIRTAZAPINE
C0049506|T121|15996|RXNORM|MIRTAZAPINE |MIRTAZAPINE
C1875508|T121||RXNORM|MONAMINE OXIDASE INHIBITOR ANTIDEPRESSANTS
C1875508|T121||RXNORM|[CN602] MONAMINE OXIDASE INHIBITOR ANTIDEPRESSANTS
C1579362|T121||RXNORM|ANTIDEPRESSANTS,OTHER
C1579362|T121||RXNORM|[CN609] ANTIDEPRESSANTS,OTHER
C2981302|T121||RXNORM|MO-1255
C2981302|T121||RXNORM|ENCYPRATE
C2981302|T121||RXNORM|CARBAMIC ACID, CYCLOPROPYL(PHENYLMETHYL)-, ETHYL ESTER
C2981302|T121||RXNORM|ETHYL N-BENZYLCYCLOPROPANECARBAMATE
C2981302|T121||RXNORM|A-19757
C2981303|T121||RXNORM|ESREBOXETINE SUCCINATE
C2981304|T121||RXNORM|FANTRIDONE HYDROCHLORIDE ANHYDROUS
C2981304|T121||RXNORM|5-(3-(DIMETHYLAMINO)PROPYL)-6(5H)-PHENANTHRIDINONE MONOHYDROCHLORIDE
C2981304|T121||RXNORM|6(5H)-PHENANTHRIDINONE, 5-(3-(DIMETHYLAMINO)PROPYL)-, MONOHYDROCHLORIDE
C0023961|T121|6465|RXNORM|LOFEPRAMINE|LOFEPRAMINE
C0023961|T121|6465|RXNORM|ETHANONE, 1-(4-CHLOROPHENYL)-2-((3-(10,11-DIHYDRO-5H-DIBENZ(B,F)AZEPIN-5-YL)PROPYL)METHYLAMINO)-|LOFEPRAMINE
C0023961|T121|6465|RXNORM|LOFEPRAMINE [CHEMICAL/INGREDIENT]|LOFEPRAMINE
C0023961|T121|6465|RXNORM|LOPRAMINE|LOFEPRAMINE
C0023961|T121|6465|RXNORM|4'-CHLORO-2-((3-(10,11-DIHYDRO-5H-DIBENZ(B,F)AZEPIN-5-YL)PROPYL)METHYLAMINO)ACETOPHENONE|LOFEPRAMINE
C0023961|T121|6465|RXNORM|LOFEPRAMINE |LOFEPRAMINE
C0023961|T121|6465|RXNORM|LOFEPRAMINE |LOFEPRAMINE
C0023330|T121|6294|RXNORM|HYDROCHLORIDE, LOFEPRAMINE|LOFEPRAMINE HYDROCHLORIDE
C0023330|T121|6294|RXNORM|ANTIDEPRESSANTS LOFEPRAMINE HYDROCHLORIDE|LOFEPRAMINE HYDROCHLORIDE
C0023330|T121|6294|RXNORM|LOFEPRAMINE HYDROCHLORIDE|LOFEPRAMINE HYDROCHLORIDE
C0023330|T121|6294|RXNORM|LOFEPRAMINE HYDROCHLORIDE |LOFEPRAMINE HYDROCHLORIDE
C0023330|T121|6294|RXNORM|LOFEPRAMINE HYDROCHLORIDE |LOFEPRAMINE HYDROCHLORIDE
C0023330|T121|6294|RXNORM|4'-CHLORO-2-((3-(10,11-DIHYDRO-5H-DIBENZ(B, F)AZEPIN-5-YL)PROPYL)METHYLAMINO)ACETOPHENONE MONOHYDROCHLORIDE|LOFEPRAMINE HYDROCHLORIDE
C0023330|T121|6294|RXNORM|ETHANONE, 1-(4-CHLOROPHENYL)-2-((3-(10,11-DIHYDRO-5H-DIBENZ(B, F)AZEPIN-5-YL)PROPYL)METHYLAMINO)-, MONOHYDROCHLORIDE|LOFEPRAMINE HYDROCHLORIDE
C0066057|T121||RXNORM|15-METHYL-10-METHYLAMINO-10,11- DIHYDRODIBENZO(B,F)-AZEPINE
C0066057|T121||RXNORM|METAPRAMINE
C0066057|T121||RXNORM|15-METHYL-10-METHYLAMINO-10,11-DIHYDRODIBENZO(B,F)- AZEPINE
C0066057|T121||RXNORM|10,11-DIHYDRO-5-METHYL-10-(METHYLAMINO)-5H-DIBENZ(B,F)AZEPINE
C0029105|T121|7674|RXNORM|OPIPRAMOL|OPIPRAMOL
C0029105|T121|7674|RXNORM|1-PIPERAZINEETHANOL, 4-(3-(5H-DIBENZ(B,F)AZEPIN-5-YL)PROPYL)-|OPIPRAMOL
C0029105|T121|7674|RXNORM|OPIPRAMOL [CHEMICAL/INGREDIENT]|OPIPRAMOL
C2983799|T121||RXNORM|ORVEPITANT
C2983799|T121||RXNORM|1-PIPERIDINECARBOXAMIDE, N-[(1R)-1-[3,5-BIS(TRIFLUOROMETHYL)PHENYL]ETHYL]-2-(4-FLUORO-2-METHYLPHENYL)-4-[(8AS)-HEXAHYDRO-6-OXOPYRROLO[1,2-A]PYRAZIN-2(1H)-YL]-N-METHYL-, (2R,4S)-
C2983800|T121||RXNORM|GW823296B
C2983800|T121||RXNORM|ORVEPITANT MALEATE
C2983846|T121||RXNORM|MELITRACEN HYDROCHLORIDE
C2983846|T121||RXNORM|U 24,973A
C2983847|T121||RXNORM|MODALINE SULFATE
C2983847|T121||RXNORM|W 3207B
C2983848|T121||RXNORM|NAPRODOXIME
C2983849|T121||RXNORM|NEMIFITIDE
C2983850|T121||RXNORM|NITRAFUDAM
C2983851|T121||RXNORM|OMILOXETINE
C1530072|T121|1086769|RXNORM|VILAZODONE|VILAZODONE
C1530072|T121|1086769|RXNORM|5-{4-[4-(5-CYANO-1H-INDOL-3-YL)BUTYL]PIPERAZIN-1-YL}BENZOFURAN-2-CARBOXAMIDE|VILAZODONE
C1530072|T121|1086769|RXNORM|VILAZODONE |VILAZODONE
C1530072|T121|1086769|RXNORM|5-(4-(4-(5-CYANO-3-INDOLYL)BUTYL)-1-PIPERAZINYL)BENZOFURAN-2-CARBOXAMIDE|VILAZODONE
C2962546|T121|1086768|RXNORM|VILAZODONE HYDROCHLORIDE|VILAZODONE HYDROCHLORIDE
C2962546|T121|1086768|RXNORM|5-{4-[4-(5-CYANO-1H-INDOL-3-YL)BUTYL]PIPERAZIN-1-YL}BENZOFURAN-2-CARBOXAMIDE HYDROCHLORIDE|VILAZODONE HYDROCHLORIDE
C2962546|T121|1086768|RXNORM|ANTIDEPRESSANTS VILAZODONE|VILAZODONE HYDROCHLORIDE
C2962546|T121|1086768|RXNORM|VILAZODONE HCL |VILAZODONE HYDROCHLORIDE
C2962546|T121|1086768|RXNORM|VILAZODONE HCL|VILAZODONE HYDROCHLORIDE
C2962546|T121|1086768|RXNORM|VILAZODONE HYDROCHLORIDE |VILAZODONE HYDROCHLORIDE
C2962546|T121|1086768|RXNORM|HCL, VILAZODONE|VILAZODONE HYDROCHLORIDE
C2962546|T121|1086768|RXNORM|HYDROCHLORIDE, VILAZODONE|VILAZODONE HYDROCHLORIDE
C2962546|T121|1086768|RXNORM|2-BENZOFURANCARBOXAMIDE, 5-(4-(4-(5-CYANO-1H-INDOL-3-YL)BUTYL)-1-PIPERAZINYL)-, HYDROCHLORIDE (1:1)|VILAZODONE HYDROCHLORIDE
C2962546|T121|1086768|RXNORM|VILAZODONE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|VILAZODONE HYDROCHLORIDE
C2698285|T121||RXNORM|AZALOXAN
C0282270|T121|82062|RXNORM|HYDROCHLORIDE, OPIPRAMOL|OPIPRAMOL HYDROCHLORIDE
C0282270|T121|82062|RXNORM|OPIPRAMOL HYDROCHLORIDE|OPIPRAMOL HYDROCHLORIDE
C0282270|T121|82062|RXNORM|OPIPRAMOL DIHYDROCHLORIDE|OPIPRAMOL HYDROCHLORIDE
C0282270|T121|82062|RXNORM|4-(3-(5H-DIBENZ(B,F)AZEPIN-5-YL)PROPYL)-1-PIPERAZINEETHANOL DIHYDROCHLORIDE|OPIPRAMOL HYDROCHLORIDE
C0282270|T121|82062|RXNORM|1-PIPERAZINEETHANOL, 4-(3-(5H-DIBENZ(B,F)AZEPIN-5-YL)PROPYL)-, DIHYDROCHLORIDE|OPIPRAMOL HYDROCHLORIDE
C0732706|T121|226942|RXNORM|LITHIUM SUCCINATE 80 MG/ML TOPICAL CREAM|LITHIUM SUCCINATE 8 % TOPICAL CREAM
C0732706|T121|226942|RXNORM|LITHIUM SUCCINATE 8 % TOPICAL CREAM|LITHIUM SUCCINATE 8 % TOPICAL CREAM
C0732706|T121|226942|RXNORM|LITHIUM SUCCINATE 8% CREAM|LITHIUM SUCCINATE 8 % TOPICAL CREAM
C0732706|T121|226942|RXNORM|LITHIUM SUCCINATE 8% CREAM |LITHIUM SUCCINATE 8 % TOPICAL CREAM
C0732706|T121|226942|RXNORM|LITHIUM SUCCINATE 8% CREAM |LITHIUM SUCCINATE 8 % TOPICAL CREAM
C0013065|T121|3634|RXNORM|DOTHIEPIN|DOTHIEPIN
C0013065|T121|3634|RXNORM|1-PROPANAMINE, 3-DIBENZO(B,E)THIEPIN-11(6H)-YLIDENE-N,N-DIMETHYL-|DOTHIEPIN
C0013065|T121|3634|RXNORM|DOTHIEPIN [CHEMICAL/INGREDIENT]|DOTHIEPIN
C0013065|T121|3634|RXNORM|DOSULEPIN|DOTHIEPIN
C0013065|T121|3634|RXNORM|DOTHIEPIN |DOTHIEPIN
C0013065|T121|3634|RXNORM|DOTHIEPIN |DOTHIEPIN
C0013065|T121|3634|RXNORM|DOSULEPIN |DOTHIEPIN
C0973506|T121||RXNORM|OTHER ANTIDEPRESSANT DRUGS 
C0973506|T121||RXNORM|OTHER ANTIDEPRESSANT DRUGS
C0973506|T121||RXNORM|OTHER ANTIDEPRESSANT DRUGS 
C0693279|T121|993506|RXNORM|BUPROPION HCL 100MG SA TAB|BUPROPION HYDROCHLORIDE 100 MG EXTENDED RELEASE ORAL TABLET
C0693279|T121|993506|RXNORM|BUPROPION HCL 100MG TAB,SA|BUPROPION HYDROCHLORIDE 100 MG EXTENDED RELEASE ORAL TABLET
C0693279|T121|993506|RXNORM|BUPROPION HCL 100MG TAB,SA [VA PRODUCT]|BUPROPION HYDROCHLORIDE 100 MG EXTENDED RELEASE ORAL TABLET
C0693279|T121|993506|RXNORM|BUPROPION HYDROCHLORIDE 100 MG EXTENDED RELEASE ORAL TABLET|BUPROPION HYDROCHLORIDE 100 MG EXTENDED RELEASE ORAL TABLET
C0693279|T121|993506|RXNORM|BUPROPION HYDROCHLORIDE 100MG M/R TABLET |BUPROPION HYDROCHLORIDE 100 MG EXTENDED RELEASE ORAL TABLET
C0693279|T121|993506|RXNORM|BUPROPION HYDROCHLORIDE 100MG M/R TABLET|BUPROPION HYDROCHLORIDE 100 MG EXTENDED RELEASE ORAL TABLET
C0162758|T121||RXNORM|SEROTONIN UPTAKE INHIBITORS
C0162758|T121||RXNORM|5 HT UPTAKE INHIBITORS
C0162758|T121||RXNORM|5 HYDROXYTRYPTAMINE UPTAKE INHIBITORS
C0162758|T121||RXNORM|INHIBITORS, 5 HT UPTAKE
C0162758|T121||RXNORM|INHIBITORS, 5 HYDROXYTRYPTAMINE UPTAKE
C0162758|T121||RXNORM|UPTAKE INHIBITORS, 5 HT
C0162758|T121||RXNORM|UPTAKE INHIBITORS, 5 HYDROXYTRYPTAMINE
C0162758|T121||RXNORM|SEROTONIN INHIBITOR
C0162758|T121||RXNORM|HT 05 UPTAKE INHIBITORS
C0162758|T121||RXNORM|SEROTONIN UPTAKE INHIB
C0162758|T121||RXNORM|5 HT UPTAKE INHIB
C0162758|T121||RXNORM|SEROTONIN REUPTAKE INHIB
C0162758|T121||RXNORM|INHIB 5 HYDROXYTRYPTAMINE UPTAKE
C0162758|T121||RXNORM|HYDROXYTRYPTAMINE UPTAKE INHIBITORS 05
C0162758|T121||RXNORM|UPTAKE INHIB SEROTONIN
C0162758|T121||RXNORM|INHIB 5 HT UPTAKE
C0162758|T121||RXNORM|UPTAKE INHIB 5 HT
C0162758|T121||RXNORM|5 HYDROXYTRYPTAMINE UPTAKE INHIB
C0162758|T121||RXNORM|REUPTAKE INHIB SEROTONIN
C0162758|T121||RXNORM|INHIB SREOTONIN REUPTAKE
C0162758|T121||RXNORM|UPTAKE INHIB 5 HYDROXYTRYPTAMINE
C0162758|T121||RXNORM|INHIB SEROTONIN UPTAKE
C0162758|T121||RXNORM|SEROTONIN REUPTAKE INHIBITOR
C0162758|T121||RXNORM|SEROTONIN UPTAKE INHIBITOR 
C0162758|T121||RXNORM|SEROTONIN UPTAKE INHIBITOR
C0162758|T121||RXNORM|SEROTONIN UPTAKE INHIBITOR 
C0162758|T121||RXNORM|UPTAKE INHIBITORS, 5-HT
C0162758|T121||RXNORM|SEROTONIN REUPTAKE INHIBITORS
C0162758|T121||RXNORM|UPTAKE INHIBITORS, 5-HYDROXYTRYPTAMINE
C0162758|T121||RXNORM|UPTAKE INHIBITORS, SEROTONIN
C0162758|T121||RXNORM|INHIBITORS, 5-HYDROXYTRYPTAMINE UPTAKE
C0162758|T121||RXNORM|INHIBITORS, 5-HT UPTAKE
C0162758|T121||RXNORM|5-HYDROXYTRYPTAMINE UPTAKE INHIBITORS
C0162758|T121||RXNORM|INHIBITORS, SEROTONIN REUPTAKE
C0162758|T121||RXNORM|REUPTAKE INHIBITORS, SEROTONIN
C0162758|T121||RXNORM|5-HT UPTAKE INHIBITORS
C0162758|T121||RXNORM|INHIBITORS, SEROTONIN UPTAKE
C0162758|T121||RXNORM|SEROTONIN UPTAKE INHIBITOR, NOS
C0486980|T121||RXNORM|HYDROXYBUPROPION
C0486980|T121||RXNORM|4-HYDROXY BUPROPION
C0486980|T121||RXNORM|HYDROXYBUPROPION 
C0068485|T121|31565|RXNORM|NEFAZODONE|NEFAZODONE
C0068485|T121|31565|RXNORM|NEFAZODONE [CHEMICAL/INGREDIENT]|NEFAZODONE
C0068485|T121|31565|RXNORM|NEFAZODONE |NEFAZODONE
C0068485|T121|31565|RXNORM|NEFAZODONE |NEFAZODONE
C0358139|T121|106343|RXNORM|LITHIUM SUCCINATE 0.08 MG/MG TOPICAL OINTMENT|LITHIUM SUCCINATE 8 % TOPICAL OINTMENT
C0358139|T121|106343|RXNORM|LITHIUM SUCCINATE 8 % TOPICAL OINTMENT|LITHIUM SUCCINATE 8 % TOPICAL OINTMENT
C0358139|T121|106343|RXNORM|LITHIUM SUCCINATE 8% OINTMENT|LITHIUM SUCCINATE 8 % TOPICAL OINTMENT
C0358139|T121|106343|RXNORM|LITHIUM SUCCINATE 8% OINTMENT |LITHIUM SUCCINATE 8 % TOPICAL OINTMENT
C0358139|T121|106343|RXNORM|LITHIUM SUCCINATE 8% OINTMENT |LITHIUM SUCCINATE 8 % TOPICAL OINTMENT
C0245561|T121|72625|RXNORM|DULOXETINE|DULOXETINE
C0245561|T121|72625|RXNORM|SELECTIVE NOREPINEPHRINE REUPTAKE INHIBITORS DULOXETINE|DULOXETINE
C0245561|T121|72625|RXNORM|DULOXETINE |DULOXETINE
C0245561|T121|72625|RXNORM|N-METHYL-3-(1-NAPHTHALENYLOXY)-3-(2-THIOPHENE)PROPANAMIDE|DULOXETINE
C0245561|T121|72625|RXNORM|N-METHYL-3-(1-NAPHTHALENYLOXY)-2-THIOPHENEPROPANAMINE|DULOXETINE
C0245561|T121|72625|RXNORM|DULOXETINE |DULOXETINE
C0245561|T121|72625|RXNORM|DULOXETINE |DULOXETINE
C0304364|T121||RXNORM|BICYCLIC ANTIDEPRESSANT 
C0304364|T121||RXNORM|BICYCLIC ANTIDEPRESSANT
C0304364|T121||RXNORM|BICYCLIC ANTIDEPRESSANT, NOS
C0700535|T121|203179|RXNORM|DOXEPIN HYDROCHLORIDE|DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|HYDROCHLORIDE, DOXEPIN|DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|DOXEPIN HYDROCHLORIDE [CHEMICAL/INGREDIENT]|DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|DOXEPIN HYDROCHLORIDE, CIS-TRANS ISOMER MIXTURE (APPROXIMATELY 1:5)|DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|DOXEPIN HYDROCHLORIDE [ANTIPRURITIC] |DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|DOXEPIN HYDROCHLORIDE |DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|DOXEPIN HYDROCHLORIDE [ANTIPRURITIC]|DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|ANTIDEPRESSANTS DOXEPIN HYDROCHLORIDE|DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|ANTIPRURITICS DOXEPIN HYDROCHLORIDE|DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|ANTIPRURITICS DOXEPIN HYDROCHLORIDE |DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|ANTIDEPRESSANTS DOXEPIN HYDROCHLORIDE |DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|DOXEPIN HYDROCHLORIDE |DOXEPIN HYDROCHLORIDE
C0700535|T121|203179|RXNORM|DOXEPIN HYDROCHLORIDE [ANTIPRURITIC] |DOXEPIN HYDROCHLORIDE
C1289960|T121||RXNORM|O-DESMETHYVENLAFAXINE 
C1289960|T121||RXNORM|O-DESMETHYVENLAFAXINE
C3650301|T121||RXNORM|ANTIDEPRESSANTS MAPROTILINE 
C3650301|T121||RXNORM|ANTIDEPRESSANTS MAPROTILINE
C3650306|T121||RXNORM|ANTIDEPRESSANTS ESCITALOPRAM
C3650306|T121||RXNORM|ANTIDEPRESSANTS ESCITALOPRAM 
C2936679|T121||RXNORM|FLUPENTIXOL, MELITRACEN DRUG COMBINATION
C2936679|T121||RXNORM|FLUPENTIXOL - MELITRACEN
C2936679|T121||RXNORM|FLUPENTIXOL + MELITRACEN 
C2936679|T121||RXNORM|FLUPENTIXOL + MELITRACEN
C2936679|T121||RXNORM|ANTIDEPRESSANTS FLUPENTIXOL + MELITRACEN
C3650307|T121||RXNORM|ANTIDEPRESSANTS DOTHIEPIN
C3650307|T121||RXNORM|ANTIDEPRESSANTS DOTHIEPIN 
C0971637|T121||RXNORM|AGOMELATINE
C0971637|T121||RXNORM|AGOMELATINE 
C0971637|T121||RXNORM|AGOMELATINE 
C1993532|T121||RXNORM|NOMIFENSINE &#X7C; BLD-SER-PLAS
C1099456|T121|321988|RXNORM|ESCITALOPRAM|ESCITALOPRAM
C1099456|T121|321988|RXNORM|S(+)-CITALOPRAM|ESCITALOPRAM
C1099456|T121|321988|RXNORM|(S)-CITALOPRAM|ESCITALOPRAM
C1099456|T121|321988|RXNORM|ESCITALOPRAM |ESCITALOPRAM
C1099456|T121|321988|RXNORM|ESCITALOPRAM |ESCITALOPRAM
C0074493|T121|36514|RXNORM|SIBUTRAMINE|SIBUTRAMINE
C0074493|T121|36514|RXNORM|SIBUTRAMINE [CHEMICAL/INGREDIENT]|SIBUTRAMINE
C0074493|T121|36514|RXNORM|SIBUTRAMINE PRODUCT |SIBUTRAMINE
C0074493|T121|36514|RXNORM|SIBUTRAMINE PRODUCT|SIBUTRAMINE
C0074493|T121|36514|RXNORM|SIBUTRAMINE |SIBUTRAMINE
C0074493|T121|36514|RXNORM|SIBUTRAMINE |SIBUTRAMINE
C1981553|T121||RXNORM|ANTIDEPRESSANTS &#X7C; GASTRIC FLUID
C1972481|T121||RXNORM|REBOXETINE &#X7C; BLD-SER-PLAS
C1981554|T121||RXNORM|ANTIDEPRESSANTS &#X7C; URINE
C1975864|T121||RXNORM|ZIMELIDINE &#X7C; BLD-SER-PLAS
C1992738|T121||RXNORM|MOCLOBEMIDE &#X7C; BLD-SER-PLAS
C1994490|T121||RXNORM|PHENELZINE &#X7C; BLD-SER-PLAS
C1981552|T121||RXNORM|ANTIDEPRESSANTS &#X7C; BLD-SER-PLAS
C0072127|T121|34604|RXNORM|1-(ALPHA-PROPYLPHENETHYL)PYRROLIDINE|PROLINTANE
C0072127|T121|34604|RXNORM|PHENYLPYRROLIDINYLPENTAN|PROLINTANE
C0072127|T121|34604|RXNORM|PROLINTANE|PROLINTANE
C0072127|T121|34604|RXNORM|PROLINTANE |PROLINTANE
C0072127|T121|34604|RXNORM|PROLINTANE |PROLINTANE
C0076652|T121|38252|RXNORM|(3-CHLORO-6-METHYL-5,5-DIOXO-6,11-DIHYDRODIBENZO(C,F)(1,2)THIAZEPIN-11-YL)-7-AMINOHEPTANOIC ACID|TIANEPTINE
C0076652|T121|38252|RXNORM|TIANEPTINE|TIANEPTINE
C0076652|T121|38252|RXNORM|TIANEPTINE |TIANEPTINE
C3847513|T121||RXNORM|VILAZODONE &#X7C; URINE
C0040098|T121||RXNORM|THYMOLEPTICS
C0040094|T121||RXNORM|THYMOANALEPTICS
C0771509|T121||RXNORM|TIANEPTINE SODIUM
C0771509|T121||RXNORM|TIANEPTINE SODIUM 
C0771509|T121||RXNORM|TIANEPTINE SODIUM 
C4038278|T121||RXNORM|CITALOPRAM+ESCITALOPRAM &#X7C; URINE
C3661282|T121|1455099|RXNORM|VORTIOXETINE|VORTIOXETINE
C3661282|T121|1455099|RXNORM|1-(2-(2,4-DIMETHYLPHENYLSULFANYL)PHENYL)PIPERAZINE|VORTIOXETINE
C3661282|T121|1455099|RXNORM|ANTIDEPRESSANTS VORTIOXETINE|VORTIOXETINE
C3661282|T121|1455099|RXNORM|VORTIOXETINE |VORTIOXETINE
C3661282|T121|1455099|RXNORM|VORTIOXETINE |VORTIOXETINE
C1742884|T121|683693|RXNORM|DESVENLAFAXINE SUCCINATE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|DESVENLAFAXINE SUCCINATE |DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|DESVENLAFAXINE SUCCINATE |DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|BUTANEDIOIC ACID, COMPOUND WITH 4-(2-(DIMETHYLAMINO)-1-(1-HYDROXYCYCLOHEXYL)ETHYL)PHENOL (1:1), MONOHYDRATE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|SUCCINATE MONOHYDRATE, O-DESMETHYLVENLAFAXINE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|MONOHYDRATE, O-DESMETHYLVENLAFAXINE SUCCINATE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|O DESMETHYLVENLAFAXINE SUCCINATE MONOHYDRATE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|SUCCINATE, DESVENLAFAXINE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|O DESMETHYLVENLAFAXINE SUCCINATE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|SUCCINATE, O-DESMETHYLVENLAFAXINE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|O-DESMETHYLVENLAFAXINE SUCCINATE MONOHYDRATE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|O-DESMETHYLVENLAFAXINE SUCCINATE|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|DESVENLAFAXINE SUCCINATE [CHEMICAL/INGREDIENT]|DESVENLAFAXINE SUCCINATE
C1742884|T121|683693|RXNORM|2-(1-HYDROXYCYCLOHEXYL)-2-((4-HYDROXYPHENYL)ETHYL)DIMETHYLAMMONIUM 3-CARBOXYPROPANOATE MONOHYDRATE|DESVENLAFAXINE SUCCINATE
C1505020|T121|476250|RXNORM|DULOXETINE HYDROCHLORIDE|DULOXETINE HYDROCHLORIDE
C1505020|T121|476250|RXNORM|DULOXETINE HYDROCHLORIDE |DULOXETINE HYDROCHLORIDE
C1505020|T121|476250|RXNORM|DULOXETINE HYDROCHLORIDE |DULOXETINE HYDROCHLORIDE
C1505020|T121|476250|RXNORM|HYDROCHLORIDE, DULOXETINE|DULOXETINE HYDROCHLORIDE
C1505020|T121|476250|RXNORM|HCL, DULOXETINE|DULOXETINE HYDROCHLORIDE
C1505020|T121|476250|RXNORM|DULOXETINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|DULOXETINE HYDROCHLORIDE
C1505020|T121|476250|RXNORM|DULOXETINE HCL|DULOXETINE HYDROCHLORIDE
C2980164|T121||RXNORM|GABOXETINE KIT
C2980164|T121||RXNORM|GABOXETINE CONVENIENCE PACK
C2980164|T121||RXNORM|ACETYLCARNITINE/CHOLINE BITARTRATE/COCOA EXTRACT/GAMMA AMINOBUTYRIC ACID/GINKGO BILOBA LEAF/GLUTAMIC ACID/GRAPE SEED EXTRACT/GRIFFONIA SEED EXTRACT/VALERIAN ROOT EXTRACT/WHEY PROTEIN HYDROLYSATE;FLUOXETINE HYDROCHLORIDE 62.5 MG; 10 MG ORAL CAPSULE [GABOXETINE]
C0041249|T121|10898|RXNORM|L TRYPTOPHAN|TRYPTOPHAN
C0041249|T121|10898|RXNORM|TRYPTOPHAN|TRYPTOPHAN
C0041249|T121|10898|RXNORM|L-TRYPTOPHAN|TRYPTOPHAN
C0041249|T121|10898|RXNORM|L-TRYPTOPHAN |TRYPTOPHAN
C0041249|T121|10898|RXNORM|LEVOTRYPTOPHAN|TRYPTOPHAN
C0041249|T121|10898|RXNORM|TRYPTOPHAN [CHEMICAL/INGREDIENT]|TRYPTOPHAN
C0041249|T121|10898|RXNORM|L-TRYPTOPHAN |TRYPTOPHAN
C0041249|T121|10898|RXNORM|TRP|TRYPTOPHAN
C0041249|T121|10898|RXNORM|(S)-2-AMINO-3-(1H-INDOL-3-YL)-PROPANOIC ACID|TRYPTOPHAN
C0041249|T121|10898|RXNORM|TRYPTOPHAN PRODUCT|TRYPTOPHAN
C0041249|T121|10898|RXNORM|L-TRYPTOPHAN |TRYPTOPHAN
C0041249|T121|10898|RXNORM|TRYPTOPHAN |TRYPTOPHAN
C0023870|T121|6448|RXNORM|LITHIUM|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM PRODUCT|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM |LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM [CHEMICAL/INGREDIENT]|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM METALLICUM|LITHIUM
C0023870|T121|6448|RXNORM|LI|LITHIUM
C0023870|T121|6448|RXNORM|LI ELEMENT|LITHIUM
C0023870|T121|6448|RXNORM|LI+ ELEMENT|LITHIUM
C0023870|T121|6448|RXNORM|LI - LITHIUM|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM |LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM |LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM, NOS|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM PRODUCT |LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM PRODUCT |LITHIUM
C0042665|T121|11196|RXNORM|VILOXAZINE|VILOXAZINE
C0042665|T121|11196|RXNORM|MORPHOLINE, 2-((2-ETHOXYPHENOXY)METHYL)-|VILOXAZINE
C0042665|T121|11196|RXNORM|VILOXAZINE [CHEMICAL/INGREDIENT]|VILOXAZINE
C0042665|T121|11196|RXNORM|VILOXAZINE |VILOXAZINE
C0042665|T121|11196|RXNORM|VILOXAZINE |VILOXAZINE
C0168388|T121|60842|RXNORM|REBOXETINE|REBOXETINE
C0168388|T121|60842|RXNORM|REBOXETINE [CHEMICAL/INGREDIENT]|REBOXETINE
C0168388|T121|60842|RXNORM|SELECTIVE NOREPINEPHRINE REUPTAKE INHIBITORS REBOXETINE|REBOXETINE
C0168388|T121|60842|RXNORM|REBOXETINE |REBOXETINE
C0168388|T121|60842|RXNORM|REBOXETINE |REBOXETINE
C0168388|T121|60842|RXNORM|REBOXETINE |REBOXETINE
C0360108|T121||RXNORM|TETRACYCLIC ANTIDEPRESSANT
C0360108|T121||RXNORM|TETRACYCLIC ANTIDEPRESSANT DRUG
C0360108|T121||RXNORM|TETRACYCLIC ANTIDEPRESSANT 
C0360108|T121||RXNORM|TETRACYCLIC ANTIDEPRESSANT 
C0360108|T121||RXNORM|TETRACYCLIC ANTIDEPRESSANT, NOS
C1271027|T121||RXNORM|TRIAZOLOPYRIDINE
C1271027|T121||RXNORM|TRIAZOLOPYRIDINE 
C1271027|T121||RXNORM|TRIAZOLOPYRIDINE 
C0012035|T121||RXNORM|DIBENZOTHIEPINS
C0012035|T121||RXNORM|DIBENZOTHIEPINS [CHEMICAL/INGREDIENT]
C0012035|T121||RXNORM|DIBENZOTHIEPIN
C0012035|T121||RXNORM|DIBENZOTHIEPIN 
C0063220|T121|1546455|RXNORM|1,3,4,6,8,13-HEXAHYDROXY-10,11-DIMETHYLPHENANTHRO(1,10,9,8-OPQRA)PERYLENE-7,14-DIONE|HYPERICIN
C0063220|T121|1546455|RXNORM|HYPERICIN|HYPERICIN
C0063220|T121|1546455|RXNORM|4,5,7,4',5',7'-HEXAHYDROXY-2,2'-DIMETHYL-MESONAPTHTODIANTHRON|HYPERICIN
C0063220|T121|1546455|RXNORM|HYPERICIN |HYPERICIN
C0066561|T121|30031|RXNORM|3-(MORPHOLINOETHYL)AMINO-4-METHYL-6-PHENYLPYRIDAZINE|MINAPRINE
C0066561|T121|30031|RXNORM|MINAPRINE|MINAPRINE
C0066561|T121|30031|RXNORM|N-(4-METHYL-6-PHENYL-3-PYRIDAZINYL)-4-MORPHOLINEETHANAMINE|MINAPRINE
C0066561|T121|30031|RXNORM|4-MORPHOLINEETHANAMINE, N-(4-METHYL-6-PHENYL-3-PYRIDAZINYL)-|MINAPRINE
C0074500|T121||RXNORM|MESOCARB
C0074500|T121||RXNORM|N-PHENYLCARBAMOYL-3-(BETA-PHENYLISOPROPYL)SYDNONIMINE
C0074500|T121||RXNORM|SIDNOCARB
C0074500|T121||RXNORM|SYDNOCARB
C0071143|T121||RXNORM|1,10-TRIMETHYLENE-8-METHYL-1,2,3,4-TETRAHYDROPYRAZINO(1,2-A)INDOLE
C0071143|T121||RXNORM|1H-PYRAZINO(3,2,1-JK)CARBAZOLE, 2,3,3A,4,5,6-HEXAHYDRO-8-METHYL-, MONOHYDROCHLORIDE
C0071143|T121||RXNORM|PIRLINDOL
C0071143|T121||RXNORM|PIRLINDOLE
C0071143|T121||RXNORM|PYRLINDOLE
C0060145|T121||RXNORM|FEMOXETINE
C0060145|T121||RXNORM|FEMOXITINE
C0060145|T121||RXNORM|PIPERIDINE, 3-((4-METHOXYPHENOXY)METHYL)-1-METHYL-4-PHENYL-, (3R-TRANS)-
C0060145|T121||RXNORM|TRANS-(+)-3-((4-METHOXYPHENOXY)METHYL)-1-METHYL-4-PHENYLPIPERIDINE
C0060145|T121||RXNORM|TRANS-3-((4-METHOXYPHENOXY)METHYL)-1-METHYL-4-PHENYLPIPERIDINE
C0076804|T121|38382|RXNORM|(3-METHYL)-3-PHENYL-5-HYDROXYMETHYL-2-OXAZOLIDINONE|TOLOXATONE
C0076804|T121|38382|RXNORM|5-(HYDROXYMETHYL)-3-(3-METHYLPHENYL)-2- OXAZOLIDINONE|TOLOXATONE
C0076804|T121|38382|RXNORM|TOLOXATONE|TOLOXATONE
C0076804|T121|38382|RXNORM|5-(HYDROXYMETHYL)-3-(3-METHYLPHENYL)-2-OXAZOLIDINONE|TOLOXATONE
C0076804|T121|38382|RXNORM|5-HYDROXYMETHYL-3-(M-TOLYL)-2-OXAZOLIDINONE|TOLOXATONE
C0076784|T121|38365|RXNORM|1-(3,4-DIMETHOXYPHENYL)-5-ETHYL-7,8-DIMETHOXY- 4-METHYL-5H-2,3-BENZODIAZEPINE|TOFISOPAM
C0076784|T121|38365|RXNORM|TOFISOPAM|TOFISOPAM
C0076784|T121|38365|RXNORM|TOFIZOPAM|TOFISOPAM
C0076784|T121|38365|RXNORM|1-(3,4-DIMETHOXYPHENYL)-5-ETHYL-7,8-DIMETHOXY-4-METHYL-5H-2,3-BENZODIAZEPINE|TOFISOPAM
C0069039|T121||RXNORM|3-(4-BROMOPHENYL)-N-METHYL-(3-PYIIDYL)ALLYLAMINE OXALATE
C0069039|T121||RXNORM|NORZIMELDINE
C0069039|T121||RXNORM|NORZIMELIDINE
C0072076|T121|34568|RXNORM|BUTANAMIDE, 4-(((4-CHLOROPHENYL)(5-FLUORO-2-HYDROXYPHENYL)METHYLENE)AMINO)-|PROGABIDE
C0072076|T121|34568|RXNORM|PROGABIDE|PROGABIDE
C0063448|T121||RXNORM|(3-INDOLYL-2-ETHYL)PIPERIDINE
C0063448|T121||RXNORM|1H-INDOLE, 3-(2-(4-PIPERIDINYL)ETHYL)-
C0063448|T121||RXNORM|4-(2-(3-INDOLYL)ETHYL)PIPERIDINE
C0063448|T121||RXNORM|INDALPINE
C0043636|T121||RXNORM|(DES-TYR(1))-GAMMA-ENDORPHIN
C0043636|T121||RXNORM|1-DE-TYR-GAMMA-ENDORPHIN
C0043636|T121||RXNORM|BETA-LIPOTROPIN(62-77)
C0043636|T121||RXNORM|BETA-LPH(62-77)
C0043636|T121||RXNORM|DTGAMMAE
C0043636|T121||RXNORM|GAMMA-ENDORPHIN, DES-TYR(1)-
C0043636|T121||RXNORM|GAMMA-ENDORPHIN, DES-TYROSINE(1)-
C0139500|T121||RXNORM|PYRO(L-ALPHA-AMINOADIPYL)-L-HISTIDYL-L-THIAZOLIDINE-4-CARBOXAMIDE
C0139500|T121||RXNORM|PYRO-AAD-HIS-TZL-NH2
C0139500|T121||RXNORM|PYRO-2-AMINOADIPYLHISTIDYLTHIAZOLIDINE-4-CARBOXYAMIDE
C0139500|T121||RXNORM|(2S)-N-((2S)-1-((4S)-4-CARBAMOYL-1,3-THIAZOLIDIN-3-YL)-3-(1H-IMIDAZOL-5-YL)-1-OXO-2-PROPANYL)-6-OXO-2-PIPERIDINECARBOXAMIDE
C0075784|T121||RXNORM|2-AMINO-6-ALLYL-5,6,7,8-TETRAHYDRO-4H-THIAZOLO-(5,4-D)AZEPIN-DIHYDROCHLORIDE
C0075784|T121||RXNORM|4H-THIAZOLO(4,5-D)AZEPIN-2-AMINE, 5,6,7,8-TETRAHYDRO-6-(2-PROPENYL)-, DIHYDROCHLORIDE
C0075784|T121||RXNORM|TALIPEXOLE
C0075784|T121||RXNORM|6-ALLYL-2-AMINO-5,6,7,8-TETRAHYDRO-4H-THIAZOLO(4,5-D)AZEPIN DIHYDROCHLORIDE
C0051086|T121||RXNORM|ALAPROCLATE
C0051086|T121||RXNORM|DL-ALANINE, 2-(4-CHLOROPHENYL)-1,1-DIMETHYLETHYL ESTER
C0063159|T121||RXNORM|HYDROXYMAPROTILIN
C0063159|T121||RXNORM|OXAPROTILINE
C0106291|T121|47111|RXNORM|1-BUTANAMINE, N-METHYL-4-(2-(PHENYLMETHYL)PHENOXY)-, HYDROCHLORIDE|BIFEMELANE
C0106291|T121|47111|RXNORM|2-(4-METHYLAMINOBUTOXY)DIPHENYLMETHANE|BIFEMELANE
C0106291|T121|47111|RXNORM|4-(2-BENZYLPHENOXY)-N-METHYLBUTYLAMINE|BIFEMELANE
C0106291|T121|47111|RXNORM|BIFEMELANE|BIFEMELANE
C0051917|T121|17939|RXNORM|1-(4-METHOXYBENZOYL)-2-PYRROLIDINONE|ANIRACETAM
C0051917|T121|17939|RXNORM|1-ANISOYL-2-PYRROLIDINONE|ANIRACETAM
C0051917|T121|17939|RXNORM|ANIRACETAM|ANIRACETAM
C0050844|T121||RXNORM|ADINAZOLAM
C0066624|T121||RXNORM|4,4-DIMETHYL-1-(4-(4-(2-PYRIMIDINYL)-1-PIPERAZINYL)BUTYL)-2,6-PIPERIDINEDIONE
C0066624|T121||RXNORM|GEPIRONE
C0075591|T121||RXNORM|SULFORIDAZINE
C0060454|T121||RXNORM|FLESINOXAN
C0060454|T121||RXNORM|P-FLUORO-N-(2-(4-(2-(HYDROXYMETHYL)-1,4-BENZODIOXAN-5-YL)-1-PIPERAZINYL)ETHYL)BENZAMIDE
C0299772|T121||RXNORM|L 701,324
C0299772|T121||RXNORM|L 701324
C0299772|T121||RXNORM|L-701,324
C0299772|T121||RXNORM|L-701324
C1445647|T121||RXNORM|PHENYLPIPERAZINE ANTIDEPRESSANT 
C1445647|T121||RXNORM|PHENYLPIPERAZINE ANTIDEPRESSANT
C0303506|T121||RXNORM|LITHIUM AND ITS DERIVATIVES
C0303506|T121||RXNORM|LITHIUM AND/OR LITHIUM COMPOUND 
C0303506|T121||RXNORM|LITHIUM AND/OR LITHIUM COMPOUND
C1881039|T121||RXNORM|HEPZIDINE
C1880846|T121||RXNORM|FOSENAZIDE
C0123216|T121||RXNORM|IFOXETINE
C0600526|T121|155137|RXNORM|SERTRALINE HYDROCHLORIDE|SERTRALINE HYDROCHLORIDE
C0600526|T121|155137|RXNORM|HYDROCHLORIDE, SERTRALINE|SERTRALINE HYDROCHLORIDE
C0600526|T121|155137|RXNORM|SERTRALINE HYDROCHLORIDE |SERTRALINE HYDROCHLORIDE
C0600526|T121|155137|RXNORM|ANTIDEPRESSANTS SERTRALINE HYDROCHLORIDE|SERTRALINE HYDROCHLORIDE
C0600526|T121|155137|RXNORM|SERTRALINE HYDROCHLORIDE (1S-CIS)-ISOMER|SERTRALINE HYDROCHLORIDE
C0600526|T121|155137|RXNORM|SERTRALINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|SERTRALINE HYDROCHLORIDE
C0600526|T121|155137|RXNORM|SERTRALINE HYDROCHLORIDE |SERTRALINE HYDROCHLORIDE
C0600526|T121|155137|RXNORM|SERTRALINE HYDROCHLORIDE |SERTRALINE HYDROCHLORIDE
C1881247|T121||RXNORM|INTRIPTYLINE
C1831797|T121||RXNORM|CASOPITANT MESYLATE
C0060394|T121||RXNORM|FIPEXIDE
C0733380|T121|227224|RXNORM|FLUOXETINE HYDROCHLORIDE|FLUOXETINE HYDROCHLORIDE
C0733380|T121|227224|RXNORM|ANTIDEPRESSANTS FLUOXETINE HYDROCHLORIDE|FLUOXETINE HYDROCHLORIDE
C0733380|T121|227224|RXNORM|FLUOXETINE HYDROCHLORIDE |FLUOXETINE HYDROCHLORIDE
C0733380|T121|227224|RXNORM|FLUOXETINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|FLUOXETINE HYDROCHLORIDE
C0733380|T121|227224|RXNORM|FLUOXETINE HCL|FLUOXETINE HYDROCHLORIDE
C0733380|T121|227224|RXNORM|FLUOXETINE HYDROCHLORIDE |FLUOXETINE HYDROCHLORIDE
C0733380|T121|227224|RXNORM|FLUOXETINE HYDROCHLORIDE [DUP] |FLUOXETINE HYDROCHLORIDE
C1880764|T121||RXNORM|FEPROSIDNINE
C1881816|T121||RXNORM|MEZEPINE
C0526501|T121|135091|RXNORM|4-AMINO-5-CHLORO-2-ETHOXY-N-((4-(4-FLUOROBENZYL)-2-MORPHOLINYL)METHYL)BENZAMIDE|MOSAPRIDE
C0526501|T121|135091|RXNORM|BENZAMIDE, 4-AMINO-5-CHLORO-2-ETHOXY-N-((4-((4-FLUOROPHENYL)METHYL)-2-MORPHOLINYL)METHYL)-, 2-HYDROXY-1,2,3-PROPANETRICARBOXYLATE (1:1)|MOSAPRIDE
C0526501|T121|135091|RXNORM|MOSAPRIDE|MOSAPRIDE
C1881248|T121||RXNORM|INTRIPTYLINE HYDROCHLORIDE
C1873234|T121||RXNORM|TESOFENSINE
C1881896|T121||RXNORM|MONOMETACRINE
C1880560|T121||RXNORM|ETACEPRIDE
C1881131|T121||RXNORM|IMAFEN HYDROCHLORIDE
C1880288|T121|734064|RXNORM|DESVENLAFAXINE|DESVENLAFAXINE
C1880288|T121|734064|RXNORM|DESVENLAFAXINE |DESVENLAFAXINE
C1880288|T121|734064|RXNORM|DESVENLAFAXINE |DESVENLAFAXINE
C1880288|T121|734064|RXNORM|O DESMETHYLVENLAFAXINE|DESVENLAFAXINE
C1880288|T121|734064|RXNORM|4-(2-(DIMETHYLAMINO)-1-(1-HYDROXYCYCLOHEXYL)ETHYL)PHENOL|DESVENLAFAXINE
C1880288|T121|734064|RXNORM|O-DESMETHYLVENLAFAXINE|DESVENLAFAXINE
C1880733|T121||RXNORM|FANTRIDONE HYDROCHLORIDE
C0065963|T121||RXNORM|MEPIPRAZOLE
C0070047|T121||RXNORM|1-BENZOYL-3-(1-(2-NAPHTHYLMETHYL)-4-PIPERIDYL)UREA
C0070047|T121||RXNORM|PANURAMINE
C1881414|T121||RXNORM|LITRACEN
C1880857|T121||RXNORM|FTORPROPAZINE
C0165077|T121||RXNORM|4-(2-NAPHTHALENYLMETHOXY)PIPERIDINE
C0165077|T121||RXNORM|LITOXETINE
C1881811|T121||RXNORM|METOXEPIN
C0066473|T121||RXNORM|1H-3,4,6A-TRIAZAFLUORANTHENE, 2,4,5,6-TETRAHYDRO-9-METHOXY-4-METHYL-
C0066473|T121||RXNORM|3-METHYL-8-METHOXY-(3H)-1,2,5,6-TETRAHYDROPYRAZINO(1,2,3-AB)-BETA-CARBOLINE
C0066473|T121||RXNORM|METRALINDOLE
C0117861|T121||RXNORM|FLEROBUTEROL
C1365510|T121|436212|RXNORM|PAROXETINE MESYLATE|PAROXETINE MESYLATE
C1365510|T121|436212|RXNORM|PAROXETINE METHANESULFONATE|PAROXETINE MESYLATE
C1365510|T121|436212|RXNORM|PIPERIDINE, 3-((1,3-BENZODIOXOL-5-YLOXY)METHYL)-4-(4-FLUOROPHENYL)-,(3S,4R)-, METHANESULFONATE|PAROXETINE MESYLATE
C1365510|T121|436212|RXNORM|PAROXETINE MESYLATE |PAROXETINE MESYLATE
C1365510|T121|436212|RXNORM|PAROXETINE MESYLATE |PAROXETINE MESYLATE
C1365510|T121|436212|RXNORM|(-)-(3S,4R)-4-(P-FLUOROPHENYL)-3-((3,4-(METHYLENEDIOXY)PHENOXY)METHYL)PIPERIDINE MESYLATE|PAROXETINE MESYLATE
C1365510|T121|436212|RXNORM|PAROXETINE MESILATE|PAROXETINE MESYLATE
C1882438|T121||RXNORM|PRAZEPINE
C1881288|T121||RXNORM|IVOQUALINE
C0078842|T121||RXNORM|4-(3-CHLOROPHENYL)-1,6,7,8-TETRAHYDRO-1,3-DIMETHYLPYRAZOLO(3,4-E)(1,4)DIAZEPINE
C0078842|T121||RXNORM|ZOMETAPINE
C0700563|T121|203204|RXNORM|BUPROPION HYDROCHLORIDE|BUPROPION HYDROCHLORIDE
C0700563|T121|203204|RXNORM|(+-)-1-(3-CHLOROPHENYL)-2-[(1,1-DIMETHYLETHYL)AMINO]-1-PROPANONE HYDROCHLORIDE|BUPROPION HYDROCHLORIDE
C0700563|T121|203204|RXNORM|ANTIDEPRESSANTS BUPROPION HYDROCHLORIDE|BUPROPION HYDROCHLORIDE
C0700563|T121|203204|RXNORM|BUPROPION HYDROCHLORIDE |BUPROPION HYDROCHLORIDE
C0700563|T121|203204|RXNORM|BUPROPION HYDROCHLORIDE [CHEMICAL/INGREDIENT]|BUPROPION HYDROCHLORIDE
C0700563|T121|203204|RXNORM|BUPROPION HYDROCHLORIDE |BUPROPION HYDROCHLORIDE
C0700563|T121|203204|RXNORM|BUPROPION HYDROCHLORIDE |BUPROPION HYDROCHLORIDE
C1170741|T121|353103|RXNORM|ATOMOXETINE HYDROCHLORIDE|ATOMOXETINE HYDROCHLORIDE
C1170741|T121|353103|RXNORM|(-)-N -METHYL-3-PHENYL-3-(O-TOLYLOXY)-PROPYLAMINE HYDROCHLORIDE|ATOMOXETINE HYDROCHLORIDE
C1170741|T121|353103|RXNORM|(-)-N-METHYL-GAMMA(2-METHYLPHENOXY)BENZENEPROPAMINE HYDROCHLORIDE|ATOMOXETINE HYDROCHLORIDE
C1170741|T121|353103|RXNORM|ATOMOXETINE HCL|ATOMOXETINE HYDROCHLORIDE
C1170741|T121|353103|RXNORM|ATOMOXETINE HCL |ATOMOXETINE HYDROCHLORIDE
C1170741|T121|353103|RXNORM|HCL, ATOMOXETINE|ATOMOXETINE HYDROCHLORIDE
C1170741|T121|353103|RXNORM|HYDROCHLORIDE, ATOMOXETINE|ATOMOXETINE HYDROCHLORIDE
C1170741|T121|353103|RXNORM|ATOMOXETINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|ATOMOXETINE HYDROCHLORIDE
C1170741|T121|353103|RXNORM|N-METHYL-GAMMA-(2-METHYLPHENOXY)BENZENEPROPANAMINE HYDROCHLORIDE|ATOMOXETINE HYDROCHLORIDE
C1170741|T121|353103|RXNORM|ATOMOXETINE HYDROCHLORIDE |ATOMOXETINE HYDROCHLORIDE
C0771310|T121|236082|RXNORM|NEFAZODONE HYDROCHLORIDE|NEFAZODONE HYDROCHLORIDE
C0771310|T121|236082|RXNORM|ANTIDEPRESSANTS NEFAZODONE HYDROCHLORIDE|NEFAZODONE HYDROCHLORIDE
C0771310|T121|236082|RXNORM|NEFAZODONE HYDROCHLORIDE |NEFAZODONE HYDROCHLORIDE
C0771310|T121|236082|RXNORM|NEFAZODONE HYDROCHLORIDE |NEFAZODONE HYDROCHLORIDE
C0771310|T121|236082|RXNORM|NEFAZODONE HYDROCHLORIDE |NEFAZODONE HYDROCHLORIDE
C0771310|T121|236082|RXNORM|NEFAZADONE HCL|NEFAZODONE HYDROCHLORIDE
C1881066|T121||RXNORM|HOMOPIPRAMOL
C1881066|T121||RXNORM|2-(4-(3-(5H-DIBENZ(B,F)AZEPIN-5-YL)PROPYL)-1,4-DIAZEPIN-1-YL)ETHANOL
C1881066|T121||RXNORM|4-(3-(5H-DIBENZ(B,F)AZEPIN-5-YL)PROPYL)HEXAHYDRO-1H-1,4-DIAZEPINE-1-ETHANOL
C0071001|T121||RXNORM|EPTASTIGMINE
C0071001|T121||RXNORM|HEPTYL PHYSOSTIGMINE
C0071001|T121||RXNORM|PHYSOSTIGMINE HEPTYL
C0071001|T121||RXNORM|PYRROLO(2,3-B)INDOL-5-OL-1,2,3,3A,8,8A-HEXAHYDRO-1,3A,8-TRIMETHYL HEPTYLCARBAMATE ESTER
C0071001|T121||RXNORM|HEPTASTIGMINE
C0071001|T121||RXNORM|HEPTYLPHYSOSTIGMINE
C0071001|T121||RXNORM|HEPTYL-PHYSOSTIGMINE
C0724555|T121|221078|RXNORM|CITALOPRAM (AS CITALOPRAM HYDROBROMIDE)|CITALOPRAM HYDROBROMIDE
C0724555|T121|221078|RXNORM|CITALOPRAM HYDROBROMIDE|CITALOPRAM HYDROBROMIDE
C0724555|T121|221078|RXNORM|(![PLUS-MINUS SIGN]!)-1-(3-DIMETHYLAMINOPROPYL)-1- (4-FLUOROPHENYL)-1,3 DIHYDROISOBENZOFURAN-5-CARBONITRILE, HBR|CITALOPRAM HYDROBROMIDE
C0724555|T121|221078|RXNORM|(±)-1-(3-DIMETHYLAMINOPROPYL)-1- (4-FLUOROPHENYL)-1,3 DIHYDROISOBENZOFURAN-5-CARBONITRILE, HBR|CITALOPRAM HYDROBROMIDE
C0724555|T121|221078|RXNORM|CITALOPRAM HYDROBROMIDE |CITALOPRAM HYDROBROMIDE
C0724555|T121|221078|RXNORM|1-[3-(DIMETHYLAMINO)PROPYL]-1-(4-FLUOROPHENYL)-1,3-DIHYDRO-5-ISOBENZOFURANCARBONITRILE MONOHYDROBROMIDE|CITALOPRAM HYDROBROMIDE
C0724555|T121|221078|RXNORM|CITALOPRAM HYDROBROMIDE |CITALOPRAM HYDROBROMIDE
C1880541|T121||RXNORM|EPROBEMIDE
C1881269|T121||RXNORM|IROLAPRIDE
C0771019|T121|235830|RXNORM|PAROXETINE HYDROCHLORIDE|PAROXETINE HYDROCHLORIDE
C0771019|T121|235830|RXNORM|PAROXETINE HYDROCHLORIDE |PAROXETINE HYDROCHLORIDE
C0771019|T121|235830|RXNORM|(-)-(3S,4R)-4-(P-FLUOROPHENYL)-3-((3,4-(METHYLENEDIOXY)PHENOXY)METHYL)PIPERIDINE HYDROCHLORIDE|PAROXETINE HYDROCHLORIDE
C0771019|T121|235830|RXNORM|PAROXETINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|PAROXETINE HYDROCHLORIDE
C0771019|T121|235830|RXNORM|HYDROCHLORIDE, PAROXETINE|PAROXETINE HYDROCHLORIDE
C0771019|T121|235830|RXNORM|PAROXETINE HYDROCHLORIDE |PAROXETINE HYDROCHLORIDE
C0771019|T121|235830|RXNORM|PAROXETINE HYDROCHLORIDE |PAROXETINE HYDROCHLORIDE
C0282369|T121|82112|RXNORM|TRAZODONE HYDROCHLORIDE|TRAZODONE HYDROCHLORIDE
C0282369|T121|82112|RXNORM|2-(3-(4-(3-CHLOROPHENYL)PIPERAZIN-1-Y)PROPYL)-1,2,4-TRIAZOLO(4,3-A)PYRIDINE-3(2H)-ONE HYDROCHLORIDE|TRAZODONE HYDROCHLORIDE
C0282369|T121|82112|RXNORM|1,2,4-TRIAZOLO(4,3-A)PYRIDIN-3(2H)-ONE, 2-(3-(4-(3-CHLOROPHENYL)-1-PIPERAZINYL)PROPYL)-, MONOHYDROCHLORIDE|TRAZODONE HYDROCHLORIDE
C0282369|T121|82112|RXNORM|TRAZODONE HYDROCHLORIDE |TRAZODONE HYDROCHLORIDE
C0282369|T121|82112|RXNORM|ANTIDEPRESSANTS TRAZODONE HYDROCHLORIDE|TRAZODONE HYDROCHLORIDE
C0282369|T121|82112|RXNORM|TRAZODONE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|TRAZODONE HYDROCHLORIDE
C0282369|T121|82112|RXNORM|TRAZODONE HYDROCHLORIDE |TRAZODONE HYDROCHLORIDE
C0282369|T121|82112|RXNORM|TRAZODONE HYDROCHLORIDE [DUP] |TRAZODONE HYDROCHLORIDE
C0208216|T121||RXNORM|3-CHLORO-5-(3-(2-OXO-1,2,3,5,6,7,8,8A-OCTAHYDROIMIDAZO(1,2-A)PYRIDINE-3-SPIRO-4'-PIPERIDINO)PROPYL)-10,11-DIHYDRO-5H-DIBENZ(B,F)AZEPINE
C0208216|T121||RXNORM|MOSAPRAMINE
C0208216|T121||RXNORM|SPIRO(IMIDAZO(1,2-A)PYRIDINE-3(2H),4'-PIPERIDIN)-2-ONE, 1'-(3-(3-CHLORO-10,11-DIHYDRO-5H-DIBENZ(B,F)AZEPIN-5-YL)PROPYL)HEXAHYDRO-, DIHYDROCHLORIDE
C0700473|T121|203143|RXNORM|FLUVOXAMINE MALEATE|FLUVOXAMINE MALEATE
C0700473|T121|203143|RXNORM|FLUVOXAMINE MALEATE |FLUVOXAMINE MALEATE
C0700473|T121|203143|RXNORM|FLUVOXAMINE MALEATE [CHEMICAL/INGREDIENT]|FLUVOXAMINE MALEATE
C0700473|T121|203143|RXNORM|FLUVOXAMINE MALEATE |FLUVOXAMINE MALEATE
C0700473|T121|203143|RXNORM|FLUVOXAMINE MALEATE, (E)-ISOMER|FLUVOXAMINE MALEATE
C0700473|T121|203143|RXNORM|FLUVOXAMINE MALEATE [DUP] |FLUVOXAMINE MALEATE
C1880815|T121||RXNORM|FLUOXETINE HYDROCHLORIDE, (R)-
C1880815|T121||RXNORM|FLUOXETINE HYDROCHLORIDE, R-
C1880815|T121||RXNORM|BENZENEPROPANAMINE, N-METHYL-GAMMA-(4-(TRIFLUOROMETHYL)PHENOXY)-, HYDROCHLORIDE (1:1), (GAMMA R)-
C0074710|T121|746741|RXNORM|2,6-BENZOTHIAZOLEDIAMINE, 4,5,6,7-TETRAHYDRO-N6-PROPYL-, (S)-|PRAMIPEXOLE
C0074710|T121|746741|RXNORM|2-AMINO-4,5,6,7-TETRAHYDRO-6-PROPYLAMINOBENZOTHIAZOLE|PRAMIPEXOLE
C0074710|T121|746741|RXNORM|PRAMIPEXOLE|PRAMIPEXOLE
C0074710|T121|746741|RXNORM|2-AMINO-6-PROPYLAMINOTETRAHYDROBENZOTHIAZOLE|PRAMIPEXOLE
C0074710|T121|746741|RXNORM|4,5,6,7-TETRAHYDRO-N6-PROPYL-2,6-BENZOTHIAZOLE-DIAMINE|PRAMIPEXOLE
C0074710|T121|746741|RXNORM|PRAMIPEXOL|PRAMIPEXOLE
C0074710|T121|746741|RXNORM|PRAMIPEXOLE |PRAMIPEXOLE
C0074710|T121|746741|RXNORM|PRAMIPEXOLE |PRAMIPEXOLE
C1882243|T121||RXNORM|OXITRIPTYLINE
C0127034|T121||RXNORM|MAROXEPIN
C0127034|T121||RXNORM|MAROXEPINE
C1882439|T121||RXNORM|PRAZITONE
C1880799|T121||RXNORM|FLUBEPRIDE
C0125988|T121|52101|RXNORM|CYCLOBENZAPRINE HYDROCHLORIDE|CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|CLOBEN|CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|3-(5H-DIBENZO(A,D)CYCLOHEPTEN-5-YLIDENE)PROPYL(DIMETHYL)AMMONIUM CHLORIDE|CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|CYCLOFLEX|CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|FR2100873|CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|FLEXIBAN|CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|1-PROPANAMINE, 3-(5H-DIBENZO(A,D)CYCLOHEPTEN-5-YLIDENE)-N,N-DIMETHYL-, HYDROCHLORIDE|CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|10,11DELTA-AMITRIPTYLINE HYDROCHLORIDE|CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|MUSCLE RELAXANTS SKELETAL CYCLOBENZAPRINE HYDROCHLORIDE|CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|CYCLOBENZAPRINE HYDROCHLORIDE |CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|CYCLOBENZAPRINE HYDROCHLORIDE |CYCLOBENZAPRINE HYDROCHLORIDE
C0125988|T121|52101|RXNORM|CYCLOBENZAPRINE HYDROCHLORIDE |CYCLOBENZAPRINE HYDROCHLORIDE
C0063841|T121||RXNORM|(4-CHLOROPHENOXY)ACETIC ACID 2-(1-METHYLETHYL)HYDRAZIDE
C0063841|T121||RXNORM|IPROCLOZIDE
C0063841|T121||RXNORM|P-(CHLOROPHENOXY)ACETIC ACID 2-ISOPROPYLHYDRAZIDE
C0606667|T121||RXNORM|PIROLAZAMIDE
C0606667|T121||RXNORM|HEXAHYDRO-ALPHA,ALPHA-DIPHENYLPYRROLO-(1,2-ALPHA)PYRAZINE-2(1H)-BUTYRAMIDE
C1170746|T121|353108|RXNORM|ESCITALOPRAM OXALATE|ESCITALOPRAM OXALATE
C1170746|T121|353108|RXNORM|5-ISOBENZOFURANCARBONITRILE, 1-(3-(DIMETHYLAMINO)PROPYL)-1-(4-FLUOROPHENYL)-1,3-DIHYDRO-,(1S)-, ETHANEDIOATE(1:1)|ESCITALOPRAM OXALATE
C1170746|T121|353108|RXNORM|ESCITALOPRAM OXALATE |ESCITALOPRAM OXALATE
C1170746|T121|353108|RXNORM|ESCITALOPRAM OXALATE |ESCITALOPRAM OXALATE
C0060188|T121||RXNORM|2-(4-CHLOROPHENYL)-4-METHYL-2,4-PENTANEDIOL
C0060188|T121||RXNORM|FENPENTADIOL
C1881130|T121||RXNORM|IMAFEN
C1882389|T121||RXNORM|PIPOFEZINE
C1881138|T121||RXNORM|IMIPRAMINOXIDE
C1880856|T121||RXNORM|FTORMETAZINE
C0088224|T121||RXNORM|1,3,4,9-TETRAHYDRO-N,N,1-TRIMETHYLINDENO(1,2-C)- PYRAN-1,ETHYLAMINE.HCL
C0088224|T121||RXNORM|PIRANDAMINE HYDROCHLORIDE
C1883593|T121||RXNORM|ZAFULEPTINE
C1883384|T121||RXNORM|TRAZOLOPRIDE
C2347566|T121||RXNORM|CASOPITANT
C2349098|T121||RXNORM|VALDIPROMIDE
C0608826|T121|161203|RXNORM|ACEPROMETAZINE|ACEPROMETAZINE
C0608826|T121|161203|RXNORM|1-(10-(2-(DIMETHYLAMINO)PROPYL)-10H-PHENOTHIAZIN- 2-YL)ETHANONE|ACEPROMETAZINE
C0050721|T121||RXNORM|2-(1-ADAMANTYLAMINO)ETHYL(P-CHLOROPHENOXY)ACETATE
C0050721|T121||RXNORM|ADAFENOXATE
C2347998|T121||RXNORM|AFALANINE
C2347998|T121||RXNORM|ACETYLPHENYLALANINE
C0051694|T121||RXNORM|AMITRIPTYLINE N-OXIDE
C0051694|T121||RXNORM|AMITRIPTYLINOXIDE
C2346789|T121||RXNORM|ANSOXETINE
C2346868|T121||RXNORM|ATIBEPRONE
C2346892|T121||RXNORM|AZALOXAN FUMARATE
C2346896|T121||RXNORM|AZIPRAMINE
C2346971|T121||RXNORM|BAZINAPRINE
C0053072|T121||RXNORM|BEFURALINE
C0053072|T121||RXNORM|N-BENZO(B)FURAN-2-YLCARBONYL-N'-BENZYLPIPERAZINE.HCL
C0053611|T121||RXNORM|1,2-ETHANEDIAMINE, N,N-DIMETHYL-N'-((3-PHENYL-1H-INDOL-1-YL)METHYL)-
C0053611|T121||RXNORM|BINEDALINE
C0053611|T121||RXNORM|BINODALINE
C0054820|T121||RXNORM|2,3-DIHYDRO-4H-1,3-BENZOXAZIN-2-ONE-3-ACETAMIDE
C0054820|T121||RXNORM|2H-1,3-BENZOXAZINE-3(4H)-ACETAMIDE, 2-OXO-
C0054820|T121||RXNORM|4H-3-METHYLCARBOXAMIDE-1,3-BENZOXAZIN-2-ONE
C0054820|T121||RXNORM|CAROXAZONE
C2348381|T121||RXNORM|EFETOZOLE
C2348443|T121||RXNORM|ENEFEXINE
C2348450|T121||RXNORM|ENPRAZEPINE
C0060170|T121||RXNORM|2-(N-BUTYL-O-CHLOROBENZIMIDOYL)-4-CHLOROPHENYL
C0060170|T121||RXNORM|FENGABINE
C0060305|T121||RXNORM|FEZOLAMINE
C0956920|T121||RXNORM|FEZOLAMINE FUMARATE
C0537150|T121||RXNORM|3ALPHA-HYDROXY-3BETA-METHYL-5ALPHA-PREGNAN-20-ONE
C0537150|T121||RXNORM|GANAXOLONE
C2347511|T121||RXNORM|PIBERALINE
C0072207|T121||RXNORM|PROPIZEPIN
C0072207|T121||RXNORM|PROPIZEPINE
C0072207|T121||RXNORM|PYRIDOBENZODIAZEPINE
C0076671|T121||RXNORM|9-ETHYL-4-FLUORO-1-METHYL-7,8,9,10-TETRAHYDROTHIENO(3,2E)PYRIDO(4,3B)INDOLE LACTATE
C0076671|T121||RXNORM|TIFLUCARBINE
C2348815|T121||RXNORM|TRAZIUM ESILATE
C0132764|T121||RXNORM|7-(1,2-DIMETHYLHEPTYL)-2,2-DIMETHYL-4-(4-PYRIDINYL)-2H-1-BENZOPYRAN-5-OL
C0132764|T121||RXNORM|NONABINE
C2347355|T121||RXNORM|NITRAFUDAM HYDROCHLORIDE
C2348183|T121||RXNORM|SEPROXETINE HYDROCHLORIDE
C2348647|T121||RXNORM|TALOPRAM HYDROCHLORIDE
C0076823|T121|38400|RXNORM|ATOMOXETINE|ATOMOXETINE
C0076823|T121|38400|RXNORM|TOMOXETINE|ATOMOXETINE
C0076823|T121|38400|RXNORM|ATOMOXETINE |ATOMOXETINE
C0076823|T121|38400|RXNORM|ATOMOXETINE |ATOMOXETINE
C0051607|T121|17698|RXNORM|10,11-DIHYDRODIBENZO(A,D)CYCLOHEPT-5-ENYL-7-AMINOHEPTANOIC ACID|AMINEPTINE
C0051607|T121|17698|RXNORM|7-((10,11-DIHYDRO-5H-DIBENZO(A,D)CYCLOHEPTEN-5-YL)AMINO)HEPTANOIC ACID|AMINEPTINE
C0051607|T121|17698|RXNORM|AMINEPTIN|AMINEPTINE
C0051607|T121|17698|RXNORM|AMINEPTINE|AMINEPTINE
C2168874|T121||RXNORM|PYRITINOL + CYPROHEPTADINE + VITAMINS 
C2168874|T121||RXNORM|PYRITINOL + CYPROHEPTADINE + VITAMINS
C0071125|T121||RXNORM|PIRANDAMINE
C0600985|T121||RXNORM|1-NAPHTHALENAMINE, 8-CHLORO-1,2,3,4-TETRAHYDRO-5-METHOXY-N,N-DIMETHYL-
C0600985|T121||RXNORM|N,N-DIMETHYL-5-METHOXY-8-CHLORO-1,2,3,4-TETRAHYDRO-1-NAPHTHYLAMINE
C0600985|T121||RXNORM|LOMETRALINE
C0888036|T121||RXNORM|LOMETRALINE HYDROCHLORIDE
C0113211|T121||RXNORM|N-DESMETHYLSERTRALINE
C0113211|T121||RXNORM|N-DEMETHYLSERTRALINE
C0113211|T121||RXNORM|DESMETHYLSERTRALINE
C0113211|T121||RXNORM|DESMETHYLSERTRALINE 
C3650305|T121||RXNORM|ANTIDEPRESSANTS FLUOXETINE
C3650305|T121||RXNORM|ANTIDEPRESSANTS FLUOXETINE 
C3650304|T121||RXNORM|ANTIDEPRESSANTS FLUVOXAMINE
C3650304|T121||RXNORM|ANTIDEPRESSANTS FLUVOXAMINE 
C3650297|T121||RXNORM|ANTIDEPRESSANTS PAROXETINE 
C3650297|T121||RXNORM|ANTIDEPRESSANTS PAROXETINE
C3650299|T121||RXNORM|ANTIDEPRESSANTS NEFAZODONE
C3650299|T121||RXNORM|ANTIDEPRESSANTS NEFAZODONE 
C0068987|T121||RXNORM|DESMETHYLFLUOXETINE
C0068987|T121||RXNORM|NORFLUOXETIN
C0068987|T121||RXNORM|NORFLUOXETINE
C0068987|T121||RXNORM|NORFLUOXETINE 
C0719199|T121|215928|RXNORM|CELEXA|CELEXA
C0719199|T121|215928|RXNORM|CITALOPRAM HYDROBROMIDE (CELEXA)|CELEXA
C0162373|T121|58827|RXNORM|PROZAC|PROZAC
C0376414|T121|114228|RXNORM|PAXIL|PAXIL
C0709644|T121|208161|RXNORM|SERTRALINE 50 MG ORAL TABLET [ZOLOFT]|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 50 MG ORAL TABLET
C0709644|T121|208161|RXNORM|ZOLOFT 50 MG ORAL TABLET|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 50 MG ORAL TABLET
C0709644|T121|208161|RXNORM|ZOLOFT 50MG TABLET|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 50 MG ORAL TABLET
C0709644|T121|208161|RXNORM|ZOLOFT, 50 MG ORAL TABLET|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 50 MG ORAL TABLET
C0709644|T121|208161|RXNORM|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 50 MG ORAL TABLET|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 50 MG ORAL TABLET
C0709644|T121|208161|RXNORM|SERTRALINE HYDROCHLORIDE 50 MG ORAL TABLET, FILM COATED [ZOLOFT]|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 50 MG ORAL TABLET
C0709644|T121|208161|RXNORM|SERTRALINE HYDROCHLORIDE 50 MG ORAL TABLET [ZOLOFT]|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 50 MG ORAL TABLET
C0709632|T121|208149|RXNORM|SERTRALINE 100 MG ORAL TABLET [ZOLOFT]|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 100 MG ORAL TABLET
C0709632|T121|208149|RXNORM|ZOLOFT 100MG TABLET|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 100 MG ORAL TABLET
C0709632|T121|208149|RXNORM|ZOLOFT, 100 MG ORAL TABLET|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 100 MG ORAL TABLET
C0709632|T121|208149|RXNORM|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 100 MG ORAL TABLET|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 100 MG ORAL TABLET
C0709632|T121|208149|RXNORM|SERTRALINE HYDROCHLORIDE 100 MG ORAL TABLET, FILM COATED [ZOLOFT]|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 100 MG ORAL TABLET
C0709632|T121|208149|RXNORM|SERTRALINE HYDROCHLORIDE 100 MG ORAL TABLET [ZOLOFT]|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 100 MG ORAL TABLET
C0709632|T121|208149|RXNORM|ZOLOFT 100 MG ORAL TABLET|ZOLOFT (AS SERTRALINE HYDROCHLORIDE) 100 MG ORAL TABLET
C0284660|T121|82728|RXNORM|ZOLOFT|ZOLOFT
C0284660|T121|82728|RXNORM|ALTRULINE|ZOLOFT
C0284660|T121|82728|RXNORM|PARKE DAVIS BRAND OF SERTRALINE HYDROCHLORIDE|ZOLOFT
C0284660|T121|82728|RXNORM|LUSTRAL|ZOLOFT
C0284660|T121|82728|RXNORM|ROERIG BRAND OF SERTRALINE HYDROCHLORIDE|ZOLOFT
C0284660|T121|82728|RXNORM|PFIZER BRAND OF SERTRALINE HYDROCHLORIDE|ZOLOFT
C0060926|T121|25480|RXNORM|1-(AMINOMETHYL)CYCLOHEXANEACETIC ACID|GABAPENTIN
C0060926|T121|25480|RXNORM|GABAPENTIN|GABAPENTIN
C0060926|T121|25480|RXNORM|GABAPENTIN |GABAPENTIN
C0060926|T121|25480|RXNORM|GABAPENTIN [CHEMICAL/INGREDIENT]|GABAPENTIN
C0060926|T121|25480|RXNORM|CONVALIS|GABAPENTIN
C0060926|T121|25480|RXNORM|GABAPENTIN |GABAPENTIN
C0060926|T121|25480|RXNORM|GABAPENTIN |GABAPENTIN
C0678176|T121|196498|RXNORM|NEURONTIN|NEURONTIN
C0657912|T121|187832|RXNORM|PREGABALIN|PREGABALIN
C0657912|T121|187832|RXNORM|3-(AMINOMETHYL)-5-METHYL-HEXANOIC ACID|PREGABALIN
C0657912|T121|187832|RXNORM|3-ISOBUTYL GABA|PREGABALIN
C0657912|T121|187832|RXNORM|PREGABALIN |PREGABALIN
C0657912|T121|187832|RXNORM|(S+)-3-ISOBUTYL GABA|PREGABALIN
C0657912|T121|187832|RXNORM|(R-)-3-ISOBUTYL GABA|PREGABALIN
C0657912|T121|187832|RXNORM|3-(AMINOMETHYL)-5-METHYLHEXANOIC ACID|PREGABALIN
C0657912|T121|187832|RXNORM|(S)-3-(AMINOMETHYL)-5-METHYLHEXANOIC ACID|PREGABALIN
C0657912|T121|187832|RXNORM|GABA, 3-ISOBUTYL|PREGABALIN
C0657912|T121|187832|RXNORM|3 ISOBUTYL GABA|PREGABALIN
C0657912|T121|187832|RXNORM|PREGABALIN [CHEMICAL/INGREDIENT]|PREGABALIN
C0657912|T121|187832|RXNORM|PREGABALIN |PREGABALIN
C0657912|T121|187832|RXNORM|PREGABALIN |PREGABALIN
C2740401|T121|898715|RXNORM|PREGABALIN 20 MG/ML ORAL SOLUTION|PREGABALIN 20 MG IN 1 ML ORAL SOLUTION
C2740401|T121|898715|RXNORM|PREGABALIN 20MG/ML ORAL SOLUTION|PREGABALIN 20 MG IN 1 ML ORAL SOLUTION
C2740401|T121|898715|RXNORM|PREGABALIN 20MG/ML ORAL SOLUTION |PREGABALIN 20 MG IN 1 ML ORAL SOLUTION
C2740401|T121|898715|RXNORM|PREGABALIN SOLN 20 MG/ML|PREGABALIN 20 MG IN 1 ML ORAL SOLUTION
C2740401|T121|898715|RXNORM|PREGABALIN 20MG ORAL SOLUTION|PREGABALIN 20 MG IN 1 ML ORAL SOLUTION
C2740401|T121|898715|RXNORM|PREGABALIN 20MG/ML SOLN,ORAL|PREGABALIN 20 MG IN 1 ML ORAL SOLUTION
C2740401|T121|898715|RXNORM|PREGABALIN 20MG/ML ORAL SOLN|PREGABALIN 20 MG IN 1 ML ORAL SOLUTION
C2740401|T121|898715|RXNORM|PREGABALIN 20MG/ML SOLN,ORAL [VA PRODUCT]|PREGABALIN 20 MG IN 1 ML ORAL SOLUTION
C1532848|T121|483446|RXNORM|PREGABALIN 200 MG ORAL CAPSULE|PREGABALIN 200 MG ORAL CAPSULE
C1532848|T121|483446|RXNORM|PREGABALIN CAP 200 MG|PREGABALIN 200 MG ORAL CAPSULE
C1532848|T121|483446|RXNORM|PREGABALIN 200MG CAP,ORAL|PREGABALIN 200 MG ORAL CAPSULE
C1532848|T121|483446|RXNORM|PREGABALIN 200MG ORAL CAP|PREGABALIN 200 MG ORAL CAPSULE
C1532848|T121|483446|RXNORM|PREGABALIN 200MG CAP,ORAL [VA PRODUCT]|PREGABALIN 200 MG ORAL CAPSULE
C1532848|T121|483446|RXNORM|PREGABALIN 200MG ORAL CAPSULE|PREGABALIN 200 MG ORAL CAPSULE
C1532848|T121|483446|RXNORM|PREGABALIN 200MG CAPSULE |PREGABALIN 200 MG ORAL CAPSULE
C1532848|T121|483446|RXNORM|PREGABALIN 200MG CAPSULE|PREGABALIN 200 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50 MG ORAL CAPSULE|PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN CAP 50 MG|PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50MG CAP,ORAL|PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50MG ORAL CAP|PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50MG CAP,UD|PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50MG CAP UD|PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50MG CAP,ORAL [VA PRODUCT]|PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50MG CAP,UD [VA PRODUCT]|PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50MG ORAL CAPSULE|PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50MG CAPSULE |PREGABALIN 50 MG ORAL CAPSULE
C1532851|T121|483448|RXNORM|PREGABALIN 50MG CAPSULE|PREGABALIN 50 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75 MG ORAL CAPSULE|PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN CAP 75 MG|PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75MG CAP,ORAL|PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75MG CAP,UD|PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75MG ORAL CAP|PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75MG CAP UD|PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75MG CAP,ORAL [VA PRODUCT]|PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75MG CAP,UD [VA PRODUCT]|PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75MG ORAL CAPSULE|PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75MG CAPSULE |PREGABALIN 75 MG ORAL CAPSULE
C1532852|T121|483450|RXNORM|PREGABALIN 75MG CAPSULE|PREGABALIN 75 MG ORAL CAPSULE
C1532849|T121|483442|RXNORM|PREGABALIN 25 MG ORAL CAPSULE|PREGABALIN 25 MG ORAL CAPSULE
C1532849|T121|483442|RXNORM|PREGABALIN CAP 25 MG|PREGABALIN 25 MG ORAL CAPSULE
C1532849|T121|483442|RXNORM|PREGABALIN 25MG CAP,ORAL|PREGABALIN 25 MG ORAL CAPSULE
C1532849|T121|483442|RXNORM|PREGABALIN 25MG ORAL CAP|PREGABALIN 25 MG ORAL CAPSULE
C1532849|T121|483442|RXNORM|PREGABALIN 25MG CAP,ORAL [VA PRODUCT]|PREGABALIN 25 MG ORAL CAPSULE
C1532849|T121|483442|RXNORM|PREGABALIN 25MG ORAL CAPSULE|PREGABALIN 25 MG ORAL CAPSULE
C1532849|T121|483442|RXNORM|PREGABALIN 25MG CAPSULE |PREGABALIN 25 MG ORAL CAPSULE
C1532849|T121|483442|RXNORM|PREGABALIN 25MG CAPSULE|PREGABALIN 25 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150 MG ORAL CAPSULE|PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN CAP 150 MG|PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150MG CAP,ORAL|PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150MG CAP UD|PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150MG ORAL CAP|PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150MG CAP,UD|PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150MG CAP,ORAL [VA PRODUCT]|PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150MG CAP,UD [VA PRODUCT]|PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150MG ORAL CAPSULE|PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150MG CAPSULE |PREGABALIN 150 MG ORAL CAPSULE
C1532847|T121|483440|RXNORM|PREGABALIN 150MG CAPSULE|PREGABALIN 150 MG ORAL CAPSULE
C0388352|T121||RXNORM|CI 1008
C0388352|T121||RXNORM|CI1008
C0388352|T121||RXNORM|1008, CI
C0388352|T121||RXNORM|CI-1008
C1972026|T121||RXNORM|PREGABALIN &#X7C; BLD-SER-PLAS
C3170841|T121||RXNORM|PREGABALIN &#X7C; URINE
C1570232|T121|593441|RXNORM|LYRICA|LYRICA
C1532846|T121|483438|RXNORM|PREGABALIN 100 MG ORAL CAPSULE|PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN CAP 100 MG|PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN 100MG CAP,ORAL|PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN 100MG CAP,UD|PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN 100MG ORAL CAP|PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN 100MG CAP UD|PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN 100MG CAP,UD [VA PRODUCT]|PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN 100MG CAP,ORAL [VA PRODUCT]|PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN 100MG ORAL CAPSULE|PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN 100MG CAPSULE |PREGABALIN 100 MG ORAL CAPSULE
C1532846|T121|483438|RXNORM|PREGABALIN 100MG CAPSULE|PREGABALIN 100 MG ORAL CAPSULE
C1532850|T121|483444|RXNORM|PREGABALIN 300 MG ORAL CAPSULE|PREGABALIN 300 MG ORAL CAPSULE
C1532850|T121|483444|RXNORM|PREGABALIN CAP 300 MG|PREGABALIN 300 MG ORAL CAPSULE
C1532850|T121|483444|RXNORM|PREGABALIN 300MG CAP,ORAL|PREGABALIN 300 MG ORAL CAPSULE
C1532850|T121|483444|RXNORM|PREGABALIN 300MG ORAL CAP|PREGABALIN 300 MG ORAL CAPSULE
C1532850|T121|483444|RXNORM|PREGABALIN 300MG CAP,ORAL [VA PRODUCT]|PREGABALIN 300 MG ORAL CAPSULE
C1532850|T121|483444|RXNORM|PREGABALIN 300MG ORAL CAPSULE|PREGABALIN 300 MG ORAL CAPSULE
C1532850|T121|483444|RXNORM|PREGABALIN 300MG CAPSULE |PREGABALIN 300 MG ORAL CAPSULE
C1532850|T121|483444|RXNORM|PREGABALIN 300MG CAPSULE|PREGABALIN 300 MG ORAL CAPSULE
C1613977|T121|577127|RXNORM|PREGABALIN 225 MG ORAL CAPSULE|PREGABALIN 225 MG ORAL CAPSULE
C1613977|T121|577127|RXNORM|PREGABALIN CAP 225 MG|PREGABALIN 225 MG ORAL CAPSULE
C1613977|T121|577127|RXNORM|PREGABALIN 225MG CAPSULE |PREGABALIN 225 MG ORAL CAPSULE
C1613977|T121|577127|RXNORM|PREGABALIN 225MG CAPSULE|PREGABALIN 225 MG ORAL CAPSULE
C1613977|T121|577127|RXNORM|PREGABALIN 225MG CAP,ORAL|PREGABALIN 225 MG ORAL CAPSULE
C1613977|T121|577127|RXNORM|PREGABALIN 225MG ORAL CAP|PREGABALIN 225 MG ORAL CAPSULE
C1613977|T121|577127|RXNORM|PREGABALIN 225MG CAP,ORAL [VA PRODUCT]|PREGABALIN 225 MG ORAL CAPSULE
C1613977|T121|577127|RXNORM|PREGABALIN 225MG ORAL CAPSULE|PREGABALIN 225 MG ORAL CAPSULE
C1955823|T121||RXNORM|PD 144723
