C0948762|T034||LNC|ABSOLUTE NEUTROPHIL COUNT
C1168174|T034||LNC|INTERPERTATION, NOT VALUE
C1262264|T034||LNC|ABSOLUTE NEUTROPHIL COUNT ABNORMAL
C1699112|T034||LNC|ABSOLUTE NEUTROPHIL COUNT INCREASED
C0362968|T034|751-8|LNC|NEUTROPHILS # BLD AUTO|NEUTROPHILS [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0948762|T034||LNC|ABSOLUTE NEUTROPHIL COUNT
C0948762|T034||LNC|ANC
C0948762|T034||LNC|BLOOD ABSOLUTE NEUTROPHIL COUNT (ANC)
C0948762|T034||LNC|BLOOD ABSOLUTE NEUTROPHIL COUNT (ANC) 
C0948762|T034||LNC|BLOOD ANC
C0948762|T034||LNC|BLOOD ABSOLUTE NEUTROPHIL COUNT
C0948762|T034||LNC|BLOOD ANC (ABSOLUTE NEUTROPHIL COUNT)
C0948762|T034||LNC|BLOOD ABSOLUTE NEUTROPHIL COUNT 
C0948762|T034||LNC|NEUTROPHILS
C0948762|T034||LNC|NEUT
C1168174|T034||LNC|DECREASED ANC
C1168174|T034||LNC|DECREASED ABSOLUTE NEUTROPHIL COUNT
C1168174|T034||LNC|ABSOLUTE NEUTROPHIL COUNT DECREASED
C1262264|T034||LNC|ABSOLUTE NEUTROPHIL COUNT ABNORMAL
C1699112|T034||LNC|ABSOLUTE NEUTROPHIL COUNT INCREASED
C0362968|T034|751-8|LNC|NEUTROPHILS|NEUTROPHILS [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0362968|T034|751-8|LNC|NEUTROPHILS VOLUME IN BLOOD BY AUTOMATED COUNT|NEUTROPHILS [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0362968|T034|751-8|LNC|NEUTROPHILS NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:WHOLE BLOOD:QUANTITATIVE:AUTOMATED COUNT|NEUTROPHILS [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0362968|T034|751-8|LNC|NEUTROPHILS NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:WHOLE BLOOD:QUANTITATIVE:AUTOMATED COUNT|NEUTROPHILS [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
