C1399448|T037||SNOMEDCT_US|BIRTH TO AN HCV-INFECTED MOTHER
C1399448|T037||SNOMEDCT_US|BORN WITH HCV
C1399448|T037||SNOMEDCT_US|MOTHER HAS HCV
C1399448|T037||SNOMEDCT_US|MOTHER HAD HCV
C1399448|T037||SNOMEDCT_US|MATERNAL; HEPATITIS, AFFECTING FETUS
C1399448|T037||SNOMEDCT_US|HEPATITIS; MATERNAL, AFFECTING FETUS
C1399448|T037||SNOMEDCT_US|MATERNAL; HEPATITIS, AFFECTING FETUS
