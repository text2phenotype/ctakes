C2367818|T061|304150|MEDCIN|HEPATITIS C TREATMENT PRESCRIBED|HEPATITIS C TREATMENT PRESCRIBED (TREATMENT)
C2367822|T061|304154|MEDCIN|PEGINTERFERON AND RIBAVIRIN THERAPY PRESCRIBED FOR HEPATITIS C|PEGINTERFERON AND RIBAVIRIN THERAPY PRESCRIBED FOR HEPATITIS C (TREATMENT)
C2750389|T061||MEDCIN|HEPATITIS C VIRUS INFECTION, RESPONSE TO THERAPY OF
C2750389|T061||MEDCIN|PREVIOUS HCV TREATMENT
C2750389|T061||MEDCIN|PREVIOUSLY TREATED FOR HCV
C2750389|T061||MEDCIN|PREVIOUS TREATMENT FOR HCV
C2750389|T061||MEDCIN|PREVIOUS HCV TREATMEN
C2367819|T061|304151|MEDCIN|ANTIVIRAL HEPATITIS C TREATMENT|ANTIVIRAL HEPATITIS C TREATMENT BEING RECEIVED (TREATMENT)
C2367819|T061|304151|MEDCIN|ANTIVIRAL HEPATITIS C TREATMENT BEING RECEIVED |ANTIVIRAL HEPATITIS C TREATMENT BEING RECEIVED (TREATMENT)
C2367819|T061|304151|MEDCIN|ANTIVIRAL HEPATITIS C TREATMENT BEING RECEIVED|ANTIVIRAL HEPATITIS C TREATMENT BEING RECEIVED (TREATMENT)
C2367822|T061|304154|MEDCIN|PEGINTERFERON|PEGINTERFERON
C2367822|T061|304154|MEDCIN|RIBAVIRIN|PEGINTERFERON
C2367822|T061|304154|MEDCIN|PEGINTERFERON AND RIBAVIRIN THERAPY PRESCRIBED FOR HEPATITIS C |PEGINTERFERON AND RIBAVIRIN THERAPY PRESCRIBED FOR HEPATITIS C (TREATMENT)
C2367822|T061|304154|MEDCIN|PEGINTERFERON AND RIBAVIRIN THERAPY PRESCRIBED FOR HEPATITIS C|PEGINTERFERON AND RIBAVIRIN THERAPY PRESCRIBED FOR HEPATITIS C (TREATMENT)
