C1274583|T053|403182006|SNOMEDCT_US|NON-PROFESSIONAL TATTOO|AMATEUR DECORATIVE TATTOO OF SKIN
C1274583|T053|403182006|SNOMEDCT_US|AMATEUR TATTOO|AMATEUR DECORATIVE TATTOO OF SKIN
C1274583|T053|403182006|SNOMEDCT_US|TATTOO DIRTY|AMATEUR DECORATIVE TATTOO OF SKIN
