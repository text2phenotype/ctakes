C0484660|T201|10466-1|LNC|ANION GAP3 SERPL-SCNC|ANION GAP 3 IN SERUM OR PLASMA
C0484683|T201|9830-1|LNC|CHOLEST/HDLC SERPL-MRTO|CHOLESTEROL.TOTAL/CHOLESTEROL IN HDL [MASS RATIO] IN SERUM OR PLASMA
C0942468|T201|26508-2|LNC|NEUTS BAND NFR BLD|BAND FORM NEUTROPHILS/100 LEUKOCYTES IN BLOOD
C0484430|T201|6690-2|LNC|WBC # BLD AUTO|LEUKOCYTES [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0942471|T201|26511-6|LNC|NEUTROPHILS NFR BLD|NEUTROPHILS/100 LEUKOCYTES IN BLOOD
C0366777|T201|4544-3|LNC|HCT VFR BLD AUTO|HCT VFR BLD AUTO
C0364121|T201|1988-5|LNC|CRP SERPL-MCNC|C REACTIVE PROTEIN [MASS/VOLUME] IN SERUM OR PLASMA
C0944746|T201|29265-6|LNC|CALCIUM ALBUM COR SERPL-SCNC|CALCIUM [MOLES/VOLUME] CORRECTED FOR ALBUMIN IN SERUM OR PLASMA
C1526484|T201|38483-4|LNC|CREAT BLD-MCNC|CREATININE [MASS/VOLUME] IN BLOOD
C0366770|T201|4537-7|LNC|ESR BLD QN WESTRGRN|ERYTHROCYTE SEDIMENTATION RATE BY WESTERGREN METHOD
C0484448|T201|10378-8|LNC|POLYCHROMASIA BLD QL SMEAR|POLYCHROMASIA [PRESENCE] IN BLOOD BY LIGHT MICROSCOPY
C0802588|T201|19773-1|LNC|RECOM F/U CVX/VAG CYTO|RECOMMENDED FOLLOW-UP [IDENTIFIER] IN CERVICAL OR VAGINAL SMEAR OR SCRAPING BY CYTO STAIN
C0484652|T201|1798-8|LNC|AMYLASE SERPL-CCNC|AMYLASE [ENZYMATIC ACTIVITY/VOLUME] IN SERUM OR PLASMA
C0363117|T201|925-8|LNC|BLD PROD DISPOSITION BPU|BLOOD PRODUCT DISPOSITION [TYPE]
C0482158|T201|933-2|LNC|BLD PROD TYP BPU|BLD PROD TYP BPU
C1315182|T201|32623-1|LNC|PMV BLD AUTO|PMV BLD AUTO
C0365091|T201|2947-0|LNC|SODIUM BLD-SCNC|SODIUM [MOLES/VOLUME] IN BLOOD
C0942474|T201|26515-7|LNC|PLATELET # BLD|PLATELETS [#/VOLUME] IN BLOOD
C1714656|T201|43304-5|LNC|C TRACH RRNA XXX QL PCR|C TRACH RRNA XXX QL NAA+PROBE
C1114891|T201|30341-2|LNC|ESR BLD QN|ESR BLD QN
C0942447|T201|26485-3|LNC|MONOCYTES NFR BLD|MONOCYTES/100 LEUKOCYTES IN BLOOD
C1954900|T201|49136-5|LNC|CK MB SERPL-RTO|CREATINE KINASE.MB/CREATINE KINASE.TOTAL [RATIO] IN SERUM OR PLASMA
C0367784|T201|3393-6|LNC|BZE UR QL|BENZOYLECGONINE [PRESENCE] IN URINE
C0364160|T201|2028-9|LNC|CO2 SERPL-SCNC|CARBON DIOXIDE, TOTAL [MOLES/VOLUME] IN SERUM OR PLASMA
C0368036|T201|5821-4|LNC|WBC #/AREA URNS HPF|WBC #/AREA URNS HPF
C0485610|T201|10701-1|LNC|O+P STL CONC|OVA AND PARASITES IDENTIFIED IN STOOL BY CONCENTRATION
C0362968|T201|751-8|LNC|NEUTROPHILS # BLD AUTO|NEUTROPHILS [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0364459|T201|2324-2|LNC|GGT SERPL-CCNC|GAMMA GLUTAMYL TRANSFERASE [ENZYMATIC ACTIVITY/VOLUME] IN SERUM OR PLASMA
C1507842|T201|35691-5|LNC|OTHER MICROORGANISM DNA XXX QL PCR|OTHER MICROORG DNA XXX QL NAA+PROBE
C0364714|T201|2571-8|LNC|TRIGL SERPL-MCNC|TRIGL SERPL-MCNC
C0364225|T201|2089-1|LNC|LDLC SERPL-MCNC|CHOLESTEROL IN LDL [MASS/VOLUME] IN SERUM OR PLASMA
C0365195|T201|3051-0|LNC|T3FREE SERPL-MCNC|TRIIODOTHYRONINE (T3) FREE [MASS/VOLUME] IN SERUM OR PLASMA
C0802583|T201|19767-3|LNC|CYTOLOGIST CVX/VAG CYTO|CYTOLOGIST WHO READ CYTO STAIN OF CERVICAL OR VAGINAL SMEAR OR SCRAPING
C0365609|T201|3377-9|LNC|BARBITURATES UR QL|BARBITURATES [PRESENCE] IN URINE
C1714740|T201|43396-1|LNC|NONHDLC SERPL-MCNC|CHOLESTEROL NON HDL [MASS/VOLUME] IN SERUM OR PLASMA
C0368555|T201|624-7|LNC|BACTERIA SPT RESP CULT|BACTERIA IDENTIFIED IN SPUTUM BY RESPIRATORY CULTURE
C1369580|T201|34714-6|LNC|INR BLD|INR BLD
C0802028|T201|19080-1|LNC|HCG SERPL-ACNC|CHORIOGONADOTROPIN [UNITS/VOLUME] IN SERUM OR PLASMA
C0942414|T201|26444-0|LNC|BASOPHILS # BLD|BASOPHILS [#/VOLUME] IN BLOOD
C0798369|T201|15198-5|LNC|MACROCYTES BLD QL AUTO|MACROCYTES [PRESENCE] IN BLOOD BY AUTOMATED COUNT
C0881426|T201|24111-7|LNC|N GONORRHOEA DNA XXX QL PCR|NEISSERIA GONORRHOEAE DNA [PRESENCE] IN UNSPECIFIED SPECIMEN BY NAA WITH PROBE DETECTION
C0368530|T201|600-7|LNC|BACTERIA BLD CULT|BACTERIA IDENTIFIED IN BLOOD BY CULTURE
C0485832|T201|8061-4|LNC|ANA SER QL|NUCLEAR AB [PRESENCE] IN SERUM
C0942419|T201|26449-9|LNC|EOSINOPHIL # BLD|EOSINOPHILS [#/VOLUME] IN BLOOD
C0365237|T201|6299-2|LNC|BUN BLD-MCNC|UREA NITROGEN [MASS/VOLUME] IN BLOOD
C0550447|T201|11558-4|LNC|PH BLD|PH BLD
C0803434|T201|20629-2|LNC|LEVOFLOXACIN SUSC ISLT|LEVOFLOXACIN [SUSCEPTIBILITY]
C1316366|T201|33903-6|LNC|KETONES UR QL|KETONES [PRESENCE] IN URINE
C0367985|T201|5770-3|LNC|BILIRUB UR QL STRIP|BILIRUB UR QL STRIP
C0877807|T201|1003-3|LNC|IAT COMP-SP REAG SERPL QL|INDIRECT ANTIGLOBULIN TEST.COMPLEMENT SPECIFIC REAGENT [PRESENCE] IN SERUM OR PLASMA
C0942461|T201|26499-4|LNC|NEUTROPHILS # BLD|NEUTROPHILS [#/VOLUME] IN BLOOD
C0364127|T201|1994-3|LNC|CA-I BLD-SCNC|CALCIUM.IONIZED [MOLES/VOLUME] IN BLOOD
C0482131|T201|883-9|LNC|ABO GROUP BLD|ABO GROUP [TYPE] IN BLOOD
C0549842|T201|11125-2|LNC|PLAT MORPH BLD|PLATELET MORPHOLOGY FINDING [IDENTIFIER] IN BLOOD
C0550528|T201|11580-8|LNC|TSH SERPL DL<=0.005 MIU/L-ACNC|THYROTROPIN:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DETECTION LIMIT <= 0.005 MIU/L
C0802579|T201|19763-2|LNC|SPECIMEN SOURCE CVX/VAG CYTO|SPECIMEN SOURCE [IDENTIFIER] IN CERVICAL OR VAGINAL SMEAR OR SCRAPING BY CYTO STAIN
C0367982|T201|5767-9|LNC|APPEARANCE UR|APPEARANCE UR
C0368020|T201|5794-3|LNC|HGB UR QL STRIP|HEMOGLOBIN [PRESENCE] IN URINE BY TEST STRIP
C0362947|T201|731-0|LNC|LYMPHOCYTES # BLD AUTO|LYMPHOCYTES [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0362981|T201|764-1|LNC|NEUTS BAND NFR BLD MANUAL|BAND FORM NEUTROPHILS/100 LEUKOCYTES IN BLOOD BY MANUAL COUNT
C0802580|T201|19764-0|LNC|STAT OF ADQ CVX/VAG CYTO-IMP|STATEMENT OF ADEQUACY [INTERPRETATION] OF CERVICAL OR VAGINAL SMEAR OR SCRAPING BY CYTO STAIN
C0803797|T201|21000-5|LNC|RDW RBC AUTO|ERYTHROCYTE DISTRIBUTION WIDTH [ENTITIC VOLUME] BY AUTOMATED COUNT
C0550221|T201|11555-0|LNC|BASE EXCESS BLD-SCNC|BASE EXCESS IN BLOOD BY CALCULATION
C0550440|T201|11556-8|LNC|PO2 BLD|PO2 BLD
C0362952|T201|736-9|LNC|LYMPHOCYTES NFR BLD AUTO|LYMPHOCYTES/100 LEUKOCYTES IN BLOOD BY AUTOMATED COUNT
C0802522|T201|19659-2|LNC|PCP UR QL SCN|PHENCYCLIDINE [PRESENCE] IN URINE BY SCREEN METHOD
C0364122|T201|1989-3|LNC|25(OH)D3 SERPL-MCNC|25(OH)D3 SERPL-MCNC
C0364874|T201|2731-8|LNC|PTH-INTACT SERPL-MCNC|PTH-INTACT SERPL-MCNC
C0364655|T201|2514-8|LNC|KETONES UR QL STRIP|KETONES [PRESENCE] IN URINE BY TEST STRIP
C0549856|T201|12258-0|LNC|SQUAMOUS URNS QL MICRO|EPITHELIAL CELLS.SQUAMOUS [PRESENCE] IN URINE SEDIMENT BY LIGHT MICROSCOPY
C0362958|T201|742-7|LNC|MONOCYTES # BLD AUTO|MONOCYTES [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0368042|T201|5803-2|LNC|PH UR STRIP|PH OF URINE BY TEST STRIP
C0362957|T201|741-9|LNC|MICROCYTES BLD QL SMEAR|MICROCYTES [PRESENCE] IN BLOOD BY LIGHT MICROSCOPY
C1831574|T201|47527-7|LNC|CYTOLOGY CVX/VAG DOC THIN PREP|CYTOLOGY REPORT OF CERVICAL OR VAGINAL SMEAR OR SCRAPING CYTO STAIN.THIN PREP
C0364207|T201|2075-0|LNC|CHLORIDE SERPL-SCNC|CHLORIDE [MOLES/VOLUME] IN SERUM OR PLASMA
C0362987|T201|770-8|LNC|NEUTROPHILS NFR BLD AUTO|NEUTROPHILS/100 LEUKOCYTES IN BLOOD BY AUTOMATED COUNT
C0368011|T201|5787-7|LNC|EPI CELLS #/AREA URNS HPF|EPI CELLS #/AREA URNS HPF
C0801991|T201|18998-5|LNC|TMP SMX SUSC ISLT|TRIMETHOPRIM+SULFAMETHOXAZOLE [SUSCEPTIBILITY]
C0365095|T201|2951-2|LNC|SODIUM SERPL-SCNC|SODIUM [MOLES/VOLUME] IN SERUM OR PLASMA
C0801308|T201|18262-6|LNC|LDLC SERPL DIRECT ASSAY-MCNC|CHOLESTEROL IN LDL [MASS/VOLUME] IN SERUM OR PLASMA BY DIRECT ASSAY
C1315522|T201|33051-4|LNC|RBC UR QL|ERYTHROCYTES [PRESENCE] IN URINE
C0365170|T201|3026-2|LNC|T4 SERPL-MCNC|THYROXINE (T4) [MASS/VOLUME] IN SERUM OR PLASMA
C0368403|T201|5195-3|LNC|HBV SURFACE AG SER QL|HEPATITIS B VIRUS SURFACE AG [PRESENCE] IN SERUM
C0798130|T201|14957-5|LNC|MICROALBUMIN UR-MCNC|MICROALBUMIN [MASS/VOLUME] IN URINE
C1114261|T201|30405-5|LNC|WBC # UR|LEUKOCYTES [#/VOLUME] IN URINE
C0803374|T201|20565-8|LNC|CO2 BLD-SCNC|CARBON DIOXIDE, TOTAL [MOLES/VOLUME] IN BLOOD
C0365253|T201|3107-0|LNC|UROBILINOGEN UR-MCNC|UROBILINOGEN:MCNC:PT:URINE:QN
C0368404|T201|5196-1|LNC|HBV SURFACE AG SER QL EIA|HEPATITIS B VIRUS SURFACE ANTIGEN:PRESENCE OR THRESHOLD:POINT IN TIME:SERUM/PLASMA:ORDINAL:ENZYME IMMUNOASSAY
C0362900|T201|711-2|LNC|EOSINOPHIL # BLD AUTO|EOSINOPHILS [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0368406|T201|5198-7|LNC|HCV AB SER EIA-ACNC|HEPATITIS C VIRUS AB [UNITS/VOLUME] IN SERUM BY IMMUNOASSAY
C0551356|T201|11572-5|LNC|RHEUMATOID FACT SER-ACNC|RHEUMATOID FACTOR:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C0364092|T201|1959-6|LNC|HCO3 BLD-SCNC|BICARBONATE [MOLES/VOLUME] IN BLOOD
C0364419|T201|2284-8|LNC|FOLATE SERPL-MCNC|FOLATE:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C0368043|T201|5804-0|LNC|PROT UR STRIP-MCNC|PROTEIN [MASS/VOLUME] IN URINE BY TEST STRIP
C0364201|T201|2069-3|LNC|CHLORIDE BLD-SCNC|CHLORIDE [MOLES/VOLUME] IN BLOOD
C0364708|T201|2093-3|LNC|CHOLEST SERPL-MCNC|CHOLESTEROL [MASS/VOLUME] IN SERUM OR PLASMA
C0364641|T201|2500-7|LNC|TIBC SERPL-MCNC|TIBC SERPL-MCNC
C1632381|T201|42931-6|LNC|C TRACH RRNA UR QL PCR|CHLAMYDIA TRACHOMATIS RRNA [PRESENCE] IN URINE BY NAA WITH PROBE DETECTION
C1953859|T201|48346-1|LNC|HIV 1+O+2 AB SERPL-ACNC|HIV 1+O+2 AB [UNITS/VOLUME] IN SERUM OR PLASMA
C0550258|T201|11054-4|LNC|LDLC/HDLC SERPL-MRTO|CHOLESTEROL IN LDL/CHOLESTEROL IN HDL [MASS RATIO] IN SERUM OR PLASMA
C0802029|T201|13362-9|LNC|COLLECT DURATION TIME UR|COLLECT DURATION TIME UR
C1714657|T201|43305-2|LNC|N GONORRHOEA RRNA XXX QL PCR|NEISSERIA GONORRHOEAE RRNA [PRESENCE] IN UNSPECIFIED SPECIMEN BY NAA WITH PROBE DETECTION
C0549795|T201|11282-1|LNC|TOTAL CELLS COUNTED BLD|TOTAL CELLS COUNTED BLD
C0362991|T201|774-0|LNC|OVALOCYTES BLD QL SMEAR|OVALOCYTES [PRESENCE] IN BLOOD BY LIGHT MICROSCOPY
C0368032|T201|5797-6|LNC|KETONES UR STRIP-MCNC|KETONES [MASS/VOLUME] IN URINE BY TEST STRIP
C0798351|T201|15180-3|LNC|HYPOCHROMIA BLD QL AUTO|HYPOCHROMIA [PRESENCE] IN BLOOD BY AUTOMATED COUNT
C2599173|T201|53925-4|LNC|C TRACH RRNA URTH QL PCR|CHLAMYDIA TRACHOMATIS RRNA [PRESENCE] IN URETHRA BY NAA WITH PROBE DETECTION
C0362994|T201|777-3|LNC|PLATELET # BLD AUTO|PLATELETS [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0482130|T201|882-1|LNC|ABO+RH GP BLD|ABO AND RH GROUP [TYPE] IN BLOOD
C0945357|T201|26464-8|LNC|WBC # BLD|LEUKOCYTES [#/VOLUME] IN BLOOD
C0363413|T201|1250-0|LNC|MAJ XM SERPL-IMP|MAJOR CROSSMATCH [INTERPRETATION]
C0362910|T201|789-8|LNC|RBC # BLD AUTO|ERYTHROCYTES [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0365160|T201|3016-3|LNC|TSH SERPL-ACNC|THYROTROPIN [UNITS/VOLUME] IN SERUM OR PLASMA
C0484424|T201|6742-1|LNC|RBC MORPH BLD|RBC MORPH BLD
C1146785|T201|31100-1|LNC|HCT VFR BLD IMPED|HCT VFR BLD IMPED
C0364104|T201|35192-4|LNC|BILIRUB INDIRECT SERPL-MCNC|BILIRUBIN.INDIRECT [MASS OR MOLES/VOLUME] IN SERUM OR PLASMA
C0364887|T201|2744-1|LNC|PH BLDA|PH BLDA
C0362908|T201|787-2|LNC|MCV RBC AUTO|MCV RBC AUTO
C0364474|T201|2336-6|LNC|GLOBULIN SER-MCNC|GLOBULIN [MASS/VOLUME] IN SERUM
C0367244|T201|6463-4|LNC|BACTERIA XXX CULT|BACTERIA IDENTIFIED IN UNSPECIFIED SPECIMEN BY CULTURE
C0364605|T201|2465-3|LNC|IGG SER-MCNC|IMMUNOGLOBULIN G:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C0803318|T201|20507-0|LNC|RPR SER QL|REAGIN AB [PRESENCE] IN SERUM BY RPR
C0802082|T201|19161-9|LNC|UROBILINOGEN UR STRIP-ACNC|UROBILINOGEN [UNITS/VOLUME] IN URINE BY TEST STRIP
C2970099|T201|60256-5|LNC|N GONORRHOEA RRNA UR QL PCR|N GONORRHOEA RRNA UR QL NAA+PROBE
C0368563|T201|630-4|LNC|BACTERIA UR CULT|BACTERIA IDENTIFIED IN URINE BY CULTURE
C0802585|T201|19769-9|LNC|PATHOLOGIST CVX/VAG CYTO|PATHOLOGIST WHO READ CYTO STAIN OF CERVICAL OR VAGINAL SMEAR OR SCRAPING
C0550349|T201|10834-0|LNC|GLOBULIN SER CALC-MCNC|GLOBULIN [MASS/VOLUME] IN SERUM BY CALCULATION
C0365392|T201|3173-2|LNC|APTT TIME BLD|APTT BLD
C0364290|T201|2157-6|LNC|CK SERPL-CCNC|CREATINE KINASE [ENZYMATIC ACTIVITY/VOLUME] IN SERUM OR PLASMA
C0362890|T201|702-1|LNC|ANISOCYTOSIS BLD QL SMEAR|ANISOCYTOSIS [PRESENCE] IN BLOOD BY LIGHT MICROSCOPY
C0482608|T201|3184-9|LNC|ACT TIME BLD|ACT BLD
C0798321|T201|15150-6|LNC|ANISOCYTOSIS BLD QL AUTO|ANISOCYTOSIS [PRESENCE] IN BLOOD BY AUTOMATED COUNT
C0362933|T201|728-6|LNC|HYPOCHROMIA BLD QL SMEAR|HYPOCHROMIA [PRESENCE] IN BLOOD BY LIGHT MICROSCOPY
C0551499|T201|12454-5|LNC|AMORPH URATE CRY URNS QL MICRO|URATE CRYSTALS AMORPHOUS [PRESENCE] IN URINE SEDIMENT BY LIGHT MICROSCOPY
C1114065|T201|30180-4|LNC|BASOPHILS NFR BLD|BASOPHILS/100 LEUKOCYTES IN BLOOD
C0362960|T201|5905-5|LNC|MONOCYTES NFR BLD AUTO|MONOCYTES/100 LEUKOCYTES IN BLOOD BY AUTOMATED COUNT
C0945354|T201|26450-7|LNC|EOSINOPHIL NFR BLD|EOSINOPHILS/100 LEUKOCYTES IN BLOOD
C0550265|T201|13458-5|LNC|VLDLC SERPL CALC-MCNC|CHOLESTEROL IN VLDL [MASS/VOLUME] IN SERUM OR PLASMA BY CALCULATION
C0801360|T201|18314-5|LNC|MORPHOLOGY BLD-IMP|MORPHOLOGY [INTERPRETATION] IN BLOOD NARRATIVE
C0362954|T201|738-5|LNC|MACROCYTES BLD QL SMEAR|MACROCYTES [PRESENCE] IN BLOOD BY LIGHT MICROSCOPY
C0368013|T201|5808-1|LNC|RBC # URNS HPF|ERYTHROCYTES [#/VOLUME] IN URINE SEDIMENT BY MICROSCOPY HIGH POWER FIELD
C0364674|T201|2532-0|LNC|LDH SERPL-CCNC|LACTATE DEHYDROGENASE [ENZYMATIC ACTIVITY/VOLUME] IN SERUM OR PLASMA
C0943165|T201|27353-2|LNC|EST. AVERAGE GLUCOSE BLD GHB EST-MCNC|GLUCOSE MEAN VALUE [MASS/VOLUME] IN BLOOD ESTIMATED FROM GLYCATED HEMOGLOBIN
C0364968|T201|2823-3|LNC|POTASSIUM SERPL-SCNC|POTASSIUM [MOLES/VOLUME] IN SERUM OR PLASMA
C0365197|T201|3053-6|LNC|T3 SERPL-MCNC|TRIIODOTHYRONINE (T3) [MASS/VOLUME] IN SERUM OR PLASMA
C0367857|T201|5671-3|LNC|LEAD BLD-MCNC|LEAD [MASS/VOLUME] IN BLOOD
C0366781|T201|4548-4|LNC|HGB A1C MFR BLD|HEMOGLOBIN A1C/HEMOGLOBIN.TOTAL IN BLOOD
C0365032|T201|2888-6|LNC|PROT UR-MCNC|PROTEIN [MASS/VOLUME] IN URINE
C0368002|T201|5778-6|LNC|COLOR UR|COLOR:TYPE:PT:URINE:NOM
C0365240|T201|3094-0|LNC|BUN SERPL-MCNC|BUN SERPL-MCNC
C1953857|T201|48345-3|LNC|HIV 1+O+2 AB SERPL QL|HIV 1+O+2 AB [PRESENCE] IN SERUM OR PLASMA
C0367235|T201|6462-6|LNC|BACTERIA WND CULT|BACTERIA IDENTIFIED IN WOUND BY CULTURE
C0550246|T201|11557-6|LNC|PCO2 BLD|PCO2 BLD
C0365243|T201|3097-3|LNC|BUN/CREAT SERPL-MRTO|UREA NITROGEN/CREATININE [MASS RATIO] IN SERUM OR PLASMA
C0366908|T201|4679-7|LNC|RETICS/100 RBC NFR|RETICULOCYTES/100 ERYTHROCYTES:NUMBER FRACTION:POINT IN TIME:WHOLE BLOOD:QUANTITATIVE
C0802148|T201|19244-3|LNC|CHARACTER UR|CHARACTER OF URINE
C0801921|T201|18928-2|LNC|GENTAMICIN SUSC ISLT|GENTAMICIN [SUSCEPTIBILITY]
C0945362|T201|26507-4|LNC|NEUTS BAND # BLD|BAND FORM NEUTROPHILS [#/VOLUME] IN BLOOD
C0367237|T201|634-6|LNC|BACTERIA XXX AEROBE CULT|BACTERIA IDENTIFIED IN UNSPECIFIED SPECIMEN BY AEROBE CULTURE
C0365194|T201|3050-2|LNC|T3RU NFR SERPL|T3RU NFR SERPL
C0362907|T201|786-4|LNC|MCHC RBC AUTO-MCNC|MCHC RBC AUTO-MCNC
C0803267|T201|20453-7|LNC|EPI CELLS URNS QL MICRO|EPITHELIAL CELLS [PRESENCE] IN URINE SEDIMENT BY LIGHT MICROSCOPY
C0364378|T201|35207-0|LNC|ESTRADIOL SERPL-MCNC|ESTRADIOL SERPL-MSCNC
C0364236|T201|2106-3|LNC|HCG PREG UR QL|HCG PREG UR QL
C1145645|T201|2703-7|LNC|PO2 BLDA|PO2 BLDA
C1114184|T201|30313-1|LNC|HGB BLDA-MCNC|HEMOGLOBIN [MASS/VOLUME] IN ARTERIAL BLOOD
C0362895|T201|707-0|LNC|BASOPHILS NFR BLD MANUAL|BASOPHILS/100 LEUKOCYTES IN BLOOD BY MANUAL COUNT
C0365000|T201|2857-1|LNC|PSA SERPL-MCNC|PROSTATE SPECIFIC AG [MASS/VOLUME] IN SERUM OR PLASMA
C1114281|T201|30428-7|LNC|MCV RBC|ERYTHROCYTE MEAN CORPUSCULAR VOLUME:ENTITIC VOLUME:POINT IN TIME:ERYTHROCYTES:QUANTITATIVE
C0803268|T201|20454-5|LNC|PROT UR QL STRIP|PROTEIN [PRESENCE] IN URINE BY TEST STRIP
C0363876|T201|1742-6|LNC|ALT SERPL-CCNC|ALANINE AMINOTRANSFERASE [ENZYMATIC ACTIVITY/VOLUME] IN SERUM OR PLASMA
C0364411|T201|2276-4|LNC|FERRITIN SERPL-MCNC|FERRITIN SERPL-MCNC
C0364221|T201|2085-9|LNC|HDLC SERPL-MCNC|HDLC SERPL-MCNC
C0484638|T201|6768-6|LNC|ALP SERPL-CCNC|ALKALINE PHOSPHATASE [ENZYMATIC ACTIVITY/VOLUME] IN SERUM OR PLASMA
C0368035|T201|5799-2|LNC|LEUKOCYTE ESTERASE UR QL STRIP|LEUKOCYTE ESTERASE UR QL STRIP
C0942446|T201|26484-6|LNC|MONOCYTES # BLD|MONOCYTES [#/VOLUME] IN BLOOD
C1315508|T201|33037-3|LNC|ANION GAP SERPL-SCNC|ANION GAP IN SERUM OR PLASMA
C0368018|T201|5792-7|LNC|GLUCOSE UR STRIP-MCNC|GLUCOSE [MASS/VOLUME] IN URINE BY TEST STRIP
C0804406|T201|21613-5|LNC|C TRACH DNA XXX QL PCR|CHLAMYDIA TRACHOMATIS DNA [PRESENCE] IN UNSPECIFIED SPECIMEN BY NAA WITH PROBE DETECTION
C0364151|T201|2019-8|LNC|PCO2 BLDA|PCO2 BLDA
C0797519|T201|14338-8|LNC|PREALB SERPL-MCNC|PREALBUMIN [MASS/VOLUME] IN SERUM OR PLASMA
C0942440|T201|26478-8|LNC|LYMPHOCYTES NFR BLD|LYMPHOCYTES/100 LEUKOCYTES IN BLOOD
C0364128|T201|1995-0|LNC|CA-I SERPL-SCNC|CALCIUM.IONIZED [MOLES/VOLUME] IN SERUM OR PLASMA
C0945446|T201|27045-4|LNC|MICROSCOPIC UR-IMP|MICROSCOPIC EXAM [INTERPRETATION] OF URINE BY CYTOLOGY
C0801328|T201|18282-4|LNC|CANNABINOIDS UR QL SCN|CANNABINOIDS [PRESENCE] IN URINE BY SCREEN METHOD
C0484447|T201|9317-9|LNC|PLATELET BLD QL SMEAR|PLATELET BLD QL SMEAR
C0362894|T201|706-2|LNC|BASOPHILS NFR BLD AUTO|BASOPHILS/100 LEUKOCYTES IN BLOOD BY AUTOMATED COUNT
C0365228|T201|3084-1|LNC|URATE SERPL-MCNC|URATE SERPL-MCNC
C0484796|T201|10501-5|LNC|LH SERPL-ACNC|LUTROPIN [UNITS/VOLUME] IN SERUM OR PLASMA
C0363081|T201|890-4|LNC|BLD GP AB SCN SERPL QL|BLOOD GROUP ANTIBODY SCREEN [PRESENCE] IN SERUM OR PLASMA
C0362961|T201|744-3|LNC|MONOCYTES NFR BLD MANUAL|MONOCYTES/100 LEUKOCYTES IN BLOOD BY MANUAL COUNT
C0367338|T201|664-3|LNC|GRAM STN XXX|MICROSCOPIC OBSERVATION [IDENTIFIER] IN UNSPECIFIED SPECIMEN BY GRAM STAIN
C0362953|T201|737-7|LNC|LYMPHOCYTES NFR BLD MANUAL|LYMPHOCYTES/100 LEUKOCYTES IN BLOOD BY MANUAL COUNT
C0482694|T201|5902-2|LNC|PT TIME PPP|COAGULATION TISSUE FACTOR INDUCED:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0550543|T201|10839-9|LNC|TROPONIN I SERPL-MCNC|TROPONIN I.CARDIAC [MASS/VOLUME] IN SERUM OR PLASMA
C0362903|T201|714-6|LNC|EOSINOPHIL NFR BLD MANUAL|EOSINOPHILS/100 LEUKOCYTES IN BLOOD BY MANUAL COUNT
C0803379|T201|20570-8|LNC|HCT VFR BLD|HCT VFR BLD
C0482705|T201|3255-7|LNC|FIBRINOGEN PPP-MCNC|FIBRINOGEN [MASS/VOLUME] IN PLATELET POOR PLASMA BY COAGULATION ASSAY
C0364639|T201|2498-4|LNC|IRON SERPL-MCNC|IRON SERPL-MCNC
C0364612|T201|2472-9|LNC|IGM SER-MCNC|IGM [MASS/VOLUME] IN SERUM OR PLASMA
C1114721|T201|30934-4|LNC|BNP SERPL-MCNC|BNP SERPL-MCNC
C0363885|T201|1751-7|LNC|ALBUMIN SERPL-MCNC|ALBUMIN [MASS/VOLUME] IN SERUM OR PLASMA
C0798152|T201|14979-9|LNC|APTT TIME PPP|APTT PPP
C0364642|T201|2501-5|LNC|UIBC SERPL-MCNC|UIBC SERPL-MCNC
C2739456|T201|56598-6|LNC|EBV EA IGM SER EIA-ACNC|EPSTEIN BARR VIRUS EARLY ANTIBODY.IMMUNOGLOBULIN M:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM:QUANTITATIVE:ENZYME IMMUNOASSAY
C0484851|T201|6598-7|LNC|TROPONIN T SERPL-MCNC|TROPONIN T.CARDIAC [MASS/VOLUME] IN SERUM OR PLASMA
C0364961|T201|6298-4|LNC|POTASSIUM BLD-SCNC|POTASSIUM [MOLES/VOLUME] IN BLOOD
C0482691|T201|6301-6|LNC|INR PPP|INR PPP
C0364489|T201|2349-9|LNC|GLUCOSE UR QL|GLUCOSE [PRESENCE] IN URINE
C0486210|T201|8247-9|LNC|MUCOUS THREADS URNS QL MICRO|MUCUS [PRESENCE] IN URINE SEDIMENT BY LIGHT MICROSCOPY
C0364856|T201|2713-6|LNC|SAO2% FROM PO2 BLD|SAO2 % BLD FROM PO2
C0362919|T201|798-9|LNC|RBC # UR AUTO|ERYTHROCYTES [#/VOLUME] IN URINE BY AUTOMATED COUNT
C0550529|T201|11579-0|LNC|TSH SERPL DL<=0.05 MIU/L-ACNC|THYROTROPIN:ARBITRARY CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE:DETECTION LIMIT <= 0.05 MIU/L
C0484485|T201|10331-7|LNC|RH BLD|RH BLD
C0364896|T201|2753-2|LNC|PH SERPL|PH OF SERUM OR PLASMA
C0365168|T201|3024-7|LNC|T4 FREE SERPL-MCNC|THYROXINE (T4) FREE [MASS/VOLUME] IN SERUM OR PLASMA
C0363126|T201|934-0|LNC|BPU ID|BPU ID
C0368061|T201|5811-5|LNC|SP GR UR STRIP|SP GR UR STRIP
C0364101|T201|35191-6|LNC|BILIRUB DIRECT SERPL-MCNC|BILIRUBIN.DIRECT [MASS OR MOLES/VOLUME] IN SERUM OR PLASMA
C0365111|T201|2965-2|LNC|SP GR UR|SP GR UR
C0364264|T201|2132-9|LNC|VIT B12 SERPL-MCNC|COBALAMINS:MCNC:PT:SER/PLAS:QN
C1146893|T201|31208-2|LNC|SPECIMEN SOURCE XXX|SPECIMEN SOURCE [IDENTIFIER] OF UNSPECIFIED SPECIMEN
C1978249|T201|50387-0|LNC|C TRACH RRNA CERVIX QL PCR|C TRACH RRNA CVX QL NAA+PROBE
C0365184|T201|3040-3|LNC|LIPASE SERPL-CCNC|LIPASE [ENZYMATIC ACTIVITY/VOLUME] IN SERUM OR PLASMA
C0803378|T201|20569-0|LNC|CK MB CFR SERPL|CK MB CFR SERPL
C0941357|T201|25162-9|LNC|HYALINE CASTS URNS QL MICRO|HYALINE CASTS [PRESENCE] IN URINE SEDIMENT BY LIGHT MICROSCOPY
C0797157|T201|13969-1|LNC|CK MB SERPL-MCNC|CREATINE KINASE.MB [MASS/VOLUME] IN SERUM OR PLASMA
C0368044|T201|5334-8|LNC|RUBV IGG SER EIA-ACNC|RUBV IGG SERPL IA-ACNC
C0942437|T201|26474-7|LNC|LYMPHOCYTES # BLD|LYMPHOCYTES [#/VOLUME] IN BLOOD
C0364227|T201|2091-7|LNC|VLDLC SERPL-MCNC|VLDLC SERPL-MCNC
C0368025|T201|5796-8|LNC|HYALINE CASTS #/AREA URNS LPF|HYALINE CASTS [#/AREA] IN URINE SEDIMENT BY MICROSCOPY LOW POWER FIELD
C0797133|T201|13945-1|LNC|RBC #/AREA URNS HPF|ERYTHROCYTES [#/AREA] IN URINE SEDIMENT BY MICROSCOPY HIGH POWER FIELD
C0362986|T201|769-0|LNC|NEUTS SEG NFR BLD MANUAL|SEGMENTED NEUTROPHILS/100 LEUKOCYTES IN BLOOD BY MANUAL COUNT
C0803224|T201|20409-9|LNC|RBC # UR STRIP|ERYTHROCYTES [#/VOLUME] IN URINE BY TEST STRIP
C0364295|T201|35204-7|LNC|CREAT UR-MCNC|CREATININE [MASS OR MOLES/VOLUME] IN URINE
C0484731|T201|2345-7|LNC|GLUCOSE SERPL-MCNC|GLUCOSE [MASS/VOLUME] IN SERUM OR PLASMA
C0803223|T201|20408-1|LNC|WBC # UR STRIP|LEUKOCYTES [#/VOLUME] IN URINE BY TEST STRIP
C0798370|T201|15199-3|LNC|MICROCYTES BLD QL AUTO|MICROCYTES [PRESENCE] IN BLOOD BY AUTOMATED COUNT
C2598074|T201|53927-0|LNC|N GONORRHOEA RRNA URTH QL PCR|NEISSERIA GONORRHOEAE RRNA [PRESENCE] IN URETHRA BY NAA WITH PROBE DETECTION
C1978250|T201|50388-8|LNC|N GONORRHOEA RRNA CERVIX QL PCR|N GONORRHOEA RRNA CVX QL NAA+PROBE
C0368040|T201|5802-4|LNC|NITRITE UR QL STRIP|NITRITE [PRESENCE] IN URINE BY TEST STRIP
C0362902|T201|713-8|LNC|EOSINOPHIL NFR BLD AUTO|EOSINOPHILS/100 LEUKOCYTES IN BLOOD BY AUTOMATED COUNT
C0364745|T201|2601-3|LNC|MAGNESIUM SERPL-SCNC|MAGNESIUM [MOLES/VOLUME] IN SERUM OR PLASMA
C0364108|T201|1975-2|LNC|BILIRUB SERPL-MCNC|BILIRUBIN.TOTAL [MASS/VOLUME] IN SERUM OR PLASMA
C0550264|T201|13457-7|LNC|LDLC SERPL CALC-MCNC|CHOLESTEROL IN LDL [MASS/VOLUME] IN SERUM OR PLASMA BY CALCULATION
C1116462|T201|30167-1|LNC|HPV I/H RISK 1 DNA CERVIX QL BDNA|HPV I/H RISK 1 DNA CVX QL PROBE+SIG AMP
C0363893|T201|1759-0|LNC|ALBUMIN/GLOB SERPL-MRTO|ALBUMIN/GLOBULIN [MASS RATIO] IN SERUM OR PLASMA
C0364479|T201|2339-0|LNC|GLUCOSE BLD-MCNC|GLUCOSE [MASS/VOLUME] IN BLOOD
C0803220|T201|20405-7|LNC|UROBILINOGEN UR STRIP-MCNC|UROBILINOGEN [MASS/VOLUME] IN URINE BY TEST STRIP
C0550795|T201|11253-2|LNC|TACROLIMUS BLD-MCNC|TACROLIMUS [MASS/VOLUME] IN BLOOD
C0802053|T201|19123-9|LNC|MAGNESIUM SERPL-MCNC|MAGNESIUM SERPL-MCNC
C0364055|T201|1920-8|LNC|AST SERPL-CCNC|ASPARTATE AMINOTRANSFERASE [ENZYMATIC ACTIVITY/VOLUME] IN SERUM OR PLASMA
C0367984|T201|5769-5|LNC|BACTERIA #/AREA URNS HPF|BACTERIA [#/AREA] IN URINE SEDIMENT BY MICROSCOPY HIGH POWER FIELD
C0362923|T201|718-7|LNC|HGB BLD-MCNC|HEMOGLOBIN [MASS/VOLUME] IN BLOOD
C0362906|T201|785-6|LNC|MCH RBC QN AUTO|MCH RBC QN AUTO
C1370010|T201|2777-1|LNC|PHOSPHATE SERPL-MCNC|PHOSPHATE [MASS/VOLUME] IN SERUM OR PLASMA
C0366106|T201|3879-4|LNC|OPIATES UR QL|OPIATES [PRESENCE] IN URINE
C0362909|T201|788-0|LNC|RDW RBC AUTO-RTO|ERYTHROCYTE DISTRIBUTION WIDTH [RATIO] BY AUTOMATED COUNT
C0362892|T201|704-7|LNC|BASOPHILS # BLD AUTO|BASOPHILS [#/VOLUME] IN BLOOD BY AUTOMATED COUNT
C0364294|T201|2160-0|LNC|CREAT SERPL-MCNC|CREAT SERPL-MCNC
C0800963|T201|17856-6|LNC|HGB A1C MFR BLD HPLC|HEMOGLOBIN A1C/HEMOGLOBIN.TOTAL IN BLOOD BY HPLC
C0368078|T201|5818-0|LNC|UROBILINOGEN UR QL STRIP|UROBILINOGEN [PRESENCE] IN URINE BY TEST STRIP
C0486204|T201|9842-6|LNC|CASTS #/AREA URNS LPF|CASTS [#/AREA] IN URINE SEDIMENT BY MICROSCOPY LOW POWER FIELD
C2360327|T201|51656-7|LNC|HCV AB S/CO FLD-RTO|HEPATITIS C VIRUS AB SIGNAL/CUTOFF IN BODY FLUID
C0365137|T201|2986-8|LNC|TESTOST SERPL-MCNC|TESTOST SERPL-MCNC
C0482602|T201|2842-3|LNC|PROLACTIN SERPL-MCNC|PROLACTIN [MASS/VOLUME] IN SERUM OR PLASMA
C0362951|T201|735-1|LNC|VARIANT LYMPHS NFR BLD MANUAL|LYMPHOCYTES.VARIANT/100 LEUKOCYTES:NUMBER FRACTION:POINT IN TIME:WHOLE BLOOD:QUANTITATIVE:MANUAL COUNT
C1147899|T201|32215-6|LNC|FTI SERPL-ACNC|THYROXINE (T4) FREE INDEX IN SERUM OR PLASMA BY CALCULATION
C0365620|T201|3390-2|LNC|BENZODIAZ UR QL|BENZODIAZEPINES [PRESENCE] IN URINE
C0364598|T201|2458-8|LNC|IGA SER-MCNC|IMMUNOGLOBULIN A:MASS CONCENTRATION:POINT IN TIME:SERUM/PLASMA:QUANTITATIVE
C0365583|T201|3349-8|LNC|AMPHETAMINES UR QL|AMPHETAMINES [PRESENCE] IN URINE
C0798132|T201|14959-1|LNC|MICROALBUMIN/CREAT UR-MRTO|MICROALBUMIN/CREATININE [MASS RATIO] IN URINE
C0551506|T201|11277-1|LNC|SQUAMOUS #/AREA URNS HPF|EPITHELIAL CELLS.SQUAMOUS [#/AREA] IN URINE SEDIMENT BY MICROSCOPY HIGH POWER FIELD
C0364111|T201|1978-6|LNC|BILIRUB UR-MCNC|BILIRUB UR-MCNC
C0798239|T201|15067-2|LNC|FSH SERPL-ACNC|FOLLITROPIN [UNITS/VOLUME] IN SERUM OR PLASMA
C0881037|T201|23658-8|LNC|OTHER ANTIBIOTIC SUSC ISLT|OTHER ANTIBIOTIC [SUSCEPTIBILITY]
