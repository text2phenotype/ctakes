ST|STREET
STR|STREET
RD|ROAD
PK|PIKE
AV|AVENUE
CRT|COURT
CT|COURT
CY|CANYON
CYN|CANYON
DR|DRIVE
LN|LANE
BLVD|BOULEVARD
CIR|CIRCLE
CR|CIRCLE
LP|LOOP
SQ|SQUARE
PL|PLACE
FWY|FREEWAY
FRWY|FREEWAY
PKWY|PARKWAY
TPK|TURNPIKE
HWY|HIGHWAY
BR|BRIDGE
TUNL|TUNNEL
TN|TUNNEL
MNT|MOUNTAIN
FY|FERRY
FRY|FERRY
JCT|JUNCTION