C0220847|T005|62944002|SNOMEDCT_US|HEPATITIS C VIRUS|HEPATITIS C VIRUS (ORGANISM)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS C|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0220847|T005|62944002|SNOMEDCT_US|HEPATITIS C VIRUS|HEPATITIS C VIRUS (ORGANISM)
C3839041|T005|702969000|SNOMEDCT_US|REACTIVATION OF HEPATITIS C VIRAL HEPATITIS|REACTIVATION OF HEPATITIS C VIRAL HEPATITIS (DISORDER)
C0369335|T005|121204002|SNOMEDCT_US|HEPATITIS C VIRUS RNA|HEPATITIS C VIRUS RNA (SUBSTANCE)
C0400914|T005|235866006|SNOMEDCT_US|ACUTE HEPATITIS C|ACUTE HEPATITIS C (DISORDER)
C0400920|T005|235872006|SNOMEDCT_US|HEPATITIS C CARRIER |HEPATITIS C CARRIER
C1112419|T005||SNOMEDCT_US|HEPATITIS C POSITIVE
C1698259|T005||SNOMEDCT_US|HCV COINFECTION
C0700073|T005|112386001|SNOMEDCT_US|VERY OLD NAME FOR HEP C|NON-A, NON-B HEPATITIS VIRUS (ORGANISM)
C0700073|T005|112386001|SNOMEDCT_US|ENTERICALLY-TRANSMITTED NON-A, NON-B HEPATITIS VIRUS ET-NANBHV|NON-A, NON-B HEPATITIS VIRUS (ORGANISM)
C0700073|T005|112386001|SNOMEDCT_US|NON-A NON-B HEPATITIS VIRUS|NON-A, NON-B HEPATITIS VIRUS (ORGANISM)
C0700073|T005|112386001|SNOMEDCT_US|NON-A, NON-B HEPATITIS VIRUS ET-NANBHV|NON-A, NON-B HEPATITIS VIRUS (ORGANISM)
C0700073|T005|112386001|SNOMEDCT_US|NON-A, NON-B HEPATITIS-ASSOCIATED VIRUS|NON-A, NON-B HEPATITIS VIRUS (ORGANISM)
C0700073|T005|112386001|SNOMEDCT_US|NON-A, NON-B HEPATITIS VIRUS|NON-A, NON-B HEPATITIS VIRUS (ORGANISM)
C0700073|T005|112386001|SNOMEDCT_US|NON-A, NON-B HEPATITIS VIRUS |NON-A, NON-B HEPATITIS VIRUS (ORGANISM)
C0079500|T005|243606007|SNOMEDCT_US|HEPACAVIRUS|GENUS HEPACIVIRUS
C0079500|T005|243606007|SNOMEDCT_US|HEPACIVIRUS|GENUS HEPACIVIRUS
C0079500|T005|243606007|SNOMEDCT_US|HEPACIVIRUSES|GENUS HEPACIVIRUS
C0079500|T005|243606007|SNOMEDCT_US|HEPATITIS C VIRUS GROUP|GENUS HEPACIVIRUS
C0079500|T005|243606007|SNOMEDCT_US|HEPATITIS C VIRUSES|GENUS HEPACIVIRUS
C0079500|T005|243606007|SNOMEDCT_US|HEPACAVIRUS |GENUS HEPACIVIRUS
C0079500|T005|243606007|SNOMEDCT_US|HEPACIVIRUS |GENUS HEPACIVIRUS
C3601684|T005||SNOMEDCT_US|UNCLASSIFIED HEPACIVIRUS
C0220847|T005|62944002|SNOMEDCT_US|HEPATITIS C VIRUS|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HEPATITIS C VIRUSES|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HEPATITIS C|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HEPATITIS C VIRUS (HCV)|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HCV|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HEPATITIS C VIRUS HCV|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HUMAN HEPATITIS C VIRUS|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HUMAN HEPATITIS C VIRUS HCV|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HUMAN HEPATITIS VIRUS C HCV|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|POST-TRANSFUSION HEPATITIS NON A NON B VIRUS|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HCV - HEPATITIS C VIRUS|HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|HEPATITIS C VIRUS |HEPATITIS C VIRUS (ORGANISM)
C0220847|T005|62944002|SNOMEDCT_US|VIRUS-HEPATITIS C|HEPATITIS C VIRUS (ORGANISM)
C3532919|T005|603422006|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 1 |HEPATITIS C VIRUS GENOTYPE 1 (ORGANISM)
C3532919|T005|603422006|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 1|HEPATITIS C VIRUS GENOTYPE 1 (ORGANISM)
C3532920|T005|603423001|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 2|HEPATITIS C VIRUS GENOTYPE 2 (ORGANISM)
C3532920|T005|603423001|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 2 |HEPATITIS C VIRUS GENOTYPE 2 (ORGANISM)
C3532921|T005|603424007|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 3 |HEPATITIS C VIRUS GENOTYPE 3 (ORGANISM)
C3532921|T005|603424007|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 3|HEPATITIS C VIRUS GENOTYPE 3 (ORGANISM)
C3532922|T005|603425008|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 4 |HEPATITIS C VIRUS GENOTYPE 4 (ORGANISM)
C3532922|T005|603425008|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 4|HEPATITIS C VIRUS GENOTYPE 4 (ORGANISM)
C3532923|T005|603426009|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 5 |HEPATITIS C VIRUS GENOTYPE 5 (ORGANISM)
C3532923|T005|603426009|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 5|HEPATITIS C VIRUS GENOTYPE 5 (ORGANISM)
C3532924|T005|603427000|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 6|HEPATITIS C VIRUS GENOTYPE 6 (ORGANISM)
C3532924|T005|603427000|SNOMEDCT_US|HEPATITIS C VIRUS GENOTYPE 6 |HEPATITIS C VIRUS GENOTYPE 6 (ORGANISM)
C3494961|T005|603418001|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 3B |HEPATITIS C VIRUS SUBTYPE 3B (ORGANISM)
C3494961|T005|603418001|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 3B|HEPATITIS C VIRUS SUBTYPE 3B (ORGANISM)
C3494962|T005|603417006|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 3A|HEPATITIS C VIRUS SUBTYPE 3A (ORGANISM)
C3494962|T005|603417006|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 3A |HEPATITIS C VIRUS SUBTYPE 3A (ORGANISM)
C3494958|T005|603420003|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 6A |HEPATITIS C VIRUS SUBTYPE 6A (ORGANISM)
C3494958|T005|603420003|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 6A|HEPATITIS C VIRUS SUBTYPE 6A (ORGANISM)
C3494966|T005|603413005|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 1A |HEPATITIS C VIRUS SUBTYPE 1A (ORGANISM)
C3494966|T005|603413005|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 1A|HEPATITIS C VIRUS SUBTYPE 1A (ORGANISM)
C3494964|T005|603415003|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 2A|HEPATITIS C VIRUS SUBTYPE 2A (ORGANISM)
C3494964|T005|603415003|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 2A |HEPATITIS C VIRUS SUBTYPE 2A (ORGANISM)
C3494959|T005|603419009|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 5A |HEPATITIS C VIRUS SUBTYPE 5A (ORGANISM)
C3494959|T005|603419009|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 5A|HEPATITIS C VIRUS SUBTYPE 5A (ORGANISM)
C3494963|T005|603416002|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 2B |HEPATITIS C VIRUS SUBTYPE 2B (ORGANISM)
C3494963|T005|603416002|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 2B|HEPATITIS C VIRUS SUBTYPE 2B (ORGANISM)
C3494965|T005|603414004|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 1B |HEPATITIS C VIRUS SUBTYPE 1B (ORGANISM)
C3494965|T005|603414004|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 1B|HEPATITIS C VIRUS SUBTYPE 1B (ORGANISM)
C3662864|T005|431831000124103|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 4|HEPATITIS C VIRUS SUBTYPE 4 (ORGANISM)
C3662864|T005|431831000124103|SNOMEDCT_US|HEPATITIS C VIRUS SUBTYPE 4 |HEPATITIS C VIRUS SUBTYPE 4 (ORGANISM)
C0524910|T005|186640001|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS C|CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|HEPATITIS C, CHRONIC|CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|CHRONIC HEPATITIS, C VIRUS|CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS C INFECTION|CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|CHRONIC HEPATITIS C INFECTION |CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|CHRONIC HEPATITIS C INFECTION|CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|CHRONIC HEPATITIS C|CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|HEPATITIS C, CHRONIC [DISEASE/FINDING]|CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS C |CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|CHRONIC HEPATITIS C |CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|CHRONIC TYPE C VIRAL HEPATITIS|CHRONIC VIRAL HEPATITIS C (DISORDER)
C0524910|T005|186640001|SNOMEDCT_US|HEPATITIS; VIRUS, CHRONIC, TYPE C|CHRONIC VIRAL HEPATITIS C (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS C|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|PT NANBH|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRAL HEPATITIS, NON-A, NON-B -RETIRED-|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRAL HEPATITIS C INFECTION|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS C INFECTION |VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS C INFECTION|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS NON-A NON-B|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|UNSPECIFIED VIRAL HEPATITIS C|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRAL HEPATITIS C NOS|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS C [DISEASE/FINDING]|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|PT-NANBH|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|PARENTERALLY-TRANSMITTED NON-A, NON-B HEPATITIS|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS, VIRAL, NON-A, NON-B, PARENTERALLY-TRANSMITTED|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|PARENTERALLY TRANSMITTED NON A, NON B HEPATITIS|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRAL HEPATITIS, NON-A, NON-B|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS C |VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRAL HEPATITIS, NON-A, NON-B |VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRAL HEPATITIS C |VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRAL HEPATITIS TYPE C |VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRAL HEPATITIS TYPE C|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|NON-A NON-B HEPATITIS|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEP NON-A NON-B|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRAL HEPATITIS C|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS (NON-A NON-B)|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|TYPE C VIRAL HEPATITIS|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS NON-A NON-B |VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS NONA NONB|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS NON A NON B|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS; VIRUS, NON-A, NON-B|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|HEPATITIS; VIRUS, TYPE C|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|NON-A NON-B-HEPATITIS|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|VIRUS; HEPATITIS, NON-A, NON-B|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|NON-A, NON-B HEPATITIS|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|NANBH|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C0019196|T005|123324009|SNOMEDCT_US|UNSPECIFIED VIRAL HEPATITIS C NOS|VIRAL HEPATITIS, NON-A, NON-B (DISORDER)
C2711110|T005|442374005|SNOMEDCT_US|HEPATITIS B AND HEPATITIS C |HEPATITIS B AND HEPATITIS C (DISORDER)
C2711110|T005|442374005|SNOMEDCT_US|HEPATITIS B AND HEPATITIS C|HEPATITIS B AND HEPATITIS C (DISORDER)
C2711110|T005|442374005|SNOMEDCT_US|HEPATITIS B AND HEPATITIS C |HEPATITIS B AND HEPATITIS C (DISORDER)
C2711110|T005|442374005|SNOMEDCT_US|HEPATITIS VIRAL B AND C|HEPATITIS B AND HEPATITIS C (DISORDER)
C1456263|T005||SNOMEDCT_US|HPT C W/O HEPAT COMA NOS
C1456263|T005||SNOMEDCT_US|UNSPECIFIED VIRAL HEPATITIS C WITHOUT HEPATIC COMA
C1456265|T005||SNOMEDCT_US|HPT C W HEPATIC COMA NOS
C1456265|T005||SNOMEDCT_US|UNSPECIFIED VIRAL HEPATITIS C WITH HEPATIC COMA
C2063424|T005||SNOMEDCT_US|CHRONIC HEPATITIS C INFECTION WITH HEPATIC COMA 
C2063424|T005||SNOMEDCT_US|HEPATITIS, C VIRUS WITH HEPATIC COMA
C2063424|T005||SNOMEDCT_US|CHRONIC VIRAL HEPATITIS C INFECTION WITH HEPATIC COMA
C2063424|T005||SNOMEDCT_US|CHRONIC HEPATITIS, C VIRUS WITH HEPATIC COMA
C2063424|T005||SNOMEDCT_US|HEPATITIS C INFECTION WITH HEPATIC COMA 
C2063424|T005||SNOMEDCT_US|HEPATITIS C INFECTION WITH HEPATIC COMA
C2063424|T005||SNOMEDCT_US|CHRONIC HEPATITIS C INFECTION WITH HEPATIC COMA
C0400914|T005|235866006|SNOMEDCT_US|ACUTE HEPATITIS C|ACUTE HEPATITIS C (DISORDER)
C0400914|T005|235866006|SNOMEDCT_US|ACUTE VIRAL HEPATITIS C INFECTION|ACUTE HEPATITIS C (DISORDER)
C0400914|T005|235866006|SNOMEDCT_US|ACUTE HEPATITIS C INFECTION |ACUTE HEPATITIS C (DISORDER)
C0400914|T005|235866006|SNOMEDCT_US|ACUTE HEPATITIS C INFECTION|ACUTE HEPATITIS C (DISORDER)
C0400914|T005|235866006|SNOMEDCT_US|ACUTE TYPE C VIRAL HEPATITIS|ACUTE HEPATITIS C (DISORDER)
C0400914|T005|235866006|SNOMEDCT_US|ACUTE HEPATITIS C NOS|ACUTE HEPATITIS C (DISORDER)
C0400914|T005|235866006|SNOMEDCT_US|HEPATITIS C, ACUTE|ACUTE HEPATITIS C (DISORDER)
C0400914|T005|235866006|SNOMEDCT_US|ACUTE HEPATITIS C |ACUTE HEPATITIS C (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|POSTTRANSFUSION HEPATITIS|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|HEPATITIS POST TRANSFUSION|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|POST TRANSFUSION HEPATITIS|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|POSTTRANSFUSION VIRAL HEPATITIS |POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|POSTTRANSFUSION VIRAL HEPATITIS|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|TRANSFUSION HEPATITIS|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|HEPATITIS; POST-TRANSFUSION|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|POST-TRANSFUSION; HEPATITIS|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|POSTTRANSFUSION HEPATITIS, NOS|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|POSTTRANSFUSION VIRAL HEPATITIS, NOS|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0520788|T005|28766006|SNOMEDCT_US|TRANSFUSION HEPATITIS, NOS|POSTTRANSFUSION VIRAL HEPATITIS (DISORDER)
C0400900|T005|186631000|SNOMEDCT_US|VIRAL HEPATITIS C WITHOUT MENTION OF HEPATIC COMA |VIRAL HEPATITIS C WITHOUT MENTION OF HEPATIC COMA (DISORDER)
C0400900|T005|186631000|SNOMEDCT_US|VIRAL HEPATITIS C WITHOUT MENTION OF HEPATIC COMA|VIRAL HEPATITIS C WITHOUT MENTION OF HEPATIC COMA (DISORDER)
C0375009|T005|435101000124104|SNOMEDCT_US|CHRNC HPT C W HEPAT COMA|CHRONIC VIRAL HEPATITIS C WITH HEPATIC COMA (DISORDER)
C0375009|T005|435101000124104|SNOMEDCT_US|CHRONIC HEPATITIS C WITH HEPATIC COMA|CHRONIC VIRAL HEPATITIS C WITH HEPATIC COMA (DISORDER)
C0375009|T005|435101000124104|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS C WITH HEPATIC COMA |CHRONIC VIRAL HEPATITIS C WITH HEPATIC COMA (DISORDER)
C0375009|T005|435101000124104|SNOMEDCT_US|CHRONIC VIRAL HEPATITIS C WITH HEPATIC COMA|CHRONIC VIRAL HEPATITIS C WITH HEPATIC COMA (DISORDER)
C3837244|T005||SNOMEDCT_US|HEPATITIS, C VIRUS - WITHOUT HEPATIC COMA
C3837244|T005||SNOMEDCT_US|HEPATITIS, C VIRUS WITHOUT HEPATIC COMA
C3837244|T005||SNOMEDCT_US|HEPATITIS, C VIRUS WITHOUT HEPATIC COMA 
C3839041|T005|702969000|SNOMEDCT_US|REACTIVATION OF HEPATITIS C VIRAL HEPATITIS |REACTIVATION OF HEPATITIS C VIRAL HEPATITIS (DISORDER)
C3839041|T005|702969000|SNOMEDCT_US|REACTIVATION OF HEPATITIS C VIRAL HEPATITIS|REACTIVATION OF HEPATITIS C VIRAL HEPATITIS (DISORDER)
C0400915|T005|186628001|SNOMEDCT_US|VIRAL HEPATITIS C WITH COMA|VIRAL HEPATITIS C WITH COMA (DISORDER)
C0400915|T005|186628001|SNOMEDCT_US|VIRAL HEPATITIS C WITH COMA |VIRAL HEPATITIS C WITH COMA (DISORDER)
C0241911|T005|235870003|SNOMEDCT_US|CHRONIC NON-A NON-B HEPATITIS|CHRONIC NON-A NON-B HEPATITIS (DISORDER)
C0241911|T005|235870003|SNOMEDCT_US|CHRONIC NON-A NON-B HEPATITIS |CHRONIC NON-A NON-B HEPATITIS (DISORDER)
C0458009|T005|278929008|SNOMEDCT_US|CONGENITAL HEPATITIS C INFECTION|CONGENITAL HEPATITIS C INFECTION (DISORDER)
C0458009|T005|278929008|SNOMEDCT_US|CONGENITAL HEPATITIS C INFECTION |CONGENITAL HEPATITIS C INFECTION (DISORDER)
C2357728|T005||SNOMEDCT_US|HEPATITIS C VIRUS RNA &#X7C; BODY FLUID
C1989118|T005||SNOMEDCT_US|HEPATITIS C VIRUS RNA &#X7C; BLD-SER-PLAS
C1989120|T005||SNOMEDCT_US|HEPATITIS C VIRUS RNA &#X7C; CEREBRAL SPINAL FLUID
C1989119|T005||SNOMEDCT_US|HEPATITIS C VIRUS RNA &#X7C; BONE MARROW
C1989121|T005||SNOMEDCT_US|HEPATITIS C VIRUS RNA &#X7C; TISSUE AND SMEARS
C1989122|T005||SNOMEDCT_US|HEPATITIS C VIRUS RNA &#X7C; XXX
C1545335|T005||SNOMEDCT_US|HIV 1+HEPATITIS C VIRUS RNA
C1545335|T005||SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS 1+HEPATITIS C VIRUS RIBONUCLEIC ACID
C2911593|T005||SNOMEDCT_US|ACUTE HEPATITIS C WITHOUT HEPATIC COMA
C1456261|T005||SNOMEDCT_US|HPT C ACUTE W HEPAT COMA
C1456261|T005||SNOMEDCT_US|ACUTE HEPATITIS C WITH HEPATIC COMA
C2215293|T005||SNOMEDCT_US|ACUTE HEPATITIS C INFECTION WITH HEPATIC COMA
C2215293|T005||SNOMEDCT_US|ACUTE HEPATITIS C INFECTION WITH HEPATIC COMA 
C2215293|T005||SNOMEDCT_US|ACUTE TYPE C VIRAL HEPATITIS WITH HEPATIC COMA
C2118423|T005||SNOMEDCT_US|ACUTE HEPATITIS C INFECTION WITH FULMINANT HEPATIC FAILURE
C2118423|T005||SNOMEDCT_US|ACUTE HEPATITIS C INFECTION WITH FULMINANT HEPATIC FAILURE 
C2118423|T005||SNOMEDCT_US|ACUTE TYPE C VIRAL HEPATITIS WITH FULMINANT HEPATIC FAILURE
C3838646|T005||SNOMEDCT_US|ACUTE HEPATITIS, C VIRUS WITHOUT HEPATIC COMA
C3838646|T005||SNOMEDCT_US|ACUTE HEPATITIS, C VIRUS WITHOUT HEPATIC COMA 
C3838646|T005||SNOMEDCT_US|HEPATITIS, C VIRUS - ACUTE WITHOUT HEPATIC COMA
C0400920|T005|235872006|SNOMEDCT_US|HEPATITIS C CARRIER |HEPATITIS C CARRIER
C0400920|T005|235872006|SNOMEDCT_US|HEPATITIS C CARRIER|HEPATITIS C CARRIER
C2025298|T005||SNOMEDCT_US|CARRYING VIRAL HEPATITIS TYPE C
C2025298|T005||SNOMEDCT_US|CARRIER OF TYPE C VIRAL HEPATITIS
C2025298|T005||SNOMEDCT_US|CARRIER OF TYPE C VIRAL HEPATITIS 
C1112419|T005||SNOMEDCT_US|HEPATITIS C POSITIVE
C1698259|T005||SNOMEDCT_US|HCV COINFECTION
