C0362625|T201|COMP|6019-4|LNC2000|Prunus dulcis Ab.IgE|Prunus dulcis Ab.IgE
C0362627|T201|COMP|6021-0|LNC2000|Malus sylvestris Ab.IgE|Malus sylvestris Ab.IgE
C0362631|T201|COMP|6025-1|LNC2000|Aspergillus fumigatus Ab.IgE|Aspergillus fumigatus Ab.IgE
C0362634|T201|COMP|6029-3|LNC2000|Aureobasidium pullulans Ab.IgE|Aureobasidium pullulans Ab.IgE
C0362640|T201|COMP|6034-3|LNC2000|Paspalum notatum Ab.IgE|Paspalum notatum Ab.IgE
C0362641|T201|COMP|6035-0|LNC2000|Musa spp Ab.IgE|Musa spp Ab.IgE
C0362642|T201|COMP|6037-6|LNC2000|Hordeum vulgare Ab.IgE|Hordeum vulgare Ab.IgE
C0362644|T201|COMP|6038-4|LNC2000|Fagus grandifolia Ab.IgE|Fagus grandifolia Ab.IgE
C0362645|T201|COMP|6039-2|LNC2000|Beef Ab.IgE|Beef Ab.IgE
C0362647|T201|COMP|6041-8|LNC2000|Cynodon dactylon Ab.IgE|Cynodon dactylon Ab.IgE
C0362656|T201|COMP|6050-9|LNC2000|Bertholletia excelsa Ab.IgE|Bertholletia excelsa Ab.IgE
C0362665|T201|COMP|6059-0|LNC2000|Candida albicans Ab.IgE|Candida albicans Ab.IgE
C0362667|T201|COMP|6061-6|LNC2000|Daucus carota Ab.IgE|Daucus carota Ab.IgE
C0362668|T201|COMP|6062-4|LNC2000|Casein Ab.IgE|Casein Ab.IgE
C0362679|T201|COMP|6073-1|LNC2000|Chocolate Ab.IgE|Chocolate Ab.IgE
C0362681|T201|COMP|6075-6|LNC2000|Cladosporium herbarum Ab.IgE|Cladosporium herbarum Ab.IgE
C0362682|T201|COMP|6076-4|LNC2000|Ruditapes spp Ab.IgE|Ruditapes spp Ab.IgE
C0362684|T201|COMP|6078-0|LNC2000|Blatella germanica Ab.IgE|Blatella germanica Ab.IgE
C0362686|T201|COMP|6081-4|LNC2000|Cocos nucifera Ab.IgE|Cocos nucifera Ab.IgE
C0362687|T201|COMP|6082-2|LNC2000|Gadus morhua Ab.IgE|Gadus morhua Ab.IgE
C0362690|T201|COMP|6085-5|LNC2000|Ambrosia elatior Ab.IgE|Ambrosia elatior Ab.IgE
C0362691|T201|COMP|6087-1|LNC2000|Zea mays Ab.IgE|Zea mays Ab.IgE
C0362694|T201|COMP|6090-5|LNC2000|Populus deltoides Ab.IgE|Populus deltoides Ab.IgE
C0362696|T201|COMP|6092-1|LNC2000|Cancer pagurus Ab.IgE|Cancer pagurus Ab.IgE
C0362699|T201|COMP|6095-4|LNC2000|Dermatophagoides farinae Ab.IgE|Dermatophagoides farinae Ab.IgE
C0362700|T201|COMP|6096-2|LNC2000|Dermatophagoides pteronyssinus Ab.IgE|Dermatophagoides pteronyssinus Ab.IgE
C0362701|T201|COMP|6098-8|LNC2000|Dog dander Ab.IgE|Dog dander Ab.IgE
C0362702|T201|COMP|6099-6|LNC2000|Dog epithelium Ab.IgE|Dog epithelium Ab.IgE
C0362708|T201|COMP|6106-9|LNC2000|Egg white Ab.IgE|Egg white Ab.IgE
C0362709|T201|COMP|6107-7|LNC2000|Egg yolk Ab.IgE|Egg yolk Ab.IgE
C0362712|T201|COMP|6110-1|LNC2000|Plantago lanceolata Ab.IgE|Plantago lanceolata Ab.IgE
C0362715|T201|COMP|6113-5|LNC2000|Eucalyptus spp Ab.IgE|Eucalyptus spp Ab.IgE
C0362727|T201|COMP|6125-9|LNC2000|Gluten Ab.IgE|Gluten Ab.IgE
C0362738|T201|COMP|6136-6|LNC2000|Corylus avellana Ab.IgE|Corylus avellana Ab.IgE
C0362739|T201|COMP|6137-4|LNC2000|Corylus avellana pollen Ab.IgE|Corylus avellana pollen Ab.IgE
C0362740|T201|COMP|6138-2|LNC2000|Setomelanomma rostrata Ab.IgE|Setomelanomma rostrata Ab.IgE
C0362752|T201|COMP|6151-5|LNC2000|Cupressus sempervirens Ab.IgE|Cupressus sempervirens Ab.IgE
C0362753|T201|COMP|6152-3|LNC2000|Sorghum halepense Ab.IgE|Sorghum halepense Ab.IgE
C0362754|T201|COMP|6153-1|LNC2000|Poa pratensis Ab.IgE|Poa pratensis Ab.IgE
C0362758|T201|COMP|6156-4|LNC2000|Chenopodium album Ab.IgE|Chenopodium album Ab.IgE
C0362759|T201|COMP|6158-0|LNC2000|Latex Ab.IgE|Latex Ab.IgE
C0362766|T201|COMP|6165-5|LNC2000|Homarus gammarus Ab.IgE|Homarus gammarus Ab.IgE
C0362775|T201|COMP|6174-7|LNC2000|Milk Ab.IgE|Milk Ab.IgE
C0362779|T201|COMP|6178-8|LNC2000|Juniperus sabinoides Ab.IgE|Juniperus sabinoides Ab.IgE
C0362783|T201|COMP|6182-0|LNC2000|Mucor racemosus Ab.IgE|Mucor racemosus Ab.IgE
C0362784|T201|COMP|6183-8|LNC2000|Artemisia vulgaris Ab.IgE|Artemisia vulgaris Ab.IgE
C0362787|T201|COMP|6186-1|LNC2000|Urtica dioica Ab.IgE|Urtica dioica Ab.IgE
C0362795|T201|COMP|6194-5|LNC2000|Citrus sinensis Ab.IgE|Citrus sinensis Ab.IgE
C0362796|T201|COMP|6195-2|LNC2000|Dactylis glomerata Ab.IgE|Dactylis glomerata Ab.IgE
C0362807|T201|COMP|6206-7|LNC2000|Arachis hypogaea Ab.IgE|Arachis hypogaea Ab.IgE
C0362813|T201|COMP|6212-5|LNC2000|Penicillium notatum Ab.IgE|Penicillium notatum Ab.IgE
C0362820|T201|COMP|6219-0|LNC2000|Pork Ab.IgE|Pork Ab.IgE
C0362823|T201|COMP|6222-4|LNC2000|Syagrus romanzoffianum Ab.IgE|Syagrus romanzoffianum Ab.IgE
C0362831|T201|COMP|6230-7|LNC2000|Oryza sativa Ab.IgE|Oryza sativa Ab.IgE
C0362834|T201|COMP|6233-1|LNC2000|Pigweed rough Ab.IgE|Pigweed rough Ab.IgE
C0362835|T201|COMP|6234-9|LNC2000|Salsola kali Ab.IgE|Salsola kali Ab.IgE
C0362838|T201|COMP|6237-2|LNC2000|Salmo salar Ab.IgE|Salmo salar Ab.IgE
C0362843|T201|COMP|6242-2|LNC2000|Sesamum indicum Ab.IgE|Sesamum indicum Ab.IgE
C0362845|T201|COMP|6244-8|LNC2000|Rumex acetosella Ab.IgE|Rumex acetosella Ab.IgE
C0362847|T201|COMP|6246-3|LNC2000|Pandalus borealis Ab.IgE|Pandalus borealis Ab.IgE
C0362853|T201|COMP|6252-1|LNC2000|Stemphylium botryosum Ab.IgE|Stemphylium botryosum Ab.IgE
C0362858|T201|COMP|6257-0|LNC2000|Fragaria vesca Ab.IgE|Fragaria vesca Ab.IgE
C0362866|T201|COMP|6265-3|LNC2000|Phleum pratense Ab.IgE|Phleum pratense Ab.IgE
C0362867|T201|COMP|6266-1|LNC2000|Lycopersicon lycopersicum Ab.IgE|Lycopersicon lycopersicum Ab.IgE
C0362871|T201|COMP|6270-3|LNC2000|Thunnus albacares Ab.IgE|Thunnus albacares Ab.IgE
C0362874|T201|COMP|6273-7|LNC2000|Juglans spp Ab.IgE|Juglans spp Ab.IgE
C0362877|T201|COMP|6276-0|LNC2000|Triticum aestivum Ab.IgE|Triticum aestivum Ab.IgE
C0362879|T201|COMP|6278-6|LNC2000|Fraxinus americana Ab.IgE|Fraxinus americana Ab.IgE
C0362887|T201|COMP|6286-9|LNC2000|Artemisia absinthium Ab.IgE|Artemisia absinthium Ab.IgE
C0362888|T201|COMP|6287-7|LNC2000|Saccharomyces cerevisiae Ab.IgE|Saccharomyces cerevisiae Ab.IgE
C0362890|T201|COMP|702-1|LNC2000|Anisocytosis|Anisocytosis
C0362891|T201|COMP|703-9|LNC2000|Basophilic stippling|Basophilic stippling
C0362892|T201|COMP|704-7|LNC2000|Basophils|Basophils
C0362894|T201|COMP|706-2|LNC2000|Basophils/100 leukocytes|Basophils/100 leukocytes
C0362895|T201|COMP|707-0|LNC2000|Basophils/100 leukocytes|Basophils/100 leukocytes
C0362896|T201|COMP|708-8|LNC2000|Blasts|Blasts
C0362897|T201|COMP|709-6|LNC2000|Blasts/100 leukocytes|Blasts/100 leukocytes
C0362898|T201|COMP|5909-7|LNC2000|Blood smear finding|Blood smear finding
C0362900|T201|COMP|711-2|LNC2000|Eosinophils|Eosinophils
C0362902|T201|COMP|713-8|LNC2000|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0362903|T201|COMP|714-6|LNC2000|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0362906|T201|COMP|785-6|LNC2000|Erythrocyte mean corpuscular hemoglobin|Erythrocyte mean corpuscular hemoglobin
C0362908|T201|COMP|787-2|LNC2000|Erythrocyte mean corpuscular volume|Erythrocyte mean corpuscular volume
C0362909|T201|COMP|788-0|LNC2000|Erythrocyte distribution width|Erythrocyte distribution width
C0362910|T201|COMP|789-8|LNC2000|Erythrocytes|Erythrocytes
C0362913|T201|COMP|792-2|LNC2000|Erythrocytes|Erythrocytes
C0362919|T201|COMP|798-9|LNC2000|Erythrocytes|Erythrocytes
C0362921|T201|COMP|716-1|LNC2000|Heinz bodies|Heinz bodies
C0362923|T201|COMP|718-7|LNC2000|Hemoglobin|Hemoglobin
C0362926|T201|COMP|721-1|LNC2000|Hemoglobin.free|Hemoglobin.free
C0362933|T201|COMP|728-6|LNC2000|Hypochromia|Hypochromia
C0362936|T201|COMP|806-0|LNC2000|Leukocytes|Leukocytes
C0362938|T201|COMP|808-6|LNC2000|Leukocytes|Leukocytes
C0362946|T201|COMP|730-2|LNC2000|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0362947|T201|COMP|731-0|LNC2000|Lymphocytes|Lymphocytes
C0362951|T201|COMP|735-1|LNC2000|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C0362952|T201|COMP|736-9|LNC2000|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0362953|T201|COMP|737-7|LNC2000|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0362954|T201|COMP|738-5|LNC2000|Macrocytes|Macrocytes
C0362955|T201|COMP|739-3|LNC2000|Metamyelocytes|Metamyelocytes
C0362956|T201|COMP|740-1|LNC2000|Metamyelocytes/100 leukocytes|Metamyelocytes/100 leukocytes
C0362957|T201|COMP|741-9|LNC2000|Microcytes|Microcytes
C0362958|T201|COMP|742-7|LNC2000|Monocytes|Monocytes
C0362959|T201|COMP|743-5|LNC2000|Monocytes|Monocytes
C0362960|T201|COMP|5905-5|LNC2000|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0362961|T201|COMP|744-3|LNC2000|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0362965|T201|COMP|748-4|LNC2000|Myelocytes|Myelocytes
C0362967|T201|COMP|749-2|LNC2000|Myelocytes/100 leukocytes|Myelocytes/100 leukocytes
C0362968|T201|COMP|751-8|LNC2000|Neutrophils|Neutrophils
C0362980|T201|COMP|763-3|LNC2000|Neutrophils.band form|Neutrophils.band form
C0362981|T201|COMP|764-1|LNC2000|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0362982|T201|COMP|765-8|LNC2000|Neutrophils.hypersegmented|Neutrophils.hypersegmented
C0362986|T201|COMP|769-0|LNC2000|Neutrophils.segmented/100 leukocytes|Neutrophils.segmented/100 leukocytes
C0362987|T201|COMP|770-8|LNC2000|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0362988|T201|COMP|771-6|LNC2000|Erythrocytes.nucleated|Erythrocytes.nucleated
C0362989|T201|COMP|772-4|LNC2000|Erythrocytes.nucleated|Erythrocytes.nucleated
C0362990|T201|COMP|773-2|LNC2000|Erythrocytes.nucleated/100 erythrocytes|Erythrocytes.nucleated/100 erythrocytes
C0362991|T201|COMP|774-0|LNC2000|Ovalocytes|Ovalocytes
C0362994|T201|COMP|777-3|LNC2000|Platelets|Platelets
C0362996|T201|COMP|5908-9|LNC2000|Platelets.giant|Platelets.giant
C0362997|T201|COMP|7791-7|LNC2000|Dacryocytes|Dacryocytes
C0362999|T201|COMP|781-5|LNC2000|Promyelocytes|Promyelocytes
C0363002|T201|COMP|800-3|LNC2000|Schistocytes|Schistocytes
C0363003|T201|COMP|801-1|LNC2000|Sickle cells|Sickle cells
C0363004|T201|COMP|802-9|LNC2000|Spherocytes|Spherocytes
C0363005|T201|COMP|803-7|LNC2000|Toxic granules|Toxic granules
C0363081|T201|COMP|890-4|LNC2000|Blood group antibody screen|Blood group antibody screen
C0363117|T201|COMP|925-8|LNC2000|Blood product disposition|Blood product disposition
C0363123|T201|COMP|931-6|LNC2000|Blood product source|Blood product source
C0363126|T201|COMP|934-0|LNC2000|Blood product unit ID|Blood product unit ID
C0363128|T201|COMP|936-5|LNC2000|Blood product unit identifier|Blood product unit identifier
C0363184|T201|COMP|1305-2|LNC2000|D Ag|D Ag
C0363413|T201|COMP|1250-0|LNC2000|Major crossmatch|Major crossmatch
C0363635|T201|COMP|1501-6|LNC2000|Glucose^1H post 100 g glucose PO|Glucose^1H post 100 g glucose PO
C0363638|T201|COMP|1504-0|LNC2000|Glucose^1H post 50 g glucose PO|Glucose^1H post 50 g glucose PO
C0363641|T201|COMP|1507-3|LNC2000|Glucose^1H post 75 g glucose PO|Glucose^1H post 75 g glucose PO
C0363647|T201|COMP|1514-9|LNC2000|Glucose^2H post 100 g glucose PO|Glucose^2H post 100 g glucose PO
C0363651|T201|COMP|1518-0|LNC2000|Glucose^2H post 75 g glucose PO|Glucose^2H post 75 g glucose PO
C0363662|T201|COMP|1530-5|LNC2000|Glucose^3H post 100 g glucose PO|Glucose^3H post 100 g glucose PO
C0363783|T201|COMP|1649-3|LNC2000|Calcitriol|Calcitriol
C0363802|T201|COMP|1668-3|LNC2000|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C0363829|T201|COMP|1695-6|LNC2000|5-Hydroxyindoleacetate|5-Hydroxyindoleacetate
C0363876|T201|COMP|1742-6|LNC2000|Alanine aminotransferase|Alanine aminotransferase
C0363880|T201|COMP|1746-7|LNC2000|Albumin|Albumin
C0363881|T201|COMP|1747-5|LNC2000|Albumin|Albumin
C0363885|T201|COMP|1751-7|LNC2000|Albumin|Albumin
C0363893|T201|COMP|1759-0|LNC2000|Albumin/Globulin|Albumin/Globulin
C0363895|T201|COMP|1761-6|LNC2000|Aldolase|Aldolase
C0363897|T201|COMP|1763-2|LNC2000|Aldosterone|Aldosterone
C0363911|T201|COMP|1777-2|LNC2000|Alkaline phosphatase.bone|Alkaline phosphatase.bone
C0363913|T201|COMP|1779-8|LNC2000|Alkaline phosphatase.liver|Alkaline phosphatase.liver
C0363929|T201|COMP|1795-4|LNC2000|Amylase|Amylase
C0363968|T201|COMP|1834-1|LNC2000|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0363983|T201|COMP|1848-1|LNC2000|Androstanolone|Androstanolone
C0363989|T201|COMP|1854-9|LNC2000|Androstenedione|Androstenedione
C0363992|T201|COMP|1857-2|LNC2000|Angiotensin converting enzyme|Angiotensin converting enzyme
C0363998|T201|COMP|1863-0|LNC2000|Anion gap 4|Anion gap 4
C0364006|T201|COMP|1871-3|LNC2000|Apolipoprotein B-100|Apolipoprotein B-100
C0364019|T201|COMP|1884-6|LNC2000|Apolipoprotein B|Apolipoprotein B
C0364055|T201|COMP|1920-8|LNC2000|Aspartate aminotransferase|Aspartate aminotransferase
C0364057|T201|COMP|1922-4|LNC2000|Base deficit|Base deficit
C0364059|T201|COMP|1924-0|LNC2000|Base deficit|Base deficit
C0364060|T201|COMP|1925-7|LNC2000|Base excess|Base excess
C0364061|T201|COMP|1926-5|LNC2000|Base excess|Base excess
C0364062|T201|COMP|1927-3|LNC2000|Base excess|Base excess
C0364085|T201|COMP|1952-1|LNC2000|Beta-2-Microglobulin|Beta-2-Microglobulin
C0364092|T201|COMP|1959-6|LNC2000|Bicarbonate|Bicarbonate
C0364093|T201|COMP|1960-4|LNC2000|Bicarbonate|Bicarbonate
C0364094|T201|COMP|1961-2|LNC2000|Bicarbonate|Bicarbonate
C0364101|T201|COMP|1968-7|LNC2000|Bilirubin.glucuronidated+Bilirubin.albumin bound|Bilirubin.glucuronidated+Bilirubin.albumin bound
C0364104|T201|COMP|1971-1|LNC2000|Bilirubin.non-glucuronidated|Bilirubin.non-glucuronidated
C0364108|T201|COMP|1975-2|LNC2000|Bilirubin|Bilirubin
C0364110|T201|COMP|1977-8|LNC2000|Bilirubin|Bilirubin
C0364111|T201|COMP|1978-6|LNC2000|Bilirubin|Bilirubin
C0364119|T201|COMP|1986-9|LNC2000|C peptide|C peptide
C0364121|T201|COMP|1988-5|LNC2000|C reactive protein|C reactive protein
C0364122|T201|COMP|1989-3|LNC2000|Calcidiol|Calcidiol
C0364123|T201|COMP|1990-1|LNC2000|Cholecalciferol|Cholecalciferol
C0364125|T201|COMP|1992-7|LNC2000|Calcitonin|Calcitonin
C0364127|T201|COMP|1994-3|LNC2000|Calcium.ionized|Calcium.ionized
C0364128|T201|COMP|1995-0|LNC2000|Calcium.ionized|Calcium.ionized
C0364139|T201|COMP|2006-5|LNC2000|Cancer Ag 125|Cancer Ag 125
C0364151|T201|COMP|2019-8|LNC2000|Carbon dioxide|Carbon dioxide
C0364153|T201|COMP|2021-4|LNC2000|Carbon dioxide|Carbon dioxide
C0364158|T201|COMP|2026-3|LNC2000|Carbon dioxide|Carbon dioxide
C0364159|T201|COMP|2027-1|LNC2000|Carbon dioxide|Carbon dioxide
C0364160|T201|COMP|2028-9|LNC2000|Carbon dioxide|Carbon dioxide
C0364162|T201|COMP|2030-5|LNC2000|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C0364164|T201|COMP|2032-1|LNC2000|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C0364171|T201|COMP|2039-6|LNC2000|Carcinoembryonic Ag|Carcinoembryonic Ag
C0364196|T201|COMP|2064-4|LNC2000|Ceruloplasmin|Ceruloplasmin
C0364201|T201|COMP|2069-3|LNC2000|Chloride|Chloride
C0364207|T201|COMP|2075-0|LNC2000|Chloride|Chloride
C0364209|T201|COMP|2077-6|LNC2000|Chloride|Chloride
C0364210|T201|COMP|2078-4|LNC2000|Chloride|Chloride
C0364221|T201|COMP|2085-9|LNC2000|Cholesterol.in HDL|Cholesterol.in HDL
C0364223|T201|COMP|2087-5|LNC2000|Cholesterol.in IDL|Cholesterol.in IDL
C0364225|T201|COMP|2089-1|LNC2000|Cholesterol.in LDL|Cholesterol.in LDL
C0364227|T201|COMP|2091-7|LNC2000|Cholesterol.in VLDL|Cholesterol.in VLDL
C0364236|T201|COMP|2106-3|LNC2000|Choriogonadotropin (pregnancy test)|Choriogonadotropin (pregnancy test)
C0364238|T201|COMP|2118-8|LNC2000|Choriogonadotropin (pregnancy test)|Choriogonadotropin (pregnancy test)
C0364244|T201|COMP|2110-5|LNC2000|Choriogonadotropin.beta subunit (pregnancy test)|Choriogonadotropin.beta subunit (pregnancy test)
C0364245|T201|COMP|2111-3|LNC2000|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0364246|T201|COMP|2112-1|LNC2000|Choriogonadotropin.beta subunit (pregnancy test)|Choriogonadotropin.beta subunit (pregnancy test)
C0364249|T201|COMP|2115-4|LNC2000|Choriogonadotropin.beta subunit.free|Choriogonadotropin.beta subunit.free
C0364264|T201|COMP|2132-9|LNC2000|Cobalamins|Cobalamins
C0364273|T201|COMP|2141-0|LNC2000|Corticotropin|Corticotropin
C0364274|T201|COMP|2142-8|LNC2000|Cortisol|Cortisol
C0364275|T201|COMP|2143-6|LNC2000|Cortisol|Cortisol
C0364279|T201|COMP|2147-7|LNC2000|Cortisol.free|Cortisol.free
C0364290|T201|COMP|2157-6|LNC2000|Creatine kinase|Creatine kinase
C0364292|T201|COMP|2159-2|LNC2000|Creatinine|Creatinine
C0364294|T201|COMP|2160-0|LNC2000|Creatinine|Creatinine
C0364295|T201|COMP|2161-8|LNC2000|Creatinine|Creatinine
C0364296|T201|COMP|2162-6|LNC2000|Creatinine|Creatinine
C0364298|T201|COMP|2164-2|LNC2000|Creatinine renal clearance|Creatinine renal clearance
C0364325|T201|COMP|2191-5|LNC2000|Dehydroepiandrosterone sulfate|Dehydroepiandrosterone sulfate
C0364327|T201|COMP|2193-1|LNC2000|Dehydroepiandrosterone|Dehydroepiandrosterone
C0364350|T201|COMP|2216-0|LNC2000|DOPamine|DOPamine
C0364351|T201|COMP|2217-8|LNC2000|DOPamine|DOPamine
C0364352|T201|COMP|2218-6|LNC2000|DOPamine|DOPamine
C0364367|T201|COMP|2232-7|LNC2000|EPINEPHrine|EPINEPHrine
C0364371|T201|COMP|2236-8|LNC2000|Calciferol|Calciferol
C0364378|T201|COMP|2243-4|LNC2000|Estradiol|Estradiol
C0364385|T201|COMP|2250-9|LNC2000|Estriol.unconjugated|Estriol.unconjugated
C0364386|T201|COMP|2251-7|LNC2000|Estriol|Estriol
C0364389|T201|COMP|2254-1|LNC2000|Estrogen|Estrogen
C0364393|T201|COMP|2258-2|LNC2000|Estrone|Estrone
C0364411|T201|COMP|2276-4|LNC2000|Ferritin|Ferritin
C0364417|T201|COMP|2282-2|LNC2000|Folate|Folate
C0364418|T201|COMP|2283-0|LNC2000|Folate|Folate
C0364419|T201|COMP|2284-8|LNC2000|Folate|Folate
C0364459|T201|COMP|2324-2|LNC2000|Gamma glutamyl transferase|Gamma glutamyl transferase
C0364471|T201|COMP|2333-3|LNC2000|Gastrin|Gastrin
C0364472|T201|COMP|2334-1|LNC2000|Hemoglobin.gastrointestinal|Hemoglobin.gastrointestinal
C0364473|T201|COMP|2335-8|LNC2000|Hemoglobin.gastrointestinal|Hemoglobin.gastrointestinal
C0364474|T201|COMP|2336-6|LNC2000|Globulin|Globulin
C0364479|T201|COMP|2339-0|LNC2000|Glucose|Glucose
C0364482|T201|COMP|2342-4|LNC2000|Glucose|Glucose
C0364484|T201|COMP|2344-0|LNC2000|Glucose|Glucose
C0364489|T201|COMP|2349-9|LNC2000|Glucose|Glucose
C0364490|T201|COMP|2350-7|LNC2000|Glucose|Glucose
C0364497|T201|COMP|2357-2|LNC2000|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C0364543|T201|COMP|2095-8|LNC2000|Cholesterol.in HDL/Cholesterol.total|Cholesterol.in HDL/Cholesterol.total
C0364569|T201|COMP|2428-1|LNC2000|Homocysteine|Homocysteine
C0364598|T201|COMP|2458-8|LNC2000|IgA|IgA
C0364604|T201|COMP|2464-6|LNC2000|IgG|IgG
C0364605|T201|COMP|2465-3|LNC2000|IgG|IgG
C0364606|T201|COMP|2466-1|LNC2000|IgG subclass 1|IgG subclass 1
C0364607|T201|COMP|2467-9|LNC2000|IgG subclass 2|IgG subclass 2
C0364608|T201|COMP|2468-7|LNC2000|IgG subclass 3|IgG subclass 3
C0364609|T201|COMP|2469-5|LNC2000|IgG subclass 4|IgG subclass 4
C0364612|T201|COMP|2472-9|LNC2000|IgM|IgM
C0364625|T201|COMP|2483-6|LNC2000|Insulin-like growth factor binding protein 3|Insulin-like growth factor binding protein 3
C0364626|T201|COMP|2484-4|LNC2000|Insulin-like growth factor-I|Insulin-like growth factor-I
C0364639|T201|COMP|2498-4|LNC2000|Iron|Iron
C0364641|T201|COMP|2500-7|LNC2000|Iron binding capacity|Iron binding capacity
C0364642|T201|COMP|2501-5|LNC2000|Iron binding capacity.unsaturated|Iron binding capacity.unsaturated
C0364643|T201|COMP|2502-3|LNC2000|Iron saturation|Iron saturation
C0364646|T201|COMP|2505-6|LNC2000|Iron/Iron binding capacity.total|Iron/Iron binding capacity.total
C0364654|T201|COMP|2513-0|LNC2000|Ketones|Ketones
C0364655|T201|COMP|2514-8|LNC2000|Ketones|Ketones
C0364659|T201|COMP|2518-9|LNC2000|Lactate|Lactate
C0364665|T201|COMP|2524-7|LNC2000|Lactate|Lactate
C0364671|T201|COMP|2529-6|LNC2000|Lactate dehydrogenase|Lactate dehydrogenase
C0364674|T201|COMP|2532-0|LNC2000|Lactate dehydrogenase|Lactate dehydrogenase
C0364708|T201|COMP|2093-3|LNC2000|Cholesterol|Cholesterol
C0364714|T201|COMP|2571-8|LNC2000|Triglyceride|Triglyceride
C0364741|T201|COMP|2597-3|LNC2000|Magnesium|Magnesium
C0364745|T201|COMP|2601-3|LNC2000|Magnesium|Magnesium
C0364749|T201|COMP|2605-4|LNC2000|Meat fibers|Meat fibers
C0364759|T201|COMP|2614-6|LNC2000|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C0364760|T201|COMP|2615-3|LNC2000|Methemoglobin/Hemoglobin.total|Methemoglobin/Hemoglobin.total
C0364783|T201|COMP|2638-5|LNC2000|Myelin basic protein|Myelin basic protein
C0364784|T201|COMP|2639-3|LNC2000|Myoglobin|Myoglobin
C0364785|T201|COMP|2640-1|LNC2000|Myoglobin|Myoglobin
C0364812|T201|COMP|2667-4|LNC2000|Norepinephrine|Norepinephrine
C0364813|T201|COMP|2668-2|LNC2000|Norepinephrine|Norepinephrine
C0364814|T201|COMP|2669-0|LNC2000|Normetanephrine|Normetanephrine
C0364816|T201|COMP|2671-6|LNC2000|Normetanephrine|Normetanephrine
C0364835|T201|COMP|2692-2|LNC2000|Osmolality|Osmolality
C0364838|T201|COMP|2695-5|LNC2000|Osmolality|Osmolality
C0364843|T201|COMP|2700-3|LNC2000|Oxalate|Oxalate
C0364844|T201|COMP|2701-1|LNC2000|Oxalate|Oxalate
C0364851|T201|COMP|2708-6|LNC2000|Oxygen saturation|Oxygen saturation
C0364856|T201|COMP|2713-6|LNC2000|Oxygen saturation|Oxygen saturation
C0364857|T201|COMP|2714-4|LNC2000|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C0364859|T201|COMP|2716-9|LNC2000|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C0364874|T201|COMP|2731-8|LNC2000|Parathyrin.intact|Parathyrin.intact
C0364885|T201|COMP|2742-5|LNC2000|Angiotensin converting enzyme|Angiotensin converting enzyme
C0364910|T201|COMP|2761-5|LNC2000|Phenylketones|Phenylketones
C0364923|T201|COMP|2778-9|LNC2000|Phosphate|Phosphate
C0364924|T201|COMP|2779-7|LNC2000|Phosphate|Phosphate
C0364961|T201|COMP|6298-4|LNC2000|Potassium|Potassium
C0364968|T201|COMP|2823-3|LNC2000|Potassium|Potassium
C0364971|T201|COMP|2828-2|LNC2000|Potassium|Potassium
C0364980|T201|COMP|2837-3|LNC2000|Pregnenolone|Pregnenolone
C0364982|T201|COMP|2839-9|LNC2000|Progesterone|Progesterone
C0365000|T201|COMP|2857-1|LNC2000|Prostate specific Ag|Prostate specific Ag
C0365005|T201|COMP|2862-1|LNC2000|Albumin|Albumin
C0365008|T201|COMP|2865-4|LNC2000|Alpha 1 globulin|Alpha 1 globulin
C0365011|T201|COMP|2868-8|LNC2000|Alpha 2 globulin|Alpha 2 globulin
C0365014|T201|COMP|2871-2|LNC2000|Beta globulin|Beta globulin
C0365016|T201|COMP|2873-8|LNC2000|Gamma globulin|Gamma globulin
C0365017|T201|COMP|2874-6|LNC2000|Gamma globulin|Gamma globulin
C0365023|T201|COMP|2880-3|LNC2000|Protein|Protein
C0365025|T201|COMP|2881-1|LNC2000|Protein|Protein
C0365029|T201|COMP|2885-2|LNC2000|Protein|Protein
C0365032|T201|COMP|2888-6|LNC2000|Protein|Protein
C0365033|T201|COMP|2889-4|LNC2000|Protein|Protein
C0365034|T201|COMP|2890-2|LNC2000|Protein/Creatinine|Protein/Creatinine
C0365036|T201|COMP|2892-8|LNC2000|Protoporphyrin.free|Protoporphyrin.free
C0365039|T201|COMP|2895-1|LNC2000|Protoporphyrin.zinc|Protoporphyrin.zinc
C0365044|T201|COMP|2900-9|LNC2000|Pyridoxine|Pyridoxine
C0365059|T201|COMP|2915-7|LNC2000|Renin|Renin
C0365067|T201|COMP|2923-1|LNC2000|Retinol|Retinol
C0365091|T201|COMP|2947-0|LNC2000|Sodium|Sodium
C0365095|T201|COMP|2951-2|LNC2000|Sodium|Sodium
C0365099|T201|COMP|2955-3|LNC2000|Sodium|Sodium
C0365100|T201|COMP|2956-1|LNC2000|Sodium|Sodium
C0365108|T201|COMP|2963-7|LNC2000|Somatotropin|Somatotropin
C0365111|T201|COMP|2965-2|LNC2000|Specific gravity|Specific gravity
C0365135|T201|COMP|2991-8|LNC2000|Testosterone.free|Testosterone.free
C0365137|T201|COMP|2986-8|LNC2000|Testosterone|Testosterone
C0365142|T201|COMP|2998-3|LNC2000|Thiamine|Thiamine
C0365143|T201|COMP|2999-1|LNC2000|Thiamine|Thiamine
C0365157|T201|COMP|3013-0|LNC2000|Thyroglobulin|Thyroglobulin
C0365160|T201|COMP|3016-3|LNC2000|Thyrotropin|Thyrotropin
C0365168|T201|COMP|3024-7|LNC2000|Thyroxine.free|Thyroxine.free
C0365170|T201|COMP|3026-2|LNC2000|Thyroxine|Thyroxine
C0365178|T201|COMP|3034-6|LNC2000|Transferrin|Transferrin
C0365184|T201|COMP|3040-3|LNC2000|Triacylglycerol lipase|Triacylglycerol lipase
C0365187|T201|COMP|3043-7|LNC2000|Triglyceride|Triglyceride
C0365194|T201|COMP|3050-2|LNC2000|Triiodothyronine resin uptake (T3RU)|Triiodothyronine resin uptake (T3RU)
C0365195|T201|COMP|3051-0|LNC2000|Triiodothyronine.free|Triiodothyronine.free
C0365196|T201|COMP|3052-8|LNC2000|Triiodothyronine.reverse|Triiodothyronine.reverse
C0365197|T201|COMP|3053-6|LNC2000|Triiodothyronine|Triiodothyronine
C0365228|T201|COMP|3084-1|LNC2000|Urate|Urate
C0365230|T201|COMP|3086-6|LNC2000|Urate|Urate
C0365231|T201|COMP|3087-4|LNC2000|Urate|Urate
C0365237|T201|COMP|6299-2|LNC2000|Urea nitrogen|Urea nitrogen
C0365239|T201|COMP|3093-2|LNC2000|Urea nitrogen|Urea nitrogen
C0365240|T201|COMP|3094-0|LNC2000|Urea nitrogen|Urea nitrogen
C0365241|T201|COMP|3095-7|LNC2000|Urea nitrogen|Urea nitrogen
C0365242|T201|COMP|3096-5|LNC2000|Urea nitrogen|Urea nitrogen
C0365243|T201|COMP|3097-3|LNC2000|Urea nitrogen/Creatinine|Urea nitrogen/Creatinine
C0365253|T201|COMP|3107-0|LNC2000|Urobilinogen|Urobilinogen
C0365268|T201|COMP|3122-9|LNC2000|Vanillylmandelate|Vanillylmandelate
C0365305|T201|COMP|3160-9|LNC2000|Specimen volume|Specimen volume
C0365312|T201|COMP|3167-4|LNC2000|Specimen volume|Specimen volume
C0365325|T201|COMP|3181-5|LNC2000|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C0365326|T201|COMP|3182-3|LNC2000|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C0365329|T201|COMP|6303-2|LNC2000|Coagulation dilute Russell viper venom induced|Coagulation dilute Russell viper venom induced
C0365392|T201|COMP|3173-2|LNC2000|Coagulation surface induced|Coagulation surface induced
C0365531|T201|COMP|3297-9|LNC2000|Acetaminophen|Acetaminophen
C0365532|T201|COMP|3298-7|LNC2000|Acetaminophen|Acetaminophen
C0365533|T201|COMP|3299-5|LNC2000|Acetaminophen|Acetaminophen
C0365583|T201|COMP|3349-8|LNC2000|Amphetamines|Amphetamines
C0365608|T201|COMP|3376-1|LNC2000|Barbiturates|Barbiturates
C0365609|T201|COMP|3377-9|LNC2000|Barbiturates|Barbiturates
C0365619|T201|COMP|3389-4|LNC2000|Benzodiazepines|Benzodiazepines
C0365620|T201|COMP|3390-2|LNC2000|Benzodiazepines|Benzodiazepines
C0365627|T201|COMP|3397-7|LNC2000|Cocaine|Cocaine
C0365644|T201|COMP|3414-0|LNC2000|Buprenorphine|Buprenorphine
C0365652|T201|COMP|3422-3|LNC2000|Caffeine|Caffeine
C0365656|T201|COMP|3426-4|LNC2000|Tetrahydrocannabinol|Tetrahydrocannabinol
C0365661|T201|COMP|3432-2|LNC2000|carBAMazepine|carBAMazepine
C0365665|T201|COMP|3436-3|LNC2000|Carboxy tetrahydrocannabinol|Carboxy tetrahydrocannabinol
C0365736|T201|COMP|3507-1|LNC2000|Codeine|Codeine
C0365749|T201|COMP|3520-4|LNC2000|cycloSPORINE|cycloSPORINE
C0365773|T201|COMP|19141-1|LNC2000|Propoxyphene|Propoxyphene
C0365774|T201|COMP|3545-1|LNC2000|Propoxyphene|Propoxyphene
C0365892|T201|COMP|3663-2|LNC2000|Gentamicin^peak|Gentamicin^peak
C0365894|T201|COMP|3665-7|LNC2000|Gentamicin^trough|Gentamicin^trough
C0365943|T201|COMP|3714-3|LNC2000|Lidocaine|Lidocaine
C0365948|T201|COMP|3719-2|LNC2000|Lithium|Lithium
C0365974|T201|COMP|3746-5|LNC2000|Meperidine|Meperidine
C0366000|T201|COMP|3773-9|LNC2000|Methadone|Methadone
C0366006|T201|COMP|3779-6|LNC2000|Methamphetamine|Methamphetamine
C0366013|T201|COMP|3786-1|LNC2000|Methaqualone|Methaqualone
C0366057|T201|COMP|3830-7|LNC2000|Morphine|Morphine
C0366081|T201|COMP|3854-7|LNC2000|Nicotine|Nicotine
C0366088|T201|COMP|3861-2|LNC2000|Nordiazepam|Nordiazepam
C0366106|T201|COMP|3879-4|LNC2000|Opiates|Opiates
C0366163|T201|COMP|3936-2|LNC2000|Phencyclidine|Phencyclidine
C0366175|T201|COMP|3948-7|LNC2000|PHENobarbital|PHENobarbital
C0366195|T201|COMP|3968-5|LNC2000|Phenytoin|Phenytoin
C0366196|T201|COMP|3969-3|LNC2000|Phenytoin.free|Phenytoin.free
C0366250|T201|COMP|4023-8|LNC2000|Salicylates|Salicylates
C0366251|T201|COMP|4024-6|LNC2000|Salicylates|Salicylates
C0366275|T201|COMP|4049-3|LNC2000|Theophylline|Theophylline
C0366283|T201|COMP|4057-6|LNC2000|Tobramycin^peak|Tobramycin^peak
C0366285|T201|COMP|4059-2|LNC2000|Tobramycin^trough|Tobramycin^trough
C0366299|T201|COMP|4073-3|LNC2000|Tricyclic antidepressants|Tricyclic antidepressants
C0366312|T201|COMP|4086-5|LNC2000|Valproate|Valproate
C0366316|T201|COMP|4090-7|LNC2000|Vancomycin^peak|Vancomycin^peak
C0366318|T201|COMP|4092-3|LNC2000|Vancomycin^trough|Vancomycin^trough
C0366702|T201|COMP|4477-6|LNC2000|Complement C1 esterase inhibitor|Complement C1 esterase inhibitor
C0366711|T201|COMP|4485-9|LNC2000|Complement C3|Complement C3
C0366727|T201|COMP|4498-2|LNC2000|Complement C4|Complement C4
C0366770|T201|COMP|4537-7|LNC2000|Erythrocyte sedimentation rate|Erythrocyte sedimentation rate
C0366775|T201|COMP|4542-7|LNC2000|Haptoglobin|Haptoglobin
C0366777|T201|COMP|4544-3|LNC2000|Hematocrit|Hematocrit
C0366778|T201|COMP|4545-0|LNC2000|Hematocrit|Hematocrit
C0366779|T201|COMP|4546-8|LNC2000|Hemoglobin A/Hemoglobin.total|Hemoglobin A/Hemoglobin.total
C0366780|T201|COMP|4547-6|LNC2000|Hemoglobin A1/Hemoglobin.total|Hemoglobin A1/Hemoglobin.total
C0366781|T201|COMP|4548-4|LNC2000|Hemoglobin A1c/Hemoglobin.total|Hemoglobin A1c/Hemoglobin.total
C0366784|T201|COMP|4551-8|LNC2000|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C0366785|T201|COMP|4552-6|LNC2000|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C0366794|T201|COMP|4563-3|LNC2000|Hemoglobin C/Hemoglobin.total|Hemoglobin C/Hemoglobin.total
C0366802|T201|COMP|4569-0|LNC2000|Hemoglobin D/Hemoglobin.total|Hemoglobin D/Hemoglobin.total
C0366806|T201|COMP|4575-7|LNC2000|Hemoglobin E/Hemoglobin.total|Hemoglobin E/Hemoglobin.total
C0366811|T201|COMP|4633-4|LNC2000|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C0366812|T201|COMP|4576-5|LNC2000|Hemoglobin F/Hemoglobin.total|Hemoglobin F/Hemoglobin.total
C0366856|T201|COMP|4621-9|LNC2000|Hemoglobin S|Hemoglobin S
C0366860|T201|COMP|4625-0|LNC2000|Hemoglobin S/Hemoglobin.total|Hemoglobin S/Hemoglobin.total
C0366908|T201|COMP|4679-7|LNC2000|Reticulocytes/100 erythrocytes|Reticulocytes/100 erythrocytes
C0367223|T201|COMP|584-3|LNC2000|Streptococcus agalactiae|Streptococcus agalactiae
C0367227|T201|COMP|5034-4|LNC2000|Streptococcus agalactiae rRNA|Streptococcus agalactiae rRNA
C0367235|T201|COMP|6462-6|LNC2000|Bacteria identified|Bacteria identified
C0367237|T201|COMP|634-6|LNC2000|Bacteria identified|Bacteria identified
C0367238|T201|COMP|635-3|LNC2000|Bacteria identified|Bacteria identified
C0367244|T201|COMP|6463-4|LNC2000|Bacteria identified|Bacteria identified
C0367245|T201|COMP|5036-9|LNC2000|Streptococcus pyogenes rRNA|Streptococcus pyogenes rRNA
C0367246|T201|COMP|546-2|LNC2000|Streptococcus.beta-hemolytic|Streptococcus.beta-hemolytic
C0367247|T201|COMP|547-0|LNC2000|Streptococcus.beta-hemolytic|Streptococcus.beta-hemolytic
C0367250|T201|COMP|5370-2|LNC2000|Streptolysin O Ab|Streptolysin O Ab
C0367268|T201|COMP|5388-4|LNC2000|Toxoplasma gondii Ab.IgG|Toxoplasma gondii Ab.IgG
C0367271|T201|COMP|5390-0|LNC2000|Toxoplasma gondii Ab.IgM|Toxoplasma gondii Ab.IgM
C0367281|T201|COMP|5393-4|LNC2000|Treponema pallidum Ab|Treponema pallidum Ab
C0367283|T201|COMP|6561-5|LNC2000|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C0367289|T201|COMP|6565-6|LNC2000|Trichomonas vaginalis|Trichomonas vaginalis
C0367301|T201|COMP|6568-0|LNC2000|Trichomonas vaginalis rRNA|Trichomonas vaginalis rRNA
C0367308|T201|COMP|5403-1|LNC2000|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0367314|T201|COMP|5404-9|LNC2000|Varicella zoster virus Ab.IgM|Varicella zoster virus Ab.IgM
C0367350|T201|COMP|673-4|LNC2000|Ova & parasites identified|Ova & parasites identified
C0367394|T201|COMP|5048-4|LNC2000|Nuclear Ab|Nuclear Ab
C0367396|T201|COMP|5076-5|LNC2000|Cardiolipin Ab.IgA|Cardiolipin Ab.IgA
C0367401|T201|COMP|5117-7|LNC2000|Cryoglobulin|Cryoglobulin
C0367402|T201|COMP|6476-6|LNC2000|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0367411|T201|COMP|5130-0|LNC2000|DNA double strand Ab|DNA double strand Ab
C0367418|T201|COMP|5170-6|LNC2000|Gliadin Ab.IgG|Gliadin Ab.IgG
C0367421|T201|COMP|533-0|LNC2000|Mycobacterium sp identified|Mycobacterium sp identified
C0367435|T201|COMP|5247-2|LNC2000|Mitochondria Ab|Mitochondria Ab
C0367444|T201|COMP|543-9|LNC2000|Mycobacterium sp identified|Mycobacterium sp identified
C0367449|T201|COMP|5297-7|LNC2000|Rheumatoid factor|Rheumatoid factor
C0367470|T201|COMP|5358-7|LNC2000|Smooth muscle Ab|Smooth muscle Ab
C0367476|T201|COMP|5255-5|LNC2000|Mycoplasma pneumoniae Ab.IgG|Mycoplasma pneumoniae Ab.IgG
C0367478|T201|COMP|5256-3|LNC2000|Mycoplasma pneumoniae Ab.IgM|Mycoplasma pneumoniae Ab.IgM
C0367512|T201|COMP|688-2|LNC2000|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367539|T201|COMP|693-2|LNC2000|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367584|T201|COMP|697-3|LNC2000|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367589|T201|COMP|698-1|LNC2000|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C0367607|T201|COMP|5028-6|LNC2000|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C0367700|T201|COMP|5568-1|LNC2000|Acetone|Acetone
C0367701|T201|COMP|5569-9|LNC2000|Acetone|Acetone
C0367720|T201|COMP|5583-0|LNC2000|Arsenic|Arsenic
C0367722|T201|COMP|5869-3|LNC2000|Parainfluenza virus 1 Ag|Parainfluenza virus 1 Ag
C0367774|T201|COMP|5273-8|LNC2000|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0367775|T201|COMP|5274-6|LNC2000|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0367784|T201|COMP|3393-6|LNC2000|Benzoylecgonine|Benzoylecgonine
C0367788|T201|COMP|5631-7|LNC2000|Copper|Copper
C0367797|T201|COMP|5640-8|LNC2000|Ethanol|Ethanol
C0367798|T201|COMP|5639-0|LNC2000|Ethanol|Ethanol
C0367801|T201|COMP|5643-2|LNC2000|Ethanol|Ethanol
C0367802|T201|COMP|5644-0|LNC2000|Ethanol|Ethanol
C0367803|T201|COMP|5645-7|LNC2000|Ethanol|Ethanol
C0367809|T201|COMP|5646-5|LNC2000|Ethylene glycol|Ethylene glycol
C0367855|T201|COMP|5669-7|LNC2000|Isopropanol|Isopropanol
C0367857|T201|COMP|5671-3|LNC2000|Lead|Lead
C0367871|T201|COMP|5685-3|LNC2000|Mercury|Mercury
C0367879|T201|COMP|5290-2|LNC2000|Reagin Ab|Reagin Ab
C0367888|T201|COMP|5292-8|LNC2000|Reagin Ab|Reagin Ab
C0367894|T201|COMP|5876-8|LNC2000|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C0367895|T201|COMP|5877-6|LNC2000|Respiratory syncytial virus Ag|Respiratory syncytial virus Ag
C0367930|T201|COMP|5724-0|LNC2000|Selenium|Selenium
C0367978|T201|COMP|5763-8|LNC2000|Zinc|Zinc
C0367981|T201|COMP|5766-1|LNC2000|Ammonium urate crystals|Ammonium urate crystals
C0367982|T201|COMP|5767-9|LNC2000|Appearance|Appearance
C0367984|T201|COMP|5769-5|LNC2000|Bacteria|Bacteria
C0367985|T201|COMP|5770-3|LNC2000|Bilirubin|Bilirubin
C0367986|T201|COMP|5771-1|LNC2000|Bilirubin crystals|Bilirubin crystals
C0367990|T201|COMP|5773-7|LNC2000|Calcium carbonate crystals|Calcium carbonate crystals
C0367994|T201|COMP|5774-5|LNC2000|Calcium oxalate crystals|Calcium oxalate crystals
C0367999|T201|COMP|5775-2|LNC2000|Calcium phosphate crystals|Calcium phosphate crystals
C0368000|T201|COMP|5776-0|LNC2000|Calcium sulfate crystals|Calcium sulfate crystals
C0368001|T201|COMP|5777-8|LNC2000|Cholesterol crystals|Cholesterol crystals
C0368002|T201|COMP|5778-6|LNC2000|Color|Color
C0368005|T201|COMP|5781-0|LNC2000|Crystals|Crystals
C0368006|T201|COMP|5782-8|LNC2000|Crystals|Crystals
C0368007|T201|COMP|5783-6|LNC2000|Crystals.unidentified|Crystals.unidentified
C0368008|T201|COMP|5784-4|LNC2000|Cystine crystals|Cystine crystals
C0368009|T201|COMP|5785-1|LNC2000|Eosinophils|Eosinophils
C0368010|T201|COMP|5786-9|LNC2000|Epithelial casts|Epithelial casts
C0368011|T201|COMP|5787-7|LNC2000|Epithelial cells|Epithelial cells
C0368012|T201|COMP|5807-3|LNC2000|Erythrocyte casts|Erythrocyte casts
C0368013|T201|COMP|5808-1|LNC2000|Erythrocytes|Erythrocytes
C0368014|T201|COMP|5788-5|LNC2000|Oval fat bodies (globules)|Oval fat bodies (globules)
C0368015|T201|COMP|5789-3|LNC2000|Fatty casts|Fatty casts
C0368017|T201|COMP|5791-9|LNC2000|Fungi.yeastlike|Fungi.yeastlike
C0368018|T201|COMP|5792-7|LNC2000|Glucose|Glucose
C0368020|T201|COMP|5794-3|LNC2000|Hemoglobin|Hemoglobin
C0368021|T201|COMP|5793-5|LNC2000|Granular casts|Granular casts
C0368022|T201|COMP|5795-0|LNC2000|Hippurate crystals|Hippurate crystals
C0368025|T201|COMP|5796-8|LNC2000|Hyaline casts|Hyaline casts
C0368028|T201|COMP|5880-0|LNC2000|Rotavirus Ag|Rotavirus Ag
C0368032|T201|COMP|5797-6|LNC2000|Ketones|Ketones
C0368033|T201|COMP|5798-4|LNC2000|Leucine crystals|Leucine crystals
C0368034|T201|COMP|5820-6|LNC2000|Leukocyte casts|Leukocyte casts
C0368035|T201|COMP|5799-2|LNC2000|Leukocyte esterase|Leukocyte esterase
C0368036|T201|COMP|5821-4|LNC2000|Leukocytes|Leukocytes
C0368039|T201|COMP|5332-2|LNC2000|Rubella virus Ab|Rubella virus Ab
C0368040|T201|COMP|5802-4|LNC2000|Nitrite|Nitrite
C0368043|T201|COMP|5804-0|LNC2000|Protein|Protein
C0368044|T201|COMP|5334-8|LNC2000|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0368045|T201|COMP|5335-5|LNC2000|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C0368058|T201|COMP|5809-9|LNC2000|Reducing substances|Reducing substances
C0368061|T201|COMP|5811-5|LNC2000|Specific gravity|Specific gravity
C0368062|T201|COMP|5812-3|LNC2000|Sulfonamide crystals|Sulfonamide crystals
C0368063|T201|COMP|5813-1|LNC2000|Trichomonas vaginalis|Trichomonas vaginalis
C0368065|T201|COMP|5814-9|LNC2000|Triple phosphate crystals|Triple phosphate crystals
C0368075|T201|COMP|5815-6|LNC2000|Tyrosine crystals|Tyrosine crystals
C0368077|T201|COMP|5817-2|LNC2000|Urate crystals|Urate crystals
C0368078|T201|COMP|5818-0|LNC2000|Urobilinogen|Urobilinogen
C0368079|T201|COMP|5819-8|LNC2000|Waxy casts|Waxy casts
C0368080|T201|COMP|5822-2|LNC2000|Yeast|Yeast
C0368096|T201|COMP|5834-7|LNC2000|Adenovirus Ag|Adenovirus Ag
C0368105|T201|COMP|5052-6|LNC2000|Aspergillus sp Ab|Aspergillus sp Ab
C0368106|T201|COMP|5053-4|LNC2000|Aspergillus sp Ab|Aspergillus sp Ab
C0368113|T201|COMP|5057-5|LNC2000|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0368123|T201|COMP|550-4|LNC2000|Bordetella pertussis Ag|Bordetella pertussis Ag
C0368129|T201|COMP|5062-5|LNC2000|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0368132|T201|COMP|5064-1|LNC2000|Borrelia burgdorferi Ab.IgM|Borrelia burgdorferi Ab.IgM
C0368136|T201|COMP|4991-6|LNC2000|Borrelia burgdorferi DNA|Borrelia burgdorferi DNA
C0368155|T201|COMP|6331-3|LNC2000|Campylobacter sp identified|Campylobacter sp identified
C0368180|T201|COMP|560-3|LNC2000|Chlamydia sp identified|Chlamydia sp identified
C0368193|T201|COMP|6349-5|LNC2000|Chlamydia trachomatis|Chlamydia trachomatis
C0368205|T201|COMP|6357-8|LNC2000|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0368206|T201|COMP|4993-2|LNC2000|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C0368219|T201|COMP|6367-7|LNC2000|Clostridium tetani Ab.IgG|Clostridium tetani Ab.IgG
C0368221|T201|COMP|5095-5|LNC2000|Coccidioides immitis Ab|Coccidioides immitis Ab
C0368222|T201|COMP|5096-3|LNC2000|Coccidioides immitis Ab|Coccidioides immitis Ab
C0368259|T201|COMP|5124-3|LNC2000|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0368261|T201|COMP|5126-8|LNC2000|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0368262|T201|COMP|5127-6|LNC2000|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0368268|T201|COMP|6379-2|LNC2000|Cytomegalovirus Ag|Cytomegalovirus Ag
C0368274|T201|COMP|5000-5|LNC2000|Cytomegalovirus DNA|Cytomegalovirus DNA
C0368278|T201|COMP|5838-8|LNC2000|Cytomegalovirus|Cytomegalovirus
C0368326|T201|COMP|5005-4|LNC2000|Epstein Barr virus DNA|Epstein Barr virus DNA
C0368356|T201|COMP|575-1|LNC2000|Fungus identified|Fungus identified
C0368362|T201|COMP|17949-9|LNC2000|Fungus identified^^^4|Fungus identified^^^4
C0368363|T201|COMP|6410-5|LNC2000|Gardnerella vaginalis rRNA|Gardnerella vaginalis rRNA
C0368366|T201|COMP|6412-1|LNC2000|Giardia lamblia Ag|Giardia lamblia Ag
C0368380|T201|COMP|6420-4|LNC2000|Helicobacter pylori Ab.IgA|Helicobacter pylori Ab.IgA
C0368381|T201|COMP|5176-3|LNC2000|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C0368382|T201|COMP|5177-1|LNC2000|Helicobacter pylori Ab.IgM|Helicobacter pylori Ab.IgM
C0368385|T201|COMP|5181-3|LNC2000|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C0368387|T201|COMP|5183-9|LNC2000|Hepatitis A virus Ab|Hepatitis A virus Ab
C0368389|T201|COMP|5185-4|LNC2000|Hepatitis B virus core Ab.IgM|Hepatitis B virus core Ab.IgM
C0368391|T201|COMP|5187-0|LNC2000|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C0368401|T201|COMP|5193-8|LNC2000|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0368402|T201|COMP|5194-6|LNC2000|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0368403|T201|COMP|5195-3|LNC2000|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C0368404|T201|COMP|5196-1|LNC2000|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C0368406|T201|COMP|5198-7|LNC2000|Hepatitis C virus Ab|Hepatitis C virus Ab
C0368407|T201|COMP|5199-5|LNC2000|Hepatitis C virus Ab|Hepatitis C virus Ab
C0368420|T201|COMP|5202-7|LNC2000|Herpes simplex virus Ab|Herpes simplex virus Ab
C0368434|T201|COMP|5859-4|LNC2000|Herpes simplex virus identified|Herpes simplex virus identified
C0368438|T201|COMP|5209-2|LNC2000|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0368444|T201|COMP|5213-4|LNC2000|Heterophile Ab|Heterophile Ab
C0368449|T201|COMP|5218-3|LNC2000|Histoplasma capsulatum Ab|Histoplasma capsulatum Ab
C0368456|T201|COMP|5221-7|LNC2000|HIV 1 Ab|HIV 1 Ab
C0368457|T201|COMP|5222-5|LNC2000|HIV 1 Ag|HIV 1 Ag
C0368473|T201|COMP|5862-8|LNC2000|Influenza virus A Ag|Influenza virus A Ag
C0368474|T201|COMP|5863-6|LNC2000|Influenza virus A Ag|Influenza virus A Ag
C0368478|T201|COMP|6437-8|LNC2000|Influenza virus A+B Ag|Influenza virus A+B Ag
C0368487|T201|COMP|5866-9|LNC2000|Influenza virus B Ag|Influenza virus B Ag
C0368497|T201|COMP|6448-5|LNC2000|Legionella pneumophila Ag|Legionella pneumophila Ag
C0368498|T201|COMP|588-4|LNC2000|Legionella pneumophila Ag|Legionella pneumophila Ag
C0368504|T201|COMP|593-4|LNC2000|Legionella sp identified|Legionella sp identified
C0368523|T201|COMP|5244-9|LNC2000|Measles virus Ab.IgG|Measles virus Ab.IgG
C0368530|T201|COMP|600-7|LNC2000|Bacteria identified|Bacteria identified
C0368531|T201|COMP|601-5|LNC2000|Fungus identified|Fungus identified
C0368536|T201|COMP|606-4|LNC2000|Bacteria identified|Bacteria identified
C0368539|T201|COMP|609-8|LNC2000|Bacteria identified|Bacteria identified
C0368540|T201|COMP|610-6|LNC2000|Bacteria identified|Bacteria identified
C0368541|T201|COMP|611-4|LNC2000|Bacteria identified|Bacteria identified
C0368555|T201|COMP|624-7|LNC2000|Bacteria identified|Bacteria identified
C0368556|T201|COMP|6460-0|LNC2000|Bacteria identified|Bacteria identified
C0368559|T201|COMP|626-2|LNC2000|Bacteria identified|Bacteria identified
C0368563|T201|COMP|630-4|LNC2000|Bacteria identified|Bacteria identified
C0368567|T201|COMP|5206-8|LNC2000|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C0369164|T201|COMP|12208-5|LNC2000|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0369741|T201|COMP|12238-2|LNC2000|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0482054|T201|COMP|6121-8|LNC2000|Fusarium moniliforme Ab.IgE|Fusarium moniliforme Ab.IgE
C0482057|T201|COMP|6208-3|LNC2000|Carya illinoinensis nut Ab.IgE|Carya illinoinensis nut Ab.IgE
C0482059|T201|COMP|6248-9|LNC2000|Glycine max Ab.IgE|Glycine max Ab.IgE
C0482130|T201|COMP|882-1|LNC2000|ABO & Rh group|ABO & Rh group
C0482131|T201|COMP|883-9|LNC2000|ABO group|ABO group
C0482158|T201|COMP|933-2|LNC2000|Blood product type|Blood product type
C0482217|T201|COMP|1006-6|LNC2000|Direct antiglobulin test.IgG specific reagent|Direct antiglobulin test.IgG specific reagent
C0482218|T201|COMP|1007-4|LNC2000|Direct antiglobulin test.poly specific reagent|Direct antiglobulin test.poly specific reagent
C0482535|T201|COMP|1521-4|LNC2000|Glucose^2H post meal|Glucose^2H post meal
C0482537|T201|COMP|1527-1|LNC2000|Glucose^30M post 75 g glucose PO|Glucose^30M post 75 g glucose PO
C0482539|T201|COMP|1549-5|LNC2000|Glucose^pre 100 g glucose PO|Glucose^pre 100 g glucose PO
C0482544|T201|COMP|1558-6|LNC2000|Glucose^post CFst|Glucose^post CFst
C0482590|T201|COMP|1721-0|LNC2000|Adenosine triphosphate|Adenosine triphosphate
C0482592|T201|COMP|1869-7|LNC2000|Apolipoprotein A-I|Apolipoprotein A-I
C0482602|T201|COMP|2842-3|LNC2000|Prolactin|Prolactin
C0482604|T201|COMP|3174-0|LNC2000|Antithrombin|Antithrombin
C0482605|T201|COMP|3175-7|LNC2000|Antithrombin Ag|Antithrombin Ag
C0482608|T201|COMP|3184-9|LNC2000|Activated clotting time|Activated clotting time
C0482611|T201|COMP|3187-2|LNC2000|Coagulation factor IX activity actual/Normal|Coagulation factor IX activity actual/Normal
C0482617|T201|COMP|3193-0|LNC2000|Coagulation factor V activity actual/Normal|Coagulation factor V activity actual/Normal
C0482622|T201|COMP|3198-9|LNC2000|Coagulation factor VII activity actual/Normal|Coagulation factor VII activity actual/Normal
C0482633|T201|COMP|3209-4|LNC2000|Coagulation factor VIII activity actual/Normal|Coagulation factor VIII activity actual/Normal
C0482641|T201|COMP|3218-5|LNC2000|Coagulation factor X activity actual/Normal|Coagulation factor X activity actual/Normal
C0482682|T201|COMP|5894-1|LNC2000|Coagulation tissue factor induced actual/Normal|Coagulation tissue factor induced actual/Normal
C0482691|T201|COMP|6301-6|LNC2000|Coagulation tissue factor induced.INR|Coagulation tissue factor induced.INR
C0482694|T201|COMP|5902-2|LNC2000|Coagulation tissue factor induced|Coagulation tissue factor induced
C0482696|T201|COMP|3243-3|LNC2000|Coagulation thrombin induced|Coagulation thrombin induced
C0482705|T201|COMP|3255-7|LNC2000|Fibrinogen|Fibrinogen
C0482708|T201|COMP|3256-5|LNC2000|Fibrinogen Ag|Fibrinogen Ag
C0482727|T201|COMP|3281-3|LNC2000|Lupus anticoagulant|Lupus anticoagulant
C0482730|T201|COMP|3284-7|LNC2000|Lupus anticoagulant neutralization.platelet|Lupus anticoagulant neutralization.platelet
C0482755|T201|COMP|6002-0|LNC2000|Platelet factor 4|Platelet factor 4
C0482759|T201|COMP|6007-9|LNC2000|Protein C|Protein C
C0482761|T201|COMP|6009-5|LNC2000|Protein C Ag|Protein C Ag
C0482769|T201|COMP|5892-5|LNC2000|Protein S|Protein S
C0482773|T201|COMP|6012-9|LNC2000|von Willebrand factor Ag|von Willebrand factor Ag
C0482780|T201|COMP|4532-8|LNC2000|Complement total hemolytic CH50|Complement total hemolytic CH50
C0482781|T201|COMP|4635-9|LNC2000|Hemoglobin.free|Hemoglobin.free
C0482909|T201|COMP|4821-5|LNC2000|HLA-B27|HLA-B27
C0483084|T201|COMP|5234-0|LNC2000|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C0483088|T201|COMP|5301-7|LNC2000|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0483090|T201|COMP|5348-8|LNC2000|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C0483092|T201|COMP|5351-2|LNC2000|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C0483093|T201|COMP|5352-0|LNC2000|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C0483094|T201|COMP|5353-8|LNC2000|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C0483095|T201|COMP|5354-6|LNC2000|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C0483097|T201|COMP|5356-1|LNC2000|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0483098|T201|COMP|5357-9|LNC2000|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0483102|T201|COMP|5381-9|LNC2000|Thyroglobulin Ab|Thyroglobulin Ab
C0483120|T201|COMP|5693-7|LNC2000|Methanol|Methanol
C0483147|T201|COMP|5116-9|LNC2000|Corynebacterium diphtheriae Ab|Corynebacterium diphtheriae Ab
C0483154|T201|COMP|5156-5|LNC2000|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0483155|T201|COMP|5157-3|LNC2000|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0483156|T201|COMP|5158-1|LNC2000|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0483157|T201|COMP|5159-9|LNC2000|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0483158|T201|COMP|5160-7|LNC2000|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0483171|T201|COMP|5191-2|LNC2000|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C0483558|T201|COMP|6998-9|LNC2000|cefTRIAXone|cefTRIAXone
C0483606|T201|COMP|7041-7|LNC2000|Penicillin G|Penicillin G
C0483607|T201|COMP|7042-5|LNC2000|Penicillin V|Penicillin V
C0483625|T201|COMP|7059-9|LNC2000|Vancomycin|Vancomycin
C0483642|T201|COMP|6020-2|LNC2000|Alternaria alternata Ab.IgE|Alternaria alternata Ab.IgE
C0483681|T201|COMP|7110-0|LNC2000|Baccharis spp Ab.IgE|Baccharis spp Ab.IgE
C0483694|T201|COMP|7124-1|LNC2000|Myrica spp pollen Ab.IgE|Myrica spp pollen Ab.IgE
C0483730|T201|COMP|7155-5|LNC2000|Acer negundo Ab.IgE|Acer negundo Ab.IgE
C0483759|T201|COMP|6718-1|LNC2000|Anacardium occidentale Ab.IgE|Anacardium occidentale Ab.IgE
C0483761|T201|COMP|6833-8|LNC2000|Cat dander Ab.IgE|Cat dander Ab.IgE
C0483846|T201|COMP|7258-7|LNC2000|Cow milk Ab.IgE|Cow milk Ab.IgE
C0483879|T201|COMP|7287-6|LNC2000|Anthemis cotula Ab.IgE|Anthemis cotula Ab.IgE
C0483884|T201|COMP|7291-8|LNC2000|Egg whole Ab.IgE|Egg whole Ab.IgE
C0483895|T201|COMP|6109-3|LNC2000|Ulmus americana Ab.IgE|Ulmus americana Ab.IgE
C0483969|T201|COMP|7369-2|LNC2000|Lolium perenne Ab.IgE|Lolium perenne Ab.IgE
C0484005|T201|COMP|6209-1|LNC2000|Carya illinoinensis tree Ab.IgE|Carya illinoinensis tree Ab.IgE
C0484006|T201|COMP|7407-0|LNC2000|Carya tomentosa Ab.IgE|Carya tomentosa Ab.IgE
C0484012|T201|COMP|7415-3|LNC2000|Cladosporium sphaerospermum Ab.IgE|Cladosporium sphaerospermum Ab.IgE
C0484045|T201|COMP|7445-0|LNC2000|Lactalbumin alpha Ab.IgE|Lactalbumin alpha Ab.IgE
C0484060|T201|COMP|6239-8|LNC2000|Atriplex lentiformis Ab.IgE|Atriplex lentiformis Ab.IgE
C0484080|T201|COMP|7477-3|LNC2000|Mangifera indica pollen Ab.IgE|Mangifera indica pollen Ab.IgE
C0484113|T201|COMP|6281-0|LNC2000|Morus alba Ab.IgE|Morus alba Ab.IgE
C0484138|T201|COMP|6189-5|LNC2000|Quercus alba Ab.IgE|Quercus alba Ab.IgE
C0484144|T201|COMP|6190-3|LNC2000|Avena sativa Ab.IgE|Avena sativa Ab.IgE
C0484162|T201|COMP|7558-0|LNC2000|Ostrea edulis Ab.IgE|Ostrea edulis Ab.IgE
C0484211|T201|COMP|6733-0|LNC2000|Pigeon serum Ab|Pigeon serum Ab
C0484222|T201|COMP|7613-3|LNC2000|Pistacia vera Ab.IgE|Pistacia vera Ab.IgE
C0484243|T201|COMP|7632-3|LNC2000|Ligustrum vulgare Ab.IgE|Ligustrum vulgare Ab.IgE
C0484303|T201|COMP|7691-9|LNC2000|Pecten spp Ab.IgE|Pecten spp Ab.IgE
C0484348|T201|COMP|6263-8|LNC2000|Platanus occidentalis Ab.IgE|Platanus occidentalis Ab.IgE
C0484399|T201|COMP|7774-3|LNC2000|Cow whey Ab.IgE|Cow whey Ab.IgE
C0484416|T201|COMP|7789-1|LNC2000|Acanthocytes|Acanthocytes
C0484419|T201|COMP|7790-9|LNC2000|Burr cells|Burr cells
C0484421|T201|COMP|7792-5|LNC2000|Dohle body|Dohle body
C0484424|T201|COMP|6742-1|LNC2000|Erythrocyte morphology finding|Erythrocyte morphology finding
C0484425|T201|COMP|6741-3|LNC2000|Erythrocytes|Erythrocytes
C0484428|T201|COMP|7793-3|LNC2000|Howell-Jolly bodies|Howell-Jolly bodies
C0484430|T201|COMP|6690-2|LNC2000|Leukocytes|Leukocytes
C0484437|T201|COMP|10328-3|LNC2000|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0484444|T201|COMP|7795-8|LNC2000|Pappenheimer bodies|Pappenheimer bodies
C0484446|T201|COMP|7796-6|LNC2000|Platelet clump|Platelet clump
C0484447|T201|COMP|9317-9|LNC2000|Platelets|Platelets
C0484448|T201|COMP|10378-8|LNC2000|Polychromasia|Polychromasia
C0484453|T201|COMP|7797-4|LNC2000|Rouleaux|Rouleaux
C0484454|T201|COMP|7798-2|LNC2000|Smudge cells|Smudge cells
C0484455|T201|COMP|10380-4|LNC2000|Stomatocytes|Stomatocytes
C0484456|T201|COMP|10381-2|LNC2000|Target cells|Target cells
C0484461|T201|COMP|10386-1|LNC2000|Albumin given|Albumin given
C0484485|T201|COMP|10331-7|LNC2000|Rh|Rh
C0484521|T201|COMP|8101-8|LNC2000|Cells.CD3+CD8+/100 cells|Cells.CD3+CD8+/100 cells
C0484536|T201|COMP|8112-5|LNC2000|Cells.CD3-CD16+CD56+/100 cells|Cells.CD3-CD16+CD56+/100 cells
C0484539|T201|COMP|8116-6|LNC2000|Cells.CD19|Cells.CD19
C0484540|T201|COMP|8117-4|LNC2000|Cells.CD19/100 cells|Cells.CD19/100 cells
C0484541|T201|COMP|9557-0|LNC2000|Cells.CD2|Cells.CD2
C0484542|T201|COMP|8118-2|LNC2000|Cells.CD2/100 cells|Cells.CD2/100 cells
C0484547|T201|COMP|8122-4|LNC2000|Cells.CD3|Cells.CD3
C0484548|T201|COMP|8123-2|LNC2000|Cells.CD3+CD4+/100 cells|Cells.CD3+CD4+/100 cells
C0484550|T201|COMP|8124-0|LNC2000|Cells.CD3/100 cells|Cells.CD3/100 cells
C0484556|T201|COMP|8130-7|LNC2000|Cells.CD45/100 cells|Cells.CD45/100 cells
C0484581|T201|COMP|10449-7|LNC2000|Glucose^1H post meal|Glucose^1H post meal
C0484638|T201|COMP|6768-6|LNC2000|Alkaline phosphatase|Alkaline phosphatase
C0484643|T201|COMP|10459-6|LNC2000|Alpha-1-Fetoprotein Ag|Alpha-1-Fetoprotein Ag
C0484652|T201|COMP|1798-8|LNC2000|Amylase|Amylase
C0484660|T201|COMP|10466-1|LNC2000|Anion gap 3|Anion gap 3
C0484664|T201|COMP|10333-3|LNC2000|Appearance|Appearance
C0484665|T201|COMP|1903-4|LNC2000|Ascorbate|Ascorbate
C0484670|T201|COMP|6873-4|LNC2000|Beta hydroxybutyrate|Beta hydroxybutyrate
C0484673|T201|COMP|6874-2|LNC2000|Calcium|Calcium
C0484675|T201|COMP|10334-1|LNC2000|Cancer Ag 125|Cancer Ag 125
C0484676|T201|COMP|6875-9|LNC2000|Cancer Ag 15-3|Cancer Ag 15-3
C0484683|T201|COMP|9830-1|LNC2000|Cholesterol.total/Cholesterol.in HDL|Cholesterol.total/Cholesterol.in HDL
C0484687|T201|COMP|9811-1|LNC2000|Chromogranin A|Chromogranin A
C0484692|T201|COMP|6687-8|LNC2000|Citrate|Citrate
C0484696|T201|COMP|10335-8|LNC2000|Color|Color
C0484704|T201|COMP|9812-9|LNC2000|Cortisol^PM trough specimen|Cortisol^PM trough specimen
C0484705|T201|COMP|9813-7|LNC2000|Cortisol^AM peak specimen|Cortisol^AM peak specimen
C0484731|T201|COMP|2345-7|LNC2000|Glucose|Glucose
C0484796|T201|COMP|10501-5|LNC2000|Lutropin|Lutropin
C0484825|T201|COMP|6942-7|LNC2000|Albumin|Albumin
C0484842|T201|COMP|6891-6|LNC2000|Testosterone.free+weakly bound/Testosterone.total|Testosterone.free+weakly bound/Testosterone.total
C0484848|T201|COMP|6892-4|LNC2000|Thyroxine.free|Thyroxine.free
C0484851|T201|COMP|6598-7|LNC2000|Troponin T.cardiac|Troponin T.cardiac
C0484858|T201|COMP|9624-8|LNC2000|Vanillylmandelate|Vanillylmandelate
C0484865|T201|COMP|6683-7|LNC2000|Coagulation reptilase induced|Coagulation reptilase induced
C0484920|T201|COMP|10535-3|LNC2000|Digoxin|Digoxin
C0484937|T201|COMP|9834-3|LNC2000|HYDROmorphone|HYDROmorphone
C0484942|T201|COMP|6901-3|LNC2000|Insulin.free|Insulin.free
C0484944|T201|COMP|6948-4|LNC2000|lamoTRIgine|lamoTRIgine
C0484950|T201|COMP|2609-6|LNC2000|Metanephrines|Metanephrines
C0485041|T201|COMP|10579-1|LNC2000|Leukocytes|Leukocytes
C0485042|T201|COMP|10580-9|LNC2000|Liquefaction|Liquefaction
C0485047|T201|COMP|10585-8|LNC2000|Round cells|Round cells
C0485049|T201|COMP|10587-4|LNC2000|Sexual abstinence duration|Sexual abstinence duration
C0485050|T201|COMP|6800-7|LNC2000|Spermatozoa.motile/100 spermatozoa|Spermatozoa.motile/100 spermatozoa
C0485056|T201|COMP|9704-8|LNC2000|Spermatozoa|Spermatozoa
C0485057|T201|COMP|9780-8|LNC2000|Spermatozoa|Spermatozoa
C0485085|T201|COMP|10622-9|LNC2000|Spermatozoa.normal/100 spermatozoa|Spermatozoa.normal/100 spermatozoa
C0485098|T201|COMP|9631-3|LNC2000|Viscosity|Viscosity
C0485107|T201|COMP|6864-3|LNC2000|Hemoglobin S|Hemoglobin S
C0485138|T201|COMP|9490-4|LNC2000|Aspergillus flavus Ab|Aspergillus flavus Ab
C0485143|T201|COMP|9632-1|LNC2000|Aspergillus fumigatus Ab|Aspergillus fumigatus Ab
C0485164|T201|COMP|9360-9|LNC2000|Bartonella quintana Ab.IgG|Bartonella quintana Ab.IgG
C0485166|T201|COMP|9361-7|LNC2000|Bartonella quintana Ab.IgM|Bartonella quintana Ab.IgM
C0485167|T201|COMP|7816-2|LNC2000|Blastomyces dermatitidis Ab|Blastomyces dermatitidis Ab
C0485173|T201|COMP|9588-5|LNC2000|Borrelia burgdorferi 18kD Ab.IgG|Borrelia burgdorferi 18kD Ab.IgG
C0485174|T201|COMP|9589-3|LNC2000|Borrelia burgdorferi 23kD Ab.IgG|Borrelia burgdorferi 23kD Ab.IgG
C0485175|T201|COMP|9598-4|LNC2000|Borrelia burgdorferi 23kD Ab.IgM|Borrelia burgdorferi 23kD Ab.IgM
C0485176|T201|COMP|9590-1|LNC2000|Borrelia burgdorferi 28kD Ab.IgG|Borrelia burgdorferi 28kD Ab.IgG
C0485177|T201|COMP|9591-9|LNC2000|Borrelia burgdorferi 30kD Ab.IgG|Borrelia burgdorferi 30kD Ab.IgG
C0485178|T201|COMP|9592-7|LNC2000|Borrelia burgdorferi 39kD Ab.IgG|Borrelia burgdorferi 39kD Ab.IgG
C0485179|T201|COMP|9599-2|LNC2000|Borrelia burgdorferi 39kD Ab.IgM|Borrelia burgdorferi 39kD Ab.IgM
C0485180|T201|COMP|9593-5|LNC2000|Borrelia burgdorferi 41kD Ab.IgG|Borrelia burgdorferi 41kD Ab.IgG
C0485181|T201|COMP|9587-7|LNC2000|Borrelia burgdorferi 41kD Ab.IgM|Borrelia burgdorferi 41kD Ab.IgM
C0485182|T201|COMP|9594-3|LNC2000|Borrelia burgdorferi 45kD Ab.IgG|Borrelia burgdorferi 45kD Ab.IgG
C0485183|T201|COMP|9595-0|LNC2000|Borrelia burgdorferi 58kD Ab.IgG|Borrelia burgdorferi 58kD Ab.IgG
C0485184|T201|COMP|9596-8|LNC2000|Borrelia burgdorferi 66kD Ab.IgG|Borrelia burgdorferi 66kD Ab.IgG
C0485185|T201|COMP|9597-6|LNC2000|Borrelia burgdorferi 93kD Ab.IgG|Borrelia burgdorferi 93kD Ab.IgG
C0485186|T201|COMP|9586-9|LNC2000|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0485187|T201|COMP|7817-0|LNC2000|Borrelia burgdorferi Ab.IgG|Borrelia burgdorferi Ab.IgG
C0485271|T201|COMP|9820-2|LNC2000|Cryptococcus sp Ag|Cryptococcus sp Ag
C0485332|T201|COMP|9783-2|LNC2000|Ehrlichia chaffeensis Ab.IgG|Ehrlichia chaffeensis Ab.IgG
C0485334|T201|COMP|9784-0|LNC2000|Ehrlichia chaffeensis Ab.IgM|Ehrlichia chaffeensis Ab.IgM
C0485349|T201|COMP|7883-2|LNC2000|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C0485352|T201|COMP|7885-7|LNC2000|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0485353|T201|COMP|7886-5|LNC2000|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0485371|T201|COMP|7893-1|LNC2000|Gliadin Ab|Gliadin Ab
C0485387|T201|COMP|7900-4|LNC2000|Helicobacter pylori Ab|Helicobacter pylori Ab
C0485388|T201|COMP|7901-2|LNC2000|Helicobacter pylori Ab.IgA|Helicobacter pylori Ab.IgA
C0485389|T201|COMP|7902-0|LNC2000|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C0485397|T201|COMP|7905-3|LNC2000|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C0485400|T201|COMP|9609-9|LNC2000|Hepatitis C virus 22-3 Ab|Hepatitis C virus 22-3 Ab
C0485401|T201|COMP|9610-7|LNC2000|Hepatitis C virus c33c Ab|Hepatitis C virus c33c Ab
C0485429|T201|COMP|7917-8|LNC2000|HIV 1 Ab|HIV 1 Ab
C0485431|T201|COMP|9661-0|LNC2000|HIV 1 gp120 Ab|HIV 1 gp120 Ab
C0485432|T201|COMP|9660-2|LNC2000|HIV 1 gp160 Ab|HIV 1 gp160 Ab
C0485433|T201|COMP|9662-8|LNC2000|HIV 1 gp41 Ab|HIV 1 gp41 Ab
C0485435|T201|COMP|9664-4|LNC2000|HIV 1 p24 Ab|HIV 1 p24 Ab
C0485438|T201|COMP|9666-9|LNC2000|HIV 1 p31 Ab|HIV 1 p31 Ab
C0485439|T201|COMP|9667-7|LNC2000|HIV 1 p51 Ab|HIV 1 p51 Ab
C0485440|T201|COMP|9668-5|LNC2000|HIV 1 p55 Ab|HIV 1 p55 Ab
C0485444|T201|COMP|7918-6|LNC2000|HIV 1+2 Ab|HIV 1+2 Ab
C0485481|T201|COMP|6604-3|LNC2000|Influenza virus identified|Influenza virus identified
C0485544|T201|COMP|9822-8|LNC2000|Bacteria identified|Bacteria identified
C0485584|T201|COMP|7966-5|LNC2000|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0485610|T201|COMP|10701-1|LNC2000|Ova & parasites identified|Ova & parasites identified
C0485613|T201|COMP|10704-5|LNC2000|Ova & parasites identified|Ova & parasites identified
C0485621|T201|COMP|7981-4|LNC2000|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0485623|T201|COMP|7983-0|LNC2000|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0485624|T201|COMP|7984-8|LNC2000|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0485669|T201|COMP|8014-3|LNC2000|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0485670|T201|COMP|8015-0|LNC2000|Rubella virus Ab.IgM|Rubella virus Ab.IgM
C0485752|T201|COMP|10728-4|LNC2000|Trichomonas sp identified|Trichomonas sp identified
C0485761|T201|COMP|8047-3|LNC2000|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0485795|T201|COMP|8251-1|LNC2000|Service comment|Service comment
C0485815|T201|COMP|9796-4|LNC2000|Color|Color
C0485816|T201|COMP|9795-6|LNC2000|Composition|Composition
C0485822|T201|COMP|9802-0|LNC2000|Size|Size
C0485824|T201|COMP|9804-6|LNC2000|Weight|Weight
C0485826|T201|COMP|9326-0|LNC2000|Phosphatidylserine Ab.IgG|Phosphatidylserine Ab.IgG
C0485827|T201|COMP|9327-8|LNC2000|Phosphatidylserine Ab.IgM|Phosphatidylserine Ab.IgM
C0485832|T201|COMP|8061-4|LNC2000|Nuclear Ab|Nuclear Ab
C0485843|T201|COMP|10362-2|LNC2000|Endomysium Ab.IgA|Endomysium Ab.IgA
C0485845|T201|COMP|6924-5|LNC2000|Gliadin Ab.IgA|Gliadin Ab.IgA
C0485848|T201|COMP|8072-1|LNC2000|Insulin Ab|Insulin Ab
C0485863|T201|COMP|6969-0|LNC2000|Myeloperoxidase Ab|Myeloperoxidase Ab
C0485869|T201|COMP|8087-9|LNC2000|Parietal cell Ab|Parietal cell Ab
C0485874|T201|COMP|6968-2|LNC2000|Proteinase 3 Ab|Proteinase 3 Ab
C0485882|T201|COMP|8091-1|LNC2000|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0485892|T201|COMP|8095-2|LNC2000|Smooth muscle Ab|Smooth muscle Ab
C0485899|T201|COMP|8098-6|LNC2000|Thyroglobulin Ab|Thyroglobulin Ab
C0486006|T201|COMP|8144-8|LNC2000|Amphetamines|Amphetamines
C0486008|T201|COMP|8146-3|LNC2000|Amphetamines|Amphetamines
C0486011|T201|COMP|8149-7|LNC2000|Amphetamines|Amphetamines
C0486015|T201|COMP|8150-5|LNC2000|Amphetamines|Amphetamines
C0486026|T201|COMP|9426-8|LNC2000|Barbiturates|Barbiturates
C0486032|T201|COMP|9428-4|LNC2000|Benzodiazepines|Benzodiazepines
C0486053|T201|COMP|8169-5|LNC2000|Tetrahydrocannabinol|Tetrahydrocannabinol
C0486087|T201|COMP|8187-7|LNC2000|Benzoylecgonine|Benzoylecgonine
C0486092|T201|COMP|8191-9|LNC2000|Cocaine|Cocaine
C0486103|T201|COMP|10366-3|LNC2000|Cotinine|Cotinine
C0486146|T201|COMP|8214-9|LNC2000|Opiates|Opiates
C0486148|T201|COMP|8216-4|LNC2000|Opiates|Opiates
C0486155|T201|COMP|8220-6|LNC2000|Opiates|Opiates
C0486170|T201|COMP|8234-7|LNC2000|Phencyclidine|Phencyclidine
C0486200|T201|COMP|8246-1|LNC2000|Amorphous sediment|Amorphous sediment
C0486201|T201|COMP|9335-1|LNC2000|Appearance|Appearance
C0486203|T201|COMP|9439-1|LNC2000|Casts|Casts
C0486204|T201|COMP|9842-6|LNC2000|Casts|Casts
C0486206|T201|COMP|6824-7|LNC2000|Color|Color
C0486208|T201|COMP|6825-4|LNC2000|Crystals|Crystals
C0486210|T201|COMP|8247-9|LNC2000|Mucus|Mucus
C0486211|T201|COMP|8248-7|LNC2000|Spermatozoa|Spermatozoa
C0486212|T201|COMP|8249-5|LNC2000|Transitional cells|Transitional cells
C0549703|T201|COMP|13183-9|LNC2000|Ulmus americana Ab.IgG|Ulmus americana Ab.IgG
C0549723|T201|COMP|11183-1|LNC2000|Macadamia spp Ab.IgE|Macadamia spp Ab.IgE
C0549788|T201|COMP|11281-3|LNC2000|Auer rods|Auer rods
C0549790|T201|COMP|12179-8|LNC2000|Basophils/100 leukocytes|Basophils/100 leukocytes
C0549795|T201|COMP|11282-1|LNC2000|Cells counted.total|Cells counted.total
C0549796|T201|COMP|11274-8|LNC2000|Elliptocytes|Elliptocytes
C0549797|T201|COMP|12209-3|LNC2000|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0549806|T201|COMP|11156-7|LNC2000|Leukocyte morphology finding|Leukocyte morphology finding
C0549811|T201|COMP|13349-6|LNC2000|Leukocytes|Leukocytes
C0549813|T201|COMP|13046-8|LNC2000|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C0549816|T201|COMP|11031-2|LNC2000|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0549818|T201|COMP|12229-1|LNC2000|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C0549819|T201|COMP|12230-9|LNC2000|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C0549823|T201|COMP|12234-1|LNC2000|Mesothelial cells/100 leukocytes|Mesothelial cells/100 leukocytes
C0549831|T201|COMP|12278-8|LNC2000|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0549840|T201|COMP|13047-6|LNC2000|Plasma cells/100 leukocytes|Plasma cells/100 leukocytes
C0549842|T201|COMP|11125-2|LNC2000|Platelet morphology finding|Platelet morphology finding
C0549853|T201|COMP|12248-1|LNC2000|Epithelial cells.renal|Epithelial cells.renal
C0549856|T201|COMP|12258-0|LNC2000|Epithelial cells.squamous|Epithelial cells.squamous
C0549857|T201|COMP|11276-3|LNC2000|Tubular cells|Tubular cells
C0549881|T201|COMP|13337-1|LNC2000|Cells.CD8+HLA-DR+/100 cells|Cells.CD8+HLA-DR+/100 cells
C0550178|T201|COMP|11034-6|LNC2000|Acetylcholine receptor binding Ab|Acetylcholine receptor binding Ab
C0550212|T201|COMP|13462-7|LNC2000|Apolipoprotein A-I/Apolipoprotein B|Apolipoprotein A-I/Apolipoprotein B
C0550213|T201|COMP|11135-1|LNC2000|Appearance|Appearance
C0550221|T201|COMP|11555-0|LNC2000|Base excess|Base excess
C0550237|T201|COMP|11039-5|LNC2000|C reactive protein|C reactive protein
C0550246|T201|COMP|11557-6|LNC2000|Carbon dioxide|Carbon dioxide
C0550258|T201|COMP|11054-4|LNC2000|Cholesterol.in LDL/Cholesterol.in HDL|Cholesterol.in LDL/Cholesterol.in HDL
C0550264|T201|COMP|13457-7|LNC2000|Cholesterol.in LDL|Cholesterol.in LDL
C0550265|T201|COMP|13458-5|LNC2000|Cholesterol.in VLDL|Cholesterol.in VLDL
C0550275|T201|COMP|11040-3|LNC2000|Cortisol.free|Cortisol.free
C0550279|T201|COMP|12187-1|LNC2000|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C0550281|T201|COMP|12190-5|LNC2000|Creatinine|Creatinine
C0550292|T201|COMP|13451-0|LNC2000|Creatinine dialysis fluid clearance|Creatinine dialysis fluid clearance
C0550311|T201|COMP|11043-7|LNC2000|Cryofibrinogen|Cryofibrinogen
C0550317|T201|COMP|12201-0|LNC2000|Cryoglobulin|Cryoglobulin
C0550339|T201|COMP|11046-0|LNC2000|EPINEPHrine|EPINEPHrine
C0550344|T201|COMP|12598-9|LNC2000|Fat.neutral|Fat.neutral
C0550345|T201|COMP|12215-0|LNC2000|Fatty acids.very long chain|Fatty acids.very long chain
C0550349|T201|COMP|10834-0|LNC2000|Globulin|Globulin
C0550398|T201|COMP|11050-2|LNC2000|Immunoglobulin light chains.kappa|Immunoglobulin light chains.kappa
C0550399|T201|COMP|11051-0|LNC2000|Immunoglobulin light chains.lambda|Immunoglobulin light chains.lambda
C0550413|T201|COMP|10835-7|LNC2000|Lipoprotein (little a)|Lipoprotein (little a)
C0550440|T201|COMP|11556-8|LNC2000|Oxygen|Oxygen
C0550441|T201|COMP|11559-2|LNC2000|Oxyhemoglobin/Hemoglobin.total|Oxyhemoglobin/Hemoglobin.total
C0550486|T201|COMP|10886-0|LNC2000|Prostate specific Ag.free|Prostate specific Ag.free
C0550489|T201|COMP|12851-2|LNC2000|Protein pattern|Protein pattern
C0550490|T201|COMP|13438-7|LNC2000|Protein pattern|Protein pattern
C0550491|T201|COMP|12782-9|LNC2000|Protein fractions.oligoclonal bands|Protein fractions.oligoclonal bands
C0550506|T201|COMP|11060-1|LNC2000|Reducing substances|Reducing substances
C0550528|T201|COMP|11580-8|LNC2000|Thyrotropin|Thyrotropin
C0550529|T201|COMP|11579-0|LNC2000|Thyrotropin|Thyrotropin
C0550543|T201|COMP|10839-9|LNC2000|Troponin I.cardiac|Troponin I.cardiac
C0550574|T201|COMP|11064-3|LNC2000|Urea nitrogen^post dialysis|Urea nitrogen^post dialysis
C0550575|T201|COMP|11065-0|LNC2000|Urea nitrogen^pre dialysis|Urea nitrogen^pre dialysis
C0550605|T201|COMP|10976-9|LNC2000|6-Monoacetylmorphine|6-Monoacetylmorphine
C0550678|T201|COMP|11235-9|LNC2000|fentaNYL|fentaNYL
C0550690|T201|COMP|12308-3|LNC2000|HYDROcodone|HYDROcodone
C0550753|T201|COMP|12361-2|LNC2000|Oxazepam|Oxazepam
C0550755|T201|COMP|10998-3|LNC2000|oxyCODONE|oxyCODONE
C0550795|T201|COMP|11253-2|LNC2000|Tacrolimus|Tacrolimus
C0550810|T201|COMP|11004-9|LNC2000|Tricyclic antidepressants|Tricyclic antidepressants
C0550833|T201|COMP|13088-0|LNC2000|Complement total hemolytic CH100|Complement total hemolytic CH100
C0550836|T201|COMP|11153-4|LNC2000|Hematocrit|Hematocrit
C0550839|T201|COMP|12710-0|LNC2000|Hemoglobin pattern|Hemoglobin pattern
C0550846|T201|COMP|12227-5|LNC2000|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C0550907|T201|COMP|11006-4|LNC2000|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0550913|T201|COMP|13502-0|LNC2000|Borrelia burgdorferi Ab.IgG band pattern|Borrelia burgdorferi Ab.IgG band pattern
C0550917|T201|COMP|13503-8|LNC2000|Borrelia burgdorferi Ab.IgM band pattern|Borrelia burgdorferi Ab.IgM band pattern
C0550950|T201|COMP|13227-4|LNC2000|Corynebacterium diphtheriae Ab.IgG|Corynebacterium diphtheriae Ab.IgG
C0551003|T201|COMP|11258-1|LNC2000|Hepatitis B virus DNA|Hepatitis B virus DNA
C0551004|T201|COMP|10900-9|LNC2000|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0551008|T201|COMP|11011-4|LNC2000|Hepatitis C virus RNA|Hepatitis C virus RNA
C0551009|T201|COMP|11259-9|LNC2000|Hepatitis C virus RNA|Hepatitis C virus RNA
C0551023|T201|COMP|13499-9|LNC2000|HIV 1 Ab band pattern|HIV 1 Ab band pattern
C0551027|T201|COMP|12859-5|LNC2000|HIV 1 p18 Ab|HIV 1 p18 Ab
C0551035|T201|COMP|12856-1|LNC2000|HIV 1 p65 Ab|HIV 1 p65 Ab
C0551049|T201|COMP|10853-0|LNC2000|Isospora belli|Isospora belli
C0551069|T201|COMP|12232-5|LNC2000|Measles virus Ag|Measles virus Ag
C0551072|T201|COMP|11261-5|LNC2000|Bacteria identified|Bacteria identified
C0551105|T201|COMP|13327-2|LNC2000|Parainfluenza virus Ag|Parainfluenza virus Ag
C0551144|T201|COMP|11266-4|LNC2000|Streptococcus agalactiae Ag|Streptococcus agalactiae Ag
C0551214|T201|COMP|13358-7|LNC2000|Collection time|Collection time
C0551231|T201|COMP|13169-8|LNC2000|Interpretation|Interpretation
C0551232|T201|COMP|13440-3|LNC2000|Interpretation|Interpretation
C0551288|T201|COMP|11013-0|LNC2000|DNA double strand Ab|DNA double strand Ab
C0551292|T201|COMP|10863-9|LNC2000|Endomysium Ab.IgA|Endomysium Ab.IgA
C0551303|T201|COMP|11565-9|LNC2000|Jo-1 extractable nuclear Ab|Jo-1 extractable nuclear Ab
C0551323|T201|COMP|13068-2|LNC2000|Nuclear Ab pattern|Nuclear Ab pattern
C0551356|T201|COMP|11572-5|LNC2000|Rheumatoid factor|Rheumatoid factor
C0551360|T201|COMP|11090-8|LNC2000|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C0551368|T201|COMP|8099-4|LNC2000|Thyroperoxidase Ab|Thyroperoxidase Ab
C0551435|T201|COMP|10912-4|LNC2000|Lead|Lead
C0551499|T201|COMP|12454-5|LNC2000|Urate crystals.amorphous|Urate crystals.amorphous
C0551505|T201|COMP|12210-1|LNC2000|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0551506|T201|COMP|11277-1|LNC2000|Epithelial cells.squamous|Epithelial cells.squamous
C0551507|T201|COMP|11279-7|LNC2000|Urine sediment comments|Urine sediment comments
C0796702|T201|COMP|13508-7|LNC2000|Hematocrit|Hematocrit
C0796708|T201|COMP|13514-5|LNC2000|Hemoglobin pattern|Hemoglobin pattern
C0796710|T201|COMP|13516-0|LNC2000|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0796711|T201|COMP|13517-8|LNC2000|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C0796712|T201|COMP|13518-6|LNC2000|Lymphocytes.variant/100 leukocytes|Lymphocytes.variant/100 leukocytes
C0796713|T201|COMP|13519-4|LNC2000|Basophils/100 leukocytes|Basophils/100 leukocytes
C0796715|T201|COMP|13522-8|LNC2000|Blasts/100 leukocytes|Blasts/100 leukocytes
C0796718|T201|COMP|13525-1|LNC2000|Nonhematic cells/100 leukocytes|Nonhematic cells/100 leukocytes
C0796720|T201|COMP|13527-7|LNC2000|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C0796722|T201|COMP|13529-3|LNC2000|Erythrocytes.nucleated|Erythrocytes.nucleated
C0796723|T201|COMP|13530-1|LNC2000|Erythrocytes.nucleated|Erythrocytes.nucleated
C0796725|T201|COMP|13532-7|LNC2000|Xanthochromia|Xanthochromia
C0796731|T201|COMP|13538-4|LNC2000|Carbon dioxide|Carbon dioxide
C0796780|T201|COMP|13589-7|LNC2000|Activated protein C resistance|Activated protein C resistance
C0796781|T201|COMP|13590-5|LNC2000|Activated protein C resistance|Activated protein C resistance
C0796789|T201|COMP|783-1|LNC2000|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C0796818|T201|COMP|13627-5|LNC2000|Erythrocytes|Erythrocytes
C0796846|T201|COMP|13655-6|LNC2000|Leukocytes|Leukocytes
C0797114|T201|COMP|13926-1|LNC2000|Glutamate decarboxylase 65 Ab|Glutamate decarboxylase 65 Ab
C0797129|T201|COMP|13941-0|LNC2000|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0797130|T201|COMP|13942-8|LNC2000|Spermatozoa.motile|Spermatozoa.motile
C0797131|T201|COMP|13943-6|LNC2000|Fructose|Fructose
C0797133|T201|COMP|13945-1|LNC2000|Erythrocytes|Erythrocytes
C0797135|T201|COMP|13947-7|LNC2000|Coccidioides immitis Ab.IgG|Coccidioides immitis Ab.IgG
C0797136|T201|COMP|13948-5|LNC2000|Coccidioides immitis Ab.IgM|Coccidioides immitis Ab.IgM
C0797138|T201|COMP|13950-1|LNC2000|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C0797139|T201|COMP|13951-9|LNC2000|Hepatitis A virus Ab|Hepatitis A virus Ab
C0797140|T201|COMP|13952-7|LNC2000|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C0797141|T201|COMP|13953-5|LNC2000|Hepatitis B virus little e Ab|Hepatitis B virus little e Ab
C0797142|T201|COMP|13954-3|LNC2000|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C0797143|T201|COMP|13955-0|LNC2000|Hepatitis C virus Ab|Hepatitis C virus Ab
C0797152|T201|COMP|13964-2|LNC2000|Methylmalonate|Methylmalonate
C0797153|T201|COMP|13965-9|LNC2000|Homocysteine|Homocysteine
C0797155|T201|COMP|13967-5|LNC2000|Sex hormone binding globulin|Sex hormone binding globulin
C0797157|T201|COMP|13969-1|LNC2000|Creatine kinase.MB|Creatine kinase.MB
C0797172|T201|COMP|13984-0|LNC2000|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0797174|T201|COMP|13986-5|LNC2000|Albumin/Protein.total|Albumin/Protein.total
C0797175|T201|COMP|13987-3|LNC2000|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0797176|T201|COMP|13988-1|LNC2000|Beta globulin/Protein.total|Beta globulin/Protein.total
C0797177|T201|COMP|13989-9|LNC2000|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0797178|T201|COMP|13990-7|LNC2000|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0797180|T201|COMP|13992-3|LNC2000|Albumin/Protein.total|Albumin/Protein.total
C0797181|T201|COMP|13993-1|LNC2000|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0797182|T201|COMP|13994-9|LNC2000|Beta globulin/Protein.total|Beta globulin/Protein.total
C0797183|T201|COMP|13995-6|LNC2000|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0797271|T201|COMP|14083-0|LNC2000|Epstein Barr virus early Ab|Epstein Barr virus early Ab
C0797301|T201|COMP|14115-0|LNC2000|Collagen crosslinked N-telopeptide/Creatinine|Collagen crosslinked N-telopeptide/Creatinine
C0797302|T201|COMP|14116-8|LNC2000|IgG synthesis rate|IgG synthesis rate
C0797303|T201|COMP|14117-6|LNC2000|IgG clearance/Albumin clearance|IgG clearance/Albumin clearance
C0797307|T201|COMP|14121-8|LNC2000|Pyruvate|Pyruvate
C0797321|T201|COMP|14135-8|LNC2000|Cells.CD3+CD8+|Cells.CD3+CD8+
C0797379|T201|COMP|14194-5|LNC2000|Spermatozoa.progressive/100 spermatozoa|Spermatozoa.progressive/100 spermatozoa
C0797381|T201|COMP|14196-0|LNC2000|Reticulocytes|Reticulocytes
C0797392|T201|COMP|14207-5|LNC2000|DNAse B Ab.Streptococcal|DNAse B Ab.Streptococcal
C0797431|T201|COMP|14246-3|LNC2000|Phosphatidylserine Ab.IgM|Phosphatidylserine Ab.IgM
C0797437|T201|COMP|14252-1|LNC2000|Smooth muscle Ab|Smooth muscle Ab
C0797462|T201|COMP|14277-8|LNC2000|Neutrophil cytoplasmic Ab.classic|Neutrophil cytoplasmic Ab.classic
C0797463|T201|COMP|14278-6|LNC2000|Neutrophil cytoplasmic Ab.perinuclear|Neutrophil cytoplasmic Ab.perinuclear
C0797468|T201|COMP|14286-9|LNC2000|Carnitine.free (C0)|Carnitine.free (C0)
C0797470|T201|COMP|14288-5|LNC2000|Carnitine|Carnitine
C0797495|T201|COMP|14314-9|LNC2000|Benzoylecgonine|Benzoylecgonine
C0797497|T201|COMP|14316-4|LNC2000|Benzodiazepines|Benzodiazepines
C0797515|T201|COMP|14334-7|LNC2000|Lithium|Lithium
C0797519|T201|COMP|14338-8|LNC2000|Prealbumin|Prealbumin
C0797640|T201|COMP|14463-4|LNC2000|Chlamydia trachomatis|Chlamydia trachomatis
C0797641|T201|COMP|14464-2|LNC2000|Chlamydia trachomatis|Chlamydia trachomatis
C0797642|T201|COMP|14465-9|LNC2000|Chlamydia trachomatis|Chlamydia trachomatis
C0797739|T201|COMP|14563-1|LNC2000|Hemoglobin.gastrointestinal^1st specimen|Hemoglobin.gastrointestinal^1st specimen
C0797740|T201|COMP|14564-9|LNC2000|Hemoglobin.gastrointestinal^2nd specimen|Hemoglobin.gastrointestinal^2nd specimen
C0797741|T201|COMP|14565-6|LNC2000|Hemoglobin.gastrointestinal^3rd specimen|Hemoglobin.gastrointestinal^3rd specimen
C0797754|T201|COMP|14578-9|LNC2000|ABO group|ABO group
C0797779|T201|COMP|14604-3|LNC2000|Blood group antibodies identified|Blood group antibodies identified
C0797786|T201|COMP|14611-8|LNC2000|Nuclear Ab pattern|Nuclear Ab pattern
C0797802|T201|COMP|14627-4|LNC2000|Bicarbonate|Bicarbonate
C0797838|T201|COMP|14664-7|LNC2000|Color|Color
C0797882|T201|COMP|14708-2|LNC2000|Endomysium Ab|Endomysium Ab
C0797899|T201|COMP|14725-6|LNC2000|Fluid|Fluid
C0798010|T201|COMP|14836-1|LNC2000|Methotrexate|Methotrexate
C0798036|T201|COMP|14862-7|LNC2000|Oxalate|Oxalate
C0798043|T201|COMP|14869-2|LNC2000|Pathologist review|Pathologist review
C0798049|T201|COMP|14875-9|LNC2000|Phenylalanine|Phenylalanine
C0798069|T201|COMP|14895-7|LNC2000|Protein pattern|Protein pattern
C0798079|T201|COMP|14906-2|LNC2000|Rh|Rh
C0798080|T201|COMP|14907-0|LNC2000|Rh|Rh
C0798085|T201|COMP|14912-0|LNC2000|Smudge cells/100 leukocytes|Smudge cells/100 leukocytes
C0798129|T201|COMP|14956-7|LNC2000|Albumin|Albumin
C0798130|T201|COMP|14957-5|LNC2000|Albumin|Albumin
C0798131|T201|COMP|14958-3|LNC2000|Albumin/Creatinine|Albumin/Creatinine
C0798132|T201|COMP|14959-1|LNC2000|Albumin/Creatinine|Albumin/Creatinine
C0798149|T201|COMP|14976-5|LNC2000|Lecithin/Sphingomyelin|Lecithin/Sphingomyelin
C0798152|T201|COMP|14979-9|LNC2000|Coagulation surface induced|Coagulation surface induced
C0798221|T201|COMP|15048-2|LNC2000|Creatine kinase.BB/Creatine kinase.total|Creatine kinase.BB/Creatine kinase.total
C0798222|T201|COMP|15049-0|LNC2000|Creatine kinase.MM/Creatine kinase.total|Creatine kinase.MM/Creatine kinase.total
C0798233|T201|COMP|15061-5|LNC2000|Erythropoietin|Erythropoietin
C0798239|T201|COMP|15067-2|LNC2000|Follitropin|Follitropin
C0798241|T201|COMP|15069-8|LNC2000|Fructosamine|Fructosamine
C0798321|T201|COMP|15150-6|LNC2000|Anisocytosis|Anisocytosis
C0798345|T201|COMP|15174-6|LNC2000|Cryoglobulin/Serum.total|Cryoglobulin/Serum.total
C0798351|T201|COMP|15180-3|LNC2000|Hypochromia|Hypochromia
C0798363|T201|COMP|15192-8|LNC2000|Lymphocytes.variant|Lymphocytes.variant
C0798368|T201|COMP|15197-7|LNC2000|Lymphocytes.clefted/100 leukocytes|Lymphocytes.clefted/100 leukocytes
C0798369|T201|COMP|15198-5|LNC2000|Macrocytes|Macrocytes
C0798370|T201|COMP|15199-3|LNC2000|Microcytes|Microcytes
C0798376|T201|COMP|15205-8|LNC2000|Rheumatoid factor|Rheumatoid factor
C0798381|T201|COMP|15210-8|LNC2000|Thyroglobulin Ab|Thyroglobulin Ab
C0798383|T201|COMP|15212-4|LNC2000|Triacylglycerol lipase|Triacylglycerol lipase
C0798453|T201|COMP|15283-5|LNC2000|Betula verrucosa Ab.IgE|Betula verrucosa Ab.IgE
C0798557|T201|COMP|15388-2|LNC2000|Mycoplasma hominis|Mycoplasma hominis
C0798579|T201|COMP|15410-4|LNC2000|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0798601|T201|COMP|15432-8|LNC2000|Testosterone.free/Testosterone.total|Testosterone.free/Testosterone.total
C0798698|T201|COMP|15530-9|LNC2000|Alternaria alternata Ab.IgE.RAST class|Alternaria alternata Ab.IgE.RAST class
C0798735|T201|COMP|15568-9|LNC2000|Glycine max Ab.IgE.RAST class|Glycine max Ab.IgE.RAST class
C0798810|T201|COMP|15643-0|LNC2000|Ruditapes spp Ab.IgE.RAST class|Ruditapes spp Ab.IgE.RAST class
C0799084|T201|COMP|15917-8|LNC2000|Arachis hypogaea Ab.IgE.RAST class|Arachis hypogaea Ab.IgE.RAST class
C0799239|T201|COMP|16074-7|LNC2000|Juglans spp Ab.IgE.RAST class|Juglans spp Ab.IgE.RAST class
C0799250|T201|COMP|16085-3|LNC2000|Triticum aestivum Ab.IgE.RAST class|Triticum aestivum Ab.IgE.RAST class
C0799282|T201|COMP|16117-4|LNC2000|Babesia microti Ab.IgG|Babesia microti Ab.IgG
C0799283|T201|COMP|16118-2|LNC2000|Babesia microti Ab.IgM|Babesia microti Ab.IgM
C0799291|T201|COMP|16126-5|LNC2000|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C0799293|T201|COMP|16128-1|LNC2000|Hepatitis C virus Ab|Hepatitis C virus Ab
C0799295|T201|COMP|16130-7|LNC2000|Herpes simplex virus 1 DNA|Herpes simplex virus 1 DNA
C0799296|T201|COMP|16131-5|LNC2000|Herpes simplex virus 2 DNA|Herpes simplex virus 2 DNA
C0799300|T201|COMP|16135-6|LNC2000|Beta 2 glycoprotein 1 Ab.IgG|Beta 2 glycoprotein 1 Ab.IgG
C0799301|T201|COMP|16136-4|LNC2000|Beta 2 glycoprotein 1 Ab.IgM|Beta 2 glycoprotein 1 Ab.IgM
C0799360|T201|COMP|16195-0|LNC2000|Benzodiazepines|Benzodiazepines
C0799366|T201|COMP|16201-6|LNC2000|Oxazepam|Oxazepam
C0799393|T201|COMP|16228-9|LNC2000|Nordiazepam|Nordiazepam
C0799414|T201|COMP|16249-5|LNC2000|oxyCODONE|oxyCODONE
C0799415|T201|COMP|16250-3|LNC2000|Codeine|Codeine
C0799416|T201|COMP|16251-1|LNC2000|Morphine|Morphine
C0799427|T201|COMP|16263-6|LNC2000|Calcium oxalate dihydrate crystals|Calcium oxalate dihydrate crystals
C0799428|T201|COMP|16264-4|LNC2000|Calcium oxalate monohydrate crystals|Calcium oxalate monohydrate crystals
C0799432|T201|COMP|16268-5|LNC2000|Calcium phosphate crystals|Calcium phosphate crystals
C0799525|T201|COMP|16362-6|LNC2000|Ammonia|Ammonia
C0800069|T201|COMP|16935-9|LNC2000|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0800113|T201|COMP|16982-1|LNC2000|HTLV I+II Ab|HTLV I+II Ab
C0800250|T201|COMP|17122-3|LNC2000|Cells.CD19+Kappa+/100 cells|Cells.CD19+Kappa+/100 cells
C0800251|T201|COMP|17123-1|LNC2000|Cells.CD19+Lambda+/100 cells|Cells.CD19+Lambda+/100 cells
C0800407|T201|COMP|17284-1|LNC2000|Mitochondria Ab|Mitochondria Ab
C0800515|T201|COMP|17395-5|LNC2000|oxyMORphone|oxyMORphone
C0800721|T201|COMP|17607-3|LNC2000|Specimen volume|Specimen volume
C0800823|T201|COMP|17713-9|LNC2000|Topiramate|Topiramate
C0800887|T201|COMP|17780-8|LNC2000|Helicobacter pylori Ag|Helicobacter pylori Ag
C0800895|T201|COMP|17788-1|LNC2000|Large unstained cells/100 leukocytes|Large unstained cells/100 leukocytes
C0800897|T201|COMP|17790-7|LNC2000|Leukocytes.left shift|Leukocytes.left shift
C0800898|T201|COMP|17791-5|LNC2000|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C0800899|T201|COMP|17792-3|LNC2000|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C0800900|T201|COMP|17793-1|LNC2000|Immunoglobulin light chains|Immunoglobulin light chains
C0800918|T201|COMP|17811-1|LNC2000|Alpha 1 globulin/Protein.total|Alpha 1 globulin/Protein.total
C0800920|T201|COMP|17813-7|LNC2000|Alpha 2 globulin/Protein.total|Alpha 2 globulin/Protein.total
C0800922|T201|COMP|17815-2|LNC2000|Beta globulin/Protein.total|Beta globulin/Protein.total
C0800924|T201|COMP|17817-8|LNC2000|Gamma globulin/Protein.total|Gamma globulin/Protein.total
C0800926|T201|COMP|17819-4|LNC2000|Albumin/Protein.total|Albumin/Protein.total
C0800949|T201|COMP|17842-6|LNC2000|Cancer Ag 27-29|Cancer Ag 27-29
C0800956|T201|COMP|17849-1|LNC2000|Reticulocytes/100 erythrocytes|Reticulocytes/100 erythrocytes
C0800957|T201|COMP|17850-9|LNC2000|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C0800958|T201|COMP|17851-7|LNC2000|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C0800959|T201|COMP|17852-5|LNC2000|Ureaplasma urealyticum|Ureaplasma urealyticum
C0800963|T201|COMP|17856-6|LNC2000|Hemoglobin A1c/Hemoglobin.total|Hemoglobin A1c/Hemoglobin.total
C0800966|T201|COMP|17859-0|LNC2000|Helicobacter pylori Ab.IgG|Helicobacter pylori Ab.IgG
C0800968|T201|COMP|17861-6|LNC2000|Calcium|Calcium
C0800969|T201|COMP|17862-4|LNC2000|Calcium|Calcium
C0800971|T201|COMP|17864-0|LNC2000|Calcium.ionized|Calcium.ionized
C0800980|T201|COMP|17898-8|LNC2000|Bacteria identified|Bacteria identified
C0801230|T201|COMP|18182-6|LNC2000|Osmolality|Osmolality
C0801308|T201|COMP|18262-6|LNC2000|Cholesterol.in LDL|Cholesterol.in LDL
C0801313|T201|COMP|18267-5|LNC2000|Cells.CD16+CD56+/100 cells|Cells.CD16+CD56+/100 cells
C0801328|T201|COMP|18282-4|LNC2000|Cannabinoids|Cannabinoids
C0801355|T201|COMP|18309-5|LNC2000|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C0801357|T201|COMP|18311-1|LNC2000|Pelger Huet cells|Pelger Huet cells
C0801358|T201|COMP|18312-9|LNC2000|Platelet satellitism|Platelet satellitism
C0801360|T201|COMP|18314-5|LNC2000|Morphology|Morphology
C0801361|T201|COMP|18319-4|LNC2000|Neutrophils.vacuolated|Neutrophils.vacuolated
C0801367|T201|COMP|18325-1|LNC2000|oxyMORphone|oxyMORphone
C0801432|T201|COMP|18390-5|LNC2000|Opiates|Opiates
C0801522|T201|COMP|18481-2|LNC2000|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C0801523|T201|COMP|18482-0|LNC2000|Yeast|Yeast
C0801528|T201|COMP|18487-9|LNC2000|Broad casts|Broad casts
C0801529|T201|COMP|18488-7|LNC2000|Calcium|Calcium
C0801853|T201|COMP|18860-7|LNC2000|Amikacin|Amikacin
C0801855|T201|COMP|18862-3|LNC2000|Amoxicillin+Clavulanate|Amoxicillin+Clavulanate
C0801857|T201|COMP|18864-9|LNC2000|Ampicillin|Ampicillin
C0801858|T201|COMP|18865-6|LNC2000|Ampicillin+Sulbactam|Ampicillin+Sulbactam
C0801861|T201|COMP|18868-0|LNC2000|Aztreonam|Aztreonam
C0801871|T201|COMP|18878-9|LNC2000|ceFAZolin|ceFAZolin
C0801872|T201|COMP|18879-7|LNC2000|Cefepime|Cefepime
C0801879|T201|COMP|18886-2|LNC2000|Cefotaxime|Cefotaxime
C0801880|T201|COMP|18887-0|LNC2000|cefoTEtan|cefoTEtan
C0801886|T201|COMP|18893-8|LNC2000|cefTAZidime|cefTAZidime
C0801888|T201|COMP|18895-3|LNC2000|cefTRIAXone|cefTRIAXone
C0801896|T201|COMP|18903-5|LNC2000|Chloramphenicol|Chloramphenicol
C0801899|T201|COMP|18906-8|LNC2000|Ciprofloxacin|Ciprofloxacin
C0801901|T201|COMP|18908-4|LNC2000|Clindamycin|Clindamycin
C0801912|T201|COMP|18919-1|LNC2000|Erythromycin|Erythromycin
C0801921|T201|COMP|18928-2|LNC2000|Gentamicin|Gentamicin
C0801922|T201|COMP|18929-0|LNC2000|Gentamicin.high potency|Gentamicin.high potency
C0801925|T201|COMP|18932-4|LNC2000|Imipenem|Imipenem
C0801936|T201|COMP|18943-1|LNC2000|Meropenem|Meropenem
C0801948|T201|COMP|18955-5|LNC2000|Nitrofurantoin|Nitrofurantoin
C0801954|T201|COMP|18961-3|LNC2000|Oxacillin|Oxacillin
C0801957|T201|COMP|18964-7|LNC2000|Penicillin|Penicillin
C0801958|T201|COMP|18965-4|LNC2000|Penicillin G|Penicillin G
C0801962|T201|COMP|18969-6|LNC2000|Piperacillin|Piperacillin
C0801963|T201|COMP|18970-4|LNC2000|Piperacillin+Tazobactam|Piperacillin+Tazobactam
C0801967|T201|COMP|18974-6|LNC2000|rifAMPin|rifAMPin
C0801976|T201|COMP|18983-7|LNC2000|Streptomycin.high potency|Streptomycin.high potency
C0801986|T201|COMP|18993-6|LNC2000|Tetracycline|Tetracycline
C0801989|T201|COMP|18996-9|LNC2000|Tobramycin|Tobramycin
C0801991|T201|COMP|18998-5|LNC2000|Trimethoprim+Sulfamethoxazole|Trimethoprim+Sulfamethoxazole
C0801993|T201|COMP|19000-9|LNC2000|Vancomycin|Vancomycin
C0802013|T201|COMP|19057-9|LNC2000|ABO & Rh group|ABO & Rh group
C0802016|T201|COMP|888-8|LNC2000|Blood group antibodies identified|Blood group antibodies identified
C0802019|T201|COMP|19066-0|LNC2000|Blood bank comment|Blood bank comment
C0802022|T201|COMP|19074-4|LNC2000|Carnitine esters|Carnitine esters
C0802023|T201|COMP|19075-1|LNC2000|Cells counted.total|Cells counted.total
C0802024|T201|COMP|19076-9|LNC2000|Cells counted.total|Cells counted.total
C0802025|T201|COMP|19077-7|LNC2000|Cells identified|Cells identified
C0802028|T201|COMP|19080-1|LNC2000|Choriogonadotropin|Choriogonadotropin
C0802029|T201|COMP|13362-9|LNC2000|Collection duration|Collection duration
C0802030|T201|COMP|19086-8|LNC2000|Collection end date|Collection end date
C0802031|T201|COMP|19087-6|LNC2000|Collection end time|Collection end time
C0802032|T201|COMP|19088-4|LNC2000|Collection start date|Collection start date
C0802033|T201|COMP|19089-2|LNC2000|Collection start time|Collection start time
C0802038|T201|COMP|19098-3|LNC2000|Erythrocytes|Erythrocytes
C0802045|T201|COMP|19107-2|LNC2000|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C0802046|T201|COMP|19108-0|LNC2000|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C0802050|T201|COMP|19113-0|LNC2000|IgE|IgE
C0802053|T201|COMP|19123-9|LNC2000|Magnesium|Magnesium
C0802055|T201|COMP|19125-4|LNC2000|Meconium|Meconium
C0802056|T201|COMP|19126-2|LNC2000|Bacteria identified|Bacteria identified
C0802058|T201|COMP|19128-8|LNC2000|Bacteria identified|Bacteria identified
C0802069|T201|COMP|19145-2|LNC2000|Reference lab test name|Reference lab test name
C0802070|T201|COMP|19146-0|LNC2000|Reference lab test results|Reference lab test results
C0802077|T201|COMP|19153-6|LNC2000|Specimen volume|Specimen volume
C0802079|T201|COMP|19157-7|LNC2000|Tube number|Tube number
C0802082|T201|COMP|19161-9|LNC2000|Urobilinogen|Urobilinogen
C0802083|T201|COMP|19162-7|LNC2000|Varicella zoster virus Ab.IgG|Varicella zoster virus Ab.IgG
C0802092|T201|COMP|19171-8|LNC2000|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0802118|T201|COMP|19201-3|LNC2000|Prostate specific Ag.free|Prostate specific Ag.free
C0802148|T201|COMP|19244-3|LNC2000|Character|Character
C0802157|T201|COMP|19254-2|LNC2000|Oxygen^^adjusted to patient's actual temperature|Oxygen^^adjusted to patient's actual temperature
C0802161|T201|COMP|19261-7|LNC2000|Amphetamines|Amphetamines
C0802169|T201|COMP|19270-8|LNC2000|Barbiturates|Barbiturates
C0802184|T201|COMP|19287-2|LNC2000|Cannabinoids tested for|Cannabinoids tested for
C0802192|T201|COMP|19295-5|LNC2000|Opiates|Opiates
C0802193|T201|COMP|19296-3|LNC2000|Opiates tested for|Opiates tested for
C0802209|T201|COMP|19312-8|LNC2000|Tricyclic antidepressants|Tricyclic antidepressants
C0802237|T201|COMP|19343-3|LNC2000|Amphetamine|Amphetamine
C0802301|T201|COMP|19415-9|LNC2000|Tetrahydrocannabinol|Tetrahydrocannabinol
C0802315|T201|COMP|19429-0|LNC2000|Propoxyphene|Propoxyphene
C0802425|T201|COMP|19550-3|LNC2000|Methadone|Methadone
C0802428|T201|COMP|19554-5|LNC2000|Methamphetamine|Methamphetamine
C0802464|T201|COMP|19593-3|LNC2000|6-Monoacetylmorphine|6-Monoacetylmorphine
C0802508|T201|COMP|19643-6|LNC2000|oxyCODONE|oxyCODONE
C0802522|T201|COMP|19659-2|LNC2000|Phencyclidine|Phencyclidine
C0802566|T201|COMP|19710-3|LNC2000|traMADol|traMADol
C0802579|T201|COMP|19763-2|LNC2000|Specimen source|Specimen source
C0802580|T201|COMP|19764-0|LNC2000|Statement of adequacy|Statement of adequacy
C0802583|T201|COMP|19767-3|LNC2000|Cytologist|Cytologist
C0802584|T201|COMP|19768-1|LNC2000|Reviewing cytologist|Reviewing cytologist
C0802585|T201|COMP|19769-9|LNC2000|Pathologist|Pathologist
C0802588|T201|COMP|19773-1|LNC2000|Recommended follow-up|Recommended follow-up
C0802589|T201|COMP|19774-9|LNC2000|Cytology study comment|Cytology study comment
C0803213|T201|COMP|20398-4|LNC2000|Nuclear Ab pattern.homogeneous|Nuclear Ab pattern.homogeneous
C0803214|T201|COMP|20399-2|LNC2000|Nuclear Ab pattern.nucleolar|Nuclear Ab pattern.nucleolar
C0803216|T201|COMP|20401-6|LNC2000|Nuclear Ab pattern.speckled|Nuclear Ab pattern.speckled
C0803217|T201|COMP|20402-4|LNC2000|Cells.CD16+CD56+|Cells.CD16+CD56+
C0803219|T201|COMP|20404-0|LNC2000|Fibronectin.fetal|Fibronectin.fetal
C0803220|T201|COMP|20405-7|LNC2000|Urobilinogen|Urobilinogen
C0803223|T201|COMP|20408-1|LNC2000|Leukocytes|Leukocytes
C0803224|T201|COMP|20409-9|LNC2000|Erythrocytes|Erythrocytes
C0803231|T201|COMP|20416-4|LNC2000|Hepatitis C virus RNA|Hepatitis C virus RNA
C0803235|T201|COMP|20420-6|LNC2000|Acid phosphatase.prostatic|Acid phosphatase.prostatic
C0803237|T201|COMP|1825-9|LNC2000|Alpha 1 antitrypsin|Alpha 1 antitrypsin
C0803238|T201|COMP|20423-0|LNC2000|Beta lactamase organism identified|Beta lactamase organism identified
C0803239|T201|COMP|20424-8|LNC2000|Cardiolipin Ab.IgG|Cardiolipin Ab.IgG
C0803240|T201|COMP|20425-5|LNC2000|Cardiolipin Ab.IgM|Cardiolipin Ab.IgM
C0803242|T201|COMP|20427-1|LNC2000|Acetylcholine receptor Ab|Acetylcholine receptor Ab
C0803251|T201|COMP|20436-2|LNC2000|Glucose^2H post dose glucose|Glucose^2H post dose glucose
C0803252|T201|COMP|20437-0|LNC2000|Glucose^3H post dose glucose|Glucose^3H post dose glucose
C0803253|T201|COMP|20438-8|LNC2000|Glucose^1H post dose glucose|Glucose^1H post dose glucose
C0803258|T201|COMP|20444-6|LNC2000|Herpes simplex virus 1+2 DNA|Herpes simplex virus 1+2 DNA
C0803260|T201|COMP|20446-1|LNC2000|Herpes simplex virus Ab.IgG|Herpes simplex virus Ab.IgG
C0803261|T201|COMP|20447-9|LNC2000|HIV 1 RNA|HIV 1 RNA
C0803262|T201|COMP|20448-7|LNC2000|Insulin|Insulin
C0803263|T201|COMP|20449-5|LNC2000|Borrelia burgdorferi Ab|Borrelia burgdorferi Ab
C0803264|T201|COMP|20450-3|LNC2000|Alpha-1-Fetoprotein|Alpha-1-Fetoprotein
C0803267|T201|COMP|20453-7|LNC2000|Epithelial cells|Epithelial cells
C0803268|T201|COMP|20454-5|LNC2000|Protein|Protein
C0803269|T201|COMP|20455-2|LNC2000|Leukocytes|Leukocytes
C0803270|T201|COMP|20456-0|LNC2000|Fungi.yeastlike|Fungi.yeastlike
C0803271|T201|COMP|20457-8|LNC2000|Fungi.filamentous|Fungi.filamentous
C0803272|T201|COMP|20458-6|LNC2000|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C0803274|T201|COMP|20460-2|LNC2000|Cefuroxime.oral|Cefuroxime.oral
C0803279|T201|COMP|20465-1|LNC2000|Choriogonadotropin|Choriogonadotropin
C0803280|T201|COMP|20466-9|LNC2000|Estriol.unconjugated|Estriol.unconjugated
C0803282|T201|COMP|20468-5|LNC2000|Thiamine|Thiamine
C0803283|T201|COMP|20469-3|LNC2000|Acetone|Acetone
C0803287|T201|COMP|20473-5|LNC2000|Polymorphonuclear cells|Polymorphonuclear cells
C0803288|T201|COMP|20474-3|LNC2000|Bacteria identified|Bacteria identified
C0803289|T201|COMP|20475-0|LNC2000|Cytomegalovirus Ab.IgG|Cytomegalovirus Ab.IgG
C0803293|T201|COMP|20479-2|LNC2000|Measles virus Ab.IgG|Measles virus Ab.IgG
C0803306|T201|COMP|20495-8|LNC2000|Gliadin Ab.IgA|Gliadin Ab.IgA
C0803307|T201|COMP|20496-6|LNC2000|Gliadin Ab.IgG|Gliadin Ab.IgG
C0803310|T201|COMP|20499-0|LNC2000|Phosphatidylglycerol/Surfactant.total|Phosphatidylglycerol/Surfactant.total
C0803316|T201|COMP|20505-4|LNC2000|Bilirubin|Bilirubin
C0803317|T201|COMP|20506-2|LNC2000|Specimen drawn from|Specimen drawn from
C0803318|T201|COMP|20507-0|LNC2000|Reagin Ab|Reagin Ab
C0803323|T201|COMP|20512-0|LNC2000|Turbidity|Turbidity
C0803324|T201|COMP|20513-8|LNC2000|Turbidity|Turbidity
C0803372|T201|COMP|20563-3|LNC2000|Carboxyhemoglobin/Hemoglobin.total|Carboxyhemoglobin/Hemoglobin.total
C0803374|T201|COMP|20565-8|LNC2000|Carbon dioxide|Carbon dioxide
C0803378|T201|COMP|20569-0|LNC2000|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C0803379|T201|COMP|20570-8|LNC2000|Hematocrit|Hematocrit
C0803382|T201|COMP|20573-2|LNC2000|Histoplasma capsulatum mycelial phase Ab|Histoplasma capsulatum mycelial phase Ab
C0803383|T201|COMP|20574-0|LNC2000|Histoplasma capsulatum yeast phase Ab|Histoplasma capsulatum yeast phase Ab
C0803387|T201|COMP|20578-1|LNC2000|Vancomycin|Vancomycin
C0803398|T201|COMP|20593-0|LNC2000|Cells.CD19/100 cells|Cells.CD19/100 cells
C0803429|T201|COMP|20624-3|LNC2000|Creatinine|Creatinine
C0803434|T201|COMP|20629-2|LNC2000|levoFLOXacin|levoFLOXacin
C0803440|T201|COMP|20636-7|LNC2000|Alanine|Alanine
C0803441|T201|COMP|20637-5|LNC2000|Arginine|Arginine
C0803442|T201|COMP|20638-3|LNC2000|Asparagine|Asparagine
C0803444|T201|COMP|20640-9|LNC2000|Citrulline|Citrulline
C0803447|T201|COMP|20643-3|LNC2000|Glutamine|Glutamine
C0803448|T201|COMP|20644-1|LNC2000|Glycine|Glycine
C0803449|T201|COMP|20645-8|LNC2000|Histidine|Histidine
C0803452|T201|COMP|20648-2|LNC2000|Isoleucine|Isoleucine
C0803453|T201|COMP|20649-0|LNC2000|Leucine|Leucine
C0803454|T201|COMP|20650-8|LNC2000|Lysine|Lysine
C0803455|T201|COMP|20651-6|LNC2000|Methionine|Methionine
C0803456|T201|COMP|20652-4|LNC2000|Ornithine|Ornithine
C0803458|T201|COMP|20655-7|LNC2000|Proline|Proline
C0803459|T201|COMP|20656-5|LNC2000|Serine|Serine
C0803460|T201|COMP|20657-3|LNC2000|Taurine|Taurine
C0803461|T201|COMP|20658-1|LNC2000|Threonine|Threonine
C0803463|T201|COMP|20660-7|LNC2000|Tyrosine|Tyrosine
C0803464|T201|COMP|20661-5|LNC2000|Valine|Valine
C0803561|T201|COMP|20761-3|LNC2000|Clostridioides difficile|Clostridioides difficile
C0803581|T201|COMP|20781-1|LNC2000|Cryptosporidium sp|Cryptosporidium sp
C0803789|T201|COMP|20991-6|LNC2000|Antithrombin|Antithrombin
C0803796|T201|COMP|20999-9|LNC2000|Cell fractions|Cell fractions
C0803797|T201|COMP|21000-5|LNC2000|Erythrocyte distribution width|Erythrocyte distribution width
C0803800|T201|COMP|21003-9|LNC2000|Fungus identified|Fungus identified
C0803816|T201|COMP|19050-4|LNC2000|Metanephrines|Metanephrines
C0803817|T201|COMP|21020-3|LNC2000|Bacteria identified|Bacteria identified
C0803820|T201|COMP|21023-7|LNC2000|Neutrophil cytoplasmic Ab|Neutrophil cytoplasmic Ab
C0803821|T201|COMP|21024-5|LNC2000|Pathologist interpretation|Pathologist interpretation
C0803823|T201|COMP|21026-0|LNC2000|Pathologist interpretation|Pathologist interpretation
C0803824|T201|COMP|21027-8|LNC2000|Platelet aggregation|Platelet aggregation
C0803828|T201|COMP|21032-8|LNC2000|Coagulation thrombin induced|Coagulation thrombin induced
C0803829|T201|COMP|21033-6|LNC2000|Yeast.budding|Yeast.budding
C0803902|T201|COMP|21108-6|LNC2000|Beta 2 glycoprotein 1 Ab.IgA|Beta 2 glycoprotein 1 Ab.IgA
C0803906|T201|COMP|21112-8|LNC2000|Birth date|Birth date
C0803971|T201|COMP|21654-9|LNC2000|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C0803984|T201|COMP|21190-4|LNC2000|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0803992|T201|COMP|21198-7|LNC2000|Choriogonadotropin.beta subunit|Choriogonadotropin.beta subunit
C0804054|T201|COMP|21260-5|LNC2000|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C0804056|T201|COMP|21262-1|LNC2000|Escherichia coli shiga-like toxin|Escherichia coli shiga-like toxin
C0804058|T201|COMP|21264-7|LNC2000|Estriol.unconjugated^^adjusted|Estriol.unconjugated^^adjusted
C0804159|T201|COMP|21365-2|LNC2000|Leptin|Leptin
C0804210|T201|COMP|21416-3|LNC2000|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C0804216|T201|COMP|21422-1|LNC2000|Normetanephrine|Normetanephrine
C0804235|T201|COMP|21441-1|LNC2000|Human papilloma virus 6+11+42+43+44 DNA|Human papilloma virus 6+11+42+43+44 DNA
C0804271|T201|COMP|6220-8|LNC2000|Solanum tuberosum Ab.IgE|Solanum tuberosum Ab.IgE
C0804276|T201|COMP|21482-5|LNC2000|Protein|Protein
C0804319|T201|COMP|21525-1|LNC2000|Sodium|Sodium
C0804343|T201|COMP|15761-0|LNC2000|Liquidambar styraciflua Ab.IgE.RAST class|Liquidambar styraciflua Ab.IgE.RAST class
C0804376|T201|COMP|21582-2|LNC2000|Tryptase|Tryptase
C0804405|T201|COMP|21612-7|LNC2000|Age|Age
C0804406|T201|COMP|21613-5|LNC2000|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C0804411|T201|COMP|21619-2|LNC2000|APOE gene targeted mutation analysis|APOE gene targeted mutation analysis
C0804457|T201|COMP|21667-1|LNC2000|F5 gene targeted mutation analysis|F5 gene targeted mutation analysis
C0804485|T201|COMP|21695-2|LNC2000|HFE gene.p.Cys282Tyr|HFE gene.p.Cys282Tyr
C0804499|T201|COMP|21709-1|LNC2000|MTHFR gene targeted mutation analysis|MTHFR gene targeted mutation analysis
C0804549|T201|COMP|21760-4|LNC2000|FRAXE gene.CGG repeats|FRAXE gene.CGG repeats
C0804609|T201|COMP|21821-4|LNC2000|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript|t(9;22)(q34.1;q11)(ABL1,BCR) fusion transcript
C0879657|T201|COMP|19734-3|LNC2000|Chicken droppings Ab.IgE|Chicken droppings Ab.IgE
C0879690|T201|COMP|22086-3|LNC2000|Aspergillus niger Ab|Aspergillus niger Ab
C0879709|T201|COMP|22110-1|LNC2000|Bartonella henselae Ab.IgG|Bartonella henselae Ab.IgG
C0879710|T201|COMP|22111-9|LNC2000|Bartonella henselae Ab.IgM|Bartonella henselae Ab.IgM
C0879728|T201|COMP|22131-7|LNC2000|Borrelia burgdorferi Ab.IgG+IgM|Borrelia burgdorferi Ab.IgG+IgM
C0879869|T201|COMP|22296-8|LNC2000|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C0879870|T201|COMP|22297-6|LNC2000|Epstein Barr virus nuclear Ab|Epstein Barr virus nuclear Ab
C0879883|T201|COMP|22310-7|LNC2000|Helicobacter pylori Ab|Helicobacter pylori Ab
C0879885|T201|COMP|22314-9|LNC2000|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C0879886|T201|COMP|22315-6|LNC2000|Hepatitis A virus Ab.IgM|Hepatitis A virus Ab.IgM
C0879891|T201|COMP|22322-2|LNC2000|Hepatitis B virus surface Ab|Hepatitis B virus surface Ab
C0879897|T201|COMP|22330-5|LNC2000|Hepatitis D virus Ab|Hepatitis D virus Ab
C0879925|T201|COMP|22362-8|LNC2000|HTLV I+II Ab|HTLV I+II Ab
C0879967|T201|COMP|22412-1|LNC2000|Saccharopolyspora rectivirgula Ab|Saccharopolyspora rectivirgula Ab
C0879970|T201|COMP|22415-4|LNC2000|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0880011|T201|COMP|22463-4|LNC2000|Reagin Ab|Reagin Ab
C0880042|T201|COMP|22496-4|LNC2000|Rubella virus Ab|Rubella virus Ab
C0880102|T201|COMP|22568-0|LNC2000|Streptolysin O Ab|Streptolysin O Ab
C0880118|T201|COMP|22587-0|LNC2000|Treponema pallidum Ab|Treponema pallidum Ab
C0880187|T201|COMP|20642-5|LNC2000|Glutamate|Glutamate
C0880263|T201|COMP|22763-7|LNC2000|Ammonia|Ammonia
C0880736|T201|COMP|23301-5|LNC2000|Mycoplasma sp DNA|Mycoplasma sp DNA
C0881021|T201|COMP|23641-4|LNC2000|Quinupristin+Dalfopristin|Quinupristin+Dalfopristin
C0881037|T201|COMP|23658-8|LNC2000|Antibiotic XXX|Antibiotic XXX
C0881125|T201|COMP|23761-0|LNC2000|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0881171|T201|COMP|23811-3|LNC2000|Alpha-1-Fetoprotein^^adjusted|Alpha-1-Fetoprotein^^adjusted
C0881199|T201|COMP|23841-0|LNC2000|Choriogonadotropin.beta subunit^^adjusted|Choriogonadotropin.beta subunit^^adjusted
C0881213|T201|COMP|23860-0|LNC2000|Erythrocytes|Erythrocytes
C0881221|T201|COMP|23870-9|LNC2000|Hepatitis C virus 100+5-1-1 Ab|Hepatitis C virus 100+5-1-1 Ab
C0881222|T201|COMP|23871-7|LNC2000|Hepatitis C virus NS5 Ab|Hepatitis C virus NS5 Ab
C0881226|T201|COMP|23876-6|LNC2000|HIV 1 RNA|HIV 1 RNA
C0881227|T201|COMP|23877-4|LNC2000|Anaplasma phagocytophilum Ab.IgG|Anaplasma phagocytophilum Ab.IgG
C0881228|T201|COMP|23878-2|LNC2000|Anaplasma phagocytophilum Ab.IgM|Anaplasma phagocytophilum Ab.IgM
C0881233|T201|COMP|23883-2|LNC2000|Inhibin A|Inhibin A
C0881253|T201|COMP|23905-3|LNC2000|Mycophenolate|Mycophenolate
C0881343|T201|COMP|24012-7|LNC2000|HIV 1 Ag|HIV 1 Ag
C0881344|T201|COMP|24013-5|LNC2000|HIV 1 RNA|HIV 1 RNA
C0881346|T201|COMP|24015-0|LNC2000|Influenza virus A+B Ag|Influenza virus A+B Ag
C0881426|T201|COMP|24111-7|LNC2000|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C0881427|T201|COMP|24113-3|LNC2000|Hepatitis B virus core Ab.IgM|Hepatitis B virus core Ab.IgM
C0881428|T201|COMP|24114-1|LNC2000|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C0881429|T201|COMP|24115-8|LNC2000|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C0881432|T201|COMP|24119-0|LNC2000|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C0881438|T201|COMP|24125-7|LNC2000|Androgen.free index|Androgen.free index
C0881452|T201|COMP|24139-8|LNC2000|Blatella germanica Ab.IgG|Blatella germanica Ab.IgG
C0881468|T201|COMP|6164-8|LNC2000|Quercus virginiana Ab.IgE|Quercus virginiana Ab.IgE
C0881590|T201|COMP|24312-1|LNC2000|Treponema pallidum Ab|Treponema pallidum Ab
C0881644|T201|COMP|24378-2|LNC2000|Platelet aggregation.EPINEPHrine induced|Platelet aggregation.EPINEPHrine induced
C0881717|T201|COMP|24467-3|LNC2000|Cells.CD3+CD4+|Cells.CD3+CD4+
C0881719|T201|COMP|24469-9|LNC2000|Hemoglobin XXX/Hemoglobin.total|Hemoglobin XXX/Hemoglobin.total
C0881724|T201|COMP|24475-6|LNC2000|F2 gene.c.20210G>A|F2 gene.c.20210G>A
C0881725|T201|COMP|24476-4|LNC2000|F2 gene targeted mutation analysis|F2 gene targeted mutation analysis
C0882250|T201|COMP|22203-4|LNC2000|Clostridium tetani Ab.IgG|Clostridium tetani Ab.IgG
C0882468|T201|COMP|24103-4|LNC2000|Plasma cells|Plasma cells
C0882469|T201|COMP|24108-3|LNC2000|Cancer Ag 19-9|Cancer Ag 19-9
C0884314|T201|COMP|24011-9|LNC2000|Hepatitis C virus Ab band pattern|Hepatitis C virus Ab band pattern
C0941344|T201|COMP|25145-4|LNC2000|Bacteria|Bacteria
C0941346|T201|COMP|25148-8|LNC2000|Calcium oxalate crystals|Calcium oxalate crystals
C0941347|T201|COMP|25149-6|LNC2000|Calcium phosphate crystals|Calcium phosphate crystals
C0941350|T201|COMP|25154-6|LNC2000|Crystals.unidentified|Crystals.unidentified
C0941352|T201|COMP|25157-9|LNC2000|Epithelial casts|Epithelial casts
C0941353|T201|COMP|25158-7|LNC2000|Oval fat bodies (globules)|Oval fat bodies (globules)
C0941355|T201|COMP|25160-3|LNC2000|Granular casts|Granular casts
C0941357|T201|COMP|25162-9|LNC2000|Hyaline casts|Hyaline casts
C0941533|T201|COMP|25383-1|LNC2000|Cow milk Ab.IgE.RAST class|Cow milk Ab.IgE.RAST class
C0941565|T201|COMP|25418-5|LNC2000|Mumps virus Ab.IgG|Mumps virus Ab.IgG
C0941572|T201|COMP|25428-4|LNC2000|Glucose|Glucose
C0941609|T201|COMP|25473-0|LNC2000|Metanephrine|Metanephrine
C0941610|T201|COMP|25474-8|LNC2000|Metanephrines|Metanephrines
C0941622|T201|COMP|25489-6|LNC2000|Normetanephrine|Normetanephrine
C0941729|T201|COMP|25630-5|LNC2000|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0941730|T201|COMP|25631-3|LNC2000|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C0941788|T201|COMP|25700-6|LNC2000|Interpretation|Interpretation
C0941896|T201|COMP|25836-8|LNC2000|HIV 1 RNA|HIV 1 RNA
C0942025|T201|COMP|25987-9|LNC2000|Testosterone.free|Testosterone.free
C0942070|T201|COMP|26043-0|LNC2000|HLA-B27|HLA-B27
C0942079|T201|COMP|26052-1|LNC2000|Epithelial cells.renal|Epithelial cells.renal
C0942414|T201|COMP|26444-0|LNC2000|Basophils|Basophils
C0942416|T201|COMP|26446-5|LNC2000|Blasts/100 leukocytes|Blasts/100 leukocytes
C0942417|T201|COMP|26447-3|LNC2000|Blasts/100 leukocytes|Blasts/100 leukocytes
C0942419|T201|COMP|26449-9|LNC2000|Eosinophils|Eosinophils
C0942420|T201|COMP|26451-5|LNC2000|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0942421|T201|COMP|26452-3|LNC2000|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0942423|T201|COMP|26454-9|LNC2000|Erythrocytes|Erythrocytes
C0942426|T201|COMP|26458-0|LNC2000|Erythrocytes|Erythrocytes
C0942431|T201|COMP|26466-3|LNC2000|Leukocytes|Leukocytes
C0942435|T201|COMP|26472-1|LNC2000|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0942436|T201|COMP|26473-9|LNC2000|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0942437|T201|COMP|26474-7|LNC2000|Lymphocytes|Lymphocytes
C0942440|T201|COMP|26478-8|LNC2000|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0942441|T201|COMP|26479-6|LNC2000|Lymphocytes/100 leukocytes|Lymphocytes/100 leukocytes
C0942446|T201|COMP|26484-6|LNC2000|Monocytes|Monocytes
C0942447|T201|COMP|26485-3|LNC2000|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0942448|T201|COMP|26486-1|LNC2000|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0942449|T201|COMP|26487-9|LNC2000|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C0942460|T201|COMP|26498-6|LNC2000|Myelocytes/100 leukocytes|Myelocytes/100 leukocytes
C0942461|T201|COMP|26499-4|LNC2000|Neutrophils|Neutrophils
C0942468|T201|COMP|26508-2|LNC2000|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0942469|T201|COMP|26509-0|LNC2000|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0942470|T201|COMP|26510-8|LNC2000|Neutrophils.band form/100 leukocytes|Neutrophils.band form/100 leukocytes
C0942471|T201|COMP|26511-6|LNC2000|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0942474|T201|COMP|26515-7|LNC2000|Platelets|Platelets
C0942476|T201|COMP|26518-1|LNC2000|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0942480|T201|COMP|26523-1|LNC2000|Promyelocytes|Promyelocytes
C0942484|T201|COMP|26528-0|LNC2000|Cortisol^1H post dose corticotropin|Cortisol^1H post dose corticotropin
C0942486|T201|COMP|26530-6|LNC2000|Cortisol^30M post dose corticotropin|Cortisol^30M post dose corticotropin
C0942549|T201|COMP|26607-2|LNC2000|Cystathionine|Cystathionine
C0942903|T201|COMP|27038-9|LNC2000|Endomysium Ab.IgA|Endomysium Ab.IgA
C0942931|T201|COMP|27071-0|LNC2000|Cells.CD45|Cells.CD45
C0943037|T201|COMP|27200-5|LNC2000|Nuclear Ab|Nuclear Ab
C0943165|T201|COMP|27353-2|LNC2000|Estimated average glucose|Estimated average glucose
C0943215|T201|COMP|27416-7|LNC2000|SCL-70 extractable nuclear Ab|SCL-70 extractable nuclear Ab
C0943506|T201|COMP|27811-9|LNC2000|Antithrombin actual/Normal|Antithrombin actual/Normal
C0943511|T201|COMP|27816-8|LNC2000|von Willebrand factor Ag actual/Normal|von Willebrand factor Ag actual/Normal
C0943513|T201|COMP|27818-4|LNC2000|Protein C actual/Normal|Protein C actual/Normal
C0943514|T201|COMP|27819-2|LNC2000|Protein C actual/Normal|Protein C actual/Normal
C0943515|T201|COMP|27820-0|LNC2000|Protein C Ag actual/Normal|Protein C Ag actual/Normal
C0943516|T201|COMP|27821-8|LNC2000|Protein S.free Ag actual/Normal|Protein S.free Ag actual/Normal
C0943517|T201|COMP|27823-4|LNC2000|Protein S Ag actual/Normal|Protein S Ag actual/Normal
C0943603|T201|COMP|27923-2|LNC2000|Ubiquinone 10|Ubiquinone 10
C0943616|T201|COMP|27939-8|LNC2000|Collagen crosslinked N-telopeptide|Collagen crosslinked N-telopeptide
C0943622|T201|COMP|27948-9|LNC2000|Herpes simplex virus 1+2 Ab.IgG|Herpes simplex virus 1+2 Ab.IgG
C0943672|T201|COMP|28005-7|LNC2000|MTHFR gene.c.677C>T|MTHFR gene.c.677C>T
C0943674|T201|COMP|28009-9|LNC2000|Specimen volume|Specimen volume
C0944135|T201|COMP|28541-1|LNC2000|Metamyelocytes/100 leukocytes|Metamyelocytes/100 leukocytes
C0944137|T201|COMP|28543-7|LNC2000|Basophils/100 leukocytes|Basophils/100 leukocytes
C0944138|T201|COMP|28545-2|LNC2000|Mucus|Mucus
C0944218|T201|COMP|28637-7|LNC2000|Base deficit|Base deficit
C0944221|T201|COMP|28640-1|LNC2000|Bicarbonate|Bicarbonate
C0944222|T201|COMP|28641-9|LNC2000|Bicarbonate|Bicarbonate
C0944223|T201|COMP|28642-7|LNC2000|Oxygen saturation|Oxygen saturation
C0944224|T201|COMP|28644-3|LNC2000|Carbon dioxide|Carbon dioxide
C0944225|T201|COMP|28645-0|LNC2000|Carbon dioxide|Carbon dioxide
C0944227|T201|COMP|28648-4|LNC2000|Oxygen|Oxygen
C0944729|T201|COMP|29247-4|LNC2000|Sirolimus|Sirolimus
C0944746|T201|COMP|29265-6|LNC2000|Calcium^^corrected for albumin|Calcium^^corrected for albumin
C0944759|T201|COMP|29280-5|LNC2000|Fibrin D-dimer|Fibrin D-dimer
C0944978|T201|COMP|29541-0|LNC2000|HIV 1 RNA|HIV 1 RNA
C0944993|T201|COMP|29559-2|LNC2000|Haemophilus ducreyi DNA|Haemophilus ducreyi DNA
C0945005|T201|COMP|29571-7|LNC2000|Phenylalanine|Phenylalanine
C0945007|T201|COMP|29573-3|LNC2000|Phenylalanine|Phenylalanine
C0945008|T201|COMP|29574-1|LNC2000|Thyrotropin|Thyrotropin
C0945009|T201|COMP|29575-8|LNC2000|Thyrotropin|Thyrotropin
C0945022|T201|COMP|29591-5|LNC2000|Enterovirus RNA|Enterovirus RNA
C0945041|T201|COMP|29615-2|LNC2000|Hepatitis B virus DNA|Hepatitis B virus DNA
C0945063|T201|COMP|29641-8|LNC2000|Neutrophil cytoplasmic Ab.atypical|Neutrophil cytoplasmic Ab.atypical
C0945079|T201|COMP|29660-8|LNC2000|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0945089|T201|COMP|29675-6|LNC2000|Parvovirus B19 Ab.IgG|Parvovirus B19 Ab.IgG
C0945181|T201|COMP|25147-0|LNC2000|Calcium carbonate crystals|Calcium carbonate crystals
C0945182|T201|COMP|25156-1|LNC2000|Eosinophils|Eosinophils
C0945223|T201|COMP|25435-9|LNC2000|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C0945272|T201|COMP|25835-0|LNC2000|HIV 1 RNA|HIV 1 RNA
C0945354|T201|COMP|26450-7|LNC2000|Eosinophils/100 leukocytes|Eosinophils/100 leukocytes
C0945355|T201|COMP|26455-6|LNC2000|Erythrocytes|Erythrocytes
C0945357|T201|COMP|26464-8|LNC2000|Leukocytes|Leukocytes
C0945359|T201|COMP|26471-3|LNC2000|Leukocytes other/100 leukocytes|Leukocytes other/100 leukocytes
C0945362|T201|COMP|26507-4|LNC2000|Neutrophils.band form|Neutrophils.band form
C0945363|T201|COMP|26512-4|LNC2000|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C0945364|T201|COMP|26517-3|LNC2000|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C0945400|T201|COMP|26760-9|LNC2000|Cannabinoids|Cannabinoids
C0945429|T201|COMP|26927-4|LNC2000|Herpes simplex virus 2 Ab.IgM|Herpes simplex virus 2 Ab.IgM
C0945446|T201|COMP|27045-4|LNC2000|Microscopic exam|Microscopic exam
C0945541|T201|COMP|27822-6|LNC2000|Protein S actual/Normal|Protein S actual/Normal
C0945637|T201|COMP|28643-5|LNC2000|Oxygen saturation|Oxygen saturation
C0945639|T201|COMP|28649-2|LNC2000|Oxygen|Oxygen
C0945742|T201|COMP|29374-6|LNC2000|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C0945763|T201|COMP|29539-4|LNC2000|HIV 1 RNA|HIV 1 RNA
C0947260|T201|COMP|28008-1|LNC2000|Cytomegalovirus DNA|Cytomegalovirus DNA
C0947495|T201|COMP|14251-3|LNC2000|Mitochondria M2 Ab.IgG|Mitochondria M2 Ab.IgG
C1113710|T201|COMP|29770-5|LNC2000|Karyotype|Karyotype
C1113711|T201|COMP|29771-3|LNC2000|Hemoglobin.gastrointestinal.lower|Hemoglobin.gastrointestinal.lower
C1113816|T201|COMP|29891-9|LNC2000|Carbon dioxide^post dose urea|Carbon dioxide^post dose urea
C1113818|T201|COMP|29893-5|LNC2000|HIV 1 Ab|HIV 1 Ab
C1113826|T201|COMP|29901-6|LNC2000|HTLV I+II Ab|HTLV I+II Ab
C1113883|T201|COMP|29967-7|LNC2000|Neutrophil cytoplasmic Ab.IgG|Neutrophil cytoplasmic Ab.IgG
C1113913|T201|COMP|30003-8|LNC2000|Albumin|Albumin
C1113982|T201|COMP|30083-0|LNC2000|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C1113987|T201|COMP|30089-7|LNC2000|Transitional cells|Transitional cells
C1113995|T201|COMP|30099-6|LNC2000|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C1114052|T201|COMP|30165-5|LNC2000|Phosphatidylcholine/Albumin|Phosphatidylcholine/Albumin
C1114053|T201|COMP|30166-3|LNC2000|Thyroid stimulating immunoglobulins actual/Normal|Thyroid stimulating immunoglobulins actual/Normal
C1114056|T201|COMP|30170-5|LNC2000|Periplaneta americana Ab.IgE|Periplaneta americana Ab.IgE
C1114065|T201|COMP|30180-4|LNC2000|Basophils/100 leukocytes|Basophils/100 leukocytes
C1114078|T201|COMP|30193-7|LNC2000|Acylcarnitine/Carnitine.free (C0)|Acylcarnitine/Carnitine.free (C0)
C1114121|T201|COMP|30243-0|LNC2000|Choriogonadotropin.intact|Choriogonadotropin.intact
C1114125|T201|COMP|30247-1|LNC2000|Cytomegalovirus DNA|Cytomegalovirus DNA
C1114184|T201|COMP|30313-1|LNC2000|Hemoglobin|Hemoglobin
C1114188|T201|COMP|30318-0|LNC2000|Base deficit|Base deficit
C1114205|T201|COMP|30339-6|LNC2000|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C1114206|T201|COMP|30340-4|LNC2000|Epstein Barr virus capsid Ab.IgM|Epstein Barr virus capsid Ab.IgM
C1114213|T201|COMP|30350-3|LNC2000|Hemoglobin|Hemoglobin
C1114223|T201|COMP|30361-0|LNC2000|HIV 2 Ab|HIV 2 Ab
C1114236|T201|COMP|30374-3|LNC2000|Basophils/100 leukocytes|Basophils/100 leukocytes
C1114238|T201|COMP|30376-8|LNC2000|Blasts|Blasts
C1114261|T201|COMP|30405-5|LNC2000|Leukocytes|Leukocytes
C1114280|T201|COMP|30427-9|LNC2000|Macrophages/100 leukocytes|Macrophages/100 leukocytes
C1114281|T201|COMP|30428-7|LNC2000|Erythrocyte mean corpuscular volume|Erythrocyte mean corpuscular volume
C1114290|T201|COMP|30437-8|LNC2000|Monocytes+Macrophages/100 leukocytes|Monocytes+Macrophages/100 leukocytes
C1114307|T201|COMP|30457-6|LNC2000|Nonhematic cells/100 leukocytes|Nonhematic cells/100 leukocytes
C1114318|T201|COMP|30471-7|LNC2000|levETIRAcetam|levETIRAcetam
C1114363|T201|COMP|30522-7|LNC2000|C reactive protein|C reactive protein
C1114365|T201|COMP|30525-0|LNC2000|Age|Age
C1114721|T201|COMP|30934-4|LNC2000|Natriuretic peptide.B|Natriuretic peptide.B
C1114799|T201|COMP|31017-7|LNC2000|Tissue transglutaminase Ab.IgA|Tissue transglutaminase Ab.IgA
C1114801|T201|COMP|31019-3|LNC2000|10-Hydroxycarbazepine|10-Hydroxycarbazepine
C1114812|T201|COMP|31032-6|LNC2000|Saccharomyces cerevisiae Ab.IgA|Saccharomyces cerevisiae Ab.IgA
C1114815|T201|COMP|31036-7|LNC2000|Gatifloxacin|Gatifloxacin
C1114843|T201|COMP|29953-7|LNC2000|Nuclear Ab|Nuclear Ab
C1114891|T201|COMP|30341-2|LNC2000|Erythrocyte sedimentation rate|Erythrocyte sedimentation rate
C1114897|T201|COMP|30394-1|LNC2000|Granulocytes|Granulocytes
C1114903|T201|COMP|30446-9|LNC2000|Myelocytes|Myelocytes
C1114906|T201|COMP|26524-9|LNC2000|Promyelocytes/100 leukocytes|Promyelocytes/100 leukocytes
C1145645|T201|COMP|2703-7|LNC2000|Oxygen|Oxygen
C1145647|T201|COMP|2705-2|LNC2000|Oxygen|Oxygen
C1145649|T201|COMP|6584-7|LNC2000|Virus identified|Virus identified
C1145650|T201|COMP|580-1|LNC2000|Fungus identified|Fungus identified
C1145656|T201|COMP|625-4|LNC2000|Bacteria identified|Bacteria identified
C1145716|T201|COMP|12195-4|LNC2000|Creatinine renal clearance/1.73 sq M|Creatinine renal clearance/1.73 sq M
C1145717|T201|COMP|17948-1|LNC2000|Fungus identified^^^3|Fungus identified^^^3
C1145718|T201|COMP|17947-3|LNC2000|Fungus identified^^^2|Fungus identified^^^2
C1145723|T201|COMP|10352-3|LNC2000|Bacteria identified|Bacteria identified
C1145728|T201|COMP|10353-1|LNC2000|Bacteria identified|Bacteria identified
C1146765|T201|COMP|31080-5|LNC2000|Cannabinoids|Cannabinoids
C1146785|T201|COMP|31100-1|LNC2000|Hematocrit|Hematocrit
C1146787|T201|COMP|31102-7|LNC2000|Protein S actual/Normal|Protein S actual/Normal
C1146797|T201|COMP|31112-6|LNC2000|Reticulocytes/100 erythrocytes|Reticulocytes/100 erythrocytes
C1146829|T201|COMP|31144-9|LNC2000|Thyroxine|Thyroxine
C1146832|T201|COMP|31147-2|LNC2000|Reagin Ab|Reagin Ab
C1146841|T201|COMP|31156-3|LNC2000|Hemoglobin Barts/Hemoglobin.total|Hemoglobin Barts/Hemoglobin.total
C1146845|T201|COMP|31160-5|LNC2000|Polymorphonuclear cells/100 leukocytes|Polymorphonuclear cells/100 leukocytes
C1146886|T201|COMP|31201-7|LNC2000|HIV 1+2 Ab|HIV 1+2 Ab
C1146889|T201|COMP|31204-1|LNC2000|Hepatitis B virus core Ab.IgM|Hepatitis B virus core Ab.IgM
C1146893|T201|COMP|31208-2|LNC2000|Specimen source|Specimen source
C1146894|T201|COMP|31209-0|LNC2000|Islet cell 512 Ab|Islet cell 512 Ab
C1147059|T201|COMP|31374-2|LNC2000|Epstein Barr virus nuclear Ab.IgG|Epstein Barr virus nuclear Ab.IgG
C1147103|T201|COMP|31418-7|LNC2000|Heterophile Ab|Heterophile Ab
C1147472|T201|COMP|31788-3|LNC2000|Cryptococcus sp Ag|Cryptococcus sp Ag
C1147481|T201|COMP|31797-4|LNC2000|Cytomegalovirus Ag|Cytomegalovirus Ag
C1147527|T201|COMP|31843-6|LNC2000|Helicobacter pylori Ag|Helicobacter pylori Ag
C1147528|T201|COMP|31844-4|LNC2000|Hepatitis B virus little e Ag|Hepatitis B virus little e Ag
C1147715|T201|COMP|32031-7|LNC2000|Phosphatidylserine Ab.IgA|Phosphatidylserine Ab.IgA
C1147716|T201|COMP|32032-5|LNC2000|Phosphatidylserine Ab.IgG|Phosphatidylserine Ab.IgG
C1147717|T201|COMP|32033-3|LNC2000|Phosphatidylserine Ab.IgM|Phosphatidylserine Ab.IgM
C1147730|T201|COMP|32046-5|LNC2000|Pregnancy associated plasma protein A|Pregnancy associated plasma protein A
C1147817|T201|COMP|32133-1|LNC2000|Lactate|Lactate
C1147824|T201|COMP|32140-6|LNC2000|Hemoglobin F|Hemoglobin F
C1147830|T201|COMP|32146-3|LNC2000|Platelets.large|Platelets.large
C1147831|T201|COMP|32147-1|LNC2000|Reducing substances|Reducing substances
C1147848|T201|COMP|32164-6|LNC2000|Cells|Cells
C1147850|T201|COMP|32166-1|LNC2000|Choriogonadotropin^^adjusted|Choriogonadotropin^^adjusted
C1147851|T201|COMP|32167-9|LNC2000|Clarity|Clarity
C1147882|T201|COMP|32198-4|LNC2000|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1147891|T201|COMP|32207-3|LNC2000|Platelet distribution width|Platelet distribution width
C1147899|T201|COMP|32215-6|LNC2000|Thyroxine free index|Thyroxine free index
C1147901|T201|COMP|32217-2|LNC2000|von Willebrand factor multimers|von Willebrand factor multimers
C1147902|T201|COMP|32218-0|LNC2000|Cyclic citrullinated peptide Ab|Cyclic citrullinated peptide Ab
C1147904|T201|COMP|32220-6|LNC2000|Liver kidney microsomal 1 Ab|Liver kidney microsomal 1 Ab
C1147968|T201|COMP|32284-2|LNC2000|BK virus DNA|BK virus DNA
C1147970|T201|COMP|32286-7|LNC2000|Hepatitis C virus genotype|Hepatitis C virus genotype
C1148040|T201|COMP|32356-8|LNC2000|Yeast|Yeast
C1148199|T201|COMP|32515-9|LNC2000|Cells.CD3+CD4+|Cells.CD3+CD4+
C1148230|T201|COMP|32546-4|LNC2000|Glucose-6-Phosphate dehydrogenase|Glucose-6-Phosphate dehydrogenase
C1148238|T201|COMP|32554-8|LNC2000|Thiamine|Thiamine
C1148269|T201|COMP|32585-2|LNC2000|Epstein Barr virus DNA|Epstein Barr virus DNA
C1153739|T201|COMP|19049-6|LNC2000|Metanephrine|Metanephrine
C1315106|T201|COMP|32632-2|LNC2000|HEXA gene targeted mutation analysis|HEXA gene targeted mutation analysis
C1315111|T201|COMP|32637-1|LNC2000|Urease|Urease
C1315147|T201|COMP|32673-6|LNC2000|Creatine kinase.MB|Creatine kinase.MB
C1315154|T201|COMP|32680-1|LNC2000|Granular casts.fine|Granular casts.fine
C1315166|T201|COMP|32693-4|LNC2000|Lactate|Lactate
C1315177|T201|COMP|32705-6|LNC2000|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C1315182|T201|COMP|32623-1|LNC2000|Platelet mean volume|Platelet mean volume
C1315235|T201|COMP|32764-3|LNC2000|Clue cells|Clue cells
C1315236|T201|COMP|32765-0|LNC2000|Yeast|Yeast
C1315237|T201|COMP|32766-8|LNC2000|Trichomonas vaginalis|Trichomonas vaginalis
C1315257|T201|COMP|32786-6|LNC2000|Thyroperoxidase Ab|Thyroperoxidase Ab
C1315258|T201|COMP|32787-4|LNC2000|Neutrophil cytoplasmic Ab.perinuclear|Neutrophil cytoplasmic Ab.perinuclear
C1315260|T201|COMP|32789-0|LNC2000|Viscosity|Viscosity
C1315325|T201|COMP|32854-2|LNC2000|17-Hydroxyprogesterone|17-Hydroxyprogesterone
C1315469|T201|COMP|32998-7|LNC2000|Tissue transglutaminase Ab.IgG|Tissue transglutaminase Ab.IgG
C1315477|T201|COMP|33006-8|LNC2000|Cytomegalovirus DNA|Cytomegalovirus DNA
C1315508|T201|COMP|33037-3|LNC2000|Anion gap|Anion gap
C1315522|T201|COMP|33051-4|LNC2000|Erythrocytes|Erythrocytes
C1315686|T201|COMP|33215-5|LNC2000|Neutrophils.agranular|Neutrophils.agranular
C1315687|T201|COMP|33216-3|LNC2000|Platelets.agranular|Platelets.agranular
C1315688|T201|COMP|33217-1|LNC2000|Spermatozoa.agglutinated|Spermatozoa.agglutinated
C1315713|T201|COMP|33242-9|LNC2000|Fungi.filamentous|Fungi.filamentous
C1315718|T201|COMP|33247-8|LNC2000|Specimen weight|Specimen weight
C1315719|T201|COMP|33248-6|LNC2000|Diabetes status|Diabetes status
C1315723|T201|COMP|33254-4|LNC2000|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1315724|T201|COMP|33255-1|LNC2000|Cell fractions|Cell fractions
C1315725|T201|COMP|33256-9|LNC2000|Leukocytes^^corrected for nucleated erythrocytes|Leukocytes^^corrected for nucleated erythrocytes
C1315757|T201|COMP|33288-2|LNC2000|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C1315801|T201|COMP|33332-8|LNC2000|Linezolid|Linezolid
C1315802|T201|COMP|33333-6|LNC2000|Colistin|Colistin
C1315827|T201|COMP|33358-3|LNC2000|Protein.monoclonal|Protein.monoclonal
C1315862|T201|COMP|33393-0|LNC2000|Granular casts.coarse|Granular casts.coarse
C1316005|T201|COMP|33536-4|LNC2000|Allergen.miscellaneous Ab.IgE.RAST class|Allergen.miscellaneous Ab.IgE.RAST class
C1316038|T201|COMP|33569-5|LNC2000|Sjogrens syndrome-A extractable nuclear Ab|Sjogrens syndrome-A extractable nuclear Ab
C1316060|T201|COMP|33593-5|LNC2000|Hemoglobin G-Coushatta/Hemoglobin.total|Hemoglobin G-Coushatta/Hemoglobin.total
C1316061|T201|COMP|33594-3|LNC2000|Platelet factor 4|Platelet factor 4
C1316094|T201|COMP|33630-5|LNC2000|HIV protease gene mutations detected|HIV protease gene mutations detected
C1316111|T201|COMP|33647-9|LNC2000|Protein.monoclonal/Protein.total|Protein.monoclonal/Protein.total
C1316182|T201|COMP|33718-8|LNC2000|Cytology report|Cytology report
C1316185|T201|COMP|33721-2|LNC2000|Pathology biopsy report|Pathology biopsy report
C1316226|T201|COMP|33762-6|LNC2000|Natriuretic peptide.B prohormone N-Terminal|Natriuretic peptide.B prohormone N-Terminal
C1316232|T201|COMP|33768-3|LNC2000|Leukocyte clumps|Leukocyte clumps
C1316237|T201|COMP|33773-3|LNC2000|Karyotype|Karyotype
C1316268|T201|COMP|33804-6|LNC2000|Erythrocyte casts|Erythrocyte casts
C1316356|T201|COMP|33893-9|LNC2000|Karyotype|Karyotype
C1316366|T201|COMP|33903-6|LNC2000|Ketones|Ketones
C1316368|T201|COMP|33905-1|LNC2000|Trichomonas sp|Trichomonas sp
C1316373|T201|COMP|33910-1|LNC2000|Rheumatoid factor|Rheumatoid factor
C1316377|T201|COMP|33914-3|LNC2000|Glomerular filtration rate/1.73 sq M.predicted|Glomerular filtration rate/1.73 sq M.predicted
C1316378|T201|COMP|33915-0|LNC2000|Anabasine|Anabasine
C1316380|T201|COMP|33917-6|LNC2000|Nornicotine|Nornicotine
C1316398|T201|COMP|33935-8|LNC2000|Cyclic citrullinated peptide Ab.IgG|Cyclic citrullinated peptide Ab.IgG
C1316407|T201|COMP|33944-0|LNC2000|Immunoglobulin light chains.lambda.free|Immunoglobulin light chains.lambda.free
C1316447|T201|COMP|33984-6|LNC2000|Coagulation factor X activity actual/Normal|Coagulation factor X activity actual/Normal
C1316611|T201|COMP|34148-7|LNC2000|Borrelia burgdorferi Ab.IgG+IgM|Borrelia burgdorferi Ab.IgG+IgM
C1316628|T201|COMP|34165-1|LNC2000|Granulocytes.immature|Granulocytes.immature
C1316903|T201|COMP|34441-6|LNC2000|Spermatozoa|Spermatozoa
C1316930|T201|COMP|34468-9|LNC2000|Clostridioides difficile toxin A+B|Clostridioides difficile toxin A+B
C1316981|T201|COMP|34519-9|LNC2000|HFE gene targeted mutation analysis|HFE gene targeted mutation analysis
C1316986|T201|COMP|34524-9|LNC2000|Neutrophils.band form|Neutrophils.band form
C1317032|T201|COMP|34571-0|LNC2000|Coagulation surface induced.lupus sensitive|Coagulation surface induced.lupus sensitive
C1369526|T201|COMP|34660-1|LNC2000|Hemoglobin A2/Hemoglobin.total|Hemoglobin A2/Hemoglobin.total
C1369527|T201|COMP|34661-9|LNC2000|Actin Ab.IgG|Actin Ab.IgG
C1369562|T201|COMP|34696-5|LNC2000|Collection method|Collection method
C1369567|T201|COMP|34701-3|LNC2000|Platelet factor 4 heparin complex induced Ab|Platelet factor 4 heparin complex induced Ab
C1369578|T201|COMP|34712-0|LNC2000|Clostridioides difficile|Clostridioides difficile
C1369579|T201|COMP|34713-8|LNC2000|Clostridioides difficile toxin A+B|Clostridioides difficile toxin A+B
C1369580|T201|COMP|34714-6|LNC2000|Coagulation tissue factor induced.INR|Coagulation tissue factor induced.INR
C1369847|T201|COMP|34985-2|LNC2000|Unidentified cells/100 leukocytes|Unidentified cells/100 leukocytes
C1369914|T201|COMP|35125-4|LNC2000|Hemoglobin Lepore/Hemoglobin.total|Hemoglobin Lepore/Hemoglobin.total
C1369915|T201|COMP|35126-2|LNC2000|Hemoglobin O-Arab/Hemoglobin.total|Hemoglobin O-Arab/Hemoglobin.total
C1369916|T201|COMP|35127-0|LNC2000|Hemoglobin A2.prime/Hemoglobin.total|Hemoglobin A2.prime/Hemoglobin.total
C1369982|T201|COMP|1974-5|LNC2000|Bilirubin|Bilirubin
C1370010|T201|COMP|2777-1|LNC2000|Phosphate|Phosphate
C1370059|T201|COMP|35270-8|LNC2000|Candida sp Ab|Candida sp Ab
C1370064|T201|COMP|35275-7|LNC2000|Measles virus Ab.IgG|Measles virus Ab.IgG
C1378285|T201|COMP|35051-2|LNC2000|Leukocytes other|Leukocytes other
C1507400|T201|COMP|35622-0|LNC2000|Nordiazepam|Nordiazepam
C1507465|T201|COMP|35331-8|LNC2000|OXcarbazepine|OXcarbazepine
C1507499|T201|COMP|35365-6|LNC2000|Vitamin D+Metabolites|Vitamin D+Metabolites
C1507517|T201|COMP|35383-9|LNC2000|Galactomannan Ag|Galactomannan Ag
C1507586|T201|COMP|35452-2|LNC2000|HIV 1 gp40 Ab|HIV 1 gp40 Ab
C1507626|T201|COMP|35492-8|LNC2000|Staphylococcus aureus.methicillin resistant DNA|Staphylococcus aureus.methicillin resistant DNA
C1507698|T201|COMP|35538-8|LNC2000|Saccharomyces cerevisiae Ab.IgG|Saccharomyces cerevisiae Ab.IgG
C1507731|T201|COMP|35571-9|LNC2000|Tyrosine|Tyrosine
C1507732|T201|COMP|35572-7|LNC2000|Phenylalanine/Tyrosine|Phenylalanine/Tyrosine
C1507751|T201|COMP|35591-7|LNC2000|Creatinine renal clearance.predicted|Creatinine renal clearance.predicted
C1507755|T201|COMP|35595-8|LNC2000|Acetaminophen|Acetaminophen
C1507757|T201|COMP|35597-4|LNC2000|Salicylates|Salicylates
C1507763|T201|COMP|35603-0|LNC2000|clonazePAM|clonazePAM
C1507814|T201|COMP|35663-4|LNC2000|Protein|Protein
C1507819|T201|COMP|35668-3|LNC2000|Gentamicin|Gentamicin
C1507821|T201|COMP|35670-9|LNC2000|Tobramycin|Tobramycin
C1507825|T201|COMP|35674-1|LNC2000|Creatinine|Creatinine
C1507826|T201|COMP|35675-8|LNC2000|Calcium|Calcium
C1507827|T201|COMP|35676-6|LNC2000|Chloride|Chloride
C1507829|T201|COMP|35678-2|LNC2000|Sodium|Sodium
C1507842|T201|COMP|35691-5|LNC2000|XXX microorganism DNA|XXX microorganism DNA
C1507883|T201|COMP|35732-7|LNC2000|Histoplasma capsulatum H Ab|Histoplasma capsulatum H Ab
C1507892|T201|COMP|35741-8|LNC2000|Prostate specific Ag|Prostate specific Ag
C1507940|T201|COMP|35789-7|LNC2000|DAPTOmycin|DAPTOmycin
C1508043|T201|COMP|36903-3|LNC2000|Chlamydia trachomatis & Neisseria gonorrhoeae DNA|Chlamydia trachomatis & Neisseria gonorrhoeae DNA
C1508044|T201|COMP|36904-1|LNC2000|Inhibin A^^adjusted|Inhibin A^^adjusted
C1508053|T201|COMP|36913-2|LNC2000|FMR1 gene targeted mutation analysis|FMR1 gene targeted mutation analysis
C1508056|T201|COMP|36916-5|LNC2000|Immunoglobulin light chains.kappa.free|Immunoglobulin light chains.kappa.free
C1508062|T201|COMP|36922-3|LNC2000|TPMT gene targeted mutation analysis|TPMT gene targeted mutation analysis
C1508100|T201|COMP|38168-1|LNC2000|Major crossmatch|Major crossmatch
C1508112|T201|COMP|38180-6|LNC2000|Hepatitis C virus RNA|Hepatitis C virus RNA
C1508141|T201|COMP|38256-4|LNC2000|Cells counted.total|Cells counted.total
C1526406|T201|COMP|38404-0|LNC2000|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C1526416|T201|COMP|38415-6|LNC2000|MTHFR gene targeted mutation analysis|MTHFR gene targeted mutation analysis
C1526477|T201|COMP|38476-8|LNC2000|Mullerian inhibiting substance|Mullerian inhibiting substance
C1526479|T201|COMP|38478-4|LNC2000|Biotinidase|Biotinidase
C1526480|T201|COMP|38479-2|LNC2000|Branched chain keto-acid dehydrogenase complex|Branched chain keto-acid dehydrogenase complex
C1526482|T201|COMP|38481-8|LNC2000|Carnitine.free (C0)|Carnitine.free (C0)
C1526484|T201|COMP|38483-4|LNC2000|Creatinine|Creatinine
C1526487|T201|COMP|38486-7|LNC2000|Homocystine|Homocystine
C1526495|T201|COMP|38494-1|LNC2000|Metanephrine.free|Metanephrine.free
C1526497|T201|COMP|38496-6|LNC2000|Retinyl palmitate|Retinyl palmitate
C1526506|T201|COMP|38505-4|LNC2000|Thyroglobulin recovery|Thyroglobulin recovery
C1526507|T201|COMP|38506-2|LNC2000|Thyroxine|Thyroxine
C1526527|T201|COMP|38526-0|LNC2000|Number of specimens tested|Number of specimens tested
C1526528|T201|COMP|38527-8|LNC2000|Number of specimens received|Number of specimens received
C1526541|T201|COMP|38540-1|LNC2000|Spermatozoa.motile/100 spermatozoa^pre washing|Spermatozoa.motile/100 spermatozoa^pre washing
C1526545|T201|COMP|38544-3|LNC2000|Spermatozoa^pre washing|Spermatozoa^pre washing
C1542992|T201|COMP|40527-4|LNC2000|Cocaine|Cocaine
C1543030|T201|COMP|38908-0|LNC2000|Poikilocytosis|Poikilocytosis
C1543117|T201|COMP|38995-7|LNC2000|Mixed cellular casts|Mixed cellular casts
C1543118|T201|COMP|38996-5|LNC2000|Neutrophils|Neutrophils
C1544439|T201|COMP|40464-0|LNC2000|Drugs identified|Drugs identified
C1544613|T201|COMP|40658-7|LNC2000|Parvovirus B19 Ab.IgM|Parvovirus B19 Ab.IgM
C1544647|T201|COMP|40692-6|LNC2000|Specimen volume^pre washing|Specimen volume^pre washing
C1544684|T201|COMP|40729-6|LNC2000|Herpes simplex virus Ab.IgM|Herpes simplex virus Ab.IgM
C1544705|T201|COMP|40750-2|LNC2000|Epstein Barr virus capsid Ab.IgG|Epstein Barr virus capsid Ab.IgG
C1544707|T201|COMP|40752-8|LNC2000|Epstein Barr virus early Ab.IgG|Epstein Barr virus early Ab.IgG
C1545091|T201|COMP|41163-7|LNC2000|Treponema pallidum DNA|Treponema pallidum DNA
C1545145|T201|COMP|41222-1|LNC2000|Yeast|Yeast
C1545197|T201|COMP|41274-2|LNC2000|Alpha-1-Fetoprotein interpretation|Alpha-1-Fetoprotein interpretation
C1624147|T201|COMP|42768-2|LNC2000|HIV 1 & 2 Ab|HIV 1 & 2 Ab
C1626279|T201|COMP|42803-7|LNC2000|Bacteria identified|Bacteria identified
C1627302|T201|COMP|42176-8|LNC2000|1,3 beta glucan|1,3 beta glucan
C1627329|T201|COMP|42810-2|LNC2000|Hemoglobin|Hemoglobin
C1627423|T201|COMP|41479-7|LNC2000|BK virus DNA|BK virus DNA
C1627424|T201|COMP|42481-2|LNC2000|Human papilloma virus 6+11+42+43+44 DNA|Human papilloma virus 6+11+42+43+44 DNA
C1628434|T201|COMP|42192-5|LNC2000|Nidus|Nidus
C1629582|T201|COMP|42216-2|LNC2000|Reference lab name|Reference lab name
C1629591|T201|COMP|42892-0|LNC2000|Citrulline|Citrulline
C1629593|T201|COMP|42906-8|LNC2000|Galactose 1 phosphate uridyl transferase|Galactose 1 phosphate uridyl transferase
C1630770|T201|COMP|42484-6|LNC2000|Protein.monoclonal/Protein.total|Protein.monoclonal/Protein.total
C1631779|T201|COMP|42247-7|LNC2000|Hemoglobin pattern|Hemoglobin pattern
C1632381|T201|COMP|42931-6|LNC2000|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1634498|T201|COMP|41499-5|LNC2000|Legionella pneumophila 1 Ag|Legionella pneumophila 1 Ag
C1637793|T201|COMP|41399-7|LNC2000|Herpes simplex virus 1+2 Ab.IgM|Herpes simplex virus 1+2 Ab.IgM
C1639534|T201|COMP|42483-8|LNC2000|Protein.monoclonal/Protein.total|Protein.monoclonal/Protein.total
C1641489|T201|COMP|41475-5|LNC2000|Rickettsia rickettsii Ab.IgM|Rickettsia rickettsii Ab.IgM
C1641490|T201|COMP|41476-3|LNC2000|Rickettsia rickettsii Ab.IgG|Rickettsia rickettsii Ab.IgG
C1642059|T201|COMP|42621-3|LNC2000|Mycoplasma hominis DNA|Mycoplasma hominis DNA
C1642549|T201|COMP|41477-1|LNC2000|Bacterial sialidase|Bacterial sialidase
C1642552|T201|COMP|41487-0|LNC2000|Cryptosporidium parvum Ag|Cryptosporidium parvum Ag
C1642559|T201|COMP|42637-9|LNC2000|Natriuretic peptide.B|Natriuretic peptide.B
C1642589|T201|COMP|41763-4|LNC2000|Rubella virus Ab.IgG|Rubella virus Ab.IgG
C1643184|T201|COMP|41480-5|LNC2000|BK virus DNA|BK virus DNA
C1645324|T201|COMP|41874-9|LNC2000|Betula populifolia Ab.IgE|Betula populifolia Ab.IgE
C1714522|T201|COMP|43180-9|LNC2000|Herpes simplex virus 2 Ab.IgG|Herpes simplex virus 2 Ab.IgG
C1714524|T201|COMP|43182-5|LNC2000|Smith extractable nuclear Ab|Smith extractable nuclear Ab
C1714656|T201|COMP|43304-5|LNC2000|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1714657|T201|COMP|43305-2|LNC2000|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1714718|T201|COMP|43371-4|LNC2000|Salmonella & Shigella sp identified|Salmonella & Shigella sp identified
C1714730|T201|COMP|43384-7|LNC2000|Neisseria sp identified|Neisseria sp identified
C1714740|T201|COMP|43396-1|LNC2000|Cholesterol.non HDL|Cholesterol.non HDL
C1714742|T201|COMP|43399-5|LNC2000|JAK2 gene.p.Val617Phe|JAK2 gene.p.Val617Phe
C1714780|T201|COMP|43441-5|LNC2000|Bacteria identified|Bacteria identified
C1715082|T201|COMP|43734-3|LNC2000|Coagulation surface induced|Coagulation surface induced
C1715279|T201|COMP|43994-3|LNC2000|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C1715280|T201|COMP|43995-0|LNC2000|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C1715592|T201|COMP|44357-2|LNC2000|Galactomannan Ag|Galactomannan Ag
C1715672|T201|COMP|44447-1|LNC2000|Beta 2 glycoprotein 1 Ab.IgA|Beta 2 glycoprotein 1 Ab.IgA
C1715673|T201|COMP|44449-7|LNC2000|Beta 2 glycoprotein 1 Ab.IgM|Beta 2 glycoprotein 1 Ab.IgM
C1715743|T201|COMP|44525-4|LNC2000|Histoplasma capsulatum Ag|Histoplasma capsulatum Ag
C1715746|T201|COMP|44528-8|LNC2000|Histoplasma capsulatum M Ab|Histoplasma capsulatum M Ab
C1715751|T201|COMP|44533-8|LNC2000|HIV 1+2 Ab|HIV 1+2 Ab
C1715754|T201|COMP|44538-7|LNC2000|HTLV I+II Ab|HTLV I+II Ab
C1715763|T201|COMP|44547-8|LNC2000|Human papilloma virus DNA|Human papilloma virus DNA
C1715875|T201|COMP|44607-0|LNC2000|HIV 1|HIV 1
C1716020|T201|COMP|44806-8|LNC2000|Chlamydia trachomatis+Neisseria gonorrhoeae DNA|Chlamydia trachomatis+Neisseria gonorrhoeae DNA
C1716241|T201|COMP|45084-1|LNC2000|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1716243|T201|COMP|45086-6|LNC2000|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C1716249|T201|COMP|45094-0|LNC2000|Chlamydia trachomatis|Chlamydia trachomatis
C1716334|T201|COMP|45197-1|LNC2000|Decanoylcarnitine (C10)|Decanoylcarnitine (C10)
C1716335|T201|COMP|45198-9|LNC2000|Decenoylcarnitine (C10:1)|Decenoylcarnitine (C10:1)
C1716336|T201|COMP|45199-7|LNC2000|Dodecanoylcarnitine (C12)|Dodecanoylcarnitine (C12)
C1716337|T201|COMP|45200-3|LNC2000|Dodecenoylcarnitine (C12:1)|Dodecenoylcarnitine (C12:1)
C1716348|T201|COMP|45211-0|LNC2000|Hexanoylcarnitine (C6)|Hexanoylcarnitine (C6)
C1716352|T201|COMP|45216-9|LNC2000|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)|Isovalerylcarnitine+Methylbutyrylcarnitine (C5)
C1716353|T201|COMP|45217-7|LNC2000|Linoleoylcarnitine (C18:2)|Linoleoylcarnitine (C18:2)
C1716358|T201|COMP|45222-7|LNC2000|Methylmalonylcarnitine (C4-DC)|Methylmalonylcarnitine (C4-DC)
C1716477|T201|COMP|45353-0|LNC2000|Date of analysis|Date of analysis
C1716512|T201|COMP|46082-4|LNC2000|Influenza virus A Ag|Influenza virus A Ag
C1716513|T201|COMP|46083-2|LNC2000|Influenza virus B Ag|Influenza virus B Ag
C1717149|T201|COMP|46128-5|LNC2000|Tissue transglutaminase Ab.IgA|Tissue transglutaminase Ab.IgA
C1717159|T201|COMP|46138-4|LNC2000|Urate crystals|Urate crystals
C1717174|T201|COMP|46154-1|LNC2000|Trichomonas vaginalis rRNA|Trichomonas vaginalis rRNA
C1717340|T201|COMP|44448-9|LNC2000|Beta 2 glycoprotein 1 Ab.IgG|Beta 2 glycoprotein 1 Ab.IgG
C1717373|T201|COMP|44877-9|LNC2000|Insulin dependent diabetes mellitus|Insulin dependent diabetes mellitus
C1717395|T201|COMP|45142-7|LNC2000|Sjogrens syndrome-B extractable nuclear Ab|Sjogrens syndrome-B extractable nuclear Ab
C1718546|T201|COMP|43583-4|LNC2000|Lipoprotein (little a)|Lipoprotein (little a)
C1765333|T201|COMP|14638-1|LNC2000|Calculus analysis|Calculus analysis
C1830059|T201|COMP|47213-4|LNC2000|Cholesterol.in LDL real size pattern|Cholesterol.in LDL real size pattern
C1830077|T201|COMP|47383-5|LNC2000|Nuclear Ab|Nuclear Ab
C1830096|T201|COMP|46266-3|LNC2000|Myeloperoxidase Ab|Myeloperoxidase Ab
C1830097|T201|COMP|46267-1|LNC2000|Proteinase 3 Ab|Proteinase 3 Ab
C1830098|T201|COMP|46268-9|LNC2000|ABO & Rh group^post transfusion reaction|ABO & Rh group^post transfusion reaction
C1830154|T201|COMP|46248-1|LNC2000|Borrelia burgdorferi Ab.IgG & IgM|Borrelia burgdorferi Ab.IgG & IgM
C1830309|T201|COMP|46420-6|LNC2000|Leukocyte clumps|Leukocyte clumps
C1830811|T201|COMP|46733-2|LNC2000|Amino acidemias|Amino acidemias
C1830813|T201|COMP|46735-7|LNC2000|Endocrine disorders|Endocrine disorders
C1830814|T201|COMP|46736-5|LNC2000|Fatty acid oxidation defects|Fatty acid oxidation defects
C1830815|T201|COMP|46737-3|LNC2000|Galactosemias|Galactosemias
C1830818|T201|COMP|46740-7|LNC2000|Hemoglobin disorders|Hemoglobin disorders
C1830822|T201|COMP|46744-9|LNC2000|Organic acidemias|Organic acidemias
C1830843|T201|COMP|46765-4|LNC2000|Sickle cell anemia|Sickle cell anemia
C1830847|T201|COMP|46769-6|LNC2000|Cystic fibrosis|Cystic fibrosis
C1831081|T201|COMP|46986-6|LNC2000|Cholesterol.in VLDL 3|Cholesterol.in VLDL 3
C1831090|T201|COMP|46994-0|LNC2000|HLA-A+B+C Ab|HLA-A+B+C Ab
C1831092|T201|COMP|46995-7|LNC2000|HLA-DP+DQ+DR Ab|HLA-DP+DQ+DR Ab
C1831099|T201|COMP|47000-5|LNC2000|Candida sp rRNA|Candida sp rRNA
C1831301|T201|COMP|47223-3|LNC2000|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C1831304|T201|COMP|47226-6|LNC2000|Fetal lung maturity|Fetal lung maturity
C1831317|T201|COMP|47238-1|LNC2000|Treponema pallidum Ab.IgG|Treponema pallidum Ab.IgG
C1831320|T201|COMP|47252-2|LNC2000|Hepatitis C virus RNA|Hepatitis C virus RNA
C1831382|T201|COMP|47320-7|LNC2000|Saccharomyces cerevisiae Ab.IgA|Saccharomyces cerevisiae Ab.IgA
C1831426|T201|COMP|47364-5|LNC2000|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C1831428|T201|COMP|47387-6|LNC2000|Neisseria gonorrhoeae DNA|Neisseria gonorrhoeae DNA
C1831486|T201|COMP|47440-3|LNC2000|Hepatitis B virus core Ab|Hepatitis B virus core Ab
C1831487|T201|COMP|47441-1|LNC2000|Hepatitis C virus Ab|Hepatitis C virus Ab
C1831574|T201|COMP|47527-7|LNC2000|Cytology report|Cytology report
C1831575|T201|COMP|47528-5|LNC2000|Cytology report|Cytology report
C1952805|T201|COMP|47562-4|LNC2000|Arginine|Arginine
C1952938|T201|COMP|47700-0|LNC2000|Methionine|Methionine
C1953090|T201|COMP|47784-4|LNC2000|Threonine|Threonine
C1953107|T201|COMP|47799-2|LNC2000|Valine|Valine
C1953409|T201|COMP|48035-0|LNC2000|Hemoglobin|Hemoglobin
C1953412|T201|COMP|48038-4|LNC2000|Pathologist interpretation|Pathologist interpretation
C1953413|T201|COMP|48039-2|LNC2000|Fibronectin.fetal|Fibronectin.fetal
C1953429|T201|COMP|48049-1|LNC2000|Eosinophils|Eosinophils
C1953430|T201|COMP|48050-9|LNC2000|Neutrophils|Neutrophils
C1953431|T201|COMP|48051-7|LNC2000|Erythrocytes|Erythrocytes
C1953433|T201|COMP|48053-3|LNC2000|Turbidity|Turbidity
C1953440|T201|COMP|48058-2|LNC2000|Fibrin D-dimer DDU|Fibrin D-dimer DDU
C1953449|T201|COMP|48065-7|LNC2000|Fibrin D-dimer FEU|Fibrin D-dimer FEU
C1953451|T201|COMP|48066-5|LNC2000|Fibrin D-dimer DDU|Fibrin D-dimer DDU
C1953564|T201|COMP|48159-8|LNC2000|Hepatitis C virus Ab Signal/Cutoff|Hepatitis C virus Ab Signal/Cutoff
C1953855|T201|COMP|48343-8|LNC2000|Hemoglobin.other/Hemoglobin.total|Hemoglobin.other/Hemoglobin.total
C1953856|T201|COMP|48344-6|LNC2000|Activated clotting time|Activated clotting time
C1953857|T201|COMP|48345-3|LNC2000|HIV 1+O+2 Ab|HIV 1+O+2 Ab
C1953859|T201|COMP|48346-1|LNC2000|HIV 1+O+2 Ab|HIV 1+O+2 Ab
C1953891|T201|COMP|48391-7|LNC2000|Carbon dioxide|Carbon dioxide
C1954123|T201|COMP|48560-7|LNC2000|Human papilloma virus genotype|Human papilloma virus genotype
C1954215|T201|COMP|48633-2|LNC2000|Trypsinogen I.free|Trypsinogen I.free
C1954294|T201|COMP|48683-7|LNC2000|Streptococcus agalactiae DNA|Streptococcus agalactiae DNA
C1954449|T201|COMP|48803-1|LNC2000|Neural tube defect risk|Neural tube defect risk
C1954772|T201|COMP|49041-7|LNC2000|Testosterone|Testosterone
C1954773|T201|COMP|49042-5|LNC2000|Testosterone.free|Testosterone.free
C1954781|T201|COMP|49047-4|LNC2000|Globulin|Globulin
C1954782|T201|COMP|49048-2|LNC2000|Protein feed time|Protein feed time
C1954784|T201|COMP|49049-0|LNC2000|Collection time|Collection time
C1954793|T201|COMP|49054-0|LNC2000|25-Hydroxycalciferol|25-Hydroxycalciferol
C1954800|T201|COMP|49058-1|LNC2000|Coagulation surface induced|Coagulation surface induced
C1954807|T201|COMP|49062-3|LNC2000|Lipid risk factors|Lipid risk factors
C1954849|T201|COMP|49090-4|LNC2000|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C1954853|T201|COMP|49092-0|LNC2000|Second trimester quad maternal screen|Second trimester quad maternal screen
C1954879|T201|COMP|49121-7|LNC2000|Erythrocyte inclusion bodies|Erythrocyte inclusion bodies
C1954900|T201|COMP|49136-5|LNC2000|Creatine kinase.MB/Creatine kinase.total|Creatine kinase.MB/Creatine kinase.total
C1955054|T201|COMP|49295-9|LNC2000|Protein pattern|Protein pattern
C1976907|T201|COMP|50194-0|LNC2000|Cholesterol.in IDL+Cholesterol.in VLDL 3|Cholesterol.in IDL+Cholesterol.in VLDL 3
C1976967|T201|COMP|49838-6|LNC2000|Neural tube defect risk|Neural tube defect risk
C1976968|T201|COMP|49839-4|LNC2000|Eosinophils|Eosinophils
C1976978|T201|COMP|49846-9|LNC2000|Hepatitis C virus core Ag|Hepatitis C virus core Ag
C1977068|T201|COMP|49578-8|LNC2000|Aminocaproate cutoff|Aminocaproate cutoff
C1977071|T201|COMP|49580-4|LNC2000|HIV 1+2 Ab|HIV 1+2 Ab
C1977072|T201|COMP|49581-2|LNC2000|Reference lab test identifier and name|Reference lab test identifier and name
C1977296|T201|COMP|49539-0|LNC2000|Cytomegalovirus Ab.IgM|Cytomegalovirus Ab.IgM
C1977297|T201|COMP|49540-8|LNC2000|Acid citrate dextrose|Acid citrate dextrose
C1977298|T201|COMP|49541-6|LNC2000|Fasting status|Fasting status
C1977299|T201|COMP|49542-4|LNC2000|Date and time of pheresis procedure|Date and time of pheresis procedure
C1977302|T201|COMP|49544-0|LNC2000|Newborn screening recommended follow-up|Newborn screening recommended follow-up
C1977318|T201|COMP|49563-0|LNC2000|Troponin I.cardiac|Troponin I.cardiac
C1977330|T201|COMP|49572-1|LNC2000|Second trimester triple maternal screen|Second trimester triple maternal screen
C1977331|T201|COMP|49573-9|LNC2000|HIV genotype|HIV genotype
C1977470|T201|COMP|49701-6|LNC2000|pH^^adjusted to patient's actual temperature|pH^^adjusted to patient's actual temperature
C1977653|T201|COMP|49835-2|LNC2000|Cells.CD19+IgD+/100 cells|Cells.CD19+IgD+/100 cells
C1977682|T201|COMP|50125-4|LNC2000|3-Hydroxypalmitoylcarnitine (C16-OH)|3-Hydroxypalmitoylcarnitine (C16-OH)
C1977965|T201|COMP|50106-4|LNC2000|3-Hydroxyisovalerylcarnitine (C5-OH)|3-Hydroxyisovalerylcarnitine (C5-OH)
C1977968|T201|COMP|50109-8|LNC2000|3-Hydroxylinoleoylcarnitine (C18:2-OH)|3-Hydroxylinoleoylcarnitine (C18:2-OH)
C1977973|T201|COMP|50113-0|LNC2000|3-Hydroxyoleoylcarnitine (C18:1-OH)|3-Hydroxyoleoylcarnitine (C18:1-OH)
C1977982|T201|COMP|50121-3|LNC2000|3-Hydroxypalmitoleylcarnitine (C16:1-OH)|3-Hydroxypalmitoleylcarnitine (C16:1-OH)
C1977985|T201|COMP|50132-0|LNC2000|3-Hydroxystearoylcarnitine (C18-OH)|3-Hydroxystearoylcarnitine (C18-OH)
C1978014|T201|COMP|50157-7|LNC2000|Acetylcarnitine (C2)|Acetylcarnitine (C2)
C1978123|T201|COMP|50281-5|LNC2000|3-Hydroxytetradecanoylcarnitine (C14-OH)|3-Hydroxytetradecanoylcarnitine (C14-OH)
C1978249|T201|COMP|50387-0|LNC2000|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C1978250|T201|COMP|50388-8|LNC2000|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C1978762|T201|COMP|50758-2|LNC2000|Herpes simplex virus 1 Ab.IgM|Herpes simplex virus 1 Ab.IgM
C1978817|T201|COMP|50970-3|LNC2000|XXX blood group Ab|XXX blood group Ab
C2359984|T201|COMP|53159-0|LNC2000|Tryptophan|Tryptophan
C2359985|T201|COMP|53160-8|LNC2000|Propionylcarnitine (C3)|Propionylcarnitine (C3)
C2359988|T201|COMP|53162-4|LNC2000|Propionylcarnitine (C3)/Carnitine.free (C0)|Propionylcarnitine (C3)/Carnitine.free (C0)
C2359990|T201|COMP|53163-2|LNC2000|Propionylcarnitine (C3)/Acetylcarnitine (C2)|Propionylcarnitine (C3)/Acetylcarnitine (C2)
C2359992|T201|COMP|53164-0|LNC2000|Propionylcarnitine (C3)/Palmitoylcarnitine (C16)|Propionylcarnitine (C3)/Palmitoylcarnitine (C16)
C2360327|T201|COMP|51656-7|LNC2000|Hepatitis C virus Ab Signal/Cutoff|Hepatitis C virus Ab Signal/Cutoff
C2360404|T201|COMP|51724-3|LNC2000|Cefuroxime|Cefuroxime
C2360474|T201|COMP|51775-5|LNC2000|Chromatin Ab|Chromatin Ab
C2360654|T201|COMP|51892-8|LNC2000|ABO group|ABO group
C2360674|T201|COMP|51916-5|LNC2000|Herpes simplex virus 1 Ab.IgG|Herpes simplex virus 1 Ab.IgG
C2360686|T201|COMP|51928-0|LNC2000|Ribonucleoprotein extractable nuclear Ab|Ribonucleoprotein extractable nuclear Ab
C2361418|T201|COMP|53398-4|LNC2000|Arginine/Phenylalanine|Arginine/Phenylalanine
C2361420|T201|COMP|53399-2|LNC2000|Citrulline/Tyrosine|Citrulline/Tyrosine
C2361550|T201|COMP|53062-6|LNC2000|Argininosuccinate|Argininosuccinate
C2361635|T201|COMP|53151-7|LNC2000|Valine/Phenylalanine|Valine/Phenylalanine
C2361637|T201|COMP|53152-5|LNC2000|Alloisoleucine+Isoleucine+Leucine+Hydroxyproline|Alloisoleucine+Isoleucine+Leucine+Hydroxyproline
C2361645|T201|COMP|53156-6|LNC2000|Methionine/Phenylalanine|Methionine/Phenylalanine
C2361647|T201|COMP|53157-4|LNC2000|Citrulline/Phenylalanine|Citrulline/Phenylalanine
C2361651|T201|COMP|53175-6|LNC2000|Octanoylcarnitine (C8)|Octanoylcarnitine (C8)
C2361652|T201|COMP|53176-4|LNC2000|Octanoylcarnitine (C8)/Acetylcarnitine (C2)|Octanoylcarnitine (C8)/Acetylcarnitine (C2)
C2361654|T201|COMP|53177-2|LNC2000|Octanoylcarnitine (C8)/Decanoylcarnitine (C10)|Octanoylcarnitine (C8)/Decanoylcarnitine (C10)
C2361664|T201|COMP|53182-2|LNC2000|3-Hydroxydecenoylcarnitine (C10:1-OH)|3-Hydroxydecenoylcarnitine (C10:1-OH)
C2361673|T201|COMP|53187-1|LNC2000|Methylglutarylcarnitine (C6-DC)|Methylglutarylcarnitine (C6-DC)
C2361675|T201|COMP|53188-9|LNC2000|3-Hydroxydodecenoylcarnitine (C12:1-OH)|3-Hydroxydodecenoylcarnitine (C12:1-OH)
C2361677|T201|COMP|53189-7|LNC2000|3-Hydroxydodecanoylcarnitine (C12-OH)|3-Hydroxydodecanoylcarnitine (C12-OH)
C2361678|T201|COMP|53190-5|LNC2000|Tetradecadienoylcarnitine (C14:2)|Tetradecadienoylcarnitine (C14:2)
C2361679|T201|COMP|53191-3|LNC2000|Tetradecenoylcarnitine (C14:1)|Tetradecenoylcarnitine (C14:1)
C2361680|T201|COMP|53192-1|LNC2000|Tetradecanoylcarnitine (C14)|Tetradecanoylcarnitine (C14)
C2361687|T201|COMP|53196-2|LNC2000|3-Hydroxytetradecadienoylcarnitine (C14:2-OH)|3-Hydroxytetradecadienoylcarnitine (C14:2-OH)
C2361689|T201|COMP|53197-0|LNC2000|3-Hydroxytetradecenoylcarnitine (C14:1-OH)|3-Hydroxytetradecenoylcarnitine (C14:1-OH)
C2361690|T201|COMP|53198-8|LNC2000|Palmitoleylcarnitine (C16:1)|Palmitoleylcarnitine (C16:1)
C2361691|T201|COMP|53199-6|LNC2000|Palmitoylcarnitine (C16)|Palmitoylcarnitine (C16)
C2361692|T201|COMP|53200-2|LNC2000|Argininosuccinate/Arginine|Argininosuccinate/Arginine
C2361696|T201|COMP|53202-8|LNC2000|Oleoylcarnitine (C18:1)|Oleoylcarnitine (C18:1)
C2361742|T201|COMP|53231-7|LNC2000|Succinylacetone|Succinylacetone
C2361760|T201|COMP|53241-6|LNC2000|Stearoylcarnitine (C18)|Stearoylcarnitine (C18)
C2361858|T201|COMP|53336-4|LNC2000|17-Hydroxyprogesterone+Androstenedione/Cortisol|17-Hydroxyprogesterone+Androstenedione/Cortisol
C2361861|T201|COMP|53338-0|LNC2000|11-Deoxycortisol|11-Deoxycortisol
C2361864|T201|COMP|53341-4|LNC2000|21-Deoxycortisol|21-Deoxycortisol
C2361866|T201|COMP|53343-0|LNC2000|Androstenedione|Androstenedione
C2361868|T201|COMP|53345-5|LNC2000|Cortisol|Cortisol
C2361870|T201|COMP|53347-1|LNC2000|11-Deoxycorticosterone|11-Deoxycorticosterone
C2363247|T201|COMP|779-9|LNC2000|Poikilocytosis|Poikilocytosis
C2363327|T201|COMP|26513-2|LNC2000|Neutrophils/100 leukocytes|Neutrophils/100 leukocytes
C2598073|T201|COMP|53926-2|LNC2000|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C2598074|T201|COMP|53927-0|LNC2000|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2598496|T201|COMP|53962-7|LNC2000|Alpha-1-Fetoprotein.tumor marker|Alpha-1-Fetoprotein.tumor marker
C2598793|T201|COMP|53879-3|LNC2000|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2599044|T201|COMP|53835-5|LNC2000|1,5-Anhydroglucitol|1,5-Anhydroglucitol
C2599173|T201|COMP|53925-4|LNC2000|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C2599234|T201|COMP|53982-5|LNC2000|Centromere protein B Ab|Centromere protein B Ab
C2599397|T201|COMP|54083-1|LNC2000|CFTR gene targeted mutation analysis|CFTR gene targeted mutation analysis
C2599398|T201|COMP|54084-9|LNC2000|Galactose|Galactose
C2599407|T201|COMP|54092-2|LNC2000|Citrulline/Arginine|Citrulline/Arginine
C2706780|T201|COMP|54218-3|LNC2000|Cells.CD3+CD4+/Cells.CD3+CD8+|Cells.CD3+CD4+/Cells.CD3+CD8+
C2734584|T201|COMP|56490-6|LNC2000|Hemoglobin.gastrointestinal.lower^2nd specimen|Hemoglobin.gastrointestinal.lower^2nd specimen
C2734585|T201|COMP|56491-4|LNC2000|Hemoglobin.gastrointestinal.lower^3rd specimen|Hemoglobin.gastrointestinal.lower^3rd specimen
C2734630|T201|COMP|56537-4|LNC2000|Tissue transglutaminase Ab.IgG|Tissue transglutaminase Ab.IgG
C2735715|T201|COMP|57288-3|LNC2000|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C2735716|T201|COMP|57289-1|LNC2000|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2736268|T201|COMP|57845-0|LNC2000|Leukocytes|Leukocytes
C2739456|T201|COMP|56598-6|LNC2000|Epstein Barr virus early Ab.IgM|Epstein Barr virus early Ab.IgM
C2923118|T201|COMP|58787-3|LNC2000|Corynebacterium diphtheriae Ab.IgG|Corynebacterium diphtheriae Ab.IgG
C2924090|T201|COMP|59841-7|LNC2000|Vendor name|Vendor name
C2926183|T201|COMP|58413-6|LNC2000|Erythrocytes.nucleated/100 leukocytes|Erythrocytes.nucleated/100 leukocytes
C2926219|T201|COMP|58448-2|LNC2000|Albumin ug/min|Albumin ug/min
C2970099|T201|COMP|60256-5|LNC2000|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C2973201|T201|COMP|62292-8|LNC2000|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3|25-Hydroxyvitamin D2+25-Hydroxyvitamin D3
C2973228|T201|COMP|62320-7|LNC2000|T-cell receptor excision circle|T-cell receptor excision circle
C2973278|T201|COMP|10329-1|LNC2000|Monocytes/100 leukocytes|Monocytes/100 leukocytes
C3173583|T201|COMP|64117-5|LNC2000|Most predominant hemoglobin|Most predominant hemoglobin
C3173585|T201|COMP|64118-3|LNC2000|Second most predominant hemoglobin|Second most predominant hemoglobin
C3173586|T201|COMP|64119-1|LNC2000|Third most predominant hemoglobin|Third most predominant hemoglobin
C3173587|T201|COMP|64120-9|LNC2000|Fourth most predominant hemoglobin|Fourth most predominant hemoglobin
C3173589|T201|COMP|64121-7|LNC2000|Fifth most predominant hemoglobin|Fifth most predominant hemoglobin
C3174659|T201|COMP|65751-0|LNC2000|Pathology biopsy report|Pathology biopsy report
C3174660|T201|COMP|65752-8|LNC2000|Pathology biopsy report|Pathology biopsy report
C3174662|T201|COMP|65754-4|LNC2000|Pathology biopsy report|Pathology biopsy report
C3174664|T201|COMP|65757-7|LNC2000|Pathology biopsy report|Pathology biopsy report
C3176086|T201|COMP|65633-0|LNC2000|Hepatitis B virus surface Ag|Hepatitis B virus surface Ag
C3262820|T201|COMP|68989-3|LNC2000|Performing laboratory|Performing laboratory
C3481505|T201|COMP|68325-0|LNC2000|Coagulation thrombin induced actual/Normal|Coagulation thrombin induced actual/Normal
C3481507|T201|COMP|68326-8|LNC2000|Coagulation reptilase induced actual/Normal|Coagulation reptilase induced actual/Normal
C3654082|T201|COMP|73970-6|LNC2000|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3654083|T201|COMP|73969-8|LNC2000|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3654084|T201|COMP|73968-0|LNC2000|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3654204|T201|COMP|73825-2|LNC2000|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3654205|T201|COMP|73824-5|LNC2000|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3654207|T201|COMP|73822-9|LNC2000|Fetal chromosome X & Y aneuploidy|Fetal chromosome X & Y aneuploidy
C3654208|T201|COMP|73821-1|LNC2000|Fetal chromosome X & Y aneuploidy risk|Fetal chromosome X & Y aneuploidy risk
C3654286|T201|COMP|73697-5|LNC2000|CCHD newborn screening protocol used|CCHD newborn screening protocol used
C3654308|T201|COMP|73967-2|LNC2000|Noninvasive prenatal fetal aneuploidy test panel|Noninvasive prenatal fetal aneuploidy test panel
C3654309|T201|COMP|73966-4|LNC2000|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3846791|T201|COMP|75217-0|LNC2000|Biotinidase|Biotinidase
C3846797|T201|COMP|75211-3|LNC2000|Propionylcarnitine (C3)+Palmitoylcarnitine (C16)|Propionylcarnitine (C3)+Palmitoylcarnitine (C16)
C3853768|T201|COMP|12286-1|LNC2000|Drugs identified|Drugs identified
C3853963|T201|COMP|75574-4|LNC2000|22q11.2 deletion prior risk|22q11.2 deletion prior risk
C3853964|T201|COMP|75568-6|LNC2000|Monosomy X prior risk|Monosomy X prior risk
C3853965|T201|COMP|75566-0|LNC2000|Monosomy X prior risk|Monosomy X prior risk
C3853966|T201|COMP|75546-2|LNC2000|Trisomy 13 prior risk|Trisomy 13 prior risk
C3853967|T201|COMP|75550-4|LNC2000|Trisomy 13 prior risk|Trisomy 13 prior risk
C3853968|T201|COMP|75556-1|LNC2000|Trisomy 18 prior risk|Trisomy 18 prior risk
C3853969|T201|COMP|75554-6|LNC2000|Trisomy 18 prior risk|Trisomy 18 prior risk
C3853970|T201|COMP|75562-9|LNC2000|Trisomy 21 prior risk|Trisomy 21 prior risk
C3853971|T201|COMP|75560-3|LNC2000|Trisomy 21 prior risk|Trisomy 21 prior risk
C3861011|T201|COMP|75599-1|LNC2000|1p36 deletion prior risk|1p36 deletion prior risk
C3864290|T201|COMP|75575-1|LNC2000|22q11.2 deletion prior risk|22q11.2 deletion prior risk
C3864940|T201|COMP|75598-3|LNC2000|1p36 deletion prior risk|1p36 deletion prior risk
C3870263|T201|COMP|75608-0|LNC2000|Citation|Citation
C3870264|T201|COMP|75607-2|LNC2000|Paternal sample received|Paternal sample received
C3870265|T201|COMP|75606-4|LNC2000|Cell-free DNA.fetal/Cell-free DNA.total|Cell-free DNA.fetal/Cell-free DNA.total
C3870266|T201|COMP|75605-6|LNC2000|Cell-free DNA.fetal/Cell-free DNA.total|Cell-free DNA.fetal/Cell-free DNA.total
C3870267|T201|COMP|75604-9|LNC2000|Fetal sex|Fetal sex
C3870269|T201|COMP|75602-3|LNC2000|Fetal 1p36 deletion risk|Fetal 1p36 deletion risk
C3870270|T201|COMP|75601-5|LNC2000|Fetal 1p36 deletion risk|Fetal 1p36 deletion risk
C3870271|T201|COMP|75600-7|LNC2000|Fetal 1p36 deletion risk|Fetal 1p36 deletion risk
C3870273|T201|COMP|75596-7|LNC2000|Fetal 5p deletion risk|Fetal 5p deletion risk
C3870274|T201|COMP|75595-9|LNC2000|Fetal 5p deletion risk|Fetal 5p deletion risk
C3870275|T201|COMP|75594-2|LNC2000|Fetal 5p deletion risk|Fetal 5p deletion risk
C3870276|T201|COMP|75593-4|LNC2000|5p deletion prior risk|5p deletion prior risk
C3870277|T201|COMP|75592-6|LNC2000|5p deletion prior risk|5p deletion prior risk
C3870279|T201|COMP|75590-0|LNC2000|Fetal Angelman syndrome risk|Fetal Angelman syndrome risk
C3870280|T201|COMP|75589-2|LNC2000|Fetal Angelman syndrome risk|Fetal Angelman syndrome risk
C3870281|T201|COMP|75588-4|LNC2000|Fetal Angelman syndrome risk|Fetal Angelman syndrome risk
C3870282|T201|COMP|75587-6|LNC2000|Angelman syndrome prior risk|Angelman syndrome prior risk
C3870283|T201|COMP|75586-8|LNC2000|Angelman syndrome prior risk|Angelman syndrome prior risk
C3870285|T201|COMP|75584-3|LNC2000|Fetal Prader-Willi syndrome risk|Fetal Prader-Willi syndrome risk
C3870291|T201|COMP|75583-5|LNC2000|Fetal Prader-Willi syndrome risk|Fetal Prader-Willi syndrome risk
C3870292|T201|COMP|75582-7|LNC2000|Fetal Prader-Willi syndrome risk|Fetal Prader-Willi syndrome risk
C3870293|T201|COMP|75581-9|LNC2000|Prader-Willi syndrome prior risk|Prader-Willi syndrome prior risk
C3870294|T201|COMP|75580-1|LNC2000|Prader-Willi syndrome prior risk|Prader-Willi syndrome prior risk
C3870296|T201|COMP|75578-5|LNC2000|Fetal 22q11.2 deletion risk|Fetal 22q11.2 deletion risk
C3870297|T201|COMP|75577-7|LNC2000|Fetal 22q11.2 deletion risk|Fetal 22q11.2 deletion risk
C3870298|T201|COMP|75576-9|LNC2000|Fetal 22q11.2 deletion risk|Fetal 22q11.2 deletion risk
C3870299|T201|COMP|75573-6|LNC2000|Genetic counselor comment on fetal Triploidy risk|Genetic counselor comment on fetal Triploidy risk
C3870300|T201|COMP|75572-8|LNC2000|Fetal triploidy risk|Fetal triploidy risk
C3870302|T201|COMP|75570-2|LNC2000|Fetal monosomy X risk|Fetal monosomy X risk
C3870303|T201|COMP|75569-4|LNC2000|Fetal monosomy X risk|Fetal monosomy X risk
C3870304|T201|COMP|75567-8|LNC2000|Fetal monosomy X risk|Fetal monosomy X risk
C3870306|T201|COMP|75564-5|LNC2000|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3870307|T201|COMP|75563-7|LNC2000|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3870308|T201|COMP|75561-1|LNC2000|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C3870310|T201|COMP|75558-7|LNC2000|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3870311|T201|COMP|75557-9|LNC2000|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3870312|T201|COMP|75555-3|LNC2000|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C3870314|T201|COMP|75552-0|LNC2000|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3870315|T201|COMP|75551-2|LNC2000|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3870317|T201|COMP|75548-8|LNC2000|Fetal trisomy 13 risk|Fetal trisomy 13 risk
C3870340|T201|COMP|75513-2|LNC2000|DRVVT with 1:1 Pooled Normal Plasma|DRVVT with 1:1 Pooled Normal Plasma
C3870341|T201|COMP|75512-4|LNC2000|DRVVT with 1:1 Pooled Normal Plasma actual/Normal|DRVVT with 1:1 Pooled Normal Plasma actual/Normal
C3870342|T201|COMP|75511-6|LNC2000|DRVVT percent correction|DRVVT percent correction
C4018866|T201|COMP|77012-3|LNC2000|Fetal chromosome 18 trisomy|Fetal chromosome 18 trisomy
C4018867|T201|COMP|77011-5|LNC2000|Fetal chromosome 21 trisomy|Fetal chromosome 21 trisomy
C4019186|T201|COMP|77013-1|LNC2000|Fetal chromosome 13 trisomy|Fetal chromosome 13 trisomy
C4037269|T201|COMP|77015-6|LNC2000|Fetal trisomy 18 risk|Fetal trisomy 18 risk
C4037270|T201|COMP|77014-9|LNC2000|Fetal trisomy 21 risk|Fetal trisomy 21 risk
C4037661|T201|COMP|77021-4|LNC2000|Fetal Y chromosome|Fetal Y chromosome
C4037662|T201|COMP|77020-6|LNC2000|Fetal Y chromosome|Fetal Y chromosome
C4069397|T201|COMP|80369-2|LNC2000|Neisseria sp identified|Neisseria sp identified
C4069398|T201|COMP|80368-4|LNC2000|Neisseria gonorrhoeae|Neisseria gonorrhoeae
C4069399|T201|COMP|80367-6|LNC2000|Chlamydia trachomatis|Chlamydia trachomatis
C4069400|T201|COMP|80366-8|LNC2000|Neisseria gonorrhoeae rRNA|Neisseria gonorrhoeae rRNA
C4069401|T201|COMP|80365-0|LNC2000|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C4069402|T201|COMP|80364-3|LNC2000|Chlamydia trachomatis rRNA|Chlamydia trachomatis rRNA
C4069403|T201|COMP|80363-5|LNC2000|Chlamydia trachomatis DNA|Chlamydia trachomatis DNA
C4069404|T201|COMP|80362-7|LNC2000|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C4069405|T201|COMP|80361-9|LNC2000|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C4069406|T201|COMP|80360-1|LNC2000|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA|Chlamydia trachomatis+Neisseria gonorrhoeae rRNA
C4071394|T201|COMP|78012-2|LNC2000|Streptococcus pyogenes Ag|Streptococcus pyogenes Ag
C4318962|T201|COMP|85954-6|LNC2000|Streptococcus pneumoniae Danish serotype 1 Ab.IgG|Streptococcus pneumoniae Danish serotype 1 Ab.IgG
C4319061|T201|COMP|86107-0|LNC2000|Streptococcus pneumoniae Danish serotype 4 Ab.IgG|Streptococcus pneumoniae Danish serotype 4 Ab.IgG
C4319115|T201|COMP|86108-8|LNC2000|Streptococcus pneumoniae Danish serotype 4 Ab.IgG|Streptococcus pneumoniae Danish serotype 4 Ab.IgG
C4483418|T201|COMP|85955-3|LNC2000|Streptococcus pneumoniae Danish serotype 1 Ab.IgG|Streptococcus pneumoniae Danish serotype 1 Ab.IgG
C4483541|T201|COMP|86080-9|LNC2000|Streptococcus pneumoniae Danish serotype 3 Ab.IgG|Streptococcus pneumoniae Danish serotype 3 Ab.IgG
C4483543|T201|COMP|86081-7|LNC2000|Streptococcus pneumoniae Danish serotype 3 Ab.IgG|Streptococcus pneumoniae Danish serotype 3 Ab.IgG
C4483631|T201|COMP|86147-6|LNC2000|Streptococcus pneumoniae Danish serotype 8 Ab.IgG|Streptococcus pneumoniae Danish serotype 8 Ab.IgG
C4483633|T201|COMP|86148-4|LNC2000|Streptococcus pneumoniae Danish serotype 8 Ab.IgG|Streptococcus pneumoniae Danish serotype 8 Ab.IgG
