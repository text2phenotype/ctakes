C0079304|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY
C0009378|T060|1007622|CPT|COLONOSCOPY|ENDOSCOPY PROCEDURES ON THE RECTUM
C0079304|T060||CPT|ESOPHAGOGASTRODUODENOSCOPIES
C0079304|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY
C0079304|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY
C0079304|T060||CPT|FIBREOPTIC OESOPHAGOGASTRODUODENOSCOPY 
C0079304|T060||CPT|FIBEROPTIC ESOPHAGOGASTRODUODENOSCOPY 
C0079304|T060||CPT|ENDOSCOPY UPPER GASTROINTESTINAL TRACT
C0079304|T060||CPT|EGD
C0079304|T060||CPT|UPPER GI ENDOSCOPY
C0079304|T060||CPT|ENDOSCOPIC EXAMINATION OF OESOPHAGUS, STOMACH AND DUODENUM
C0079304|T060||CPT|ENDOSCOPIC EXAMINATION OF ESOPHAGUS, STOMACH AND DUODENUM 
C0079304|T060||CPT|COMBINED UPPER GI ENDOSCOPY
C0079304|T060||CPT|OGD - ESOPHAGOGASTRODUODENOSCOPY
C0079304|T060||CPT|OGD - OESOPHAGOGASTRODUODENOSCOPY
C0079304|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY 
C0079304|T060||CPT|ENDOSCOPIC EXAMINATION OF UPPER GI TRACT
C0079304|T060||CPT|FIBREOPTIC OESOPHAGOGASTRODUODENOSCOPY
C0079304|T060||CPT|FIBEROPTIC ESOPHAGOGASTRODUODENOSCOPY
C0079304|T060||CPT|ENDOSCOPIC EXAMINATION OF ESOPHAGUS, STOMACH AND DUODENUM
C0079304|T060||CPT|UPPER GASTROINTESTINAL ENDOSCOPY
C0079304|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY PROCEDURES
C0079304|T060||CPT|DIAGNOSTIC ESOPHAGOGASTRODUODENOSCOPY 
C0079304|T060||CPT|DIAGNOSTIC ESOPHAGOGASTRODUODENOSCOPY
C0079304|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY 
C0079304|T060||CPT|UPPER GASTROINTESTINAL TRACT ENDOSCOPY
C0079304|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY 
C0472993|T060||CPT|FIBEROPTIC ENDOSCOPIC SNARE RESECTION OF LESION OF ESOPHAGUS
C0472993|T060||CPT|FIBREOPTIC ENDOSCOPIC SNARE RESECTION OF LESION OF OESOPHAGUS
C0472993|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND SNARE RESECTION
C0472993|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY AND SNARE RESECTION
C0472993|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND SNARE RESECTION 
C0472984|T060||CPT|FIBEROPTIC ENDOSCOPIC LASER DESTRUCTION OF LESION OF ESOPHAGUS
C0472984|T060||CPT|FIBREOPTIC ENDOSCOPIC LASER DESTRUCTION OF LESION OF OESOPHAGUS
C0472984|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND LASER
C0472984|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY AND LASER
C0472984|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND LASER 
C0472981|T060||CPT|FIBEROPTIC ENDOSCOPIC CAUTERIZATION OF LESION OF ESOPHAGUS
C0472981|T060||CPT|FIBREOPTIC ENDOSCOPIC CAUTERISATION OF LESION OF OESOPHAGUS
C0472981|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY AND CAUTERISATION
C0472981|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND CAUTERIZATION
C0472981|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND CAUTERIZATION 
C0472989|T060||CPT|FIBEROPTIC ENDOSCOPIC INJECTION SCLEROTHERAPY TO ESOPHAGEAL VARICES
C0472989|T060||CPT|FIBREOPTIC ENDOSCOPIC INJECTION SCLEROTHERAPY TO OESOPHAGEAL VARICES
C0472989|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES
C0472989|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES
C0472989|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES 
C0472952|T060||CPT|FIBEROPTIC ENDOSCOPIC BANDING OF ESOPHAGEAL VARICES
C0472952|T060||CPT|FIBREOPTIC ENDOSCOPIC BANDING OF OESOPHAGEAL VARICES
C0472952|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND BANDING OF ESOPHAGEAL VARICES
C0472952|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY AND BANDING OF OESOPHAGEAL VARICES
C0472952|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND BANDING OF ESOPHAGEAL VARICES 
C0472966|T060||CPT|FIBEROPTIC ENDOSCOPIC REMOVAL OF FOREIGN BODY FROM ESOPHAGUS
C0472966|T060||CPT|FIBREOPTIC ENDOSCOPIC REMOVAL OF FOREIGN BODY FROM OESOPHAGUS
C0472966|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND REMOVAL OF FOREIGN BODY
C0472966|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY AND REMOVAL OF FOREIGN BODY
C0472966|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND REMOVAL OF FOREIGN BODY 
C0472973|T060||CPT|FIBEROPTIC ENDOSCOPIC BALLOON DILATION OF ESOPHAGUS
C0472973|T060||CPT|FIBREOPTIC ENDOSCOPIC BALLOON DILATION OF OESOPHAGUS
C0472973|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND BALLOON DILATATION
C0472973|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY AND BALLOON DILATATION
C0472973|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND BALLOON DILATATION 
C0472962|T060||CPT|DIAGNOSTIC FIBEROPTIC ENDOSCOPIC EXAMINATION OF ESOPHAGUS AND BIOPSY OF LESION OF ESOPHAGUS
C0472962|T060||CPT|DIAGNOSTIC FIBREOPTIC ENDOSCOPIC EXAMINATION OF OESOPHAGUS AND BIOPSY OF LESION OF OESOPHAGUS
C0472962|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND BIOPSY
C0472962|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY AND BIOPSY
C0472962|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND BIOPSY 
C0472992|T060||CPT|ENDOSCOPIC SNARE RESECTION OF LESION OF ESOPHAGUS USING RIGID ESOPHAGOSCOPE
C0472992|T060||CPT|ENDOSCOPIC SNARE RESECTION OF LESION OF OESOPHAGUS USING RIGID OESOPHAGOSCOPE
C0472992|T060||CPT|RIGID ESOPHAGOSCOPY AND SNARE RESECTION
C0472992|T060||CPT|RIGID OESOPHAGOSCOPY AND SNARE RESECTION
C0472992|T060||CPT|RIGID ESOPHAGOSCOPY AND SNARE RESECTION 
C0472983|T060||CPT|ENDOSCOPIC LASER DESTRUCTION OF LESION OF ESOPHAGUS USING RIGID ESOPHAGOSCOPE
C0472983|T060||CPT|ENDOSCOPIC LASER DESTRUCTION OF LESION OF OESOPHAGUS USING RIGID OESOPHAGOSCOPE
C0472983|T060||CPT|RIGID ESOPHAGOSCOPY AND LASER
C0472983|T060||CPT|RIGID OESOPHAGOSCOPY AND LASER
C0472983|T060||CPT|RIGID ESOPHAGOSCOPY AND LASER 
C0472980|T060||CPT|ENDOSCOPIC CAUTERISATION OF LESION OF OESOPHAGUS USING RIGID OESOPHAGOSCOPE
C0472980|T060||CPT|ENDOSCOPIC CAUTERIZATION OF LESION OF ESOPHAGUS USING RIGID ESOPHAGOSCOPE
C0472980|T060||CPT|RIGID OESOPHAGOSCOPY AND CAUTERISATION
C0472980|T060||CPT|RIGID ESOPHAGOSCOPY AND CAUTERIZATION
C0472980|T060||CPT|RIGID ESOPHAGOSCOPY AND CAUTERIZATION 
C0472988|T060||CPT|ENDOSCOPIC INJECTION SCLEROTHERAPY TO VARICES OF ESOPHAGUS USING RIGID ESOPHAGOSCOPE
C0472988|T060||CPT|ENDOSCOPIC INJECTION SCLEROTHERAPY TO VARICES OF OESOPHAGUS USING RIGID OESOPHAGOSCOPE
C0472988|T060||CPT|RIGID ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES
C0472988|T060||CPT|RIGID OESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES
C0472988|T060||CPT|RIGID ESOPHAGOSCOPY AND INJECTION SCLEROTHERAPY OF VARICES 
C0472951|T060||CPT|RIGID ESOPHAGOSCOPIC BANDING OF ESOPHAGEAL VARICES
C0472951|T060||CPT|RIGID OESOPHAGOSCOPIC BANDING OF OESOPHAGEAL VARICES
C0472951|T060||CPT|RIGID ESOPHAGOSCOPY AND BANDING OF ESOPHAGEAL VARICES
C0472951|T060||CPT|RIGID OESOPHAGOSCOPY AND BANDING OF OESOPHAGEAL VARICES
C0472951|T060||CPT|RIGID ESOPHAGOSCOPY AND BANDING OF ESOPHAGEAL VARICES 
C0472965|T060||CPT|RIGID ESOPHAGOSCOPY WITH REMOVAL OF FOREIGN BODY
C0472965|T060||CPT|ESOPHAGOSCOPY FOREIGN BODY REMOVAL
C0472965|T060||CPT|RIGID ESOPHAGOSCOPY WITH FOREIGN BODY REMOVAL 
C0472965|T060||CPT|RIGID ESOPHAGOSCOPY WITH FOREIGN BODY REMOVAL
C0472965|T060||CPT|ENDOSCOPIC REMOVAL OF FOREIGN BODY FROM ESOPHAGUS USING RIGID ESOPHAGOSCOPE
C0472965|T060||CPT|ENDOSCOPIC REMOVAL OF FOREIGN BODY FROM OESOPHAGUS USING RIGID OESOPHAGOSCOPE
C0472965|T060||CPT|RIGID ESOPHAGOSCOPY AND REMOVAL OF FOREIGN BODY
C0472965|T060||CPT|RIGID OESOPHAGOSCOPY AND REMOVAL OF FOREIGN BODY
C0472965|T060||CPT|RIGID ESOPHAGOSCOPY AND REMOVAL OF FOREIGN BODY 
C0472972|T060||CPT|ENDOSCOPIC BALLOON DILATION OF ESOPHAGUS USING RIGID ESOPHAGOSCOPE
C0472972|T060||CPT|ENDOSCOPIC BALLOON DILATION OF OESOPHAGUS USING RIGID OESOPHAGOSCOPE
C0472972|T060||CPT|RIGID ESOPHAGOSCOPY AND BALLOON DILATATION
C0472972|T060||CPT|RIGID OESOPHAGOSCOPY AND BALLOON DILATATION
C0472972|T060||CPT|RIGID ESOPHAGOSCOPY AND BALLOON DILATATION 
C0472961|T060||CPT|RIGID ESOPHAGOSCOPY WITH BIOPSY
C0472961|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF ESOPHAGUS AND BIOPSY OF LESION OF ESOPHAGUS USING RIGID ESOPHAGOSCOPE
C0472961|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF OESOPHAGUS AND BIOPSY OF LESION OF OESOPHAGUS USING RIGID OESOPHAGOSCOPE
C0472961|T060||CPT|RIGID ESOPHAGOSCOPY AND BIOPSY
C0472961|T060||CPT|RIGID OESOPHAGOSCOPY AND BIOPSY
C0472961|T060||CPT|RIGID ESOPHAGOSCOPY AND BIOPSY 
C0472857|T060||CPT|FIBEROPTIC ENDOSCOPIC EXAMINATION OF UPPER GASTROINTESTINAL TRACT AND BIOPSY OF LESION OF UPPER GASTROINTESTINAL TRACT
C0472857|T060||CPT|FIBREOPTIC ENDOSCOPIC EXAMINATION OF UPPER GASTROINTESTINAL TRACT AND BIOPSY OF LESION OF UPPER GASTROINTESTINAL TRACT
C0472857|T060||CPT|FIBEROPTIC ENDOSCOPIC EXAMINATION OF UPPER GASTROINTESTINAL TRACT AND BIOPSY OF LESION OF UPPER GASTROINTESTINAL TRACT 
C0399776|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF DUODENUM NOS 
C0399776|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF DUODENUM NOS
C0399776|T060||CPT|DIAGNOSTIC DUODENOSCOPY
C0399776|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF DUODENUM
C0399776|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF DUODENUM 
C0192310|T060||CPT|ESOPHAGOSCOPY FOR REMOVAL OF POLYPOID LESION
C0192310|T060||CPT|OESOPHAGOSCOPY FOR REMOVAL OF POLYPOID LESION
C0192310|T060||CPT|ESOPHAGOSCOPY FOR REMOVAL OF POLYPOID LESION 
C0475192|T060||CPT|FIBEROPTIC ENDOSCOPIC INSERTION OF TUBAL PROSTHESIS INTO ESOPHAGUS
C0475192|T060||CPT|FIBREOPTIC ENDOSCOPIC INSERTION OF TUBAL PROSTHESIS INTO OESOPHAGUS
C0475192|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND INSERTION OF TUBE PROSTHESIS
C0475192|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY AND INSERTION OF TUBE PROSTHESIS
C0475192|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY AND INSERTION OF TUBE PROSTHESIS 
C0472996|T060||CPT|ENDOSCOPIC INSERTION OF TUBAL PROSTHESIS INTO ESOPHAGUS USING RIGID ESOPHAGOSCOPE
C0472996|T060||CPT|ENDOSCOPIC INSERTION OF TUBAL PROSTHESIS INTO OESOPHAGUS USING RIGID OESOPHAGOSCOPE
C0472996|T060||CPT|RIGID ESOPHAGOSCOPY AND INSERTION OF TUBE PROSTHESIS
C0472996|T060||CPT|RIGID OESOPHAGOSCOPY AND INSERTION OF TUBE PROSTHESIS
C0472996|T060||CPT|RIGID ESOPHAGOSCOPY AND INSERTION OF TUBE PROSTHESIS 
C0472855|T060||CPT|DIAGNOSTIC FIBEROPTIC ENDOSCOPIC EXAMINATION OF UPPER GASTROINTESTINAL TRACT NOS
C0472855|T060||CPT|DIAGNOSTIC FIBREOPTIC ENDOSCOPIC EXAMINATION OF UPPER GASTROINTESTINAL TRACT NOS
C0472855|T060||CPT|DIAGNOSTIC FIBEROPTIC ENDOSCOPIC EXAMINATION OF UPPER GASTROINTESTINAL TRACT NOS 
C0472855|T060||CPT|DIAGNOSTIC FIBREOPTIC ENDOSCOPIC EXAMINATION OF UPPER GASTROINTESTINAL TRACT
C0472855|T060||CPT|DIAGNOSTIC FIBEROPTIC ENDOSCOPIC EXAMINATION OF UPPER GASTROINTESTINAL TRACT
C0472855|T060||CPT|DIAGNOSTIC FIBEROPTIC ENDOSCOPIC EXAMINATION OF UPPER GASTROINTESTINAL TRACT 
C0192317|T060||CPT|ESOPHAGOSCOPY FOR DIRECT DILATION
C0192317|T060||CPT|OESOPHAGOSCOPY FOR DIRECT DILATION
C0192317|T060||CPT|ESOPHAGOSCOPY FOR DIRECT DILATION 
C0192467|T060||CPT|UPPER GASTROINTESTINAL ENDOSCOPY WITH DIRECTED PLACEMENT OF PERCUTANEOUS GASTROSTOMY-TUBE 
C0192467|T060||CPT|UPPER GASTROINTESTINAL ENDOSCOPY WITH DIRECTED PLACEMENT OF PERCUTANEOUS GASTROSTOMY-TUBE
C0192467|T060||CPT|UPPER GI ENDOSCOPY WITH DIRECTED PLACEMENT OF PERCUTANEOUS GASTROSTOMY-TUBE
C0192467|T060||CPT|UPPER GASTROINTESTINAL ENDOSCOPY WITH DIRECTED PLACEMENT OF PERCUTANEOUS GASTROSTOMY TUBE
C0192467|T060||CPT|UPPER GASTROINTESTINAL ENDOSCOPY FOR DIRECTED PLACEMENT OF PERCUTANEOUS GASTROSTOMY TUBE
C0192467|T060||CPT|UPPER GASTROINTESTINAL ENDOSCOPY FOR DIRECTED PLACEMENT OF PERCUTANEOUS GASTROSTOMY TUBE 
C2733057|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH ENDOSCOPIC ULTRASOUND OF UPPER GASTROINTESTINAL TRACT 
C2733057|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH ENDOSCOPIC ULTRASOUND OF UPPER GASTROINTESTINAL TRACT
C2733057|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY WITH ENDOSCOPIC ULTRASOUND OF UPPER GASTROINTESTINAL TRACT
C2733463|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH DIRECTED SUBMUCOSAL INJECTION 
C2733463|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY WITH DIRECTED SUBMUCOSAL INJECTION
C2733463|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH DIRECTED SUBMUCOSAL INJECTION
C0192318|T060|43226|CPT|ESOPHAGOSCOPY FOR INSERTION OF WIRE TO GUIDE DILATION|ESOPH ENDOSCOPY DILATION
C0192318|T060|43226|CPT|ESOPH ENDOSCOPY DILATION|ESOPH ENDOSCOPY DILATION
C0192318|T060|43226|CPT|ESOPHAGOSCOPY, FLEXIBLE, TRANSORAL; WITH INSERTION OF GUIDE WIRE FOLLOWED BY PASSAGE OF DILATOR(S) OVER GUIDE WIRE|ESOPH ENDOSCOPY DILATION
C0192318|T060|43226|CPT|ESOPHAGOSCOPY FLEXIBLE GUIDE WIRE DILATION|ESOPH ENDOSCOPY DILATION
C0192318|T060|43226|CPT|OESOPHAGOSCOPY FOR INSERTION OF WIRE TO GUIDE DILATION|ESOPH ENDOSCOPY DILATION
C0192318|T060|43226|CPT|ESOPHAGOSCOPY FOR INSERTION OF WIRE TO GUIDE DILATION |ESOPH ENDOSCOPY DILATION
C0192312|T060||CPT|FB - ESOPHOSCOPY AND REMOVAL OF FOREIGN BODY
C0192312|T060||CPT|FB - ESOPHAGOSCOPY AND REMOVAL OF FOREIGN BODY
C0192312|T060||CPT|ESOPHAGOSCOPY FOR REMOVAL OF FOREIGN BODY
C0192312|T060||CPT|REMOV INTRALUM ESOPH FB
C0192312|T060||CPT|ENDOSCOPIC REMOVAL OF INTRALUMINAL FOREIGN BODY FROM ESOPHAGUS WITHOUT INCISION
C0192312|T060||CPT|ENDOSCOPIC REMOVAL OF INTRALUMINAL FOREIGN BODY FROM OESOPHAGUS WITHOUT INCISION
C0192312|T060||CPT|OESOPHAGOSCOPY FOR REMOVAL OF FOREIGN BODY
C0192312|T060||CPT|ESOPHAGOSCOPY AND REMOVAL OF FOREIGN BODY
C0192312|T060||CPT|FB - OESOPHOSCOPY AND REMOVAL OF FOREIGN BODY
C0192312|T060||CPT|OESOPHAGOSCOPY AND REMOVAL OF FOREIGN BODY
C0192312|T060||CPT|ESOPHAGOSCOPY FOR REMOVAL OF FOREIGN BODY 
C0192312|T060||CPT|REMOVAL OF INTRALUMINAL FOREIGN BODY FROM ESOPHAGUS WITHOUT INCISION
C0192316|T060||CPT|ESOPHAGOSCOPY FOR INJECTION OF ESOPHAGEAL VARICES
C0192316|T060||CPT|INJECTION OF SCLEROSING AGENT INTO ESOPHAGEAL VARICES BY ENDOSCOPY
C0192316|T060||CPT|ENDOSCOPIC INJECTION OF ESOPHAGEAL VARICES
C0192316|T060||CPT|INJECTION OF ESOPHAGEAL VARICES BY ENDOSCOPY
C0192316|T060||CPT|INJECTION OF VARICOSE VEINS OF ESOPHAGUS BY ENDOSCOPY
C0192316|T060||CPT|ENDOSCOPIC INJECTION OF OESOPHAGEAL VARICES
C0192316|T060||CPT|INJECTION OF OESOPHAGEAL VARICES BY ENDOSCOPY
C0192316|T060||CPT|INJECTION OF SCLEROSING AGENT INTO OESOPHAGEAL VARICES BY ENDOSCOPY
C0192316|T060||CPT|INJECTION OF VARICOSE VEINS OF OESOPHAGUS BY ENDOSCOPY
C0192316|T060||CPT|OESOPHAGOSCOPY FOR INJECTION OF OESOPHAGEAL VARICES
C0192316|T060||CPT|ESOPHAGOSCOPY FOR INJECTION OF ESOPHAGEAL VARICES 
C0192316|T060||CPT|INJECTION OF ESOPHAGEAL VARICES BY ENDOSCOPIC APPROACH
C2732453|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH INSERTION OF GUIDE WIRE AND DILATION OF ESOPHAGUS 
C2732453|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY WITH INSERTION OF GUIDE WIRE AND DILATION OF OESOPHAGUS
C2732453|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH INSERTION OF GUIDE WIRE AND DILATION OF ESOPHAGUS
C2122145|T060||CPT|FIBEROPTIC DUODENOSCOPY 
C2122145|T060||CPT|FIBEROPTIC DUODENOSCOPY
C2122145|T060||CPT|FIBEROPTIC EXAMINATIONS DUODENOSCOPY
C0472844|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY 
C0472844|T060||CPT|FIBEROPTIC EXAMINATIONS ESOPHAGOSCOPY
C0472844|T060||CPT|FIBEROPTIC ESOPHAGOSCOPY
C0472844|T060||CPT|FIBREOPTIC OESOPHAGOSCOPY
C0472844|T060||CPT|FLEXIBLE ESOPHAGOSCOPY
C0472844|T060||CPT|FLEXIBLE OESOPHAGOSCOPY
C0017195|T060||CPT|GASTROSCOPIES
C0017195|T060||CPT|GASTROSCOPY
C0017195|T060||CPT|FIBEROPTIC EXAMINATIONS GASTROSCOPY
C0017195|T060||CPT|GASTROSCOPY 
C0017195|T060||CPT|ENDOSCOPY OF STOMACH
C0017195|T060||CPT|ENDOSCOPY OF STOMACH 
C0017195|T060||CPT|UPPER ENDOSCOPY
C0017195|T060||CPT|ENDOSCOPY OF STOMACH, NOS
C0017195|T060||CPT|GASTROSCOPY, NOS
C2207161|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY W/ DIRECTED SUBMUCOUSAL INJECTION
C2207161|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH DIRECTED SUBMUCOUSAL INJECTION 
C2207161|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH DIRECTED SUBMUCOUSAL INJECTION
C2207161|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH DIRECTED SUBMUCOUSAL INJECTION(S)
C0192674|T060|43239|CPT|ESOPHAGOGASTRODUODENOSCOPY WITH BIOPSY |BIOPSY OF THE ESOPHAGUS, STOMACH, AND/OR UPPER SMALL BOWEL USING AN ENDOSCOPE
C0192674|T060|43239|CPT|ESOPHAGOGASTRODUODENOSCOPY WITH BIOPSY|BIOPSY OF THE ESOPHAGUS, STOMACH, AND/OR UPPER SMALL BOWEL USING AN ENDOSCOPE
C0192674|T060|43239|CPT|UPPER GASTROINTESTINAL ENDOSCOPY WITH BIOPSY|BIOPSY OF THE ESOPHAGUS, STOMACH, AND/OR UPPER SMALL BOWEL USING AN ENDOSCOPE
C0192674|T060|43239|CPT|BIOPSY OF THE ESOPHAGUS, STOMACH, AND/OR UPPER SMALL BOWEL USING AN ENDOSCOPE|BIOPSY OF THE ESOPHAGUS, STOMACH, AND/OR UPPER SMALL BOWEL USING AN ENDOSCOPE
C0192674|T060|43239|CPT|UPPER GASTROINTESTINAL ENDOSCOPY; BIOPSY|BIOPSY OF THE ESOPHAGUS, STOMACH, AND/OR UPPER SMALL BOWEL USING AN ENDOSCOPE
C0399616|T060||CPT|GASTRESOPHAGOSCOPY VIA GASTROTOMY
C0399616|T060||CPT|GASTROESOPHAGOSCOPY VIA GASTROTOMY
C0399616|T060||CPT|GASTROOESOPHAGOSCOPY VIA GASTROTOMY
C0399616|T060||CPT|ESOPHAGOGASTROSCOPY VIA GASTROTOMY
C0399616|T060||CPT|OESOPHAGOGASTROSCOPY VIA GASTROTOMY
C0399616|T060||CPT|OESOPHAGOGASTROSCOPY VIA GASTROTOMY 
C0399616|T060||CPT|ESOPHAGOGASTROSCOPY VIA GASTROTOMY 
C0192470|T060||CPT|ESOPHAGOGASTROSCOPY THROUGH STOMA
C0192470|T060||CPT|OESOPHAGOGASTROSCOPY THROUGH STOMA
C0192470|T060||CPT|ESOPHAGOGASTROSCOPY THROUGH STOMA 
C0472851|T060||CPT|RIGID ESOPHAGOSCOPY 
C0472851|T060||CPT|RIGID ESOPHAGOSCOPY
C0472851|T060||CPT|RIGID OESOPHAGOSCOPY
C0472851|T060||CPT|RIGID ESOPHAGOSCOPY 
C0192656|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY THROUGH STOMA
C0192656|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY THROUGH STOMA
C0192656|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY THROUGH STOMA 
C0192656|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY THROUGH STOMA  [AMBIGUOUS]
C2960085|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF POLYP OF ESOPHAGUS
C2960085|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF POLYP OF OESOPHAGUS
C2960085|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND POLYPECTOMY OF OESOPHAGUS
C2960085|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND POLYPECTOMY OF ESOPHAGUS
C2960085|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF POLYP OF ESOPHAGUS 
C2960784|T060||CPT|ENDOSCOPY AND BIOPSY OF UPPER GASTROINTESTINAL TRACT 
C2960784|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND BIOPSY
C2960784|T060||CPT|ENDOSCOPY AND BIOPSY OF UPPER GASTROINTESTINAL TRACT
C2960784|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND BIOPSY
C2959366|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND DILATION OF ESOPHAGEAL STRICTURE 
C2959366|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND DILATION OF OESOPHAGEAL STRICTURE
C2959366|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND DILATION OF ESOPHAGEAL STRICTURE
C2959366|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND DILATION OF ESOPHAGEAL STRICTURE
C2959366|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND DILATION OF OESOPHAGEAL STRICTURE
C2959746|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND MUCOSECTOMY OF DUODENUM
C2959746|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF MUCOSA OF DUODENUM 
C2959746|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND MUCOSECTOMY OF DUODENUM
C2959746|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF MUCOSA OF DUODENUM
C2960325|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF MUCOSA OF STOMACH 
C2960325|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF MUCOSA OF STOMACH
C2960325|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND MUCOSECTOMY OF STOMACH
C2960325|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND MUCOSECTOMY OF STOMACH
C2959681|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF POLYP OF DUODENUM
C2959681|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND POLYPECTOMY OF DUODENUM
C2959681|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF POLYP OF DUODENUM 
C2959681|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND POLYPECTOMY OF DUODENUM
C2959668|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND REMOVAL OF FOREIGN BODY FROM ESOPHAGUS
C2959668|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND REMOVAL OF FOREIGN BODY FROM ESOPHAGUS 
C2959668|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND REMOVAL OF FOREIGN BODY FROM OESOPHAGUS
C2959668|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND REMOVAL OF FOREIGN BODY FROM OESOPHAGUS
C2959668|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND REMOVAL OF FOREIGN BODY FROM ESOPHAGUS
C2960120|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND INSERTION OF OESOPHAGEAL STENT
C2960120|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INSERTION OF ESOPHAGEAL STENT
C2960120|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INSERTION OF OESOPHAGEAL STENT
C2960120|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND INSERTION OF ESOPHAGEAL STENT
C2960120|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INSERTION OF ESOPHAGEAL STENT 
C2960528|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND DILATION OF GASTRIC CARDIA
C2960528|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND DILATION OF GASTRIC CARDIA
C2960528|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND DILATION OF GASTRIC CARDIA
C2960528|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND DILATION OF GASTRIC CARDIA 
C2960061|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND TATTOOING 
C2960061|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND TATTOOING
C2960061|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND TATTOOING
C2960061|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND TATTOOING
C2959967|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND DILATION OF GASTRIC STOMA
C2959967|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND DILATION OF GASTRIC STOMA 
C2960407|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND INJECTION OF GASTRIC VARICES
C2960407|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INJECTION OF VARIX OF STOMACH 
C2960407|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND INJECTION OF GASTRIC VARICES
C2960407|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INJECTION OF GASTRIC VARICES
C2960407|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INJECTION OF VARIX OF STOMACH
C2959433|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF MUCOSA OF ESOPHAGUS 
C2959433|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF MUCOSA OF OESOPHAGUS
C2959433|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND MUCOSECTOMY OF ESOPHAGUS
C2959433|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF MUCOSA OF ESOPHAGUS
C2959433|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND MUCOSECTOMY OF OESOPHAGUS
C2960354|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF POLYP OF STOMACH 
C2960354|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND POLYPECTOMY OF STOMACH
C2960354|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND EXCISION OF POLYP OF STOMACH
C2960354|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND POLYPECTOMY OF STOMACH
C2959632|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF ESOPHAGUS 
C2959632|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND BANDING OF ESOPHAGEAL VARICES
C2959632|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF OESOPHAGUS
C2959632|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF ESOPHAGEAL VARICES
C2959632|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF OESOPHAGEAL VARICES
C2959632|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF ESOPHAGUS
C2959632|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND BANDING OF OESOPHAGEAL VARICES
C2959721|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INJECTION OF VARIX OF ESOPHAGUS 
C2959721|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND INJECTION OF ESOPHAGEAL VARICES
C2959721|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INJECTION OF ESOPHAGEAL VARICES
C2959721|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INJECTION OF VARIX OF OESOPHAGUS
C2959721|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INJECTION OF OESOPHAGEAL VARICES
C2959721|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND INJECTION OF VARIX OF ESOPHAGUS
C2959721|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND INJECTION OF OESOPHAGEAL VARICES
C2959927|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND BANDING OF GASTRIC VARICES
C2959927|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF STOMACH
C2959927|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF GASTRIC VARICES
C2959927|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND BANDING OF VARIX OF STOMACH 
C2959927|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND BANDING OF GASTRIC VARICES
C2960375|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND LIGATION OF DUODENAL VARICES
C2960375|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND LIGATION OF DUODENAL VARICES
C2960375|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND LIGATION OF VARIX OF DUODENUM 
C2960375|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND LIGATION OF VARIX OF DUODENUM
C2960375|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND LIGATION OF DUODENAL VARICES
C0014873|T060||CPT|ESOPHAGOSCOPIES
C0014873|T060||CPT|ESOPHAGOSCOPY
C0014873|T060||CPT|OESOPHAGOSCOPY
C0014873|T060||CPT|ESOPHAGOSCOPY 
C0014873|T060||CPT|ENDOSCOPY PROCEDURES ON THE ESOPHAGUS
C0014873|T060||CPT|ENDOSCOPIC EXAMINATION OF ESOPHAGUS
C0014873|T060||CPT|ENDOSCOPIC EXAMINATION OF OESOPHAGUS
C0014873|T060||CPT|ENDOSCOPY OF ESOPHAGUS 
C0014873|T060||CPT|ENDOSCOPY OF ESOPHAGUS
C0014873|T060||CPT|ENDOSCOPY OF OESOPHAGUS
C0014873|T060||CPT|ENDOSCOPY OF ESOPHAGUS, NOS
C0014873|T060||CPT|ESOPHAGOSCOPY, NOS
C0014873|T060||CPT|OESOPHAGOSCOPY, NOS
C0192471|T060||CPT|ESOPHAGOGASTROSCOPY OPERATIVE
C0192471|T060||CPT|ESOPHAGOGASTROSCOPY OPERATIVE 
C0192471|T060||CPT|OPERATIVE ESOPHAGOGASTROSCOPY
C0192471|T060||CPT|OPERATIVE OESOPHAGOGASTROSCOPY
C0192471|T060||CPT|OPERATIVE ESOPHAGOGASTROSCOPY 
C0013301|T060||CPT|DUODENOSCOPIES
C0013301|T060||CPT|DUODENOSCOPY
C0013301|T060||CPT|DUODENOSCOPY 
C0013301|T060||CPT|ENDOSCOPY OF DUODENUM
C0013301|T060||CPT|DUODENOSCOPY, NOS
C0013301|T060||CPT|ENDOSCOPY OF DUODENUM, NOS
C0192655|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY OPERATIVE
C0192655|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY OPERATIVE 
C0192655|T060||CPT|OPERATIVE ESOPHAGOGASTRODUODENOSCOPY
C0192655|T060||CPT|OPERATIVE OESOPHAGOGASTRODUODENOSCOPY
C0192655|T060||CPT|OPERATIVE ESOPHAGOGASTRODUODENOSCOPY 
C2095043|T060||CPT|UPPER GASTROINTESTINAL ENDOSCOPY, SIMPLE PRIMARY EXAM
C2095043|T060||CPT|UPPER GASTROINTESTINAL ENDOSCOPY, SIMPLE PRIMARY EXAM 
C2095043|T060||CPT|UPPER GI ENDOSCOPY, SIMPLE PRIMARY EXAM
C2095643|T060|43235|CPT|UPPER GASTROINTESTINAL ENDOSCOPY |DIAGNOSTIC UPPER GASTROINTESTINAL ENDOSCOPY
C2095643|T060|43235|CPT|UPPER GI ENDOSCOPY DIAGNOSTIC|DIAGNOSTIC UPPER GASTROINTESTINAL ENDOSCOPY
C2095643|T060|43235|CPT|UPPER GASTROINTESTINAL DIAGNOSTIC ENDOSCOPY|DIAGNOSTIC UPPER GASTROINTESTINAL ENDOSCOPY
C2095643|T060|43235|CPT|UPPER GASTROINTESTINAL DIAGNOSTIC ENDOSCOPY |DIAGNOSTIC UPPER GASTROINTESTINAL ENDOSCOPY
C2095643|T060|43235|CPT|DIAGNOSTIC UPPER GASTROINTESTINAL ENDOSCOPY|DIAGNOSTIC UPPER GASTROINTESTINAL ENDOSCOPY
C3507762|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH OPTIC ENDOMICROSCOPY
C3507762|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH OPTIC ENDOMICROSCOPY 
C0192466|T060||CPT|OESOPHAGOGASTROSCOPY
C0192466|T060||CPT|ESOPHAGOGASTROSCOPY
C0192466|T060||CPT|ENDOSCOPIC EXAMINATION OF ESOPHAGUS AND STOMACH
C0192466|T060||CPT|ENDOSCOPIC EXAMINATION OF OESOPHAGUS AND STOMACH
C0192466|T060||CPT|ESOPHAGOGASTROSCOPY 
C0192466|T060||CPT|ESOPHAGOGASTROSCOPY 
C3694781|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY TRANSORAL FLEX W/ OPTIC ENDOMICROSCOPY 
C3694781|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY TRANSORAL FLEX W/ OPTIC ENDOMICROSCOPY
C3694780|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY TRANSORAL FLEXIBLE 
C3694780|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY TRANSORAL FLEXIBLE
C3694780|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY, FLEXIBLE, TRANSORAL
C4038699|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY AND DILATATION OF DUODENUM
C4038699|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND DILATATION OF DUODENUM 
C4038699|T060||CPT|ENDOSCOPY OF UPPER GASTROINTESTINAL TRACT AND DILATATION OF DUODENUM
C4038699|T060||CPT|OESOPHAGOGASTRODUODENOSCOPY AND DILATATION OF DUODENUM
C4065150|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH ESOPHAGOGASTRIC FUNDOPLASTY
C4065150|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH ESOPHAGOGASTRIC FUNDOPLASTY 
C0810405|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY (EGD) WITH BIOPSY
C0176784|T060||CPT|EGD WITH CLOSED BIOPSY
C0176784|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY [EGD] WITH CLOSED BIOPSY
C0176784|T060||CPT|ESOPHAGOGASTRODUODENOSCOPY WITH CLOSED BIOPSY
C0176784|T060||CPT|BIOPSY OF ONE OR MORE SITES INVOLVING ESOPHAGUS, STOMACH AND/OR DUODENUM
C0399617|T060||CPT|DIAGNOSTIC GASTROSCOPY VIA STOMA
C0399617|T060||CPT|DIAGNOSTIC GASTROSCOPY VIA STOMA 
C0009556|T060||CPT|COMPLETE COLONOSCOPY
C0009556|T060||CPT|COMPLETE COLONOSCOPY 
C0009556|T060||CPT|TOTAL COLONOSCOPY
C0009556|T060||CPT|TOTAL COLONOSCOPY 
C0192910|T060|44390|CPT|COLONOSCOPY STOMA W/RMVL FOREIGN BODY|COLONOSCOPY STOMA W/RMVL FOREIGN BODY
C0192910|T060|44390|CPT|COLONOSCOPY THROUGH STOMA WITH REMOVAL OF FOREIGN BODY|COLONOSCOPY STOMA W/RMVL FOREIGN BODY
C0192910|T060|44390|CPT|RETIRED PROCEDURE  [P1-57731]|COLONOSCOPY STOMA W/RMVL FOREIGN BODY
C0192910|T060|44390|CPT|RETIRED PROCEDURE [P1-57731]|COLONOSCOPY STOMA W/RMVL FOREIGN BODY
C0192910|T060|44390|CPT|COLONOSCOPY THROUGH STOMA; WITH REMOVAL OF FOREIGN BODY(S)|COLONOSCOPY STOMA W/RMVL FOREIGN BODY
C0192910|T060|44390|CPT|COLONOSCOPY FOR FOREIGN BODY|COLONOSCOPY STOMA W/RMVL FOREIGN BODY
C0016234|T060||CPT|FLEXIBLE FIBEROPTIC SIGMOIDOSCOPY
C0016234|T060||CPT|FIBEROPTIC EXAMINATIONS SIGMOIDOSCOPY
C0016234|T060||CPT|FIBEROPTIC SIGMOIDOSCOPY 
C0016234|T060||CPT|FIBEROPTIC SIGMOIDOSCOPY
C0016234|T060||CPT|FIBEROPTIC SIGMOIDOSCOPY 
C0016234|T060||CPT|FLEXIBLE SIGMOIDOSCOPY
C0016234|T060||CPT|SIGMOIDOSCOPY, FLEXIBLE
C0016234|T060||CPT|FIBREOPTIC SIGMOIDOSCOPY
C0016234|T060||CPT|FS - FLEXIBLE SIGMOIDOSCOPY
C0016234|T060||CPT|FOS - FIBEROPTIC SIGMOIDOSCOPY
C0016234|T060||CPT|FOS - FIBREOPTIC SIGMOIDOSCOPY
C0016234|T060||CPT|FLEXIBLE FIBEROPTIC SIGMOIDOSCOPY 
C0016234|T060||CPT|FLEXIBLE FIBREOPTIC SIGMOIDOSCOPY
C0372134|T060|45379|CPT|FLEXIBLE COLONOSCOPY PROXIMAL TO SPLENIC FLEXURE WITH REMOVAL OF FOREIGN BODY|COLONOSCOPY W/FB REMOVAL
C0372134|T060|45379|CPT|COLONOSCOPY, FLEXIBLE; WITH REMOVAL OF FOREIGN BODY(S)|COLONOSCOPY W/FB REMOVAL
C0372134|T060|45379|CPT|COLONOSCOPY FLX W/REMOVAL OF FOREIGN BODY(S)|COLONOSCOPY W/FB REMOVAL
C0372134|T060|45379|CPT|COLONOSCOPY W/FB REMOVAL|COLONOSCOPY W/FB REMOVAL
C0192899|T060||CPT|COLONOSCOPY WITH RIGID SIGMOIDOSCOPE THROUGH COLOTOMY 
C0192899|T060||CPT|COLONOSCOPY WITH RIGID SIGMOIDOSCOPE THROUGH COLOTOMY
C0192901|T060||CPT|COLONOSCOPY (FIBEROPTIC) WITH BIOPSY
C0192901|T060||CPT|FIBEROPTIC COLONOSCOPY WITH BIOPSY 
C0192901|T060||CPT|FIBEROPTIC COLONOSCOPY WITH BIOPSY
C0192901|T060||CPT|FIBREOPTIC COLONOSCOPY WITH BIOPSY
C0192909|T060||CPT|FIBEROPTIC COLONOSCOPY VIA COLOSTOMY 
C0192909|T060||CPT|FIBEROPTIC COLONOSCOPY VIA COLOSTOMY
C0192909|T060||CPT|FIBEROPTIC EXAMINATIONS COLONOSCOPY VIA COLOSTOMY
C0192909|T060||CPT|FIBEROPTIC COLONOSCOPY THROUGH COLOSTOMY
C0192909|T060||CPT|ENDOSCOPY OF COLON THROUGH ARTIFICIAL STOMA
C0192909|T060||CPT|COLONOSCOPY THROUGH ARTIFICIAL STOMA
C0192909|T060||CPT|FIBEROPTIC COLONOSCOPY THROUGH COLOSTOMY 
C0192909|T060||CPT|FIBREOPTIC COLONOSCOPY THROUGH COLOSTOMY
C0037075|T060||CPT|PROCTOSIGMOIDOSCOPIES
C0037075|T060||CPT|PROCTOSIGMOIDOSCOPY
C0037075|T060||CPT|SIGMOIDOSCOPIES
C0037075|T060||CPT|SIGMOIDOSCOPY
C0037075|T060||CPT|SIGMOIDOSCOPY 
C0037075|T060||CPT|SIGGY - SIGMOIDOSCOPY
C0037075|T060||CPT|SIGY - SIGMOIDOSCOPY
C0037075|T060||CPT|SIGMOIDOSCOPY, NOS
C0009378|T060|1007622|CPT|COLONOSCOPIES|ENDOSCOPY PROCEDURES ON THE RECTUM
C0009378|T060|1007622|CPT|COLONOSCOPY|ENDOSCOPY PROCEDURES ON THE RECTUM
C0009378|T060|1007622|CPT|COLONOSCOPY |ENDOSCOPY PROCEDURES ON THE RECTUM
C0009378|T060|1007622|CPT|COLONOSCOPY |ENDOSCOPY PROCEDURES ON THE RECTUM
C0009378|T060|1007622|CPT|ENDOSCOPY PROCEDURES ON THE RECTUM|ENDOSCOPY PROCEDURES ON THE RECTUM
C0009378|T060|1007622|CPT|ENDOSCOPIC EXAMINATION OF COLON|ENDOSCOPY PROCEDURES ON THE RECTUM
C0009378|T060|1007622|CPT|ENDOSCOPY OF COLON|ENDOSCOPY PROCEDURES ON THE RECTUM
C0009378|T060|1007622|CPT|COLONOSCOPY, NOS|ENDOSCOPY PROCEDURES ON THE RECTUM
C0009378|T060|1007622|CPT|ENDOSCOPY OF COLON, NOS|ENDOSCOPY PROCEDURES ON THE RECTUM
C0009378|T060|1007622|CPT|COLONOSCOPY [AMBIGUOUS]|ENDOSCOPY PROCEDURES ON THE RECTUM
C0751041|T060||CPT|SURG PROCEDURES COLONOSCOPIC
C0751041|T060||CPT|SURG COLONOSCOPIC
C0751041|T060||CPT|COLONOSCOPIC SURG PROCEDURES
C0751041|T060||CPT|COLONOSCOPIC SURG
C0751041|T060||CPT|COLONOSCOPIC SURGICAL PROCEDURE
C0751041|T060||CPT|PROCEDURE, COLONOSCOPIC SURGICAL
C0751041|T060||CPT|PROCEDURES, COLONOSCOPIC SURGICAL
C0751041|T060||CPT|SURGICAL PROCEDURE, COLONOSCOPIC
C0751041|T060||CPT|COLONOSCOPIC SURGERIES
C0751041|T060||CPT|SURGERIES, COLONOSCOPIC
C0751041|T060||CPT|COLONOSCOPIC SURGERY
C0751041|T060||CPT|SURGICAL PROCEDURES, COLONOSCOPIC
C0751041|T060||CPT|SURGERY, COLONOSCOPIC
C0751041|T060||CPT|COLONOSCOPIC SURGICAL PROCEDURES
C2732814|T060||CPT|COLONOSCOPY THROUGH COLOSTOMY WITH ENDOSCOPIC BIOPSY OF COLON
C2732814|T060||CPT|COLONOSCOPY THROUGH COLOSTOMY WITH ENDOSCOPIC BIOPSY OF COLON 
C2732814|T060||CPT|COLONOSCOPY VIA COLOSTOMY WITH ENDOSCOPIC BIOPSY 
C2732814|T060||CPT|COLONOSCOPY VIA COLOSTOMY WITH ENDOSCOPIC BIOPSY
C1882982|T060||CPT|SCREENING COLONOSCOPY
C1882982|T060||CPT|SCREENING COLONOSCOPY 
C1882982|T060||CPT|SCREENING COLONOSCOPY NOS
C2960146|T060||CPT|COLONOSCOPY AND EXCISION OF MUCOSA OF COLON
C2960146|T060||CPT|COLONOSCOPY AND EXCISION OF MUCOSA OF COLON 
C2960146|T060||CPT|COLONOSCOPY AND COLONIC MUCOSECTOMY
C2960146|T060||CPT|COLONOSCOPY WITH EXCISION OF MUCOSA OF COLON 
C2960146|T060||CPT|COLONOSCOPY WITH EXCISION OF MUCOSA OF COLON
C2960408|T060||CPT|COLONOSCOPY AND BIOPSY OF COLON 
C2960408|T060||CPT|COLONOSCOPY AND BIOPSY OF COLON
C2960062|T060||CPT|COLONOSCOPY AND TATTOOING 
C2960062|T060||CPT|COLONOSCOPY AND TATTOOING
C2960062|T060||CPT|COLONOSCOPY (FIBEROPTIC) WITH TATTOOING 
C2960062|T060||CPT|COLONOSCOPY (FIBEROPTIC) WITH TATTOOING
C3274817|T060||CPT|INDEX COLONOSCOPY
C3274817|T060||CPT|BASELINE COLONOSCOPY
C0399623|T060||CPT|INTRAOPERATIVE COLONOSCOPY
C0399623|T060||CPT|INTRAOPERATIVE COLONOSCOPY 
C0399623|T060||CPT|TRANSAB LG BOWEL ENDOSC
C0399623|T060||CPT|OPERATIVE ENDOSCOPY OF COLON
C0399623|T060||CPT|OPERATIVE COLONOSCOPY
C0399623|T060||CPT|TRANSABDOMINAL ENDOSCOPY OF LARGE INTESTINE
C0399623|T060||CPT|INTRAOPERATIVE ENDOSCOPY OF LARGE INTESTINE
C1298662|T060||CPT|ENDOSCOPIC INSERTION OF TEMPORARY COLONIC STENT 
C1298662|T060||CPT|ENDOSCOPIC INSERTION OF TEMPORARY COLONIC STENT
C0585464|T060||CPT|LAPAROSCOPIC RIGHT HEMICOLECTOMY
C0585464|T060||CPT|LAP RIGHT HEMICOLECTOMY
C0585464|T060||CPT|LAPAROSCOPIC-ASSISTED RIGHT COLECTOMY
C0585464|T060||CPT|LAPAROSCOPIC-ASSISTED RIGHT COLECTOMY 
C1298663|T060||CPT|ENDOSCOPIC INSERTION OF PERMANENT COLONIC STENT 
C1298663|T060||CPT|ENDOSCOPIC INSERTION OF PERMANENT COLONIC STENT
C0192929|T060||CPT|PROCTOSIGMOIDOSCOPY WITH BIOPSY
C0192929|T060||CPT|PROCTOSIGMOIDOSCOPY WITH BIOPSY 
C0035622|T060||CPT|RIGID PROCTOSIGMOIDOSCOPY 
C0035622|T060||CPT|RIGID PROCTOSIGMOIDOSCOPY
C0035622|T060||CPT|RIGID PROCTOSIGMOIDOSCPY
C0035622|T060||CPT|PROCTOSIGMOIDOSCOPY.RIGID
C0035622|T060||CPT|PROCTOSIGMOIDOSCOPY, RIGID
C0035622|T060||CPT|RIGID PROCTOSIGMOIDOSCOPY 
C0192927|T060||CPT|PROCTOSIGMOIDOSCOPY BY TRANSABDOMINAL APPROACH
C0192927|T060||CPT|PROCTOSIGMOIDOSCOPY BY TRANSABDOMINAL APPROACH 
C0578726|T060||CPT|ENDOSCOPIC BIOPSY OF LESION OF COLON
C0578726|T060||CPT|ENDOSCOPIC BIOPSY OF LESION OF COLON 
C0192933|T060||CPT|PROCTOSIGMOIDOSCOPY FOR DILATION
C0192933|T060||CPT|PROCTOSIGMOIDOSCOPY FOR DILATION 
C0521258|T060||CPT|LAPAROSCOPIC-ASSISTED LEFT COLECTOMY
C0521258|T060||CPT|LAPAROSCOPIC-ASSISTED LEFT COLECTOMY 
C0192900|T060||CPT|FIBEROPTIC COLONOSCOPY
C0192900|T060||CPT|FIBEROPTIC COLONOSCOPY, NOS
C0192900|T060||CPT|FIBREOPTIC COLONOSCOPY, NOS
C0192900|T060||CPT|FIBEROPTIC COLONOSCOPY 
C0192900|T060||CPT|FIBREOPTIC COLONOSCOPY
C0192900|T060||CPT|COLONOSCOPY 
C0192900|T060||CPT|FIBEROPTIC COLONOSCOPY  [AMBIGUOUS]
C0192900|T060||CPT|FLEXIBLE FIBEROPTIC COLONOSCOPY
C2095474|T060||CPT|COMPLETE COLONOSCOPY OF HEPATIC FLEXURE 
C2095474|T060||CPT|COMPLETE COLONOSCOPY OF HEPATIC FLEXURE
C2095866|T060||CPT|COMPLETE COLONOSCOPY OF SIGMOID COLON WITH DILATION 
C2095866|T060||CPT|COMPLETE COLONOSCOPY OF SIGMOID COLON WITH DILATION
C2095475|T060||CPT|COMPLETE COLONOSCOPY OF TRANSVERSE COLON 
C2095475|T060||CPT|COMPLETE COLONOSCOPY OF TRANSVERSE COLON
C2095473|T060||CPT|COMPLETE COLONOSCOPY OF ASCENDING COLON
C2095473|T060||CPT|COMPLETE COLONOSCOPY OF ASCENDING COLON 
C2095478|T060||CPT|COMPLETE COLONOSCOPY OF SIGMOID COLON
C2095478|T060||CPT|COMPLETE COLONOSCOPY OF SIGMOID COLON 
C2095476|T060||CPT|COMPLETE COLONOSCOPY OF SPLENIC FLEXURE 
C2095476|T060||CPT|COMPLETE COLONOSCOPY OF SPLENIC FLEXURE
C2095477|T060||CPT|COMPLETE COLONOSCOPY OF DESCENDING COLON
C2095477|T060||CPT|COMPLETE COLONOSCOPY OF DESCENDING COLON 
C0588165|T060||CPT|CHECK COLONOSCOPY 
C0588165|T060||CPT|CHECK COLONOSCOPY
C0588165|T060||CPT|COLONOSCOPY CHECK
C0588165|T060||CPT|CHECK COLONOSCOPY 
C0554063|T060||CPT|THERAPEUTIC COLONOSCOPY
C0554063|T060||CPT|COLONOSCOPY THERAPEUTIC
C0554063|T060||CPT|THERAPEUTIC COLONOSCOPY 
C0554063|T060||CPT|THERAPEUTIC COLONOSCOPY 
C0399622|T060||CPT|OPEN COLONOSCOPY 
C0399622|T060||CPT|OPEN COLONOSCOPY
C0399622|T060||CPT|OPEN COLONOSCOPY 
C3869456|T060|1022231|CPT|COLONOSCOPY, FLEXIBLE|COLONOSCOPY, FLEXIBLE
C4040527|T060||CPT|COLONOSCOPY AND DILATATION OF STRICTURE OF COLON
C4040527|T060||CPT|COLONOSCOPY AND DILATATION OF STRICTURE OF COLON 
C4039452|T060||CPT|COLONOSCOPY USING X-RAY GUIDANCE
C4039452|T060||CPT|COLONOSCOPY USING X-RAY GUIDANCE 
C4038675|T060||CPT|COLONOSCOPY USING FLUOROSCOPIC GUIDANCE
C4038675|T060||CPT|FLUOROSCOPY GUIDED COLONOSCOPY
C4038675|T060||CPT|COLONOSCOPY USING FLUOROSCOPIC GUIDANCE 
C0400018|T060||CPT|DIAGNOSTIC COLONOSCOPY
C0400018|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION ON COLON
C0400018|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF COLON NOS
C0400018|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF COLON NOS 
C0400018|T060||CPT|DIAGNOSTIC ENDOSCOPY OF COLON
C0400018|T060||CPT|COLON ENDOSCOPY 
C0400018|T060||CPT|DIAGNOSTIC ENDOSCOPY OF COLON 
C0400018|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION ON COLON 
C0399625|T060||CPT|COLONOSCOPY (FIBEROPTIC) LIMITED
C0399625|T060||CPT|LIMITED COLONOSCOPY (FIBEROPTIC) 
C0399625|T060||CPT|LIMITED COLONOSCOPY (FIBEROPTIC)
C0399625|T060||CPT|LIMITED COLONOSCOPY
C0399625|T060||CPT|LIMITED COLONOSCOPY 
C0863836|T060||CPT|ENDOSCOPY OF DESCENDING COLON
C1960976|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF COLONIC POUCH AND BIOPSY OF COLONIC POUCH USING FIBEROPTIC SIGMOIDOSCOPE 
C1960976|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF COLONIC POUCH AND BIOPSY OF COLONIC POUCH USING FIBEROPTIC SIGMOIDOSCOPE
C1960976|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF COLONIC POUCH AND BIOPSY OF COLONIC POUCH USING FIBREOPTIC SIGMOIDOSCOPE
C1960975|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF COLONIC POUCH AND BIOPSY OF COLONIC POUCH USING COLONOSCOPE 
C1960975|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF COLONIC POUCH AND BIOPSY OF COLONIC POUCH USING COLONOSCOPE
C1960975|T060||CPT|COLONOSCOPY (FIBEROPTIC) OF COLONIC POUCH WITH BIOPSY
C1960975|T060||CPT|COLONOSCOPY (FIBEROPTIC) OF COLONIC POUCH WITH BIOPSY 
C1960974|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF COLONIC POUCH AND BIOPSY OF COLONIC POUCH USING RIGID SIGMOIDOSCOPE 
C1960974|T060||CPT|DIAGNOSTIC ENDOSCOPIC EXAMINATION OF COLONIC POUCH AND BIOPSY OF COLONIC POUCH USING RIGID SIGMOIDOSCOPE
