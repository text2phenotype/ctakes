C1849687|T033||SNOMEDCT_US|LIVER BIOPSY SHOWS NORMAL NUMBERS OF ENLARGED PEROXISOMES
C1856310|T033||SNOMEDCT_US|LIVER BIOPSY SHOWS DIFFUSE INTERSTITIAL FIBROSIS
C1857356|T033||SNOMEDCT_US|LIVER BIOPSY SHOWS INCREASED LIPID DROPLETS (MICROVESICULAR STEATOSIS)
C1857367|T033||SNOMEDCT_US|LIVER BIOPSY SHOWS INCREASED LIPID DROPLETS AND ABNORMAL MITOCHONDRIA
C2021366|T033||SNOMEDCT_US|LIVER BIOPSY IRON (UG/100 MG OF DRY WEIGHT)
# C2368138|T033||SNOMEDCT_US|NOT THE SAME
C2674614|T033||SNOMEDCT_US|LIVER BIOPSY SHOWS RED AUTOFLUORESCENCE AND NEEDLE-LIKE CYTOPLASMIC INCLUSION BODIES
C2748696|T033||SNOMEDCT_US|LIVER BIOPSY SHOWS DUCTAL PROLIFERATION
C2751577|T033||SNOMEDCT_US|LIVER BIOPSY DURING ACUTE EPISODE SHOWS VARIABLE PORTAL AND SINUSOIDAL FIBROSIS
C3277942|T033||SNOMEDCT_US|LIVER BIOPSY SHOWS PORTAL AND/OR BRIDGING FIBROSIS
C4273160|T033||SNOMEDCT_US|BILE DUCT BIOPSY SHOWED PAUCITY OF DUCTS
C3899974|T033||SNOMEDCT_US|BCLC STAGE
C3897124|T033||SNOMEDCT_US|BCLC STAGE A HEPATOCELLULAR CARCINOMA
C3897124|T033||SNOMEDCT_US|BCLC STAGE A
C3898888|T033||SNOMEDCT_US|HCC BY BCLC STAGE
C3898888|T033||SNOMEDCT_US|BCLC HEPATOCELLULAR CARCINOMA
C3898888|T033||SNOMEDCT_US|BCLC STAGE HEPATOCELLULAR CARCINOMA
C3898888|T033||SNOMEDCT_US|HEPATOCELLULAR CARCINOMA BY BCLC STAGE
C3899975|T033||SNOMEDCT_US|BCLC STAGE D HEPATOCELLULAR CARCINOMA
C3899975|T033||SNOMEDCT_US|BCLC STAGE D HCC
C3899977|T033||SNOMEDCT_US|BCLC STAGE C HEPATOCELLULAR CARCINOMA
C3899975|T033||SNOMEDCT_US|BCLC STAGE C HCC
C3899979|T033||SNOMEDCT_US|BCLC STAGE B HEPATOCELLULAR CARCINOMA
C3899975|T033||SNOMEDCT_US|BCLC STAGE B HCC
C3899981|T033||SNOMEDCT_US|BCLC STAGE A ADULT HEPATOCELLULAR CARCINOMA
C3899975|T033||SNOMEDCT_US|BCLC STAGE A HCC
C3899982|T033||SNOMEDCT_US|BCLC STAGE 0 HEPATOCELLULAR CARCINOMA
C3899975|T033||SNOMEDCT_US|BCLC STAGE 0 HCC
C3899976|T033||SNOMEDCT_US|BCLC STAGE D ADULT HEPATOCELLULAR CARCINOMA
C3899976|T033||SNOMEDCT_US|BCLC STAGE D ADULT HCC
C3899978|T033||SNOMEDCT_US|BCLC STAGE C ADULT HEPATOCELLULAR CARCINOMA
C3899978|T033||SNOMEDCT_US|BCLC STAGE C ADULT HCC
C3899980|T033||SNOMEDCT_US|BCLC STAGE B ADULT HEPATOCELLULAR CARCINOMA
C3899980|T033||SNOMEDCT_US|BCLC STAGE B ADULT HCC
C3899983|T033||SNOMEDCT_US|BCLC STAGE 0 ADULT HEPATOCELLULAR CARCINOMA
C3899983|T033||SNOMEDCT_US|BCLC STAGE 0 ADULT HCC
C3550399|T033||SNOMEDCT_US|INCREASED IRON DEPOSITION SEEN ON LIVER BIOPSY
C4020697|T033||SNOMEDCT_US|GIANT CELL HEPATITIS ON LIVER BIOPSY
C4314030|T033||SNOMEDCT_US|DUCTAL REACTION SEEN ON LIVER BIOPSY
C1847706|T033||SNOMEDCT_US|ABSENCE OF BETA-UREIDOPROPIONASE ACTIVITY AND PROTEIN IN LIVER BIOPSY
C3899981|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE A ADULT HEPATOCELLULAR CARCINOMA
C3899981|T033||SNOMEDCT_US|BCLC STAGE A ADULT HEPATOCELLULAR CARCINOMA
C3899982|T033||SNOMEDCT_US|BCLC STAGE 0 HEPATOCELLULAR CARCINOMA
C3899982|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE 0 HEPATOCELLULAR CARCINOMA
C3897124|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE A HEPATOCELLULAR CARCINOMA
C3897124|T033||SNOMEDCT_US|BCLC STAGE A HEPATOCELLULAR CARCINOMA
C3899975|T033||SNOMEDCT_US|BCLC STAGE D HEPATOCELLULAR CARCINOMA
C3899975|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE D HEPATOCELLULAR CARCINOMA
C3899977|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE C HEPATOCELLULAR CARCINOMA
C3899977|T033||SNOMEDCT_US|BCLC STAGE C HEPATOCELLULAR CARCINOMA
C3899979|T033||SNOMEDCT_US|BCLC STAGE B HEPATOCELLULAR CARCINOMA
C3899979|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE B HEPATOCELLULAR CARCINOMA
C3899976|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE D ADULT HEPATOCELLULAR CARCINOMA
C3899976|T033||SNOMEDCT_US|BCLC STAGE D ADULT HEPATOCELLULAR CARCINOMA
C3899978|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE C ADULT HEPATOCELLULAR CARCINOMA
C3899978|T033||SNOMEDCT_US|BCLC STAGE C ADULT HEPATOCELLULAR CARCINOMA
C3899980|T033||SNOMEDCT_US|BCLC STAGE B ADULT HEPATOCELLULAR CARCINOMA
C3899980|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE B ADULT HEPATOCELLULAR CARCINOMA
C3899983|T033||SNOMEDCT_US|BARCELONA CLINIC LIVER CANCER STAGE 0 ADULT HEPATOCELLULAR CARCINOMA
C3899983|T033||SNOMEDCT_US|BCLC STAGE 0 ADULT HEPATOCELLULAR CARCINOMA
