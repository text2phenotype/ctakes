# CUI|TUI|CODE|SAB|TEXT|PREF_TEXT
C0000001|T059|1|TEST_VOCAB1|ONE|NUMBER ONE
C0000002|T053|2|TEST_VOCAB2|TWO|NUMBER TWO
C0000003|T034|3|TEST_VOCAB3|THREE|NUMBER THREE
C0000004|T047|4|TEST_VOCAB4|FOUR|NUMBER FOUR
C0000005|T048|5|TEST_VOCAB5|FIVE|NUMBER FIVE