C0150055|T184||CHV|CHRONIC PAIN
C0150055|T184||CHV|CHRONIC PAIN 
C0232491|T184||CHV|CHRONIC ABDOMINAL PAIN
C0457949|T184|0000047258|CHV|CHRONIC LOW BACK PAIN|BACK PAIN LOWER BACK CHRONIC
C0743541|T184||CHV|CHRONIC EPIGASTRIC PAIN
C0267515|T184||CHV|CHRONIC IDIOPATHIC ANAL PAIN
C0267515|T184||CHV|CHRONIC IDIOPATHIC ANAL PAIN 
C2316723|T184||CHV|CHRONIC PAIN DUE TO INJURY 
C2316723|T184||CHV|CHRONIC PAIN DUE TO INJURY
C2316650|T184||CHV|CHRONIC PAIN IN FACE 
C2316650|T184||CHV|CHRONIC FACIAL PAIN
C2316650|T184||CHV|CHRONIC PAIN IN FACE
C0150055|T184||CHV|CHRONIC PAIN
C0150055|T184||CHV|CHRONIC PAIN 
C0150055|T184||CHV|RNDX CHRONIC PAIN 
C0150055|T184||CHV|RNDX CHRONIC PAIN
C0150055|T184||CHV|PAIN;CHRONIC
C0150055|T184||CHV|CHRONIC PAINS
C0150055|T184||CHV|PAINS, CHRONIC
C0150055|T184||CHV|CHRONIC PAIN [DISEASE/FINDING]
C0150055|T184||CHV|PAIN, CHRONIC
C0150055|T184||CHV|CHRONIC PAIN 
C0150055|T184||CHV|CHRONIC; PAIN
C0150055|T184||CHV|PAIN; CHRONIC
C1719393|T184||CHV|CHRONIC PAIN DUE TO TRAUMA
C1719393|T184||CHV|CHRONIC PAIN DUE TO TRAUMA 
C1719393|T184||CHV|CHRONC PAIN D/T TRAUMA
C0404484|T184|0000032600|CHV|CHRONIC PAIN IN FEMALE PELVIS|CHRONIC PELVIC PAIN
C0404484|T184|0000032600|CHV|CHRONIC PELVIC PAIN OF FEMALE |CHRONIC PELVIC PAIN
C0404484|T184|0000032600|CHV|CHRONIC PAIN IN FEMALE PELVIS |CHRONIC PELVIC PAIN
C0404484|T184|0000032600|CHV|CHRONIC PELVIC PAIN|CHRONIC PELVIC PAIN
C0404484|T184|0000032600|CHV|CHRONIC PELVIC PAIN OF FEMALE|CHRONIC PELVIC PAIN
C3178789|T184||CHV|PAINS, WIDESPREAD CHRONIC
C3178789|T184||CHV|CHRONIC PAIN, WIDESPREAD
C3178789|T184||CHV|WIDESPREAD CHRONIC PAINS
C3178789|T184||CHV|PAIN, WIDESPREAD CHRONIC
C3178789|T184||CHV|CHRONIC PAINS, WIDESPREAD
C3178789|T184||CHV|PAIN AMPLIFICATION SYNDROME
C3178789|T184||CHV|AMPLIFIED MUSCULOSKELETAL PAIN SYNDROME
C3178789|T184||CHV|CHRONIC WIDESPREAD PAIN
C3178789|T184||CHV|WIDESPREAD CHRONIC PAIN
C3714625|T184||CHV|NEUROPATHIC PAIN
C3714625|T184||CHV|NEUROPATHIC PAIN 
C0478148|T184||CHV|OTHER CHRONIC PAIN
C0478148|T184||CHV|CHRONIC PAIN NEC
C0478148|T184||CHV|[X]OTHER CHRONIC PAIN
C0478148|T184||CHV|OTHER CHRONIC PAIN 
C0478148|T184||CHV|[X]OTHER CHRONIC PAIN 
C0478148|T184||CHV|[X]OTHER CHRONIC PAIN (CONTEXT-DEPENDENT CATEGORY)
C1740831|T184||CHV|CHRONIC CHEST PAIN
C1740831|T184||CHV|CHRONIC CHEST PAIN 
C3649719|T184||CHV|CHRONIC POST-PROCEDURAL PAIN
C3649719|T184||CHV|CHRONIC POST-PROCEDURAL PAIN 
C3649719|T184||CHV|CHRONIC PAIN POST-PROCEDURAAL
C3662083|T184||CHV|CHRONIC PAIN IN MALE PELVIS 
C3662083|T184||CHV|CHRONIC PAIN IN MALE PELVIS
C3662095|T184||CHV|CHRONIC PAIN IN COCCYX FOR MORE THAN THREE MONTHS 
C3662095|T184||CHV|CHRONIC PAIN IN COCCYX FOR MORE THAN THREE MONTHS
C3662064|T184||CHV|CHRONIC NONMALIGNANT PAIN
C3662064|T184||CHV|CHRONIC NONMALIGNANT PAIN 
C3662093|T184||CHV|CHRONIC PAIN DUE TO MALIGNANCY
C3662093|T184||CHV|CHRONIC PAIN DUE TO MALIGNANCY 
C3662084|T184||CHV|CHRONIC THORACIC BACK PAIN 
C3662084|T184||CHV|CHRONIC THORACIC BACK PAIN
C2074900|T184||CHV|CHRONIC POSTOPERATIVE PAIN 
C2074900|T184||CHV|CHRONIC POSTOPERATIVE PAIN
C2074900|T184||CHV|CHRONIC POSTOPERATIVE PAIN 
C0746815|T184|0000047879|CHV|CHRONIC NECK PAIN |CHRONIC CERVICAL PAIN
C0746815|T184|0000047879|CHV|CHRONIC NECK PAIN|CHRONIC CERVICAL PAIN
C0231385|T184||CHV|ALTERATION IN COMFORT: CHRONIC PAIN
C0231385|T184||CHV|ALTERATION IN COMFORT: CHRONIC PAIN 
C0232491|T184||CHV|ABDOMINAL PAIN CHRONIC / CONSTANT
C0232491|T184||CHV|CHRONIC ABDOMINAL PAIN
C0232491|T184||CHV|CHRONIC ABDOMINAL PAIN 
C0232491|T184||CHV|CHRONIC/CONSTANT ABDOMINAL PAIN
C0232491|T184||CHV|CHRONIC ABDOMINAL PAIN 
C0686729|T184||CHV|GENERALIZED CHRONIC BODY ACHES
C0686729|T184||CHV|GENERALIZED CHRONIC BODY PAINS
C0686729|T184||CHV|GENERALISED CHRONIC BODY ACHES
C0686729|T184||CHV|GENERALISED CHRONIC BODY PAINS
C0686729|T184||CHV|GENERALIZED CHRONIC BODY PAINS 
C1333034|T184||CHV|CHRONIC CANCER PAIN
C1719710|T184||CHV|CHRONIC POST-THORACOTOMY PAIN
C1719710|T184||CHV|CHRONIC POST-THORACOTOMY PAIN 
C1719710|T184||CHV|CHRON POST-THORACOT PAIN
C1719394|T184||CHV|OTHER CHRONIC POSTOPERATIVE PAIN
C1719394|T184||CHV|CHRONIC POSTOP PAIN NEC
C1960183|T184||CHV|CHRONIC VAGINAL PAIN
C1960183|T184||CHV|CHRONIC VAGINAL PAIN 
C1960183|T184||CHV|CHRONIC PAIN IN VAGINA
C0476481|T184||CHV|CHRONIC INTRACTABLE PAIN
C0476481|T184||CHV|[D]CHRONIC INTRACTABLE PAIN (CONTEXT-DEPENDENT CATEGORY)
C0476481|T184||CHV|[D]CHRONIC INTRACTABLE PAIN 
C0476481|T184||CHV|[D]CHRONIC INTRACTABLE PAIN
C0476481|T184||CHV|CHRONIC INTRACTABLE PAIN 
C0476481|T184||CHV|PAIN; CHRONIC, INTRACTABLE
C2919655|T184||CHV|ACUTE EXACERBATION OF CHRONIC ABDOMINAL PAIN 
C2919655|T184||CHV|ACUTE EXACERBATION OF CHRONIC ABDOMINAL PAIN
C2074609|T184||CHV|CHRONIC ABDOMINAL PAIN FOR MORE THAN THREE MONTHS 
C2074609|T184||CHV|CHRONIC / CONSTANT ABDOMINAL PAIN FOR MORE THAN 3 MONTHS
C2074609|T184||CHV|CHRONIC ABDOMINAL PAIN FOR MORE THAN THREE MONTHS
C2074609|T184||CHV|CHRONIC/CONSTANT ABDOMINAL PAIN FOR MORE THAN THREE MONTHS
C0400882|T184||CHV|CHRONIC NONSPECIFIC ABDOMINAL PAIN
C0400882|T184||CHV|CHRONIC NONSPECIFIC ABDOMINAL PAIN 
C0457949|T184|0000047258|CHV|LOWER BACK PAIN CHRONIC|BACK PAIN LOWER BACK CHRONIC
C0457949|T184|0000047258|CHV|CHRONIC LOWER BACK PAIN |BACK PAIN LOWER BACK CHRONIC
C0457949|T184|0000047258|CHV|CHRONIC LOWER BACK PAIN|BACK PAIN LOWER BACK CHRONIC
C0457949|T184|0000047258|CHV|PAIN;BACK LOW;CHRONIC|BACK PAIN LOWER BACK CHRONIC
C0457949|T184|0000047258|CHV|CHRONIC LOW BACK PAIN |BACK PAIN LOWER BACK CHRONIC
C0457949|T184|0000047258|CHV|CHRONIC LOW BACK PAIN|BACK PAIN LOWER BACK CHRONIC
C0457949|T184|0000047258|CHV|CLBP - CHRONIC LOW BACK PAIN|BACK PAIN LOWER BACK CHRONIC
C0457949|T184|0000047258|CHV|CHRONIC LOW BACK PAIN |BACK PAIN LOWER BACK CHRONIC
C0743541|T184||CHV|CHRONIC EPIGASTRIC PAIN
