C0004002|T034||LNC|ASPARTATE TRANSAMINASE
C0201899|T034||LNC|ASPARTATE AMINOTRANSFERASE MEASUREMENT
C0684153|T034||LNC|GLUTAMATE OXALOACETATE TRANS 002
C0684153|T034||LNC|ASPARTATE AMINOTRANSFERASE, MITOCHONDRIAL [CHEMICAL/INGREDIENT]
C0684153|T034||LNC|LIVER SPECIFIC AST, BUT NOT THE MOST COMMONLY MEASURED ??INCLUDE?
C0684153|T034||LNC|ASPARTATE AMINOTRANSFERASE, MITOCHONDRIAL
C0684153|T034||LNC|AMINOTRANSFERASE, MITOCHONDRIAL ASPARTATE
C0684153|T034||LNC|GLUTAMATE OXALOACETATE TRANSAMINASE 2
C0684153|T034||LNC|MITOCHONDRIAL ASPARTATE AMINOTRANSFERASE
C0684153|T034||LNC|OXALOACETATE TRANSAMINASE-2, GLUTAMATE
C0684153|T034||LNC|TRANSAMINASE-2, GLUTAMATE OXALOACETATE
C0684153|T034||LNC|EC 2.6.1.1
C0684153|T034||LNC|ASPARTATE AMINOTRANSFERASE 2
C0684153|T034||LNC|MASPAT
C0684153|T034||LNC|TRANSAMINASE A
C0684153|T034||LNC|GOT2
C0684153|T034||LNC|MITOCHONDRIAL GLUTAMIC-OXALOACETIC TRANSAMINASE 2
C0949643|T034||LNC|EC 2.6.1.1
C0949643|T034||LNC|TRANSAMINASE A
C0004002|T034||LNC|AMINOTRANSFERASE, ASPARTATE
C0004002|T034||LNC|AMINOTRANSFERASE, L-ASPARTATE-2-OXOGLUTARATE
C0004002|T034||LNC|APOAMINOTRANSFERASE, ASPARTATE
C0004002|T034||LNC|ASPARTATE AMINOTRANSFERASE
C0004002|T034||LNC|ASPARTATE TRANSAMINASE
C0004002|T034||LNC|GLUTAMIC-OXALOACETIC TRANSAMINASE
C0004002|T034||LNC|TRANSAMINASE, ASPARTATE
C0004002|T034||LNC|TRANSAMINASE, GLUTAMATE-ASPARTATE
C0004002|T034||LNC|TRANSAMINASE, GLUTAMIC-OXALOACETIC
C0004002|T034||LNC|GLUTAMATE ASPARTATE TRANSAMINASE
C0004002|T034||LNC|GLUTAMIC OXALOACETIC TRANSAMINASE
C0004002|T034||LNC|L ASPARTATE 2 OXOGLUTARATE AMINOTRANSFERASE
C0004002|T034||LNC|L-ASPARTATE:2-OXOGLUTARATE AMINOTRANSAMINASE
C0004002|T034||LNC|GLUTAMIC OXALOACETIC TRANS 000
C0004002|T034||LNC|TRANSAMINASE A
C0004002|T034||LNC|GLUTAMIC ASPARTIC TRANSAMINASE
C0004002|T034||LNC|ASPARTATE AMINOTRANSFERASES
C0004002|T034||LNC|GLUTAMATE-ASPARTATE TRANSAMINASE
C0004002|T034||LNC|L-ASPARTATE-2-OXOGLUTARATE AMINOTRANSFERASE
C0004002|T034||LNC|ASPARTATE APOAMINOTRANSFERASE
C0004002|T034||LNC|ASPARTATE AMINOTRANSFERASES [CHEMICAL/INGREDIENT]
C0004002|T034||LNC|AMINOTRANSFERASES, ASPARTATE
C0004002|T034||LNC|ASAT - ASPARTATE AMINOTRANSFERASE
C0004002|T034||LNC|AST - ASPARTATE TRANSAMINASE
# C0004002|T034||LNC|GOT
C0004002|T034||LNC|GLUTAMATE OXALOACETATE TRANSAMINASE
C0004002|T034||LNC|GLUTAMIC-ASPARTIC TRANSAMINASE
C0004002|T034||LNC|L-ASPARTATE:2-OXOGLUTARATE AMINOTRANSFERASE
C0004002|T034||LNC|ASPARTATE AMINOTRANSFERASE 
C1981801|T034|LP45656-3|LNC|ASPARTATE AMINOTRANSFERASE &#X7C; BLD-SER-PLAS|ASPARTATE AMINOTRANSFERASE &#X7C; BLD-SER-PLAS
C0201899|T034||LNC|SERUM SGOT
C0201899|T034||LNC|SERUM AST
C0201899|T034||LNC|ASPARTATE AMINOTRANSFERASE
# C0201899|T034||LNC|GOT
C0201899|T034||LNC|AST
C0201899|T034||LNC|ASPARTATE AMINOTRANSFERASE MEASUREMENT
C0201899|T034||LNC|TRANSFERASE; ASPARTATE AMINO (AST) (SGOT)
C0201899|T034||LNC|TRANSFERASE ASPARTATE AMINO AST SGOT
C0201899|T034||LNC|LIVER ENZYME (SGOT), LEVEL
C0201899|T034||LNC|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T034||LNC|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE (AST) (SGOT)
C0201899|T034||LNC|AST - ASPARTATE TRANSAM SGOT (& LEVEL) 
C0201899|T034||LNC|AST - ASPARTATE TRANSAM SGOT (& LEVEL)
C0201899|T034||LNC|TRANSFERASE (AST) (SGOT)
C0201899|T034||LNC|SGOT
C0201899|T034||LNC|ASPT
C0201899|T034||LNC|ASPARTATE TRANSFERASE
C0201899|T034||LNC|ASP TRANSFERASE
C0201899|T034||LNC|SERUM GLUTAMIC-OXALOACETIC TRANSFERASE
C0201899|T034||LNC|GLUTAMIC-OXALOACETIC TRANSFERASE
C0201899|T034||LNC|SERUM ASPARTATE TRANSAMINASE TEST
C0201899|T034||LNC|AST MEASUREMENT
C0201899|T034||LNC|GLUTAMIC OXALOACETIC TRANSAMINASE MEASUREMENT
C0201899|T034||LNC|GOT MEASUREMENT
C0201899|T034||LNC|SGOT MEASUREMENT
C0201899|T034||LNC|ASPARTATE AMINOTRANSFERASE MEASUREMENT 
C1261155|T034||LNC|AST SERUM MEASUREMENT 
C1261155|T034||LNC|SERUM ASPARTATE TRANSAMINASE MEASUREMENT
C1261155|T034||LNC|SERUM ASPARTATE AMINOTRANSFERASE MEASUREMENT
C1261155|T034||LNC|SERUM SGOT MEASUREMENT
C1261155|T034||LNC|AST SERUM LEVEL
C1261155|T034||LNC|AST SERUM LEVEL 
C1261155|T034||LNC|ASPARTATE AMINOTRANSFERASE (AST) SERUM MEASUREMENT 
C1261155|T034||LNC|ASPARTATE AMINOTRANSFERASE SERUM MEASUREMENT 
C1261155|T034||LNC|ASPARTATE AMINOTRANSFERASE (AST) SERUM MEASUREMENT
C1261155|T034||LNC|ASPARTATE AMINOTRANSFERASE SERUM MEASUREMENT
C1261155|T034||LNC|AST SERUM MEASUREMENT
C1278050|T034||LNC|PLASMA ASPARTATE TRANSAMINASE LEVEL 
C1278050|T034||LNC|PLASMA ASPARTATE TRANSAMINASE LEVEL
C1278050|T034||LNC|PLASMA ASPARTATE TRANSAMINASE MEASUREMENT 
C1278050|T034||LNC|PLASMA ASPARTATE TRANSAMINASE MEASUREMENT
