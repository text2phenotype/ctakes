C1953564|T034|48159-8|LNC|HEP C VIRUS AB|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|HCV AB|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|HCV ANTIBODIES|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|HCV ANTIBODY TEST|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|HEPATITIS C VIRUS (HCV) ANTIBODY|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|HEPATITIS C VIRUS AB|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|HEPATITIS C VIRUS AB SIGNAL|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|HEPATITIS C VIRUS ANTIBODY SIGNAL|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|HEPATITIS C VIRUS ANTIBODY TEST|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|TEST 140659|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|LOINC 48159-8|HCV AB S/CO SERPL IA
C1953564|T034|48159-8|LNC|LNC 48159-8|HCV AB S/CO SERPL IA
