C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC PANEL|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC CHEMICAL PANEL|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|BLOOD TEST, COMPREHENSIVE GROUP OF BLOOD CHEMICALS|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC PANEL |COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC CHEM PANEL|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHEN METABOLIC PANEL|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C2041458|T059||CPT|BLOOD CHEMISTRY TEST PANELS 
C2041458|T059||CPT|BLOOD CHEMISTRY TEST PANELS
C0438930|T059||CPT|CHEM. METABOLIC FUNCTION TESTS
C0438930|T059||CPT|CHEM. METABOLIC FUNCTION TESTS 
C0201838|T059|1011249|CPT|ALBUMIN MEASUREMENT|ALBUMIN
C0201838|T059|1011249|CPT|TEST;ALBUMIN|ALBUMIN
C0201838|T059|1011249|CPT|MEASUREMENT OF ALBUMIN|ALBUMIN
C0201838|T059|1011249|CPT|ALBUMIN|ALBUMIN
C0201838|T059|1011249|CPT|ALB|ALBUMIN
C0201838|T059|1011249|CPT|MICROALBUMIN|ALBUMIN
C0201838|T059|1011249|CPT|ALBUMIN MEASUREMENT |ALBUMIN
C0201838|T059|1011249|CPT|ALBUMIN TEST|ALBUMIN
C0201925|T059|82310|CPT|CALCIUM; TOTAL|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM MEASUREMENT|ASSAY OF CALCIUM
# C0201925|T059|82310|CPT|CA|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM TOTAL|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|MEASUREMENT OF CALCIUM|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM LEVEL|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|LAB-BASED CHEM MEASUREMENTS CALCIUM|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|MEASUREMENT OF CALCIUM |ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CA++|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM MEASUREMENT |ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM MEASUREMENT, NOS|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|ASSAY OF CALCIUM|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM TOTAL EACH TEST|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CA TOT EA.TST|ASSAY OF CALCIUM
C0337438|T059|1011445|CPT|GLUCOSE|GLUCOSE
C0337438|T059|1011445|CPT|GLUCOSE MEASUREMENT|GLUCOSE
C0337438|T059|1011445|CPT|TEST;GLUCOSE|GLUCOSE
C0337438|T059|1011445|CPT|MEASUREMENT OF GLUCOSE|GLUCOSE
C0337438|T059|1011445|CPT|GLUC|GLUCOSE
C0337438|T059|1011445|CPT|GLUCOSE MEASUREMENT |GLUCOSE
C0337438|T059|1011445|CPT|GLUCOSE MEASUREMENT, NOS|GLUCOSE
C0337438|T059|1011445|CPT|GLUCOSE TEST|GLUCOSE
C0201850|T059|84075|CPT|ALKALINE PHOSPHATASE MEASUREMENT|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|PHOSPHATASE, ALKALINE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALP|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|TEST;ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|MEASUREMENT OF ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ASSAY OF PHOSPHATASE ALKALINE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALK PHOSPH|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALK PHOS|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALKALINE PHOSPHATASE MEASUREMENT |ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ASSAY ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALKALINE PHOSPHATASE TEST|ASSAY OF PHOSPHATASE ALKALINE
C0201952|T059|1011335|CPT|CHLORIDE MEASUREMENT|CHLORIDE
C0201952|T059|1011335|CPT|MEASUREMENT OF CHLORIDE|CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE|CHLORIDE
C0201952|T059|1011335|CPT|CL|CHLORIDE
C0201952|T059|1011335|CPT|CL-|CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE MEASUREMENT |CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE MEASUREMENT, NOS|CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE EACH TEST|CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE EA.TST|CHLORIDE
C0201975|T059|82565|CPT|CREATININE MEASUREMENT|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE; BLOOD|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|BLOOD CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|TEST;CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE BLOOD|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|BLOOD CREATININE LEVEL|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|MEASUREMENT OF CREATININE|BLOOD CREATININE LEVEL
# C0201975|T059|82565|CPT|CR|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|LAB-BASED CHEM MEASUREMENTS CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|MEASUREMENT OF CREATININE |BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREAT|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|BLOOD CREATININE LEVEL |BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE MEASUREMENT |BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE MEASUREMENT, NOS|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|ASSAY OF CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE TEST|BLOOD CREATININE LEVEL
C0201930|T059|82374|CPT|CARBON DIOXIDE CONTENT MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CO2 CONTENT MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|PCO2, BLOOD|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CO<SUB>2</SUB> CONTENT MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|PCO<SUB>2</SUB>, BLOOD|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE (BICARBONATE)|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|ASSAY BLOOD CARBON DIOXIDE|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE BICARBONATE|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|MEASUREMENT OF CARBON DIOXIDE|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CO2|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|PCO>2<, BLOOD|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CO>2< CONTENT MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE CONTENT MEASUREMENT |ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE MEASUREMENT |ASSAY BLOOD CARBON DIOXIDE
C0005845|T059|84520|CPT|BLOOD UREA NITROGEN|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BUN|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|NITROGEN, BLOOD UREA|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|UREA NITROGEN, BLOOD|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA NITROGEN MEASUREMENT|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|UREA NITROGEN; QUANTITATIVE|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BUN LEVEL|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|MEASUREMENT OF BLOOD UREA NITROGEN (BUN)|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|ASSAY OF UREA NITROGEN QUANTITATIVE|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|MEASUREMENT OF UREA NITROGEN (BUN)|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|UREA - BLOOD|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA |ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA NITROGEN MEASUREMENT |ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BUN MEASUREMENT|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA MEASUREMENT |ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA MEASUREMENT|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA NITROGEN MEASUREMENT |ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|ASSAY OF UREA NITROGEN|ASSAY OF UREA NITROGEN QUANTITATIVE
C0200379|T059|80050|CPT|GENERAL HEALTH PANEL|GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)
C0200379|T059|80050|CPT|GENERAL HEALTH PANEL |GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)
C0200379|T059|80050|CPT|GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)|GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)
C0200379|T059|80050|CPT|GENERAL HEALTH PANEL, NOS|GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)
C0201836|T059|84460|CPT|ALANINE AMINOTRANSFERASE MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALANINE AMINOTRANSFERASE|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
# C0201836|T059|84460|CPT|ALT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|TRANSFERASE; ALANINE AMINO (ALT) (SGPT)|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|TEST;ALANINE AMINOTRANSFERASE|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|TRANSFERASE ALANINE AMINO ALT SGPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|LIVER ENZYME (SGPT), LEVEL|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALANINE AMINO (ALT) (SGPT)|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|SGPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|GLUTAMIC-PYRUVATE TRANSAMINASE|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|GPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|GPT MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|GLUTAMIC PYRUVATE TRANSAMINASE MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|SGPT MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALT MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALANINE AMINOTRANSFERASE MEASUREMENT |MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALANINE AMINOTRANSFERASE TEST|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201913|T059|1011294|CPT|BILIRUBIN; TOTAL|BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN MEASUREMENT|BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN TOTAL|BILIRUBIN
C0201913|T059|1011294|CPT|MEASUREMENT OF TOTAL BILIRUBIN|BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN|BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN (& LEVEL) |BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN, TOTAL MEASUREMENT|BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN, TOTAL MEASUREMENT |BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN (& LEVEL)|BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN|BILIRUBIN
C0201913|T059|1011294|CPT|BILI|BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN LEVEL|BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN, TOTAL MEASUREMENT  [AMBIGUOUS]|BILIRUBIN
C0523465|T059|82040|CPT|SERUM ALBUMIN|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN MEASUREMENT|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN SERUM PLASMA/WHOLE BLOOD|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN; SERUM, PLASMA OR WHOLE BLOOD|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN MEASUREMENT |ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|MEASUREMENT OF ALBUMIN IN SERUM|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN (& LEVEL) |ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN - SERUM|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN (& LEVEL)|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN TEST|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN MEASUREMENT, SERUM|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN LEVEL|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SA - SERUM ALBUMIN|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN MEASUREMENT, SERUM |ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ASSAY OF SERUM ALBUMIN|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523658|T059|82947|CPT|ASSAY GLUCOSE BLOOD QUANT|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T059|82947|CPT|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T059|82947|CPT|GLUCOSE QUANTITATIVE BLOOD XCPT REAGENT STRIP|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T059|82947|CPT|GLUCOSE MEASUREMENT, QUANTITATIVE|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T059|82947|CPT|GLUCOSE MEASUREMENT, QUANTITATIVE |GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0201899|T059|80076|CPT|SERUM SGOT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SERUM AST|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPARTATE AMINOTRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
# C0201899|T059|80076|CPT|GOT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
# C0201899|T059|80076|CPT|AST|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPARTATE AMINOTRANSFERASE MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|TRANSFERASE; ASPARTATE AMINO (AST) (SGOT)|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|TRANSFERASE ASPARTATE AMINO AST SGOT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|LIVER ENZYME (SGOT), LEVEL|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE (AST) (SGOT)|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|AST - ASPARTATE TRANSAM SGOT (& LEVEL) |MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|AST - ASPARTATE TRANSAM SGOT (& LEVEL)|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|TRANSFERASE (AST) (SGOT)|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SGOT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPARTATE TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASP TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SERUM GLUTAMIC-OXALOACETIC TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|GLUTAMIC-OXALOACETIC TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SERUM ASPARTATE TRANSAMINASE TEST|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|AST MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|GLUTAMIC OXALOACETIC TRANSAMINASE MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|GOT MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SGOT MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPARTATE AMINOTRANSFERASE MEASUREMENT |MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0391938|T059|82435|CPT|CHLORIDE; BLOOD|CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE|CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE LEVEL|CHLORIDE BLD
C0391938|T059|82435|CPT|MEASUREMENT OF CHLORIDE IN BLOOD|CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE LEVEL |CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE LEVEL |CHLORIDE BLD
C0391938|T059|82435|CPT|CHLORIDE MEASUREMENT, BLOOD|CHLORIDE BLD
C0391938|T059|82435|CPT|CHLORIDE MEASUREMENT, BLOOD |CHLORIDE BLD
C0391938|T059|82435|CPT|ASSAY OF BLOOD CHLORIDE|CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE LEVEL MEASUREMENT|CHLORIDE BLD
C0391938|T059|82435|CPT|CHLORIDE BLD|CHLORIDE BLD
C0523891|T059|84295|CPT|SERUM SODIUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM NA+|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM MEASUREMENT|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM MEASUREMENT |SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM; SERUM, PLASMA OR WHOLE BLOOD|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM SERUM PLASMA OR WHOLE BLOOD|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|MEASUREMENT OF SODIUM IN SERUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM (& LEVEL) |SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM (& LEVEL)|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM - SERUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM ION TEST|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM MEASUREMENT, SERUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM LEVEL|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM MEASUREMENT, SERUM |SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|ASSAY OF SERUM SODIUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM EACH TEST|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM EA.TST|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM K+|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM MEASUREMENT|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM MEASUREMENT |POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|POTASSIUM LEVEL|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|POTASSIUM SERUM PLASMA/WHOLE BLOOD|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|POTASSIUM; SERUM, PLASMA OR WHOLE BLOOD|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|MEASUREMENT OF POTASSIUM IN SERUM|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|POTASSIUM - SERUM|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM (& LEVEL) |POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM (& LEVEL)|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM LEVEL|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM MEASUREMENT |POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|ASSAY OF SERUM POTASSIUM|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0373708|T059|84155|CPT|PROTEIN, TOTAL, EXCEPT BY REFRACTOMETRY; SERUM, PLASMA OR WHOLE BLOOD|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD
C0373708|T059|84155|CPT|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD
C0373708|T059|84155|CPT|ASSAY OF PROTEIN SERUM|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD
C4048459|T059|80055|CPT|OBSTETRIC PANEL|OBSTETRIC PANEL
C4048459|T059|80055|CPT|OBSTETRIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) HEPATITIS B SURFACE ANTIGEN (HBSAG) (87340) ANTIBODY, RUBELLA (86762) SYPHILIS TEST, NON-TREPONEMAL ANTIBODY; QUALITATIVE (EG, VDRL, RPR, ART) (86592) ANTIBODY SCREEN, RBC, EACH SERUM TECHNIQUE (86850) BLOOD TYPING, ABO (86900) AND BLOOD TYPING, RH (D) (86901)|OBSTETRIC PANEL
C0812553|T059|80074|CPT|ACUTE HEPATITIS PANEL|ACUTE HEPATITIS PANEL
C0812553|T059|80074|CPT|ACUTE HEPATITIS PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: HEPATITIS A ANTIBODY (HAAB), IGM ANTIBODY (86709) HEPATITIS B CORE ANTIBODY (HBCAB), IGM ANTIBODY (86705) HEPATITIS B SURFACE ANTIGEN (HBSAG) (87340) HEPATITIS C ANTIBODY (86803)|ACUTE HEPATITIS PANEL
C0519824|T059|80051|CPT|ELECTROLYTE PANEL|ELECTROLYTE PANEL
C0519824|T059|80051|CPT|ELECTROLYTES PANEL|ELECTROLYTE PANEL
C0519824|T059|80051|CPT|ELECTROLYTE PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) POTASSIUM (84132) SODIUM (84295)|ELECTROLYTE PANEL
C0519824|T059|80051|CPT|BLOOD ELECTROLYTE PANEL|ELECTROLYTE PANEL
C0519824|T059|80051|CPT|BLOOD ELECTROLYTE PANEL |ELECTROLYTE PANEL
C1964052|T059|80047|CPT|BASIC METABOLIC PANEL CALCIUM IONIZED|METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|METABOLIC PANEL IONIZED CA|METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|BMP WITH IONIZED CALCIUM|METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|BASIC METABOLIC PANEL WITH IONIZED CALCIUM |METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|BASIC METABOLIC PANEL WITH IONIZED CALCIUM|METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|BASIC METABOLIC PANEL (CALCIUM, IONIZED) THIS PANEL MUST INCLUDE THE FOLLOWING: CALCIUM, IONIZED (82330) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) POTASSIUM (84132) SODIUM (84295) UREA NITROGEN (BUN) (84520)|METABOLIC PANEL IONIZED CA
C0200382|T059|80061|CPT|LIPID PANEL|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|LIPIDS TEST PANEL|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|LIPID PANEL |LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|BLOOD TEST, LIPIDS (CHOLESTEROL AND TRIGLYCERIDES)|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|LIPID PANEL |LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0519823|T059|80048|CPT|METABOLIC PANEL TOTAL CA|BASIC METABOLIC PANEL CALCIUM TOTAL
C0519823|T059|80048|CPT|BASIC METABOLIC PANEL CALCIUM TOTAL|BASIC METABOLIC PANEL CALCIUM TOTAL
C0519823|T059|80048|CPT|BASIC METABOLIC PANEL (CALCIUM, TOTAL) THIS PANEL MUST INCLUDE THE FOLLOWING: CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) POTASSIUM (84132) SODIUM (84295) UREA NITROGEN (BUN) (84520)|BASIC METABOLIC PANEL CALCIUM TOTAL
C0374833|T059|1011137|CPT|ORGAN OR DISEASE ORIENTED PANELS|ORGAN OR DISEASE ORIENTED PANELS
C0812554|T059|80076|CPT|HEPATIC FUNCTION PANEL|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)
C0812554|T059|80076|CPT|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)
C0812554|T059|80076|CPT|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT)|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)
C0812554|T059|80076|CPT|LIVER FUNCTION BLOOD TEST PANEL|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)
C0812552|T059|80069|CPT|RENAL FUNCTION PANEL |RENAL FUNCTION PANEL
C0812552|T059|80069|CPT|RENAL FUNCTION PANEL|RENAL FUNCTION PANEL
C0812552|T059|80069|CPT|RENAL FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHORUS INORGANIC (PHOSPHATE) (84100) POTASSIUM (84132) SODIUM (84295) UREA NITROGEN (BUN) (84520)|RENAL FUNCTION PANEL
C0812552|T059|80069|CPT|KIDNEY FUNCTION BLOOD TEST PANEL|RENAL FUNCTION PANEL
C0430174|T059||CPT|METABOLIC FUNCTION TESTED
C0430174|T059||CPT|METABOLIC FUNCTION TEST NOS 
C0430174|T059||CPT|METABOLIC FUNCTION TEST NOS
C0430174|T059||CPT|METABOLIC FUNCTION TESTED 
C0430174|T059||CPT|METABOLIC FUNCTION TEST
C0430174|T059||CPT|METABOLIC FUNCTION TEST 
C0430174|T059||CPT|METABOLIC FUNCTION TESTED 
C4050228|T059|80081|CPT|OBSTETRIC PANEL|OBSTETRIC PANEL
C4050228|T059|80081|CPT|OBSTETRIC PANEL (INCLUDES HIV TESTING) THIS PANEL MUST INCLUDE THE FOLLOWING: BLOOD COUNT, COMPLETE (CBC), AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) HEPATITIS B SURFACE ANTIGEN (HBSAG) (87340) HIV-1 ANTIGEN(S), WITH HIV-1 AND HIV-2 ANTIBODIES, SINGLE RESULT (87389) ANTIBODY, RUBELLA (86762) SYPHILIS TEST, NON-TREPONEMAL ANTIBODY; QUALITATIVE (EG, VDRL, RPR, ART) (86592) ANTIBODY SCREEN, RBC, EACH SERUM TECHNIQUE (86850) BLOOD TYPING, ABO (86900) AND BLOOD TYPING, RH (D) (86901)|OBSTETRIC PANEL
C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC PANEL|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC CHEMICAL PANEL|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|BLOOD TEST, COMPREHENSIVE GROUP OF BLOOD CHEMICALS|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC PANEL |COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHENSIVE METABOLIC CHEM PANEL|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519825|T059|80053|CPT|COMPREHEN METABOLIC PANEL|COMPREHENSIVE METABOLIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHATASE, ALKALINE (84075) POTASSIUM (84132) PROTEIN, TOTAL (84155) SODIUM (84295) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450) UREA NITROGEN (BUN) (84520)
C0519824|T059|80051|CPT|ELECTROLYTE PANEL|ELECTROLYTE PANEL
C0519824|T059|80051|CPT|ELECTROLYTES PANEL|ELECTROLYTE PANEL
C0519824|T059|80051|CPT|ELECTROLYTE PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) POTASSIUM (84132) SODIUM (84295)|ELECTROLYTE PANEL
C0519824|T059|80051|CPT|BLOOD ELECTROLYTE PANEL|ELECTROLYTE PANEL
C0519824|T059|80051|CPT|BLOOD ELECTROLYTE PANEL |ELECTROLYTE PANEL
C0812552|T059|80069|CPT|RENAL FUNCTION PANEL |RENAL FUNCTION PANEL
C0812552|T059|80069|CPT|RENAL FUNCTION PANEL|RENAL FUNCTION PANEL
C0812552|T059|80069|CPT|RENAL FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) PHOSPHORUS INORGANIC (PHOSPHATE) (84100) POTASSIUM (84132) SODIUM (84295) UREA NITROGEN (BUN) (84520)|RENAL FUNCTION PANEL
C0812552|T059|80069|CPT|KIDNEY FUNCTION BLOOD TEST PANEL|RENAL FUNCTION PANEL
C2010717|T059||CPT|GENERAL HEALTH TEST PANEL 
C2010717|T059||CPT|GENERAL HEALTH TEST PANEL
C0023901|T059||CPT|FUNCTION TEST, LIVER
C0023901|T059||CPT|FUNCTION TESTS, LIVER
C0023901|T059||CPT|LIVER FUNCTION TEST
C0023901|T059||CPT|LIVER FUNCTION TESTS
C0023901|T059||CPT|TEST, LIVER FUNCTION
C0023901|T059||CPT|TESTS, LIVER FUNCTION
C0023901|T059||CPT|HEPATIC FUNCTION PANEL
C0023901|T059||CPT|HEPATIC FUNCTION PANEL 
C0023901|T059||CPT|LIVER FUNCTION ANALYSES
C0023901|T059||CPT|LFTS
C0023901|T059||CPT|LFT
C0023901|T059||CPT|LIVER STUDY
C0023901|T059||CPT|TEST;LIVER FUNCTION
C0023901|T059||CPT|LIVER FUNCTION TESTS NOS
C0023901|T059||CPT|LIVER FUNCTION TESTS (& [GENERAL])
C0023901|T059||CPT|LIVER FUNCT. TEST -GEN.
C0023901|T059||CPT|LIVER FUNCTION TESTS (& GENERAL)
C0023901|T059||CPT|LIVER FUNCTION TESTS (& [GENERAL]) 
C0023901|T059||CPT|LIVER FUNCTION TESTS 
C0023901|T059||CPT|LIVER FUNCTION TESTS (& GENERAL) 
C0023901|T059||CPT|LIVER FUNCTION TESTS NOS 
C0023901|T059||CPT|LIVER FUNCTION TESTS - GENERAL
C0023901|T059||CPT|LFT - LIVER FUNCTION TEST
C0023901|T059||CPT|HEPATIC FUNCTION PANEL 
C0023901|T059||CPT|LIVER FUNCTION TESTS - GENERAL 
C0023901|T059||CPT|LFT'S
C2030682|T059||CPT|HEPATITIS SCREEN PANEL 
C2030682|T059||CPT|HEPATITIS SCREEN PANEL
C0200382|T059|80061|CPT|LIPID PANEL|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|LIPIDS TEST PANEL|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|LIPID PANEL |LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|BLOOD TEST, LIPIDS (CHOLESTEROL AND TRIGLYCERIDES)|LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C0200382|T059|80061|CPT|LIPID PANEL |LIPID PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: CHOLESTEROL, SERUM, TOTAL (82465) LIPOPROTEIN, DIRECT MEASUREMENT, HIGH DENSITY CHOLESTEROL (HDL CHOLESTEROL) (83718) TRIGLYCERIDES (84478)
C2041460|T059||CPT|ARTHRITIS TEST PANEL
C2041460|T059||CPT|ARTHRITIS TEST PANEL 
C2041461|T059||CPT|TORCH ANTIBODY PANEL 
C2041461|T059||CPT|TORCH ANTIBODY PANEL
C0027617|T059||CPT|NEONATAL SCREENING
C0027617|T059||CPT|NEONATAL SCREENINGS
C0027617|T059||CPT|NEWBORN INFANT SCREENINGS
C0027617|T059||CPT|SCREENING, NEONATAL
C0027617|T059||CPT|SCREENING, NEWBORN INFANT
C0027617|T059||CPT|SCREENINGS, NEONATAL
C0027617|T059||CPT|SCREENINGS, NEWBORN INFANT
C0027617|T059||CPT|NEWBORN SCREEN 
C0027617|T059||CPT|NEWBORN SCREEN
C0027617|T059||CPT|NEWBORN ASSESSMENT
C0027617|T059||CPT|NEWBORN SCREENING
C0027617|T059||CPT|SCREENING, NEWBORN
C0027617|T059||CPT|INFANT, NEWBORN, SCREENING
C0027617|T059||CPT|NEWBORN INFANT SCREENING
C0027617|T059||CPT|NEONATAL SCREENING 
C0027617|T059||CPT|NEONATAL SCREENING, NOS
C0027617|T059||CPT|NEONATAL SCREENING TEST
C2210821|T059||CPT|BASIC THYROID PANEL
C2210821|T059||CPT|BASIC THYROID PANEL 
C2106943|T059||CPT|COMPREHENSIVE THYROID PANEL 
C2106943|T059||CPT|COMPREHENSIVE THYROID PANEL
C2237045|T059|80047|CPT|CHEM 7|BLOOD TEST, BASIC GROUP OF BLOOD CHEMICALS
C2237045|T059|80047|CPT|SMAC 7|BLOOD TEST, BASIC GROUP OF BLOOD CHEMICALS
C2237045|T059|80047|CPT|BASIC METABOLIC PANEL|BLOOD TEST, BASIC GROUP OF BLOOD CHEMICALS
C2237045|T059|80047|CPT|BASIC METABOLIC PANEL |BLOOD TEST, BASIC GROUP OF BLOOD CHEMICALS
C2237045|T059|80047|CPT|BMP (BASIC METABOLIC PANEL)|BLOOD TEST, BASIC GROUP OF BLOOD CHEMICALS
C2237045|T059|80047|CPT|BLOOD TEST, BASIC GROUP OF BLOOD CHEMICALS|BLOOD TEST, BASIC GROUP OF BLOOD CHEMICALS
C1315055|T059||CPT|CARDIAC STUDIES ORDER SET
C1315055|T059||CPT|CARDIAC PANEL 
C1315055|T059||CPT|CARDIAC PANEL
C1315055|T059||CPT|PANEL.CARDIAC
C3836618|T059||CPT|OBSTETRIC 1996 PANEL IN SERUM AND BLOOD 
C3836618|T059||CPT|OBSTETRIC 1996 PANEL IN SERUM AND BLOOD
C4064645|T059||CPT|MATERNAL SERUM OR PLASMA SCREENING
C4064645|T059||CPT|MATERNAL SERUM OR PLASMA SCREENING 
C2122148|T059||CPT|BASIC METABOLIC CHEM PANEL
C2122148|T059||CPT|BASIC METABOLIC CHEMISTRY PANEL
C2122148|T059||CPT|BASIC METABOLIC CHEM PANEL 
C0438930|T059||CPT|CHEM. METABOLIC FUNCTION TESTS
C0438930|T059||CPT|CHEM. METABOLIC FUNCTION TESTS 
C0523464|T059||CPT|ALBUMIN RENAL CLEARANCE MEASUREMENT
C0523464|T059||CPT|ALBUMIN RENAL CLEARANCE MEASUREMENT 
C0201837|T059||CPT|ALBUMIN/GLOBULIN RATIO
C0201837|T059||CPT|ALBUMIN GLOBULIN RATIO
C0201837|T059||CPT|A/G RATIO
C0201837|T059||CPT|ALBUMIN/GLOBULIN RATIO 
C0523465|T059|82040|CPT|SERUM ALBUMIN|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN MEASUREMENT|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN SERUM PLASMA/WHOLE BLOOD|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN; SERUM, PLASMA OR WHOLE BLOOD|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN MEASUREMENT |ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|MEASUREMENT OF ALBUMIN IN SERUM|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN (& LEVEL) |ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN - SERUM|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN (& LEVEL)|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN TEST|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN MEASUREMENT, SERUM|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SERUM ALBUMIN LEVEL|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|SA - SERUM ALBUMIN|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ALBUMIN MEASUREMENT, SERUM |ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|T059|82040|CPT|ASSAY OF SERUM ALBUMIN|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0201838|T059|1011249|CPT|ALBUMIN MEASUREMENT|ALBUMIN
C0201838|T059|1011249|CPT|TEST;ALBUMIN|ALBUMIN
C0201838|T059|1011249|CPT|MEASUREMENT OF ALBUMIN|ALBUMIN
C0201838|T059|1011249|CPT|ALBUMIN|ALBUMIN
C0201838|T059|1011249|CPT|ALB|ALBUMIN
C0201838|T059|1011249|CPT|MICROALBUMIN|ALBUMIN
C0201838|T059|1011249|CPT|ALBUMIN MEASUREMENT |ALBUMIN
C0201838|T059|1011249|CPT|ALBUMIN TEST|ALBUMIN
C1278236|T059||CPT|24 HOUR URINE ALBUMIN OUTPUT
C1278236|T059||CPT|24 HOUR URINE ALBUMIN OUTPUT 
C1278236|T059||CPT|24 HOUR URINE ALBUMIN OUTPUT MEASUREMENT 
C1278236|T059||CPT|24 HOUR URINE ALBUMIN OUTPUT MEASUREMENT
C0523466|T059|82042|CPT|ALBUMIN; URINE OR OTHER SOURCE, QUANTITATIVE, EACH SPECIMEN|OTHER SOURCE ALBUMIN QUAN EA
C0523466|T059|82042|CPT|ALBUMIN URINE/OTHER SOURCE QUAN EACH SPECIMEN|OTHER SOURCE ALBUMIN QUAN EA
C0523466|T059|82042|CPT|ALBUMIN MEASUREMENT, URINE, QUANTITATIVE|OTHER SOURCE ALBUMIN QUAN EA
C0523466|T059|82042|CPT|ALBUMIN MEASUREMENT, URINE, QUANTITATIVE |OTHER SOURCE ALBUMIN QUAN EA
C0523466|T059|82042|CPT|ASSAY OF URINE ALBUMIN|OTHER SOURCE ALBUMIN QUAN EA
C0373533|T059|82044|CPT|ALBUMIN; URINE, MICROALBUMIN, SEMIQUANTITATIVE (EG, REAGENT STRIP ASSAY)|UR ALBUMIN SEMIQUANTITATIVE
C0373533|T059|82044|CPT|MICROALBUMIN SEMIQUANT|UR ALBUMIN SEMIQUANTITATIVE
C0373533|T059|82044|CPT|ALBUMIN URINE MICROALBUMIN SEMIQUANTITATIVE|UR ALBUMIN SEMIQUANTITATIVE
C0373533|T059|82044|CPT|SEMIQUANTITATIVE ANALYSIS OF MICROALBUMIN IN URINE|UR ALBUMIN SEMIQUANTITATIVE
C1504155|T059|82045|CPT|SERUM ALBUMIN ISCHEMIA MODIFIED |ALBUMIN; ISCHEMIA MODIFIED
C1504155|T059|82045|CPT|SERUM ALBUMIN ISCHEMIA MODIFIED|ALBUMIN; ISCHEMIA MODIFIED
C1504155|T059|82045|CPT|ISCHEMIA-MODIFIED SERUM ALBUMIN|ALBUMIN; ISCHEMIA MODIFIED
C1504155|T059|82045|CPT|ALBUMIN ISCHEMIA MODIFIED|ALBUMIN; ISCHEMIA MODIFIED
C1504155|T059|82045|CPT|SERUM ALBUMIN ISCHEMIA MODIFIED LAB PROCEDURE|ALBUMIN; ISCHEMIA MODIFIED
C1504155|T059|82045|CPT|ALBUMIN; ISCHEMIA MODIFIED|ALBUMIN; ISCHEMIA MODIFIED
C0373532|T059|82043|CPT|ALBUMIN; URINE, MICROALBUMIN, QUANTITATIVE|UR ALBUMIN QUANTITATIVE
C0373532|T059|82043|CPT|MICROALBUMIN QUANTITATIVE|UR ALBUMIN QUANTITATIVE
C0373532|T059|82043|CPT|ALBUMIN URINE MICROALBUMIN QUANTIATIVE|UR ALBUMIN QUANTITATIVE
C0523674|T059||CPT|ALBGLYCA
C0523674|T059||CPT|GLYCATED ALBUMIN
C0523674|T059||CPT|GLYCATED ALBUMIN MEASUREMENT
C0523674|T059||CPT|GLYCATED ALBUMIN MEASUREMENT 
C1278275|T059||CPT|CEREBROSPINAL FLUID ALBUMIN LEVEL
C1278275|T059||CPT|CEREBROSPINAL FLUID ALBUMIN LEVEL 
C1278275|T059||CPT|CEREBROSPINAL FLUID ALBUMIN MEASUREMENT 
C1278275|T059||CPT|CEREBROSPINAL FLUID ALBUMIN MEASUREMENT
C0428520|T059||CPT|FLUID SAMPLE ALBUMIN LEVEL
C0428520|T059||CPT|FLUID SAMPLE ALBUMIN MEASUREMENT 
C0428520|T059||CPT|FLUID SAMPLE ALBUMIN MEASUREMENT
C0428623|T059||CPT|ALBUMIN/IMMUNOGLOBULIN G RATIO
C0428623|T059||CPT|IGG - ALBUMIN/IMMUNOGLOBULIN G RATIO
C0428623|T059||CPT|ALBUMIN/IMMUNOGLOBULIN G RATIO MEASUREMENT 
C0428623|T059||CPT|ALBUMIN/IMMUNOGLOBULIN G RATIO MEASUREMENT
C1272106|T059||CPT|PLASMA ALBUMIN LEVEL 
C1272106|T059||CPT|PLASMA ALBUMIN LEVEL
C1273508|T059||CPT|SERUM PREALBUMIN LEVEL
C1273508|T059||CPT|SERUM PREALBUMIN LEVEL 
C1318429|T059||CPT|MEASUREMENT OF ALBUMIN IN URINE
C1318429|T059||CPT|URINE ALBUMIN (& LEVEL) 
C1318429|T059||CPT|URINE ALBUMIN (& LEVEL)
C1318429|T059||CPT|URINE ALBUMIN LEVEL
C1318429|T059||CPT|URINE ALBUMIN MEASUREMENT 
C1318429|T059||CPT|URINE ALBUMIN MEASUREMENT
C0523463|T059||CPT|CSF ALBUMIN/PLASMA ALBUMIN RATIO MEASUREMENT 
C0523463|T059||CPT|CEREBROSPINAL FLUID ALBUMIN/PLASMA ALBUMIN RATIO MEASUREMENT 
C0523463|T059||CPT|CEREBROSPINAL FLUID ALBUMIN/PLASMA ALBUMIN RATIO MEASUREMENT
C0523463|T059||CPT|CSF ALBUMIN/PLASMA ALBUMIN RATIO MEASUREMENT
C0025634|T059|83857|CPT|METHEMALBUMIN|METHEMALBUMIN (PROTEIN) LEVEL
C0025634|T059|83857|CPT|METHEMALBUMIN ASSAY|METHEMALBUMIN (PROTEIN) LEVEL
C0025634|T059|83857|CPT|METHEMALBUMIN (PROTEIN) LEVEL|METHEMALBUMIN (PROTEIN) LEVEL
C0025634|T059|83857|CPT|MEASUREMENT OF METHEMALBUMIN|METHEMALBUMIN (PROTEIN) LEVEL
C0025634|T059|83857|CPT|METHEMALBUMIN MEASUREMENT|METHEMALBUMIN (PROTEIN) LEVEL
C0025634|T059|83857|CPT|METHAEMALBUMIN MEASUREMENT|METHEMALBUMIN (PROTEIN) LEVEL
C0025634|T059|83857|CPT|METHEMALBUMIN MEASUREMENT |METHEMALBUMIN (PROTEIN) LEVEL
C0025634|T059|83857|CPT|ASSAY OF METHEMALBUMIN|METHEMALBUMIN (PROTEIN) LEVEL
C1293929|T059||CPT|MEASUREMENT OF RATIO OF ANALYTE TO ALBUMIN 
C1293929|T059||CPT|MEASUREMENT OF RATIO OF ANALYTE TO ALBUMIN
C0201925|T059|82310|CPT|CALCIUM; TOTAL|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM MEASUREMENT|ASSAY OF CALCIUM
# C0201925|T059|82310|CPT|CA|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM TOTAL|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|MEASUREMENT OF CALCIUM|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM LEVEL|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|LAB-BASED CHEM MEASUREMENTS CALCIUM|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|MEASUREMENT OF CALCIUM |ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CA++|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM MEASUREMENT |ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM MEASUREMENT, NOS|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|ASSAY OF CALCIUM|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CALCIUM TOTAL EACH TEST|ASSAY OF CALCIUM
C0201925|T059|82310|CPT|CA TOT EA.TST|ASSAY OF CALCIUM
C0728876|T059||CPT|SERUM CALCIUM
C0728876|T059||CPT|SERUM CA++
C0728876|T059||CPT|SERUM CALCIUM MEASUREMENT
C0728876|T059||CPT|SERUM CALCIUM (& LEVEL) 
C0728876|T059||CPT|SERUM CALCIUM (& LEVEL)
C0728876|T059||CPT|CALCIUM - SERUM
C0728876|T059||CPT|SERUM CALCIUM TEST
C0728876|T059||CPT|SERUM CALCIUM LEVEL
C0728876|T059||CPT|SERUM CALCIUM MEASUREMENT 
C0428303|T059|82340|CPT|URINE CALCIUM|URINE CALCIUM LEVEL
C0428303|T059|82340|CPT|URINE CALCIUM MEASUREMENT|URINE CALCIUM LEVEL
C0428303|T059|82340|CPT|URINE CALCIUM MEASUREMENT |URINE CALCIUM LEVEL
C0428303|T059|82340|CPT|URINE CALCIUM LEVEL|URINE CALCIUM LEVEL
C0428303|T059|82340|CPT|CALCIUM - URINE|URINE CALCIUM LEVEL
C0428303|T059|82340|CPT|URINE CALCIUM (& LEVEL) |URINE CALCIUM LEVEL
C0428303|T059|82340|CPT|URINE CALCIUM (& LEVEL)|URINE CALCIUM LEVEL
C0428303|T059|82340|CPT|URINE CALCIUM TEST|URINE CALCIUM LEVEL
C0428303|T059|82340|CPT|CALCIUM MEASUREMENT, URINE|URINE CALCIUM LEVEL
C0428303|T059|82340|CPT|CALCIUM MEASUREMENT, URINE |URINE CALCIUM LEVEL
C0430040|T059||CPT|CALCIUM PROFILE
C0430040|T059||CPT|CALCIUM PROFILE 
C1278284|T059||CPT|CALCULUS CALCIUM CONTENT
C1278284|T059||CPT|CALCULUS CALCIUM CONTENT 
C1278284|T059||CPT|CALCULUS CALCIUM CONTENT MEASUREMENT 
C1278284|T059||CPT|CALCULUS CALCIUM CONTENT MEASUREMENT
C1271835|T059||CPT|FLUID SAMPLE CALCIUM LEVEL 
C1271835|T059||CPT|FLUID SAMPLE CALCIUM LEVEL
C2711247|T059||CPT|CALCULATION OF IONIZED CALCIUM CONCENTRATION
C2711247|T059||CPT|CALCULATION OF IONISED CALCIUM CONCENTRATION
C2711247|T059||CPT|CALCULATION OF IONIZED CALCIUM CONCENTRATION 
C2732404|T059||CPT|CORRECTED MEASUREMENT OF CALCIUM
C2732404|T059||CPT|CORRECTED MEASUREMENT OF CALCIUM 
C2732404|T059||CPT|CALCIUM CORRECTED
C2732404|T059||CPT|CACR
C2732404|T059||CPT|CALCIUM CORRECTED MEASUREMENT
C3272884|T059||CPT|CALCIUM CLEARANCE MEASUREMENT
C3272884|T059||CPT|CALCIUM CLEARANCE
C3272884|T059||CPT|CACLR
C0201927|T059|80047|CPT|MEASUREMENT OF SERUM IONIZED CALCIUM|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|MEASUREMENT OF SERUM IONISED CALCIUM|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|SERUM IONIZED CALCIUM MEASUREMENT|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|SERUM IONISED CALCIUM MEASUREMENT |MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|MEASUREMENT OF SERUM IONIZED CALCIUM |MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|SERUM IONIZED CALCIUM MEASUREMENT |MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|IONIZED CALCIUM LEVEL|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|IONIZED CALCIUM MEASUREMENT|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|MEASUREMENT OF IONIZED CALCIUM|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|SERUM IONISED CALCIUM LEVEL |MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|SERUM IONISED CALCIUM LEVEL|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|CALCIUM, SERUM, IONIZED MEASUREMENT|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|CALCIUM, SERUM, IONIZED MEASUREMENT |MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|CALCIUM, SERUM, IONISED MEASUREMENT|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|CAION|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|CALCIUM, IONIZED|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|SERUM IONIZED CALCIUM LEVEL|MEASUREMENT OF IONIZED CALCIUM
C0201927|T059|80047|CPT|SERUM IONISED CALCIUM MEASUREMENT|MEASUREMENT OF IONIZED CALCIUM
C0373563|T059|82340|CPT|CALCIUM; URINE QUANTITATIVE, TIMED SPECIMEN|ASSAY OF CALCIUM IN URINE
C0373563|T059|82340|CPT|CALCIUM URINE QUANTITATIVE TIMED SPECIMEN|ASSAY OF CALCIUM IN URINE
C0373563|T059|82340|CPT|ASSAY OF CALCIUM IN URINE|ASSAY OF CALCIUM IN URINE
C0523539|T059|82331|CPT|CALCIUM; AFTER CALCIUM INFUSION TEST|MEASUREMENT OF CALCIUM AFTER CALCIUM INFUSION TEST
C0523539|T059|82331|CPT|CALCIUM CHALLENGE TESTS |MEASUREMENT OF CALCIUM AFTER CALCIUM INFUSION TEST
C0523539|T059|82331|CPT|CALCIUM AFTER CALCIUM INFUSION TEST|MEASUREMENT OF CALCIUM AFTER CALCIUM INFUSION TEST
C0523539|T059|82331|CPT|MEASUREMENT OF CALCIUM AFTER CALCIUM INFUSION TEST|MEASUREMENT OF CALCIUM AFTER CALCIUM INFUSION TEST
C0523539|T059|82331|CPT|CALCIUM CHALLENGE TESTS|MEASUREMENT OF CALCIUM AFTER CALCIUM INFUSION TEST
C0523539|T059|82331|CPT|CALCIUM MEASUREMENT AFTER CALCIUM INFUSION|MEASUREMENT OF CALCIUM AFTER CALCIUM INFUSION TEST
C0523539|T059|82331|CPT|CALCIUM INFUSION TEST|MEASUREMENT OF CALCIUM AFTER CALCIUM INFUSION TEST
C0489943|T059|82330|CPT|CALCIUM; IONIZED|ASSAY OF CALCIUM
C0489943|T059|82330|CPT|IONIZED CALCIUM ASSAY|ASSAY OF CALCIUM
C0489943|T059|82330|CPT|CALCIUM IONIZED|ASSAY OF CALCIUM
C0489943|T059|82330|CPT|IONIZED CALCIUM|ASSAY OF CALCIUM
C0489943|T059|82330|CPT|CALCIUM IONISED|ASSAY OF CALCIUM
C0489943|T059|82330|CPT|ASSAY OF CALCIUM|ASSAY OF CALCIUM
C0489943|T059|82330|CPT|CALCIUM IONIZED EACH TEST|ASSAY OF CALCIUM
C0489943|T059|82330|CPT|CA IONIZED EA.TST|ASSAY OF CALCIUM
C3830083|T059||CPT|FECA
C3830083|T059||CPT|FRACTIONAL EXCRETION OF CALCIUM
C3830083|T059||CPT|FRACTIONAL EXCRETION OF CA
C3830083|T059||CPT|FRACTIONAL CALCIUM EXCRETION
C0201928|T059||CPT|CALCIUM EXCRETION, 2-HOUR COLLECTION, FASTING, URINE
C0201928|T059||CPT|CALCIUM EXCRETION, 2-HOUR COLLECTION, FASTING, URINE 
C0278369|T059||CPT|CALCIUM MEASUREMENT IN 24 HOUR EXCRETION IN FECES
C0278369|T059||CPT|CALCIUM MEASUREMENT IN 24 HOUR EXCRETION IN FAECES
C0278369|T059||CPT|CALCIUM MEASUREMENT IN 24 HOUR EXCRETION IN FECES 
C0278369|T059||CPT|CALCIUM MEASUREMENT, 24H STOOL
C0278369|T059||CPT|CALCIUM TOTAL MEASUREMENT, 24 HOUR EXCRETION IN STOOL
C0729820|T059||CPT|BLOOD CALCIUM
C0729820|T059||CPT|BLOOD CALCIUM LEVEL
C0729820|T059||CPT|BLOOD CALCIUM LEVEL 
C0729820|T059||CPT|BLOOD CALCIUM MEASUREMENT 
C0729820|T059||CPT|CALCIUM BLOOD
C0729820|T059||CPT|BLOOD CALCIUM MEASUREMENT
C0729820|T059||CPT|BLOOD CALCIUM MEASUREMENT 
C0428613|T059||CPT|CALCIUM TO CREATININE RATIO MEASUREMENT
C0428613|T059||CPT|CALCIUM/CREATININE RATIO
C0428613|T059||CPT|CALCIUM/CREATININE RATIO 
C0428613|T059||CPT|CACREAT
C0428613|T059||CPT|CALCIUM/CREATININE
C0428613|T059||CPT|CALCIUM/CREATININE RATIO MEASUREMENT 
C0428613|T059||CPT|CALCIUM/CREATININE RATIO MEASUREMENT
C0523660|T059||CPT|GLUCOSE MEASUREMENT, POST GLUCOSE DOSE
C0523660|T059||CPT|GLUCOSE MEASUREMENT, POST GLUCOSE DOSE 
C0337438|T059|1011445|CPT|GLUCOSE|GLUCOSE
C0337438|T059|1011445|CPT|GLUCOSE MEASUREMENT|GLUCOSE
C0337438|T059|1011445|CPT|TEST;GLUCOSE|GLUCOSE
C0337438|T059|1011445|CPT|MEASUREMENT OF GLUCOSE|GLUCOSE
C0337438|T059|1011445|CPT|GLUC|GLUCOSE
C0337438|T059|1011445|CPT|GLUCOSE MEASUREMENT |GLUCOSE
C0337438|T059|1011445|CPT|GLUCOSE MEASUREMENT, NOS|GLUCOSE
C0337438|T059|1011445|CPT|GLUCOSE TEST|GLUCOSE
C0392201|T059|82947|CPT|BLOOD GLUCOSE|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|BLOOD GLUCOSE TESTS |BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|BLOOD GLUCOSE TESTS|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|BLOOD GLUCOSE MEASUREMENT|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|BLOOD GLUCOSE LEVEL|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|BLOOD GLUCOSE MEASUREMENT |BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|BLOOD GLUCOSE (SUGAR) LEVEL|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|MEASUREMENT OF GLUCOSE IN BLOOD|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|BLOOD SUGAR|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|GLUCOSE MEASUREMENT, BLOOD|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|BLOOD SUGAR LEVEL|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|BS - BLOOD GLUCOSE LEVEL|BLOOD GLUCOSE (SUGAR) LEVEL
C0392201|T059|82947|CPT|GLUCOSE MEASUREMENT, BLOOD |BLOOD GLUCOSE (SUGAR) LEVEL
C0202048|T059||CPT|GLUCOSE MEASUREMENT BY MONITORING DEVICE
C0202048|T059||CPT|GLUCOSE MEASUREMENT BY MONITORING DEVICE 
C0202048|T059||CPT|GLUCOSE MEASUREMENT BY MONITORING DEVICE  [AMBIGUOUS]
C2732668|T059||CPT|UREA, ELECTROLYTES AND GLUCOSE MEASUREMENT
C2732668|T059||CPT|MEASUREMENT OF UREA, SODIUM, POTASSIUM, CHLORIDE, BICARBONATE AND GLUCOSE 
C2732668|T059||CPT|MEASUREMENT OF UREA, SODIUM, POTASSIUM, CHLORIDE, BICARBONATE AND GLUCOSE
C2732640|T059||CPT|CALCULATION OF ESTIMATED AVERAGE GLUCOSE BASED ON HEMOGLOBIN A1C 
C2732640|T059||CPT|CALCULATION OF ESTIMATED AVERAGE GLUCOSE BASED ON HEMOGLOBIN A1C
C2732640|T059||CPT|ESTIMATED AVERAGE GLUCOSE MEASUREMENT
C2732640|T059||CPT|CALCULATION OF ESTIMATED AVERAGE GLUCOSE BASED ON HAEMOGLOBIN A1C
C0204885|T059||CPT|WARD GLUCOMETER TEST
C0204885|T059||CPT|WARD GLUCOMETER TEST 
C0202040|T059||CPT|CEREBROSPINAL FLUID GLUCOSE 
C0202040|T059||CPT|CEREBROSPINAL FLUID GLUCOSE
C0202040|T059||CPT|CSF GLUCOSE
C0202040|T059||CPT|GLUCOSE CSF
C0202040|T059||CPT|GLUCOSE MEASUREMENT, CEREBROSPINAL FLUID
C0202040|T059||CPT|GLUCOSE MEASUREMENT, CEREBROSPINAL FLUID 
C0202040|T059||CPT|GLUCOSE MEASUREMENT, CSF 
C0202040|T059||CPT|CSF GLUCOSE TEST
C0202040|T059||CPT|GLUCOSE MEASUREMENT, CSF
C1271625|T059||CPT|URINE CLINITEST
C1271625|T059||CPT|URINE CLINITEST 
C0202041|T059||CPT|SERUM GLUCOSE
C0202041|T059||CPT|SERUM GLUCOSE MEASUREMENT
C0202041|T059||CPT|SERUM GLUCOSE TEST
C0202041|T059||CPT|GLUCOSE MEASUREMENT, SERUM
C0202041|T059||CPT|GLUCOSE MEASUREMENT, SERUM 
C0202042|T059||CPT|PLASMA GLUCOSE MEASUREMENT
C0202042|T059||CPT|PLASMA GLUCOSE MEASUREMENT 
C0202042|T059||CPT|PLASMA GLUCOSE
C0202042|T059||CPT|PLASMA GLUCOSE LEVEL
C0202042|T059||CPT|PLASMA GLUCOSE LEVEL 
C0202042|T059||CPT|GLUCOSE MEASUREMENT, PLASMA
C0202042|T059||CPT|GLUCOSE MEASUREMENT, PLASMA 
C0523655|T059||CPT|GLUCOSE CEREBROSPINAL FLUID/GLUCOSE PLASMA RATIO MEASUREMENT 
C0523655|T059||CPT|GLUCOSE CEREBROSPINAL FLUID/GLUCOSE PLASMA RATIO MEASUREMENT
C0523655|T059||CPT|GLUCOSE CSF/GLUCOSE PLASMA RATIO MEASUREMENT 
C0523655|T059||CPT|GLUCOSE CSF/GLUCOSE PLASMA RATIO MEASUREMENT
C0004076|T059||CPT|URINE GLUCOSE
C0004076|T059||CPT|GLUCOSE MEASUREMENT, URINE
C0004076|T059||CPT|URINE GLUCOSE MEASUREMENT 
C0004076|T059||CPT|URINE GLUCOSE MEASUREMENT
C0004076|T059||CPT|GLUCOSE URINE
C0004076|T059||CPT|URINE SCREEN FOR SUGAR (& [GLUCOSE]) 
C0004076|T059||CPT|SUGAR - URINE TEST (& GLUCOSE)
C0004076|T059||CPT|URINE GLUCOSE TEST NOS
C0004076|T059||CPT|URINE GLUCOSE TEST NOS 
C0004076|T059||CPT|SUGAR - URINE TEST (& GLUCOSE) 
C0004076|T059||CPT|URINE TEST FOR GLUCOSE 
C0004076|T059||CPT|URINE SCREEN FOR SUGAR (& [GLUCOSE])
C0004076|T059||CPT|URINE TEST FOR GLUCOSE
C0004076|T059||CPT|GLUCOSE - URINE TEST
C0004076|T059||CPT|SUGAR - URINE TEST
C0004076|T059||CPT|URINE GLUCOSE TEST
C0004076|T059||CPT|GLUCOSE MEASUREMENT, URINE 
C0373621|T059|82950|CPT|GLUCOSE TEST; POST GLUCOSE DOSE (INCLUDES GLUCOSE)|BLOOD GLUCOSE (SUGAR) LEVEL AFTER RECEIVING DOSE OF GLUCOSE
C0373621|T059|82950|CPT|GLUCOSE; POST GLUCOSE DOSE (INCLUDES GLUCOSE)|BLOOD GLUCOSE (SUGAR) LEVEL AFTER RECEIVING DOSE OF GLUCOSE
C0373621|T059|82950|CPT|GLUCOSE POST GLUCOSE DOSE|BLOOD GLUCOSE (SUGAR) LEVEL AFTER RECEIVING DOSE OF GLUCOSE
C0373621|T059|82950|CPT|BLOOD GLUCOSE (SUGAR) LEVEL AFTER RECEIVING DOSE OF GLUCOSE|BLOOD GLUCOSE (SUGAR) LEVEL AFTER RECEIVING DOSE OF GLUCOSE
C0373621|T059|82950|CPT|MEASUREMENT OF GLUCOSE AFTER GLUCOSE DOSE|BLOOD GLUCOSE (SUGAR) LEVEL AFTER RECEIVING DOSE OF GLUCOSE
C0373621|T059|82950|CPT|GLUCOSE TEST|BLOOD GLUCOSE (SUGAR) LEVEL AFTER RECEIVING DOSE OF GLUCOSE
C0523658|T059|82947|CPT|ASSAY GLUCOSE BLOOD QUANT|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T059|82947|CPT|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T059|82947|CPT|GLUCOSE QUANTITATIVE BLOOD XCPT REAGENT STRIP|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T059|82947|CPT|GLUCOSE MEASUREMENT, QUANTITATIVE|GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0523658|T059|82947|CPT|GLUCOSE MEASUREMENT, QUANTITATIVE |GLUCOSE; QUANTITATIVE, BLOOD (EXCEPT REAGENT STRIP)
C0373622|T059|82951|CPT|GLUCOSE; TOLERANCE TEST (GTT), 3 SPECIMENS (INCLUDES GLUCOSE)|GLUCOSE TOLERANCE TEST GTT 3 SPECIMENS
C0373622|T059|82951|CPT|GLUCOSE TOLERANCE TEST GTT 3 SPECIMENS|GLUCOSE TOLERANCE TEST GTT 3 SPECIMENS
C0373622|T059|82951|CPT|GLUCOSE TOLERANCE TEST (GTT)|GLUCOSE TOLERANCE TEST GTT 3 SPECIMENS
C0373623|T059|82952|CPT|GLUCOSE TOLERANCE EA ADDL BEYOND 3 SPECIMENS|GLUCOSE TOLERANCE EA ADDL BEYOND 3 SPECIMENS
C0373623|T059|82952|CPT|GLUCOSE; TOLERANCE TEST, EACH ADDITIONAL BEYOND 3 SPECIMENS (LIST SEPARATELY IN ADDITION TO CODE FOR PRIMARY PROCEDURE)|GLUCOSE TOLERANCE EA ADDL BEYOND 3 SPECIMENS
C0373623|T059|82952|CPT|GTT-ADDED SAMPLES|GLUCOSE TOLERANCE EA ADDL BEYOND 3 SPECIMENS
C0373620|T059|82948|CPT|GLUCOSE; BLOOD, REAGENT STRIP|MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP
C0373620|T059|82948|CPT|BLOOD GLUCOSE DETERMINATION BY REAGENT STRIP |MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP
C0373620|T059|82948|CPT|BLOOD GLUCOSE DETERMINATION BY REAGENT STRIP|MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP
C0373620|T059|82948|CPT|BLOOD GLUCOSE LEVEL BY REAGENT STRIP|MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP
C0373620|T059|82948|CPT|GLUCOSE BLOOD REAGENT STRIP|MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP
C0373620|T059|82948|CPT|BLOOD GLUCOSE (SUGAR) MEASUREMENT USING REAGENT STRIP|MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP
C0373620|T059|82948|CPT|MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP|MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP
C0373620|T059|82948|CPT|REAGENT STRIP/BLOOD GLUCOSE|MEASUREMENT OF GLUCOSE IN BLOOD USING REAGENT STRIP
C4064987|T059||CPT|GLUCOSE IN SERUM OR PLASMA 
C4064987|T059||CPT|GLUCOSE IN SERUM OR PLASMA
C0202045|T059||CPT|GLUCOSE MEASUREMENT, FASTING
C0202045|T059||CPT|GLUCOSE MEASUREMENT, FASTING 
C0202045|T059||CPT|FASTING GLUCOSE TEST
C0202045|T059||CPT|TEST;GLUCOSE;FASTING
C0202046|T059||CPT|GLUCOSE MEASUREMENT, RANDOM
C0202046|T059||CPT|GLUCOSE MEASUREMENT, RANDOM 
C0202046|T059||CPT|RANDOM GLUCOSE TEST
C0202046|T059||CPT|TEST;GLUCOSE;RANDOM
C0017741|T059|82951|CPT|GLUCOSE TOLERANCE TEST|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|GLUCOSE TOLERANCE TESTS|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|TEST;GLUCOSE TOLERANCE|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|GLUCOSE TOLERANCE TEST (GTT)|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|GLUCOSE TOLERANCE TEST NOS|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|GLUCOSE TOLERANCE TEST NOS |BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|GTT|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|GTT - GLUCOSE TOLERANCE TEST|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|OGTT - ORAL GLUCOSE TOLERANCE TEST|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|GLUCOSE CHALLENGE TEST|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|GLUCOSE TOLERANCE TEST |BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0017741|T059|82951|CPT|GLUCOSE TOLERANCE TEST, NOS|BLOOD GLUCOSE (SUGAR) TOLERANCE TEST
C0523657|T059||CPT|GLUCOSE MEASUREMENT, TOLBUTAMIDE TOLERANCE TEST
C0523657|T059||CPT|GLUCOSE MEASUREMENT, TOLBUTAMIDE TOLERANCE TEST 
C1272314|T059||CPT|FECAL CLINITEST 
C1272314|T059||CPT|FAECAL CLINITEST 
C1272314|T059||CPT|FAECAL CLINITEST
C1272314|T059||CPT|FECAL CLINITEST
C0427743|T059||CPT|GLUCOSE CONCENTRATION
C0427743|T059||CPT|GLUCOSE CONCENTRATION, TEST STRIP MEASUREMENT 
C0427743|T059||CPT|GLUCOSE CONCENTRATION, TEST STRIP MEASUREMENT
C1295145|T059||CPT|GLUCOSE MEASUREMENT ESTIMATED FROM GLYCATED HAEMOGLOBIN
C1295145|T059||CPT|GLUCOSE MEASUREMENT ESTIMATED FROM GLYCATED HEMOGLOBIN 
C1295145|T059||CPT|GLUCOSE MEASUREMENT ESTIMATED FROM GLYCATED HEMOGLOBIN
C0428549|T059||CPT|FLUID SAMPLE GLUCOSE MEASUREMENT
C0428549|T059||CPT|BODY FLUID GLUCOSE MEASUREMENT 
C0428549|T059||CPT|BODY FLUID GLUCOSE
C0428549|T059||CPT|BODY FLUID GLUCOSE MEASUREMENT
C0428549|T059||CPT|MEASUREMENT OF GLUCOSE IN BODY FLUID
C0428549|T059||CPT|BODY FLUID GLUCOSE TEST
C0428549|T059||CPT|FLUID SAMPLE GLUCOSE LEVEL
C0428549|T059||CPT|FLUID SAMPLE GLUCOSE MEASUREMENT 
C0428549|T059||CPT|GLUCOSE MEASUREMENT, BODY FLUID
C1319276|T059||CPT|FAECAL GLUCOSE LEVEL
C1319276|T059||CPT|FAECAL GLUCOSE MEASUREMENT
C1319276|T059||CPT|FECAL GLUCOSE LEVEL 
C1319276|T059||CPT|FECAL GLUCOSE LEVEL
C1319276|T059||CPT|FECAL GLUCOSE MEASUREMENT
C0201850|T059|84075|CPT|ALKALINE PHOSPHATASE MEASUREMENT|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|PHOSPHATASE, ALKALINE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALP|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|TEST;ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|MEASUREMENT OF ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ASSAY OF PHOSPHATASE ALKALINE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALK PHOSPH|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALK PHOS|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALKALINE PHOSPHATASE MEASUREMENT |ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ASSAY ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE
C0201850|T059|84075|CPT|ALKALINE PHOSPHATASE TEST|ASSAY OF PHOSPHATASE ALKALINE
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE
C0036776|T059||CPT|SAP
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE MEASUREMENT
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE MEASUREMENT 
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE (& LEVEL)
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE (& LEVEL) 
C0036776|T059||CPT|ALK. PHOSPHATASE -SERUM
C0036776|T059||CPT|ALKALINE PHOSPHATASE (& LEVEL (& SERUM))
C0036776|T059||CPT|PHOSPH.- ALK. - SERUM
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE NOS
C0036776|T059||CPT|ALKALINE PHOSPHATASE (& LEVEL (& SERUM)) 
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE NOS 
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE TEST
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE LEVEL
C0036776|T059||CPT|SERUM ALKALINE PHOSPHATASE MEASUREMENT 
C1293930|T059||CPT|MEASUREMENT OF RATIO OF ANALYTE TO ALKALINE PHOSPHATASE 
C1293930|T059||CPT|MEASUREMENT OF RATIO OF ANALYTE TO ALKALINE PHOSPHATASE
C0201851|T059|84080|CPT|PHOSPHATASE, ALKALINE; ISOENZYMES|ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES
C0201851|T059|84080|CPT|MEASUREMENT OF ALKALINE PHOSPHATASE ISOENZYMES|ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES
C0201851|T059|84080|CPT|ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES|ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES
C0201851|T059|84080|CPT|ALKALINE PHOSPHATASE ISOENZYMES MEASUREMENT|ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES
C0201851|T059|84080|CPT|ALKALINE PHOSPHATASE ISOENZYMES MEASUREMENT |ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES
C0201851|T059|84080|CPT|ASSAY ALKALINE PHOSPHATASES|ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES
C0201855|T059|84078|CPT|ALKALINE PHOSPHATASE, HEAT STABLE MEASUREMENT|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C0201855|T059|84078|CPT|PHOSPHATASE, ALKALINE; HEAT STABLE (TOTAL NOT INCLUDED)|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C0201855|T059|84078|CPT|MEASUREMENT OF HEAT STABLE ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C0201855|T059|84078|CPT|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C0201855|T059|84078|CPT|THERMOSTABLE ALKALINE PHOSPHATASE MEASUREMENT|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C0201855|T059|84078|CPT|ALKALINE PHOSPHATASE, HEAT STABLE MEASUREMENT |ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C0201855|T059|84078|CPT|ASSAY ALKALINE PHOSPHATASE|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C2984961|T059||CPT|BONE SPECIFIC ALKALINE PHOSPHATASE MEASUREMENT
C2984961|T059||CPT|BONE ALKALINE PHOSPHATASE MEASUREMENT
C2984961|T059||CPT|BONE SPECIFIC ALKALINE PHOSPHATASE
C2984961|T059||CPT|ALPBS
C2984961|T059||CPT|BONE ALP MEASUREMENT
C3898585|T059||CPT|LIVER SPECIFIC ALKALINE PHOSPHATASE MEASUREMENT
C3898585|T059||CPT|ALPLS
C3898585|T059||CPT|LIVER SPECIFIC ALKALINE PHOSPHATASE
C3898710|T059||CPT|INTESTINAL SPECIFIC ALKALINE PHOSPHATASE
C3898710|T059||CPT|ALPIS
C3898710|T059||CPT|INTESTINAL SPECIFIC ALKALINE PHOSPHATASE MEASUREMENT
C0200697|T059||CPT|LEUKOCYTE ALKALINE PHOSPHATASE LEVEL
C0200697|T059||CPT|LEUCOCYTE ALKALINE PHOSPHATASE LEVEL
C0200697|T059||CPT|LEUCOCYTE ALKALINE PHOSPHATASE LEVEL 
C0200697|T059||CPT|LEUKOCYTE ALKALINE PHOSPHATASE SCORE
C0200697|T059||CPT|LEUCOCYTE ALKALINE PHOSPHATASE SCORE
C0200697|T059||CPT|LEUKOCYTE ALKALINE PHOSPHATASE SCORE 
C0200697|T059||CPT|LEUKOCYTE ALKALINE PHOSPHATASE SCORE (OBSERVABLE ENTITY)
C0200697|T059||CPT|NEUTROPHIL ALKALINE PHOSPHATASE SCORE
C0200697|T059||CPT|LAP SCORE
C0200697|T059||CPT|LAP - NEUTROPHIL ALKALINE PHOSPHATASE SCORE
C0200697|T059||CPT|LAP - NEUTROPHIL ALKALINE PHOSPHATASE SCORE MEASUREMENT
C0201852|T059||CPT|PLACENTAL ALKALINE PHOSPHATASE MEASUREMENT
C0201852|T059||CPT|PLAP MEASUREMENT
C0201852|T059||CPT|PLACENTAL ALKALINE PHOSPHATASE MEASUREMENT 
C0201853|T059||CPT|INTESTINAL ALKALINE PHOSPHATASE MEASUREMENT
C0201853|T059||CPT|IAP MEASUREMENT
C0201853|T059||CPT|INTESTINAL ALKALINE PHOSPHATASE MEASUREMENT 
C0201854|T059||CPT|GERM CELL ALKALINE PHOSPHATASE MEASUREMENT
C0201854|T059||CPT|GCAP MEASUREMENT
C0201854|T059||CPT|GERM CELL ALKALINE PHOSPHATASE MEASUREMENT 
C0428333|T059||CPT|FLUID SAMPLE ALKALINE PHOSPHATASE LEVEL
C0428333|T059||CPT|FLUID SAMPLE ALKALINE PHOSPHATASE MEASUREMENT 
C0428333|T059||CPT|FLUID SAMPLE ALKALINE PHOSPHATASE MEASUREMENT
C1272113|T059||CPT|PLASMA ALKALINE PHOSPHATASE LEVEL 
C1272113|T059||CPT|PLASMA ALKALINE PHOSPHATASE LEVEL
C0391938|T059|82435|CPT|CHLORIDE; BLOOD|CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE|CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE LEVEL|CHLORIDE BLD
C0391938|T059|82435|CPT|MEASUREMENT OF CHLORIDE IN BLOOD|CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE LEVEL |CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE LEVEL |CHLORIDE BLD
C0391938|T059|82435|CPT|CHLORIDE MEASUREMENT, BLOOD|CHLORIDE BLD
C0391938|T059|82435|CPT|CHLORIDE MEASUREMENT, BLOOD |CHLORIDE BLD
C0391938|T059|82435|CPT|ASSAY OF BLOOD CHLORIDE|CHLORIDE BLD
C0391938|T059|82435|CPT|BLOOD CHLORIDE LEVEL MEASUREMENT|CHLORIDE BLD
C0391938|T059|82435|CPT|CHLORIDE BLD|CHLORIDE BLD
C1317978|T059|82438|CPT|SERUM CHLORIDE MEASUREMENT|CHLORIDE LEVEL
C1317978|T059|82438|CPT|SERUM CHLORIDE MEASUREMENT |CHLORIDE LEVEL
C1317978|T059|82438|CPT|CHLORIDE LEVEL|CHLORIDE LEVEL
C1317978|T059|82438|CPT|SERUM CHLORIDE (& LEVEL)|CHLORIDE LEVEL
C1317978|T059|82438|CPT|SERUM CHLORIDE (& LEVEL) |CHLORIDE LEVEL
C1317978|T059|82438|CPT|SERUM CHLORIDE LEVEL|CHLORIDE LEVEL
C1317978|T059|82438|CPT|SERUM CHLORIDE MEASUREMENT |CHLORIDE LEVEL
C2711521|T059||CPT|MEASUREMENT OF CHLORIDE IN STOOL SPECIMEN 
C2711521|T059||CPT|MEASUREMENT OF CHLORIDE IN STOOL SPECIMEN
C2732591|T059||CPT|UREA, ELECTROLYTES AND CREATININE MEASUREMENT
C2732591|T059||CPT|MEASUREMENT OF UREA, SODIUM, POTASSIUM, CHLORIDE, BICARBONATE AND CREATININE
C2732591|T059||CPT|MEASUREMENT OF UREA, SODIUM, POTASSIUM, CHLORIDE, BICARBONATE AND CREATININE 
C2732591|T059||CPT|LAB-BASED CHEM MEASURE UREA, NA, POTASSIUM CHLORIDE, BICARBONATE, CREATININE
C2732591|T059||CPT|MEASUREMENT OF UREA, SODIUM, POTASSIUM CHLORIDE, BICARBONATE, AND CREATININE
C2732591|T059||CPT|MEASUREMENT OF UREA, SODIUM, POTASSIUM CHLORIDE, BICARBONATE, AND CREATININE 
C0729818|T059||CPT|BLOOD CHLORIDE LEVEL RESULT
C0428295|T059||CPT|SWEAT TEST FOR CHLORIDE 
C0428295|T059||CPT|SWEAT TEST FOR CHLORIDE
C0428295|T059||CPT|SWEAT CHLORIDE (& LEVEL) 
C0428295|T059||CPT|SWEAT CHLORIDE (& LEVEL)
C0428295|T059||CPT|SWEAT CHLORIDE
C0428295|T059||CPT|SWEAT CHLORIDE TEST
C0428295|T059||CPT|CHLORIDE SWEAT TEST
C0428295|T059||CPT|CYSTIC FIBROSIS SWEAT TEST
C0428295|T059||CPT|CHLORIDE MEASUREMENT, SWEAT
C0428295|T059||CPT|SWEAT CHLORIDE LEVEL
C0428295|T059||CPT|CYSTIC FIBROSIS SWEAT TEST 
C0201953|T059|82436|CPT|CHLORIDE; URINE|URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|URINE CHLORIDE MEASUREMENT |URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|URINE CHLORIDE MEASUREMENT|URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|URINE CHLORIDE|URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|URINE CHLORIDE LEVEL|URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|MEASUREMENT OF CHLORIDE IN URINE|URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|URINE CHLORIDE LEVEL |URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|URINE CHLORIDE TEST|URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|CHLORIDE MEASUREMENT, URINE|URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|CHLORIDE MEASUREMENT, URINE |URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|ASSAY OF URINE CHLORIDE|URINE CHLORIDE LEVEL
C0201953|T059|82436|CPT|CHLORIDE URINE|URINE CHLORIDE LEVEL
C0373575|T059|82438|CPT|CHLORIDE; OTHER SOURCE|ASSAY OTHER FLUID CHLORIDES
C0373575|T059|82438|CPT|ASSAY OTHER FLUID CHLORIDES|ASSAY OTHER FLUID CHLORIDES
C0373575|T059|82438|CPT|CHLORIDE OTHER SOURCE|ASSAY OTHER FLUID CHLORIDES
C3830082|T059||CPT|FRACTIONAL EXCRETION OF CHLORIDE
C3830082|T059||CPT|FRACTIONAL CHLORIDE EXCRETION
C3830082|T059||CPT|FECL
C3830082|T059||CPT|FRACTIONAL EXCRETION OF CL
C0201952|T059|1011335|CPT|CHLORIDE MEASUREMENT|CHLORIDE
C0201952|T059|1011335|CPT|MEASUREMENT OF CHLORIDE|CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE|CHLORIDE
C0201952|T059|1011335|CPT|CL|CHLORIDE
C0201952|T059|1011335|CPT|CL-|CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE MEASUREMENT |CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE MEASUREMENT, NOS|CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE EACH TEST|CHLORIDE
C0201952|T059|1011335|CPT|CHLORIDE EA.TST|CHLORIDE
C0428297|T059||CPT|CSF CHLORIDE MEASUREMENT 
C0428297|T059||CPT|CSF: CHLORIDE LEVEL NOS 
C0428297|T059||CPT|CEREBROSPINAL FLUID CHLORIDE MEASUREMENT 
C0428297|T059||CPT|CEREBROSPINAL FLUID CHLORIDE MEASUREMENT
C0428297|T059||CPT|CSF CL
C0428297|T059||CPT|CSF CHLORIDE
C0428297|T059||CPT|CSF CHLORIDE LEVEL
C0428297|T059||CPT|CEREBROSPINAL FLUID CHLORIDE MEASUREMENT 
C0428297|T059||CPT|CEREBROSPINAL FLUID: CHLORIDE LEVEL NOS 
C0428297|T059||CPT|CEREBROSPINAL FLUID: CHLORIDE LEVEL NOS
C0428297|T059||CPT|CSF: CHLORIDE LEVEL NOS
C0428297|T059||CPT|CSF CHLORIDE TEST
C0428297|T059||CPT|CSF: CHLORIDE LEVEL
C0428297|T059||CPT|CSF CHLORIDE MEASUREMENT
C0428296|T059||CPT|BODY FLUID CHLORIDE TEST
C0428296|T059||CPT|FLUID SAMPLE CHLORIDE
C0428296|T059||CPT|FLUID SAMPLE CHLORIDE LEVEL
C0428296|T059||CPT|CHLORIDE MEASUREMENT, BODY FLUID 
C0428296|T059||CPT|CHLORIDE MEASUREMENT, BODY FLUID
C0428296|T059||CPT|BODY FLUID CHLORIDE MEASUREMENT
C0428296|T059||CPT|CHLORIDE MEASUREMENT, BODY FLUID, NOS
C1276037|T059||CPT|PLASMA CHLORIDE LEVEL
C1276037|T059||CPT|PLASMA CHLORIDE MEASUREMENT 
C1276037|T059||CPT|PLASMA CHLORIDE MEASUREMENT
C0430179|T059||CPT|SWEAT TEST
C0430179|T059||CPT|SWEAT TEST NOS
C0430179|T059||CPT|SWEAT TEST 
C0430179|T059||CPT|SWEAT TEST NOS 
C0430179|T059||CPT|SWEAT TESTS
C0430179|T059||CPT|SWEAT TESTS 
C0430179|T059||CPT|SWEAT SCREENING TEST
C0201975|T059|82565|CPT|CREATININE MEASUREMENT|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE; BLOOD|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|BLOOD CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|TEST;CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE BLOOD|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|BLOOD CREATININE LEVEL|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|MEASUREMENT OF CREATININE|BLOOD CREATININE LEVEL
# C0201975|T059|82565|CPT|CR|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|LAB-BASED CHEM MEASUREMENTS CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|MEASUREMENT OF CREATININE |BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREAT|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|BLOOD CREATININE LEVEL |BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE MEASUREMENT |BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE MEASUREMENT, NOS|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|ASSAY OF CREATININE|BLOOD CREATININE LEVEL
C0201975|T059|82565|CPT|CREATININE TEST|BLOOD CREATININE LEVEL
C2981749|T059||CPT|URINARY CREATININE ASSAY
C2981751|T059||CPT|SERUM CREATININE ASSAY
C0201976|T059||CPT|SERUM CREATININE
C0201976|T059||CPT|SERUM CREATININE MEASUREMENT
C0201976|T059||CPT|CREATININE MEASUREMENT, SERUM 
C0201976|T059||CPT|SERUM CREATININE LEVEL
C0201976|T059||CPT|SERUM CREATININE MEASUREMENT 
C0201976|T059||CPT|CREATININE.SERUM
C0201976|T059||CPT|SERUM CREATININE (& LEVEL) 
C0201976|T059||CPT|CREATININE - SERUM
C0201976|T059||CPT|SERUM CREATININE NOS 
C0201976|T059||CPT|SERUM CREATININE NOS
C0201976|T059||CPT|SERUM CREATININE (& LEVEL)
C0201976|T059||CPT|SERUM CREATININE TEST
C0201976|T059||CPT|CREATININE MEASUREMENT, SERUM
C1278055|T059||CPT|PLASMA CREATININE MEASUREMENT
C1278055|T059||CPT|PLASMA CREATININE LEVEL
C1278055|T059||CPT|PLASMA CREATININE LEVEL 
C1278055|T059||CPT|PLASMA CREATININE
C1278055|T059||CPT|PLASMA CREATININE MEASUREMENT 
C1278055|T059||CPT|PLASMA CREATININE MEASUREMENT 
C1318439|T059||CPT|URINE CREATININE MEASUREMENT
C1318439|T059||CPT|URINE CREATININE MEASUREMENT 
C1318439|T059||CPT|URINE CREATININE
C1318439|T059||CPT|CREATININE LEVEL
C1318439|T059||CPT|CREATININE URINE
C1318439|T059||CPT|URINE CREATININE (& LEVEL) 
C1318439|T059||CPT|URINE CREATININE (& LEVEL)
C1318439|T059||CPT|CREATININE - URINE
C1318439|T059||CPT|CREATININE MEASUREMENT, URINE
C1318439|T059||CPT|URINE CREATININE MEASUREMENT 
C1318439|T059||CPT|URINE CREATININE LEVEL
C0201977|T059||CPT|URINE CREATININE 12-HOUR
C0201977|T059||CPT|12-HOUR URINE CREATININE MEASUREMENT
C0201977|T059||CPT|12-HOUR URINE CREATININE MEASUREMENT 
C0201977|T059||CPT|12-HOUR CREATININE LEVEL
C0201977|T059||CPT|CREATININE MEASUREMENT, 12 HOUR URINE
C0201977|T059||CPT|CREATININE MEASUREMENT, 12 HOUR URINE 
C3694999|T059||CPT|CREATININE CONCENTRATION (SERUM OR PLASMA)
C3694999|T059||CPT|SERUM OR PLASMA CREATININE CONCENTRATION 
C3694999|T059||CPT|SERUM OR PLASMA CREATININE CONCENTRATION
C3694393|T059||CPT|LAB-BASED CHEM MEASUREMENTS CREATININE CLEARANCE - GLOMERULAR FILTRATION 
C3694393|T059||CPT|LAB-BASED CHEM MEASUREMENTS CREATININE CLEARANCE - GLOMERULAR FILTRATION
C0373594|T059|82570|CPT|CREATININE; OTHER SOURCE|ASSAY OF URINE CREATININE
C0373594|T059|82570|CPT|CREATININE OTHER SOURCE|ASSAY OF URINE CREATININE
C0373594|T059|82570|CPT|ASSAY OF URINE CREATININE|ASSAY OF URINE CREATININE
C0373595|T059|82575|CPT|CREATININE; CLEARANCE|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE RENAL CLEARANCE|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|MEASUREMENT OF RENAL CLEARANCE OF CREATININE|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE CLEARANCE TEST|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE CLEARANCE TEST |CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|MEASUREMENT OF RENAL CLEARANCE OF CREATININE |CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE CLEARANCE MEASUREMENT|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE RENAL CLEARANCE MEASUREMENT |CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE CLEARANCE-GLOM FILT|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE CLEARANCE STUDY |CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE RENAL CLEARANCE MEASUREMENT|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE CLEARANCE|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE CLEARANCE STUDY|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATCLR|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|RENAL FUNCTION CREATININE CLEARANCE|CREATININE CLEARANCE TEST
C0373595|T059|82575|CPT|CREATININE RENAL CLEARANCE |CREATININE CLEARANCE TEST
C0428279|T059||CPT|FINDING OF CREATININE LEVEL
C0428279|T059||CPT|LAB-BASED CHEM MEASUREMENTS CREATININE LEVEL FINDING
C0428279|T059||CPT|CREATININE LEVEL FINDING 
C0428279|T059||CPT|CREATININE LEVEL FINDING
C0428279|T059||CPT|CREATININE LEVEL
C0428279|T059||CPT|CREATININE LEVEL - FINDING
C0428279|T059||CPT|FINDING OF CREATININE LEVEL 
C0523586|T059||CPT|CREATININE CHALLENGE TESTS
C0523586|T059||CPT|CREATININE CHALLENGE TESTS 
C1278053|T059||CPT|CORRECTED PLASMA CREATININE LEVEL
C1278053|T059||CPT|CORRECTED PLASMA CREATININE LEVEL 
C1278053|T059||CPT|CORRECTED PLASMA CREATININE MEASUREMENT 
C1278053|T059||CPT|CORRECTED PLASMA CREATININE MEASUREMENT
C1261396|T059||CPT|FLUID SAMPLE CREATININE MEASUREMENT
C1261396|T059||CPT|BODY FLUID CREATININE TEST
C1261396|T059||CPT|CREATININE MEASUREMENT, BODY FLUID
C1261396|T059||CPT|FLUID SAMPLE CREATININE MEASUREMENT 
C1261396|T059||CPT|FLUID SAMPLE CREATININE LEVEL
C1293927|T059||CPT|MEASUREMENT OF RATIO OF ANALYTE TO CREATININE 
C1293927|T059||CPT|MEASUREMENT OF RATIO OF ANALYTE TO CREATININE
C1446045|T059||CPT|5-HYDROXYINDOLEACETIC ACID/CREATININE RATIO MEASUREMENT 
C1446045|T059||CPT|5-HYDROXYINDOLEACETIC ACID/CREATININE RATIO MEASUREMENT
C1446045|T059||CPT|5HIAA/CREATININE RATIO
C1446063|T059||CPT|AMINOLAEVULINIC ACID / CREATININE RATIO MEASUREMENT
C1446063|T059||CPT|AMINOLAEVULINIC ACID/CREATININE RATIO MEASUREMENT
C1446063|T059||CPT|AMINOLEVULINIC ACID / CREATININE RATIO MEASUREMENT
C1446063|T059||CPT|AMINOLEVULINIC ACID/CREATININE RATIO MEASUREMENT 
C1446063|T059||CPT|AMINOLEVULINIC ACID/CREATININE RATIO MEASUREMENT
C1446063|T059||CPT|ALA/CREATININE RATIO
C1446080|T059||CPT|MAGNESIUM TO CREATININE RATIO MEASUREMENT
C1446080|T059||CPT|MAGNESIUM/CREATININE
C1446080|T059||CPT|MGCREAT
C1446080|T059||CPT|MAGNESIUM / CREATININE RATIO MEASUREMENT 
C1446080|T059||CPT|MAGNESIUM / CREATININE RATIO MEASUREMENT
C1446080|T059||CPT|MAGNESIUM/CREATININE RATIO
C1446178|T059||CPT|RETINOL BINDING PROTEIN / CREATININE RATIO MEASUREMENT 
C1446178|T059||CPT|RETINOL BINDING PROTEIN / CREATININE RATIO MEASUREMENT
C1531635|T059||CPT|CITRATE:CREATININE RATIO 
C1531635|T059||CPT|CITRATE:CREATININE RATIO
C1531635|T059||CPT|MEASUREMENT OF RATIO OF CITRATE TO CREATININE 
C1531635|T059||CPT|MEASUREMENT OF RATIO OF CITRATE TO CREATININE
C1531635|T059||CPT|MEAUSREMENT OF RATIO OF CITRATE TO CREATININE
C1531635|T059||CPT|MEAUSREMENT OF RATIO OF CITRATE TO CREATININE 
C1531635|T059||CPT|CITRATE/CREATININE
C1531635|T059||CPT|CITRATE TO CREATININE RATIO MEASUREMENT
C1531635|T059||CPT|CITRIC ACID/CREATININE
C1531635|T059||CPT|CITCREAT
C0596252|T059||CPT|CARBON DIOXIDE FIXATION
C0596253|T059||CPT|CARBON DIOXIDE TENSION
C0596254|T059||CPT|CARBON DIOXIDE TRANSPORT
C0201930|T059|82374|CPT|CARBON DIOXIDE CONTENT MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CO2 CONTENT MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|PCO2, BLOOD|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CO<SUB>2</SUB> CONTENT MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|PCO<SUB>2</SUB>, BLOOD|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE (BICARBONATE)|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|ASSAY BLOOD CARBON DIOXIDE|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE BICARBONATE|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|MEASUREMENT OF CARBON DIOXIDE|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CO2|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|PCO>2<, BLOOD|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CO>2< CONTENT MEASUREMENT|ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE CONTENT MEASUREMENT |ASSAY BLOOD CARBON DIOXIDE
C0201930|T059|82374|CPT|CARBON DIOXIDE MEASUREMENT |ASSAY BLOOD CARBON DIOXIDE
C2144939|T059||CPT|SERUM TOTAL CO2
C2144939|T059||CPT|SERUM TOTAL CO2 
C2144939|T059||CPT|TOTAL CO2 CONTENT
C0201931|T059||CPT|PARTIAL PRESSURE OF CARBON DIOXIDE MEASUREMENT
C0201931|T059||CPT|CARBON DIOXIDE MEASUREMENT, PARTIAL PRESSURE
C0201931|T059||CPT|PCO2
C0201931|T059||CPT|PARTIAL PRESSURE CARBON DIOXIDE
C0201931|T059||CPT|PACO2 MEASUREMENT
C0201931|T059||CPT|CARBON DIOXIDE MEASUREMENT, PARTIAL PRESSURE 
C0005845|T059|84520|CPT|BLOOD UREA NITROGEN|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BUN|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|NITROGEN, BLOOD UREA|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|UREA NITROGEN, BLOOD|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA NITROGEN MEASUREMENT|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|UREA NITROGEN; QUANTITATIVE|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BUN LEVEL|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|MEASUREMENT OF BLOOD UREA NITROGEN (BUN)|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|ASSAY OF UREA NITROGEN QUANTITATIVE|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|MEASUREMENT OF UREA NITROGEN (BUN)|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|UREA - BLOOD|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA |ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA NITROGEN MEASUREMENT |ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BUN MEASUREMENT|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA MEASUREMENT |ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA MEASUREMENT|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|BLOOD UREA NITROGEN MEASUREMENT |ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|T059|84520|CPT|ASSAY OF UREA NITROGEN|ASSAY OF UREA NITROGEN QUANTITATIVE
C0455273|T059||CPT|SERUM UREA LEVEL
C0455273|T059||CPT|SERUM UREA LEVEL 
C0455273|T059||CPT|SERUM UREA MEASUREMENT 
C0455273|T059||CPT|SERUM UREA MEASUREMENT
C0729828|T059||CPT|PLASMA UREA LEVEL
C0729828|T059||CPT|PLASMA UREA LEVEL 
C0729828|T059||CPT|PLASMA UREA MEASUREMENT 
C0729828|T059||CPT|PLASMA UREA MEASUREMENT
C0201922|T059||CPT|BUN/CREATININE RATIO 
C0201922|T059||CPT|BLOOD UREA NITROGEN (BUN)/CREATININE RATIO
C0201922|T059||CPT|BLOOD UREA NITROGEN/CREATININE RATIO 
C0201922|T059||CPT|BLOOD UREA NITROGEN/CREATININE RATIO
C0201922|T059||CPT|BLOOD UREA NITROGEN (BUN)/CREATININE RATIO 
C0201922|T059||CPT|BUN/CREATININE RATIO
C0201922|T059||CPT|BUN/CREATININE RATIO 
C0201922|T059||CPT|UREA NITROGEN/CREATININE RATIO, SERUM
C2208743|T059||CPT|SERUM BUN/CREATININE RATIO
C2208743|T059||CPT|SERUM BUN/CREATININE RATIO 
C2097174|T059||CPT|BUN USING REAGENT STRIP 
C2097174|T059||CPT|BUN USING REAGENT STRIP
C2097174|T059||CPT|BUN BY REAGENT STRIP
C2097689|T059||CPT|BUN WAS OBTAINED PRE-PROCEDURE
C2097689|T059||CPT|BUN WAS OBTAINED PRE-PROCEDURE 
C2097689|T059||CPT|A BUN LEVEL WAS OBTAINED PRE-PROCEDURE
C0729816|T059|84132|CPT|BLOOD POTASSIUM LEVEL|BLOOD POTASSIUM LEVEL
C0729816|T059|84132|CPT|BLOOD POTASSIUM LEVEL |BLOOD POTASSIUM LEVEL
C0729816|T059|84132|CPT|BLOOD POTASSIUM MEASUREMENT |BLOOD POTASSIUM LEVEL
C0729816|T059|84132|CPT|BLOOD POTASSIUM MEASUREMENT|BLOOD POTASSIUM LEVEL
C4027477|T059||CPT|UREA NITROGEN LEVEL IN SERUM OR PLASMA 
C4027477|T059||CPT|UREA NITROGEN LEVEL IN SERUM OR PLASMA
C0200379|T059|80050|CPT|GENERAL HEALTH PANEL|GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)
C0200379|T059|80050|CPT|GENERAL HEALTH PANEL |GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)
C0200379|T059|80050|CPT|GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)|GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)
C0200379|T059|80050|CPT|GENERAL HEALTH PANEL, NOS|GENERAL HEALTH PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: COMPREHENSIVE METABOLIC PANEL (80053) BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) THYROID STIMULATING HORMONE (TSH) (84443)
C0201836|T059|84460|CPT|ALANINE AMINOTRANSFERASE MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALANINE AMINOTRANSFERASE|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
# C0201836|T059|84460|CPT|ALT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|TRANSFERASE; ALANINE AMINO (ALT) (SGPT)|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|TEST;ALANINE AMINOTRANSFERASE|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|TRANSFERASE ALANINE AMINO ALT SGPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|LIVER ENZYME (SGPT), LEVEL|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALANINE AMINO (ALT) (SGPT)|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|SGPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|GLUTAMIC-PYRUVATE TRANSAMINASE|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|GPT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|GPT MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|GLUTAMIC PYRUVATE TRANSAMINASE MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|SGPT MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALT MEASUREMENT|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALANINE AMINOTRANSFERASE MEASUREMENT |MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C0201836|T059|84460|CPT|ALANINE AMINOTRANSFERASE TEST|MEASUREMENT OF ALANINE AMINO TRANSFERASE (ALT) (SGPT)
C1883008|T059||CPT|SERUM ALANINE AMINOTRANSFERASE MEASUREMENT
C1883008|T059||CPT|SERUM SGPT MEASUREMENT
C1883008|T059||CPT|SERUM ALANINE TRANSAMINASE MEASUREMENT
C1883008|T059||CPT|SERUM ALANINE AMINOTRANSFERASE MEASUREMENT 
C1883008|T059||CPT|ALT (SGPT) LEVEL
C0428324|T059||CPT|ALANINE TRANSAMINASE LEVEL
C0428324|T059||CPT|ALANINE TRANSAMINASE LEVEL 
C0428325|T059||CPT|ALT/SGPT SERUM LEVEL
C0428325|T059||CPT|ALT/SGPT SERUM LEVEL 
C0523461|T059||CPT|ALT MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE 
C0523461|T059||CPT|ALANINE AMINOTRANSFERASE (ALT) MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE
C0523461|T059||CPT|ALANINE AMINOTRANSFERASE MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE 
C0523461|T059||CPT|ALANINE AMINOTRANSFERASE (ALT) MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE 
C0523461|T059||CPT|ALANINE AMINOTRANSFERASE MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE
C0523461|T059||CPT|ALT MEASUREMENT, METHOD WITH PYRIDOXAL-5'-PHOSPHATE
C0523462|T059||CPT|ALT MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE 
C0523462|T059||CPT|ALANINE AMINOTRANSFERASE (ALT) MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE
C0523462|T059||CPT|ALANINE AMINOTRANSFERASE MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE 
C0523462|T059||CPT|ALANINE AMINOTRANSFERASE MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE
C0523462|T059||CPT|ALANINE AMINOTRANSFERASE (ALT) MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE 
C0523462|T059||CPT|ALT MEASUREMENT, METHOD WITHOUT PYRIDOXAL-5'-PHOSPHATE
C0428326|T059||CPT|SERUM GLUTAMIC OXALOACETIC TRANSAMINASE (SGPT) - BLOOD MEASUREMENT 
C0428326|T059||CPT|SERUM GLUTAMIC OXALOACETIC TRANSAMINASE (SGPT) - BLOOD MEASUREMENT
C0428326|T059||CPT|SGPT - BLOOD MEASUREMENT 
C0428326|T059||CPT|SGPT - BLOOD LEVEL
C0428326|T059||CPT|SGPT - BLOOD MEASUREMENT
C0428327|T059||CPT|ALT - BLOOD MEASUREMENT 
C0428327|T059||CPT|ALANINE AMINOTRANSFERASE (ALT) - BLOOD MEASUREMENT
C0428327|T059||CPT|LIVER ENZYMES (& BLOOD LEVEL [ALT] OR [SGPT])
C0428327|T059||CPT|LIVER ENZYMES (& BLOOD LEVEL [ALT] OR [SGPT]) 
C0428327|T059||CPT|SGPT - BLOOD LEVEL
C0428327|T059||CPT|ALT - BLOOD LEVEL
C0428327|T059||CPT|ALANINE AMINOTRANSFERASE - BLOOD MEASUREMENT
C0428327|T059||CPT|ALANINE AMINOTRANSFERASE (ALT) - BLOOD MEASUREMENT 
C0428327|T059||CPT|ALANINE AMINOTRANSFERASE - BLOOD MEASUREMENT 
C0428327|T059||CPT|ALT - BLOOD MEASUREMENT
C0428327|T059||CPT|ALT BLOOD MEASUREMENT
C0042040|T059||CPT|URINE BILIRUBIN TESTS
C0042040|T059||CPT|BILIRUBIN URINE
C0042040|T059||CPT|URINE BILIRUBIN TEST
C0042040|T059||CPT|BILIRUBIN MEASUREMENT, URINE
C0042040|T059||CPT|URINE BILIRUBIN
C0042040|T059||CPT|URINE BILIRUBIN LEVEL
C0042040|T059||CPT|BILIRUBIN MEASUREMENT, URINE 
C0702270|T059||CPT|AMNIOTIC FLUID BILIRUBIN TEST
C0702270|T059||CPT|BILIRUBIN MEASUREMENT, AMNIOTIC FLUID
C0702270|T059||CPT|BILIRUBIN MEASUREMENT, AMNIOTIC FLUID 
C1278039|T059||CPT|SERUM TOTAL BILIRUBIN
C1278039|T059||CPT|SERUM TOTAL BILIRUBIN MEASUREMENT
C1278039|T059||CPT|TOTAL SERUM BILIRUBIN LEVEL
C1278039|T059||CPT|SERUM TOTAL BILIRUBIN MEASUREMENT 
C1278039|T059||CPT|SERUM TOTAL BILIRUBIN LEVEL
C1278039|T059||CPT|SERUM TOTAL BILIRUBIN LEVEL 
C1278039|T059||CPT|SERUM BILIRUBIN TOTAL
C1278039|T059||CPT|SERUM TOTAL BILIRUBIN MEASUREMENT 
C2711150|T059||CPT|MEASUREMENT OF TOTAL BILIRUBIN IN CORD BLOOD SPECIMEN 
C2711150|T059||CPT|MEASUREMENT OF TOTAL BILIRUBIN IN CORD BLOOD SPECIMEN
C0201913|T059|1011294|CPT|BILIRUBIN; TOTAL|BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN MEASUREMENT|BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN TOTAL|BILIRUBIN
C0201913|T059|1011294|CPT|MEASUREMENT OF TOTAL BILIRUBIN|BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN|BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN (& LEVEL) |BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN, TOTAL MEASUREMENT|BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN, TOTAL MEASUREMENT |BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN (& LEVEL)|BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN|BILIRUBIN
C0201913|T059|1011294|CPT|BILI|BILIRUBIN
C0201913|T059|1011294|CPT|TOTAL BILIRUBIN LEVEL|BILIRUBIN
C0201913|T059|1011294|CPT|BILIRUBIN, TOTAL MEASUREMENT  [AMBIGUOUS]|BILIRUBIN
C0373554|T059|82252|CPT|BILIRUBIN; FECES, QUALITATIVE|FECAL BILIRUBIN TEST
C0373554|T059|82252|CPT|BILIRUBIN FECES QUALITATIVE|FECAL BILIRUBIN TEST
C0373554|T059|82252|CPT|FECAL BILIRUBIN TEST|FECAL BILIRUBIN TEST
C0697273|T059||CPT|BILIRUBIN; DIRECT
C0697273|T059||CPT|BILIRUBIN CONJUGATED
C0697273|T059||CPT|BILIRUBIN DIRECT
C0697273|T059||CPT|CONJUGATED BILIRUBIN TEST
C1278036|T059||CPT|PLASMA TOTAL BILIRUBIN LEVEL 
C1278036|T059||CPT|PLASMA TOTAL BILIRUBIN LEVEL
C1278036|T059||CPT|PLASMA BILIRUBIN TOTAL
C1278036|T059||CPT|PLASMA TOTAL BILIRUBIN TEST
C1278036|T059||CPT|PLASMA TOTAL BILIRUBIN MEASUREMENT 
C1278036|T059||CPT|PLASMA TOTAL BILIRUBIN MEASUREMENT
C0201917|T059||CPT|BABY BILIRUBIN MEASUREMENT
C0201917|T059||CPT|BILIRUBIN, NEONATAL MEASUREMENT
C0201917|T059||CPT|BILIRUBIN, NEONATAL MEASUREMENT 
C0201917|T059||CPT|TOTAL BILIRUBIN, NEONATAL MEASUREMENT
C0201917|T059||CPT|MICROBILIRUBIN MEASUREMENT
C0201917|T059||CPT|TOTAL BILIRUBIN, NEONATAL MEASUREMENT 
C0428441|T059||CPT|BILIRUBIN
C0428441|T059||CPT|SERUM BILIRUBIN MEASUREMENT 
C0428441|T059||CPT|SERUM BILIRUBIN (& LEVEL) 
C0428441|T059||CPT|BILIRUBIN - SERUM
C0428441|T059||CPT|SERUM BILIRUBIN NOS 
C0428441|T059||CPT|SERUM BILIRUBIN NOS
C0428441|T059||CPT|SERUM BILIRUBIN LEVEL
C0428441|T059||CPT|SERUM BILIRUBIN (& LEVEL)
C0428441|T059||CPT|SERUM BILIRUBIN
C0428441|T059||CPT|SB - SERUM BILIRUBIN
C0428441|T059||CPT|SERUM BILIRUBIN MEASUREMENT 
C0428441|T059||CPT|SERUM BILIRUBIN MEASUREMENT
C1278064|T059||CPT|SERUM METHAEMALBUMIN LEVEL 
C1278064|T059||CPT|SERUM METHAEMALBUMIN LEVEL
C1278064|T059||CPT|SERUM METHEMALBUMIN LEVEL
C1278064|T059||CPT|SERUM METHAEMALBUMIN MEASUREMENT
C1278064|T059||CPT|SERUM METHEMALBUMIN MEASUREMENT 
C1278064|T059||CPT|SERUM METHEMALBUMIN MEASUREMENT
C2711642|T059||CPT|MEASUREMENT OF ALBUMIN GRADIENT BETWEEN SERUM SPECIMEN AND ASCITIC FLUID SPECIMEN 
C2711642|T059||CPT|MEASUREMENT OF ALBUMIN GRADIENT BETWEEN SERUM SPECIMEN AND ASCITIC FLUID SPECIMEN
C2711642|T059||CPT|SERUM ASCITES ALBUMIN GRADIENT
C2097241|T059||CPT|SERUM ALBUMIN/GLOBULIN RATIO 
C2097241|T059||CPT|SERUM ALBUMIN/GLOBULIN RATIO
C2097241|T059||CPT|ALBUMIN/GLOBULIN RATIO
C2097242|T059||CPT|SERUM ALBUMIN-GLOBULIN CAPACITY 
C2097242|T059||CPT|SERUM ALBUMIN-GLOBULIN CAPACITY
C2097242|T059||CPT|ALBUMIN-GLOBULIN CAPACITY
C2732844|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN SERUM OR PLASMA SPECIMEN 120 MINUTES AFTER 75 GRAM ORAL GLUCOSE CHALLENGE 
C2732844|T059||CPT|QUANTITATIVE MEASUREMENT OF GLUCOSE IN SERUM OR PLASMA SPECIMEN 120 MINUTES AFTER 75 GRAM ORAL GLUCOSE CHALLENGE
C2732844|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN SERUM OR PLASMA SPECIMEN 120 MINUTES AFTER 75 GRAM ORAL GLUCOSE CHALLENGE
C2733143|T059||CPT|QUANTITATIVE MEASUREMENT OF SUBSTANCE RATE OF GLUCOSE EXCRETION IN URINE SPECIMEN
C2733143|T059||CPT|QUANTITATIVE MEASUREMENT OF SUBSTANCE RATE OF GLUCOSE EXCRETION IN URINE
C2733143|T059||CPT|QUANTITATIVE MEASUREMENT OF SUBSTANCE RATE OF GLUCOSE EXCRETION IN URINE SPECIMEN 
C2732700|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN PERICARDIAL FLUID SPECIMEN 
C2732700|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN PERICARDIAL FLUID SPECIMEN
C2732700|T059||CPT|QUANTITATIVE MEASUREMENT OF GLUCOSE IN PERICARDIAL FLUID SPECIMEN
C2732794|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN 1 HOUR POSTPRANDIAL URINE SPECIMEN 
C2732794|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN 1 HOUR POSTPRANDIAL URINE SPECIMEN
C2732794|T059||CPT|QUANTITATIVE MEASUREMENT OF GLUCOSE IN 1 HOUR POSTPRANDIAL URINE SPECIMEN
C2732897|T059||CPT|QUANTITATIVE MEASUREMENT OF GLUCOSE IN PERITONEAL DIALYSIS FLUID SPECIMEN
C2732897|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN PERITONEAL DIALYSIS FLUID SPECIMEN
C2732897|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN PERITONEAL DIALYSIS FLUID SPECIMEN 
C2732804|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN SYNOVIAL FLUID SPECIMEN
C2732804|T059||CPT|QUANTITATIVE MEASUREMENT OF GLUCOSE IN SYNOVIAL FLUID SPECIMEN
C2732804|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN SYNOVIAL FLUID SPECIMEN 
C2733070|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN SERUM OR PLASMA SPECIMEN 6 HOURS AFTER GLUCOSE CHALLENGE
C2733070|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN SERUM OR PLASMA SPECIMEN 6 HOURS AFTER GLUCOSE CHALLENGE 
C2733070|T059||CPT|QUANTITATIVE MEASUREMENT OF GLUCOSE IN SERUM OR PLASMA SPECIMEN 6 HOURS AFTER GLUCOSE CHALLENGE
C2732796|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS RATE OF EXCRETION OF GLUCOSE IN 24 HOUR URINE SPECIMEN
C2732796|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS RATE OF EXCRETION OF GLUCOSE IN 24 HOUR URINE SPECIMEN 
C2732796|T059||CPT|QUANTITATIVE MEASUREMENT OF GLUCOSE IN 24 HOUR URINE SPECIMEN
C2732716|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN POSTCALORIE FASTING SERUM OR PLASMA SPECIMEN
C2732716|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN POSTCALORIE FASTING SERUM OR PLASMA
C2732716|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN POSTCALORIE FASTING SERUM OR PLASMA SPECIMEN 
C2732249|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN PLEURAL FLUID SPECIMEN 
C2732249|T059||CPT|QUANTITATIVE MEASUREMENT OF MASS CONCENTRATION OF GLUCOSE IN PLEURAL FLUID SPECIMEN
C2732249|T059||CPT|QUANTITATIVE MEASUREMENT OF GLUCOSE IN PLEURAL FLUID SPECIMEN
C0201899|T059|80076|CPT|SERUM SGOT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SERUM AST|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPARTATE AMINOTRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
# C0201899|T059|80076|CPT|GOT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
# C0201899|T059|80076|CPT|AST|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPARTATE AMINOTRANSFERASE MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|TRANSFERASE; ASPARTATE AMINO (AST) (SGOT)|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|TRANSFERASE ASPARTATE AMINO AST SGOT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|LIVER ENZYME (SGOT), LEVEL|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE (AST) (SGOT)|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|AST - ASPARTATE TRANSAM SGOT (& LEVEL) |MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|AST - ASPARTATE TRANSAM SGOT (& LEVEL)|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|TRANSFERASE (AST) (SGOT)|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SGOT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPARTATE TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASP TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SERUM GLUTAMIC-OXALOACETIC TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|GLUTAMIC-OXALOACETIC TRANSFERASE|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SERUM ASPARTATE TRANSAMINASE TEST|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|AST MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|GLUTAMIC OXALOACETIC TRANSAMINASE MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|GOT MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|SGOT MEASUREMENT|MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C0201899|T059|80076|CPT|ASPARTATE AMINOTRANSFERASE MEASUREMENT |MEASUREMENT OF ASPARTATE AMINO TRANSFERASE
C1261155|T059||CPT|AST SERUM MEASUREMENT 
C1261155|T059||CPT|SERUM ASPARTATE TRANSAMINASE MEASUREMENT
C1261155|T059||CPT|SERUM ASPARTATE AMINOTRANSFERASE MEASUREMENT
C1261155|T059||CPT|SERUM SGOT MEASUREMENT
C1261155|T059||CPT|AST SERUM LEVEL
C1261155|T059||CPT|AST SERUM LEVEL 
C1261155|T059||CPT|ASPARTATE AMINOTRANSFERASE (AST) SERUM MEASUREMENT 
C1261155|T059||CPT|ASPARTATE AMINOTRANSFERASE SERUM MEASUREMENT 
C1261155|T059||CPT|ASPARTATE AMINOTRANSFERASE (AST) SERUM MEASUREMENT
C1261155|T059||CPT|ASPARTATE AMINOTRANSFERASE SERUM MEASUREMENT
C1261155|T059||CPT|AST SERUM MEASUREMENT
C0523517|T059||CPT|ASPARTATE AMINO TRANSFERASE/ALANINE AMINO TRANSFERASE RATIO MEASUREMENT
C0523517|T059||CPT|ASPARTATE AMINO TRANSFERASE/ALANINE AMINO TRANSFERASE RATIO MEASUREMENT 
C1278050|T059||CPT|PLASMA ASPARTATE TRANSAMINASE LEVEL 
C1278050|T059||CPT|PLASMA ASPARTATE TRANSAMINASE LEVEL
C1278050|T059||CPT|PLASMA ASPARTATE TRANSAMINASE MEASUREMENT 
C1278050|T059||CPT|PLASMA ASPARTATE TRANSAMINASE MEASUREMENT
C0523891|T059|84295|CPT|SERUM SODIUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM NA+|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM MEASUREMENT|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM MEASUREMENT |SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM; SERUM, PLASMA OR WHOLE BLOOD|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM SERUM PLASMA OR WHOLE BLOOD|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|MEASUREMENT OF SODIUM IN SERUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM (& LEVEL) |SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM (& LEVEL)|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM - SERUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM ION TEST|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM MEASUREMENT, SERUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM LEVEL|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SODIUM MEASUREMENT, SERUM |SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|ASSAY OF SERUM SODIUM|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM EACH TEST|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C0523891|T059|84295|CPT|SERUM SODIUM EA.TST|SODIUM; SERUM, PLASMA OR WHOLE BLOOD
C2016757|T059||CPT|SODIUM MEASUREMENT FROM OTHER SOURCE 
C2016757|T059||CPT|SODIUM MEASUREMENT FROM OTHER SOURCE
C2016757|T059||CPT|SODIUM LEVEL FROM SOURCE OTHER THAN URINE
C2702997|T059|84295|CPT|WHOLE BLOOD SODIUM MEASUREMENT |MEASUREMENT OF SODIUM IN WHOLE BLOOD
C2702997|T059|84295|CPT|WHOLE BLOOD SODIUM MEASUREMENT|MEASUREMENT OF SODIUM IN WHOLE BLOOD
C2702997|T059|84295|CPT|MEASUREMENT OF SODIUM IN WHOLE BLOOD|MEASUREMENT OF SODIUM IN WHOLE BLOOD
C3161784|T059||CPT|SERUM SODIUM AFTER FLUDROCORTISONE
C3161784|T059||CPT|SERUM SODIUM AFTER FLUDROCORTISONE 
C3161785|T059||CPT|SERUM SODIUM AFTER DEMECLOCYLINE
C3161785|T059||CPT|SERUM SODIUM AFTER DEMECLOCYLINE 
C0302353|T059|84132|CPT|SERUM K+|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM MEASUREMENT|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM MEASUREMENT |POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|POTASSIUM LEVEL|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|POTASSIUM SERUM PLASMA/WHOLE BLOOD|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|POTASSIUM; SERUM, PLASMA OR WHOLE BLOOD|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|MEASUREMENT OF POTASSIUM IN SERUM|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|POTASSIUM - SERUM|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM (& LEVEL) |POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM (& LEVEL)|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM LEVEL|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|SERUM POTASSIUM MEASUREMENT |POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|T059|84132|CPT|ASSAY OF SERUM POTASSIUM|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0553704|T059||CPT|POTASSIUM, INCREASED LEVEL
C0553704|T059||CPT|SERUM POTASIUM INCREASED
C0553704|T059||CPT|SERUM POTASSIUM INCREASED
C0553704|T059||CPT|POTASSIUM SERUM INCREASED
C2229880|T059||CPT|SERUM TOTAL BODY POTASSIUM MEASUREMENT
C2229880|T059||CPT|SERUM TOTAL BODY POTASSIUM MEASUREMENT 
C2229880|T059||CPT|TOTAL BODY POTASSIUM LEVEL
C0373708|T059|84155|CPT|PROTEIN, TOTAL, EXCEPT BY REFRACTOMETRY; SERUM, PLASMA OR WHOLE BLOOD|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD
C0373708|T059|84155|CPT|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD
C0373708|T059|84155|CPT|ASSAY OF PROTEIN SERUM|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD
C4048459|T059|80055|CPT|OBSTETRIC PANEL|OBSTETRIC PANEL
C4048459|T059|80055|CPT|OBSTETRIC PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: BLOOD COUNT, COMPLETE (CBC), AUTOMATED AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) HEPATITIS B SURFACE ANTIGEN (HBSAG) (87340) ANTIBODY, RUBELLA (86762) SYPHILIS TEST, NON-TREPONEMAL ANTIBODY; QUALITATIVE (EG, VDRL, RPR, ART) (86592) ANTIBODY SCREEN, RBC, EACH SERUM TECHNIQUE (86850) BLOOD TYPING, ABO (86900) AND BLOOD TYPING, RH (D) (86901)|OBSTETRIC PANEL
C0812553|T059|80074|CPT|ACUTE HEPATITIS PANEL|ACUTE HEPATITIS PANEL
C0812553|T059|80074|CPT|ACUTE HEPATITIS PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: HEPATITIS A ANTIBODY (HAAB), IGM ANTIBODY (86709) HEPATITIS B CORE ANTIBODY (HBCAB), IGM ANTIBODY (86705) HEPATITIS B SURFACE ANTIGEN (HBSAG) (87340) HEPATITIS C ANTIBODY (86803)|ACUTE HEPATITIS PANEL
C1964052|T059|80047|CPT|BASIC METABOLIC PANEL CALCIUM IONIZED|METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|METABOLIC PANEL IONIZED CA|METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|BMP WITH IONIZED CALCIUM|METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|BASIC METABOLIC PANEL WITH IONIZED CALCIUM |METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|BASIC METABOLIC PANEL WITH IONIZED CALCIUM|METABOLIC PANEL IONIZED CA
C1964052|T059|80047|CPT|BASIC METABOLIC PANEL (CALCIUM, IONIZED) THIS PANEL MUST INCLUDE THE FOLLOWING: CALCIUM, IONIZED (82330) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) POTASSIUM (84132) SODIUM (84295) UREA NITROGEN (BUN) (84520)|METABOLIC PANEL IONIZED CA
C3836932|T059||CPT|LIPIDS TEST PANEL SERUM OR PLASMA
C3836932|T059||CPT|LIPIDS TEST PANEL SERUM OR PLASMA 
C0430044|T059||CPT|FASTING LIPID PANEL 
C0430044|T059||CPT|FASTING LIPID PANEL
C0430044|T059||CPT|LIPIDS TEST PANEL FASTING
C0430044|T059||CPT|FASTING LIPID PROFILE
C0430044|T059||CPT|FLP - FASTING LIPID PROFILE
C0430044|T059||CPT|FASTING LIPID PROFILE 
C0523942|T059||CPT|TRIGLYCERIDE AND ESTER IN HDL MEASUREMENT 
C0523942|T059||CPT|TRIGLYCERIDE AND ESTER IN HIGH DENSITY LIPOPROTEIN MEASUREMENT 
C0523942|T059||CPT|TRIGLYCERIDE AND ESTER IN HIGH DENSITY LIPOPROTEIN MEASUREMENT
C0523942|T059||CPT|TRIGLYCERIDE AND ESTER IN HDL MEASUREMENT
C0523943|T059||CPT|TRIGLYCERIDE AND ESTER IN INTERMEDIATE DENSITY LIPOPROTEIN MEASUREMENT 
C0523943|T059||CPT|TRIGLYCERIDE AND ESTER IN IDL MEASUREMENT 
C0523943|T059||CPT|TRIGLYCERIDE AND ESTER IN INTERMEDIATE DENSITY LIPOPROTEIN MEASUREMENT
C0523943|T059||CPT|TRIGLYCERIDE AND ESTER IN IDL MEASUREMENT
C0523944|T059||CPT|TRIGLYCERIDE AND ESTER IN LOW DENSITY LIPOPROTEIN MEASUREMENT
C0523944|T059||CPT|TRIGLYCERIDE AND ESTER IN LDL MEASUREMENT 
C0523944|T059||CPT|TRIGLYCERIDE AND ESTER IN LOW DENSITY LIPOPROTEIN MEASUREMENT 
C0523944|T059||CPT|TRIGLYCERIDE AND ESTER IN LDL MEASUREMENT
C0523945|T059||CPT|TRIGLYCERIDE AND ESTER IN VLDL MEASUREMENT 
C0523945|T059||CPT|TRIGLYCERIDE AND ESTER IN VERY LOW DENSITY LIPOPROTEIN MEASUREMENT
C0523945|T059||CPT|TRIGLYCERIDE AND ESTER IN VERY LOW DENSITY LIPOPROTEIN MEASUREMENT 
C0523945|T059||CPT|TRIGLYCERIDE AND ESTER IN VLDL MEASUREMENT
C0519823|T059|80048|CPT|METABOLIC PANEL TOTAL CA|BASIC METABOLIC PANEL CALCIUM TOTAL
C0519823|T059|80048|CPT|BASIC METABOLIC PANEL CALCIUM TOTAL|BASIC METABOLIC PANEL CALCIUM TOTAL
C0519823|T059|80048|CPT|BASIC METABOLIC PANEL (CALCIUM, TOTAL) THIS PANEL MUST INCLUDE THE FOLLOWING: CALCIUM, TOTAL (82310) CARBON DIOXIDE (BICARBONATE) (82374) CHLORIDE (82435) CREATININE (82565) GLUCOSE (82947) POTASSIUM (84132) SODIUM (84295) UREA NITROGEN (BUN) (84520)|BASIC METABOLIC PANEL CALCIUM TOTAL
C0812554|T059|80076|CPT|HEPATIC FUNCTION PANEL|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)
C0812554|T059|80076|CPT|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)
C0812554|T059|80076|CPT|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT)|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)
C0812554|T059|80076|CPT|LIVER FUNCTION BLOOD TEST PANEL|HEPATIC FUNCTION PANEL THIS PANEL MUST INCLUDE THE FOLLOWING: ALBUMIN (82040) BILIRUBIN, TOTAL (82247) BILIRUBIN, DIRECT (82248) PHOSPHATASE, ALKALINE (84075) PROTEIN, TOTAL (84155) TRANSFERASE, ALANINE AMINO (ALT) (SGPT) (84460) TRANSFERASE, ASPARTATE AMINO (AST) (SGOT) (84450)
C4050228|T059|80081|CPT|OBSTETRIC PANEL|OBSTETRIC PANEL
C4050228|T059|80081|CPT|OBSTETRIC PANEL (INCLUDES HIV TESTING) THIS PANEL MUST INCLUDE THE FOLLOWING: BLOOD COUNT, COMPLETE (CBC), AND AUTOMATED DIFFERENTIAL WBC COUNT (85025 OR 85027 AND 85004) OR BLOOD COUNT, COMPLETE (CBC), AUTOMATED (85027) AND APPROPRIATE MANUAL DIFFERENTIAL WBC COUNT (85007 OR 85009) HEPATITIS B SURFACE ANTIGEN (HBSAG) (87340) HIV-1 ANTIGEN(S), WITH HIV-1 AND HIV-2 ANTIBODIES, SINGLE RESULT (87389) ANTIBODY, RUBELLA (86762) SYPHILIS TEST, NON-TREPONEMAL ANTIBODY; QUALITATIVE (EG, VDRL, RPR, ART) (86592) ANTIBODY SCREEN, RBC, EACH SERUM TECHNIQUE (86850) BLOOD TYPING, ABO (86900) AND BLOOD TYPING, RH (D) (86901)|OBSTETRIC PANEL
C0430174|T059||CPT|METABOLIC FUNCTION TESTED
C0430174|T059||CPT|METABOLIC FUNCTION TEST NOS 
C0430174|T059||CPT|METABOLIC FUNCTION TEST NOS
C0430174|T059||CPT|METABOLIC FUNCTION TESTED 
C0430174|T059||CPT|METABOLIC FUNCTION TEST
C0430174|T059||CPT|METABOLIC FUNCTION TEST 
C0430174|T059||CPT|METABOLIC FUNCTION TESTED 
C2368348|T059||CPT|BASIC METABOLIC PANEL AND RENAL FUNCTION TESTS 
C2368348|T059||CPT|BASIC METABOLIC PANEL AND RENAL FUNCTION TESTS
C0430175|T059||CPT|CHEM. METAB. FUNCTION TEST NOS
C0430175|T059||CPT|CHEM. METAB. FUNCTION TEST NOS 
C0006779|T059||CPT|CALORIMETRY
C0006779|T059||CPT|CALORIMETRY 
C0204047|T059||CPT|ISCHAEMIC FOREARM EXERCISE TEST
C0204047|T059||CPT|ISCHAEMIC FOREARM EXERCISE TEST 
C0204047|T059||CPT|ISCHEMIC FOREARM EXERCISE TEST
C0204047|T059||CPT|ISCHAEMIC FOREARM EXERCISE TEST [AMBIGUOUS]
C0204047|T059||CPT|ISCHEMIC FOREARM EXERCISE TEST 
C0204047|T059||CPT|ISCHEMIC FOREARM EXERCISE TEST (REGIME/THERAPY)
C0204048|T059||CPT|ISCHEMIC LIMB EXERCISE WITH ELECTROMYOGRAPHY AND LACTIC ACID DETERMINATION 
C0204048|T059||CPT|ISCHEMIC LIMB EXERCISE WITH ELECTROMYOGRAPHY AND LACTIC ACID DETERMINATION
C0204048|T059||CPT|ISCHEMIC LIMB EXERCISE WITH EMG AND LACTIC ACID DETERMINATION
C0204048|T059||CPT|ISCHAEMIC LIMB EXERCISE WITH EMG AND LACTIC ACID DETERMINATION
C0204048|T059||CPT|ISCHEMIC LIMB EXERCISE WITH EMG AND LACTIC ACID DETERMINATION 
C0204048|T059||CPT|ISCHEMIC LIMB EXERCISE WITH EMG AND LACTIC ACID DETERMINATION (REGIME/THERAPY)
C1283822|T059||CPT|ISCHAEMIC LACTATE TEST
C1283822|T059||CPT|ISCHEMIC LACTATE TEST
C1283822|T059||CPT|ISCHEMIC LACTATE TEST 
C0430180|T059||CPT|BODY WATER TEST
C0430180|T059||CPT|BODY WATER TEST 
C0430177|T059||CPT|FLUSH PROVOCATION TEST
C0430177|T059||CPT|FLUSH PROVOCATION TEST 
C0430603|T059||CPT|METABOLIC FUNCTION NOT TESTED 
C0430603|T059||CPT|METABOLIC FUNCTION NOT TESTED 
C0430603|T059||CPT|METABOLIC FUNCTION NOT TESTED
C0430178|T059||CPT|NICOTINIC ACID LOADING TEST
C0430178|T059||CPT|NICOTINIC ACID LOADING TEST 
C0430176|T059||CPT|NITROGEN BALANCE TEST
C0430176|T059||CPT|NITROGEN BALANCE TEST 
C1273413|T059||CPT|ENDOCRINE STUDIES
C1273413|T059||CPT|ENDOCRINE STUDIES 
