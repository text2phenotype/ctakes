C0427512|T034|365630000|SNOMEDCT_US|FINDING OF WHITE BLOOD CELL NUMBER|WHITE BLOOD CELL NUMBER - FINDING
C0023516|T034|272170001|SNOMEDCT_US|LEUKOCYTES|WHITE BLOOD CELL (CELL)
C0023508|T034|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT PROCEDURE|WHITE BLOOD CELL COUNT - OBSERVATION
C0427512|T034|365630000|SNOMEDCT_US|WHITE BLOOD CELL COUNT LABORATORY RESULT|WHITE BLOOD CELL NUMBER - FINDING
C1271681|T034|391558003|SNOMEDCT_US|TOTAL WHITE BLOOD COUNT|TOTAL WHITE BLOOD CELL COUNT (PROCEDURE)
C1820736|T034||SNOMEDCT_US|ABSOLUTE WHITE BLOOD COUNT
C1821144|T034||SNOMEDCT_US|WHITE BLOOD COUNT
C4055603|T034||SNOMEDCT_US|APACHE II - WHITE BLOOD COUNT
C0162401|T034|142925001|SNOMEDCT_US|DIFFERENTIAL WHITE BLOOD CELL COUNT PROCEDURE|DIFF. WHITE CELL COUNT NOS (PROCEDURE)
C0427547|T034|165510005|SNOMEDCT_US|TOTAL WHITE CELL COUNT MEASUREMENT|TOTAL WHITE CELL COUNT NOS (PROCEDURE)
C1318024|T034||SNOMEDCT_US|TOTAL WHITE CELL COUNT RESULT
C2186576|T034||SNOMEDCT_US|REPORTED WHITE BLOOD CELL COUNT
C3495375|T034||SNOMEDCT_US|BLOOD COUNT; LEUKOCYTE (WBC), AUTOMATED
C3525788|T034||SNOMEDCT_US|MANUAL WHITE BLOOD CELL (WBC) COUNT
C0023516|T034|272170001|SNOMEDCT_US|LEUKOCYTE|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WBC|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|LEUKOCYTES|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|BLOOD CELL, WHITE|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WHITE BLOOD CELL|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|CORPUSCLE, WHITE BLOOD|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|BLOOD CORPUSCLE, WHITE|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|CORPUSCLES, WHITE BLOOD|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WHITE BLOOD CORPUSCLE|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WBC (WHITE BLOOD CELL)|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WHITE BLOOD CELL (CELL)|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|LEUCOCYTES|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WHITE BLOOD CELLS|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WHITE BLOOD CORPUSCLES|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|BLOOD CORPUSCLES, WHITE|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|BLOOD CELLS, WHITE|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|LEUCOCYTE|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WBC - WHITE BLOOD CELL|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|LEUKOCYTE (CELL)|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|LEUKOCYTE, NOS|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WHITE BLOOD CELL, NOS|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|RETICULOENDOTHELIAL SYSTEM, LEUKOCYTES|WHITE BLOOD CELL (CELL)
C0023516|T034|272170001|SNOMEDCT_US|WHITE CELL|WHITE BLOOD CELL (CELL)
C2358187|T034||SNOMEDCT_US|LEUKOCYTES &#X7C; BLOOD PRODUCT UNIT &#X7C; BLD-SER-PLAS
C1991552|T034||SNOMEDCT_US|LEUKOCYTES &#X7C; BLD-SER-PLAS
C0803389|T034||SNOMEDCT_US|LEUKOCYTES:NCNC:PT:XXX:QN:AUTOMATED COUNT
C0803389|T034||SNOMEDCT_US|LEUKOCYTES [#/VOLUME] IN UNSPECIFIED SPECIMEN BY AUTOMATED COUNT
C0803389|T034||SNOMEDCT_US|WBC # XXX AUTO
C0803389|T034||SNOMEDCT_US|LEUKOCYTES:NUMBER CONCENTRATION (COUNT/VOL):POINT IN TIME:TO BE SPECIFIED IN ANOTHER PART OF THE MESSAGE:QUANTITATIVE:AUTOMATED COUNT
C1254480|T034||SNOMEDCT_US|WHOLE BLOOD TOTAL LEUKOCYTE COUNT
C0023508|T034|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|COUNT, LEUKOCYTE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|COUNTS, LEUKOCYTE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|LEUKOCYTE COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|LEUKOCYTE COUNTS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|LEUKOCYTE NUMBERS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|NUMBER, LEUKOCYTE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|NUMBERS, LEUKOCYTE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT PROCEDURE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|LEUKOCYTE COUNT |WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WBC COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT |WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|LEUKOCYTES|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WHITE BLOOD CELLS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WBC|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WHITE CELLS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|LEUKOCYTE COUNT NOS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT NOS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WHITE BLOOD CELL ANALYSIS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|LEUCOCYTE COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|LEUKOCYTE NUMBER|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|BLOOD CELL COUNT, WHITE|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WHOLE BLOOD LEUKOCYTE COUNTS|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WBC - WHITE BLOOD CELL COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WCC - WHITE BLOOD CELL COUNT|WHITE BLOOD CELL COUNT - OBSERVATION
C0023508|T034|767002|SNOMEDCT_US|WHITE BLOOD CELL COUNT - OBSERVATION|WHITE BLOOD CELL COUNT - OBSERVATION
C3495375|T034||SNOMEDCT_US|BLOOD COUNT LEUKOCYTE WBC AUTOMATED
C3495375|T034||SNOMEDCT_US|AUTOMATED WHITE BLOOD CELL COUNT
C3495375|T034||SNOMEDCT_US|AUTOMATED WHITE BLOOD CELL (WBC) COUNT
C3495375|T034||SNOMEDCT_US|BLOOD COUNT; LEUKOCYTE (WBC), AUTOMATED
C3495375|T034||SNOMEDCT_US|AUTOMATED LEUKOCYTE COUNT
C0427547|T034|165510005|SNOMEDCT_US|TOTAL WHITE CELL COUNT NOS|TOTAL WHITE CELL COUNT NOS (PROCEDURE)
C0427547|T034|165510005|SNOMEDCT_US|TOTAL WHITE CELL COUNT NOS |TOTAL WHITE CELL COUNT NOS (PROCEDURE)
C0427547|T034|165510005|SNOMEDCT_US|TOTAL WHITE CELL COUNT MEASUREMENT|TOTAL WHITE CELL COUNT NOS (PROCEDURE)
C1271682|T034|390136004|SNOMEDCT_US|TOTAL WBC (IMM) |TOTAL WBC (IMM) (PROCEDURE)
C1271682|T034|390136004|SNOMEDCT_US|TOTAL WBC (IMM)|TOTAL WBC (IMM) (PROCEDURE)
C1271681|T034|391558003|SNOMEDCT_US|TOTAL WHITE BLOOD CELL COUNT |TOTAL WHITE BLOOD CELL COUNT (PROCEDURE)
C1271681|T034|391558003|SNOMEDCT_US|TOTAL WHITE BLOOD COUNT |TOTAL WHITE BLOOD CELL COUNT (PROCEDURE)
C1271681|T034|391558003|SNOMEDCT_US|TOTAL WHITE BLOOD CELL COUNT|TOTAL WHITE BLOOD CELL COUNT (PROCEDURE)
C1271681|T034|391558003|SNOMEDCT_US|TOTAL WHITE BLOOD COUNT|TOTAL WHITE BLOOD CELL COUNT (PROCEDURE)
