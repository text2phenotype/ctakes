C0010054|T047|443502000|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISEASE|DISORDER OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ARTERIOSCLEROSES, CORONARY|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ARTERIOSCLEROSES|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ATHEROSCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ATHEROSCLEROTIC HEART DISEASE|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS |ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ASHD - ATHEROSCLEROTIC HEART DISEASE|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY |ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CARDIAC SCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY (ARTERY) ATHEROSCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY (ARTERY) SCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|DISEASE;ATHEROSCLEROTIC;HEART|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ATHEROSCLEROTIC HEART DISEASE NOS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ATHEROSCLEROSIS, CORONARY|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ARTERIOSCLEROSIS, CORONARY|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY |ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ATHEROSCLEROSIS CORONARY ARTERY|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ATHEROSCLEROSIS |ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY SCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ARTERIOSCLEROTIC HEART DISEASE|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ASHD|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ARTHEROSCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ARTERY SCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ARTERY ATHEROSCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ARTERIOSCLEROSIS CORONARY ARTERY|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CARDIAC; SCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY; ARTERIOSCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY; SCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|DISEASE (OR DISORDER); ARTERIOSCLEROTIC, CORONARY (ARTERY)|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|DISEASE (OR DISORDER); ARTERIOSCLEROTIC, HEART|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|HEART; ARTERIOSCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|SCLEROSIS; CARDIAC|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|SCLEROSIS; CORONARY|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ARTERIOSCLEROSIS; CORONARY (ARTERY)|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ARTERIOSCLEROSIS; CORONARY|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ARTERIOSCLEROSIS; HEART|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|ATHEROSCLEROSES, CORONARY|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ATHEROSCLEROSES|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS |ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0010054|T047|443502000|SNOMEDCT_US|CORONARY ARTERY ARTERIOSCLEROSIS|ATHEROSCLEROSIS OF CORONARY ARTERY (DISORDER)
C0002963|T047|87343002|SNOMEDCT_US|THIS IS VASOSPASM NOT BLOCKED ARTERIES - WILL INCLUDE FOR NOW, SINCE WE ARE GOING FOR INCLUSIVITY, BUT DOCTORS WILL MOSTLY CONSIDER THIS A FALSE POSITIVE FOR CAD|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|ANGINA PECTORIS, VARIANT|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|PRINZMETALS ANGINA|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|VARIANT ANGINA PECTORIS|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|ANGINA, PRINZMETAL'S|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|PRINZMETAL'S ANGINA|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|VARIANT ANGINA|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|PRINZMENTAL ANGINA|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|PRINZMETAL'S ANGINA |PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|ANGINA PECTORIS, VARIANT [DISEASE/FINDING]|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|ANGINA, PRINZMETAL|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|VASOSPASTIC ANGINA|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|CORONARY ARTERY SPASM ANGINA|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|PRINZMETAL ANGINA |PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|PRINZMETAL; ANGINA|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|ANGINA PECTORIS; VARIANT|PRINZMENTAL ANGINA
C0002963|T047|87343002|SNOMEDCT_US|VARIANT; ANGINA|PRINZMENTAL ANGINA
C0596384|T047||SNOMEDCT_US|CORONARY FIBROSIS
C0178570|T047||SNOMEDCT_US|CORONARY OCCLUSION/THROMBOSIS
C0542269|T047|314207007|SNOMEDCT_US|NON-Q WAVE MYOCARDIAL INFARCTION NOS|NON-Q WAVE MYOCARDIAL INFARCTION (DISORDER)
C0542269|T047|314207007|SNOMEDCT_US|NON-Q WAVE MYOCARDIAL INFARCTION|NON-Q WAVE MYOCARDIAL INFARCTION (DISORDER)
C0542269|T047|314207007|SNOMEDCT_US|ACUTE NON-Q-WAVE MYOCARDIAL INFARCTION|NON-Q WAVE MYOCARDIAL INFARCTION (DISORDER)
C0542269|T047|314207007|SNOMEDCT_US|ACUTE NON-Q-WAVE MYOCARDIAL INFARCTION |NON-Q WAVE MYOCARDIAL INFARCTION (DISORDER)
C0542269|T047|314207007|SNOMEDCT_US|SUBENDOCARDIAL NON-Q-WAVE MYOCARDIAL INFARCTION ACUTE|NON-Q WAVE MYOCARDIAL INFARCTION (DISORDER)
C0542269|T047|314207007|SNOMEDCT_US|NON-Q WAVE MYOCARDIAL INFARCTION |NON-Q WAVE MYOCARDIAL INFARCTION (DISORDER)
C0542060|T047||SNOMEDCT_US|ISCHEMIA CORONARY ARTERY ORIGIN
C0542060|T047||SNOMEDCT_US|ISCHAEMIA CORONARY ARTERY ORIGIN
C0542060|T047||SNOMEDCT_US|ISCHEMIA; CORONARY
C0856737|T047||SNOMEDCT_US|SINGLE VESSEL DISEASE
C0856738|T047||SNOMEDCT_US|TRIPLE VESSEL DISEASE
C0856739|T047||SNOMEDCT_US|LEFT MAIN STEM DISEASE
C0856740|T047||SNOMEDCT_US|MAIN STEM DISEASE
C0857530|T047||SNOMEDCT_US|RIGHT MAIN STEM DISEASE
C0375265|T047||SNOMEDCT_US|COR ATH BYPASS GRAFT NOS
C0375265|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF UNSPECIFIED BYPASS GRAFT
C0375265|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF BYPASS GRAFT
C0375265|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF BYPASS GRAFT
C0375265|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF BYPASS GRAFT NOS
C0340285|T047|233817007|SNOMEDCT_US|3-VESSEL CORONARY ARTERY STENOSIS |TRIPLE VESSEL DISEASE OF THE HEART (DISORDER)
C0340285|T047|233817007|SNOMEDCT_US|3-VESSEL CORONARY ARTERY STENOSIS|TRIPLE VESSEL DISEASE OF THE HEART (DISORDER)
C0340285|T047|233817007|SNOMEDCT_US|TRIPLE VESSEL CORONARY ARTERY DISEASE |TRIPLE VESSEL DISEASE OF THE HEART (DISORDER)
C0340285|T047|233817007|SNOMEDCT_US|TRIPLE VESSEL CORONARY ARTERY DISEASE|TRIPLE VESSEL DISEASE OF THE HEART (DISORDER)
C0340285|T047|233817007|SNOMEDCT_US|TRIPLE VESSEL DISEASE OF THE HEART|TRIPLE VESSEL DISEASE OF THE HEART (DISORDER)
C0340285|T047|233817007|SNOMEDCT_US|ARTERIOSCLEROSIS CORONARY ARTERY TRIPLE VESSEL DISEASE|TRIPLE VESSEL DISEASE OF THE HEART (DISORDER)
C0340285|T047|233817007|SNOMEDCT_US|TRIPLE VESSEL DISEASE OF HEART|TRIPLE VESSEL DISEASE OF THE HEART (DISORDER)
C0340285|T047|233817007|SNOMEDCT_US|TRIPLE VESSEL DISEASE OF HEART |TRIPLE VESSEL DISEASE OF THE HEART (DISORDER)
C0340285|T047|233817007|SNOMEDCT_US|TRIPLE VESSEL DISEASE OF THE HEART |TRIPLE VESSEL DISEASE OF THE HEART (DISORDER)
C2366973|T047||SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS DUE TO LIPID-RICH PLAQUE
C2366973|T047||SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS DUE TO LIPID-RICH PLAQUE 
C2062869|T047||SNOMEDCT_US|ASYMPTOMATIC CORONARY ARTERIOSCLEROSIS 
C2062869|T047||SNOMEDCT_US|ASYMPTOMATIC CORONARY ARTERIOSCLEROSIS
C0685094|T047|92517006|SNOMEDCT_US|CALCIFIC CORONARY ARTERIOSCLEROSIS|CALCIFIC CORONARY ARTERIOSCLEROSIS (DISORDER)
C0685094|T047|92517006|SNOMEDCT_US|CALCIFIC CORONARY ARTERIOSCLEROSIS |CALCIFIC CORONARY ARTERIOSCLEROSIS (DISORDER)
C0685094|T047|92517006|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS DUE TO CALCIFIED CORONARY LESION|CALCIFIC CORONARY ARTERIOSCLEROSIS (DISORDER)
C0685094|T047|92517006|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS DUE TO CALCIFIED CORONARY LESION |CALCIFIC CORONARY ARTERIOSCLEROSIS (DISORDER)
C0685094|T047|92517006|SNOMEDCT_US|CALCIFIC CORONARY ARTERIOSCLEROSIS |CALCIFIC CORONARY ARTERIOSCLEROSIS (DISORDER)
C2321373|T047||SNOMEDCT_US|PROGRESSIVE CORONARY ARTERY DISEASE
C2321373|T047||SNOMEDCT_US|PROGRESSIVE CORONARY ARTERY DISEASE 
C2321817|T047||SNOMEDCT_US|SAMPLE TEMPLATE CORONARY ARTERY DISEASE
C2321817|T047||SNOMEDCT_US|SAMPLE TEMPLATE CORONARY ARTERY DISEASE 
C1997154|T047|427919004|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS DUE TO RADIATION|CORONARY ARTERIOSCLEROSIS DUE TO RADIATION (DISORDER)
C1997154|T047|427919004|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS DUE TO RADIATION |CORONARY ARTERIOSCLEROSIS DUE TO RADIATION (DISORDER)
C1997154|T047|427919004|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS CAUSED BY RADIATION|CORONARY ARTERIOSCLEROSIS DUE TO RADIATION (DISORDER)
C1997154|T047|427919004|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS CAUSED BY RADIATION |CORONARY ARTERIOSCLEROSIS DUE TO RADIATION (DISORDER)
C1997154|T047|427919004|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS DUE TO RADIATION |CORONARY ARTERIOSCLEROSIS DUE TO RADIATION (DISORDER)
C3472163|T047|1641000119107|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS IN NATIVE ARTERY |CORONARY ARTERIOSCLEROSIS IN NATIVE ARTERY (DISORDER)
C3472163|T047|1641000119107|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS IN NATIVE ARTERY|CORONARY ARTERIOSCLEROSIS IN NATIVE ARTERY (DISORDER)
C3472163|T047|1641000119107|SNOMEDCT_US|ARTERIOSCLEROSIS CORONARY IN NATIVE ARTERY|CORONARY ARTERIOSCLEROSIS IN NATIVE ARTERY (DISORDER)
C3472163|T047|1641000119107|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS IN NATIVE ARTERY |CORONARY ARTERIOSCLEROSIS IN NATIVE ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CAD|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISEASE|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|ARTERY DISEASES, CORONARY|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISEASES|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISEASE, CORONARY ARTERY|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|ARTERY DISEASE, CORONARY|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISEASES, CORONARY ARTERY|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DIS|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CAD (CORONARY ARTERY DISEASE)|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISORDER OF CORONARY ARTERIES |DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISEASE |DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISORDER OF CORONARY ARTERIES|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISORDERS|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY DISEASE|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISEASE [DISEASE/FINDING]|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISEASE |DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISEASE OF THE CORONARY ARTERIES|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CAD - CORONARY ARTERY DISEASE|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY HEART DISEASE|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISORDER|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISEASE CORONARY ARTERY|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISORDER CORONARY ARTERY|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISORDER (NOS)|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISEASE NOS|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CARDIO/PULM: CORONARY ARTERY DISEASE|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY (ARTERY); DISEASE|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISEASE (OR DISORDER); ARTERY, CORONARY|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISEASE (OR DISORDER); CORONARY (ARTERY)|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISEASE (OR DISORDER); HEART, ARTERY, ARTERIAL|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|ARTERY; DISORDER, CORONARY|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|CORONARY ARTERY DISEASE, NOS|DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISORDER OF CORONARY ARTERY |DISORDER OF CORONARY ARTERY (DISORDER)
C1956346|T047|414024009|SNOMEDCT_US|DISORDER OF CORONARY ARTERY|DISORDER OF CORONARY ARTERY (DISORDER)
C0948089|T047|394659003|SNOMEDCT_US|ACUTE CORONARY SYNDROME|ACS - ACUTE CORONARY SYNDROME
C0948089|T047|394659003|SNOMEDCT_US|CORONARY SYNDROMES, ACUTE|ACS - ACUTE CORONARY SYNDROME
C0948089|T047|394659003|SNOMEDCT_US|SYNDROMES, ACUTE CORONARY|ACS - ACUTE CORONARY SYNDROME
C0948089|T047|394659003|SNOMEDCT_US|ACUTE CORONARY SYNDROMES|ACS - ACUTE CORONARY SYNDROME
C0948089|T047|394659003|SNOMEDCT_US|SYNDROME, ACUTE CORONARY|ACS - ACUTE CORONARY SYNDROME
C0948089|T047|394659003|SNOMEDCT_US|CORONARY SYNDROME, ACUTE|ACS - ACUTE CORONARY SYNDROME
C0948089|T047|394659003|SNOMEDCT_US|ACUTE CORONARY SYNDROME [DISEASE/FINDING]|ACS - ACUTE CORONARY SYNDROME
C0948089|T047|394659003|SNOMEDCT_US|ACUTE CORONARY SYNDROME |ACS - ACUTE CORONARY SYNDROME
C0948089|T047|394659003|SNOMEDCT_US|ACUTE CORONARY SYNDROME |ACS - ACUTE CORONARY SYNDROME
C0948089|T047|394659003|SNOMEDCT_US|ACS - ACUTE CORONARY SYNDROME|ACS - ACUTE CORONARY SYNDROME
C0340325|T047|194821006|SNOMEDCT_US|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0340325|T047|194821006|SNOMEDCT_US|ABORTED MYOCARDIAL INFARCTION|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0340325|T047|194821006|SNOMEDCT_US|MI - MYOCARDIAL INFARCTION ABORTED|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0340325|T047|194821006|SNOMEDCT_US|ABORTED MYOCARDIAL INFARCTION |CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0340325|T047|194821006|SNOMEDCT_US|CORONARY THROMBOSIS NOT LEADING TO MYOCARDIAL INFARCTION|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0340325|T047|194821006|SNOMEDCT_US|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION |CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0340325|T047|194821006|SNOMEDCT_US|CORONARY; THROMBOSIS, NOT RESULTING IN INFARCTION|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0340325|T047|194821006|SNOMEDCT_US|THROMBOEMBOLISM; CORONARY, NOT RESULTING IN INFARCTION|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0340325|T047|194821006|SNOMEDCT_US|THROMBOSIS; CARDIAC, NOT RESULTING IN INFARCTION|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0340325|T047|194821006|SNOMEDCT_US|THROMBOSIS; CORONARY, NOT RESULTING IN INFARCTION|CORONARY THROMBOSIS NOT RESULTING IN MYOCARDIAL INFARCTION (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PECTORIS|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|STENOCARDIAS|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PECTORIS, UNSPECIFIED|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|STENOCARDIA|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PECTORIS |ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINAL SYNDROME|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|CARDIAC ANGINA|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA OF EFFORT|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ISCHEMIC CHEST PAIN|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA NOS|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PECTORIS [DISEASE/FINDING]|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGOR PECTORIS|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|PAIN;ANGINA|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PECTORIS |ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA |ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PECTORIS NOS|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|STENOCARDIA |ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PECTORIS NOS |ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ISCHAEMIC CHEST PAIN|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ISCHAEMIC CHEST PAIN |ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|CHEST PAIN - CARDIAC|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|CHEST PAIN ISCHEMIC|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ISCHEMIC CHEST PAIN |ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINAL DISCOMFORT|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA SYNDROME|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINAL PAIN|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|CARDIO/PULM: ANGINA|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ISCHAEMIC HEART DISEASE - ANGINA|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ISCHEMIC HEART DISEASE - ANGINA|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|AP - ANGINA PECTORIS|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ISCHEMIC CHEST PAIN |ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|CHEST; PAIN, ISCHEMIC|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|PAIN; CHEST, ISCHEMIC|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|SYNDROME; ANGINAL|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINAL; SYNDROME|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PECTORIS, NOS|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA, NOS|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PECTORIS  [AMBIGUOUS]|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA, CARDIAC|ISCHAEMIC CHEST PAIN (DISORDER)
C0002962|T047|194835008|SNOMEDCT_US|ANGINA PAIN|ISCHAEMIC CHEST PAIN (DISORDER)
C0264692|T047|82522008|SNOMEDCT_US|ISCHEMIC CONTRACTURE OF LEFT VENTRICLE SYNDROME|ISCHEMIC CONTRACTURE OF LEFT VENTRICLE SYNDROME (DISORDER)
C0264692|T047|82522008|SNOMEDCT_US|STONE HEART SYNDROME|ISCHEMIC CONTRACTURE OF LEFT VENTRICLE SYNDROME (DISORDER)
C0264692|T047|82522008|SNOMEDCT_US|ISCHAEMIC CONTRACTURE OF LEFT VENTRICLE SYNDROME|ISCHEMIC CONTRACTURE OF LEFT VENTRICLE SYNDROME (DISORDER)
C0264692|T047|82522008|SNOMEDCT_US|ISCHEMIC CONTRACTURE OF LEFT VENTRICLE SYNDROME |ISCHEMIC CONTRACTURE OF LEFT VENTRICLE SYNDROME (DISORDER)
C1510446|T047|413439005|SNOMEDCT_US|ACUTE ISCHAEMIC HEART DISEASE, UNSPECIFIED|ACUTE ISCHEMIC HEART DISEASE (DISORDER)
C1510446|T047|413439005|SNOMEDCT_US|ACUTE ISCHEMIC HEART DISEASE, UNSPECIFIED|ACUTE ISCHEMIC HEART DISEASE (DISORDER)
C1510446|T047|413439005|SNOMEDCT_US|ACUTE ISCHEMIC HEART DISEASE |ACUTE ISCHEMIC HEART DISEASE (DISORDER)
C1510446|T047|413439005|SNOMEDCT_US|ACUTE ISCHEMIC HEART DISEASE|ACUTE ISCHEMIC HEART DISEASE (DISORDER)
C1510446|T047|413439005|SNOMEDCT_US|ACUTE ISCHEMIC HEART DISEASE |ACUTE ISCHEMIC HEART DISEASE (DISORDER)
C1510446|T047|413439005|SNOMEDCT_US|ACUTE ISCHAEMIC HEART DISEASE|ACUTE ISCHEMIC HEART DISEASE (DISORDER)
C0264684|T047|62827000|SNOMEDCT_US|ARTERITIS CORONARY|CORONARY ARTERITIS (DISORDER)
C0264684|T047|62827000|SNOMEDCT_US|CORONARY ARTERITIS|CORONARY ARTERITIS (DISORDER)
C0264684|T047|62827000|SNOMEDCT_US|CORONARY ENDARTERITIS|CORONARY ARTERITIS (DISORDER)
C0264684|T047|62827000|SNOMEDCT_US|CORONARY ARTERITIS |CORONARY ARTERITIS (DISORDER)
C0264684|T047|62827000|SNOMEDCT_US|CORONARY; ARTERITIS|CORONARY ARTERITIS (DISORDER)
C0264684|T047|62827000|SNOMEDCT_US|ARTERITIS; CORONARY|CORONARY ARTERITIS (DISORDER)
C0264684|T047|62827000|SNOMEDCT_US|CORONARY ARTERY ARTERITIS OR ENDARTERITIS|CORONARY ARTERITIS (DISORDER)
C0264684|T047|62827000|SNOMEDCT_US|CORONARY ARTERITIS OR ENDARTERITIS|CORONARY ARTERITIS (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|DRESSLER'S SYNDROME|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|POSTMYOCARDIAL INFARCTION SYNDROME|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|DRESSLER'S SYNDROME |POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|POST MI SYNDROME|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|DRESSLERS SYNDROME|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|POST MYOCARDIAL INFARCTION SYNDROME|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|POSTMYOCARDIAL INFARCTION PERICARDITIS|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|POST-MYOCARDIAL INFARCTION SYNDROME|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|POSTMYOCARDIAL INFARCTION SYNDROME |POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|POSTMYOCARDIAL INFARCTION; SYNDROME|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|SYNDROME; POSTMYOCARDIAL INFARCTION|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|DRESSLER|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C0152107|T047|66189004|SNOMEDCT_US|POSTMYOCARDIAL INFARCT SYNDROM|POSTMYOCARDIAL INFARCTION SYNDROME (DISORDER)
C1279369|T047|315348000|SNOMEDCT_US|ASYMPTOMATIC CORONARY HEART DISEASE |ASYMPTOMATIC CORONARY HEART DISEASE (DISORDER)
C1279369|T047|315348000|SNOMEDCT_US|ASYMPTOMATIC CORONARY HEART DISEASE|ASYMPTOMATIC CORONARY HEART DISEASE (DISORDER)
C0264695|T047|46109009|SNOMEDCT_US|SUBENDOCARDIAL ISCHAEMIA|SUBENDOCARDIAL ISCHEMIA (DISORDER)
C0264695|T047|46109009|SNOMEDCT_US|SUBENDOCARDIAL ISCHEMIA |SUBENDOCARDIAL ISCHEMIA (DISORDER)
C0264695|T047|46109009|SNOMEDCT_US|SUBENDOCARDIAL ISCHEMIA|SUBENDOCARDIAL ISCHEMIA (DISORDER)
C0264695|T047|46109009|SNOMEDCT_US|SUBENDOCARDIAL ISCHEMIA |SUBENDOCARDIAL ISCHEMIA (DISORDER)
C0264695|T047|46109009|SNOMEDCT_US|ISCHEMIA; SUBENDOCARDIAL|SUBENDOCARDIAL ISCHEMIA (DISORDER)
C0264687|T047|59062007|SNOMEDCT_US|CORONARY STRICTIRE|CORONARY STRICTURE (DISORDER)
C0264687|T047|59062007|SNOMEDCT_US|CORONARY STRICTIRE |CORONARY STRICTURE (DISORDER)
C0264687|T047|59062007|SNOMEDCT_US|CORONARY STRICTURE|CORONARY STRICTURE (DISORDER)
C0264687|T047|59062007|SNOMEDCT_US|CORONARY STRICTURE |CORONARY STRICTURE (DISORDER)
C0264687|T047|59062007|SNOMEDCT_US|CORONARY; STRICTURE|CORONARY STRICTURE (DISORDER)
C0264687|T047|59062007|SNOMEDCT_US|STRICTURE; CORONARY ARTERY|CORONARY STRICTURE (DISORDER)
C0264687|T047|59062007|SNOMEDCT_US|STRICTURE; CORONARY|CORONARY STRICTURE (DISORDER)
C0264687|T047|59062007|SNOMEDCT_US|CORONARY ARTERY STRICTURE|CORONARY STRICTURE (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|DISEASE, ISCHEMIC HEART|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|DISEASES, ISCHEMIC HEART|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|HEART DISEASES, ISCHEMIC|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIC HEART DISEASES|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIAL ISCHEMIA|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIAS, MYOCARDIAL|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIAL ISCHEMIAS|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHAEMIC HEART DISEASES|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIAL ISCHAEMIA|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIC HEART DISEASE|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|HEART DIS ISCHEMIC|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIC HEART DIS|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIAL ISCHEMIA |MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|HEART DISEASE, ISCHEMIC|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIA, MYOCARDIAL|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIAL ISCHEMIA [DISEASE/FINDING]|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|DISEASE;ISCHAEMIC HEART|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIAL ISCHEMIA/HYPOXIA|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIC HEART DISEASES (I20-I25)|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHAEMIC HEART DISEASE |MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|CARDIAC ISCHAEMIA|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHAEMIC HEART DISEASE|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHAEMIC HEART DISEASE NOS|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIC HEART DISEASE NOS|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|IHD - ISCHEMIC HEART DISEASE|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIC HEART DISEASE NOS |MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIAL ISCHAEMIA |MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|IHD - ISCHAEMIC HEART DISEASE|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIC HEART DISEASE |MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|CARDIAC ISCHEMIA|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHAEMIC HEART DISEASE NOS |MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIC HEART DISEASE |MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHAEMIA MYOCARDIAL|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIA MYOCARDIAL|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIA; HEART|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIA; MYOCARDIAL|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIUM; ISCHEMIC|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHEMIC HEART DISEASE, NOS|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|ISCHAEMIC HEART DISEASE, NOS|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIAL ISCHEMIA, NOS|MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|MYOCARDIAL ISCHEMIA |MYOCARDIAL ISCHEMIA (DISORDER)
C0151744|T047|414795007|SNOMEDCT_US|DISEASE;ISCHEMIC HEART|MYOCARDIAL ISCHEMIA (DISORDER)
C0340287|T047|194877008|SNOMEDCT_US|OTHER SPECIFIED ISCHAEMIC HEART DISEASE|OTHER SPECIFIED ISCHEMIC HEART DISEASE (DISORDER)
C0340287|T047|194877008|SNOMEDCT_US|OTHER SPECIFIED ISCHEMIC HEART DISEASE|OTHER SPECIFIED ISCHEMIC HEART DISEASE (DISORDER)
C0340287|T047|194877008|SNOMEDCT_US|OTHER SPECIFIED ISCHEMIC HEART DISEASE |OTHER SPECIFIED ISCHEMIC HEART DISEASE (DISORDER)
C0349466|T047|276516009|SNOMEDCT_US|MYOCARDIAL ISCHEMIA OF NEWBORN|MYOCARDIAL ISCHEMIA OF NEWBORN (DISORDER)
C0349466|T047|276516009|SNOMEDCT_US|MYOCARDIAL ISCHEMIA OF NEWBORN |MYOCARDIAL ISCHEMIA OF NEWBORN (DISORDER)
C0349466|T047|276516009|SNOMEDCT_US|MYOCARDIAL ISCHAEMIA OF NEWBORN|MYOCARDIAL ISCHEMIA OF NEWBORN (DISORDER)
C0349466|T047|276516009|SNOMEDCT_US|MYOCARDIAL ISCHEMIA OF NEWBORN |MYOCARDIAL ISCHEMIA OF NEWBORN (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE FORMS OF ISCHEMIC HEART DISEASE|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE FORMS OF ISCHAEMIC HEART DISEASE|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|AC ISCHEMIC HRT DIS NEC|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE FORMS OF ISCHEMIC HEART DISEASE, OTHER|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE ISCHEMIC HEART DISEASE|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE NOS|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE ISCHEMIC HEART DISEASE |OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE |OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE ISCHEMIC HEART DISEASE NOS|OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C0340283|T047|194822004|SNOMEDCT_US|OTHER ACUTE AND SUBACUTE ISCHEMIC HEART DISEASE NOS |OTHER ACUTE AND SUBACUTE ISCHAEMIC HEART DISEASE (DISORDER)
C1533195|T047|413844008|SNOMEDCT_US|CHRONIC CORONARY INSUFFICIENCY|CHRONIC CORONARY INSUFFICIENCY
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSMS, CARDIAC|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSMS, HEART|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|CARDIAC ANEURYSMS|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|HEART ANEURYSM|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|HEART ANEURYSMS|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM OF HEART|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM, CARDIAC|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM, HEART|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|CARDIAC ANEURYSM|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|HEART ANEURYSM [DISEASE/FINDING]|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM;CARDIAC|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM OF HEART NOS|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM OF HEART |ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM OF HEART NOS |ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|CARDIAC; ANEURYSM|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|HEART; ANEURYSM|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM; CARDIAC|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM; HEART|ANEURYSM OF HEART (DISORDER)
C0018789|T047|65340007|SNOMEDCT_US|ANEURYSM OF HEART, NOS|ANEURYSM OF HEART (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|CORONARY THROMBOSES|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|CORONARY THROMBOSIS|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|THROMBOSES, CORONARY|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|CORONARY ARTERY THROMBOSIS|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|CORONARY ARTERY THROMBOSIS |CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|CORONARY (ARTERY) THROMBOSIS|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|CORONARY THROMBOSIS [DISEASE/FINDING]|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|THROMBOSIS, CORONARY|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|THROMBOSIS;ARTERY;CORONARY|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|CORONARY ARTERY THROMBOSIS |CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|CT - CORONARY THROMBOSIS|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|THROMBOSIS - CORONARY|CORONARY ARTERY THROMBOSIS (DISORDER)
C0010072|T047|398274000|SNOMEDCT_US|THROMBOSIS CORONARY|CORONARY ARTERY THROMBOSIS (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|CORONARY (ARTERY) ATHEROMA|CORONARY ARTERY ATHEROMA (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|CORONARY ATHEROMA|CORONARY ARTERY ATHEROMA (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|CORONARY ARTERY ATHEROMA |CORONARY ARTERY ATHEROMA (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|CORONARY ARTERY ATHEROMA|CORONARY ARTERY ATHEROMA (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|ATHEROMA CORONARY ARTERY|CORONARY ARTERY ATHEROMA (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|CORONARY ARTERY ATHEROMA |CORONARY ARTERY ATHEROMA (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|ATHEROMA; CORONARY|CORONARY ARTERY ATHEROMA (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|ATHEROMA; HEART|CORONARY ARTERY ATHEROMA (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|CORONARY; ATHEROMA|CORONARY ARTERY ATHEROMA (DISORDER)
C0264683|T047|67682002|SNOMEDCT_US|HEART; ATHEROMA|CORONARY ARTERY ATHEROMA (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER FORMS OF CHRONIC ISCHEMIC HEART DISEASE|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER FORMS OF CHRONIC ISCHAEMIC HEART DISEASE|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER FORMS OF CHRONIC ISCHEMIC HEART DISEASE, OTHER|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER FORMS OF CHRONIC ISCHAEMIC HEART DISEASE, OTHER|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|[X]OTHER FORMS OF CHRONIC ISCHAEMIC HEART DISEASE|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|[X]OTHER FORMS OF CHRONIC ISCHEMIC HEART DISEASE |OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER CHRONIC ISCHAEMIC HEART DISEASE|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|[X]OTHER FORMS OF CHRONIC ISCHEMIC HEART DISEASE|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER CHRONIC ISCHAEMIC HEART DISEASE NOS|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER CHRONIC ISCHEMIC HEART DISEASE|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER CHRONIC ISCHEMIC HEART DISEASE |OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0155669|T047|194854008|SNOMEDCT_US|OTHER CHRONIC ISCHEMIC HEART DISEASE NOS |OTHER CHRONIC ISCHEMIC HEART DISEASE NOS (DISORDER)
C0348589|T047|195542009|SNOMEDCT_US|OTHER CURRENT COMPLICATIONS FOLLOWING ACUTE MYOCARDIAL INFARCTION|[X]OTHER CURRENT COMPLICATIONS FOLLOWING ACUTE MYOCARDIAL INFARCTION (DISORDER)
C0348589|T047|195542009|SNOMEDCT_US|OTH CURRENT COMPLICATIONS FOLLOWING AMI|[X]OTHER CURRENT COMPLICATIONS FOLLOWING ACUTE MYOCARDIAL INFARCTION (DISORDER)
C0348589|T047|195542009|SNOMEDCT_US|[X]OTHER CURRENT COMPLICATIONS FOLLOWING ACUTE MYOCARDIAL INFARCTION |[X]OTHER CURRENT COMPLICATIONS FOLLOWING ACUTE MYOCARDIAL INFARCTION (DISORDER)
C0348589|T047|195542009|SNOMEDCT_US|[X]OTHER CURRENT COMPLICATIONS FOLLOWING ACUTE MYOCARDIAL INFARCTION|[X]OTHER CURRENT COMPLICATIONS FOLLOWING ACUTE MYOCARDIAL INFARCTION (DISORDER)
C0009693|T047|42866003|SNOMEDCT_US|CONGENITAL CORONARY ARTERY SCLEROSIS|CONGENITAL CORONARY ARTERY SCLEROSIS (DISORDER)
C0009693|T047|42866003|SNOMEDCT_US|CONGENITAL CORONARY ARTERY SCLEROSIS |CONGENITAL CORONARY ARTERY SCLEROSIS (DISORDER)
C0340291|T047|233823002|SNOMEDCT_US|SILENT MYOCARDIAL ISCHAEMIA|SILENT MYOCARDIAL ISCHEMIA (DISORDER)
C0340291|T047|233823002|SNOMEDCT_US|SILENT MYOCARDIAL ISCHEMIA|SILENT MYOCARDIAL ISCHEMIA (DISORDER)
C0340291|T047|233823002|SNOMEDCT_US|SILENT MYOCARDIAL ISCHEMIA |SILENT MYOCARDIAL ISCHEMIA (DISORDER)
C0340291|T047|233823002|SNOMEDCT_US|SILENT MYOCARDIAL ISCHAEMIA |SILENT MYOCARDIAL ISCHEMIA (DISORDER)
C0340291|T047|233823002|SNOMEDCT_US|SILENT MYOCARDIAL ISCHEMIA |SILENT MYOCARDIAL ISCHEMIA (DISORDER)
C0340291|T047|233823002|SNOMEDCT_US|ASYMPTOMATIC ISCHAEMIA|SILENT MYOCARDIAL ISCHEMIA (DISORDER)
C0340291|T047|233823002|SNOMEDCT_US|ASYMPTOMATIC ISCHEMIA|SILENT MYOCARDIAL ISCHEMIA (DISORDER)
C0340291|T047|233823002|SNOMEDCT_US|ISCHEMIA; MYOCARDIAL, SUBCLINICAL|SILENT MYOCARDIAL ISCHEMIA (DISORDER)
C0581375|T047|194843003|SNOMEDCT_US|2-VESSEL CORONARY ARTERY STENOSIS |DOUBLE CORONARY VESSEL DISEASE (DISORDER)
C0581375|T047|194843003|SNOMEDCT_US|2-VESSEL CORONARY ARTERY STENOSIS|DOUBLE CORONARY VESSEL DISEASE (DISORDER)
C0581375|T047|194843003|SNOMEDCT_US|TWO VESSEL CORONARY DISEASE|DOUBLE CORONARY VESSEL DISEASE (DISORDER)
C0581375|T047|194843003|SNOMEDCT_US|DOUBLE VESSEL CORONARY ARTERY DISEASE|DOUBLE CORONARY VESSEL DISEASE (DISORDER)
C0581375|T047|194843003|SNOMEDCT_US|DOUBLE VESSEL CORONARY ARTERY DISEASE |DOUBLE CORONARY VESSEL DISEASE (DISORDER)
C0581375|T047|194843003|SNOMEDCT_US|TWO VESSEL DISEASE|DOUBLE CORONARY VESSEL DISEASE (DISORDER)
C0581375|T047|194843003|SNOMEDCT_US|DOUBLE CORONARY VESSEL DISEASE|DOUBLE CORONARY VESSEL DISEASE (DISORDER)
C0581375|T047|194843003|SNOMEDCT_US|TWO CORONARY VESSEL DISEASE|DOUBLE CORONARY VESSEL DISEASE (DISORDER)
C0581375|T047|194843003|SNOMEDCT_US|DOUBLE CORONARY VESSEL DISEASE |DOUBLE CORONARY VESSEL DISEASE (DISORDER)
C0581374|T047|194842008|SNOMEDCT_US|SINGLE VESSEL CORONARY ARTERY STENOSIS|SINGLE CORONARY VESSEL DISEASE (DISORDER)
C0581374|T047|194842008|SNOMEDCT_US|SINGLE VESSEL CORONARY ARTERY STENOSIS |SINGLE CORONARY VESSEL DISEASE (DISORDER)
C0581374|T047|194842008|SNOMEDCT_US|SINGLE VESSEL CORONARY ARTERY DISEASE |SINGLE CORONARY VESSEL DISEASE (DISORDER)
C0581374|T047|194842008|SNOMEDCT_US|SINGLE VESSEL CORONARY ARTERY DISEASE|SINGLE CORONARY VESSEL DISEASE (DISORDER)
C0581374|T047|194842008|SNOMEDCT_US|SINGLE CORONARY VESSEL DISEASE|SINGLE CORONARY VESSEL DISEASE (DISORDER)
C0581374|T047|194842008|SNOMEDCT_US|SINGLE CORONARY VESSEL DISEASE |SINGLE CORONARY VESSEL DISEASE (DISORDER)
C0264696|T047|194824003|SNOMEDCT_US|MICROINFARCTION OF HEART|MICROINFARCTION OF HEART (DISORDER)
C0264696|T047|194824003|SNOMEDCT_US|MICROINFARCTION OF HEART |MICROINFARCTION OF HEART (DISORDER)
C0264696|T047|194824003|SNOMEDCT_US|MICROINFARCT OF HEART |MICROINFARCTION OF HEART (DISORDER)
C0264696|T047|194824003|SNOMEDCT_US|MICROINFARCT OF HEART|MICROINFARCTION OF HEART (DISORDER)
C0264696|T047|194824003|SNOMEDCT_US|MICROINFARCT OF HEART |MICROINFARCTION OF HEART (DISORDER)
C0264696|T047|194824003|SNOMEDCT_US|MICROINFARCT; HEART|MICROINFARCTION OF HEART (DISORDER)
C0349780|T047|281091000|SNOMEDCT_US|ISCHEMIC MYOCARDIAL DYSFUNCTION |ISCHEMIC MYOCARDIAL DYSFUNCTION (DISORDER)
C0349780|T047|281091000|SNOMEDCT_US|ISCHEMIC MYOCARDIAL DYSFUNCTION|ISCHEMIC MYOCARDIAL DYSFUNCTION (DISORDER)
C0349780|T047|281091000|SNOMEDCT_US|ISCHAEMIC MYOCARDIAL DYSFUNCTION|ISCHEMIC MYOCARDIAL DYSFUNCTION (DISORDER)
C0349780|T047|281091000|SNOMEDCT_US|ISCHEMIC MYOCARDIAL DYSFUNCTION |ISCHEMIC MYOCARDIAL DYSFUNCTION (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHEMIC HEART DISEASE|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHEMIC HEART DISEASE, UNSPECIFIED|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHAEMIC HEART DISEASE|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHAEMIC HEART DISEASE, UNSPECIFIED|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC MYOCARDIAL ISCHEMIA|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC MYOCARDIAL ISCHEMIA |CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHR ISCHEMIC HRT DIS NOS|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|ISCHEMIC HEART DISEASE (CHRONIC) NOS|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|ISCHAEMIA;MYOCARDIAL;CHRONIC|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHEMIC HEART DISEASE |CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHR. ISCHEMIC HEART DIS. NOS|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHAEMIC HEART DISEASE NOS|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHEMIC HEART DISEASE NOS|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHEMIC HEART DISEASE |CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHEMIC HEART DISEASE NOS |CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC MYOCARDIAL ISCHAEMIA|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHR. ISCHAEMIC HEART DIS. NOS|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC MYOCARDIAL ISCHAEMIA |CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC ISCHAEMIC HEART DISEASE NOS |CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|CHRONIC MYOCARDIAL ISCHEMIA |CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|DISEASE;ISCHAEM HEART;CHRONIC|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C0264694|T047|413844008|SNOMEDCT_US|ISCHEMIA;MYOCARDIAL;CHRONIC|CHRONIC MYOCARDIAL ISCHEMIA (DISORDER)
C3650149|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF OTHER CORONARY VESSELS 
C3650149|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF OTHER CORONARY VESSELS
C3650188|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY WITH UNSTABLE ANGINA PECTORIS 
C3650188|T047||SNOMEDCT_US|ATHEROSCLEROSIS CORONARY ARTERY WITH UNSTABLE ANGINA PECTORIS
C3650188|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY WITH UNSTABLE ANGINA PECTORIS
C3650187|T047|451041000124103|SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY WITHOUT ANGINA PECTORIS|ATHEROSCLEROSIS OF CORONARY ARTERY WITHOUT ANGINA PECTORIS (DISORDER)
C3650187|T047|451041000124103|SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY WITHOUT ANGINA PECTORIS |ATHEROSCLEROSIS OF CORONARY ARTERY WITHOUT ANGINA PECTORIS (DISORDER)
C3650187|T047|451041000124103|SNOMEDCT_US|ATHEROSCLEROSIS CORONARY ARTERY WITHOUT ANGINA PECTORIS|ATHEROSCLEROSIS OF CORONARY ARTERY WITHOUT ANGINA PECTORIS (DISORDER)
C2882208|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF OTHER CORONARY VESSELS WITHOUT ANGINA PECTORIS
C2882208|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF OTHER CORONARY VESSELS WITHOUT ANGINA PECTORIS 
C3650190|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY WITH ANGINA PECTORIS
C3650190|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY WITH ANGINA PECTORIS 
C3650190|T047||SNOMEDCT_US|ATHEROSCLEROSIS CORONARY ARTERY WITH ANGINA PECTORIS
C3650189|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY WITH ANGINA PECTORIS WITH DOCUMENTED SPASM
C3650189|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY WITH ANGINA PECTORIS WITH DOCUMENTED SPASM 
C3650189|T047||SNOMEDCT_US|ATHEROSCLEROSIS CORONARY ARTERY WITH ANGINA PECTORIS WITH DOCUMENTED SPASM
C2349509|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS DUE TO LIPID RICH PLAQUE
C2349509|T047||SNOMEDCT_US|COR ATH D/T LPD RCH PLAQ
C2349509|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS DUE TO LIPID-RICH PLAQUE
C2349509|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS DUE TO LIPID-RICH PLAQUE 
C3161090|T047||SNOMEDCT_US|COR ATH D/T CALC COR LSN
C3161090|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS DUE TO CALCIFIED CORONARY LESION
C3161090|T047||SNOMEDCT_US|ATHEROSCLEROSIS DUE CALCIFIED CORONARY LESION
C3161090|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS DUE CALCIFIED CORONARY LESION
C3161090|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS DUE TO CALCIFIED CORONARY LESION 
C1867743|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE, PREMATURE
C1867743|T047||SNOMEDCT_US|PREMATURE CORONARY HEART DISEASE
C1867743|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE PREMATURE
C1867743|T047||SNOMEDCT_US|PREMATURE CORONARY HEART DISEASE 
C1867743|T047||SNOMEDCT_US|PREMATURE CORONARY ARTERY DISEASE
C1997109|T047|429673002|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT|ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT (DISORDER)
C1997109|T047|429673002|SNOMEDCT_US|ARTERIOSCLEROSIS IN CORONARY ARTERY BYPASS GRAFT|ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT (DISORDER)
C1997109|T047|429673002|SNOMEDCT_US|ARTERIOSCLEROSIS IN CORONARY ARTERY BYPASS GRAFT |ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT (DISORDER)
C1997109|T047|429673002|SNOMEDCT_US|ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT |ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT (DISORDER)
C1997109|T047|429673002|SNOMEDCT_US|ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT|ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT (DISORDER)
C1997109|T047|429673002|SNOMEDCT_US|ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT |ARTERIOSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT (DISORDER)
C1996973|T047|429245005|SNOMEDCT_US|RECURRENT CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS TRANSLUMINAL CORONARY ANGIOPLASTY |RECURRENT CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS TRANSLUMINAL CORONARY ANGIOPLASTY (DISORDER)
C1996973|T047|429245005|SNOMEDCT_US|RECURRENT CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS TRANSLUMINAL CORONARY ANGIOPLASTY|RECURRENT CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS TRANSLUMINAL CORONARY ANGIOPLASTY (DISORDER)
C1996973|T047|429245005|SNOMEDCT_US|RECURRENT CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS TRANSLUMINAL CORONARY ANGIOPLASTY |RECURRENT CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS TRANSLUMINAL CORONARY ANGIOPLASTY (DISORDER)
C1996973|T047|429245005|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS RECURRENT AFTER PERCUTANEOUS TRANSLUMINAL ANGIOPLASTY|RECURRENT CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS TRANSLUMINAL CORONARY ANGIOPLASTY (DISORDER)
C1842247|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE, AUTOSOMAL DOMINANT, 1
C1842247|T047||SNOMEDCT_US|ADCAD1
C1842247|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE WITH MYOCARDIAL INFARCTION
C1842247|T047||SNOMEDCT_US|CAD AUTOSOMAL DOMINANT 1 
C1842247|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE AUTOSOMAL DOMINANT 1
C1842247|T047||SNOMEDCT_US|CAD AUTOSOMAL DOMINANT 1
C1842247|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE, AUTOSOMAL DOMINANT 1
C1842247|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE/MYOCARDIAL INFARCTION
C1970440|T047||SNOMEDCT_US|ADCAD2
C1970440|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE, AUTOSOMAL DOMINANT 2
C1970440|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE, AUTOSOMAL DOMINANT 2 
C1970440|T047||SNOMEDCT_US|CAD AUTOSOMAL DOMINANT 2 
C1970440|T047||SNOMEDCT_US|CAD AUTOSOMAL DOMINANT 2
C1970440|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE AUTOSOMAL DOMINANT 2
C4039929|T047|11018701000119109|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS CORONARY ANGIOPLASTY|CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS CORONARY ANGIOPLASTY (DISORDER)
C4039929|T047|11018701000119109|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS CORONARY ANGIOPLASTY |CORONARY ARTERIOSCLEROSIS AFTER PERCUTANEOUS CORONARY ANGIOPLASTY (DISORDER)
C4074915|T047|139011000119104|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS FOLLOWING CORONARY ARTERY BYPASS GRAFT |CORONARY ARTERIOSCLEROSIS FOLLOWING CORONARY ARTERY BYPASS GRAFT (DISORDER)
C4074915|T047|139011000119104|SNOMEDCT_US|CORONARY ARTERIOSCLEROSIS FOLLOWING CORONARY ARTERY BYPASS GRAFT|CORONARY ARTERIOSCLEROSIS FOLLOWING CORONARY ARTERY BYPASS GRAFT (DISORDER)
C0340326|T047|233844002|SNOMEDCT_US|ACCELERATED CORONARY ARTERY DISEASE IN TRANSPLANTED HEART |ACCELERATED CORONARY ARTERY DISEASE IN TRANSPLANTED HEART (DISORDER)
C0340326|T047|233844002|SNOMEDCT_US|CORONARY ARTERY DISEASE IN TRANSPLANTED HEART ACCELERATED|ACCELERATED CORONARY ARTERY DISEASE IN TRANSPLANTED HEART (DISORDER)
C0340326|T047|233844002|SNOMEDCT_US|ACCELERATED CORONARY ARTERY DISEASE IN TRANSPLANTED HEART|ACCELERATED CORONARY ARTERY DISEASE IN TRANSPLANTED HEART (DISORDER)
C0340326|T047|233844002|SNOMEDCT_US|ACCELERATED CORONARY ARTERY DISEASE IN TRANSPLANTED HEART |ACCELERATED CORONARY ARTERY DISEASE IN TRANSPLANTED HEART (DISORDER)
C1299432|T047|371803003|SNOMEDCT_US|MULTI VESSEL CORONARY ARTERY DISEASE|MULTI VESSEL CORONARY ARTERY DISEASE (DISORDER)
C1299432|T047|371803003|SNOMEDCT_US|MULTI VESSEL CORONARY ARTERY DISEASE |MULTI VESSEL CORONARY ARTERY DISEASE (DISORDER)
C1299432|T047|371803003|SNOMEDCT_US|MULTI VESSEL CORONARY ARTERY DISEASE |MULTI VESSEL CORONARY ARTERY DISEASE (DISORDER)
C1299433|T047|371804009|SNOMEDCT_US|LEFT MAIN CORONARY ARTERY DISEASE |LEFT MAIN CORONARY ARTERY DISEASE (DISORDER)
C1299433|T047|371804009|SNOMEDCT_US|LEFT MAIN CORONARY ARTERY DISEASE|LEFT MAIN CORONARY ARTERY DISEASE (DISORDER)
C1299433|T047|371804009|SNOMEDCT_US|CORONARY ARTERY DISEASE LEFT MAIN|LEFT MAIN CORONARY ARTERY DISEASE (DISORDER)
C1299433|T047|371804009|SNOMEDCT_US|LEFT MAIN CORONARY ARTERY DISEASE |LEFT MAIN CORONARY ARTERY DISEASE (DISORDER)
C1299434|T047|371805005|SNOMEDCT_US|CORONARY ARTERY DISEASE OF SIGNIFICANT BYPASS GRAFT|SIGNIFICANT CORONARY BYPASS GRAFT DISEASE (DISORDER)
C1299434|T047|371805005|SNOMEDCT_US|SIGNIFICANT CORONARY BYPASS GRAFT DISEASE |SIGNIFICANT CORONARY BYPASS GRAFT DISEASE (DISORDER)
C1299434|T047|371805005|SNOMEDCT_US|SIGNIFICANT CORONARY BYPASS GRAFT DISEASE|SIGNIFICANT CORONARY BYPASS GRAFT DISEASE (DISORDER)
C1299434|T047|371805005|SNOMEDCT_US|SIGNIFICANT CORONARY BYPASS GRAFT DISEASE |SIGNIFICANT CORONARY BYPASS GRAFT DISEASE (DISORDER)
C1384784|T047||SNOMEDCT_US|A.CORONARIA; OBSTRUCTION
C1384784|T047||SNOMEDCT_US|OBSTRUCTION; CORONARY ARTERY
C1384785|T047||SNOMEDCT_US|A.CORONARIA; STRICTURE, CORONARY
C0242231|T047|233970002|SNOMEDCT_US|CORONARY STENOSIS|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|STENOSES, CORONARY|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|STENOSIS, CORONARY|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|CORONARY ARTERY STENOSIS|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|CORONARY ARTERY STENOSIS |CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|CORONARY STENOSIS [DISEASE/FINDING]|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|CORONARY STENOSES|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|ARTERY STENOSES, CORONARY|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|ARTERY STENOSIS, CORONARY|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|CORONARY ARTERY STENOSES|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|STENOSES, CORONARY ARTERY|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|STENOSIS, CORONARY ARTERY|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|NARROW CORONARY ARTERIES|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|CORONARY ARTERIES--STENOSIS|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|CORONARY ARTERY STENOSIS |CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|CORONARY; STENOSIS|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|A.CORONARIA; NARROWING|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|NARROWING; CORONARY ARTERY|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|STENOSIS; ARTERY, CORONARY|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|STENOSIS; CORONARY|CORONARY ARTERY STENOSIS (DISORDER)
C0242231|T047|233970002|SNOMEDCT_US|ARTERY; STENOSIS, CORONARY|CORONARY ARTERY STENOSIS (DISORDER)
C1384962|T047||SNOMEDCT_US|DISEASE (OR DISORDER); HEART, ARTERIOSCLEROTIC OR SCLEROTIC (SENILE)
C1388510|T047||SNOMEDCT_US|CARDIAC; ARTERIOSCLEROSIS
C1388510|T047||SNOMEDCT_US|ARTERIOSCLEROSIS; CARDIAC
C1388511|T047||SNOMEDCT_US|ARTERIOSCLEROSIS; CARDIOMYOPATHY
C1388512|T047||SNOMEDCT_US|ARTERIOSCLEROSIS; CARDIOPATHY
C1404464|T047||SNOMEDCT_US|ATHEROMA; MYOCARDIAL
C1404464|T047||SNOMEDCT_US|MYOCARDIUM; ATHEROMA
C1391994|T047||SNOMEDCT_US|CARDIOMYOPATHY; ARTERIOSCLEROTIC
C1392010|T047||SNOMEDCT_US|CARDIOPATHY; ARTERIOSCLEROTIC
C1392034|T047||SNOMEDCT_US|CARDIOSCLEROSIS
C1394006|T047||SNOMEDCT_US|CORONARY; OBSTRUCTION
C1394006|T047||SNOMEDCT_US|OBSTRUCTION; CORONARY
C1399178|T047||SNOMEDCT_US|CARDIAC; OSSIFICATION
C1399178|T047||SNOMEDCT_US|CORONARY; OSSIFICATION
C1399178|T047||SNOMEDCT_US|HEART; OSSIFICATION
C1399178|T047||SNOMEDCT_US|OSSIFICATION; CARDIAC
C1399178|T047||SNOMEDCT_US|OSSIFICATION; CORONARY
C1399178|T047||SNOMEDCT_US|OSSIFICATION; HEART
C1394968|T047||SNOMEDCT_US|DEGENERATION; HEART, ATHEROMATOUS
C1394968|T047||SNOMEDCT_US|HEART; DEGENERATION, ATHEROMATOUS
C1399129|T047||SNOMEDCT_US|HEART; DISEASE, ARTERY, ARTERIAL
C1399130|T047||SNOMEDCT_US|HEART; DISEASE, ARTERIOSCLEROTIC OR SCLEROTIC (SENILE)
C1328505|T047||SNOMEDCT_US|MYOCARDIAL SCLEROSIS
C1328505|T047||SNOMEDCT_US|MYOCARDIUM; SCLEROSIS
C1328505|T047||SNOMEDCT_US|SCLEROSIS; MYOCARDIAL
C1636672|T047|420006002|SNOMEDCT_US|CORONARY ARTERY DISEASE OBLITERATIVE|OBLITERATIVE CORONARY ARTERY DISEASE (DISORDER)
C1636672|T047|420006002|SNOMEDCT_US|OBLITERATIVE CORONARY ARTERY DISEASE |OBLITERATIVE CORONARY ARTERY DISEASE (DISORDER)
C1636672|T047|420006002|SNOMEDCT_US|OBLITERATIVE CORONARY ARTERY DISEASE|OBLITERATIVE CORONARY ARTERY DISEASE (DISORDER)
C1636672|T047|420006002|SNOMEDCT_US|OBLITERATIVE CORONARY ARTERY DISEASE |OBLITERATIVE CORONARY ARTERY DISEASE (DISORDER)
C0837136|T047||SNOMEDCT_US|CRN ATH NONATLG BLG GRFT
C0837136|T047||SNOMEDCT_US|ATHEROSCLEROTIC HEART DISEASE, OF NONAUTOLOGOUS BYPASS GRAFT
C0837136|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF NONAUTOLOGOUS BIOLOGICAL BYPASS GRAFT
C0837134|T047||SNOMEDCT_US|CRNRY ATHRSCL NATVE VSSL
C0837134|T047||SNOMEDCT_US|ATHEROSCLEROTIC HEART DISEASE OF NATIVE CORONARY ARTERY
C0837134|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF NATIVE CORONARY ARTERY
C0837133|T047||SNOMEDCT_US|COR ATH UNSP VSL NTV/GFT
C0837133|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF UNSPECIFIED TYPE OF VESSEL, NATIVE OR GRAFT
C0837135|T047||SNOMEDCT_US|CRN ATH ATLG VN BPS GRFT
C0837135|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF AUTOLOGOUS VEIN BYPASS GRAFT
C0837135|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF AUTOLOGOUS BIOLOGICAL BYPASS GRAFT
C1456095|T047||SNOMEDCT_US|COR ATH BPS GRAFT TP HRT
C1456095|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF BYPASS GRAFT (ARTERY) (VEIN) OF TRANSPLANTED HEART
C0375264|T047||SNOMEDCT_US|COR ATH ARTRY BYPAS GRFT
C0375264|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT NOS
C0375264|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT 
C0375264|T047||SNOMEDCT_US|ATHEROSCLEROSIS OF CORONARY ARTERY BYPASS GRAFT
C0375264|T047||SNOMEDCT_US|ATHEROSCLEROSIS CORONARY ARTERY BYPASS GRAFT
C0375264|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF ARTERY BYPASS GRAFT
C1135190|T047||SNOMEDCT_US|COR ATH NATV ART TP HRT
C1135190|T047||SNOMEDCT_US|CORONARY ATHEROSCLEROSIS OF NATIVE CORONARY ARTERY OF TRANSPLANTED HEART
C0852153|T047||SNOMEDCT_US|CORONARY ARTERY DISORDERS NEC
C0852149|T047||SNOMEDCT_US|ISCHAEMIC CORONARY ARTERY DISORDERS
C0852149|T047||SNOMEDCT_US|ISCHEMIC CORONARY ARTERY DISORDERS
C2584623|T047|440444007|SNOMEDCT_US|FURCATION LESION OF CORONARY ARTERY|FURCATION LESION OF CORONARY ARTERY (DISORDER)
C2584623|T047|440444007|SNOMEDCT_US|FURCATION LESION OF CORONARY ARTERY |FURCATION LESION OF CORONARY ARTERY (DISORDER)
C2711976|T047|442298000|SNOMEDCT_US|FRACTURE OF STENT OF CORONARY ARTERY |FRACTURE OF STENT OF CORONARY ARTERY (DISORDER)
C2711976|T047|442298000|SNOMEDCT_US|FRACTURE OF STENT OF CORONARY ARTERY|FRACTURE OF STENT OF CORONARY ARTERY (DISORDER)
C1611184|T047|445512009|SNOMEDCT_US|CORONARY ARTERY CALCIFICATION|CALCIFICATION OF CORONARY ARTERY (DISORDER)
C1611184|T047|445512009|SNOMEDCT_US|CALCIFICATION OF CORONARY ARTERY |CALCIFICATION OF CORONARY ARTERY (DISORDER)
C1611184|T047|445512009|SNOMEDCT_US|CALCIFICATION OF CORONARY ARTERY|CALCIFICATION OF CORONARY ARTERY (DISORDER)
C2062867|T047||SNOMEDCT_US|REBOUND ANGINA DUE TO BETA BLOCKER WITHDRAWAL
C2062867|T047||SNOMEDCT_US|BETA-BLOCKER WITHDRAWAL (REBOUND ANGINA)
C2062867|T047||SNOMEDCT_US|REBOUND ANGINA DUE TO BETA BLOCKER WITHDRAWAL 
C0003851|T047|361133006|SNOMEDCT_US|ARTERIOSCLEROSIS OBLITERANS|ARTERIOSCLEROSIS OBLITERANS (DISORDER)
C0003851|T047|361133006|SNOMEDCT_US|OBLITERANS, ARTERIOSCLEROSIS|ARTERIOSCLEROSIS OBLITERANS (DISORDER)
C0003851|T047|361133006|SNOMEDCT_US|ARTERIOSCLEROSIS OBLITERANS |ARTERIOSCLEROSIS OBLITERANS (DISORDER)
C0003851|T047|361133006|SNOMEDCT_US|ARTERIOSCLEROSIS OBLITERANS [DISEASE/FINDING]|ARTERIOSCLEROSIS OBLITERANS (DISORDER)
C0003851|T047|361133006|SNOMEDCT_US|ARTERIOSCLEROSIS OBLITERANS |ARTERIOSCLEROSIS OBLITERANS (DISORDER)
C0003851|T047|361133006|SNOMEDCT_US|ARTERIOSCLEROSIS OBLITERANS  [AMBIGUOUS]|ARTERIOSCLEROSIS OBLITERANS (DISORDER)
C0264686|T047|29899005|SNOMEDCT_US|CORONARY ARTERY EMBOLISM|CORONARY ARTERY EMBOLISM (DISORDER)
C0264686|T047|29899005|SNOMEDCT_US|CORONARY ARTERY EMBOLISM |CORONARY ARTERY EMBOLISM (DISORDER)
C0264686|T047|29899005|SNOMEDCT_US|CORONARY (ARTERY) EMBOLISM|CORONARY ARTERY EMBOLISM (DISORDER)
C0264686|T047|29899005|SNOMEDCT_US|EMBOLISM;ARTERY;CORONARY|CORONARY ARTERY EMBOLISM (DISORDER)
C0264686|T047|29899005|SNOMEDCT_US|CORONARY EMBOLISM|CORONARY ARTERY EMBOLISM (DISORDER)
C0264686|T047|29899005|SNOMEDCT_US|EMBOLUS CORONARY ARTERY|CORONARY ARTERY EMBOLISM (DISORDER)
C0264686|T047|29899005|SNOMEDCT_US|CORONARY EMBOLUS|CORONARY ARTERY EMBOLISM (DISORDER)
C0264686|T047|29899005|SNOMEDCT_US|CORONARY ARTERY EMBOLISM |CORONARY ARTERY EMBOLISM (DISORDER)
C2049072|T047||SNOMEDCT_US|INDUCED CPK ELEVATION
C2049072|T047||SNOMEDCT_US|INDUCED CPK ELEVATION 
C2024793|T047||SNOMEDCT_US|CARDIAC WALL MOTION DYSFUNCTION 
C2024793|T047||SNOMEDCT_US|CARDIAC WALL MOTION DYSFUNCTION
C0010073|T047|23687008|SNOMEDCT_US|SAME PRINCIPLES AS PRINZMETAL ANGINA - FALSE POSITIVE IN THE STRICTEST SENSE OF CAD, BUT INCLUDING FOR NOW|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|ARTERY VASOSPASMS, CORONARY|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY ARTERY VASOSPASMS|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY VASOSPASM|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY VASOSPASMS|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|VASOSPASM, CORONARY|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|VASOSPASM, CORONARY ARTERY|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|VASOSPASMS, CORONARY|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|VASOSPASMS, CORONARY ARTERY|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY ARTERY SPASM|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY ARTERY SPASM |CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|ARTERIOSPASM CORONARY|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY VASOSPASM [DISEASE/FINDING]|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY ARTERY VASOSPASM|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|SPASM;ARTERY;CORONARY|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY SPASM|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY VASCULAR SPASM|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|SPASM CORONARY ARTERY|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY ARTERY SPASM |CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|CORONARY; SPASM|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|A.CORONARIA; SPASM|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|SPASM; CORONARY ARTERY|CORONARY ARTERY SPASM (DISORDER)
C0010073|T047|23687008|SNOMEDCT_US|SPASM; CORONARY|CORONARY ARTERY SPASM (DISORDER)
C0428837|T047|251032001|SNOMEDCT_US|CORONARY COLLATERAL CIRCULATION |CORONARY ARTERY COLLATERALS (FINDING)
C0428837|T047|251032001|SNOMEDCT_US|CORONARY COLLATERAL CIRCULATION|CORONARY ARTERY COLLATERALS (FINDING)
C0428837|T047|251032001|SNOMEDCT_US|CORONARY ARTERY COLLATERALS|CORONARY ARTERY COLLATERALS (FINDING)
C0428837|T047|251032001|SNOMEDCT_US|CORONARY ARTERY COLLATERALS |CORONARY ARTERY COLLATERALS (FINDING)
C2063730|T047||SNOMEDCT_US|SEPERATE BUT RELATED
C2063730|T047||SNOMEDCT_US|CORONARY ECTASIA 
C2063731|T047||SNOMEDCT_US|CONGENITAL DISEASE
C2063731|T047||SNOMEDCT_US|CORONARY OSTIAL MEMBRANE 
C0428830|T047|251024009|SNOMEDCT_US|CORONARY BYPASS GRAFT STENOSIS |CORONARY GRAFT STENOSIS (DISORDER)
C0428830|T047|251024009|SNOMEDCT_US|CORONARY BYPASS GRAFT STENOSIS|CORONARY GRAFT STENOSIS (DISORDER)
C0428830|T047|251024009|SNOMEDCT_US|CORONARY GRAFT STENOSIS|CORONARY GRAFT STENOSIS (DISORDER)
C0428830|T047|251024009|SNOMEDCT_US|CORONARY GRAFT; STENOSIS|CORONARY GRAFT STENOSIS (DISORDER)
C0428830|T047|251024009|SNOMEDCT_US|STENOSIS; CORONARY GRAFT|CORONARY GRAFT STENOSIS (DISORDER)
C0428830|T047|251024009|SNOMEDCT_US|CORONARY GRAFT STENOSIS |CORONARY GRAFT STENOSIS (DISORDER)
C0428830|T047|251024009|SNOMEDCT_US|CORONARY GRAFT STENOSIS |CORONARY GRAFT STENOSIS (DISORDER)
C0349781|T047|281093002|SNOMEDCT_US|HIBERNATING MYOCARDIUM |HIBERNATING MYOCARDIUM (DISORDER)
C0349781|T047|281093002|SNOMEDCT_US|HIBERNATING MYOCARDIUM|HIBERNATING MYOCARDIUM (DISORDER)
C0349781|T047|281093002|SNOMEDCT_US|HIBERNATING MYOCARDIUM |HIBERNATING MYOCARDIUM (DISORDER)
C1299451|T047|371823002|SNOMEDCT_US|POST-ANGIOPLASTY CORONARY|PATIENT POST ANGIOPLASTY (FINDING)
C1299451|T047|371823002|SNOMEDCT_US|POST CORONARY ANGIOPLASTY |PATIENT POST ANGIOPLASTY (FINDING)
C1299451|T047|371823002|SNOMEDCT_US|POST CORONARY ANGIOPLASTY|PATIENT POST ANGIOPLASTY (FINDING)
C1299451|T047|371823002|SNOMEDCT_US|POST-ANGIOPLASTY|PATIENT POST ANGIOPLASTY (FINDING)
C1299451|T047|371823002|SNOMEDCT_US|PATIENT POST ANGIOPLASTY |PATIENT POST ANGIOPLASTY (FINDING)
C1299451|T047|371823002|SNOMEDCT_US|PATIENT POST ANGIOPLASTY|PATIENT POST ANGIOPLASTY (FINDING)
C3665365|T047|39468009|SNOMEDCT_US|ASCVD (ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE)|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|ARTERIOSCLEROTIC CV DISEASE|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|CARDIOVASCULAR DEGENERATION WITH ARTERIOSCLEROSIS|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|CARDIOVASCULAR SCLEROSIS WITH ARTERIOSCLEROSIS|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|CARDIOVASCULAR ARTERIOSCLEROSIS UNSPECIFIED|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|CARDIOVASCULAR ARTERIOSCLEROSIS|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|CARDIOVASCULAR DISEASE WITH ARTERIOSCLEROSIS|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|CARDIOVASCULAR ARTERIOSCLEROSIS UNSPECIFIED |ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE |ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (ASCVD)|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (ASCVD) |ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE, NOS|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|CARDIOVASCULAR; ARTERIOSCLEROSIS|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|DISEASE (OR DISORDER); ARTERIOSCLEROTIC, CARDIOVASCULAR|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C3665365|T047|39468009|SNOMEDCT_US|ARTERIOSCLEROSIS; CARDIOVASCULAR|ARTERIOSCLEROTIC CARDIOVASCULAR DISEASE (DISORDER)
C2957458|T047||SNOMEDCT_US|NATIVE CORONARY ARTERY STENOSIS
C2957458|T047||SNOMEDCT_US|NATIVE CORONARY ARTERY STENOSIS 
C0340664|T047|234010000|SNOMEDCT_US|CORONARY ARTERY PERFORATION|CORONARY ARTERY PERFORATION (DISORDER)
C0340664|T047|234010000|SNOMEDCT_US|CORONARY ARTERY PERFORATION |CORONARY ARTERY PERFORATION (DISORDER)
C0347699|T047|262941008|SNOMEDCT_US|TRANSECTION OF CORONARY ARTERY|TRANSECTION OF CORONARY ARTERY (DISORDER)
C0347699|T047|262941008|SNOMEDCT_US|TRANSECTION OF CORONARY ARTERY |TRANSECTION OF CORONARY ARTERY (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|GREY AREA DIAGNOSIS BUT UNCOMMON SO DON'T EXPECT TOO MANY FALSE POSITIVES|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CONGENITAL ANOMALY OF CORONARY ARTERY|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY ARTERY ANOMALY|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY ARTERY ANOMALY, CONGENITAL|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY ARTERY ANOMALY NOS|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY ARTERY ABNORMALITY |CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY ARTERY ABNORMALITY|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY ARTERY ANOMALY NOS |CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY ARTERIES--ABNORMALITIES|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|ABNORMALITY OF THE CORONARY ARTERIES|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CONGENITAL CORONARY ARTERY MALFORMATION NOS|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CONGENITAL CORONARY ARTERY MALFORMATION|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CONGENITAL ANOMALY OF CORONARY ARTERY |CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY ARTERY; ANOMALY|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY; ARTERY, ANOMALY|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|DEFORMITY; ARTERY, CORONARY, CONGENITAL|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|A.CORONARIA; ANOMALY|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|ANOMALY; CORONARY ARTERY|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|ARTERY; DEFORMITY, CORONARY, CONGENITAL|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CONGENITAL ANOMALY OF CORONARY ARTERY, NOS|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0158623|T047|204380003|SNOMEDCT_US|CORONARY ARTERY ABNORMALITY [AMBIGUOUS]|CORONARY ARTERY ANOMALY NOS (DISORDER)
C0392158|T047|70390005|SNOMEDCT_US|DISSECTING ANEURYSM OF CORONARY ARTERY|DISSECTING ANEURYSM OF CORONARY ARTERY (DISORDER)
C0392158|T047|70390005|SNOMEDCT_US|DISSECTING CORONARY ARTERY ANEURYSM|DISSECTING ANEURYSM OF CORONARY ARTERY (DISORDER)
C0392158|T047|70390005|SNOMEDCT_US|CORONARY ARTERY ANEURYSM AND DISSECTION|DISSECTING ANEURYSM OF CORONARY ARTERY (DISORDER)
C0392158|T047|70390005|SNOMEDCT_US|ANEURYSM DISSECTING CORONARY ARTERY|DISSECTING ANEURYSM OF CORONARY ARTERY (DISORDER)
C0392158|T047|70390005|SNOMEDCT_US|DISSECTING ANEURYSM OF CORONARY ARTERY |DISSECTING ANEURYSM OF CORONARY ARTERY (DISORDER)
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSMS, CORONARY|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|CORONARY ANEURYSM|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|CORONARY ANEURYSMS|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|CORONARY ARTERY ANEURYSM|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSM OF CORONARY ARTERY |ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSM OF CORONARY ARTERY|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSM CORONARY VESSEL|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|CORONARY ANEURYSM [DISEASE/FINDING]|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSM, CORONARY|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSM;ARTERY;CORONARY|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSMAL LESION OF CORONARY ARTERY|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSMAL LESION OF CORONARY ARTERY |ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSM OF CORONARY VESSELS|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSM OF CORONARY VESSELS |ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|CORONARY; ANEURYSM|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ANEURYSM; CORONARY|ANEURYSMAL LESION OF CORONARY ARTERY
C0010051|T047|50570003|SNOMEDCT_US|ARTERIOVENOUS ANEURYSM OF CORONARY VESSELS|ANEURYSMAL LESION OF CORONARY ARTERY
C0265899|T047|5230009|SNOMEDCT_US|CONGENITAL ABSENCE OF CORONARY ARTERY |CONGENITAL ABSENCE OF CORONARY ARTERY (DISORDER)
C0265899|T047|5230009|SNOMEDCT_US|CONGENITAL ABSENCE OF CORONARY ARTERY|CONGENITAL ABSENCE OF CORONARY ARTERY (DISORDER)
C0265899|T047|5230009|SNOMEDCT_US|ABSENCE; ARTERY, CORONARY|CONGENITAL ABSENCE OF CORONARY ARTERY (DISORDER)
C0265899|T047|5230009|SNOMEDCT_US|ARTERY; ABSENCE, CORONARY|CONGENITAL ABSENCE OF CORONARY ARTERY (DISORDER)
C0265899|T047|5230009|SNOMEDCT_US|CORONARY ARTERY, ABSENCE|CONGENITAL ABSENCE OF CORONARY ARTERY (DISORDER)
C0340648|T047|732230001|SNOMEDCT_US|CORONARY ARTERY DISSECTION|DISSECTION OF CORONARY ARTERY (DISORDER)
C0340648|T047|732230001|SNOMEDCT_US|DISSECTION OF CORONARY ARTERY|DISSECTION OF CORONARY ARTERY (DISORDER)
C0340648|T047|732230001|SNOMEDCT_US|DISSECTION OF CORONARY ARTERY |DISSECTION OF CORONARY ARTERY (DISORDER)
C0340648|T047|732230001|SNOMEDCT_US|DISSECTION COR ARTERY|DISSECTION OF CORONARY ARTERY (DISORDER)
C0340648|T047|732230001|SNOMEDCT_US|CORONARY ARTERY DISSECTION |DISSECTION OF CORONARY ARTERY (DISORDER)
C0343692|T047|240567009|SNOMEDCT_US|SYPHILITIC CORONARY ARTERY DISEASE|SYPHILITIC CORONARY ARTERY DISEASE (DISORDER)
C0343692|T047|240567009|SNOMEDCT_US|SYPHILIS CARDIOVASCULAR CORONARY ARTERY|SYPHILITIC CORONARY ARTERY DISEASE (DISORDER)
C0343692|T047|240567009|SNOMEDCT_US|SYPHILITIC CORONARY ARTERY DISEASE |SYPHILITIC CORONARY ARTERY DISEASE (DISORDER)
C0343692|T047|240567009|SNOMEDCT_US|LATE QUATERNARY SYPHILITIC CORONARY ARTERY DISEASE|SYPHILITIC CORONARY ARTERY DISEASE (DISORDER)
C0343692|T047|240567009|SNOMEDCT_US|SYPHILITIC CORONARY ARTERY DISEASE |SYPHILITIC CORONARY ARTERY DISEASE (DISORDER)
C2939120|T047|11433004|SNOMEDCT_US|CORONARY ARTERY FISTULA|CONGENITAL CORONARY ARTERY FISTULA (DISORDER)
C2939120|T047|11433004|SNOMEDCT_US|CONGENITAL CORONARY ARTERY FISTULA|CONGENITAL CORONARY ARTERY FISTULA (DISORDER)
C2939120|T047|11433004|SNOMEDCT_US|CONGENITAL CORONARY ARTERY FISTULA |CONGENITAL CORONARY ARTERY FISTULA (DISORDER)
C0519097|T047|297160003|SNOMEDCT_US|ANEURYSM OF LEFT VENTRICLE|LEFT VENTRICULAR ANEURYSM (DISORDER)
C0519097|T047|297160003|SNOMEDCT_US|ANEURYSM OF LEFT VENTRICLE |LEFT VENTRICULAR ANEURYSM (DISORDER)
C0519097|T047|297160003|SNOMEDCT_US|LEFT VENTRICULAR ANEURYSM|LEFT VENTRICULAR ANEURYSM (DISORDER)
C0519097|T047|297160003|SNOMEDCT_US|LEFT VENTRICULAR ANEURYSM |LEFT VENTRICULAR ANEURYSM (DISORDER)
C0519097|T047|297160003|SNOMEDCT_US|LV WALL ANEURYSMAL|LEFT VENTRICULAR ANEURYSM (DISORDER)
C0519097|T047|297160003|SNOMEDCT_US|LEFT VENTRICULAR WALL ANEURYSMAL|LEFT VENTRICULAR ANEURYSM (DISORDER)
C0519097|T047|297160003|SNOMEDCT_US|LVA - LEFT VENTRICULAR ANEURYSM|LEFT VENTRICULAR ANEURYSM (DISORDER)
C0340678|T047|234029006|SNOMEDCT_US|CORONARY STEAL SYNDROME|CORONARY STEAL SYNDROME (DISORDER)
C0340678|T047|234029006|SNOMEDCT_US|CORONARY STEAL SYNDROME |CORONARY STEAL SYNDROME (DISORDER)
C0264688|T047|28931004|SNOMEDCT_US|CORONARY (ARTERY) RUPTURE|CORONARY ARTERY RUPTURE (DISORDER)
C0264688|T047|28931004|SNOMEDCT_US|RUPTURE;ARTERY;CORONARY|CORONARY ARTERY RUPTURE (DISORDER)
C0264688|T047|28931004|SNOMEDCT_US|CORONARY ARTERY RUPTURE|CORONARY ARTERY RUPTURE (DISORDER)
C0264688|T047|28931004|SNOMEDCT_US|CORONARY ARTERY RUPTURE |CORONARY ARTERY RUPTURE (DISORDER)
C0264699|T047|62695002|SNOMEDCT_US|ACUTE ANTEROSEPTAL MYOCARDIAL INFARCTION |ACUTE ANTEROSEPTAL MYOCARDIAL INFARCTION (DISORDER)
C0264699|T047|62695002|SNOMEDCT_US|ACUTE ANTEROSEPTAL MYOCARDIAL INFARCTION|ACUTE ANTEROSEPTAL MYOCARDIAL INFARCTION (DISORDER)
C0264699|T047|62695002|SNOMEDCT_US|ACUTE ANTERO SEPTAL MYOCARDIAL INFARCTION|ACUTE ANTEROSEPTAL MYOCARDIAL INFARCTION (DISORDER)
C0264699|T047|62695002|SNOMEDCT_US|ACUTE ANTEROSEPTAL MYOCARDIAL INFARCTION |ACUTE ANTEROSEPTAL MYOCARDIAL INFARCTION (DISORDER)
C0264699|T047|62695002|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION, ANTEROSEPTAL|ACUTE ANTEROSEPTAL MYOCARDIAL INFARCTION (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL |ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|ACUTE INFERIOR WALL MI|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|ACUTE INFERIOR MYOCARDIAL INFARCTION|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF DIAPHRAGMATIC WALL|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL |ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL, NOS|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|INFARCTION, DIAPHRAGMATIC WALL NOS|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION, DIAPHRAGMATIC WALL NOS|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0264700|T047|73795002|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION, INFERIOR WALL NOS|ACUTE MYOCARDIAL INFARCTION OF INFERIOR WALL (DISORDER)
C0345117|T047|253709000|SNOMEDCT_US|ABNORMAL CORONARY ORIFICE |ABNORMAL CORONARY ORIFICE (DISORDER)
C0345117|T047|253709000|SNOMEDCT_US|ABNORMAL CORONARY ORIFICE|ABNORMAL CORONARY ORIFICE (DISORDER)
C0340892|T047|213037002|SNOMEDCT_US|MECHANICAL COMPLICATION OF CORONARY BYPASS|MECHANICAL COMPLICATION OF CORONARY BYPASS (DISORDER)
C0340892|T047|213037002|SNOMEDCT_US|MECHANICAL COMPLICATION OF CORONARY BYPASS |MECHANICAL COMPLICATION OF CORONARY BYPASS (DISORDER)
C0275847|T047|62207008|SNOMEDCT_US|SYPHILITIC OSTIAL CORONARY ARTERY DISEASE|SYPHILITIC OSTIAL CORONARY DISEASE (DISORDER)
C0275847|T047|62207008|SNOMEDCT_US|SYPHILIS CARDIOVASCULAR CORONARY ARTERY OSTIAL|SYPHILITIC OSTIAL CORONARY DISEASE (DISORDER)
C0275847|T047|62207008|SNOMEDCT_US|SYPHILITIC OSTIAL CORONARY ARTERY DISEASE |SYPHILITIC OSTIAL CORONARY DISEASE (DISORDER)
C0275847|T047|62207008|SNOMEDCT_US|SYPHILITIC OSTIAL CORONARY DISEASE|SYPHILITIC OSTIAL CORONARY DISEASE (DISORDER)
C0275847|T047|62207008|SNOMEDCT_US|SYPHILITIC OSTIAL CORONARY DISEASE |SYPHILITIC OSTIAL CORONARY DISEASE (DISORDER)
C0221359|T047|75398000|SNOMEDCT_US|ANOMALOUS ORIGIN OF CORONARY ARTERY |ANOMALOUS ORIGIN OF CORONARY ARTERY (DISORDER)
C0221359|T047|75398000|SNOMEDCT_US|ANOMALOUS ORIGIN OF CORONARY ARTERY|ANOMALOUS ORIGIN OF CORONARY ARTERY (DISORDER)
C0221359|T047|75398000|SNOMEDCT_US|CONGENITAL ANOMALY OF CORONARY ARTERY OF ANOMALOUS ORIGIN|ANOMALOUS ORIGIN OF CORONARY ARTERY (DISORDER)
C0221359|T047|75398000|SNOMEDCT_US|ANOMALOUS CORONARY ARTERY ORIGIN|ANOMALOUS ORIGIN OF CORONARY ARTERY (DISORDER)
C0221359|T047|75398000|SNOMEDCT_US|ANOMALOUS ORIGIN OF CORONARY ARTERY |ANOMALOUS ORIGIN OF CORONARY ARTERY (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY OCCLUSION|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY ARTERY OCCLUSION|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|OCCLUSIONS, CORONARY|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY OCCLUSIONS|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|OCCLUSION, CORONARY|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY (ARTERY) OCCLUSION|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY OCCLUSION [DISEASE/FINDING]|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|OCCLUSION;CORONARY|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY ARTERY OCCLUSION |CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|OCCLUSION CORONARY|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|OCCLUSION CORONARY ARTERY|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY ARTERY OCCLUDED|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY OCCLUSION |CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY OCCLUSION, NOS|CORONARY OCCLUSION (DISORDER)
C0151814|T047|63739005|SNOMEDCT_US|CORONARY OCCLUSION NOS|CORONARY OCCLUSION (DISORDER)
C0340297|T047|79009004|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF SEPTAL WALL |ACUTE MYOCARDIAL INFARCTION OF SEPTUM (DISORDER)
C0340297|T047|79009004|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF SEPTAL WALL|ACUTE MYOCARDIAL INFARCTION OF SEPTUM (DISORDER)
C0340297|T047|79009004|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF SEPTUM|ACUTE MYOCARDIAL INFARCTION OF SEPTUM (DISORDER)
C0340297|T047|79009004|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF SEPTUM ALONE|ACUTE MYOCARDIAL INFARCTION OF SEPTUM (DISORDER)
C0340297|T047|79009004|SNOMEDCT_US|ACUTE SEPTAL INFARCTION|ACUTE MYOCARDIAL INFARCTION OF SEPTUM (DISORDER)
C0340297|T047|79009004|SNOMEDCT_US|ACUTE MYOCARDIAL INFARCTION OF SEPTUM |ACUTE MYOCARDIAL INFARCTION OF SEPTUM (DISORDER)
C0340297|T047|79009004|SNOMEDCT_US|INFARCTION OF SEPTUM ALONE|ACUTE MYOCARDIAL INFARCTION OF SEPTUM (DISORDER)
C3695002|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE IN TRANSPLANTED HEART 
C3695002|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE IN TRANSPLANTED HEART
C3697310|T047|699257002|SNOMEDCT_US|INCREASE IN VELOCITY OF CORONARY ARTERY OF FETUS|INCREASE IN VELOCITY OF CORONARY ARTERY OF FETUS (DISORDER)
C3697310|T047|699257002|SNOMEDCT_US|INCREASE IN VELOCITY OF CORONARY ARTERY OF FETUS |INCREASE IN VELOCITY OF CORONARY ARTERY OF FETUS (DISORDER)
C1834751|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE, DEVELOPMENT OF, IN HIV
C1859728|T047||SNOMEDCT_US|CORONARY SCLEROSIS, MEDIAL, OF INFANCY
C2063729|T047||SNOMEDCT_US|MULTIPLE CORONARY ANEURYSMS
C2063729|T047||SNOMEDCT_US|MULTIPLE CORONARY ANEURYSMS 
C0027051|T047|22298006|SNOMEDCT_US|INFARCTIONS, MYOCARDIAL|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTION|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTIONS|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCTS, MYOCARDIAL|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTS|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCT, MYOCARDIAL|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCTION, MYOCARDIAL|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MI|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTION (MI)|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|HEART ATTACK|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|CARDIAC INFARCTION|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTION [DISEASE/FINDING]|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCT|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCTION;HEART|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCTION;MYOCARDIAL|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|ATTACK - HEART|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MI - MYOCARDIAL INFARCTION|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTION |MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|CARDIAC INFARCT|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTION |MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|-- HEART ATTACK|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|CARDIOVASCULAR STROKES|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|STROKE, CARDIOVASCULAR|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|STROKES, CARDIOVASCULAR|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|CARDIOVASCULAR STROKE|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MI, MYOCARDIAL INFARCTION|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTION, (MI)|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCTION (MI), MYOCARDIAL|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|HEART ATTACKS|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|ATTACK CORONARY|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|ATTACK HEART (NOS)|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCT MYOCARDIAL|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|CARDIO/PULM: MYOCARDIAL INFARCTION|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCTION OF HEART|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|CARDIAC; INFARCTION|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCTION; MYOCARDIAL|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|CARDIAC INFARCTION, NOS|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|HEART ATTACK, NOS|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCTION OF HEART, NOS|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTION, NOS|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|INFARCTIONS (MYOCARDIAL)|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|MYOCARDIAL INFARCTION NOS|MYOCARDIAL INFARCTION (DISORDER)
C0027051|T047|22298006|SNOMEDCT_US|HEART INFARCTION|MYOCARDIAL INFARCTION (DISORDER)
C3165030|T047|448478000|SNOMEDCT_US|SYSTEMIC TO PULMONARY COLLATERAL FROM CORONARY ARTERY|SYSTEMIC TO PULMONARY COLLATERAL FROM CORONARY ARTERY
C3165030|T047|448478000|SNOMEDCT_US|SYSTEMIC TO PULMONARY COLLATERAL ARTERY FROM CORONARY ARTERY |SYSTEMIC TO PULMONARY COLLATERAL FROM CORONARY ARTERY
C3165030|T047|448478000|SNOMEDCT_US|SYSTEMIC TO PULMONARY COLLATERAL FROM CORONARY ARTERY |SYSTEMIC TO PULMONARY COLLATERAL FROM CORONARY ARTERY
C3165030|T047|448478000|SNOMEDCT_US|SYSTEMIC TO PULMONARY COLLATERAL ARTERY FROM CORONARY ARTERY|SYSTEMIC TO PULMONARY COLLATERAL FROM CORONARY ARTERY
C4020725|T047||SNOMEDCT_US|NON-OCCLUSIVE CORONARY ARTERY DISEASE
C4020725|T047||SNOMEDCT_US|NONOCCLUSIVE CORONARY ARTERY DISEASE
C4020725|T047||SNOMEDCT_US|NON-OCCLUSIVE CORONARY ARTERY STENOSIS
C2676505|T047||SNOMEDCT_US|POST-ANGIOPLASTY CORONARY ARTERY RESTENOSIS
C4047786|T047|19830001000004106|SNOMEDCT_US|THROMBOSIS OF LEFT CIRCUMFLEX ARTERY|THROMBOSIS OF LEFT CIRCUMFLEX ARTERY (DISORDER)
C4047786|T047|19830001000004106|SNOMEDCT_US|THROMBOSIS OF LEFT CIRCUMFLEX ARTERY |THROMBOSIS OF LEFT CIRCUMFLEX ARTERY (DISORDER)
C4075502|T047|714180007|SNOMEDCT_US|ABNORMAL OSTIUM OF CORONARY ARTERY|ABNORMAL OSTIUM OF CORONARY ARTERY (DISORDER)
C4075502|T047|714180007|SNOMEDCT_US|ABNORMAL OSTIUM OF CORONARY ARTERY |ABNORMAL OSTIUM OF CORONARY ARTERY (DISORDER)
C1299363|T047|371894001|SNOMEDCT_US|BIFURCATION LESION OF CORONARY ARTERY|BIFURCATION LESION OF CORONARY ARTERY (DISORDER)
C1299363|T047|371894001|SNOMEDCT_US|BIFURCATION LESION OF CORONARY ARTERY |BIFURCATION LESION OF CORONARY ARTERY (DISORDER)
C1299363|T047|371894001|SNOMEDCT_US|BIFURCATION LESION OF CORONARY ARTERY |BIFURCATION LESION OF CORONARY ARTERY (DISORDER)
C0265898|T047|373093003|SNOMEDCT_US|CORONARY ARTERY FISTULA|CORONARY ARTERY FISTULA (DISORDER)
C0265898|T047|373093003|SNOMEDCT_US|CORONARY ARTERY FISTULA |CORONARY ARTERY FISTULA (DISORDER)
