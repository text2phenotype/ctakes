C0982429|T121|1313771|RXNORM|TEA-DODECYLBENZENESULFONATE|TRIETHANOLAMINE DODECYLBENZENESULFONATE
C0067870|T109|1313770|RXNORM|N-BUTYL ACRYLATE|N-BUTYL ACRYLATE
C3257527|T121|1426332|RXNORM|MANGO EXTRACT|MANGIFERA INDICA (MANGO) FRUIT EXTRACT
C0936105|T121|282427|RXNORM|AMITRIPTYLINE / PERPHENAZINE|AMITRIPTYLINE / PERPHENAZINE
C3541952|T109|1426336|RXNORM|PHENOXYACETATE|PHENOXYACETATE
C0220874|T109|1426331|RXNORM|MALEATE|MALEATE
C0771904|T121|1426339|RXNORM|POLIFEPROSAN 20|POLIFEPROSAN 20
C3256060|T121|1307836|RXNORM|MELISSA OFFICINALIS LEAF EXTRACT|MELISSA OFFICINALIS LEAF EXTRACT
C2929085|T121|1008178|RXNORM|TOLNAFTATE / TRICLOSAN|TOLNAFTATE / TRICLOSAN
C2929086|T121|1008179|RXNORM|CHLORZOXAZONE / FLUFENAMIC ACID|CHLORZOXAZONE / FLUFENAMIC ACID
C3555482|T121|1420957|RXNORM|ALOE ANDONGENSIS LEAF EXTRACT|ALOE ANDONGENSIS LEAF EXTRACT
C2929079|T121|1008172|RXNORM|CODEINE / PHENYLTOLOXAMINE|CODEINE / PHENYLTOLOXAMINE
C2929080|T121|1008173|RXNORM|ANISE OIL / THYME PREPARATION|ANISE OIL / THYME PREPARATION
C2929077|T121|1008170|RXNORM|IBUPROFEN / NIACIN|IBUPROFEN / NIACIN
C2929078|T121|1008171|RXNORM|LAURETH-9 / ZINC OXIDE|POLIDOCANOL / ZINC OXIDE
C2929083|T121|1008176|RXNORM|ERGOTAMINE / PROPYPHENAZONE|ERGOTAMINE / PROPYPHENAZONE
C2929084|T121|1008177|RXNORM|COUMARIN / TROXERUTIN|COUMARIN / TROXERUTIN
C2929081|T121|1008174|RXNORM|ADRENAL CORTEX EXTRACT / ROSEMARY OIL|ADRENAL CORTEX EXTRACT / ROSEMARY OIL
C2929082|T121|1008175|RXNORM|BUTALAMINE / PAPAVERINE|BUTALAMINE / PAPAVERINE
C3256865|T121|1307653|RXNORM|PRUNUS MUME FLOWER EXTRACT|PRUNUS MUME FLOWER EXTRACT
C3256213|T121|1307655|RXNORM|CURCUMA LONGA LEAF EXTRACT|CURCUMA LONGA LEAF EXTRACT
C3255687|T121|1307659|RXNORM|LIGUSTICUM TENUISSIMUM ROOT EXTRACT|LIGUSTICUM TENUISSIMUM ROOT EXTRACT
C3256567|T121|1307658|RXNORM|THYMUS VULGARIS LEAF EXTRACT|THYMUS VULGARIS LEAF EXTRACT
C3255623|T130|1310562|RXNORM|FD &C YELLOW #6 ALUMINUM LAKE|FD &C YELLOW #6 ALUMINUM LAKE
C2183732|T121|813715|RXNORM|ACETAMINOPHEN / DIPHENHYDRAMINE / PHENYLPROPANOLAMINE|ACETAMINOPHEN / DIPHENHYDRAMINE / PHENYLPROPANOLAMINE
C0060435|T121|25060|RXNORM|FLAVODIC ACID|FLAVODIC ACID
C1720359|T121|645244|RXNORM|DESOXIMETASONE / SALICYLIC ACID|DESOXIMETASONE / SALICYLIC ACID
C1720293|T121|645247|RXNORM|DEXTROMETHORPHAN / MENTHOL|DEXTROMETHORPHAN / MENTHOL
C3256712|T109|1426389|RXNORM|OLDENLANDIA DIFFUSA EXTRACT|OLDENLANDIA DIFFUSA EXTRACT
C0770355|T121|235389|RXNORM|MESTRANOL / NORETHYNODREL|MESTRANOL / NORETHYNODREL
C1719967|T121|645246|RXNORM|DEXTROMETHORPHAN / DIPHENHYDRAMINE|DEXTROMETHORPHAN / DIPHENHYDRAMINE
C2740965|T129|900045|RXNORM|OREGON ASH POLLEN EXTRACT|FRAXINUS LATIFOLIA POLLEN EXTRACT
C1828708|T121|1363571|RXNORM|1,2-OCTANEDIOL|1,2-OCTANEDIOL
C3855140|T109|1547472|RXNORM|CORYDALIS BUNGEANA WHOLE EXTRACT|CORYDALIS BUNGEANA WHOLE EXTRACT
C2350383|T121|816249|RXNORM|PENTASTARCH|PENTASTARCH
C3643373|T109|1421429|RXNORM|ADANSONIA DIGITATA SEED OIL|ADANSONIA DIGITATA SEED OIL
C3645051|T109|1426388|RXNORM|MESYLATE|MESYLATE
C1875213|T121|689436|RXNORM|GLYCERIN / PROPYLENE GLYCOL|GLYCERIN / PROPYLENE GLYCOL
C2727890|T129|350173|RXNORM|HOUSE FLY ALLERGENIC EXTRACT|MUSCA DOMESTICA ALLERGENIC EXTRACT
C1875214|T121|689438|RXNORM|GLYCERIN / SALICYLIC ACID|GLYCERIN / SALICYLIC ACID
C2356045|T121|802646|RXNORM|METFORMIN / REPAGLINIDE|METFORMIN / REPAGLINIDE
C2701991|T109|853112|RXNORM|MOMORDICAE|MOMORDICAE
C0060692|T125|25284|RXNORM|FOSFESTROL|FOSFESTROL
C2057476|T121|822000|RXNORM|CARISOPRODOL / DEXAMETHASONE / TENOXICAM|CARISOPRODOL / DEXAMETHASONE / TENOXICAM
C0074750|T197|36702|RXNORM|SODIUM PERBORATE|SODIUM PERBORATE
C0001268|T195|270|RXNORM|SPECTINOMYCIN|SPECTINOMYCIN
C3497613|T121|1314266|RXNORM|ARACHIDYL BEHENATE|ARACHIDYL BEHENATE
C0001275|T121|272|RXNORM|ACTIVATED CHARCOAL|MEDICINAL CHARCOAL
C0001275|T121|272|RXNORM|ACTIVATED CHARCOAL|MEDICINAL CHARCOAL
C0074748|T197|36700|RXNORM|SODIUM NITRATE|SODIUM NITRATE
C0915142|T121|279950|RXNORM|PARECOXIB|PARECOXIB
C3555481|T121|1420958|RXNORM|ARALIA CORDATA ROOT EXTRACT|ARALIA CORDATA ROOT EXTRACT
C3555480|T121|1420959|RXNORM|CNIDIUM OFFICINALE WHOLE EXTRACT|CNIDIUM OFFICINALE WHOLE EXTRACT
C0026917|T007|1320629|RXNORM|MYCOBACTERIUM BOVIS|MYCOBACTERIUM BOVIS
C0057362|T121|22483|RXNORM|DEMEGESTONE|DEMEGESTONE
C0733397|T121|227239|RXNORM|MASOPROCOL|MASOPROCOL
C0002728|T109|1368128|RXNORM|AMYLOPECTIN|AMYLOPECTIN
C0298499|T121|1368129|RXNORM|APAFLURANE|APAFLURANE
C3818809|T121|1489919|RXNORM|PPG-1-PEG-9 LAURYL GLYCOL ETHER|PPG-1-PEG-9 LAURYL GLYCOL ETHER
C2353443|T109|1489918|RXNORM|METAFLUMIZONE|METAFLUMIZONE
C0318115|T007|1489917|RXNORM|STAPHYLOCOCCUS SIMULANS|STAPHYLOCOCCUS SIMULANS
C0318114|T007|1489916|RXNORM|STAPHYLOCOCCUS HAEMOLYTICUS|STAPHYLOCOCCUS HAEMOLYTICUS
C0038174|T007|1489915|RXNORM|STAPHYLOCOCCUS EPIDERMIDIS|STAPHYLOCOCCUS EPIDERMIDIS
C3817397|T121|1489914|RXNORM|ELOSULFASE ALFA|ELOSULFASE ALFA
C0000378|T123|1489913|RXNORM|DROXIDOPA|DROXIDOPA
C3485673|T121|1368127|RXNORM|AMNIOTIC FLUID (BOVINE)|AMNIOTIC FLUID (BOVINE)
C0050587|T131|1368125|RXNORM|ACRYLAMIDE|ACRYLAMIDE
C2183093|T121|819018|RXNORM|CARBOCYSTEINE / DEXTROMETHORPHAN|CARBOCYSTEINE / DEXTROMETHORPHAN
C0035167|T121|9259|RXNORM|RESCINNAMINE|RESCINNAMINE
C0036078|T121|9524|RXNORM|SULFASALAZINE|SULFASALAZINE
C0036079|T121|9525|RXNORM|SALICYLIC ACID|SALICYLIC ACID
C0036079|T121|9525|RXNORM|SALICYLIC ACID|SALICYLIC ACID
C0036079|T121|9525|RXNORM|SALICYLIC ACID|SALICYLIC ACID
C0771169|T121|235961|RXNORM|FEDRILATE|FEDRILATE
C1654081|T122|1311163|RXNORM|CARBOMER 1342|CARBOMER COPOLYMER TYPE B (ALLYL PENTAERYTHRITOL CROSSLINKED)
C0041249|T123|10898|RXNORM|TRYPTOPHAN|TRYPTOPHAN
C3535835|T121|1370659|RXNORM|DODECYLBENZENESULFONATE|DODECYLBENZENESULFONATE
C3535819|T121|1370658|RXNORM|COCOATE|COCOATE
C0105205|T121|46795|RXNORM|BARBEXACLONE|BARBEXACLONE
C3535838|T121|1370655|RXNORM|C14 OLEFIN SULFONATE|C14 OLEFIN SULFONATE
C3535839|T121|1370654|RXNORM|C12-15 PARETH-15 SULFONATE|C12-15 PARETH-15 SULFONATE
C3535836|T197|1370657|RXNORM|COCO-SULFATE|COCO-SULFATE
C3535837|T121|1370656|RXNORM|CASEINATE|CASEINATE
C3535842|T121|1370651|RXNORM|OLEAMIDO MIPA-SULFOSUCCINATE|OLEAMIDO MIPA-SULFOSUCCINATE
C3535843|T121|1370650|RXNORM|OLEAMIDO MEA-SULFOSUCCINATE|OLEAMIDO MEA-SULFOSUCCINATE
C3535840|T121|1370653|RXNORM|C12-14 OLEFIN SULFONATE|C12-14 OLEFIN SULFONATE
C3535841|T121|1370652|RXNORM|C12 OLEFIN SULFONATE|C12 OLEFIN SULFONATE
C1445763|T121|466529|RXNORM|CHLORPHENIRAMINE / GUAIFENESIN / HYDROCODONE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / GUAIFENESIN / HYDROCODONE / PSEUDOEPHEDRINE
C2114805|T121|816721|RXNORM|PHOLCODINE / PROMETHAZINE|PHOLCODINE / PROMETHAZINE
C2047218|T121|816726|RXNORM|INSULIN LISPRO / INSULIN, PROTAMINE LISPRO, HUMAN|INSULIN LISPRO / INSULIN, PROTAMINE LISPRO, HUMAN
C2741499|T129|901317|RXNORM|SPINACH ALLERGENIC EXTRACT|SPINACIA OLERACEA ALLERGENIC EXTRACT
C1445756|T121|466522|RXNORM|DIPHENHYDRAMINE / ZINC ACETATE|DIPHENHYDRAMINE / ZINC ACETATE
C3696421|T121|1484756|RXNORM|NOVOBIOCIN / PENICILLIN G|NOVOBIOCIN / PENICILLIN G
C1445758|T121|466524|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / DOXYLAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / DEXTROMETHORPHAN / DOXYLAMINE / PSEUDOEPHEDRINE
C3832607|T109|1539194|RXNORM|SCROPHULARIA BUEGERIANA ROOT EXTRACT|SCROPHULARIA BUEGERIANA ROOT EXTRACT
C3486792|T121|1311410|RXNORM|MAITAKE EXTRACT|MAITAKE EXTRACT
C2079437|T121|821005|RXNORM|ETHAMBUTOL / ISONIAZID|ETHAMBUTOL / ISONIAZID
C3486538|T121|1306291|RXNORM|COBICISTAT / ELVITEGRAVIR / EMTRICITABINE / TENOFOVIR DISOPROXIL|COBICISTAT / ELVITEGRAVIR / EMTRICITABINE / TENOFOVIR DISOPROXIL
C0525227|T121|134615|RXNORM|BRIMONIDINE|BRIMONIDINE
C0525227|T121|134615|RXNORM|BRIMONIDINE|BRIMONIDINE
C3855209|T121|1547556|RXNORM|SPHAERANTHUS INDICUS FLOWERING TOP EXTRACT|SPHAERANTHUS INDICUS FLOWERING TOP EXTRACT
C1445182|T130|465953|RXNORM|CAT DANDER EXTRACT|FELIS CATUS DANDER EXTRACT
C3855208|T121|1547555|RXNORM|CYTISUS SCOPARIUS FLOWER EXTRACT|CYTISUS SCOPARIUS FLOWER EXTRACT
C3255208|T126|1431738|RXNORM|ASPARAGINASE ERWINIA CHRYSANTHEMI|ASPARAGINASE ERWINIA CHRYSANTHEMI
C3474129|T121|1314262|RXNORM|ACHYRANTHES JAPONICA WHOLE EXTRACT|ACHYRANTHES JAPONICA WHOLE EXTRACT
C1533699|T129|1294580|RXNORM|GEMTUZUMAB OZOGAMICIN|GEMTUZUMAB OZOGAMICIN
C0962432|T121|1547558|RXNORM|THREONATE|THREONATE
C3855211|T109|1547559|RXNORM|GENTIANA MANSHURICA WHOLE EXTRACT|GENTIANA MANSHURICA WHOLE EXTRACT
C1874613|T121|690647|RXNORM|BROMPHENIRAMINE / CODEINE / PHENYLEPHRINE|BROMPHENIRAMINE / CODEINE / PHENYLEPHRINE
C1719893|T121|645045|RXNORM|CALAMINE / ZINC OXIDE|CALAMINE / ZINC OXIDE
C0178474|T121|618257|RXNORM|AMINOBUTYRATE|AMINOBUTYRATE
C1874609|T121|690642|RXNORM|BRILLIANT GREEN / GENTIAN VIOLET / PROFLAVINE|BRILLIANT GREEN / GENTIAN VIOLET / PROFLAVINE
C0076107|T121|37798|RXNORM|TERAZOSIN|TERAZOSIN
C1433702|T122|1431309|RXNORM|POLYGLYCERYL-6-DIOLEATE|POLYGLYCERYL-6-DIOLEATE
C0086761|T130|42837|RXNORM|P-AMINOHIPPURATE|P-AMINOHIPPURATE
C3538462|T121|1372879|RXNORM|BRILLIANT GREEN / COD LIVER OIL / GENTIAN VIOLET|BRILLIANT GREEN / COD LIVER OIL / GENTIAN VIOLET
C1640726|T121|645048|RXNORM|CALCIUM CARBONATE / SIMETHICONE|CALCIUM CARBONATE / SIMETHICONE
C0012547|T129|3510|RXNORM|DIPHTHERIA ANTITOXIN|DIPHTHERIA IMMUNOGLOBULIN
C1565316|T121|596205|RXNORM|RAMELTEON|RAMELTEON
C3256781|T121|1314302|RXNORM|LARIX SIBIRICA WOOD EXTRACT|LARIX SIBIRICA WOOD EXTRACT
C0009279|T121|2685|RXNORM|COLESTIPOL|COLESTIPOL
C1876049|T121|692863|RXNORM|IODINE POVACRYLEX|IODINE POVACRYLEX
C3486071|T121|1326501|RXNORM|CARBO ANIMALIS PREPARATION|CARBO ANIMALIS PREPARATION
C0009262|T121|2683|RXNORM|COLCHICINE|COLCHICINE
C2929669|T121|1008770|RXNORM|BENDROFLUMETHIAZIDE / PAPAVERINE / RAUWOLFIA PREPARATION|BENDROFLUMETHIAZIDE / PAPAVERINE / RAUWOLFIA PREPARATION
C2929670|T121|1008771|RXNORM|ALANINE / ARGININE / CALCIUM ACETATE / CYSTEINE / GLYCERIN / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM ACETATE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM ACETATE / SODIUM CHLORIDE|ALANINE / ARGININE / CALCIUM ACETATE / CYSTEINE / GLYCERIN / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM ACETATE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / VALINE
C2929671|T121|1008772|RXNORM|BOX ELDER MAPLE POLLEN EXTRACT / HARD MAPLE POLLEN EXTRACT / RED MAPLE POLLEN EXTRACT|BOX ELDER MAPLE POLLEN EXTRACT / HARD MAPLE POLLEN EXTRACT / RED MAPLE POLLEN EXTRACT
C2929672|T121|1008773|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / FOLIC ACID / ST. JOHN'S WORT EXTRACT|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / FOLIC ACID / ST. JOHN'S WORT EXTRACT
C2929673|T121|1008774|RXNORM|CITICOLINE / ERGOLOID MESYLATES, USP|CITICOLINE / ERGOLOID MESYLATES, USP
C2929674|T121|1008775|RXNORM|EVENING PRIMROSE OIL / GAMMA LINOLEIC ACID|EVENING PRIMROSE OIL / GAMMA LINOLEIC ACID
C2929675|T121|1008776|RXNORM|BELLADONNA EXTRACT, USP / CHLORPHENIRAMINE / EPHEDRINE / PHENOBARBITAL|BELLADONNA EXTRACT, USP / CHLORPHENIRAMINE / EPHEDRINE / PHENOBARBITAL
C0242531|T121|71535|RXNORM|VECURONIUM|VECURONIUM
C2929678|T121|1008779|RXNORM|GLYCERIN / LACTATE / PETROLATUM|GLYCERIN / LACTATE / PETROLATUM
C0012201|T121|3389|RXNORM|DIETHYLPROPION|DIETHYLPROPION
C0000608|T121|99|RXNORM|6-AMINOCAPROIC ACID|6-AMINOCAPROIC ACID
C2075008|T121|818150|RXNORM|ALGINIC ACID / CIMETIDINE|ALGINIC ACID / CIMETIDINE
C0001134|T197|236|RXNORM|FRUIT EXTRACTS|ACIDULATED PHOSPHATE FLUORIDE
C0000578|T123|94|RXNORM|5-HYDROXYTRYPTOPHAN|5-HYDROXYTRYPTOPHAN
C3178623|T121|1368878|RXNORM|ISOCETETH 20|ISOCETETH 20
C3486826|T197|1358876|RXNORM|SILVER CATION|SILVER CATION
C2928911|T121|1007999|RXNORM|CARBOCYSTEINE / PROMETHAZINE|CARBOCYSTEINE / PROMETHAZINE
C2928910|T121|1007998|RXNORM|CARBOCYSTEINE / OXOLAMINE|CARBOCYSTEINE / OXOLAMINE
C0019351|T005|1318479|RXNORM|HUMAN HERPESVIRUS 2|HUMAN HERPESVIRUS 2
C2928907|T121|1007995|RXNORM|CALCIUM CHLORIDE / GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE|CALCIUM CHLORIDE / GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE
C2928906|T121|1007994|RXNORM|GLUCOSE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE|GLUCOSE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE
C2928909|T121|1007997|RXNORM|BIOTIN / CHROMIUM PICOLINATE|BIOTIN / CHROMIUM PICOLINATE
C2928908|T121|1007996|RXNORM|FLORFENICOL / FLUNIXIN|FLORFENICOL / FLUNIXIN
C2928903|T121|1007991|RXNORM|BIOTIN / CYSTEINE / SILICON DIOXIDE|BIOTIN / CYSTEINE / SILICON DIOXIDE
C2928902|T121|1007990|RXNORM|ALLANTOIN / CAMPHOR / MENTHOL / PHENOL|ALLANTOIN / CAMPHOR / MENTHOL / PHENOL
C2928905|T121|1007993|RXNORM|ASCORBIC ACID / BUTCHER'S BROOM PREPARATION / HESPERIDIN|ASCORBIC ACID / BUTCHER'S BROOM PREPARATION / HESPERIDIN
C2928904|T121|1007992|RXNORM|BENZOCAINE / ETHANOL / METHYLBENZETHONIUM|BENZOCAINE / ETHANOL / METHYLBENZETHONIUM
C3488182|T129|1310455|RXNORM|AGKISTRODON CONTORTRIX VENOM|COPPERHEAD VENOM
C3488214|T131|1310457|RXNORM|HELODERMA HORRIDUM VENOM|HELODERMA HORRIDUM VENOM
C3486775|T121|1310108|RXNORM|POPULUS TREMULOIDES LEAF EXTRACT|POPULUS TREMULOIDES LEAF EXTRACT
C3486308|T121|1310107|RXNORM|PINUS DENSIFLORA BARK EXTRACT|PINUS DENSIFLORA BARK EXTRACT
C3486774|T121|1310106|RXNORM|POPULUS TREMULOIDES BARK EXTRACT|POPULUS TREMULOIDES BARK EXTRACT
C3486305|T121|1310105|RXNORM|CITRUS BERGAMIA LEAF EXTRACT|CITRUS BERGAMIA LEAF EXTRACT
C3486069|T121|1310103|RXNORM|TRILLIUM ERECTUM ROOT EXTRACT|TRILLIUM ERECTUM ROOT EXTRACT
C3485067|T121|1310102|RXNORM|AGROSTIS GIGANTEA TOP EXTRACT|AGROSTIS GIGANTEA TOP EXTRACT
C3486066|T121|1310101|RXNORM|PAEONIA OFFICINALIS ROOT EXTRACT|PAEONIA OFFICINALIS ROOT EXTRACT
C3486773|T121|1310100|RXNORM|POPULUS TREMULA FLOWERING TOP EXTRACT|POPULUS TREMULA FLOWERING TOP EXTRACT
C0939804|T121|285155|RXNORM|KELP PREPARATION|KELP PREPARATION
C0939806|T121|285157|RXNORM|MATRICARIA RECUTITA EXTRACT|MATRICARIA CHAMOMILLA EXTRACT
C0317625|T007|285156|RXNORM|LACTOBACILLUS REUTERI|LACTOBACILLUS REUTERI
C3497966|T121|1311508|RXNORM|ORIGANUM VULGARE SUBSP. HIRTUM FLOWER EXTRACT|ORIGANUM VULGARE SUBSP. HIRTUM FLOWER EXTRACT
C3488923|T121|1311509|RXNORM|PAULLINIA CUPANA SEED EXTRACT|PAULLINIA CUPANA SEED EXTRACT
C0939802|T121|285153|RXNORM|GELSEMIUM SEMPERVIRENS PREPARATION|GELSEMIUM SEMPERVIRENS PREPARATION
C0939801|T109|285152|RXNORM|EUPATORIUM PERFOLIATUM PREPARATION|EUPATORIUM PERFOLIATUM PREPARATION
C0002367|T196|1311504|RXNORM|ALUMINUM|ALUMINUM
C2697513|T121|1311505|RXNORM|GLYCYRRHIZIN, AMMONIATED|GLYCYRRHIZIN, AMMONIATED
C0017986|T121|1311506|RXNORM|GLYCYRRHETINIC ACID|GLYCYRRHETINIC ACID
C0094910|T121|1311507|RXNORM|ENZACAMENE|ENZACAMENE
C1337345|T121|1311500|RXNORM|MEBROFENIN|MEBROFENIN
C3257441|T121|1311501|RXNORM|ROSA CANINA FRUIT EXTRACT|ROSA CANINA FRUIT EXTRACT
C2928117|T121|1007195|RXNORM|MYRTOL / OXYTETRACYCLINE|MYRTOL / OXYTETRACYCLINE
C2928116|T121|1007194|RXNORM|ALLANTOIN / CLIOQUINOL / PHENOL|ALLANTOIN / CLIOQUINOL / PHENOL
C2928119|T121|1007197|RXNORM|HYDROCORTISONE / METRONIDAZOLE / MICONAZOLE|HYDROCORTISONE / METRONIDAZOLE / MICONAZOLE
C0717449|T121|214257|RXNORM|ASPIRIN / PENTAZOCINE|ASPIRIN / PENTAZOCINE
C2928113|T121|1007191|RXNORM|PASSION FLOWER EXTRACT / VALERIAN ROOT EXTRACT|PASSION FLOWER EXTRACT / VALERIAN ROOT EXTRACT
C2928112|T121|1007190|RXNORM|CHOLINE / INOSITOL / LYSINE / METHIONINE / VITAMIN B 12|CHOLINE / INOSITOL / LYSINE / METHIONINE / VITAMIN B 12
C3665259|T121|1435633|RXNORM|DYCLONINE / PHENOL|DYCLONINE / PHENOL
C2928121|T121|1007199|RXNORM|HALCINONIDE / NEOMYCIN|HALCINONIDE / NEOMYCIN
C2928120|T121|1007198|RXNORM|DIPYRONE / PROPINOX|DIPYRONE / PROPINOX
C3665262|T121|1435637|RXNORM|ZANTHOXYLUM PIPERITUM FRUIT RIND EXTRACT|ZANTHOXYLUM PIPERITUM FRUIT RIND EXTRACT
C3503281|T121|1370574|RXNORM|VALERATE|VALERATE
C0114771|T121|49247|RXNORM|DOFETILIDE|DOFETILIDE
C2364549|T129|805549|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007 (H1N1) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007 (H1N1) STRAIN
C2701140|T129|851894|RXNORM|IODINE BUSH POLLEN EXTRACT|ALLENROLFEA OCCIDENTALIS POLLEN EXTRACT
C0206461|T121|67109|RXNORM|DALTEPARIN|DALTEPARIN
C0206460|T121|67108|RXNORM|ENOXAPARIN|ENOXAPARIN
C0982042|T121|314521|RXNORM|BENZOXIQUINE|BENZOXIQUINE
C0981927|T129|314411|RXNORM|MONILIA SITOPHILA EXTRACT|CHRYSONILIA SITOPHILA EXTRACT
C2194307|T121|816825|RXNORM|CAFFEINE / DIPYRONE / ERGOTAMINE|CAFFEINE / DIPYRONE / ERGOTAMINE
C1273169|T121|388499|RXNORM|INDAPAMIDE / PERINDOPRIL|INDAPAMIDE / PERINDOPRIL
C0719741|T121|216449|RXNORM|DENATURED ETHANOL|DENATURED ETHANOL
C2216439|T121|815062|RXNORM|MAGNESIUM ASPARTATE / POTASSIUM ASPARTATE|MAGNESIUM ASPARTATE / POTASSIUM ASPARTATE
C0068746|T121|31786|RXNORM|NIFURZIDE|NIFURZIDE
C2928293|T121|1007371|RXNORM|CHROMIUM PICOLINATE / GRAPEFRUIT EXTRACT / LIPOTROPIC AGENTS|CHROMIUM PICOLINATE / GRAPEFRUIT EXTRACT / LIPOTROPIC AGENTS
C2928292|T121|1007370|RXNORM|COENZYME Q10 / GARLIC PREPARATION / HAWTHORN PREPARATION / VITAMIN E|COENZYME Q10 / GARLIC PREPARATION / HAWTHORN PREPARATION / VITAMIN E
C2928295|T121|1007373|RXNORM|IBUPROFEN / VITAMIN B 12|IBUPROFEN / VITAMIN B 12
C2928294|T121|1007372|RXNORM|POTASSIUM GLUCONATE / VITAMIN B6|POTASSIUM GLUCONATE / VITAMIN B6
C2928297|T121|1007375|RXNORM|MENTHOL / METHYL SALICYLATE / METHYLNICOTINATE|MENTHOL / METHYL SALICYLATE / METHYLNICOTINATE
C2928296|T121|1007374|RXNORM|HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / PHENYL SALICYLATE / SODIUM PHOSPHATE, MONOBASIC|HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / PHENYL SALICYLATE / SODIUM PHOSPHATE, MONOBASIC
C2928299|T121|1007377|RXNORM|ECHINACEA ROOT EXTRACT / ECHINACEA, AERIAL PARTS|ECHINACEA ROOT EXTRACT / ECHINACEA, AERIAL PARTS
C2928298|T121|1007376|RXNORM|PENTOXIFYLLINE / PROCYANIDOLIC OLIGOMER|PENTOXIFYLLINE / PROCYANIDOLIC OLIGOMER
C2928301|T121|1007379|RXNORM|ALUMINUM HYDROXIDE / BISMUTH SUBNITRATE / MAGNESIUM HYDROXIDE|ALUMINUM HYDROXIDE / BISMUTH SUBNITRATE / MAGNESIUM HYDROXIDE
C2928300|T121|1007378|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL / VITAMIN K 1|CALCIUM CARBONATE / CHOLECALCIFEROL / VITAMIN K 1
C2364524|T129|857917|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007, IVR-148 (H1N1) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007, IVR-148 (H1N1) STRAIN
C0162969|T121|59038|RXNORM|CHITOSAN|CHITOSAN
C0771458|T121|236206|RXNORM|DIISOPROMINE|DIISOPROMINE
C1120952|T125|326374|RXNORM|NORELGESTROMIN|NORELGESTROMIN
C2728174|T129|1011412|RXNORM|TANGERINE ALLERGENIC EXTRACT|TANGERINE ALLERGENIC EXTRACT
C0766108|T121|233603|RXNORM|CLEVIDIPINE|CLEVIDIPINE
C2728178|T129|1011418|RXNORM|WATERCRESS ALLERGENIC EXTRACT|WATERCRESS ALLERGENIC EXTRACT
C0002412|T121|623|RXNORM|AMBENONIUM|AMBENONIUM
C0244713|T129|72257|RXNORM|INTERFERON BETA-1B|INTERFERON BETA-1B
C0256089|T121|76887|RXNORM|QUINAGOLIDE|QUINAGOLIDE
C3848704|T121|1545902|RXNORM|NALOXONE / OXYCODONE|NALOXONE / OXYCODONE
C1377670|T121|446248|RXNORM|MELITRACEN|MELITRACEN
C0012341|T121|3435|RXNORM|IODOQUINOL|IODOQUINOL
C0012341|T121|3435|RXNORM|IODOQUINOL|IODOQUINOL
C0035924|T005|1365969|RXNORM|RUBELLA VIRUS|RUBELLA VIRUS
C0002436|T195|627|RXNORM|AMDINOCILLIN PIVOXIL|AMDINOCILLIN PIVOXIL
C0030903|T121|8015|RXNORM|PENTYLENETETRAZOLE|PENTAETRAZOL
C0030899|T121|8013|RXNORM|PENTOXIFYLLINE|PENTOXIFYLLINE
C0030896|T195|8011|RXNORM|PENTOSTATIN|PENTOSTATIN
C0030895|T121|8010|RXNORM|SODIUM STIBOGLUCONATE|SODIUM STIBOGLUCONATE
C0028158|T196|7456|RXNORM|NITROGEN|NITROGEN
C0028156|T121|7454|RXNORM|NITROFURANTOIN|NITROFURANTOIN
C0028157|T121|7455|RXNORM|NITROFURAZONE|NITROFURAZONE
C1874396|T121|689609|RXNORM|ATROPINE / MEPERIDINE|ATROPINE / MEPERIDINE
C1874395|T121|689608|RXNORM|ATROPINE / KAOLIN / PHENOBARBITAL|ATROPINE / KAOLIN / PHENOBARBITAL
C1874393|T121|689606|RXNORM|ATROPINE / HYOSCYAMINE / PHENOBARBITAL / SCOPOLAMINE|ATROPINE / HYOSCYAMINE / PHENOBARBITAL / SCOPOLAMINE
C3463993|T129|1299981|RXNORM|SIBERIAN ELM POLLEN EXTRACT|ULMUS PUMILA POLLEN EXTRACT
C0851344|T121|258494|RXNORM|EXEMESTANE|EXEMESTANE
C3474021|T121|1299989|RXNORM|AMERICAN ELM POLLEN EXTRACT / SIBERIAN ELM POLLEN EXTRACT|AMERICAN ELM POLLEN EXTRACT / SIBERIAN ELM POLLEN EXTRACT
C0007010|T196|2032|RXNORM|CARBON BLACK|CARBON BLACK
C3499505|T109|1312365|RXNORM|CHRYSANTHELLUM INDICUM FLOWER OIL|CHRYSANTHELLUM INDICUM FLOWER OIL
C1445771|T121|466537|RXNORM|MENTHOL / METHYL SALICYLATE|MENTHOL / METHYL SALICYLATE
C0057269|T130|1312367|RXNORM|DEHYDROACETIC ACID|DEHYDROACETIC ACID
C3499506|T121|1312366|RXNORM|CITRIC ACID ACETATE|CITRIC ACID ACETATE
C1451179|T109|1312361|RXNORM|CETEARYL ISONONANOATE|CETEARYL ISONONANOATE
C1686337|T109|1312360|RXNORM|C10-18 TRIGLYCERIDES|C10-18 TRIGLYCERIDES
C3541343|T121|1421430|RXNORM|SALMON PREPARATION|SALMON PREPARATION
C0650224|T131|1312362|RXNORM|CHLOROMETHYL METHYL ETHER|CHLOROMETHYL METHYL ETHER
C0700602|T121|203219|RXNORM|EVENING PRIMROSE OIL|EVENING PRIMROSE OIL
C0663344|T121|190410|RXNORM|FLUCLORONIDE|FLUCLORONIDE
C3256459|T121|1312369|RXNORM|TUSSILAGO FARFARA EXTRACT|TUSSILAGO FARFARA EXTRACT
C3256383|T121|1312368|RXNORM|TRIDECETH-9|TRIDECETH-9
C3541336|T109|1421438|RXNORM|PACIFIC COD PREPARATION|PACIFIC COD PREPARATION
C0064567|T121|28381|RXNORM|LACHESINE|LACHESINE
C2928769|T121|1007855|RXNORM|HISTIDINE / ZINC SULFATE|HISTIDINE / ZINC SULFATE
C2727871|T129|889602|RXNORM|NORTHERN PIKE ALLERGENIC EXTRACT|NORTHERN PIKE ALLERGENIC EXTRACT
C0064568|T121|28382|RXNORM|LACIDIPINE|LACIDIPINE
C0718013|T121|214791|RXNORM|POTASSIUM BICARBONATE / SODIUM BICARBONATE|POTASSIUM BICARBONATE / SODIUM BICARBONATE
C0718016|T121|214793|RXNORM|POTASSIUM IODIDE / THEOPHYLLINE|POTASSIUM IODIDE / THEOPHYLLINE
C0718014|T121|214792|RXNORM|POTASSIUM CHLORIDE / SODIUM CHLORIDE|POTASSIUM CHLORIDE / SODIUM CHLORIDE
C0718014|T121|214792|RXNORM|POTASSIUM CHLORIDE / SODIUM CHLORIDE|POTASSIUM CHLORIDE / SODIUM CHLORIDE
C0057577|T121|22672|RXNORM|DETOMIDINE|DETOMIDINE
C2928123|T121|1007201|RXNORM|4-CYMENE / CHLORPROETHAZINE|4-CYMENE / CHLORPROETHAZINE
C0120446|T123|50675|RXNORM|GUANIDINE|GUANIDINE
C0056592|T121|1311216|RXNORM|CUPRIC ACETATE|CUPRIC ACETATE
C0391001|T129|120608|RXNORM|PEGINTERFERON ALFA-2A|PEGINTERFERON ALFA-2A
C0724689|T129|221158|RXNORM|S TYPHI (TY-2 STRAIN)|S TYPHI (TY-2 STRAIN)
C3855876|T109|1549224|RXNORM|CITRUS MAXIMA FRUIT OIL|CITRUS MAXIMA FRUIT OIL
C2980958|T121|1094282|RXNORM|MILBEMYCIN OXIME / SPINOSAD|MILBEMYCIN OXIME / SPINOSAD
C2740841|T129|899873|RXNORM|PAPRIKA ALLERGENIC EXTRACT|PAPRIKA ALLERGENIC EXTRACT
C2740844|T129|899877|RXNORM|PARSLEY ALLERGENIC EXTRACT|PARSLEY ALLERGENIC EXTRACT
C0048220|T121|15002|RXNORM|4-CYMENE|4-CYMENE
C0717737|T121|214535|RXNORM|ENALAPRIL / FELODIPINE|ENALAPRIL / FELODIPINE
C2047880|T121|818715|RXNORM|IDEBENONE / VITAMIN E|IDEBENONE / VITAMIN E
C0717738|T121|214536|RXNORM|ENALAPRIL / HYDROCHLOROTHIAZIDE|ENALAPRIL / HYDROCHLOROTHIAZIDE
C0717439|T121|214247|RXNORM|ASCORBIC ACID / FERROUS FUMARATE|ASCORBIC ACID / FERROUS FUMARATE
C0063757|T130|27729|RXNORM|IODIXANOL|IODIXANOL
C0717441|T121|214249|RXNORM|ASPIRIN / BUTALBITAL|ASPIRIN / BUTALBITAL
C0717440|T121|214248|RXNORM|ASCORBIC ACID / FERROUS SULFATE|ASCORBIC ACID / FERROUS SULFATE
C0717741|T121|214539|RXNORM|EPHEDRINE / POTASSIUM IODIDE|EPHEDRINE / POTASSIUM IODIDE
C0717740|T121|214538|RXNORM|EPHEDRINE / GUAIFENESIN|EPHEDRINE / GUAIFENESIN
C0055923|T195|21272|RXNORM|CLOMOCYCLINE|CLOMOCYCLINE
C0031849|T121|8299|RXNORM|PHYSOSTIGMINE|PHYSOSTIGMINE
C0031849|T121|8299|RXNORM|PHYSOSTIGMINE|PHYSOSTIGMINE
C0257928|T197|77754|RXNORM|FERUMOXSIL|FERUMOXSIL
C0001771|T130|397|RXNORM|AGAR|AGAR
C0032493|T121|8521|RXNORM|COW SKIN EXTRACT|POLYGELINE
C1700730|T109|1552337|RXNORM|NETUPITANT|NETUPITANT
C2701705|T129|852634|RXNORM|ALFALFA POLLEN EXTRACT|MEDICAGO SATIVA POLLEN EXTRACT
C0081002|T121|40450|RXNORM|PIDOTIMOD|PIDOTIMOD
C3255918|T109|1306153|RXNORM|CITRUS AURANTIUM LEAFY TWIG OIL|CITRUS AURANTIUM LEAFY TWIG OIL
C0062168|T130|1364568|RXNORM|N-(HYDROXYETHYL)ETHYLENEDIAMINETRIACETIC ACID|N-(HYDROXYETHYL)ETHYLENEDIAMINETRIACETIC ACID
C0068881|T121|31901|RXNORM|NITROXOLINE|NITROXOLINE
C0043031|T131|11289|RXNORM|WARFARIN|WARFARIN
C3245116|T121|1190311|RXNORM|CHLOPHEDIANOL / CHLORCYCLIZINE / PHENYLEPHRINE|CHLOPHEDIANOL / CHLORCYCLIZINE / PHENYLEPHRINE
C0051522|T197|17621|RXNORM|ALUMINUM SULFATE|ALUMINUM SULFATE
C0051522|T197|17621|RXNORM|ALUMINUM SULFATE|ALUMINUM SULFATE
C0051528|T121|17627|RXNORM|ALVERINE|ALVERINE
C0064961|T121|28701|RXNORM|LIDAMIDINE|LIDAMIDINE
C3832720|T109|1539416|RXNORM|TREMELLA FUCIFORMIS WHOLE EXTRACT|TREMELLA FUCIFORMIS WHOLE EXTRACT
C0013547|T121|3743|RXNORM|ECONAZOLE|ECONAZOLE
C1095911|T121|1441652|RXNORM|WHEAT PREPARATION|WHEAT PREPARATION
C3832721|T109|1539417|RXNORM|OXALIS CORNICULATA WHOLE EXTRACT|OXALIS CORNICULATA WHOLE EXTRACT
C3818774|T121|1492184|RXNORM|TILIA AMERICANA FLOWER EXTRACT|TILIA AMERICANA FLOWER EXTRACT
C0082500|T109|1426475|RXNORM|ETHYL SEBACATE|DIETHYL SEBACATE
C3255931|T121|1426474|RXNORM|DIACETYLATED MONOGLYCERIDES|ACETYLATED MONOGLYCERIDES
C3257080|T109|1426473|RXNORM|LIME EXTRACT|LIME EXTRACT
C0075491|T120|1426472|RXNORM|SUDAN III|D&C RED NO. 17
C3255678|T109|1426471|RXNORM|HEXANOYL DIPEPTIDE-3 NORLEUCINE ACETATE|HEXANOYL DIPEPTIDE-3 NORLEUCINE ACETATE
C0113723|T122|1426470|RXNORM|DICHLOROFLUOROMETHANE|DICHLOROMONOFLUOROMETHANE
C3832724|T109|1539420|RXNORM|ROSA DAMASCENA FLOWER WAX|ROSA DAMASCENA FLOWER WAX
C2701587|T129|852450|RXNORM|WHITE ASH POLLEN EXTRACT|FRAXINUS AMERICANA POLLEN EXTRACT
C3813720|T121|1539415|RXNORM|TAGETES ERECTA WHOLE EXTRACT|TAGETES ERECTA WHOLE EXTRACT
C3488089|T197|1311377|RXNORM|POTASSIUM SILICATE|POTASSIUM SILICATE
C3818773|T109|1492189|RXNORM|PEG-80 GLYCERYL COCOATE|PEG-80 GLYCERYL COCOATE
C3497038|T121|1426479|RXNORM|MENTHONE 1,2-GLYCEROL KETAL, (-)-|MENTHONE 1,2-GLYCEROL KETAL, (-)-
C0982245|T121|1426478|RXNORM|LANOLIN ALCOHOLS|LANOLIN ALCOHOLS
C3255952|T109|1309488|RXNORM|MALVA SYLVESTRIS FLOWERING TOP EXTRACT|HIGH MALLOW FLOWERING TOP EXTRACT
C3255785|T109|1309489|RXNORM|OCIMUM BASILICUM FLOWERING TOP EXTRACT|OCIMUM BASILICUM FLOWERING TOP EXTRACT
C0893761|T121|623400|RXNORM|LACOSAMIDE|LACOSAMIDE
C0770947|T121|235776|RXNORM|POTASSIUM HYDROXYQUINOLINE SULFATE|POTASSIUM HYDROXYQUINOLINE SULFATE
C3504647|T121|1356342|RXNORM|EUCALYPTOL / THYMOL|EUCALYPTOL / THYMOL
C3858059|T121|1550699|RXNORM|KENTUCKY BLUEGRASS POLLEN EXTRACT / ORCHARD GRASS POLLEN EXTRACT / PERENNIAL RYE GRASS POLLEN EXTRACT / SWEET VERNAL GRASS POLLEN EXTRACT / TIMOTHY GRASS POLLEN EXTRACT|KENTUCKY BLUEGRASS POLLEN EXTRACT / ORCHARD GRASS POLLEN EXTRACT / PERENNIAL RYE GRASS POLLEN EXTRACT / SWEET VERNAL GRASS POLLEN EXTRACT / TIMOTHY GRASS POLLEN EXTRACT
C3255935|T109|1309481|RXNORM|HYDROGENATED MENHADEN OIL|HYDROGENATED MENHADEN OIL
C3488965|T121|1309483|RXNORM|ULMUS PROCERA FLOWERING TWIG EXTRACT|ULMUS PROCERA FLOWERING TWIG EXTRACT
C3488971|T121|1309484|RXNORM|ULMUS RUBRA BARK EXTRACT|ULMUS RUBRA BARK EXTRACT
C3488980|T121|1309485|RXNORM|VITIS VINIFERA FLOWERING TOP EXTRACT|VITIS VINIFERA FLOWERING TOP EXTRACT
C3256815|T109|1309486|RXNORM|VITIS VINIFERA FRUIT OIL|VITIS VINIFERA FRUIT OIL
C3255851|T109|1309487|RXNORM|MACHILUS THUNBERGII BARK EXTRACT|MACHILUS THUNBERGII BARK EXTRACT
C3489010|T121|1338938|RXNORM|PYRROLE|PYRROLE
C2741301|T129|900788|RXNORM|MAPLE LEAF SYCAMORE POLLEN EXTRACT|PLANTUS HYBRIDA POLLEN EXTRACT
C0148398|T121|57954|RXNORM|VINBURNINE|VINBURNINE
C2001271|T121|787390|RXNORM|TAPENTADOL|TAPENTADOL
C2722027|T129|895582|RXNORM|AVOCADO ALLERGENIC EXTRACT|PERSEA GRATISSIMA ALLERGENIC EXTRACT
C3833115|T121|1540525|RXNORM|AMINOETHYLPHOSPHINIC ACID|AMINOETHYLPHOSPHINIC ACID
C0039854|T195|10463|RXNORM|THIAMPHENICOL|THIAMPHENICOL
C0125995|T121|52103|RXNORM|LITHIUM ACETATE|LITHIUM ACETATE
C0041984|T121|11017|RXNORM|URIDINE|URIDINE
C3205299|T121|1150462|RXNORM|DIMETHICONE / LANOLIN / ZINC OXIDE|DIMETHICONE / LANOLIN / ZINC OXIDE
C3255872|T109|1367148|RXNORM|STEARETH-15|STEARETH-15
C0125997|T121|52105|RXNORM|LITHIUM CITRATE|LITHIUM CITRATE
C2827228|T130|1367145|RXNORM|LAURETH-2|LAURETH-2
C3255705|T109|1367144|RXNORM|NEOPENTYL GLYCOL DICAPRATE|NEOPENTYL GLYCOL DICAPRATE
C3255871|T109|1367147|RXNORM|STEARETH-10|STEARETH-10
C2699492|T121|1367146|RXNORM|SORBITAN|SORBITAN
C2826070|T121|1367141|RXNORM|POVIDONE K25|POVIDONE K25
C3205330|T121|1367143|RXNORM|POLYQUATERNIUM-10 (400 CPS AT 2%)|POLYQUATERNIUM-10 (400 CPS AT 2%)
C3159526|T122|1367142|RXNORM|POLYSILICONE-15|POLYSILICONE-15
C2146622|T121|817356|RXNORM|ACETAMINOPHEN / CODEINE / IBUPROFEN|ACETAMINOPHEN / CODEINE / IBUPROFEN
C0061008|T130|25544|RXNORM|GALLIUM NITRATE|GALLIUM NITRATE
C3488556|T121|1309737|RXNORM|VERATRUM VIRIDE ROOT EXTRACT|VERATRUM VIRIDE ROOT EXTRACT
C1874541|T121|710957|RXNORM|BETA CAROTENE / VITAMIN A|BETA CAROTENE / VITAMIN A
C2345399|T121|1376148|RXNORM|GAMMA-UNDECALACTONE|GAMMA-UNDECALACTONE
C3488427|T121|1309738|RXNORM|COCHLEARIA OFFICINALIS FLOWERING TOP EXTRACT|COCHLEARIA OFFICINALIS FLOWERING TOP EXTRACT
C3488050|T121|1309739|RXNORM|CENTAURIUM ERYTHRAEA FLOWER EXTRACT|CENTAURIUM ERYTHRAEA FLOWER EXTRACT
C0000992|T121|173|RXNORM|ACETOHEXAMIDE|ACETOHEXAMIDE
C1965461|T121|730907|RXNORM|VITIS EXTRACT|VITIS EXTRACT
C0789408|T129|248123|RXNORM|CAT HAIR EXTRACT|FELIS CATUS HAIR EXTRACT
C0071755|T197|34300|RXNORM|POTASSIUM CARBONATE|POTASSIUM CARBONATE
C1576662|T121|485853|RXNORM|SENNA LEAF EXTRACT|SENNA LEAF EXTRACT
C0103045|T121|46303|RXNORM|AMISULPRIDE|AMISULPRIDE
C0103049|T121|46307|RXNORM|AMLEXANOX|AMLEXANOX
C2928304|T121|1007382|RXNORM|SODIUM BITARTRATE / SODIUM PERBORATE|SODIUM BITARTRATE / SODIUM PERBORATE
C0059792|T130|1540523|RXNORM|ETHYLBENZENE|ETHYLBENZENE
C0085174|T121|42331|RXNORM|MISOPROSTOL|MISOPROSTOL
C0085173|T121|42330|RXNORM|TERFENADINE|TERFENADINE
C0085176|T121|42333|RXNORM|TRIMETREXATE|TRIMETREXATE
C3855139|T109|1547471|RXNORM|CELOSIA CRISTATA FLOWER EXTRACT|CELOSIA CRISTATA FLOWER EXTRACT
C3256058|T109|1307888|RXNORM|MELALEUCA QUINQUENERVIA LEAF OIL|MELALEUCA QUINQUENERVIA LEAF OIL
C1165265|T121|349656|RXNORM|GINSENOSIDE|GINSENOSIDE
C0752270|T121|228041|RXNORM|ECHINACEA PREPARATION|ECHINACEA PREPARATION
C0524639|T125|134404|RXNORM|UROFOLLITROPIN|UROFOLLITROPIN
C3257435|T121|1307886|RXNORM|LAVANDULA ANGUSTIFOLIA FLOWER EXTRACT|LAVANDULA ANGUSTIFOLIA FLOWER EXTRACT
C3255728|T121|1307887|RXNORM|HAMAMELIS VIRGINIANA LEAF EXTRACT|HAMAMELIS VIRGINIANA LEAF EXTRACT
C0039623|T121|10390|RXNORM|TETRABENAZINE|TETRABENAZINE
C0039629|T121|10391|RXNORM|TETRACAINE|TETRACAINE
C0039629|T121|10391|RXNORM|TETRACAINE|TETRACAINE
C0039629|T121|10391|RXNORM|TETRACAINE|TETRACAINE
C0014448|T120|1310593|RXNORM|EOSINE YELLOWISH|D&C RED NO. 22
C0032479|T121|1310594|RXNORM|POLYETHYLENE GLYCOL 4000|POLYETHYLENE GLYCOL 4000
C0039644|T195|10395|RXNORM|TETRACYCLINE|TETRACYCLINE
C0039644|T195|10395|RXNORM|TETRACYCLINE|TETRACYCLINE
C0039644|T195|10395|RXNORM|TETRACYCLINE|TETRACYCLINE
C0039644|T195|10395|RXNORM|TETRACYCLINE|TETRACYCLINE
C1337247|T121|1310598|RXNORM|POLYETHYLENE GLYCOL 600|POLYETHYLENE GLYCOL 600
C3256296|T121|1310599|RXNORM|CARBOMER COPOLYMER TYPE A|CARBOMER COPOLYMER TYPE A (ALLYL PENTAERYTHRITOL CROSSLINKED)
C3855138|T109|1547470|RXNORM|BRUCEA JAVANICA WHOLE EXTRACT|BRUCEA JAVANICA WHOLE EXTRACT
C0031376|T121|8119|RXNORM|PHENAZOCINE|PHENAZOCINE
C1601139|T121|539399|RXNORM|FERRIC HEXACYANOFERRATE|FERRIC HEXACYANOFERRATE
C3542908|T109|1376501|RXNORM|HUPERZIA SERRATA EXTRACT|HUPERZIA SERRATA EXTRACT
C0027235|T121|7213|RXNORM|IPRATROPIUM|IPRATROPIUM
C0027235|T121|7213|RXNORM|IPRATROPIUM|IPRATROPIUM
C1562066|T121|597159|RXNORM|NAPHAZOLINE / PHENIRAMINE|NAPHAZOLINE / PHENIRAMINE
C2927833|T121|1006909|RXNORM|SHARK CARTILAGE EXTRACT / SQUALENE|SHARK CARTILAGE EXTRACT / SQUALENE
C2927832|T121|1006908|RXNORM|TESTOSTERONE 17-PHENYLPROPIONATE / TESTOSTERONE DECANOATE / TESTOSTERONE ISOCAPROATE / TESTOSTERONE PROPIONATE|TESTOSTERONE 17-PHENYLPROPIONATE / TESTOSTERONE DECANOATE / TESTOSTERONE ISOCAPROATE / TESTOSTERONE PROPIONATE
C0022949|T123|6211|RXNORM|LACTOSE|LACTOSE
C2929914|T121|1009019|RXNORM|CHLORHEXIDINE / COAL TAR|CHLORHEXIDINE / COAL TAR
C2927825|T121|1006901|RXNORM|CASCARA SAGRADA / DEHYDROCHOLATE|CASCARA SAGRADA / DEHYDROCHOLATE
C2927824|T121|1006900|RXNORM|GLUTAMATE / MAGNESIUM CITRATE|GLUTAMATE / MAGNESIUM CITRATE
C2927827|T121|1006903|RXNORM|PANCREATIN / VITAMIN B6|PANCREATIN / VITAMIN B6
C1966230|T121|1009015|RXNORM|AMLODIPINE / OLMESARTAN|AMLODIPINE / OLMESARTAN
C2929907|T121|1009012|RXNORM|ETHANOL / SULFUR / ZINC OXIDE / ZINC SULFATE|ETHANOL / SULFUR / ZINC OXIDE / ZINC SULFATE
C2927828|T121|1006904|RXNORM|HEPARINOIDS / HYALURONIDASE|HEPARINOIDS / HYALURONIDASE
C2927831|T121|1006907|RXNORM|ETHANOL / GLUCOSE|ETHANOL / GLUCOSE
C0022957|T121|6218|RXNORM|LACTULOSE|LACTULOSE
C0025616|T125|6818|RXNORM|METHANDROSTENOLONE|METHANDROSTENOLONE
C0025605|T121|6813|RXNORM|METHADONE|METHADONE
C0025603|T195|6812|RXNORM|METHACYCLINE|METHACYCLINE
C0025607|T121|6814|RXNORM|METHADYL ACETATE|METHADYL ACETATE
C0025615|T125|6817|RXNORM|METHANDRIOL|METHANDRIOL
C0025611|T131|6816|RXNORM|METHAMPHETAMINE|METHAMPHETAMINE
C0040160|T125|10579|RXNORM|THYROTROPIN|THYROTROPIN
C0982291|T121|1425924|RXNORM|MYRISTYL MYRISTATE|MYRISTYL MYRISTATE
C3256308|T121|1425926|RXNORM|MODIFIED CORN STARCH (1-OCTENYL SUCCINIC ANHYDRIDE)|MODIFIED CORN STARCH (1-OCTENYL SUCCINIC ANHYDRIDE)
C3256458|T121|1425927|RXNORM|TROPAEOLUM MAJUS EXTRACT|TROPAEOLUM MAJUS EXTRACT
C1455035|T125|475230|RXNORM|DEGARELIX|DEGARELIX
C0040134|T125|10572|RXNORM|THYROID (USP)|THYROID (USP)
C2365115|T109|1425923|RXNORM|MYRISTYL LAURATE|MYRISTYL LAURATE
C0064080|T109|1362928|RXNORM|ISOSTEARYL ALCOHOL|ISOSTEARYL ALCOHOL
C0066255|T109|1362929|RXNORM|METHYL ISOBUTYL KETONE|METHYL ISOBUTYL KETONE
C0058163|T130|1362925|RXNORM|DIISOPROPYLAMINE|DIISOPROPYLAMINE
C0058252|T131|1362926|RXNORM|DIMETHYLAMPHETAMINE|DIMETHYLAMPHETAMINE
C0058632|T121|1362927|RXNORM|DODECYL SULFATE|LAURYL SULFATE
C0063348|T116|1362920|RXNORM|PENTIGIDE|PENTIGIDE
C0057934|T109|1362921|RXNORM|DIETHYL PHTHALATE|DIETHYL PHTHALATE
C0142928|T121|1311370|RXNORM|SODIUM SUCCINATE|SODIUM SUCCINATE
C0051244|T121|17384|RXNORM|ALUMINUM HYDROXIDE / MAGNESIUM CARBONATE|ALUMINUM HYDROXIDE / MAGNESIUM CARBONATE
C0001134|T197|236|RXNORM|HEPARIN, BOVINE|ACIDULATED PHOSPHATE FLUORIDE
C0445746|T007|1310846|RXNORM|PROTEUS INCONSTANS|PROTEUS INCONSTANS
C0314879|T007|1310844|RXNORM|BACILLUS COAGULANS|BACILLUS COAGULANS
C0317592|T007|1310845|RXNORM|LACTOBACILLUS HELVETICUS|LACTOBACILLUS HELVETICUS
C2093587|T129|852074|RXNORM|WING SCALE POLLEN EXTRACT|ATRIPLEX CANESCENS POLLEN EXTRACT
C0331721|T007|1310848|RXNORM|APHANIZOMENON FLOS-AQUAE|APHANIZOMENON FLOS-AQUAE
C0071120|T121|33758|RXNORM|PIPOXOLAN|PIPOXOLAN
C0072171|T121|34644|RXNORM|PROPENTOFYLLINE|PROPENTOFYLLINE
C0771394|T197|1427203|RXNORM|ALUMINUM SODIUM SILICATE|SODIUM ALUMINIUM SILICATE
C0007267|T123|1362697|RXNORM|CARNOSINE|CARNOSINE
C0006632|T196|1362694|RXNORM|CADMIUM|CADMIUM
C0002620|T197|1362695|RXNORM|AMMONIUM SULFATE|AMMONIUM SULFATE
C0063127|T122|1362692|RXNORM|2-HYDROXYETHYL METHACRYLATE|2-HYDROXYETHYL METHACRYLATE
C3484565|T121|1427206|RXNORM|LACHNANTHES CAROLINIANA EXTRACT|LACHNANTHES CAROLINIANA EXTRACT
C0443371|T109|1362691|RXNORM|1-BUTENE|1-BUTENE
C0318389|T005|1427209|RXNORM|HUMAN COXSACKIEVIRUS B1|HUMAN COXSACKIEVIRUS B1
C3486816|T121|1427208|RXNORM|OVEMOTIDE|OVEMOTIDE
C0008238|T131|1362698|RXNORM|CHLOROFORM|CHLOROFORM
C0021223|T196|1362699|RXNORM|INDIUM|INDIUM
C2216441|T121|1008699|RXNORM|MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE|MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE
C2216441|T121|1008699|RXNORM|MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE|MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE
C3153362|T121|1099032|RXNORM|BIOTIN / DEXPANTHENOL / NIACINAMIDE / ZINC PYRITHIONE|BIOTIN / DEXPANTHENOL / NIACINAMIDE / ZINC PYRITHIONE
C3497970|T121|1311615|RXNORM|KIGELIA AFRICANA FRUIT EXTRACT|KIGELIA AFRICANA FRUIT EXTRACT
C2929593|T121|1008693|RXNORM|PHENOLPHTHALEIN / RHUBARB PREPARATION|PHENOLPHTHALEIN / RHUBARB PREPARATION
C2929592|T121|1008692|RXNORM|ESTRADIOL / ESTRIOL / LEVONORGESTREL|ESTRADIOL / ESTRIOL / LEVONORGESTREL
C2929591|T121|1008691|RXNORM|CAFFEINE / DIMENHYDRINATE / SCOPOLAMINE|CAFFEINE / DIMENHYDRINATE / SCOPOLAMINE
C2929590|T121|1008690|RXNORM|ALLOBARBITAL / AMINOPYRINE|ALLOBARBITAL / AMINOPYRINE
C2929596|T121|1008696|RXNORM|DALTEPARIN / DIHYDROERGOTAMINE|DALTEPARIN / DIHYDROERGOTAMINE
C2929595|T121|1008695|RXNORM|ARGININE / CALCIUM CARBONATE|ARGININE / CALCIUM CARBONATE
C2929594|T121|1008694|RXNORM|METHENAMINE / SULFUR|METHENAMINE / SULFUR
C3265534|T121|1371995|RXNORM|LAMINARIA ANGUSTATA EXTRACT|LAMINARIA ANGUSTATA EXTRACT
C2948080|T121|1371994|RXNORM|SYNTHETIC CAMPHOR|SYNTHETIC CAMPHOR
C3495097|T121|1371997|RXNORM|STELLARIA MEDIA EXTRACT|STELLARIA MEDIA EXTRACT
C0771636|T121|1371996|RXNORM|VIOLA TRICOLOR EXTRACT|VIOLA TRICOLOR EXTRACT
C3486717|T121|1355830|RXNORM|PROTORTONIA CACTI PREPARATION|PROTORTONIA CACTI PREPARATION
C3486746|T121|1355831|RXNORM|CLEMATIS VITALBA FLOWER EXTRACT|CLEMATIS VITALBA FLOWER EXTRACT
C3486778|T121|1355832|RXNORM|DRYOPTERIS FILIX-MAS ROOT EXTRACT|DRYOPTERIS FILIX-MAS ROOT EXTRACT
C3486840|T121|1355833|RXNORM|PASSIFLORA INCARNATA FLOWER EXTRACT|PASSIFLORA INCARNATA FLOWER EXTRACT
C3465257|T121|1311610|RXNORM|INONOTUS OBLIQUUS FRUITING BODY EXTRACT|INONOTUS OBLIQUUS FRUITING BODY EXTRACT
C0006230|T121|1760|RXNORM|BROMOCRIPTINE|BROMOCRIPTINE
C0075206|T121|37071|RXNORM|STEARYL ALCOHOL|STEARYL ALCOHOL
C3486813|T121|1371999|RXNORM|ONOPORDUM EXTRACT|ONOPORDUM EXTRACT
C0006246|T121|1767|RXNORM|BROMPHENIRAMINE|BROMPHENIRAMINE
C3265002|T168|1311611|RXNORM|AVOCADO OIL|AVOCADO OIL
C3700907|T109|1485540|RXNORM|MYRISTAMIDOPROPYLAMINE OXIDE|MYRISTAMIDOPROPYLAMINE OXIDE
C0066040|T121|29590|RXNORM|METACLAZEPAM HYDROCHLORIDE|METACLAZEPAM HYDROCHLORIDE
C3700906|T109|1485541|RXNORM|C12-20 ACID PEG-8 ESTER|C12-20 ACID PEG-8 ESTER
C2722028|T129|891830|RXNORM|BANANA ALLERGENIC EXTRACT|BANANA ALLERGENIC EXTRACT
C3818690|T109|1537318|RXNORM|C24-28 OLEFIN|C24-28 OLEFIN
C2978518|T121|1089042|RXNORM|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE
C2929429|T121|1008525|RXNORM|CHLOPHEDIANOL / GUAIACOL ETHYLGLYCOLATE / OXATOMIDE|CHLOPHEDIANOL / GUAIACOL ETHYLGLYCOLATE / OXATOMIDE
C2929428|T121|1008524|RXNORM|AMYLMETACRESOL / DICHLOROBENZYL ALCOHOL / MENTHOL|AMYLMETACRESOL / DICHLOROBENZYL ALCOHOL / MENTHOL
C2929424|T121|1008520|RXNORM|MEGLUMINE BENZOATE / POLYSORBATES|MEGLUMINE BENZOATE / POLYSORBATES
C2929427|T121|1008523|RXNORM|AMBROXOL / CHLOPHEDIANOL|AMBROXOL / CHLOPHEDIANOL
C2929426|T121|1008522|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL / FOLIC ACID / HYDROXOCOBALAMIN|CALCIUM CARBONATE / CHOLECALCIFEROL / FOLIC ACID / HYDROXOCOBALAMIN
C3700892|T121|1486677|RXNORM|BLACK MUSTARD SEED EXTRACT|BLACK MUSTARD SEED EXTRACT
C2929433|T121|1008529|RXNORM|BELLADONNA EXTRACT, USP / CHLORPHENIRAMINE / PHENIRAMINE / PHENYLPROPANOLAMINE|BELLADONNA EXTRACT, USP / CHLORPHENIRAMINE / PHENIRAMINE / PHENYLPROPANOLAMINE
C2929432|T121|1008528|RXNORM|BORAGE OIL / GAMMA-LINOLENATE|BORAGE OIL / GAMMA-LINOLENATE
C1720044|T121|645566|RXNORM|BENDROFLUMETHIAZIDE / PROPRANOLOL|BENDROFLUMETHIAZIDE / PROPRANOLOL
C1719890|T121|645567|RXNORM|BENDROFLUMETHIAZIDE / TIMOLOL|BENDROFLUMETHIAZIDE / TIMOLOL
C0108342|T121|47686|RXNORM|CARBAMIDE PEROXIDE|CARBAMIDE PEROXIDE
C0108342|T121|47686|RXNORM|CARBAMIDE PEROXIDE|CARBAMIDE PEROXIDE
C0108342|T121|47686|RXNORM|CARBAMIDE PEROXIDE|CARBAMIDE PEROXIDE
C0005404|T123|1540|RXNORM|BILE SALTS|BILE SALTS
C0002586|T121|695|RXNORM|AMINOPYRINE|AMINOPYRINE
C3256285|T121|1311618|RXNORM|LEMON PEEL WAX|LEMON PEEL WAX
C3486783|T121|1311248|RXNORM|SUS SCROFA CARTILAGE PREPARATION|PORCINE CARTILAGE PREPARATION
C0042285|T123|11115|RXNORM|VALINE|VALINE
C3715229|T109|1541719|RXNORM|JASMINUM OFFICINALE WHOLE EXTRACT|JASMINUM OFFICINALE WHOLE EXTRACT
C0282097|T121|1311619|RXNORM|CETEARETH 20|CETEARETH 20
C3256622|T121|1312620|RXNORM|ISOPROPYL STEARATE|ISOPROPYL STEARATE
C2928725|T121|1007810|RXNORM|DODECYL SULFATE / OXYQUINOLINE|DODECYL SULFATE / OXYQUINOLINE
C3281930|T109|1312622|RXNORM|LIGUSTICUM WALLICHII WHOLE EXTRACT|LIGUSTICUM WALLICHII WHOLE EXTRACT
C2928726|T121|1007811|RXNORM|ESTROGENS, CONJUGATED (USP) / PHENOBARBITAL|ESTROGENS, CONJUGATED (USP) / PHENOBARBITAL
C0033254|T121|8718|RXNORM|PROCYCLIDINE|PROCYCLIDINE
C3254760|T121|1232311|RXNORM|SALIX NIGRA BARK EXTRACT|SALIX NIGRA BARK EXTRACT
C0304889|T127|91473|RXNORM|HALIBUT LIVER OIL|HALIBUT LIVER OIL
C0068495|T121|31575|RXNORM|MENFEGOL|MENFEGOL
C3665208|T121|1435521|RXNORM|PEG-150-DECYL ALCOHOL-SMDI COPOLYMER (1350 MPA.S AT 3%)|PEG-150-DECYL ALCOHOL-SMDI COPOLYMER (1350 MPA.S AT 3%)
C0066803|T121|30225|RXNORM|MORNIFLUMATE|MORNIFLUMATE
C0070034|T121|32863|RXNORM|PANTETHINE|PANTETHINE
C2344295|T129|798266|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18 VACCINE
C3665209|T121|1435523|RXNORM|MIMOSA PUDICA LEAF EXTRACT|MIMOSA PUDICA LEAF EXTRACT
C0163061|T121|59082|RXNORM|MYRTECAINE|MYRTECAINE
C0083858|T129|798264|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 16 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 16 VACCINE
C0010725|T121|997602|RXNORM|CITICOLINE|CITICOLINE
C2701190|T129|851955|RXNORM|SANDBUR RAGWEED POLLEN EXTRACT|AMBROSIA CHAMISSONIS POLLEN EXTRACT
C3700991|T121|1486415|RXNORM|COCONUT OIL / LINSEED OIL|COCONUT OIL / LINSEED OIL
C2938117|T129|1011627|RXNORM|SAGE LEAF ALLERGENIC EXTRACT|SALVIA OFFICINALIS ALLERGENIC EXTRACT
C0076784|T121|38365|RXNORM|TOFISOPAM|TOFISOPAM
C2342462|T121|792786|RXNORM|METHSCOPOLAMINE / PHENYLEPHRINE|METHSCOPOLAMINE / PHENYLEPHRINE
C3530615|T109|1426914|RXNORM|POLYQUATERNIUM-28 (1100000 MW)|POLYQUATERNIUM-28 (1100000 MW)
C3257696|T109|1426915|RXNORM|GLYCERYL 1,2-DIOLEATE|GLYCERYL 1,2-DIOLEATE
C0040892|T204|1426916|RXNORM|TRICHINELLA SPIRALIS|TRICHINELLA SPIRALIS
C3257019|T109|1426917|RXNORM|PORPHYRA YEZOENSIS EXTRACT|PORPHYRA YEZOENSIS EXTRACT
C0017911|T123|1426910|RXNORM|GLYCOGEN|GLYCOGEN
C0026783|T005|1426911|RXNORM|MUMPS VIRUS|MUMPS VIRUS
C3257529|T109|1426912|RXNORM|PISUM SATIVUM (PEA) EXTRACT|PISUM SATIVUM (PEA) EXTRACT
C0070422|T109|1426913|RXNORM|PERILLALDEHYDE|PERILLALDEHYDE
C3256868|T109|1426918|RXNORM|PSEUDEVERNIA FURFURACEA EXTRACT|PSEUDEVERNIA FURFURACEA EXTRACT
C3500341|T121|1314244|RXNORM|AVENA SATIVA WHOLE EXTRACT|AVENA SATIVA WHOLE EXTRACT
C1874605|T121|690637|RXNORM|BORIC ACID / ZINC OXIDE|BORIC ACID / ZINC OXIDE
C1959625|T121|704942|RXNORM|LEVISTICUM OFFICINALE LEAF EXTRACT|LEVISTICUM OFFICINALE LEAF EXTRACT
C0373704|T125|114052|RXNORM|PREGNENOLONE|PREGNENOLONE
C3282849|T122|1313719|RXNORM|POLYACRYLAMIDE (10000 MW)|POLYACRYLAMIDE (10000 MW)
C2826071|T122|1313718|RXNORM|POVIDONE K25-28|POVIDONE K25-28
C3485670|T121|1426649|RXNORM|POLYQUATERNIUM-39 (35-35-30 ACRYLIC ACID-ACRYLAMIDE-DADMAC; 1500000 MW)|POLYQUATERNIUM-39 (35-35-30 ACRYLIC ACID-ACRYLAMIDE-DADMAC; 1500000 MW)
C0164311|T116|1426644|RXNORM|ECTOINE|ECTOINE
C3255940|T121|1313712|RXNORM|HYDROLYZED GLYCOSAMINOGLYCANS (BOVINE; 50000 MW)|HYDROLYZED GLYCOSAMINOGLYCANS (BOVINE; 50000 MW)
C3255800|T121|1313711|RXNORM|POLOXAMER 335|POLOXAMER 335
C3255764|T121|1313710|RXNORM|ETHYLENE-VINYL ACETATE COPOLYMER (15% VINYL ACETATE)|ETHYLENE-VINYL ACETATE COPOLYMER (15% VINYL ACETATE)
C3530632|T121|1364991|RXNORM|TRIFOLIUM PRATENSE LEAF EXTRACT|TRIFOLIUM PRATENSE LEAF EXTRACT
C3530631|T121|1364990|RXNORM|ROSMARINUS OFFICINALIS WHOLE EXTRACT|ROSMARINUS OFFICINALIS WHOLE EXTRACT
C0127429|T130|52527|RXNORM|MEGLUMINE IOTROXINATE|MEGLUMINE IOTROXINATE
C0166532|T121|60451|RXNORM|DELMOPINOL|DELMOPINOL
C2928336|T121|1007414|RXNORM|GOTU KOLA EXTRACT / NITROFURANTOIN|GOTU KOLA EXTRACT / NITROFURANTOIN
C2928337|T121|1007415|RXNORM|ALOE EXTRACT / BUCKTHORN PREPARATION / PHENOLPHTHALEIN|ALOE EXTRACT / BUCKTHORN PREPARATION / PHENOLPHTHALEIN
C2928338|T121|1007416|RXNORM|AMOXICILLIN / PROBENECID|AMOXICILLIN / PROBENECID
C2928339|T121|1007417|RXNORM|METHYL SALICYLATE / NIACIN|METHYL SALICYLATE / NIACIN
C2928332|T121|1007410|RXNORM|CARISOPRODOL / IBUPROFEN|CARISOPRODOL / IBUPROFEN
C2928333|T121|1007411|RXNORM|CHLORPROPAMIDE / METFORMIN|CHLORPROPAMIDE / METFORMIN
C2928334|T121|1007412|RXNORM|AMBROXOL / DOXYCYCLINE|AMBROXOL / DOXYCYCLINE
C2928335|T121|1007413|RXNORM|SODIUM FLUORIDE / XYLITOL|SODIUM FLUORIDE / XYLITOL
C3256663|T121|1307675|RXNORM|ASPARAGUS COCHINCHINESIS TUBER EXTRACT|ASPARAGUS COCHINCHINESIS TUBER EXTRACT
C3475162|T121|1302826|RXNORM|PHENTERMINE / TOPIRAMATE|PHENTERMINE / TOPIRAMATE
C3256499|T121|1307677|RXNORM|ARCTIUM LAPPA FRUIT EXTRACT|ARCTIUM LAPPA FRUIT EXTRACT
C2827601|T168|1307676|RXNORM|HYDROGENATED PALM OIL|HYDROGENATED PALM OIL
C2928340|T121|1007418|RXNORM|GLUCOSAMINE / SHARK CARTILAGE EXTRACT|GLUCOSAMINE / SHARK CARTILAGE EXTRACT
C2928341|T121|1007419|RXNORM|ALOE VERA PREPARATION / DEXPANTHENOL|ALOE VERA PREPARATION / DEXPANTHENOL
C3256911|T121|1307673|RXNORM|ECHINACEA ANGUSTIFOLIA LEAF EXTRACT|ECHINACEA ANGUSTIFOLIA LEAF EXTRACT
C3256244|T109|1307672|RXNORM|PERILLA FRUTESCENS LEAF OIL|PERILLA FRUTESCENS LEAF OIL
C1874655|T121|691015|RXNORM|CALCIUM CARBONATE / MAGNESIUM HYDROXIDE / SIMETHICONE|CALCIUM CARBONATE / MAGNESIUM HYDROXIDE / SIMETHICONE
C1874654|T121|691014|RXNORM|CALCIUM CARBONATE / MAGNESIUM HYDROXIDE / PHENOBARBITAL|CALCIUM CARBONATE / MAGNESIUM HYDROXIDE / PHENOBARBITAL
C1874657|T121|691017|RXNORM|CALCIUM CARBONATE / PECTIN|CALCIUM CARBONATE / PECTIN
C1874657|T121|691017|RXNORM|CALCIUM CARBONATE / PECTIN|CALCIUM CARBONATE / PECTIN
C0040217|T121|1535217|RXNORM|TILETAMINE|TILETAMINE
C1874651|T121|691010|RXNORM|CALCIUM CARBONATE / MAGNESIUM CARBONATE / MAGNESIUM OXIDE|CALCIUM CARBONATE / MAGNESIUM CARBONATE / MAGNESIUM OXIDE
C1874653|T121|691012|RXNORM|CALCIUM CARBONATE / MAGNESIUM CARBONATE / VITAMIN D|CALCIUM CARBONATE / MAGNESIUM CARBONATE / VITAMIN D
C1609931|T129|1535218|RXNORM|SILTUXIMAB|SILTUXIMAB
C1874658|T121|691018|RXNORM|CALCIUM CARBONATE / PHENOBARBITAL|CALCIUM CARBONATE / PHENOBARBITAL
C0717833|T121|214627|RXNORM|HYDROCODONE / IBUPROFEN|HYDROCODONE / IBUPROFEN
C0061246|T121|25734|RXNORM|GESTODENE|GESTODENE
C3500337|T121|1314236|RXNORM|AMMONIAC|AMMONIAC
C3179929|T121|1248798|RXNORM|PEGINESATIDE|PEGINESATIDE
C2973895|T121|1440051|RXNORM|LIXISENATIDE|LIXISENATIDE
C3854887|T109|1546869|RXNORM|SUS SCROFA LIGAMENT PREPARATION|SUS SCROFA LIGAMENT PREPARATION
C3854886|T109|1546868|RXNORM|BOS TAURUS MAMMARY GLAND PREPARATION|BOS TAURUS MAMMARY GLAND PREPARATION
C0025497|T121|6779|RXNORM|MESORIDAZINE|MESORIDAZINE
C3853864|T109|1546861|RXNORM|ACMELLA OLERACEA WHOLE EXTRACT|ACMELLA OLERACEA WHOLE EXTRACT
C3854881|T109|1546863|RXNORM|ARTEMISIA TRIDENTATA TOP OIL|ARTEMISIA TRIDENTATA TOP OIL
C3854880|T109|1546862|RXNORM|ADONIS VERNALIS FLOWERING TOP EXTRACT|ADONIS VERNALIS FLOWERING TOP EXTRACT
C3854883|T109|1546865|RXNORM|SPARGANIUM STOLONIFERUM ROOT EXTRACT|SPARGANIUM STOLONIFERUM ROOT EXTRACT
C3854882|T109|1546864|RXNORM|CYNANCHUM PANICULATUM ROOT EXTRACT|CYNANCHUM PANICULATUM ROOT EXTRACT
C3854885|T109|1546867|RXNORM|ENTADA PHASEOLOIDES WHOLE EXTRACT|ENTADA PHASEOLOIDES WHOLE EXTRACT
C3854884|T109|1546866|RXNORM|TINOSPORA CAPILLIPES ROOT EXTRACT|TINOSPORA CAPILLIPES ROOT EXTRACT
C1874826|T121|689410|RXNORM|CHLORPHENIRAMINE / HYDROCORTISONE / PHENIRAMINE / PYRILAMINE|CHLORPHENIRAMINE / HYDROCORTISONE / PHENIRAMINE / PYRILAMINE
C3538557|T121|1373039|RXNORM|RHEUM OFFICINALE STEM EXTRACT|RHEUM OFFICINALE STEM EXTRACT
C3538552|T121|1373032|RXNORM|MIRABILIS JALAPA FLOWERING TOP EXTRACT|MIRABILIS JALAPA FLOWERING TOP EXTRACT
C1273021|T121|388458|RXNORM|CETYL DIMETHICONE|CETYL DIMETHICONE
C0037854|T121|9968|RXNORM|SPERMACETI|SPERMACETI
C3538554|T121|1373036|RXNORM|PETIVERIA ALLIACEA WHOLE EXTRACT|PETIVERIA ALLIACEA WHOLE EXTRACT
C0907828|T121|1366840|RXNORM|COCOYL ISETHIONATE|COCOYL ISETHIONATE
C0354652|T121|104486|RXNORM|NICOFURANOSE|NICOFURANOSE
C0301382|T121|89791|RXNORM|GITALIN|GITALIN
C0589330|T197|150596|RXNORM|COPPER CHLORIDE|COPPER CHLORIDE
C0022059|T121|5981|RXNORM|IPRONIAZID|IPRONIAZID
C3496089|T129|1314927|RXNORM|SALSOLA TRAGUS POLLEN EXTRACT|PRICKLY RUSSIAN THISTLE
C0050451|T121|16728|RXNORM|ACETOHYDROXAMIC ACID|ACETOHYDROXAMIC ACID
C0359620|T121|710303|RXNORM|CODEINE / IBUPROFEN|CODEINE / IBUPROFEN
C0759933|T121|231049|RXNORM|ELETRIPTAN|ELETRIPTAN
C0593879|T121|153153|RXNORM|ATENOLOL / BENDROFLUMETHIAZIDE|ATENOLOL / BENDROFLUMETHIAZIDE
C2702428|T129|1306108|RXNORM|SILVER BIRCH POLLEN ALLERGENIC EXTRACT|BETULA PENDULA POLLEN ALLERGENIC EXTRACT
C2955387|T121|1050086|RXNORM|CAMPHOR / MENTHOL / PETROLATUM|CAMPHOR / MENTHOL / PETROLATUM
C0028042|T131|1306107|RXNORM|NICOTINE BITARTRATE|NICOTINE BITARTRATE
C1337344|T121|1306100|RXNORM|BICISATE|BICISATE
C0086154|T121|1427193|RXNORM|DIETHYLDITHIOCARBAMATE|DIETHYLDITHIOCARBAMATE
C2106307|T121|818560|RXNORM|CODEINE / DIPHENHYDRAMINE|CODEINE / DIPHENHYDRAMINE
C0036023|T121|9509|RXNORM|SACCHARIN|SACCHARIN
C3645277|T121|1427197|RXNORM|DODECYL-2-N,N-DIMETHYLAMINOPROPIONATE|DODECYL-2-N,N-DIMETHYLAMINOPROPIONATE
C3489290|T197|1427195|RXNORM|EGG SHELL, COOKED|EGG SHELL, COOKED
C3695976|T109|1483423|RXNORM|EUCALYPTUS RADIATA LEAF OIL|EUCALYPTUS RADIATA LEAF OIL
C1177210|T197|1427198|RXNORM|CUPRIC CATION|CU 2+
C3695974|T121|1483425|RXNORM|LAVANDULA DENTATA WHOLE EXTRACT|LAVANDULA DENTATA WHOLE EXTRACT
C3695975|T121|1483424|RXNORM|CUPRESSUS SEMPERVIRENS WHOLE EXTRACT|CUPRESSUS SEMPERVIRENS WHOLE EXTRACT
C0036002|T123|9504|RXNORM|S-ADENOSYLMETHIONINE|S-ADENOSYLMETHIONINE
C1445742|T121|466508|RXNORM|STARCH / ZINC OXIDE|STARCH / ZINC OXIDE
C0289313|T121|84108|RXNORM|ROSIGLITAZONE|ROSIGLITAZONE
C2701825|T129|852844|RXNORM|CHINESE ELM POLLEN EXTRACT|ULMUS PARVIFOLIA POLLEN EXTRACT
C3848617|T121|1544248|RXNORM|MYRISTICA FRAGRANS WHOLE EXTRACT|MYRISTICA FRAGRANS WHOLE EXTRACT
C3848618|T121|1544247|RXNORM|IMPERATORIA OSTRUTHIA ROOT EXTRACT|IMPERATORIA OSTRUTHIA ROOT EXTRACT
C3848619|T121|1544246|RXNORM|CENTAURIUM ERYTHRAEA FLOWERING TOP EXTRACT|CENTAURIUM ERYTHRAEA FLOWERING TOP EXTRACT
C3848620|T121|1544245|RXNORM|BOS TAURUS SOMATIC NERVE PREPARATION|BOS TAURUS SOMATIC NERVE PREPARATION
C2702414|T129|901337|RXNORM|RICE ALLERGENIC EXTRACT|RICE ALLERGENIC EXTRACT
C0060231|T197|1594675|RXNORM|FERRIC CITRATE|FERRIC CITRATE
C3645278|T127|1427200|RXNORM|ASCORBYL TOCOPHERYL PHOSPHATE|ASCORBYL TOCOPHERYL PHOSPHATE
C2937591|T121|1009466|RXNORM|CARBETAPENTANE / DEXCHLORPHENIRAMINE / PHENYLEPHRINE|CARBETAPENTANE / DEXCHLORPHENIRAMINE / PHENYLEPHRINE
C0025179|T121|6704|RXNORM|MEGLUMINE|MEGLUMINE
C2741496|T129|901313|RXNORM|SPEARMINT ALLERGENIC EXTRACT|MENTHA VIRIDIS ALLERGENIC EXTRACT
C0075474|T109|1363646|RXNORM|SUCROSE ACETATE ISOBUTYRATE|SUCROSE ACETATE ISOBUTYRATE
C0075475|T121|1363647|RXNORM|SUCROSE MONOLAURATE|SUCROSE MONOLAURATE
C0075083|T130|1363644|RXNORM|SQUALANE|SQUALANE
C0075245|T121|1363645|RXNORM|STEVIOL|STEVIOL
C0074917|T121|1363643|RXNORM|SORBITAN TRIOLEATE|SORBITAN TRIOLEATE
C0097513|T121|45045|RXNORM|AVOBENZONE|AVOBENZONE
C0073689|T197|1367087|RXNORM|RUBIDIUM CHLORIDE|RUBIDIUM CHLORIDE
C0132776|T121|53750|RXNORM|NONOXYNOL-9|NONOXYNOL-9
C0040869|T121|10763|RXNORM|TRIAMTERENE|TRIAMTERENE
C0040879|T121|10767|RXNORM|TRIAZOLAM|TRIAZOLAM
C0302933|T196|90249|RXNORM|NATURAL GRAPHITE|NATURAL GRAPHITE
C3527695|T121|1360737|RXNORM|CHLOPHEDIANOL / PHENYLEPHRINE / THONZYLAMINE|CHLOPHEDIANOL / PHENYLEPHRINE / THONZYLAMINE
C3666986|T121|1438113|RXNORM|OSTREA EDULIS SHELL PREPARATION|OSTREA EDULIS SHELL PREPARATION
C2929657|T121|1008758|RXNORM|PHOLCODINE / PROMETHAZINE / PSEUDOEPHEDRINE|PHOLCODINE / PROMETHAZINE / PSEUDOEPHEDRINE
C2929658|T121|1008759|RXNORM|PHOLCODINE / SQUILL EXTRACT|PHOLCODINE / SQUILL EXTRACT
C0053122|T130|18896|RXNORM|BENTIROMIDE|BENTIROMIDE
C2929651|T121|1008752|RXNORM|PSEUDOEPHEDRINE / TRIPELENNAMINE|PSEUDOEPHEDRINE / TRIPELENNAMINE
C2929652|T121|1008753|RXNORM|DEXCHLORPHENIRAMINE / HYDROCODONE|DEXCHLORPHENIRAMINE / HYDROCODONE
C2929649|T121|1008750|RXNORM|HEPATITIS A VACCINE, INACTIVATED / HEPATITIS B VACCINE|HEPATITIS A VACCINE, INACTIVATED / HEPATITIS B SURFACE ANTIGEN VACCINE
C2929655|T121|1008756|RXNORM|BROMPHENIRAMINE / DEXTROMETHORPHAN|BROMPHENIRAMINE / DEXTROMETHORPHAN
C2929656|T121|1008757|RXNORM|LACTATE / PEPSIN A|LACTATE / PEPSIN A
C2929653|T121|1008754|RXNORM|GUAIACOLSULFONATE / SODIUM CITRATE|GUAIACOLSULFONATE / SODIUM CITRATE
C2929654|T121|1008755|RXNORM|ALANINE / ARGININE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE|ALANINE / ARGININE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE
C0077089|T121|38623|RXNORM|TRIETHANOLAMINE|TRIETHANOLAMINE
C0077091|T121|38624|RXNORM|TRIETHANOLAMINE POLYPEPTIDE OLEATE CONDENSATE|TRIETHANOLAMINE POLYPEPTIDE OLEATE CONDENSATE
C2609465|T121|1423345|RXNORM|TRIBULUS|TRIBULUS
C2747183|T129|905088|RXNORM|ACROTHECIUM ROBUSTUM ALLERGENIC EXTRACT|ACROTHECIUM ROBUSTUM ALLERGENIC EXTRACT
C1874002|T121|690195|RXNORM|ACETIC ACID / ALUMINUM SULFATE|ACETIC ACID / ALUMINUM SULFATE
C0077388|T121|38876|RXNORM|TROPATEPINE|TROPATEPINE
C0607428|T197|1363426|RXNORM|BORON NITRIDE|BORON NITRIDE
C2987417|T121|1364347|RXNORM|PONATINIB|PONATINIB
C0772394|T121|237057|RXNORM|LEPIRUDIN|LEPIRUDIN
C0772395|T121|237058|RXNORM|THONZONIUM|THONZONIUM
C0358595|T121|106642|RXNORM|DIMETHICONE / PIPENZOLATE|DIMETHICONE / PIPENZOLATE
C3848702|T121|1546166|RXNORM|APROLIUM|APROLIUM
C3486526|T121|1310128|RXNORM|COFFEA ARABICA SEED, ROASTED, EXTRACT|COFFEA ARABICA SEED, ROASTED, EXTRACT
C3651701|T109|1431715|RXNORM|SUNFLOWER SEED OIL GLYCERETH-8 ESTERS|SUNFLOWER SEED OIL GLYCERETH-8 ESTERS
C2930451|T121|1028612|RXNORM|PYRIDOXINE / THIAMINE / VITAMIN B 12|PYRIDOXINE / THIAMINE / VITAMIN B 12
C0007886|T196|1310121|RXNORM|CESIUM|CESIUM
C3497577|T121|1310120|RXNORM|BERBERIS VULGARIS ROOT EXTRACT|BERBERIS VULGARIS ROOT EXTRACT
C0016330|T196|1310123|RXNORM|FLUORINE|FLUORINE
C0008209|T196|1310122|RXNORM|CHLORINE|CHLORINE
C0016980|T196|1310124|RXNORM|GALLIUM|GALLIUM
C3486525|T109|1310127|RXNORM|CITRUS PARADISI FRUIT OIL|CITRUS PARADISI FRUIT OIL
C3486523|T121|1310126|RXNORM|BACOPA MONNIERA LEAF EXTRACT|BACOPA MONNIERA LEAF EXTRACT
C1621234|T129|612937|RXNORM|INTERFERON ALFA-N3|INTERFERON ALFA-N3
C1721300|T121|662019|RXNORM|PRALATREXATE|PRALATREXATE
C2702350|T129|892503|RXNORM|TUNA ALLERGENIC EXTRACT|TUNA ALLERGENIC EXTRACT
C2346726|T196|1546162|RXNORM|ALUMINUM CATION|ALUMINUM CATION
C2702310|T129|892507|RXNORM|ALMOND ALLERGENIC EXTRACT|ALMOND ALLERGENIC EXTRACT
C3651696|T109|1428861|RXNORM|BASIC YELLOW 57|BASIC YELLOW 57
C1702916|T121|618371|RXNORM|PENTETATE|PENTETATE
C0873197|T121|285170|RXNORM|YELLOWJACKET VENOM PROTEIN|YELLOW JACKET VENOM PROTEIN
C2928100|T121|1007178|RXNORM|COAL TAR / DODECYL SULFATE|COAL TAR / DODECYL SULFATE
C2928099|T121|1007177|RXNORM|PETROLEUM PREPARATION / PIPERONYL BUTOXIDE / PYRETHRINS|PETROLEUM PREPARATION / PIPERONYL BUTOXIDE / PYRETHRINS
C2928098|T121|1007176|RXNORM|BETA SITOSTEROL / GUGGUL LIPIDS|BETA SITOSTEROL / GUGGUL LIPIDS
C2928096|T121|1007174|RXNORM|CHLORHEXIDINE / SODIUM FLUORIDE|CHLORHEXIDINE / SODIUM FLUORIDE
C2928095|T121|1007173|RXNORM|FOLIC ACID / INTRINSIC FACTOR / VITAMIN B 12|FOLIC ACID / INTRINSIC FACTOR / VITAMIN B 12
C2928094|T121|1007172|RXNORM|ARNICA EXTRACT / ETHANOL|ARNICA EXTRACT / ETHANOL
C2928093|T121|1007171|RXNORM|ACETAMINOPHEN / CAFFEINE / HYOSCYAMUS EXTRACT|ACETAMINOPHEN / CAFFEINE / HYOSCYAMUS EXTRACT
C2928092|T121|1007170|RXNORM|PETROLATUM / SALICYLIC ACID|PETROLATUM / SALICYLIC ACID
C1874340|T121|689256|RXNORM|ASCORBIC ACID / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PYRILAMINE|ASCORBIC ACID / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PYRILAMINE
C0038702|T195|10184|RXNORM|SULFANILAMIDE|SULFANILAMIDE
C0002575|T121|689|RXNORM|ASCORBIC ACID / BIOFLAVONOIDS|AMINOPHYLLINE
C0038693|T195|10181|RXNORM|SULFAMETHOXYPYRIDAZINE|SULFAMETHOXYPYRIDAZINE
C0301249|T168|1309229|RXNORM|CINNAMON OIL|CINNAMON OIL
C0038700|T121|10183|RXNORM|SULFAMOXOLE|SULFAMOXOLE
C0304115|T109|1309224|RXNORM|SANDALWOOD OIL|SANDALWOOD OIL
C0982446|T109|1309225|RXNORM|HYDROGENATED VEGETABLE OIL|HYDROGENATED VEGETABLE OIL
C0439963|T121|1309226|RXNORM|CHAMOMILE EXTRACT|CHAMOMILE EXTRACT
C1721515|T109|1309227|RXNORM|CINNAMON OIL, LEAF|CINNAMON OIL, LEAF
C2699024|T121|1309220|RXNORM|REHMANNIA GLUTINOSA ROOT EXTRACT|REHMANNIA GLUTINOSA ROOT EXTRACT
C0038710|T195|10188|RXNORM|SULFAPYRIDINE|SULFAPYRIDINE
C1509841|T168|1309222|RXNORM|HYDROGENATED SOYBEAN OIL|HYDROGENATED SOYBEAN OIL
C0073354|T109|1309223|RXNORM|RICE BRAN OIL|RICE BRAN OIL
C0066226|T121|29742|RXNORM|METHYL ANTHRANILATE|METHYL ANTHRANILATE
C0982025|T121|314504|RXNORM|ANTI-INHIBITOR COAGULANT COMPLEX|FACTOR VIII INHIBITOR BYPASSING ACTIVITY
C0913469|T125|278739|RXNORM|PEGVISOMANT|PEGVISOMANT
C0066230|T131|29746|RXNORM|METHYL BROMIDE|METHYL BROMIDE
C0598549|T121|637485|RXNORM|IOPANOATE|IOPANOATE
C1611934|T121|857974|RXNORM|SAXAGLIPTIN|SAXAGLIPTIN
C0003995|T123|1157|RXNORM|ASPARAGINE|ASPARAGINE
C0003993|T126|1156|RXNORM|ASPARAGINASE|ASPARAGINASE
C0003968|T127|1151|RXNORM|ASCORBIC ACID|ASCORBIC ACID
C0075821|T130|37578|RXNORM|TARTARIC ACID|TARTARIC ACID
C2349153|T121|1592898|RXNORM|ROSA ARKANSANA ROOT EXTRACT|ROSA ARKANSANA ROOT EXTRACT
C2928241|T121|1007319|RXNORM|CHLOROQUINE / PROGUANIL|CHLOROQUINE / PROGUANIL
C2928240|T121|1007318|RXNORM|MENTHOL / SELENIUM SULFIDE|MENTHOL / SELENIUM SULFIDE
C2928235|T121|1007313|RXNORM|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2928234|T121|1007312|RXNORM|BENZOCAINE / GLYCERIN|BENZOCAINE / GLYCERIN
C2928233|T121|1007311|RXNORM|BENZOCAINE / GLYCERIN / MENTHOL|BENZOCAINE / GLYCERIN / MENTHOL
C2928232|T121|1007310|RXNORM|ASCORBIC ACID / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / VITAMIN B 12|ASCORBIC ACID / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / VITAMIN B 12
C2928239|T121|1007317|RXNORM|ASCORBIC ACID / FERROUS SULFATE / VITAMIN A / VITAMIN D|ASCORBIC ACID / FERROUS SULFATE / VITAMIN A / VITAMIN D
C2928238|T121|1007316|RXNORM|DEXPANTHENOL / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC SULFATE|DEXPANTHENOL / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC SULFATE
C2928237|T121|1007315|RXNORM|GLYCINE / SODIUM CHLORIDE|GLYCINE / SODIUM CHLORIDE
C2928236|T121|1007314|RXNORM|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / SODIUM PHOSPHATE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / SODIUM PHOSPHATE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C3819181|T121|1491503|RXNORM|KETOPROFEN / LIDOCAINE|KETOPROFEN / LIDOCAINE
C0062961|T121|1374845|RXNORM|TRAMIPROSATE|TRAMIPROSATE
C3555516|T122|1374847|RXNORM|BEHENYL OLIVATE|BEHENYL OLIVATE
C0054483|T197|1311526|RXNORM|CALCIUM SILICATE|CALCIUM SILICATE
C0059459|T121|24263|RXNORM|EPOMEDIOL|EPOMEDIOL
C0003999|T121|1311524|RXNORM|ASPARTAME|ASPARTAME
C0068700|T121|31748|RXNORM|NICORANDIL|NICORANDIL
C0081959|T195|1311521|RXNORM|CEFTIOFUR|CEFTIOFUR
C2928128|T121|1007206|RXNORM|MAGNESIUM CHLORIDE / TUBOCURARINE|MAGNESIUM CHLORIDE / TUBOCURARINE
C3256027|T109|1311528|RXNORM|COCAMIDOPROPYL PG-DIMONIUM CHLORIDE PHOSPHATE|COCAMIDOPROPYL PROPYLENE GLYCOL-DIMONIUM CHLORIDE PHOSPHATE
C3488588|T121|1311529|RXNORM|COFFEA ARABICA FRUIT EXTRACT|COFFEA ARABICA FRUIT EXTRACT
C3486222|T121|1352519|RXNORM|NASTURTIUM OFFICINALE EXTRACT|NASTURTIUM OFFICINALE EXTRACT
C0873198|T121|259525|RXNORM|APIS MELLIFERA VEN PROTEIN|APIS MELLIFERA VEN PROTEIN
C3475362|T121|1356150|RXNORM|TRIOCTYLDODECYL CITRATE|TRIOCTYLDODECYL CITRATE
C3486579|T197|1313314|RXNORM|ANTIMONY ARSENATE|ANTIMONY ARSENATE
C0717569|T121|214372|RXNORM|CHARCOAL / SIMETHICONE|CHARCOAL / SIMETHICONE
C0982374|T109|1356151|RXNORM|RICE BRAN|RICE BRAN
C1874411|T121|689625|RXNORM|BACITRACIN / LIDOCAINE / POLYMYXIN B|BACITRACIN / LIDOCAINE / POLYMYXIN B
C1874409|T121|689623|RXNORM|BACITRACIN / HYDROCORTISONE / NEOMYCIN / POLYMYXIN B|BACITRACIN / HYDROCORTISONE / NEOMYCIN / POLYMYXIN B
C1874409|T121|689623|RXNORM|BACITRACIN / HYDROCORTISONE / NEOMYCIN / POLYMYXIN B|BACITRACIN / HYDROCORTISONE / NEOMYCIN / POLYMYXIN B
C3668711|T121|1441299|RXNORM|AMANITA PHALLOIDES WHOLE EXTRACT|AMANITA PHALLOIDES WHOLE EXTRACT
C0072032|T121|34530|RXNORM|PROCATEROL|PROCATEROL
C1874414|T121|689629|RXNORM|BACITRACIN / POLYMYXIN B / PRAMOXINE|BACITRACIN / POLYMYXIN B / PRAMOXINE
C0119394|T121|50470|RXNORM|GLUCEPTATE|GLUCEPTATE
C3498054|T127|1313966|RXNORM|5-METHYLTETRAHYDROFOLIC ACID|5-METHYLTETRAHYDROFOLIC ACID
C3496683|T121|1306926|RXNORM|ALLANTOIN / PETROLATUM / ZINC OXIDE|ALLANTOIN / PETROLATUM / ZINC OXIDE
C3710164|T121|1489157|RXNORM|BENZALKONIUM / BENZYL ALCOHOL|BENZALKONIUM / BENZYL ALCOHOL
C2348066|T121|1546356|RXNORM|DABIGATRAN|DABIGATRAN
C3538243|T109|1538275|RXNORM|SCHIZOCHYTRIUM DHA OIL|ALGAL OIL
C1719979|T121|645049|RXNORM|CALCIUM CARBONATE / KAOLIN|CALCIUM CARBONATE / KAOLIN
C0071849|T121|1088591|RXNORM|PREGNA-4,17-DIENE-3,16-DIONE|PREGNA-4,17-DIENE-3,16-DIONE
C0076096|T121|37790|RXNORM|TENOXICAM|TENOXICAM
C2978280|T121|1088594|RXNORM|ASCORBIC ACID / CHROMIUM POLYNICOTINATE / NIACINAMIDE / OAT BRAN / PHYTOSTEROLS / PREGNA-4,17-DIENE-3,16-DIONE|ASCORBIC ACID / CHROMIUM POLYNICOTINATE / NIACINAMIDE / OAT BRAN / PHYTOSTEROLS / PREGNA-4,17-DIENE-3,16-DIONE
C3700879|T121|1486881|RXNORM|CEDRUS DEODARA WOOD EXTRACT|CEDRUS DEODARA WOOD EXTRACT
C0142916|T121|56513|RXNORM|SODIUM PROPIONATE|SODIUM PROPIONATE
C3643661|T121|1421450|RXNORM|BRIMONIDINE / BRINZOLAMIDE|BRIMONIDINE / BRINZOLAMIDE
C0057558|T125|22656|RXNORM|DESOGESTREL|DESOGESTREL
C2194073|T121|816243|RXNORM|BISMUTH CARBONATE / SIMETHICONE|BISMUTH CARBONATE / SIMETHICONE
C3499522|T121|1312389|RXNORM|MYRISTOYL TETRAPEPTIDE-4|MYRISTOYL TETRAPEPTIDE-4
C3499521|T121|1312388|RXNORM|MELANIN SYNTHETIC (TYROSINE, PEROXIDE)|MELANIN SYNTHETIC (TYROSINE, PEROXIDE)
C3499520|T121|1312387|RXNORM|DIMETHICONE-DIENE DIMETHICONE CROSSPOLYMER|DIMETHICONE-DIENE DIMETHICONE CROSSPOLYMER
C3651783|T121|1428416|RXNORM|ASARUM CANADENSE ROOT EXTRACT|ASARUM CANADENSE ROOT EXTRACT
C3651784|T121|1428415|RXNORM|ALNUS SERRULATA BARK EXTRACT|ALNUS SERRULATA BARK EXTRACT
C1375516|T005|1312384|RXNORM|MEASLES VIRUS PREPARATION|MEASLES VIRUS PREPARATION
C3256089|T109|1312383|RXNORM|QUERCUS ALBA EXTRACT|QUERCUS ALBA EXTRACT
C3499518|T121|1312382|RXNORM|QUERCUS RUBRA BARK EXTRACT|QUERCUS RUBRA BARK EXTRACT
C0070914|T197|1312381|RXNORM|PHOSPHORAMIDIC ACID|PHOSPHORAMIDIC ACID
C3499517|T121|1312380|RXNORM|ATROPA BELLADONNA FRUITING TOP EXTRACT|ATROPA BELLADONNA FRUITING TOP EXTRACT
C0033056|T121|8673|RXNORM|SACCHAROMYCES CEREVISIAE EXTRACT|FEPRAZONE
C3192967|T121|1148112|RXNORM|DOG HAIR EXTRACT / ENGLISH PLANTAIN POLLEN EXTRACT|DOG HAIR EXTRACT / ENGLISH PLANTAIN POLLEN EXTRACT
C0057239|T121|22380|RXNORM|DECANOIC ACID|DECANOIC ACID
C3834070|T122|1541747|RXNORM|POLYGLYCERYL-10 HEXAOLEATE|POLYGLYCERYL-10 HEXAOLEATE
C3700900|T109|1486086|RXNORM|ARNICA MONTANA FLOWER WATER|ARNICA MONTANA FLOWER WATER
C2728175|T129|973880|RXNORM|FIG ALLERGENIC EXTRACT|FICUS CARICA ALLERGENIC EXTRACT
C0046882|T121|13982|RXNORM|TIRATRICOL|TIRATRICOL
C0064906|T121|28656|RXNORM|NAFARELIN|NAFARELIN
C3538401|T116|1372682|RXNORM|POLY(N-ACETYL, N-ARGINYL)GLUCOSAMINE (50000-80000 MW)|POLY(N-ACETYL, N-ARGINYL)GLUCOSAMINE (50000-80000 MW)
C0058389|T121|23386|RXNORM|DIPHENYLPYRALINE|DIPHENYLPYRALINE
C2081462|T121|815628|RXNORM|ASCORBIC ACID / PIROXICAM|ASCORBIC ACID / PIROXICAM
C2064850|T121|818771|RXNORM|CITRIC ACID / POTASSIUM BICARBONATE / SODIUM BICARBONATE|CITRIC ACID / POTASSIUM BICARBONATE / SODIUM BICARBONATE
C0056831|T121|22033|RXNORM|CYCLOTHIAZIDE|CYCLOTHIAZIDE
C2825682|T121|1242806|RXNORM|INGENOL MEBUTATE|INGENOL MEBUTATE
C0717720|T121|214519|RXNORM|DOCUSATE / FERROUS FUMARATE|DOCUSATE / FERROUS FUMARATE
C0056835|T121|22037|RXNORM|CYCRIMINE|CYCRIMINE
C2146631|T121|816029|RXNORM|ACETAMINOPHEN / SCOPOLAMINE|ACETAMINOPHEN / SCOPOLAMINE
C0066033|T121|29584|RXNORM|MESULFEN|MESULFEN
C0717713|T121|214512|RXNORM|DIPHENHYDRAMINE / PSEUDOEPHEDRINE|DIPHENHYDRAMINE / PSEUDOEPHEDRINE
C0388753|T121|119565|RXNORM|TOLTERODINE|TOLTERODINE
C3651794|T121|1428027|RXNORM|CALENDULA OFFICINALIS WHOLE EXTRACT|CALENDULA OFFICINALIS WHOLE EXTRACT
C0246719|T121|73056|RXNORM|RISEDRONATE|RISEDRONATE
C2701689|T129|852613|RXNORM|WINTERFAT POLLEN EXTRACT|KRASCHENINNIKOVIA LANATA POLLEN EXTRACT
C2701693|T121|852617|RXNORM|KARAYA GUM EXTRACT|KARAYA GUM EXTRACT
C3486595|T121|1348450|RXNORM|AILANTHUS ALTISSIMA FLOWERING TWIG EXTRACT|AILANTHUS ALTISSIMA FLOWERING TWIG EXTRACT
C2929896|T121|1009001|RXNORM|DIHYDROXYALUMINUM SODIUM CARBONATE / SIMETHICONE|DIHYDROXYALUMINUM SODIUM CARBONATE / SIMETHICONE
C3486668|T121|1348452|RXNORM|IMPATIENS GLANDULIFERA FLOWER EXTRACT|IMPATIENS GLANDULIFERA FLOWER EXTRACT
C3464497|T121|1292422|RXNORM|VARICELLA-ZOSTER VIRUS VACCINE LIVE (OKA-MERCK) STRAIN|VARICELLA-ZOSTER VIRUS VACCINE LIVE (OKA-MERCK) STRAIN
C3486697|T121|1348454|RXNORM|ACONITUM FEROX ROOT EXTRACT|ACONITUM FEROX ROOT EXTRACT
C3488382|T121|1348455|RXNORM|TAENIA SOLIUM PREPARATION|TAENIA SOLIUM PREPARATION
C2928950|T121|1008039|RXNORM|ASCORBIC ACID / FERROUS BISGLYCINATE / POLYSACCHARIDE IRON COMPLEX|ASCORBIC ACID / FERROUS BISGLYCINATE / POLYSACCHARIDE IRON COMPLEX
C2928949|T121|1008038|RXNORM|CRANBERRY PREPARATION / EVENING PRIMROSE EXTRACT / GAMMA-LINOLENATE / LINOLEATE|CRANBERRY PREPARATION / EVENING PRIMROSE EXTRACT / GAMMA-LINOLENATE / LINOLEATE
C0101303|T122|1364500|RXNORM|ACRYLATE|ACRYLATE
C2928947|T121|1008036|RXNORM|PHENOLPHTHALEIN / SENNOSIDES, USP|PHENOLPHTHALEIN / SENNOSIDES, USP
C2928946|T121|1008035|RXNORM|CALCIUM CITRATE / CHOLECALCIFEROL / MAGNESIUM CITRATE|CALCIUM CITRATE / CHOLECALCIFEROL / MAGNESIUM CITRATE
C2928945|T121|1008034|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP A CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP C CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP W-135 CAPSUL|NEISSERIA MENINGITIDIS SEROGROUP A CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP C CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP W-135 CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP Y CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE
C2928945|T121|1008034|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP A CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP C CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP W-135 CAPSUL|NEISSERIA MENINGITIDIS SEROGROUP A CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP C CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP W-135 CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP Y CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE
C1664205|T195|1364504|RXNORM|BEDAQUILINE|BEDAQUILINE
C2928943|T121|1008032|RXNORM|MELATONIN / THEANINE|MELATONIN / THEANINE
C2928942|T121|1008031|RXNORM|CHYMOSIN / PEPSIN A|CHYMOSIN / PEPSIN A
C2928941|T121|1008030|RXNORM|DIPROPIZINE / GUAIACOL ETHYLGLYCOLATE|DIPROPIZINE / GUAIACOL ETHYLGLYCOLATE
C2347977|T121|1322046|RXNORM|ROSE PETAL EXTRACT|ROSA RUGOSA FLOWER EXTRACT
C2709752|T129|854948|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 19F VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 19F VACCINE
C0875913|T121|261407|RXNORM|BUTABARBITAL / HYOSCYAMINE / PHENAZOPYRIDINE|BUTABARBITAL / HYOSCYAMINE / PHENAZOPYRIDINE
C0040077|T123|1372538|RXNORM|THYMIDINE|DEOXYRIBOSYLTHYMINE
C0018321|T114|1372539|RXNORM|GUANINE|GUANINE
C0005011|T121|1372|RXNORM|ASCORBIC ACID / BUTCHER'S BROOM PREPARATION / CITRUS BIOFLAVONOIDS / DIOSMIN / RUTIN|BENORILATE
C0054129|T121|19768|RXNORM|BROMOPRIDE|BROMOPRIDE
C2709750|T129|854946|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 19A VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 19A VACCINE
C2081466|T121|815961|RXNORM|PIROXICAM / PREDNISONE|PIROXICAM / PREDNISONE
C2709748|T129|854944|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 18C VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 18C VACCINE
C2929899|T121|1009004|RXNORM|CETYLPYRIDINIUM / ZINC CHLORIDE|CETYLPYRIDINIUM / ZINC CHLORIDE
C0057074|T120|1310601|RXNORM|D.C. RED NO. 33|D.C. RED NO. 33
C0051510|T121|17609|RXNORM|ALUMINUM ACETATE|ALUMINUM ACETATE
C0051209|T121|17354|RXNORM|ALLOIN|ALLOIN
C2701595|T129|852479|RXNORM|HORSE SKIN EXTRACT|HORSE SKIN EXTRACT
C0007551|T195|2183|RXNORM|CEFONICID|CEFONICID
C2929904|T121|1009009|RXNORM|CLOFIBRATE / NICOTINYL ALCOHOL|CLOFIBRATE / NICOTINYL ALCOHOL
C0007546|T195|2180|RXNORM|CEFAZOLIN|CEFAZOLIN
C0007555|T195|2187|RXNORM|CEFOTETAN|CEFOTETAN
C0007554|T195|2186|RXNORM|CEFOTAXIME|CEFOTAXIME
C3255755|T121|1426457|RXNORM|ETHYL ACRYLATE AND METHYL METHACRYLATE COPOLYMER (2:1; 750000 MW)|ETHYL ACRYLATE AND METHYL METHACRYLATE COPOLYMER (2:1; 750000 MW)
C0007552|T195|2184|RXNORM|CEFOPERAZONE|CEFOPERAZONE
C3555513|T121|1375414|RXNORM|C20-40 PARETH-3|C20-40 PARETH-3
C0728747|T129|224905|RXNORM|TRASTUZUMAB|TRASTUZUMAB
C0007556|T195|2188|RXNORM|CEFOTIAM|CEFOTIAM
C0016860|T121|4603|RXNORM|FUROSEMIDE|FUROSEMIDE
C0016855|T195|4601|RXNORM|FURAZOLIDONE|FURAZOLIDONE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT,CLADOSPORIUM CLADOSPORIS|PRASTERONE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, COMMON SAGEBRUSH|PRASTERONE
C0885057|T121|265647|RXNORM|GARLIC PREPARATION|GARLIC PREPARATION
C2093618|T129|905301|RXNORM|ARABIC GUM ALLERGENIC EXTRACT|ARABIC GUM ALLERGENIC EXTRACT
C2928420|T121|1007498|RXNORM|CALCIUM CARBONATE / PSYLLIUM|CALCIUM CARBONATE / PSYLLIUM
C3700988|T121|1487171|RXNORM|LUFENURON / MILBEMYCIN OXIME|LUFENURON / MILBEMYCIN OXIME
C0071330|T121|968170|RXNORM|POLIDOCANOL|POLIDOCANOL
C0059774|T109|1546209|RXNORM|ETHYL METHYLPHENYLGLYCIDATE|ETHYL METHYLPHENYLGLYCIDATE
C0213404|T121|69036|RXNORM|RUFINAMIDE|RUFINAMIDE
C0806919|T121|257844|RXNORM|MEFENAMATE|MEFENAMATE
C0000956|T121|154|RXNORM|ACENOCOUMAROL|ACENOCOUMAROL
C3282697|T121|1252020|RXNORM|DODECYLBENZENESULFONIC ACID / HYDROGEN PEROXIDE / LACTATE|DODECYLBENZENESULFONIC ACID / HYDROGEN PEROXIDE / LACTATE
C0055445|T121|20861|RXNORM|CHLOROPYRAMINE|CHLOROPYRAMINE
C0051224|T120|1310600|RXNORM|ALLURA RED AC DYE|ALLURA RED AC DYE
C0031412|T121|8134|RXNORM|PHENOBARBITAL|PHENOBARBITAL
C0057749|T121|1310602|RXNORM|DIAZOLIDINYLUREA|DIAZOLIDINYLUREA
C0069414|T121|1310603|RXNORM|OLEYL ALCOHOL|OLEYL ALCOHOL
C0772270|T130|1310605|RXNORM|BRILLIANT BLUE FCF|BRILLIANT BLUE FCF
C0071444|T122|1424562|RXNORM|POLY(LACTIDE)|POLY(LACTIDE)
C2142865|T121|817379|RXNORM|ACETAMINOPHEN / CODEINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / CODEINE / PSEUDOEPHEDRINE
C3152849|T121|1098207|RXNORM|EUROPEAN RABBIT HAIR EXTRACT / EUROPEAN RABBIT SKIN EXTRACT|EUROPEAN RABBIT HAIR EXTRACT / EUROPEAN RABBIT SKIN EXTRACT
C0041037|T121|10826|RXNORM|TRIMETAZIDINE|TRIMETAZIDINE
C1445178|T129|1192987|RXNORM|PARAKEET FEATHER ALLERGENIC EXTRACT|MELOPSITTACUS UNDULATUS FEATHER ALLERGENIC EXTRACT
C3818788|T109|1491737|RXNORM|ELAEIS OLEIFERA SEED OIL|ELAEIS OLEIFERA SEED OIL
C3282703|T121|1252026|RXNORM|HEPTANOIC ACID / IODINE|HEPTANOIC ACID / IODINE
C1562545|T121|597501|RXNORM|DESLORATADINE / PSEUDOEPHEDRINE|DESLORATADINE / PSEUDOEPHEDRINE
C2928413|T121|1007491|RXNORM|PHENYLBUTAZONE / SALICYLAMIDE|PHENYLBUTAZONE / SALICYLAMIDE
C2929677|T121|1008778|RXNORM|GLYCERIN / PARAFFIN|GLYCERIN / PARAFFIN
C0022860|T121|6185|RXNORM|LABETALOL|LABETALOL
C1874366|T121|689516|RXNORM|ASPIRIN / CAFFEINE / IPECAC / OPIUM|ASPIRIN / CAFFEINE / IPECAC / OPIUM
C0031408|T121|8132|RXNORM|PHENIRAMINE|PHENIRAMINE
C3153291|T121|1098874|RXNORM|DOCOSAHEXAENOATE / PHOSPHATIDYLSERINE|DOCOSAHEXAENOATE / PHOSPHATIDYLSERINE
C2701557|T129|852386|RXNORM|EUCALYPTUS GLOBULUS POLLEN EXTRACT|EUCALYPTUS GLOBULUS POLLEN EXTRACT
C1572554|T121|485876|RXNORM|BETA SITOSTEROL / ZINC CITRATE|BETA SITOSTEROL / ZINC CITRATE
C2928415|T121|1007493|RXNORM|ENTEROCOCCUS FAECALIS / ESCHERICHIA COLI|ENTEROCOCCUS FAECALIS / ESCHERICHIA COLI
C0085149|T121|42316|RXNORM|TACROLIMUS|TACROLIMUS
C0085149|T121|42316|RXNORM|TACROLIMUS|TACROLIMUS
C0528166|T121|135775|RXNORM|ZOLMITRIPTAN|ZOLMITRIPTAN
C1874363|T121|689513|RXNORM|ASPIRIN / CAFFEINE / DIHYDROCODEINE / PROMETHAZINE|ASPIRIN / CAFFEINE / DIHYDROCODEINE / PROMETHAZINE
C0300205|T121|1005921|RXNORM|ULIPRISTAL|ULIPRISTAL
C0110038|T195|48203|RXNORM|CLAVULANATE|CLAVULANATE
C3857946|T121|1552449|RXNORM|BOS TAURUS LIGAMENT PREPARATION|BOS TAURUS LIGAMENT PREPARATION
C2927383|T129|1005929|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-CALIFORNIA-07-2009 X-179A (H1N1) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-CALIFORNIA-07-2009 X-179A (H1N1) STRAIN
C0027329|T121|7236|RXNORM|NAFRONYL|NAFRONYL
C0982304|T129|314753|RXNORM|ORRIS ALLERGENIC EXTRACT|ORRIS ALLERGENIC EXTRACT
C3663000|T122|1432298|RXNORM|OLEYL ERUCATE|OLEYL ERUCATE
C2343876|T168|1432299|RXNORM|POPPY SEED OIL|POPPY SEED OIL
C2194285|T121|812823|RXNORM|CLOBUTINOL / METAPROTERENOL|CLOBUTINOL / METAPROTERENOL
C0027324|T195|7233|RXNORM|NAFCILLIN|NAFCILLIN
C0039600|T125|10378|RXNORM|TESTOLACTONE|TESTOLACTONE
C0039601|T125|10379|RXNORM|TESTOSTERONE|TESTOSTERONE
C3662996|T121|1432292|RXNORM|ELAEIS GUINEENSIS FRUIT EXTRACT|ELAEIS GUINEENSIS FRUIT EXTRACT
C2987605|T129|1432293|RXNORM|DALOTUZUMAB|DALOTUZUMAB
C3500809|T121|1356107|RXNORM|BENZALKONIUM / HEXYLRESORCINOL / ZINC CHLORIDE|BENZALKONIUM / HEXYLRESORCINOL / ZINC CHLORIDE
C3500803|T121|1356101|RXNORM|ALLANTOIN / CAMPHOR / HEXYLRESORCINOL / MENTHOL|ALLANTOIN / CAMPHOR / HEXYLRESORCINOL / MENTHOL
C3662999|T109|1432297|RXNORM|GLYCERYL CITRATE|MONOGLYCERIDE CITRATE
C0027348|T121|7238|RXNORM|NALBUPHINE|NALBUPHINE
C3662997|T121|1432295|RXNORM|CITRONELLOL ACETATE, (R)-|CITRONELLOL ACETATE, (R)-
C2927886|T121|1006963|RXNORM|NEOSTIGMINE / PILOCARPINE|NEOSTIGMINE / PILOCARPINE
C2927884|T121|1006961|RXNORM|ALLANTOIN / ICHTHAMMOL|ALLANTOIN / ICHTHAMMOL
C2927883|T121|1006960|RXNORM|MEFRUSIDE / RESERPINE|MEFRUSIDE / RESERPINE
C2927890|T121|1006967|RXNORM|MAGNESIUM OXIDE / MAGNESIUM SULFATE|MAGNESIUM OXIDE / MAGNESIUM SULFATE
C2927889|T121|1006966|RXNORM|LIDOCAINE / METHYLBENZETHONIUM|LIDOCAINE / METHYLBENZETHONIUM
C2927888|T121|1006965|RXNORM|BETA CAROTENE / VITAMIN E|BETA CAROTENE / VITAMIN E
C2927887|T121|1006964|RXNORM|MAGNESIUM GLUCONATE / POTASSIUM TARTRATE|MAGNESIUM GLUCONATE / POTASSIUM TARTRATE
C2702420|T129|1294630|RXNORM|METRICUS PAPER WASP VENOM PROTEIN|POLISTES METRICUS VENOM
C2927892|T121|1006969|RXNORM|CALCIUM GLUCONATE / CALCIUM LEVULINATE|CALCIUM GLUCONATE / CALCIUM LEVULINATE
C2927891|T121|1006968|RXNORM|CYSTEINE / METHIONINE|CYSTEINE / METHIONINE
C0133860|T123|1495153|RXNORM|FATTY ACIDS, OMEGA-6|FATTY ACIDS, OMEGA-6
C0051839|T121|17881|RXNORM|ANETHOLE|ANETHOLE
C2929973|T121|1009078|RXNORM|DIPYRONE / TROSPIUM|DIPYRONE / TROSPIUM
C2929974|T121|1009079|RXNORM|IDEBENONE / NIMODIPINE|IDEBENONE / NIMODIPINE
C3668770|T121|1441397|RXNORM|ASCORBIC ACID / COLLAGEN|ASCORBIC ACID / COLLAGEN
C3668765|T121|1441391|RXNORM|BAZEDOXIFENE / ESTROGENS, CONJUGATED (USP)|BAZEDOXIFENE / ESTROGENS, CONJUGATED (USP)
C2929965|T121|1009070|RXNORM|ALOE EXTRACT / PHENOLPHTHALEIN|ALOE EXTRACT / PHENOLPHTHALEIN
C2929966|T121|1009071|RXNORM|CYCLANDELATE / ETOFYLLINE|CYCLANDELATE / ETOFYLLINE
C2929967|T121|1009072|RXNORM|GLUCOSE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE|GLUCOSE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE
C1145701|T195|236594|RXNORM|AMPHOTERICIN B LIPOSOMAL|AMPHOTERICIN B LIPOSOMAL
C2929969|T121|1009074|RXNORM|AMMONIUM CHLORIDE / LICORICE ROOT EXTRACT|AMMONIUM CHLORIDE / LICORICE ROOT EXTRACT
C2929970|T121|1009075|RXNORM|HYDROCORTISONE / ZINC SULFATE|HYDROCORTISONE / ZINC SULFATE
C2929971|T121|1009076|RXNORM|CHLORDIAZEPOXIDE / PENTAERYTHRITOL|CHLORDIAZEPOXIDE / PENTAERYTHRITOL
C2929972|T121|1009077|RXNORM|PETROLATUM / ZINC OXIDE|PETROLATUM / ZINC OXIDE
C1874818|T121|689396|RXNORM|CHLORPHENIRAMINE / EPHEDRINE / GUAIFENESIN / PHENOBARBITAL / THEOPHYLLINE|CHLORPHENIRAMINE / EPHEDRINE / GUAIFENESIN / PHENOBARBITAL / THEOPHYLLINE
C1874817|T121|689395|RXNORM|CHLORPHENIRAMINE / EPHEDRINE / GUAIFENESIN / HYDROIODIC ACID|CHLORPHENIRAMINE / EPHEDRINE / GUAIFENESIN / HYDROIODIC ACID
C2742627|T121|689394|RXNORM|CHLORPHENIRAMINE / EPHEDRINE|CHLORPHENIRAMINE / EPHEDRINE
C1874814|T121|689391|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE
C3644810|T121|1425901|RXNORM|APHLOIA THEIFORMIS LEAF EXTRACT|APHLOIA THEIFORMIS LEAF EXTRACT
C0030073|T121|7814|RXNORM|OXYMORPHONE|OXYMORPHONE
C3256283|T109|1425909|RXNORM|CAPRYLIC-CAPRIC DIGLYCEROL SUCCINATE|CAPRYLIC-CAPRIC DIGLYCEROL SUCCINATE
C0036228|T123|1362906|RXNORM|SARCOSINE|SARCOSINE
C0053296|T109|1362907|RXNORM|BENZYL SALICYLATE|BENZYL SALICYLATE
C0017984|T123|1362904|RXNORM|GLYCYLGLYCINE|GLYCYLGLYCINE
C0034632|T109|1362905|RXNORM|RAFFINOSE|RAFFINOSE
C0012456|T130|1362902|RXNORM|DIMYRISTOYLPHOSPHATIDYLCHOLINE|DIMYRISTOYLPHOSPHATIDYLCHOLINE
C0015637|T121|1362903|RXNORM|FARNESOL|FARNESOL
C0006506|T131|1362900|RXNORM|BUTYLATED HYDROXYANISOLE|BUTYLATED HYDROXYANISOLE
C0006716|T197|1362901|RXNORM|CALCIUM PYROPHOSPHATE|CALCIUM PYROPHOSPHATE
C0037107|T196|9774|RXNORM|SILICON|SILICON
C0039955|T121|10510|RXNORM|THIOTHIXENE|THIOTHIXENE
C0037098|T197|9771|RXNORM|SILICON DIOXIDE|SILICON DIOXIDE
C0039962|T131|10517|RXNORM|THIRAM|THIRAM
C0054273|T121|1362908|RXNORM|BUTYL ACETATE|BUTYL ACETATE
C0054720|T122|1362909|RXNORM|CARBOMER-940|CARBOMER-940
C0048197|T121|14982|RXNORM|PARACHLOROPHENOL|PARACHLOROPHENOL
C0076681|T195|38278|RXNORM|TILMICOSIN|TILMICOSIN
C0022942|T123|1425933|RXNORM|LACTOFERRIN|LACTOFERRIN
C0056077|T123|21406|RXNORM|COENZYME Q10|COENZYME Q10
C3497034|T121|1308407|RXNORM|ALCLOXA / CHLOROXYLENOL|ALCLOXA / CHLOROXYLENOL
C3541367|T121|1433212|RXNORM|LEVOMILNACIPRAN|LEVOMILNACIPRAN
C3668630|T121|1441178|RXNORM|ALLANTOIN / ZINC OXIDE|ALLANTOIN / ZINC OXIDE
C2731513|T129|895503|RXNORM|DOMESTIC GOAT HAIR EXTRACT|CAPRA HIRCUS HAIR EXTRACT
C0666079|T121|191566|RXNORM|CLIMBAZOLE|CLIMBAZOLE
C2702399|T129|895507|RXNORM|GUINEA PIG HAIR EXTRACT|CAVIA PORCELLUS HAIR EXTRACT
C2929768|T121|1008870|RXNORM|ECHINACEA PURPUREA EXTRACT / EUCALYPTUS OIL / MENTHOL|ECHINACEA PURPUREA EXTRACT / EUCALYPTUS OIL / MENTHOL
C2985211|T121|1368879|RXNORM|ISOPROPYLPARABEN|ISOPROPYLPARABEN
C1636150|T121|608253|RXNORM|BETAMETHASONE / NEOMYCIN|BETAMETHASONE / NEOMYCIN
C0078792|T121|39952|RXNORM|ZINC PYRITHIONE|ZINC PYRITHIONE
C2741547|T129|901390|RXNORM|COMMON CARP ALLERGENIC EXTRACT|CYPRINUS CARPIO ALLERGENIC EXTRACT
C3464060|T121|1427229|RXNORM|HYDROLYSED MARINE COLLAGEN (ENZYMATIC; 2000 MW)|HYDROLYSED MARINE COLLAGEN (ENZYMATIC; 2000 MW)
C0030082|T121|7818|RXNORM|OXYPHENONIUM|OXYPHENONIUM
C2742211|T109|1427225|RXNORM|FLORBETAPIR|FLORBETAPIR
C3472775|T122|1427227|RXNORM|PPG-1 TRIDECETH-6|PPG-1 TRIDECETH-6
C3473983|T121|1427226|RXNORM|ISOPROPYL LAUROYL SARCOSINATE|ISOPROPYL LAUROYL SARCOSINATE
C3465213|T121|1427221|RXNORM|SARDINE, UNSPECIFIED PREPARATION|SARDINE, UNSPECIFIED PREPARATION
C3465039|T109|1427220|RXNORM|PICHIA JADINII EXTRACT|CYBERLINDNERA JADINII EXTRACT
C0030520|T125|1427222|RXNORM|PARATHYROID HORMONE|PARATHYROID HORMONE
C0006020|T197|1700|RXNORM|BORIC ACID|HYDROGEN BORATE
C0006020|T197|1700|RXNORM|BORIC ACID|HYDROGEN BORATE
C0006020|T197|1700|RXNORM|BORIC ACID|HYDROGEN BORATE
C0025698|T121|1305751|RXNORM|METHYL CHLORIDE|METHYL CHLORIDE
C3667709|T121|1439947|RXNORM|ACETIC ACID / CHLORHEXIDINE / KETOCONAZOLE|ACETIC ACID / CHLORHEXIDINE / KETOCONAZOLE
C0006030|T196|1705|RXNORM|BORON|BORON
C2826072|T121|1305758|RXNORM|POVIDONE K29-32|POVIDONE K29-32
C1572787|T121|1314380|RXNORM|POLOXAMER 182|POLOXAMER 182
C1364953|T121|1314382|RXNORM|POLYETHYLENE GLYCOL 1500|POLYETHYLENE GLYCOL 1500
C0141951|T121|1314385|RXNORM|SEMDURAMICIN|SEMDURAMICIN
C0030775|T121|1314384|RXNORM|POLYETHYLENE GLYCOL 6000|POLYETHYLENE GLYCOL 6000
C3255607|T109|1314386|RXNORM|PSEUDOPTEROGORGIA ELISABETHAE EXTRACT|PSEUDOPTEROGORGIA ELISABETHAE EXTRACT
C3848574|T196|1546270|RXNORM|RADIUM CATION|RADIUM CATION
C0026560|T121|1368870|RXNORM|MORPHOLINE|MORPHOLINE
C2347051|T197|1546272|RXNORM|MANGANESE CATION (2+)|MANGANESE CATION (2+)
C3848572|T196|1546273|RXNORM|FLUORIDE ION F-18|FLUORIDE ION F-18
C3848571|T196|1546274|RXNORM|BROMIDE ION|BROMIDE ION
C3848570|T196|1546275|RXNORM|IODIDE ION|IODIDE ION
C3282699|T121|1355818|RXNORM|RANUNCULUS FICARIA EXTRACT|RANUNCULUS FICARIA EXTRACT
C0040087|T123|1368871|RXNORM|THYMINE|THYMINE
C3848568|T196|1546278|RXNORM|STRONTIUM CATION|STRONTIUM CATION
C2713885|T109|1546279|RXNORM|OSELTAMIVIR CARBOXYLATE|OSELTAMIVIR CARBOXYLATE
C0009063|T007|1318475|RXNORM|CLOSTRIDIUM PERFRINGENS|CLOSTRIDIUM PERFRINGENS
C2080536|T121|814051|RXNORM|NOSCAPINE / PHENYLEPHRINE|NOSCAPINE / PHENYLEPHRINE
C0008151|T007|1318474|RXNORM|CHLAMYDIA TRACHOMATIS|CHLAMYDIA TRACHOMATIS
C3834085|T197|1541729|RXNORM|MAMMAL BONE, FOSSILIZED|MAMMAL BONE, FOSSILIZED
C3834086|T109|1541728|RXNORM|ERUCA VESICARIA SUBSP. SATIVA LEAF EXTRACT|ERUCA VESICARIA SUBSP. SATIVA LEAF EXTRACT
C3834087|T109|1541727|RXNORM|BRASSICA OLERACEA VAR. ITALICA WHOLE EXTRACT|BRASSICA OLERACEA VAR. ITALICA WHOLE EXTRACT
C0058243|T130|1368874|RXNORM|DIMETHYLACETAMIDE|N,N-DIMETHYLACETAMIDE
C0879427|T129|263034|RXNORM|PANITUMUMAB|PANITUMUMAB
C3834090|T109|1541724|RXNORM|TRITICUM POLONICUM SEED EXTRACT|TRITICUM POLONICUM SEED EXTRACT
C3834091|T109|1541723|RXNORM|PINUS DENSIFLORA LEAF EXTRACT|PINUS DENSIFLORA LEAF EXTRACT
C3834092|T109|1541722|RXNORM|LAWSONIA INERMIS WHOLE EXTRACT|LAWSONIA INERMIS WHOLE EXTRACT
C3714981|T122|1541721|RXNORM|SESAMUM INDICUM WHOLE EXTRACT|SESAMUM INDICUM WHOLE EXTRACT
C0061223|T121|1368875|RXNORM|GERANIOL|GERANIOL
C0133689|T121|54034|RXNORM|OCTOXYNOL-9|OCTOXYNOL-9
C0002268|T126|259351|RXNORM|ALPHA-D-GALACTOSIDASE ENZYME|ALPHA-D-GALACTOSIDASE ENZYME
C0033399|T121|8742|RXNORM|PROMAZINE|PROMAZINE
C0061300|T121|1368876|RXNORM|GLAUCINE|GLAUCINE
C0042338|T005|11131|RXNORM|HUMAN HERPESVIRUS 3|HUMAN HERPESVIRUS 3
C0006305|T007|1318470|RXNORM|BRUCELLA MELITENSIS|BRUCELLA MELITENSIS
C0073371|T195|35616|RXNORM|RIFAMYCIN SV|RIFAMYCIN
C2194314|T121|815452|RXNORM|CLONIXIN / CYPROHEPTADINE / ERGOTAMINE|CLONIXIN / CYPROHEPTADINE / ERGOTAMINE
C0010654|T123|3024|RXNORM|CYSTEINE|CYSTEINE
C0010648|T121|3022|RXNORM|CYSTEAMINE|CYSTEAMINE
C0010648|T121|3022|RXNORM|CYSTEAMINE|CYSTEAMINE
C0010648|T121|3022|RXNORM|CYSTEAMINE|CYSTEAMINE
C3499830|T121|1312979|RXNORM|CHOLECALCIFEROL / POLYSACCHARIDE IRON COMPLEX|CHOLECALCIFEROL / POLYSACCHARIDE IRON COMPLEX
C0063123|T121|1312602|RXNORM|HYDROXYCITRIC ACID|HYDROXYCITRIC ACID
C0770967|T121|1312975|RXNORM|AMMONIUM STEARATE|AMMONIUM STEARATE
C3474468|T121|1312600|RXNORM|HYDROLYSED BOVINE COLLAGEN (ENZYMATIC; 2000-5000 MW)|HYDROLYSED BOVINE COLLAGEN (ENZYMATIC; 2000-5000 MW)
C3257697|T121|1312601|RXNORM|HYDROLYZED ELASTIN, BOVINE, ALKALINE (1000 MW)|HYDROLYZED ELASTIN, BOVINE, ALKALINE (1000 MW)
C3484464|T121|1334747|RXNORM|FUCUS VESICULOSUS EXTRACT|BLADDERWRACK EXTRACT
C0071778|T197|34322|RXNORM|POTASSIUM PHOSPHATE|POTASSIUM PHOSPHATE
C0033321|T121|8730|RXNORM|PROGLUMIDE|PROGLUMIDE
C3700400|T121|1486436|RXNORM|DAPAGLIFLOZIN / METFORMIN|DAPAGLIFLOZIN / METFORMIN
C0068475|T121|31555|RXNORM|NEBIVOLOL|NEBIVOLOL
C0067794|T123|31005|RXNORM|N-ACETYLTYROSINE|N-ACETYLTYROSINE
C3485056|T131|1310456|RXNORM|CROTALUS HORRIDUS HORRIDUS VENOM|CROTALUS HORRIDUS HORRIDUS VENOM
C0015205|T130|4191|RXNORM|EVANS BLUE|EVANS BLUE
C0053838|T121|1310459|RXNORM|BLACK WIDOW SPIDER VENOM|LATRODECTUS MACTANS VENOM
C0205996|T195|66958|RXNORM|PRISTINAMYCIN|PRISTINAMYCIN
C0120077|T121|50598|RXNORM|GOLD KERATINATE|GOLD KERATINATE
C3489013|T123|1310458|RXNORM|LACHESIS MUTA VENOM|LACHESIS MUTA VENOM
C0071968|T121|34479|RXNORM|PRIDINOL|PRIDINOL
C2928700|T121|1007785|RXNORM|FENTANYL / SODIUM CHLORIDE|FENTANYL / SODIUM CHLORIDE
C2928701|T121|1007786|RXNORM|ERGOLOID MESYLATES, USP / FLUNARIZINE|ERGOLOID MESYLATES, USP / FLUNARIZINE
C2928702|T121|1007787|RXNORM|BELLADONNA EXTRACT, USP / METHENAMINE / SALICYLAMIDE|BELLADONNA EXTRACT, USP / METHENAMINE / SALICYLAMIDE
C2928695|T121|1007780|RXNORM|COENZYME Q10 / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / VITAMIN E|COENZYME Q10 / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / VITAMIN E
C0304520|T121|91235|RXNORM|DIGITALIS PREPARATION|DIGITALIS PREPARATION
C2928697|T121|1007782|RXNORM|ASCORBIC ACID / DOCOSAHEXAENOATE / LUTEIN|ASCORBIC ACID / DOCOSAHEXAENOATE / LUTEIN
C2928698|T121|1007783|RXNORM|FLUDROCORTISONE / HEXAMIDINE / SELENIUM SULFIDE|FLUDROCORTISONE / HEXAMIDINE / SELENIUM SULFIDE
C0076808|T121|38386|RXNORM|TOLRESTAT|TOLRESTAT
C2928703|T121|1007788|RXNORM|BENZALKONIUM / GLYCERIN|BENZALKONIUM / GLYCERIN
C2928704|T121|1007789|RXNORM|GLYCERIN / THYMOL|GLYCERIN / THYMOL
C0076804|T121|38382|RXNORM|TOLOXATONE|TOLOXATONE
C0071626|T121|34188|RXNORM|POLYNOXYLIN|POLYNOXYLIN
C2607686|T197|1426938|RXNORM|TETRAARSENIC TETRASULFIDE|TETRAARSENIC TETRASULFIDE
C3282456|T121|1426939|RXNORM|PEG-PPG-20-15 DIMETHICONE|PEG-PPG-20-15 DIMETHICONE
C1619966|T121|614391|RXNORM|ABATACEPT|ABATACEPT
C3282783|T121|1426937|RXNORM|LAURYL AMINOPROPYLGLYCINE|LAURYL AMINOPROPYLGLYCINE
C0668557|T121|1426934|RXNORM|SCLAREOLIDE|SCLAREOLIDE
C3281456|T121|1426935|RXNORM|PEG-10 GLYCERYL STEARATE|PEG-10 GLYCERYL STEARATE
C1509560|T121|476818|RXNORM|MAGNESIUM GLYCINATE|MAGNESIUM GLYCINATE
C0043850|T123|1426933|RXNORM|1,2-DISTEAROYLLECITHIN|1,2-DISTEAROYLLECITHIN
C0062921|T109|1426930|RXNORM|HOMARINE|HOMARINE
C0590743|T121|151195|RXNORM|ATENOLOL / CHLORTHALIDONE|ATENOLOL / CHLORTHALIDONE
C0590742|T121|151194|RXNORM|HYDROFLUMETHIAZIDE / SPIRONOLACTONE|HYDROFLUMETHIAZIDE / SPIRONOLACTONE
C2936929|T121|151196|RXNORM|ACETAMINOPHEN / DIHYDROCODEINE|ACETAMINOPHEN / DIHYDROCODEINE
C3556192|T121|1420991|RXNORM|ALLANTOIN / DIPHENHYDRAMINE|ALLANTOIN / DIPHENHYDRAMINE
C1700683|T121|616739|RXNORM|ROTIGOTINE|ROTIGOTINE
C0070824|T130|33504|RXNORM|PHOSPHOCELLULOSE|PHOSPHOCELLULOSE
C3818701|T122|1535932|RXNORM|AMODIMETHICONE (1300 CST)|AMODIMETHICONE (1300 CST)
C0031977|T121|8351|RXNORM|PIRACETAM|PIRACETAM
C0939799|T121|285151|RXNORM|CONIUM MACULATUM PREPARATION|CONIUM MACULATUM PREPARATION
C0058231|T121|23247|RXNORM|METHYLSULFONYLMETHANE|METHYLSULFONYLMETHANE
C1874688|T121|691179|RXNORM|CAMPHOR / EUCALYPTUS OIL / MENTHOL / METHYL SALICYLATE|CAMPHOR / EUCALYPTUS OIL / MENTHOL / METHYL SALICYLATE
C0529572|T130|136300|RXNORM|CAPROMAB PENDETIDE|CAPROMAB PENDETIDE
C0023831|T123|6436|RXNORM|LIPOTROPIC AGENTS|LIPOTROPIC AGENTS
C2728180|T129|1011043|RXNORM|HORSERADISH ALLERGENIC EXTRACT|HORSERADISH ALLERGENIC EXTRACT
C0031566|T130|8196|RXNORM|PHLOROGLUCINOL|PHLOROGLUCINOL
C2928360|T121|1007438|RXNORM|NIACINAMIDE / PROTHIONAMIDE|NIACINAMIDE / PROTHIONAMIDE
C2928361|T121|1007439|RXNORM|COENZYME Q10 / RIBOFLAVIN|COENZYME Q10 / RIBOFLAVIN
C2928358|T121|1007436|RXNORM|FLUOCORTIN BUTYL ESTER / ISOCONAZOLE|FLUOCORTIN BUTYL ESTER / ISOCONAZOLE
C2928359|T121|1007437|RXNORM|ANTIPYRINE / CAFFEINE / QUININE|ANTIPYRINE / CAFFEINE / QUININE
C2928356|T121|1007434|RXNORM|AMYLOCAINE / LINDANE|AMYLOCAINE / LINDANE
C3152894|T121|1098264|RXNORM|RED OAK POLLEN EXTRACT / WHITE OAK POLLEN EXTRACT|RED OAK POLLEN EXTRACT / WHITE OAK POLLEN EXTRACT
C0795623|T129|253174|RXNORM|HEPATITIS A VACCINE, INACTIVATED|HEPATITIS A VACCINE, INACTIVATED
C2928355|T121|1007433|RXNORM|COAL TAR / FLUMETHASONE / SALICYLIC ACID|COAL TAR / FLUMETHASONE / SALICYLIC ACID
C2928352|T121|1007430|RXNORM|ETHACRIDINE / LIDOCAINE|ETHACRIDINE / LIDOCAINE
C2928353|T121|1007431|RXNORM|SODIUM CHLORIDE / UREA|SODIUM CHLORIDE / UREA
C0078049|T129|39385|RXNORM|VARICELLA-ZOSTER IMMUNE GLOBULIN|HUMAN VARICELLA-ZOSTER IMMUNE GLOBULIN
C1874674|T121|691038|RXNORM|CALCIUM UNDECYLENATE / ZINC UNDECYLENATE|CALCIUM UNDECYLENATE / ZINC UNDECYLENATE
C1169997|T121|352372|RXNORM|DEXMETHYLPHENIDATE|DEXMETHYLPHENIDATE
C1169995|T121|352370|RXNORM|DEXCHLORPHENIRAMINE / PSEUDOEPHEDRINE|DEXCHLORPHENIRAMINE / PSEUDOEPHEDRINE
C2928956|T121|1008045|RXNORM|BELLADONNA EXTRACT, USP / PHENOBARBITAL|BELLADONNA EXTRACT, USP / PHENOBARBITAL
C1170002|T121|352376|RXNORM|ETHINYL ESTRADIOL / ETONOGESTREL|ETHINYL ESTRADIOL / ETONOGESTREL
C1170003|T121|352377|RXNORM|ETHINYL ESTRADIOL / NORELGESTROMIN|ETHINYL ESTRADIOL / NORELGESTROMIN
C1170000|T121|352374|RXNORM|DROTRECOGIN ALFA|DROTRECOGIN ALFA
C1170001|T121|352375|RXNORM|EPROSARTAN / HYDROCHLOROTHIAZIDE|EPROSARTAN / HYDROCHLOROTHIAZIDE
C3485470|T121|1307102|RXNORM|ALLYL SUCROSE|ALLYL SUCROSE
C0939808|T121|285159|RXNORM|PASSION FLOWER EXTRACT|PASSION FLOWER EXTRACT
C3255231|T121|1236450|RXNORM|CHLOPHEDIANOL / CHLORCYCLIZINE|CHLOPHEDIANOL / CHLORCYCLIZINE
C1827938|T121|687148|RXNORM|COAL TAR / LECITHIN|COAL TAR / LECITHIN
C1828401|T121|687144|RXNORM|CLINDAMYCIN / TRETINOIN|CLINDAMYCIN / TRETINOIN
C0220918|T121|1307106|RXNORM|SUCCINATE|SUCCINATE
C0025382|T121|6758|RXNORM|MEPHOBARBITAL|MEPHOBARBITAL
C0025384|T121|6759|RXNORM|MEPIVACAINE|MEPIVACAINE
C3665263|T121|1435638|RXNORM|STROPHANTHUS GRATUS SEED EXTRACT|STROPHANTHUS GRATUS SEED EXTRACT
C0028127|T121|7441|RXNORM|NITRENDIPINE|NITRENDIPINE
C0025368|T121|6750|RXNORM|MENTHOL|MENTHOL
C0025368|T121|6750|RXNORM|MENTHOL|MENTHOL
C0025368|T121|6750|RXNORM|MENTHOL|MENTHOL
C0025368|T121|6750|RXNORM|MENTHOL|MENTHOL
C0025380|T121|6756|RXNORM|MEPHENTERMINE|MEPHENTERMINE
C0025381|T121|6757|RXNORM|MEPHENYTOIN|MEPHENYTOIN
C0025376|T121|6754|RXNORM|MEPERIDINE|MEPERIDINE
C0025379|T121|6755|RXNORM|MEPHENESIN|MEPHENESIN
C3496935|T109|1313735|RXNORM|BEHENETH-25|BEHENETH-25
C3497835|T121|1313734|RXNORM|ARISAEMA DRACONTIUM ROOT EXTRACT|ARISAEMA DRACONTIUM ROOT EXTRACT
C2348056|T130|1313737|RXNORM|D&C BROWN NO. 1|D&C BROWN NO. 1
C2928118|T121|1007196|RXNORM|PANTOTHENIC ACID / THIOPHENE|PANTOTHENIC ACID / THIOPHENE
C3265001|T121|1313731|RXNORM|1-EICOSENE|1-EICOSENE
C0037707|T121|9947|RXNORM|SOTALOL|SOTALOL
C0724511|T007|221050|RXNORM|BCG, LIVE, TICE STRAIN|BCG, LIVE, TICE STRAIN
C0037688|T121|9945|RXNORM|SORBITOL|SORBITOL
C0037688|T121|9945|RXNORM|SORBITOL|SORBITOL
C2701474|T129|852281|RXNORM|HAZELNUT POLLEN EXTRACT|CORYLUS AMERICANA POLLEN EXTRACT
C0037732|T168|9949|RXNORM|SOYBEAN OIL|SOYBEAN OIL
C3465011|T122|1313739|RXNORM|DIETHYLENE GLYCOL ADIPATE|DIETHYLENE GLYCOL ADIPATE
C3256908|T121|1313738|RXNORM|DECYLOXAZOLIDINONE|DECYLOXAZOLIDINONE
C0893383|T197|272758|RXNORM|GALLIUM 67 CITRATE|GALLIUM (67GA) CITRATE
C0053289|T131|19044|RXNORM|BENZYL BENZOATE|BENZYL BENZOATE
C0028126|T121|7440|RXNORM|NITRAZEPAM|NITRAZEPAM
C3486396|T121|1355184|RXNORM|COLCHICUM AUTUMNALE BULB EXTRACT|COLCHICUM AUTUMNALE BULB EXTRACT
C1302022|T121|392483|RXNORM|BENZOYL PEROXIDE / SULFUR|BENZOYL PEROXIDE / SULFUR
C3855877|T121|1549225|RXNORM|IMPATIENS BALSAMINA FLOWER EXTRACT|IMPATIENS BALSAMINA FLOWER EXTRACT
C0991869|T121|1427008|RXNORM|PROPYLENE GLYCOL DIACETATE|PROPYLENE GLYCOL DIACETATE
C0717339|T121|214160|RXNORM|ASPIRIN / BUTALBITAL / CAFFEINE / CODEINE|ASPIRIN / BUTALBITAL / CAFFEINE / CODEINE
C0086605|T127|42781|RXNORM|VITAMIN K 2|VITAMIN K 2
C0001134|T197|236|RXNORM|ACIDULATED PHOSPHATE FLUORIDE|ACIDULATED PHOSPHATE FLUORIDE
C1370128|T123|618453|RXNORM|GAMMA-LINOLENATE|GAMMA-LINOLENATE
C3256397|T109|1306124|RXNORM|ALPHA, ALPHA-DIMETHYLBENZYL ALCOHOL|ALPHA, ALPHA-DIMETHYLBENZYL ALCOHOL
C2827077|T126|1306125|RXNORM|ALPHA-AMYLASE A TYPE 1-2|ALPHA-AMYLASE A TYPE 1-2
C2980836|T129|1306122|RXNORM|MYCOGONE NIGRA ALLERGENIC EXTRACT|MYCOGONE NIGRA ALLERGENIC EXTRACT
C3191342|T121|1306120|RXNORM|PLATYCLADUS ORIENTALIS SEED EXTRACT|PLATYCLADUS ORIENTALIS SEED EXTRACT
C2825121|T121|1306128|RXNORM|ALOE VERA LEAF EXTRACT|ALOE VERA LEAF EXTRACT
C0063986|T121|27929|RXNORM|LANATOSIDE C|LANATOSIDE C
C2747077|T129|904815|RXNORM|WHITE SEEDLESS GRAPE ALLERGENIC EXTRACT|WHITE SEEDLESS GRAPE ALLERGENIC EXTRACT
C0050846|T130|17050|RXNORM|ADIPIC ACID|ADIPIC ACID
C0048070|T109|1426595|RXNORM|4-ANISIC ACID|P-ANISIC ACID
C3255855|T109|1426596|RXNORM|PALMITOYL PENTAPEPTIDE-4|PALMITOYL PENTAPEPTIDE-3
C3536965|T196|1426598|RXNORM|SULFATE ION|SULFATE ION
C0072487|T121|1362689|RXNORM|PROTOCATECHUALDEHYDE|PROTOCATECHUALDEHYDE
C0056643|T121|21877|RXNORM|CYAMEMAZINE|CYAMEMAZINE
C0015041|T121|1314353|RXNORM|ETHOPABATE|ETHOPABATE
C0041196|T109|1368873|RXNORM|TROPOLONE|TROPOLONE
C0075333|T197|37175|RXNORM|STRONTIUM CHLORIDE|STRONTIUM CHLORIDE
C0063828|T130|27792|RXNORM|IOVERSOL|IOVERSOL
C2741523|T129|901351|RXNORM|FLAXSEED ALLERGENIC EXTRACT|LINUM USITATISSIMUM ALLERGENIC EXTRACT
C1874618|T121|690812|RXNORM|BROMPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE|BROMPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C1874619|T121|690813|RXNORM|BROMPHENIRAMINE / PHENYLEPHRINE / PHENYLTOLOXAMINE|BROMPHENIRAMINE / PHENYLEPHRINE / PHENYLTOLOXAMINE
C1948068|T121|1543543|RXNORM|BELINOSTAT|BELINOSTAT
C1874617|T121|690811|RXNORM|BROMPHENIRAMINE / GUAIFENESIN / PSEUDOEPHEDRINE|BROMPHENIRAMINE / GUAIFENESIN / PSEUDOEPHEDRINE
C3666505|T121|1437220|RXNORM|BETULA PUBESCENS FLOWER BUD EXTRACT|BETULA PUBESCENS FLOWER BUD EXTRACT
C0030637|T007|1437221|RXNORM|PASTEURELLA MULTOCIDA|PASTEURELLA MULTOCIDA
C3643356|T122|1421900|RXNORM|POLYQUATERNIUM-39 (31-40-29 ACRYLIC ACID-ACRYLAMIDE-DADMAC; 1500000 MW)|POLYQUATERNIUM-39 (31-40-29 ACRYLIC ACID-ACRYLAMIDE-DADMAC; 1500000 MW)
C0071142|T195|1367292|RXNORM|PIRLIMYCIN|PIRLIMYCIN
C0771997|T121|236693|RXNORM|CALCIUM SACCHARATE|CALCIUM SACCHARATE
C0015051|T130|1314354|RXNORM|ETHOXYQUIN|ETHOXYQUIN
C2168863|T121|817555|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN / PYRILAMINE / SODIUM CITRATE|DEXTROMETHORPHAN / GUAIFENESIN / PYRILAMINE / SODIUM CITRATE
C0059747|T121|1314355|RXNORM|ETHYL ACETATE|ETHYL ACETATE
C3281333|T109|1370778|RXNORM|ORANGE PEEL EXTRACT|ORANGE PEEL EXTRACT
C3265530|T121|1370779|RXNORM|SOYBEAN GERM EXTRACT|SOYBEAN GERM EXTRACT
C0008742|T126|2530|RXNORM|CHYMOTRYPSIN|CHYMOTRYPSIN
C0008742|T126|2530|RXNORM|CHYMOTRYPSIN|CHYMOTRYPSIN
C0146011|T121|57258|RXNORM|TIZANIDINE|TIZANIDINE
C0663241|T121|190376|RXNORM|LINEZOLID|LINEZOLID
C2937575|T121|1009447|RXNORM|WASABI PREPARATION|WASABI PREPARATION
C3864851|T109|1595299|RXNORM|SACCHARIN N-(2-ACETIC ACID ETHYL ESTER)|SACCHARIN N-(2-ACETIC ACID ETHYL ESTER)
C0884979|T121|265576|RXNORM|ESCHSCHOLZIA CALIFORNICA EXTRACT|ESCHSCHOLZIA CALIFORNICA EXTRACT
C2981068|T121|1309779|RXNORM|BAPTISIA TINCTORIA ROOT EXTRACT|BAPTISIA TINCTORIA ROOT EXTRACT
C0116190|T121|49626|RXNORM|ENOXIMONE|ENOXIMONE
C1874577|T121|690608|RXNORM|BISMUTH SUBNITRATE / CALCIUM CARBONATE / MAGNESIUM CARBONATE|BISMUTH SUBNITRATE / CALCIUM CARBONATE / MAGNESIUM CARBONATE
C0446075|T004|1328760|RXNORM|PENICILLIUM GLABRUM|PENICILLIUM GLABRUM
C0077316|T121|38810|RXNORM|TRITOQUALINE|TRITOQUALINE
C0209337|T121|68139|RXNORM|ROCURONIUM|ROCURONIUM
C3484415|T121|1309677|RXNORM|DELPHINIUM STAPHISAGRIA SEED EXTRACT|DELPHINIUM STAPHISAGRIA SEED EXTRACT
C3488332|T121|1309676|RXNORM|BRYONIA ALBA ROOT EXTRACT|BRYONIA ALBA ROOT EXTRACT
C1509628|T121|1363622|RXNORM|PEG-8 DISTEARATE|PEG-8 DISTEARATE
C3256081|T121|1363623|RXNORM|PEG-8 LAURATE|PEG-8 LAURATE
C3489392|T121|1309673|RXNORM|TOXICODENDRON PUBESCENS LEAF EXTRACT|EASTERN POISON OAK LEAF EXTRACT
C3486850|T121|1309672|RXNORM|ARTEMISIA MARITIMA FLOWER EXTRACT|ARTEMISIA MARITIMA FLOWER EXTRACT
C1365471|T121|1363626|RXNORM|QUATERNIUM-52|QUATERNIUM-52
C1365469|T121|1309670|RXNORM|SARSAPARILLA ROOT EXTRACT|SARSAPARILLA ROOT EXTRACT
C0622779|T109|1363628|RXNORM|BUTYL STEARATE|BUTYL STEARATE
C3162624|T121|1370776|RXNORM|SWERTIA JAPONICA EXTRACT|SWERTIA JAPONICA EXTRACT
C3484421|T121|1309678|RXNORM|STRYCHNOS NUX-VOMICA SEED EXTRACT|STRYCHNOS NUX-VOMICA SEED EXTRACT
C1874895|T121|689891|RXNORM|CODEINE / GUAIFENESIN / PHENIRAMINE|CODEINE / GUAIFENESIN / PHENIRAMINE
C0961781|T121|299081|RXNORM|SPINOSAD|SPINOSAD
C0070325|T168|33094|RXNORM|PEPPERMINT OIL|PEPPERMINT OIL
C0048038|T121|14845|RXNORM|APRACLONIDINE|APRACLONIDINE
C0071081|T121|33724|RXNORM|PINAVERIUM|PINAVERIUM
C0070324|T121|33093|RXNORM|PEPPERMINT PREPARATION|PEPPERMINT PREPARATION
C0077072|T121|38609|RXNORM|TRICLOCARBAN|TRICLOCARBAN
C2961699|T121|1053363|RXNORM|BENZOCAINE / PETROLATUM|BENZOCAINE / PETROLATUM
C2702412|T129|995703|RXNORM|DENDRYPHIELLA VINOSA ALLERGENIC EXTRACT|DENDRYPHIELLA VINOSA ALLERGENIC EXTRACT
C3692846|T121|1442703|RXNORM|GLEDITSIA SINENSIS WHOLE EXTRACT|GLEDITSIA SINENSIS WHOLE EXTRACT
C2701669|T129|852593|RXNORM|BURNING BUSH POLLEN EXTRACT|BASSIA SCOPARIA POLLEN EXTRACT
C3486825|T121|1310141|RXNORM|EPIMEDIUM GRANDIFLORUM FLOWERING TOP EXTRACT|EPIMEDIUM GRANDIFLORUM FLOWERING TOP EXTRACT
C2955005|T121|1310140|RXNORM|GLECHOMA HEDERACEA EXTRACT|GLECHOMA HEDERACEA EXTRACT
C0631907|T109|1442707|RXNORM|HYDROXYPROPYL-ALPHA-CYCLODEXTRIN|HYDROXYPROPYL-ALPHA-CYCLODEXTRIN
C3692849|T121|1442706|RXNORM|SOPHORA FLAVESCENS WHOLE EXTRACT|SOPHORA FLAVESCENS WHOLE EXTRACT
C3692848|T121|1442705|RXNORM|SANGUISORBA OFFICINALIS WHOLE EXTRACT|SANGUISORBA OFFICINALIS WHOLE EXTRACT
C3692847|T121|1442704|RXNORM|RHEUM PALMATUM WHOLE EXTRACT|RHEUM PALMATUM WHOLE EXTRACT
C0006220|T121|1753|RXNORM|BROMHEXINE|BROMHEXINE
C3486837|T121|1310148|RXNORM|WYETHIA HELENIOIDES ROOT EXTRACT|WYETHIA HELENIOIDES ROOT EXTRACT
C2948818|T121|1044981|RXNORM|BIOTIN / NICOTINAMIDE ADENINE DINUCLEOTIDE (NAD) / PANTHENOL / ZINC PYRITHIONE|BIOTIN / NICOTINAMIDE ADENINE DINUCLEOTIDE (NAD) / PANTHENOL / ZINC PYRITHIONE
C0056059|T109|1305724|RXNORM|COCO DIETHANOLAMIDE|COCO DIETHANOLAMIDE
C0909381|T121|275891|RXNORM|VALGANCICLOVIR|VALGANCICLOVIR
C0058410|T121|23405|RXNORM|DIPIPANONE|DIPIPANONE
C3486642|T109|1355829|RXNORM|MANUKA OIL|MANUKA OIL
C0073992|T121|36117|RXNORM|SALMETEROL|SALMETEROL
C0453256|T121|125918|RXNORM|FENNEL SEED PREPARATION|FENNEL SEED PREPARATION
C2723353|T121|866645|RXNORM|TITANIUM DIOXIDE / ZINC OXIDE|TITANIUM DIOXIDE / ZINC OXIDE
C2702415|T129|892569|RXNORM|PEA ALLERGENIC EXTRACT|PEA ALLERGENIC EXTRACT
C3282045|T168|1309939|RXNORM|SORGHUM BICOLOR STEM JUICE EXTRACT|SORGHUM BICOLOR STEM JUICE
C3666147|T121|1435859|RXNORM|CYCLOPIA INTERMEDIA LEAF EXTRACT|CYCLOPIA INTERMEDIA LEAF EXTRACT
C3488910|T109|1435858|RXNORM|CETEARYL OLIVATE|CETEARYL OLIVATE
C2702370|T129|892561|RXNORM|LOBSTER ALLERGENIC EXTRACT|LOBSTER, UNSPECIFIED ALLERGENIC EXTRACT
C1999375|T121|1116632|RXNORM|TICAGRELOR|TICAGRELOR
C0207012|T109|1309206|RXNORM|MYRRH OIL|MYRRH OIL
C2928080|T121|1007158|RXNORM|CLONIXIN / CYCLOBENZAPRINE|CLONIXIN / CYCLOBENZAPRINE
C0790018|T121|1309204|RXNORM|DILL SEED OIL|DILL SEED OIL
C3848539|T196|1546398|RXNORM|SELENITE ION|SELENITE ION
C0054599|T168|1309202|RXNORM|CANOLA OIL|CANOLA OIL
C3256122|T109|1309203|RXNORM|BIXA ORELLANA SEED EXTRACT|BIXA ORELLANA SEED EXTRACT
C3255988|T109|1309200|RXNORM|ANGELICA ACUTILOBA ROOT EXTRACT|ANGELICA ACUTILOBA ROOT EXTRACT
C2365869|T109|1309201|RXNORM|BLACK PEPPER OIL|BLACK PEPPER OIL
C0700599|T121|203218|RXNORM|PYRIMETHAMINE / SULFADOXINE|PYRIMETHAMINE / SULFADOXINE
C2928072|T121|1007150|RXNORM|FLUMETHASONE / SALICYLIC ACID|FLUMETHASONE / SALICYLIC ACID
C2928075|T121|1007153|RXNORM|ASTEMIZOLE / CETRIMIDE / OXYMETAZOLINE|ASTEMIZOLE / CETRIMIDE / OXYMETAZOLINE
C2928074|T121|1007152|RXNORM|COENZYME Q10 / GINKGO BILOBA EXTRACT|COENZYME Q10 / GINKGO BILOBA EXTRACT
C2928077|T121|1007155|RXNORM|BENZOCAINE / LINDANE|BENZOCAINE / LINDANE
C2928076|T121|1007154|RXNORM|ECHINACEA PREPARATION / GOLDEN SEAL ROOT EXTRACT|ECHINACEA PREPARATION / GOLDEN SEAL ROOT EXTRACT
C2928079|T121|1007157|RXNORM|GUAIFENESIN / MENTHOL|GUAIFENESIN / MENTHOL
C2928078|T121|1007156|RXNORM|ANTIPYRINE / EPHEDRINE|ANTIPYRINE / EPHEDRINE
C0035608|T195|9384|RXNORM|RIFAMPIN|RIFAMPIN
C2344070|T129|797633|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP W-135 CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE|NEISSERIA MENINGITIDIS SEROGROUP W-135 CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE
C0035629|T121|9386|RXNORM|RIMANTADINE|RIMANTADINE
C2142867|T121|816433|RXNORM|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE
C3488990|T109|1353891|RXNORM|APRICOT EXTRACT|APRICOT EXTRACT
C1874777|T121|689279|RXNORM|CETYLPYRIDINIUM / CHLOROXYLENOL / TRIACETIN|CETYLPYRIDINIUM / CHLOROXYLENOL / TRIACETIN
C0035633|T121|9388|RXNORM|RIMITEROL|RIMITEROL
C2193958|T121|814268|RXNORM|CODEINE / EPHEDRINE / PYRILAMINE|CODEINE / EPHEDRINE / PYRILAMINE
C3495504|T121|1370787|RXNORM|OKRA EXTRACT|OKRA EXTRACT
C3484582|T121|1370786|RXNORM|VIOLA ODORATA EXTRACT|VIOLA ODORATA EXTRACT
C3474467|T109|1370785|RXNORM|GUM TALHA EXTRACT|GUM TALHA EXTRACT
C3256731|T109|1370783|RXNORM|SEAWEED EXTRACT|SEAWEED EXTRACT
C2827346|T121|1370781|RXNORM|WHEAT GLUTEN EXTRACT|WHEAT GLUTEN EXTRACT
C0910089|T109|1362577|RXNORM|1,2,6-HEXANETRIOL|1,2,6-HEXANETRIOL
C3486749|T121|1309932|RXNORM|DAPHNE ODORA BARK EXTRACT|DAPHNE ODORA BARK EXTRACT
C3535621|T121|1370789|RXNORM|MONOETHANOLAMINE LAURYL SULFATE|MONOETHANOLAMINE LAURYL SULFATE
C2928761|T121|1007847|RXNORM|ATTAPULGITE / PECTIN|ATTAPULGITE / PECTIN
C2928760|T121|1007846|RXNORM|CARBETAPENTANE / GUAIACOLSULFONIC ACID / PHENYLEPHRINE / PHENYLPROPANOLAMINE|CARBETAPENTANE / GUAIACOLSULFONIC ACID / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C2928259|T121|1007337|RXNORM|ASPIRIN / ISOSORBIDE|ASPIRIN / ISOSORBIDE
C2928258|T121|1007336|RXNORM|DEXCHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE / PYRILAMINE|DEXCHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE / PYRILAMINE
C2928757|T121|1007843|RXNORM|CHOLINE / INOSITOL|CHOLINE / INOSITOL
C2928756|T121|1007842|RXNORM|MENTHOL / PECTIN|MENTHOL / PECTIN
C2928254|T121|1007332|RXNORM|BENZYDAMINE / HEXETIDINE|BENZYDAMINE / HEXETIDINE
C3509937|T121|1370569|RXNORM|DIMERCAPTOSUCCINATE|DIMERCAPTOSUCCINATE
C2928261|T121|1007339|RXNORM|BETAMETHASONE / FUSIDATE|BETAMETHASONE / FUSIDATE
C2928260|T121|1007338|RXNORM|GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM CHLORIDE|GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM CHLORIDE
C2928763|T121|1007849|RXNORM|TRIAMCINOLONE / UREA|TRIAMCINOLONE / UREA
C2928762|T121|1007848|RXNORM|BENZOCAINE / METHYLCELLULOSE|BENZOCAINE / METHYLCELLULOSE
C3485035|T121|1304093|RXNORM|CITRIC ACID / MAGNESIUM OXIDE / PICOSULFATE SODIUM|CITRIC ACID / MAGNESIUM OXIDE / PICOSULFATE SODIUM
C2948051|T121|1043299|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / CHOLECALCIFEROL / DOCOSAHEXAENOATE / DOCUSATE / FERROUS FUMARATE / FOLIC ACID / PYRIDOXINE / TRICALCIUM PHOSPHATE|ALPHA TOCOPHEROL / ASCORBIC ACID / CHOLECALCIFEROL / DOCOSAHEXAENOATE / DOCUSATE / FERROUS FUMARATE / FOLIC ACID / PYRIDOXINE / TRICALCIUM PHOSPHATE
C1690512|T121|771220|RXNORM|CALCIUM GLUBIONATE / CALCIUM LACTOBIONATE|CALCIUM GLUBIONATE / CALCIUM LACTOBIONATE
C2718384|T129|857919|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-URUGUAY-716-2007, NYMC X-175C (H3N2) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-URUGUAY-716-2007, NYMC X-175C (H3N2) STRAIN
C0026933|T195|7145|RXNORM|MYCOPHENOLIC ACID|MYCOPHENOLIC ACID
C1120106|T195|325642|RXNORM|ERTAPENEM|ERTAPENEM
C0014838|T121|4065|RXNORM|ESCIN|ESCIN
C1120110|T121|325646|RXNORM|ALISKIREN|ALISKIREN
C0052940|T121|18747|RXNORM|BALSALAZIDE|BALSALAZIDE
C3486646|T121|1311541|RXNORM|ARONIA MELANOCARPA FRUIT EXTRACT|ARONIA MELANOCARPA FRUIT EXTRACT
C3500343|T121|1314246|RXNORM|DIMETHICONOL (100000 CST)|DIMETHICONOL (100000 CST)
C3255680|T121|1311543|RXNORM|HIBISCUS SABDARIFFA CALYX EXTRACT|HIBISCUS SABDARIFFA CALYX EXTRACT
C3500339|T129|1314240|RXNORM|INTERFERON GAMMA-1A|INTERFERON GAMMA-1A
C0068122|T121|1311545|RXNORM|N-METHYLEPHEDRINE|N-METHYLEPHEDRINE
C3255683|T109|1311546|RXNORM|HIPPOPHAE RHAMNOIDES FRUIT EXTRACT|HIPPOPHAE RHAMNOIDES FRUIT EXTRACT
C3486706|T121|1311547|RXNORM|HORDEUM VULGARE TOP EXTRACT|HORDEUM VULGARE TOP EXTRACT
C0020388|T123|1311548|RXNORM|HYDROXYPROLINE|HYDROXYPROLINE
C3488962|T168|1311549|RXNORM|ARONIA MELANOCARPA FRUIT JUICE|ARONIA MELANOCARPA FRUIT JUICE
C2726141|T129|967033|RXNORM|CANDIDA TROPICALIS ALLERGENIC EXTRACT|CANDIDA TROPICALIS ALLERGENIC EXTRACT
C3256878|T109|1314249|RXNORM|XYLITYLGLUCOSIDE|XYLITYLGLUCOSIDE
C0031013|T121|8050|RXNORM|PERHEXILINE|PERHEXILINE
C1699926|T129|1012892|RXNORM|FINGOLIMOD|FINGOLIMOD
C0939237|T121|284640|RXNORM|LOPINAVIR / RITONAVIR|LOPINAVIR / RITONAVIR
C0939238|T121|284641|RXNORM|NAPROXEN / PSEUDOEPHEDRINE|NAPROXEN / PSEUDOEPHEDRINE
C3535643|T121|1370192|RXNORM|POLYETHYLENE GLYCOL 4000000|POLYETHYLENE GLYCOL 4000000
C0359047|T121|106986|RXNORM|HYDROCORTISONE / OXYTETRACYCLINE|HYDROCORTISONE / OXYTETRACYCLINE
C0359048|T121|106987|RXNORM|CLIOQUINOL / HYDROCORTISONE|CLIOQUINOL / HYDROCORTISONE
C0359045|T121|106984|RXNORM|HYDROCORTISONE / NYSTATIN|HYDROCORTISONE / NYSTATIN
C1874834|T121|689641|RXNORM|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE
C0359177|T197|107056|RXNORM|FERROUS PHOSPHATE|FERROUS PHOSPHATE
C1874835|T121|689642|RXNORM|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PYRILAMINE|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PYRILAMINE
C0359163|T129|107051|RXNORM|HORSE ANTIHUMAN THYMOCYTE GAMMA GLOBULIN|HORSE ANTIHUMAN THYMOCYTE GAMMA GLOBULIN
C3256277|T109|1306948|RXNORM|BUTYLOCTYL SALICYLATE|BUTYLOCTYL SALICYLATE
C3484652|T121|1303322|RXNORM|CORNSTARCH / LANOLIN / ZINC OXIDE|CORNSTARCH / LANOLIN / ZINC OXIDE
C3651796|T121|1427411|RXNORM|BUTYLENE GLYCOL DICAPRYLATE|BUTYLENE GLYCOL DICAPRYLATE
C3531466|T109|1366994|RXNORM|POLYISOBUTYLENE (200000 MW)|POLYISOBUTYLENE (200000 MW)
C3255657|T109|1306940|RXNORM|CETYL PEG-PPG-10-1 DIMETHICONE (HLB 1.5)|CETYL PEG-PPG-10-1 DIMETHICONE (HLB 2)
C3255658|T109|1306941|RXNORM|CETYL PEG-PPG-10-1 DIMETHICONE (HLB 5)|CETYL PEG-PPG-10-1 DIMETHICONE (HLB 5)
C3255738|T109|1306942|RXNORM|BARLEY BRAN|BARLEY BRAN
C3255751|T109|1306943|RXNORM|CHITOSAN OLIGOSACCHARIDE|CHITOSAN OLIGOSACCHARIDE
C3255986|T109|1306944|RXNORM|AMMONIUM LAURETH-5 SULFATE|AMMONIUM LAURETH-5 SULFATE
C3256032|T121|1306945|RXNORM|DIETHYLHEXYL ADIPATE|DIETHYLHEXYL ADIPATE
C3256113|T197|1306946|RXNORM|BROWN IRON OXIDE|BROWN IRON OXIDE
C3256131|T109|1306947|RXNORM|COCAMINE OXIDE|COCAMINE OXIDE
C3190049|T121|1144134|RXNORM|BILBERRY EXTRACT / VITAMIN A / VITAMIN E|BILBERRY EXTRACT / VITAMIN A / VITAMIN E
C2701317|T129|852114|RXNORM|CULTIVATED OAT POLLEN EXTRACT|AVENA SATIVA POLLEN EXTRACT
C2243105|T121|815024|RXNORM|ESTRADIOL / PROGESTERONE|ESTRADIOL / PROGESTERONE
C3531464|T109|1366991|RXNORM|HEXADECYL POVIDONE (4 HEXADECYL BRANCHES-REPEAT)|HEXADECYL POVIDONE (4 HEXADECYL BRANCHES-REPEAT)
C3540667|T121|1421478|RXNORM|LIMULUS POLYPHEMUS EXTRACT|LIMULUS POLYPHEMUS EXTRACT
C0717976|T121|214758|RXNORM|PHENAZOPYRIDINE / SULFISOXAZOLE|PHENAZOPYRIDINE / SULFISOXAZOLE
C1656475|T121|607596|RXNORM|CARBETAPENTANE / PHENYLEPHRINE|CARBETAPENTANE / PHENYLEPHRINE
C3205023|T122|1366992|RXNORM|PEG-8 & SMDI COPOLYMER|PEG-8 & SMDI COPOLYMER
C3859729|T121|1593743|RXNORM|CHOLECALCIFEROL / FOLIC ACID|CHOLECALCIFEROL / FOLIC ACID
C0057293|T121|22427|RXNORM|DEHYDROSANOL|DEHYDROSANOL
C3859731|T123|1593745|RXNORM|COLLAGEN ALPHA-1(III) (HUMAN)|COLLAGEN ALPHA-1(III) (HUMAN)
C0246269|T121|1148138|RXNORM|ICATIBANT|ICATIBANT
C3535910|T121|1369590|RXNORM|PENTETATE CALCIUM|PENTETATE CALCIUM
C0011795|T121|3274|RXNORM|DEXTRAN 70|DEXTRAN HM
C3256737|T121|1307579|RXNORM|URTICA DIOICA ROOT EXTRACT|URTICA DIOICA ROOT EXTRACT
C2701321|T129|852118|RXNORM|JOHNSON GRASS SMUT POLLEN EXTRACT|JOHNSON GRASS SMUT POLLEN EXTRACT
C3715099|T196|1544139|RXNORM|CARBONATE ION|CARBONATE ION
C3256384|T121|1371366|RXNORM|TRIDECYL ALCOHOL|TRIDECANOL
C3537723|T121|1371367|RXNORM|GLYCYRRHIZIN, AMMONIATED PENTAHYDRATE|GLYCYRRHIZIN, AMMONIATED PENTAHYDRATE
C3537721|T121|1371364|RXNORM|CHLORHEXIDINE / KETOCONAZOLE|CHLORHEXIDINE / KETOCONAZOLE
C3537717|T121|1371360|RXNORM|KETOCONAZOLE / LACTATE / SALICYLIC ACID|KETOCONAZOLE / LACTATE / SALICYLIC ACID
C2728189|T129|1011017|RXNORM|POPPY SEED ALLERGENIC EXTRACT|POPPY SEED ALLERGENIC EXTRACT
C0947610|T121|287516|RXNORM|WATERCRESS PREPARATION|WATERCRESS PREPARATION
C0947608|T121|287515|RXNORM|SOYBEAN PREPARATION|SOYBEAN PREPARATION
C0246631|T121|73032|RXNORM|REMIFENTANIL|REMIFENTANIL
C2926844|T121|1001434|RXNORM|CAFFEINE / MAGNESIUM SALICYLATE|CAFFEINE / MAGNESIUM SALICYLATE
C0077266|T197|1364529|RXNORM|TRIPHOSPHORIC ACID|TRIPHOSPHORIC ACID
C0061938|T121|26296|RXNORM|GUANADREL|GUANADREL
C2928929|T121|1008018|RXNORM|CHOLINE / INOSITOL / NIACIN|CHOLINE / INOSITOL / NIACIN
C2709770|T129|854966|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 6B VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 6B VACCINE
C2709764|T129|854960|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 33F VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 33F VACCINE
C0042845|T127|11248|RXNORM|VITAMIN B 12|VITAMIN B 12
C2709766|T129|854962|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 4 VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 4 VACCINE
C2928922|T121|1008011|RXNORM|ERGOCALCIFEROL / ZINC OXIDE|ERGOCALCIFEROL / ZINC OXIDE
C2928921|T121|1008010|RXNORM|POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC|POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC
C2928924|T121|1008013|RXNORM|MAGNESIUM MALATE / MALIC ACID / VITAMIN B6|MAGNESIUM MALATE / MALIC ACID / VITAMIN B6
C0042839|T127|11246|RXNORM|VITAMIN A|VITAMIN A
C0042839|T127|11246|RXNORM|VITAMIN A|VITAMIN A
C2928926|T121|1008015|RXNORM|ASCORBIC ACID / BETA CAROTENE / CALCIUM CARBONATE, PRECIPITATED / CHOLECALCIFEROL / FOLIC ACID / IRON CARBONYL / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / BETA CAROTENE / CALCIUM CARBONATE, PRECIPITATED / CHOLECALCIFEROL / FOLIC ACID / IRON CARBONYL / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN E / ZINC OXIDE
C2928925|T121|1008014|RXNORM|GARLIC PREPARATION / GUGULU EXTRACT / NIACIN|GARLIC PREPARATION / GUGULU EXTRACT / NIACIN
C2928928|T121|1008017|RXNORM|NIACIN / ZINC CITRATE|NIACIN / ZINC CITRATE
C2928927|T121|1008016|RXNORM|DIMETHICONE / MINERAL OIL|DIMETHICONE / MINERAL OIL
C0123931|T121|51499|RXNORM|IRINOTECAN|IRINOTECAN
C0002575|T121|689|RXNORM|AMINOPHYLLINE|AMINOPHYLLINE
C0070093|T125|32915|RXNORM|TERIPARATIDE|TERIPARATIDE
C0795597|T121|968804|RXNORM|CYTARABINE LIPOSOME|CYTARABINE LIPOSOME
C0030077|T121|7815|RXNORM|OXYPERTINE|OXYPERTINE
C0981834|T129|852496|RXNORM|ARIZONA ASH POLLEN EXTRACT|FRAXINUS VELUTINA POLLEN EXTRACT
C0134110|T121|1482634|RXNORM|ORNITHINE ALPHA-KETOGLUTARATE|ORNITHINE OXOGLUTARATE
C0771276|T121|1482633|RXNORM|ARGININE PYROGLUTAMATE|ARGININE PYROGLUTAMATE
C0051235|T121|17376|RXNORM|ALLYL SULFIDE|ALLYL SULFIDE
C0126789|T121|52364|RXNORM|MAGNESIUM SALICYLATE|MAGNESIUM SALICYLATE
C1329985|T121|404780|RXNORM|BROMPHENIRAMINE / HYDROCODONE / PSEUDOEPHEDRINE|BROMPHENIRAMINE / HYDROCODONE / PSEUDOEPHEDRINE
C3488432|T121|1426439|RXNORM|EUROPEAN FLOUNDER PREPARATION|EUROPEAN FLOUNDER PREPARATION
C3488431|T121|1426438|RXNORM|EDIBLE OYSTER PREPARATION|EDIBLE OYSTER PREPARATION
C1329990|T121|404785|RXNORM|CARBETAPENTANE / PHENYLEPHRINE / PYRILAMINE|CARBETAPENTANE / PHENYLEPHRINE / PYRILAMINE
C3256708|T109|1309449|RXNORM|OENOTHERA BIENNIS FLOWER EXTRACT|OENOTHERA BIENNIS FLOWER EXTRACT
C1329991|T121|404786|RXNORM|CARBIDOPA / ENTACAPONE / LEVODOPA|CARBIDOPA / ENTACAPONE / LEVODOPA
C1329994|T121|404789|RXNORM|CHLORPHENIRAMINE / IBUPROFEN / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / IBUPROFEN / PSEUDOEPHEDRINE
C3256700|T109|1309445|RXNORM|MYRTUS COMMUNIS LEAF EXTRACT|MYRTUS COMMUNIS LEAF EXTRACT
C3256784|T109|1309446|RXNORM|NARCISSUS PSEUDONARCISSUS FLOWER EXTRACT|NARCISSUS PSEUDONARCISSUS FLOWER EXTRACT
C3255703|T109|1309447|RXNORM|NELUMBO NUCIFERA FLOWER EXTRACT|NELUMBO NUCIFERA FLOWER EXTRACT
C3255947|T109|1309440|RXNORM|MAGNOLIA OBOVATA BARK EXTRACT|MAGNOLIA OBOVATA BARK EXTRACT
C3256419|T121|1309441|RXNORM|MAHONIA AQUIFOLIUM ROOT EXTRACT|BERBERIS AQUIFOLIUM ROOT EXTRACT
C3256366|T109|1309442|RXNORM|MORINGA OLEIFERA SEED EXTRACT|MORINGA OLEIFERA SEED EXTRACT
C3256367|T109|1309443|RXNORM|MORINGA OLEIFERA SEED OIL|MORINGA OLEIFERA SEED OIL
C3555489|T121|1376341|RXNORM|3-(3,4-METHYLENEDIOXYPHENYL)-2-METHYLPROPANAL|3-(3,4-METHYLENEDIOXYPHENYL)-2-METHYLPROPANAL
C2741277|T129|900743|RXNORM|WESTERN WHITE PINE POLLEN EXTRACT|PINUS MONTICOLA POLLEN EXTRACT
C0717481|T121|214287|RXNORM|BENAZEPRIL / HYDROCHLOROTHIAZIDE|BENAZEPRIL / HYDROCHLOROTHIAZIDE
C3857965|T109|1551309|RXNORM|ORCHIS MASCULA FLOWER EXTRACT|ORCHIS MASCULA FLOWER EXTRACT
C3256184|T121|1307314|RXNORM|ROBUSTA COFFEE BEAN EXTRACT|ROBUSTA COFFEE BEAN EXTRACT
C0030776|T122|1307312|RXNORM|POLYETHYLENE GLYCOL 8000|POLYETHYLENE GLYCOL 8000
C2827307|T121|1307313|RXNORM|POLYETHYLENE GLYCOL 800|POLYETHYLENE GLYCOL 800
C2827099|T121|1307310|RXNORM|CAPRYLIC(CAPRIC MONO)DIGLCYERIDES|CAPRYLIC(CAPRIC MONO)DIGLCYERIDES
C0717482|T121|214288|RXNORM|BENDROFLUMETHIAZIDE / NADOLOL|BENDROFLUMETHIAZIDE / NADOLOL
C2194179|T121|813631|RXNORM|ALLOPURINOL / BENZBROMARONE|ALLOPURINOL / BENZBROMARONE
C3535922|T121|1370012|RXNORM|CHOLECALCIFEROL / MAGNESIUM OXIDE / TURMERIC EXTRACT|CHOLECALCIFEROL / MAGNESIUM OXIDE / TURMERIC EXTRACT
C0074281|T197|36345|RXNORM|SELENIUM SULFIDE|SELENIUM SULFIDE
C0074280|T197|36344|RXNORM|SELENIOUS ACID|SELENIOUS ACID
C0767550|T121|1368877|RXNORM|ILOMASTAT|ILOMASTAT
C3700984|T121|1487006|RXNORM|OCLACITINIB|OCLACITINIB
C0085259|T195|42372|RXNORM|MUPIROCIN|MUPIROCIN
C0085259|T195|42372|RXNORM|MUPIROCIN|MUPIROCIN
C0085272|T125|42375|RXNORM|LEUPROLIDE|LEUPROLIDE
C0050403|T121|16689|RXNORM|ACECLOFENAC|ACECLOFENAC
C2730230|T129|892620|RXNORM|EGG YOLK (CHICKEN) ALLERGENIC EXTRACT|EGG YOLK (CHICKEN) ALLERGENIC EXTRACT
C2016119|T121|820527|RXNORM|ACETAMINOPHEN / OXATOMIDE / PHENYLEPHRINE|ACETAMINOPHEN / OXATOMIDE / PHENYLEPHRINE
C0050393|T121|16681|RXNORM|ACARBOSE|ACARBOSE
C0079441|T123|1370419|RXNORM|TRANSFORMING GROWTH FACTOR BETA 2|TRANSFORMING GROWTH FACTOR BETA 2
C0077027|T121|1370418|RXNORM|TRICAINE|TRICAINE
C3180892|T121|1373206|RXNORM|4-TERT-BUTYLCYCLOHEXANOL|4-TERT-BUTYLCYCLOHEXANOL
C3538629|T121|1373205|RXNORM|APIS CERANA WORKER SECRETION PREPARATION|APIS CERANA WORKER SECRETION PREPARATION
C0982358|T121|1373204|RXNORM|PPG-20 METHYL GLUCOSE ETHER DISTEARATE|PPG-20 METHYL GLUCOSE ETHER DISTEARATE
C0017814|T130|4888|RXNORM|GLUTARAL|GLUTARAL
C0039468|T121|10355|RXNORM|TEMAZEPAM|TEMAZEPAM
C2929802|T121|1008905|RXNORM|CHROMIC CHLORIDE / COPPER SULFATE / MANGANESE SULFATE / ZINC SULFATE|CHROMIC CHLORIDE / COPPER SULFATE / MANGANESE SULFATE / ZINC SULFATE
C2929801|T121|1008904|RXNORM|ALANINE / GLUTAMATE / GLYCINE / THIAMINE|ALANINE / GLUTAMATE / GLYCINE / THIAMINE
C0009316|T195|2709|RXNORM|COLISTIN|COLISTIN
C0009315|T195|2708|RXNORM|COLISTIMETHATE|COLISTIMETHATE
C2929798|T121|1008901|RXNORM|CHLORPHENIRAMINE / PSEUDOEPHEDRINE / SCOPOLAMINE|CHLORPHENIRAMINE / PSEUDOEPHEDRINE / SCOPOLAMINE
C2929797|T121|1008900|RXNORM|BETAMETHASONE / SULFACETAMIDE|BETAMETHASONE / SULFACETAMIDE
C0012145|T125|3368|RXNORM|DIENESTROL|DIENESTROL
C0220578|T121|70561|RXNORM|PALONOSETRON|PALONOSETRON
C0017797|T123|4885|RXNORM|GLUTAMINE|GLUTAMINE
C2929806|T121|1008909|RXNORM|CHLORZOXAZONE / CLONIXIN|CHLORZOXAZONE / CLONIXIN
C2929805|T121|1008908|RXNORM|ALTHIAZIDE / SPIRONOLACTONE|ALTHIAZIDE / SPIRONOLACTONE
C0030771|T195|7960|RXNORM|PEFLOXACIN|PEFLOXACIN
C0040610|T121|10689|RXNORM|TRAMADOL|TRAMADOL
C0030800|T121|7966|RXNORM|PEMOLINE|PEMOLINE
C0982328|T197|314774|RXNORM|PENTETATE PENTASODIUM|PENTETATE PENTASODIUM
C0982330|T121|314776|RXNORM|PEPTONE,DRIED|PEPTONE,DRIED
C2929947|T121|1009052|RXNORM|MAGNESIUM CITRATE / POTASSIUM CITRATE|MAGNESIUM CITRATE / POTASSIUM CITRATE
C2929948|T121|1009053|RXNORM|ACETAMINOPHEN / BENZYDAMINE / TETRACYCLINE|ACETAMINOPHEN / BENZYDAMINE / TETRACYCLINE
C2929945|T121|1009050|RXNORM|CALCIUM CARBONATE / PYROGLUTAMATE|CALCIUM CARBONATE / PYROGLUTAMATE
C2929946|T121|1009051|RXNORM|CAMPHOR / METHYLNICOTINATE|CAMPHOR / METHYLNICOTINATE
C2927872|T121|1006949|RXNORM|ACTIVATED CHARCOAL / BILE SALTS / PANCREATIN|ACTIVATED CHARCOAL / BILE SALTS / PANCREATIN
C2927871|T121|1006948|RXNORM|ASCORBIC ACID / NIACINAMIDE / VITAMIN A|ASCORBIC ACID / NIACINAMIDE / VITAMIN A
C2929949|T121|1009054|RXNORM|AJMALINE / ALMITRINE|AJMALINE / ALMITRINE
C2929950|T121|1009055|RXNORM|SAW PALMETTO FRUIT EXTRACT / ZINC PICOLINATE|SAW PALMETTO FRUIT EXTRACT / ZINC PICOLINATE
C2927868|T121|1006945|RXNORM|CALCIUM PHOSPHATE / PROCYANIDOLIC OLIGOMER|CALCIUM PHOSPHATE / PROCYANIDOLIC OLIGOMER
C2927867|T121|1006944|RXNORM|CHLORAMPHENICOL / NAPHAZOLINE / NEOMYCIN|CHLORAMPHENICOL / NAPHAZOLINE / NEOMYCIN
C2927870|T121|1006947|RXNORM|ASCORBIC ACID / ECHINACEA PREPARATION / GOLDEN SEAL ROOT|ASCORBIC ACID / ECHINACEA PREPARATION / GOLDEN SEAL ROOT
C2929954|T121|1009059|RXNORM|FRANGULA PREPARATION / KARAYA GUM|FRANGULA PREPARATION / KARAYA GUM
C2927864|T121|1006941|RXNORM|GLYCOLATE / LACTATE|GLYCOLATE / LACTATE
C2927863|T121|1006940|RXNORM|SIBERIAN GINSENG ROOT / ST. JOHN'S WORT EXTRACT|SIBERIAN GINSENG ROOT / ST. JOHN'S WORT EXTRACT
C2927866|T121|1006943|RXNORM|CHROMIC SULFATE / ZINC SULFATE|CHROMIC SULFATE / ZINC SULFATE
C2927865|T121|1006942|RXNORM|GLUTAMINE / TYROSINE|GLUTAMINE / TYROSINE
C3818747|T109|1494846|RXNORM|MOSCHUS BEREZOVSKII MUSK SAC RESIN|MOSCHUS BEREZOVSKII MUSK SAC RESIN
C3818748|T109|1494845|RXNORM|METHACRYLIC ACID - ETHYL ACRYLATE COPOLYMER (4500 MPA.S)|METHACRYLIC ACID - ETHYL ACRYLATE COPOLYMER (4500 MPA.S)
C3668750|T121|1441375|RXNORM|CHLOPHEDIANOL / DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE|CHLOPHEDIANOL / DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE
C3244837|T121|1189803|RXNORM|SIMVASTATIN / SITAGLIPTIN|SIMVASTATIN / SITAGLIPTIN
C0763533|T121|232540|RXNORM|RED YEAST RICE|RED YEAST RICE
C3255672|T121|1310088|RXNORM|ERIOBOTRYA JAPONICA LEAF EXTRACT|ERIOBOTRYA JAPONICA LEAF EXTRACT
C3485574|T121|1310087|RXNORM|POLYGALA SENEGA ROOT EXTRACT|POLYGALA SENEGA ROOT EXTRACT
C3486756|T121|1310084|RXNORM|PINUS SYLVESTRIS FLOWERING TOP EXTRACT|PINUS SYLVESTRIS FLOWERING TOP EXTRACT
C3255666|T121|1310085|RXNORM|ENTADA PHASEOLOIDES LEAF EXTRACT|ENTADA PHASEOLOIDES LEAF EXTRACT
C3255617|T121|1310082|RXNORM|TRICHOSANTHES KIRILOWII ROOT EXTRACT|TRICHOSANTHES KIRILOWII ROOT EXTRACT
C3255665|T121|1310083|RXNORM|ELEUTHEROCOCCUS NODIFLORUS ROOT BARK EXTRACT|ELEUTHEROCOCCUS NODIFLORUS ROOT BARK EXTRACT
C3485015|T121|1310080|RXNORM|PLANTAGO MAJOR SEED EXTRACT|PLANTAGO MAJOR SEED EXTRACT
C3486755|T121|1310081|RXNORM|PILOCARPUS JABORANDI LEAF EXTRACT|PILOCARPUS JABORANDI LEAF EXTRACT
C0537439|T129|139896|RXNORM|ENFUVIRTIDE|ENFUVIRTIDE
C0030909|T126|8016|RXNORM|PEPSIN A|PEPSIN A
C2929402|T121|1008498|RXNORM|DANTHRON / DOCUSATE / PANTOTHENATE|DANTHRON / DOCUSATE / PANTOTHENATE
C0012471|T125|3477|RXNORM|DINOPROST|DINOPROST
C2725884|T129|895527|RXNORM|EUROPEAN RABBIT HAIR EXTRACT|ORYCTOLAGUS CUNICULUS HAIR EXTRACT
C3255039|T121|1235990|RXNORM|GLYCINE / LICORICE|GLYCINE / LICORICE
C0033743|T121|8886|RXNORM|PROTRIPTYLINE|PROTRIPTYLINE
C0012472|T125|3478|RXNORM|DINOPROSTONE|DINOPROSTONE
C2929399|T121|1008495|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP A OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP C OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP W-135 OLIGOSACCHARIDE DIPHTH|NEISSERIA MENINGITIDIS SEROGROUP A OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP C OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP W-135 OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / NEISSERIA MENINGITIDIS SEROGROUP Y OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C3255744|T121|1311376|RXNORM|CHAMAEMELUM NOBILE EXTRACT|CHAMAEMELUM NOBILE EXTRACT
C0055134|T197|20599|RXNORM|CESIUM CHLORIDE|CESIUM CHLORIDE
C2756160|T129|967529|RXNORM|RHODOTORULA MUCILAGINOSA EXTRACT|RHODOTORULA MUCILAGINOSA EXTRACT
C0022611|T121|1311375|RXNORM|KEROSENE|KEROSENE
C3194750|T121|1117114|RXNORM|BIOTIN / NIACINAMIDE / PANTHENOL / ZINC PYRITHIONE|BIOTIN / NIACINAMIDE / PANTHENOL / ZINC PYRITHIONE
C4082272|T195|26397|RXNORM|HABEKACIN|ARBEKACIN
C0079083|T121|40048|RXNORM|CARBOPLATIN|CARBOPLATIN
C2025214|T121|818929|RXNORM|CARISOPRODOL / NAPROXEN|CARISOPRODOL / NAPROXEN
C0040815|T123|1311373|RXNORM|TREHALOSE|TREHALOSE
C2606556|T121|1442132|RXNORM|MACITENTAN|MACITENTAN
C0178485|T123|1368625|RXNORM|ARACHIDONATE|ARACHIDONATE
C2929559|T121|1008659|RXNORM|HYDROCHLOROTHIAZIDE / MEPINDOLOL|HYDROCHLOROTHIAZIDE / MEPINDOLOL
C2929558|T121|1008658|RXNORM|DIETHYLAMINE SALICYLATE / METHYL SALICYLATE / NIACIN|DIETHYLAMINE SALICYLATE / METHYL SALICYLATE / NIACIN
C2929557|T121|1008657|RXNORM|INDOMETHACIN / LAURETH-9|INDOMETHACIN / POLIDOCANOL
C2929556|T121|1008656|RXNORM|ANTHRALIN / UREA|ANTHRALIN / UREA
C2929555|T121|1008655|RXNORM|NIACIN / PROCAINE / SALICYLAMIDE|NIACIN / PROCAINE / SALICYLAMIDE
C2929554|T121|1008654|RXNORM|FLUPREDNIDENE / SALICYLIC ACID|FLUPREDNIDENE / SALICYLIC ACID
C2929553|T121|1008653|RXNORM|ETHYL HEXYL SALICYLATE / TITANIUM DIOXIDE|ETHYL HEXYL SALICYLATE / TITANIUM DIOXIDE
C2929552|T121|1008652|RXNORM|CLOTRIMAZOLE / ZINC OXIDE|CLOTRIMAZOLE / ZINC OXIDE
C2929551|T121|1008651|RXNORM|BETAMETHASONE / DICLOFENAC / VITAMIN B 12|BETAMETHASONE / DICLOFENAC / VITAMIN B 12
C2929550|T121|1008650|RXNORM|AMINACRINE / LIDOCAINE|AMINACRINE / LIDOCAINE
C3666235|T121|1435991|RXNORM|C18-C21 ALKANE|C18-C21 ALKANE
C0006819|T007|1435992|RXNORM|CAMPYLOBACTER JEJUNI|CAMPYLOBACTER JEJUNI
C1874068|T121|690018|RXNORM|ALLANTOIN / CAMPHOR / PHENOL|ALLANTOIN / CAMPHOR / PHENOL
C3535911|T121|1368950|RXNORM|EDETATE CALCIUM|EDETATE CALCIUM
C1874066|T121|690016|RXNORM|ALLANTOIN / AMINACRINE / SULFISOXAZOLE|ALLANTOIN / AMINACRINE / SULFISOXAZOLE
C1874065|T121|690015|RXNORM|ALLANTOIN / AMINACRINE / SULFANILAMIDE|ALLANTOIN / AMINACRINE / SULFANILAMIDE
C3538176|T121|1372310|RXNORM|GLYCERYL 1-DIACETYLTARTARATE 2,3-STEARATE|GLYCERYL 1-DIACETYLTARTARATE 2,3-STEARATE
C2722018|T129|974650|RXNORM|BLACK OLIVE ALLERGENIC EXTRACT|OLEA EUROPAEA ALLERGENIC EXTRACT
C3818818|T109|1489549|RXNORM|PEG-40 SORBITAN STEARATE|PEG-40 SORBITAN STEARATE
C3834100|T109|1541709|RXNORM|MALLOTUS JAPONICUS FLOWER OIL|MALLOTUS JAPONICUS FLOWER OIL
C3834101|T109|1541708|RXNORM|ARCTIUM LAPPA FRUIT OIL|ARCTIUM LAPPA FRUIT OIL
C0981957|T130|851914|RXNORM|RED ALDER POLLEN EXTRACT|ALNUS RUBRA POLLEN EXTRACT
C2701152|T129|851910|RXNORM|WHITE ALDER POLLEN EXTRACT|ALNUS RHOMBIFOLIA POLLEN EXTRACT
C2929855|T121|1008959|RXNORM|THIOCTATE / VITAMIN B 12|THIOCTATE / VITAMIN B 12
C0879399|T129|263010|RXNORM|TOSITUMOMAB|TOSITUMOMAB
C0026402|T196|7024|RXNORM|MOLYBDENUM|MOLYBDENUM
C2684345|T129|851918|RXNORM|MEADOW FESCUE GRASS POLLEN EXTRACT|FESTUCA PRATENSIS POLLEN EXTRACT
C3695947|T121|1484855|RXNORM|CANNABIS SATIVA SUBSP. FLOWERING TOP EXTRACT|CANNABIS SATIVA SUBSP. FLOWERING TOP EXTRACT
C3695948|T121|1484854|RXNORM|CANNAVIS SATIVA SUSP. INDICA TOP EXTRACT|CANNAVIS SATIVA SUSP. INDICA TOP EXTRACT
C0010590|T195|3007|RXNORM|CYCLOSERINE|CYCLOSERINE
C3488088|T121|1311288|RXNORM|MEPHITIS MEPHITIS ANAL GLAND FLUID PREPARATION|MEPHITIS MEPHITIS ANAL GLAND FLUID PREPARATION
C0010582|T121|3001|RXNORM|CYCLOPENTOLATE|CYCLOPENTOLATE
C0010581|T121|3000|RXNORM|CYCLOPENTHIAZIDE|CYCLOPENTHIAZIDE
C3695949|T109|1484853|RXNORM|HUMAN DANDER PREPARATION|HUMAN DANDER PREPARATION
C0010583|T121|3002|RXNORM|CYCLOPHOSPHAMIDE|CYCLOPHOSPHAMIDE
C0392418|T197|1311283|RXNORM|MERCUROUS IODIDE PREPARATION|MERCUROUS IODIDE PREPARATION
C0038411|T007|1311281|RXNORM|STREPTOCOCCUS PYOGENES|STREPTOCOCCUS PYOGENES
C0032207|T196|1311280|RXNORM|PLATINUM|PLATINUM
C0006668|T125|1311287|RXNORM|CALCITONIN|CALCITONIN
C0010592|T121|3008|RXNORM|CYCLOSPORINE|CYCLOSPORINE
C0010592|T121|3008|RXNORM|CYCLOSPORINE|CYCLOSPORINE
C3497929|T121|1311285|RXNORM|ERSOFERMIN|ERSOFERMIN
C2347235|T121|1307954|RXNORM|SANGUISORBA OFFICINALIS ROOT EXTRACT|GREAT BURNET ROOT EXTRACT
C3255786|T121|1307955|RXNORM|OLEA EUROPAEA LEAF EXTRACT|OLEA EUROPAEA LEAF EXTRACT
C0005575|T127|1588|RXNORM|BIOTIN|BIOTIN
C0005578|T121|1589|RXNORM|BIPERIDEN|BIPERIDEN
C3255847|T109|1307951|RXNORM|LEVANT COTTONSEED OIL|LEVANT COTTONSEED OIL
C2347335|T121|1307952|RXNORM|AZADIRACHTA INDICA FLOWER EXTRACT|NEEM EXTRACT
C3488983|T121|1307953|RXNORM|LESSER GALANGAL ROOT EXTRACT|LESSER GALANGAL ROOT EXTRACT
C2726146|T129|1192729|RXNORM|COLLETOTRICHUM COCCODES ALLERGENIC EXTRACT|COLLETOTRICHUM COCCODES ALLERGENIC EXTRACT
C3695929|T109|1485183|RXNORM|PEG-30 CASTOR OIL|PEG-30 CASTOR OIL
C3695928|T122|1485184|RXNORM|C12-15 PARETH-3|C12-15 PARETH-3
C3651787|T121|1428219|RXNORM|EUONYMUS ATROPURPUREUS BRANCH BARK-ROOT BARK EXTRACT|EUONYMUS ATROPURPUREUS BRANCH BARK-ROOT BARK EXTRACT
C2726811|T109|1363620|RXNORM|PEG-75 STEARATE|PEG-75 STEARATE
C3528797|T121|1363381|RXNORM|ALUMINUM MAGNESIUM SILICATE / CALCIUM CARBONATE / SODIUM BICARBONATE|ALUMINUM MAGNESIUM SILICATE / CALCIUM CARBONATE / SODIUM BICARBONATE
C3474075|T121|1358954|RXNORM|LILIUM LANCIFOLIUM WHOLE EXTRACT|LILIUM LANCIFOLIUM WHOLE EXTRACT
C1998239|T121|758660|RXNORM|LAMIVUDINE / NEVIRAPINE / STAVUDINE|LAMIVUDINE / NEVIRAPINE / STAVUDINE
C1719900|T121|644637|RXNORM|ALLANTOIN / LIDOCAINE|ALLANTOIN / LIDOCAINE
C0452457|T168|1358955|RXNORM|LEMON JUICE|LEMON JUICE
C3497908|T121|1313239|RXNORM|ISOCETYL MYRISTATE|ISOCETYL MYRISTATE
C0034504|T123|9100|RXNORM|RACEMETHIONINE|RACEMETHIONINE
C0020823|T121|5657|RXNORM|IFOSFAMIDE|IFOSFAMIDE
C3651727|T121|1430129|RXNORM|NICOTIANA TABACUM WHOLE EXTRACT|NICOTIANA TABACUM WHOLE EXTRACT
C0020811|T121|5653|RXNORM|IDOXURIDINE|IDOXURIDINE
C0020789|T121|5650|RXNORM|IDARUBICIN|IDARUBICIN
C0286079|T121|83171|RXNORM|CIDOFOVIR|CIDOFOVIR
C0719838|T121||RXNORM|GLUCOSE / POTASSIUM CHLORIDE
C0244994|T168|72385|RXNORM|WHEAT GERM OIL|WHEAT GERM OIL
C3153839|T121|1100261|RXNORM|ASCORBIC ACID / CALCIUM CITRATE / CHOLECALCIFEROL / FOLIC ACID / IRON CARBONYL / PYRIDOXINE|ASCORBIC ACID / CALCIUM CITRATE / CHOLECALCIFEROL / FOLIC ACID / IRON CARBONYL / PYRIDOXINE
C3486388|T121|1350209|RXNORM|FRANGULA PURSHIANA BARK EXTRACT|FRANGULA PURSHIANA BARK EXTRACT
C0677829|T121|196319|RXNORM|PALIFERMIN|PALIFERMIN
C3643367|T109|1421436|RXNORM|ZINGIBER MOUTANUM FLOWERING TOP EXTRACT|ZINGIBER MOUTANUM FLOWERING TOP EXTRACT
C2194181|T121|815923|RXNORM|ALLOPURINOL / PROBENECID|ALLOPURINOL / PROBENECID
C0877804|T121|262272|RXNORM|CLOTRIMAZOLE / HYDROCORTISONE|CLOTRIMAZOLE / HYDROCORTISONE
C3643366|T109|1421437|RXNORM|PPG-2 HYDROXYETHYL COCAMIDE|PPG-2 HYDROXYETHYL COCAMIDE
C3488587|T121|1358958|RXNORM|CITRULLUS COLOCYNTHIS FRUIT EXTRACT|CITRULLUS COLOCYNTHIS FRUIT EXTRACT
C3486687|T121|1351001|RXNORM|HELLEBORUS EXTRACT|STINKING HELLEBORE ROOT EXTRACT
C3486594|T121|1351000|RXNORM|AETHUSA CYNAPIUM EXTRACT|POISON PARSLEY EXTRACT
C3488433|T121|1351003|RXNORM|GALIUM ODORATUM EXTRACT|GALIUM ODORATUM EXTRACT
C3486751|T121|1351002|RXNORM|LEONURUS CARDIACA EXTRACT|LEONURUS CARDIACA EXTRACT
C3643368|T109|1421435|RXNORM|CRINUM ASIATICUM WHOLE EXTRACT|CRINUM ASIATICUM WHOLE EXTRACT
C3643371|T109|1421432|RXNORM|BARLERIA PRIONITIS WHOLE EXTRACT|BARLERIA PRIONITIS WHOLE EXTRACT
C2364526|T129|805524|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED, B-FLORIDA-4-2006-LIKE VIRUS (B-FLORIDA-4-2006) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED, B-FLORIDA-4-2006-LIKE VIRUS (B-FLORIDA-4-2006) STRAIN
C3700897|T121|1486503|RXNORM|WHITE MUSTARD SEED EXTRACT|WHITE MUSTARD SEED EXTRACT
C3643370|T109|1421433|RXNORM|CAJANIUS CAJAN LEAF EXTRACT|CAJANIUS CAJAN LEAF EXTRACT
C2928380|T121|1007458|RXNORM|OXYQUINOLINE / SODIUM TARTRATE|OXYQUINOLINE / SODIUM TARTRATE
C2928381|T121|1007459|RXNORM|ARGININE / MALATE|ARGININE / MALATE
C0016294|T125|4458|RXNORM|FLUMETHASONE|FLUMETASONE
C2928372|T121|1007450|RXNORM|AMINOPHYLLINE / PAPAVERINE / PHENOBARBITAL|AMINOPHYLLINE / PAPAVERINE / PHENOBARBITAL
C2928373|T121|1007451|RXNORM|MAGNESIUM OXIDE / ZINC OXIDE|MAGNESIUM OXIDE / ZINC OXIDE
C2928374|T121|1007452|RXNORM|MECHLORETHAMINE / QUININE / TERPIN HYDRATE|MECHLORETHAMINE / QUININE / TERPIN HYDRATE
C2928375|T121|1007453|RXNORM|ALGINIC ACID / CALCIUM CARBONATE|ALGINIC ACID / CALCIUM CARBONATE
C2928376|T121|1007454|RXNORM|COAL TAR / FLUOCINOLONE|COAL TAR / FLUOCINOLONE
C2928377|T121|1007455|RXNORM|ASCORBIC ACID / ZINC ACETATE|ASCORBIC ACID / ZINC ACETATE
C2928378|T121|1007456|RXNORM|ANETHOLE / CHOLINE|ANETHOLE / CHOLINE
C2928379|T121|1007457|RXNORM|PANTOTHENIC ACID / SIMETHICONE|PANTOTHENIC ACID / SIMETHICONE
C0754188|T121|228656|RXNORM|AMPRENAVIR|AMPRENAVIR
C1509852|T121|479542|RXNORM|ASTRAGALUS ROOT EXTRACT|ASTRAGALUS ROOT EXTRACT
C0029983|T195|7773|RXNORM|OXACILLIN|OXACILLIN
C2741351|T129|901011|RXNORM|POST OAK POLLEN EXTRACT|QUERCUS STELLATA POLLEN EXTRACT
C0043513|T121|1535252|RXNORM|ZOLAZEPAM|ZOLAZEPAM
C0029995|T125|7779|RXNORM|OXANDROLONE|OXANDROLONE
C0029994|T121|7778|RXNORM|OXAMNIQUINE|OXAMNIQUINE
C0041030|T121|10824|RXNORM|METIPRANOLOL|METIPRANOLOL
C0053799|T121|19484|RXNORM|BISOPROLOL|BISOPROLOL
C0605193|T121|158507|RXNORM|FENBUTRAZATE|FENBUTRAZATE
C1719818|T121|758886|RXNORM|SALICYLIC ACID / ZINC OXIDE|SALICYLIC ACID / ZINC OXIDE
C0072238|T121|34706|RXNORM|PROPYLPARABEN|PROPYLPARABEN
C0031866|T123|8310|RXNORM|PHYTOSTEROLS|PHYTOSTEROLS
C0676831|T129|196102|RXNORM|BASILIXIMAB|BASILIXIMAB
C0288495|T121|83885|RXNORM|PROXIBARBAL|PROXIBARBAL
C0262964|T195|78903|RXNORM|CAPREOMYCIN|CAPREOMYCIN
C0262960|T195|78902|RXNORM|SULFACYTINE|SULFACYTINE
C0939867|T121|259314|RXNORM|BLACK PEPPER PREPARATION|BLACK PEPPER PREPARATION
C0262965|T121|78904|RXNORM|CHLORMADINONE|CHLORMADINONE
C1875227|T121|689455|RXNORM|GUAIFENESIN / HYDROCODONE / PHENINDAMINE|GUAIFENESIN / HYDROCODONE / PHENINDAMINE
C0771199|T121|235987|RXNORM|COBALT GLUCONATE|COBALT GLUCONATE
C1875226|T121|689453|RXNORM|GUAIACOL / METHYL SALICYLATE|GUAIACOL / METHYL SALICYLATE
C1875229|T121|689458|RXNORM|GUAIFENESIN / HYDROCODONE / PHENYLPROPANOLAMINE / SALICYLAMIDE|GUAIFENESIN / HYDROCODONE / PHENYLPROPANOLAMINE / SALICYLAMIDE
C0724549|T121|221072|RXNORM|CERIVASTATIN SODIUM|CERIVASTATIN SODIUM
C0072916|T121|35255|RXNORM|CISAPRIDE|CISAPRIDE
C0001981|T121|460|RXNORM|ALCURONIUM|ALCURONIUM
C3256229|T109|1426607|RXNORM|DIPENTAERYTHRITYL HEXACAPRYLATE|DIPENTAERYTHRITYL HEXACAPRYLATE
C0010558|T130|1426609|RXNORM|CYCLODEXTRINS|CYCLODEXTRINS
C0314976|T007|100213|RXNORM|BIFIDOBACTERIUM INFANTIS|BIFIDOBACTERIUM INFANTIS
C3486647|T129|1313283|RXNORM|ASPERGILLUS NIGER IMMUNOSERUM RABBIT|ASPERGILLUS NIGER IMMUNOSERUM RABBIT
C0939879|T121|1307767|RXNORM|LAVENDER EXTRACT|LAVANDULA ANGUSTIFOLIA SUBSP. ANGUSTIFOLIA FLOWERING TOP EXTRACT
C3256759|T121|1307766|RXNORM|CAPRYLYL GLUCOSIDE|CAPRYLYL GLUCOSIDE
C0068322|T109|1307764|RXNORM|1-VINYL-2-PYRROLIDONE|1-VINYL-2-PYRROLIDONE
C3255675|T121|1307763|RXNORM|HELIANTHUS ANNUUS SEEDCAKE EXTRACT|HELIANTHUS ANNUUS SEEDCAKE EXTRACT
C3256409|T121|1307762|RXNORM|ANHYDROXYLITOL|ANHYDROXYLITOL
C3256480|T109|1307761|RXNORM|1-DECENE|1-DECENE
C3256808|T121|1307760|RXNORM|SIMMONDSIA CHINENSIS SEED WAX EXTRACT|SIMMONDSIA CHINENSIS SEED WAX EXTRACT
C0022092|T121|5992|RXNORM|IRON-DEXTRAN COMPLEX|IRON-DEXTRAN COMPLEX
C2739945|T129|897499|RXNORM|SCOTCH BROOM POLLEN EXTRACT|CYTISUS SCOPARIUS POLLEN EXTRACT
C3256536|T121|1307769|RXNORM|FENUGREEK LEAF EXTRACT|FENUGREEK LEAF EXTRACT
C3256132|T109|1307768|RXNORM|COCCINIA GRANDIS FRUIT EXTRACT|COCCINIA GRANDIS FRUIT EXTRACT
C0172467|T121|61686|RXNORM|CLOSTEBOL|CLOSTEBOL
C0022432|T109|6086|RXNORM|JUNIPER TAR|JUNIPER TAR
C0022419|T195|6084|RXNORM|JOSAMYCIN|JOSAMYCIN
C0022431|T121|6085|RXNORM|JUNIPERUS COMMUNIS WHOLE EXTRACT|JUNIPERUS COMMUNIS WHOLE EXTRACT
C0057002|T129|22178|RXNORM|CYTOMEGALOVIRUS IMMUNE GLOBULIN|CYTOMEGALOVIRUS IMMUNE GLOBULIN
C2930113|T121|1000104|RXNORM|INCOBOTULINUMTOXIN A|INCOBOTULINUMTOXINA
C3256153|T109|1306144|RXNORM|CRANBERRY SEED OIL|CRANBERRY SEED OIL
C3256209|T109|1306145|RXNORM|CUCUMBER FRUIT OIL|CUCUMBER FRUIT OIL
C3256220|T109|1306146|RXNORM|CYMBOPOGON SCHOENANTHUS OIL|CYMBOPOGON SCHOENANTHUS OIL
C3255749|T109|1306148|RXNORM|CHINESE CINNAMON LEAF OIL|CHINESE CINNAMON LEAF OIL
C3255913|T109|1306149|RXNORM|CITRUS AURANTIFOLIA SEED OIL|CITRUS AURANTIFOLIA SEED OIL
C0063866|T121|27824|RXNORM|IRON SORBITEX|IRON SORBITEX
C0389169|T195|119771|RXNORM|DORIPENEM|DORIPENEM
C0008232|T121|2378|RXNORM|CHLOROBUTANOL|CHLOROBUTANOL
C0719082|T121|215815|RXNORM|CALAMINE / PHENOL|CALAMINE / PHENOL
C3256895|T121|1307640|RXNORM|AZADIRACHTA INDICA LEAF EXTRACT|AZADIRACHTA INDICA LEAF EXTRACT
C3256507|T121|1307641|RXNORM|BORAGO OFFICINALIS SEED EXTRACT|BORAGO OFFICINALIS SEED EXTRACT
C0063867|T121|27825|RXNORM|IRON SUCCINYL MILK PROTEIN COMPLEX|IRON SUCCINYL MILK PROTEIN COMPLEX
C3486713|T121|1311117|RXNORM|MAMMAL LIVER PREPARATION|MAMMAL LIVER PREPARATION
C3464706|T121|1307642|RXNORM|AVERRHOA CARAMBOLA LEAF EXTRACT|AVERRHOA CARAMBOLA LEAF EXTRACT
C1874634|T121|690832|RXNORM|CAFFEINE / PHENACETIN / SALICYLAMIDE / STYRAMATE|CAFFEINE / PHENACETIN / SALICYLAMIDE / STYRAMATE
C3464214|T121|1307643|RXNORM|WITHANIA SOMNIFERA FLOWER EXTRACT|WITHANIA SOMNIFERA FLOWER EXTRACT
C1874636|T121|690835|RXNORM|CALAMINE / CAMPHOR / DIPHENHYDRAMINE|CALAMINE / CAMPHOR / DIPHENHYDRAMINE
C1874637|T121|690836|RXNORM|CALAMINE / CAMPHOR / PRAMOXINE|CALAMINE / CAMPHOR / PRAMOXINE
C0013136|T121|3648|RXNORM|DROPERIDOL|DROPERIDOL
C3465270|T121|1307644|RXNORM|ECLIPTA PROSTRATA LEAF EXTRACT|ECLIPTA PROSTRATA LEAF EXTRACT
C0013092|T121|3642|RXNORM|DOXYLAMINE|DOXYLAMINE
C2926870|T121|1001472|RXNORM|DUTASTERIDE / TAMSULOSIN|DUTASTERIDE / TAMSULOSIN
C0013090|T195|3640|RXNORM|DOXYCYCLINE|DOXYCYCLINE
C0008806|T121|2550|RXNORM|CINOXACIN|CINOXACIN
C0008809|T121|2551|RXNORM|CIPROFLOXACIN|CIPROFLOXACIN
C0008809|T121|2551|RXNORM|CIPROFLOXACIN|CIPROFLOXACIN
C0008809|T121|2551|RXNORM|CIPROFLOXACIN|CIPROFLOXACIN
C3818684|T109|1537909|RXNORM|POLYGLUCOSE SORBITOL CARBOXYMETHYL ETHER|POLYGLUCOSE SORBITOL CARBOXYMETHYL ETHER
C0008838|T197|2555|RXNORM|CISPLATIN|CISPLATIN
C0008845|T121|2556|RXNORM|CITALOPRAM|CITALOPRAM
C3256181|T121|1307647|RXNORM|QUERCUS ROBUR TWIG BARK EXTRACT|QUERCUS ROBUR TWIG BARK EXTRACT
C2701808|T129|852806|RXNORM|SALT CEDAR POLLEN EXTRACT|TAMARIX GALLICA POLLEN EXTRACT
C0043611|T121|11476|RXNORM|TILUDRONIC ACID|TILUDRONIC ACID
C1720377|T121|645114|RXNORM|MICONAZOLE / PETROLATUM / ZINC OXIDE|MICONAZOLE / PETROLATUM / ZINC OXIDE
C0043603|T121|11473|RXNORM|PAMIDRONATE|PAMIDRONATE
C0770575|T121|235494|RXNORM|POTASSIUM CITRATE / SODIUM CITRATE|POTASSIUM CITRATE / SODIUM CITRATE
C1684405|T121|623033|RXNORM|LUBIPROSTONE|LUBIPROSTONE
C2927813|T121|1006889|RXNORM|DIMETHICONE / MENTHOL / PRAMOXINE|DIMETHICONE / MENTHOL / PRAMOXINE
C2740624|T129|899424|RXNORM|GRAPEFRUIT ALLERGENIC EXTRACT|CITRUS PARADISI ALLERGENIC EXTRACT
C2026329|T121|1006881|RXNORM|BROMHEXINE / CEPHALEXIN|BROMHEXINE / CEPHALEXIN
C2927806|T121|1006882|RXNORM|TRICLOSAN / VITAMIN E|TRICLOSAN / VITAMIN E
C2927807|T121|1006883|RXNORM|PIRENZEPINE / RANITIDINE|PIRENZEPINE / RANITIDINE
C2927808|T121|1006884|RXNORM|CARBOXYMETHYLCELLULOSE / DANTHRON / POLOXAMER|CARBOXYMETHYLCELLULOSE / DANTHRON / POLOXAMER
C2927809|T121|1006885|RXNORM|BROMHEXINE / ERYTHROMYCIN|BROMHEXINE / ERYTHROMYCIN
C2927810|T121|1006886|RXNORM|PHENYLEPHRINE / ZINC OXIDE|PHENYLEPHRINE / ZINC OXIDE
C0663182|T129|190353|RXNORM|DACLIZUMAB|DACLIZUMAB
C3834064|T109|1541886|RXNORM|PEG-8 PROPYLHEPTYL ETHER|PEG-8 PROPYLHEPTYL ETHER
C3715225|T109|1541884|RXNORM|GARDENIA JASMINOIDES WHOLE EXTRACT|GARDENIA JASMINOIDES WHOLE EXTRACT
C3834065|T109|1541885|RXNORM|PPG-26|PPG-26
C3715198|T109|1541882|RXNORM|ARTEMISIA VULGARIS WHOLE EXTRACT|ARTEMISIA VULGARIS WHOLE EXTRACT
C3834066|T109|1541883|RXNORM|CNIDIUM OFFICINALE ROOT OIL|CNIDIUM OFFICINALE ROOT OIL
C3834067|T109|1541881|RXNORM|ANGELICA GIGAS ROOT OIL|ANGELICA GIGAS ROOT OIL
C0050962|T121|17145|RXNORM|MONOBENZONE|MONOBENZONE
C0046237|T121|1363608|RXNORM|HYDROXYPROPYLBETADEX (0.58-0.68 MS)|HYDROXYPROPYLBETADEX (0.58-0.68 MS)
C2346446|T121|1363609|RXNORM|HYPNEA MUSCIFORMIS EXTRACT|HYPNEA MUSCIFORMIS EXTRACT
C0060583|T121|25193|RXNORM|FLUPIRTINE|FLUPIRTINE
C0016157|T121|4419|RXNORM|FISH OILS|FISH OILS
C3256041|T109|1363602|RXNORM|DIISOSTEARYL MALATE|DIISOSTEARYL MALATE
C3256042|T109|1363603|RXNORM|DILSEA CARNOSA EXTRACT|DILSEA CARNOSA EXTRACT
C0627405|T130|1363600|RXNORM|DIISOPROPYL ADIPATE|DIISOPROPYL ADIPATE
C0164628|T121|1363601|RXNORM|DIISOPROPYL SEBACATE|DIISOPROPYL SEBACATE
C3256047|T121|1363606|RXNORM|HYDROXYMETHYL CELLULOSE|HYDROXYMETHYL CELLULOSE
C3257245|T121|1363607|RXNORM|HYDROXYPROPYL CORN STARCH (5% SUBSTITUTION BY WEIGHT)|HYDROXYPROPYL CORN STARCH (5% SUBSTITUTION BY WEIGHT)
C3256045|T121|1363604|RXNORM|HYDROXYETHYL CELLULOSE (3000 CPS AT 1%)|HYDROXYETHYL CELLULOSE (3000 CPS AT 1%)
C3257244|T121|1363605|RXNORM|HYDROXYETHYL UREA|HYDROXYETHYL UREA
C3154026|T121|1100741|RXNORM|CALCIUM CHLORIDE / ICODEXTRIN / LACTATE / MAGNESIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CHLORIDE / ICODEXTRIN / LACTATE / MAGNESIUM CHLORIDE / SODIUM CHLORIDE
C0770213|T125|235279|RXNORM|INSULIN, PROTAMINE ZINC, PORK|INSULIN, PROTAMINE ZINC, PORK
C0770209|T125|235278|RXNORM|INSULIN, PROTAMINE ZINC, BEEF|INSULIN, PROTAMINE ZINC, BEEF
C0770201|T125|235275|RXNORM|INSULIN, REGULAR, BEEF-PORK|INSULIN, REGULAR, BEEF-PORK
C0770199|T197|235273|RXNORM|CALCIUM IODIDE|CALCIUM IODIDE
C0770198|T121|235272|RXNORM|IRON,PEPTONIZED|IRON,PEPTONIZED
C0770197|T197|235271|RXNORM|FERROUS CACODYLATE|FERROUS CACODYLATE
C0890177|T121|1368896|RXNORM|LINALOOL, (+-)-|LINALOOL, (+-)-
C3256558|T109|1368894|RXNORM|POLYETHYLENE GLYCOL 35000|POLYETHYLENE GLYCOL 35000
C3256634|T109|1368895|RXNORM|POLYISOBUTYLENE (1000 MW)|POLYISOBUTYLENE (1000 MW)
C3256107|T109|1368892|RXNORM|HYPROMELLOSE PHTHALATE (31% PHTHALATE, 40 CST)|HYPROMELLOSE PHTHALATE (31% PHTHALATE, 40 CST)
C3256555|T109|1368893|RXNORM|POLYETHYLENE GLYCOL 14000|POLYETHYLENE GLYCOL 14000
C2702386|T129|1297529|RXNORM|EASTERN YELLOWJACKET VENOM PROTEIN|VESPULA MACULIFRONS VENOM PROTEIN
C3256106|T109|1368891|RXNORM|HYPROMELLOSE PHTHALATE (31% PHTHALATE, 170 CST)|HYPROMELLOSE PHTHALATE (31% PHTHALATE, 170 CST)
C2702389|T129|1297527|RXNORM|COMMON WASP VENOM PROTEIN|VESPULA VULGARIS VENOM PROTEIN
C0440460|T129|1297525|RXNORM|BALD-FACED HORNET VENOM PROTEIN|DOLICHOVESPULA MACULATA VENOM PROTEIN
C0074445|T122|1368898|RXNORM|SHELLAC|SHELLAC
C1814800|T121|1364386|RXNORM|OCTYLDODECYL NEOPENTANOATE|OCTYLDODECYL NEOPENTANOATE
C1743069|T121|1364387|RXNORM|O-CYMEN-5-OL|O-CYMEN-5-OL
C0032397|T109|1364384|RXNORM|POLOXAMER 338|POLOXAMER 338
C1695071|T121|1364385|RXNORM|CERAMIDE 1|CERAMIDE 1
C1615089|T121|1364382|RXNORM|LAURYL GLUCOSIDE|LAURYL GLUCOSIDE
C0032476|T109|1364383|RXNORM|POLYETHYLENE GLYCOL 2000|POLYETHYLENE GLYCOL 2000
C1576833|T121|1364380|RXNORM|POLYGLYCERYL-3 DIISOSTEARATE|POLYGLYCERYL-3 DIISOSTEARATE
C1576843|T121|1364381|RXNORM|CETYL RICINOLEATE|CETYL RICINOLEATE
C1875540|T121|705034|RXNORM|NITROGEN / OXYGEN|NITROGEN / OXYGEN
C3643656|T121|1423473|RXNORM|HEPTANOIC ACID / LACTATE|HEPTANOIC ACID / LACTATE
C1875535|T121|705033|RXNORM|NIACIN / RIBOFLAVIN / THIAMINE|NIACIN / RIBOFLAVIN / THIAMINE
C3818792|T121|1491001|RXNORM|ISOBORNYL METHACRYLATE|ISOBORNYL METHACRYLATE
C3818791|T122|1491002|RXNORM|CETYL DIMETHICONE 45|CETYL DIMETHICONE 45
C1365976|T121|1310168|RXNORM|QUASSIA AMARA WOOD EXTRACT|QUASSIA
C0057803|T109|1491007|RXNORM|DIBUTYL MALEATE|DIBUTYL MALEATE
C3818790|T109|1491008|RXNORM|AMINOMETHYLPROPANOL (PERFLUORO-C6-C12 ETHYL)PHOSPHATE|AMINOMETHYLPROPANOL (PERFLUORO-C6-C12 ETHYL)PHOSPHATE
C1696547|T121|616877|RXNORM|MECASERMIN RINFABATE|MECASERMIN RINFABATE
C3487980|T121|1310167|RXNORM|TABEBUIA IMPETIGINOSA BARK EXTRACT|HANDROANTHUS IMPETIGINOSUS BARK EXTRACT
C3249216|T121|1234471|RXNORM|ASCORBIC ACID / CHOLECALCIFEROL / NIACIN / RIBOFLAVIN / SODIUM FLUORIDE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN E|ASCORBIC ACID / CHOLECALCIFEROL / NIACIN / RIBOFLAVIN / SODIUM FLUORIDE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN E
C3487973|T121|1310161|RXNORM|JUNIPERUS SABINA LEAF|JUNIPERUS SABINA LEAF
C0874161|T121|260101|RXNORM|OSELTAMIVIR|OSELTAMIVIR
C3486620|T121|1310162|RXNORM|CHRYSANTHELLUM INDICUM SUBSP. AFROAMERICANUM EXTRACT|CHRYSANTHELLUM INDICUM SUBSP. AFROAMERICANUM EXTRACT
C0066249|T109|1313237|RXNORM|METHYL HEPTINE CARBONATE|METHYL HEPTINE CARBONATE
C0453273|T121|125933|RXNORM|CRANBERRY PREPARATION|CRANBERRY PREPARATION
C0063865|T121|27823|RXNORM|IRON PROTEIN SUCCINYLATE|IRON PROTEIN SUCCINYLATE
C3194707|T121|1116982|RXNORM|AMERICAN HOUSE DUST MITE EXTRACT / EUROPEAN HOUSE DUST MITE EXTRACT|AMERICAN HOUSE DUST MITE EXTRACT / EUROPEAN HOUSE DUST MITE EXTRACT
C2364551|T129|805551|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-URUGUAY-716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-URUGUAY-716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN
C2928055|T121|1007133|RXNORM|COAL TAR / SALICYLIC ACID / SULFUR,COLLOIDAL|COAL TAR / SALICYLIC ACID / SULFUR,COLLOIDAL
C2928054|T121|1007132|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 11 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 16 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 6 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 11 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 16 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 6 VACCINE
C2928053|T121|1007131|RXNORM|MECLIZINE / VITAMIN B6|MECLIZINE / VITAMIN B6
C2928052|T121|1007130|RXNORM|ACETAMINOPHEN / DEXBROMPHENIRAMINE / PHENYLEPHRINE|ACETAMINOPHEN / DEXBROMPHENIRAMINE / PHENYLEPHRINE
C2928059|T121|1007137|RXNORM|BEE POLLEN / KOREAN GINSENG PREPARATION / ROYAL JELLY|BEE POLLEN / KOREAN GINSENG PREPARATION / ROYAL JELLY
C2928058|T121|1007136|RXNORM|PASSIFLORA INCARNATA EXTRACT / VALERIAN ROOT EXTRACT|PASSIFLORA INCARNATA EXTRACT / VALERIAN ROOT EXTRACT
C2928057|T121|1007135|RXNORM|DYCLONINE / MENTHOL|DYCLONINE / MENTHOL
C2928056|T121|1007134|RXNORM|ESTROGENS, CONJUGATED (USP) / METHYLTESTOSTERONE|ESTROGENS, CONJUGATED (USP) / METHYLTESTOSTERONE
C2928061|T121|1007139|RXNORM|BELLADONNA ALKALOIDS / CAFFEINE|BELLADONNA ALKALOIDS / CAFFEINE
C2928060|T121|1007138|RXNORM|PHENYLEPHRINE / SHARK LIVER OIL|PHENYLEPHRINE / SHARK LIVER OIL
C2710480|T109|1309260|RXNORM|THEOBROMA GRANDIFLORUM SEED EXTRACT|THEOBROMA GRANDIFLORUM SEED EXTRACT
C3535896|T121|1370584|RXNORM|MYRISTOYL GLUTAMATE|MYRISTOYL GLUTAMATE
C0164674|T126|59768|RXNORM|PEGADEMASE BOVINE|PEGADEMASE
C0885824|T121|317687|RXNORM|THUJA OCCIDENTALIS PREPARATION|THUJA OCCIDENTALIS PREPARATION
C0164662|T121|59763|RXNORM|STAVUDINE|STAVUDINE
C0982068|T121|314546|RXNORM|CERIUM OXALATE|CERIUM OXALATE
C0068314|T195|31435|RXNORM|VALRUBICIN|VALRUBICIN
C0068314|T195|31435|RXNORM|VALRUBICIN|VALRUBICIN
C0065636|T130|29256|RXNORM|MANDELIC ACID|MANDELIC ACID
C0056603|T197|21842|RXNORM|CUPROUS OXIDE|CUPROUS OXIDE
C2928775|T121|1007861|RXNORM|BANANA EXTRACT / POTASSIUM / WATERMELON PREPARATION|BANANA EXTRACT / POTASSIUM / WATERMELON PREPARATION
C2928774|T121|1007860|RXNORM|PHENYLEHRINE / ZINC SULFATE|PHENYLEHRINE / ZINC SULFATE
C2928777|T121|1007863|RXNORM|BROMHEXINE / OXELADIN|BROMHEXINE / OXELADIN
C2928776|T121|1007862|RXNORM|GINKGO BILOBA LEAF EXTRACT / VINCAMINE|GINKGO BILOBA LEAF EXTRACT / VINCAMINE
C2928605|T121|1007689|RXNORM|CHYMOTRYPSIN / PAPAIN / TRYPSIN|CHYMOTRYPSIN / PAPAIN / TRYPSIN
C2928604|T121|1007688|RXNORM|CYPROHEPTADINE / VITAMIN B 12|CYPROHEPTADINE / VITAMIN B 12
C2928780|T121|1007866|RXNORM|CHLOROPHYLLIN / SOYBEAN OIL|CHLOROPHYLLIN / SOYBEAN OIL
C2928601|T121|1007685|RXNORM|EUCALYPTUS EXTRACT / MENTHOL|EUCALYPTUS EXTRACT / MENTHOL
C2928600|T121|1007684|RXNORM|GLYCOL SALICYLATE / NONIVAMIDE / SALICYLIC ACID|GLYCOL SALICYLATE / NONIVAMIDE / SALICYLIC ACID
C2928603|T121|1007687|RXNORM|DEQUALINIUM / TETRACAINE|DEQUALINIUM / TETRACAINE
C2928602|T121|1007686|RXNORM|CHLORPHENIRAMINE / CHLORTHENOXAZIN|CHLORPHENIRAMINE / CHLORTHENOXAZIN
C2928597|T121|1007681|RXNORM|ACETAMINOPHEN / PROPYPHENAZONE|ACETAMINOPHEN / PROPYPHENAZONE
C2928599|T121|1007683|RXNORM|HYDROCORTISONE / LIDOCAINE / PROCYANIDOLIC OLIGOMER|HYDROCORTISONE / LIDOCAINE / PROCYANIDOLIC OLIGOMER
C2928598|T121|1007682|RXNORM|CHLORHEXIDINE / FELYPRESSIN|CHLORHEXIDINE / FELYPRESSIN
C3700908|T109|1485539|RXNORM|LAURAMIDOPROPYL DIMETHYLAMINE|LAURAMIDOPROPYL DIMETHYLAMINE
C3700909|T109|1485538|RXNORM|ERODIUM STEPHANIANUM TOP EXTRACT|ERODIUM STEPHANIANUM TOP EXTRACT
C3531069|T168|1366027|RXNORM|CARROT JUICE|CARROT JUICE
C2954288|T121|1047471|RXNORM|FLUNIXIN / OXYTETRACYCLINE|FLUNIXIN / OXYTETRACYCLINE
C1875504|T121|691286|RXNORM|MINERAL OIL / PETROLATUM|MINERAL OIL / PETROLATUM
C1875504|T121|691286|RXNORM|MINERAL OIL / PETROLATUM|MINERAL OIL / PETROLATUM
C0300903|T195|995897|RXNORM|ORBIFLOXACIN|ORBIFLOXACIN
C3700910|T109|1485537|RXNORM|PERIPLOCA SEPIUM ROOT BARK EXTRACT|PERIPLOCA SEPIUM ROOT BARK EXTRACT
C0031562|T123|1362735|RXNORM|PHLORHIZIN|PHLORHIZIN
C0046056|T130|1362737|RXNORM|FLUORODEOXYGLUCOSE F18|FLUDEOXYGLUCOSE (18F)
C0046563|T121|1362739|RXNORM|2-TERT-BUTYLHYDROQUINONE|2-TERT-BUTYLHYDROQUINONE
C0046404|T121|1362738|RXNORM|2-N-OCTYL-4-ISOTHIAZOLIN-3-ONE|OCTHILINONE
C0070895|T121|33562|RXNORM|FOSCARNET|FOSCARNET
C0981864|T129|892547|RXNORM|CORN ALLERGENIC EXTRACT|ZEA MAYS ALLERGENIC EXTRACT
C3474011|T109|1314268|RXNORM|ASCORBYL METHYLSILANOL PECTINATE|ASCORBYL METHYLSILANOL PECTINATE
C3496661|T121|1314269|RXNORM|BIS-PEG-18 METHYL ETHER DIMETHYL SILANE|BIS-PEG-18 METHYL ETHER DIMETHYL SILANE
C3474464|T121|1311562|RXNORM|BIDENS BIPINNATA TOP EXTRACT|BIDENS BIPINNATA TOP EXTRACT
C0030866|T109|1311563|RXNORM|PENTANE|PENTANE
C0068988|T121|1311560|RXNORM|NORFLURANE|NORFLURANE
C2961394|T121|1311561|RXNORM|OCIMUM TENUIFLORUM TOP EXTRACT|OCIMUM TENUIFLORUM TOP EXTRACT
C0301527|T121|89903|RXNORM|POTASSIUM GLUCONATE|POTASSIUM GLUCONATE
C0075618|T121|1311567|RXNORM|SULISOBENZONE|SULISOBENZONE
C0982053|T121|1311564|RXNORM|CANDELILLA WAX|CANDELILLA WAX
C0033472|T131|1311565|RXNORM|PROPIOLACTONE|PROPIOLACTONE
C0066561|T121|30031|RXNORM|MINAPRINE|MINAPRINE
C0379881|T195|115552|RXNORM|TROVAFLOXACIN|TROVAFLOXACIN
C1959878|T121|729743|RXNORM|SODIUM FLUORIDE / TRICLOSAN|SODIUM FLUORIDE / TRICLOSAN
C0031184|T121|8076|RXNORM|PERPHENAZINE|PERPHENAZINE
C3710173|T121|1489196|RXNORM|BETAINE SALICYLATE|BETAINE SALICYLATE
C2929368|T121|1008464|RXNORM|AMINOPHYLLINE / PROMETHAZINE|AMINOPHYLLINE / PROMETHAZINE
C2929369|T121|1008465|RXNORM|RESERPINE / XIPAMIDE|RESERPINE / XIPAMIDE
C2929370|T121|1008466|RXNORM|ALANINE / ARGININE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / PROLINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / PROLINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929371|T121|1008467|RXNORM|CRANBERRY PREPARATION / MILK THISTLE EXTRACT|CRANBERRY PREPARATION / MILK THISTLE EXTRACT
C2929364|T121|1008460|RXNORM|ETHANOLAMINE / FRAMYCETIN|ETHANOLAMINE / FRAMYCETIN
C2929365|T121|1008461|RXNORM|BACITRACIN / BENZOCAINE / TYROTHRICIN|BACITRACIN / BENZOCAINE / TYROTHRICIN
C2929366|T121|1008462|RXNORM|DIBUCAINE / PHENYLBUTAZONE|DIBUCAINE / PHENYLBUTAZONE
C2929367|T121|1008463|RXNORM|METOPROLOL / NIFEDIPINE|METOPROLOL / NIFEDIPINE
C2740787|T129|899724|RXNORM|CLOVE ALLERGENIC EXTRACT|CLOVE ALLERGENIC EXTRACT
C2929372|T121|1008468|RXNORM|ASCORBIC ACID / CALCIUM SULFATE / CHOLECALCIFEROL / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / KELP PREPARATION / MAGNESIUM OXIDE / MAGNESIUM SULFATE / NIACINAMIDE / POTASSIUM SULFATE / PYRIDOXINE / RIBOFLAVIN / VITAMIN A / VITAMIN B 12 / ZINC SULFATE|ASCORBIC ACID / CALCIUM SULFATE / CHOLECALCIFEROL / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / KELP PREPARATION / MAGNESIUM OXIDE / MAGNESIUM SULFATE / NIACINAMIDE / POTASSIUM SULFATE / PYRIDOXINE / RIBOFLAVIN / VITAMIN A / VITAMIN B 12 / ZINC SULFATE
C0360534|T121|108088|RXNORM|ALCLOMETASONE|ALCLOMETASONE
C0003818|T196|1111|RXNORM|ARSENIC|ARSENIC
C2006144|T121|813927|RXNORM|CALCIUM LACTATE / THIAMINE|CALCIUM LACTATE / THIAMINE
C2080534|T121|815008|RXNORM|NAPHAZOLINE / PHENYLEPHRINE|NAPHAZOLINE / PHENYLEPHRINE
C3819174|T121|1534422|RXNORM|ASPIRIN / CARBIDOPA|ASPIRIN / CARBIDOPA
C1720618|T121|645422|RXNORM|AMMONIUM CHLORIDE / CAFFEINE|AMMONIUM CHLORIDE / CAFFEINE
C3486712|T109|1352522|RXNORM|HYPERICUM OIL|HYPERICUM OIL
C0109105|T121|47907|RXNORM|CETALKONIUM CHLORIDE|CETALKONIUM CHLORIDE
C3486605|T121|1352520|RXNORM|GUAIACUM OFFICINALE RESIN EXTRACT|GUAIACUM OFFICINALE RESIN
C2073890|T121|815003|RXNORM|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / PSEUDOEPHEDRINE
C1436328|T121|461016|RXNORM|ESZOPICLONE|ESZOPICLONE
C2194002|T121|815321|RXNORM|DYPHYLLINE / POTASSIUM IODIDE|DYPHYLLINE / POTASSIUM IODIDE
C3253985|T121|1433868|RXNORM|DOLUTEGRAVIR|DOLUTEGRAVIR
C3281540|T121|1249101|RXNORM|BISMUTH SUBSALICYLATE / KAOLIN|BISMUTH SUBSALICYLATE / KAOLIN
C2740859|T129|899895|RXNORM|PINEAPPLE ALLERGENIC EXTRACT|ACCA SELLOWIANA ALLERGENIC EXTRACT
C0022124|T130|1364896|RXNORM|ISETHIONIC ACID|ISETHIONIC ACID
C0014834|T007|350202|RXNORM|ESCHERICHIA COLI|ESCHERICHIA COLI
C1874413|T121|692572|RXNORM|BACITRACIN / NEOMYCIN / POLYMYXIN B|BACITRACIN / NEOMYCIN / POLYMYXIN B
C1874413|T121|692572|RXNORM|BACITRACIN / NEOMYCIN / POLYMYXIN B|BACITRACIN / NEOMYCIN / POLYMYXIN B
C0062212|T121|26506|RXNORM|HEME ARGINATE|HEME ARGINATE
C1874408|T121|692570|RXNORM|BACITRACIN / DIPERODON / NEOMYCIN / POLYMYXIN B|BACITRACIN / DIPERODON / NEOMYCIN / POLYMYXIN B
C3256766|T121|1311596|RXNORM|GLEDITSIA SINENSIS FRUIT EXTRACT|GLEDITSIA SINENSIS FRUIT EXTRACT
C3486695|T121|1311595|RXNORM|GARCINIA CAMBOGIA FRUIT EXTRACT|GARCINIA GUMMI-GUTTA FRUIT EXTRACT
C0244656|T121|72236|RXNORM|FOSPHENYTOIN|FOSPHENYTOIN
C0076612|T121|38221|RXNORM|THYMALFASIN|THYMALFASIN
C0058263|T121|1311593|RXNORM|DIMETHYLDODECYLBENZYLAMMONIUM|BENZODODECINIUM
C3475281|T109|1313736|RXNORM|C12-14 PARETH-12|C12-14 PARETH-12
C0016778|T121|4582|RXNORM|TEGAFUR|TEGAFUR
C3537684|T121|1371300|RXNORM|CHICKORY ROOT EXTRACT|CHICORY ROOT EXTRACT
C1508750|T121|480639|RXNORM|ALVIMOPAN|ALVIMOPAN
C3537686|T121|1371302|RXNORM|PTYCHOPETALUM OLACOIDES WOOD EXTRACT|PTYCHOPETALUM OLACOIDES WOOD EXTRACT
C3537687|T121|1371303|RXNORM|PEG-9 POLYDIMETHYLSILOXYETHYL DIMETHICONE|PEG-9 POLYDIMETHYLSILOXYETHYL DIMETHICONE
C0981992|T129|852659|RXNORM|WESTERN WHEATGRASS POLLEN EXTRACT|PASCOPYRUM SMITHII POLLEN EXTRACT
C3537689|T130|1371306|RXNORM|C.I. FOOD YELLOW 3 (FREE ACID)|C.I. FOOD YELLOW 3 (FREE ACID)
C0051466|T121|1371307|RXNORM|ALPHA-TERPINEOL|ALPHA-TERPINEOL
C3537690|T116|1371308|RXNORM|ALUMINUM HYDROXYIDE-GLYCINE (2:1)|ALUMINUM HYDROXYIDE-GLYCINE (2:1)
C2701327|T129|852124|RXNORM|FIVEHORN SMOTHERWEED POLLEN EXTRACT|BASSIA HYSSOPIFOLIA POLLEN EXTRACT
C3256617|T121|1311590|RXNORM|FORSYTHIA SUSPENSA FRUIT EXTRACT|FORSYTHIA SUSPENSA FRUIT EXTRACT
C0035976|T121|9500|RXNORM|RUTIN|RUTIN
C2701713|T129|852653|RXNORM|EUROPEAN OLIVE POLLEN EXTRACT|OLEA EUROPAEA POLLEN EXTRACT
C2928982|T121|1008072|RXNORM|CHLORAMPHENICOL / COLLAGENASE|CHLORAMPHENICOL / COLLAGENASE
C2928981|T121|1008071|RXNORM|FUMARATE / NICKEL SULFATE / POTASSIUM BROMIDE|FUMARATE / NICKEL SULFATE / POTASSIUM BROMIDE
C2928980|T121|1008070|RXNORM|CAPSAICIN / TURPENTINE|CAPSAICIN / TURPENTINE
C2928986|T121|1008077|RXNORM|ALUMINUM HYDROXIDE / MAGNESIUM OXIDE|ALUMINUM HYDROXIDE / MAGNESIUM OXIDE
C2928985|T121|1008076|RXNORM|BENZOCAINE / PYRILAMINE|BENZOCAINE / PYRILAMINE
C0376160|T121|114176|RXNORM|ZUCLOPENTHIXOL|ZUCLOPENTHIXOL
C2193830|T121|1008074|RXNORM|AMPICILLIN / CARBOCYSTEINE|AMPICILLIN / CARBOCYSTEINE
C2928988|T121|1008079|RXNORM|HOMATROPINE / IBUPROFEN|HOMATROPINE / IBUPROFEN
C2928987|T121|1008078|RXNORM|RACEPINEPHRINE / ZINC CHLORIDE|RACEPINEPHRINE / ZINC CHLORIDE
C2347624|T121|1369713|RXNORM|POMALIDOMIDE|POMALIDOMIDE
C3855347|T121|1547755|RXNORM|STEPHANIA TETRANDRA ROOT EXTRACT|STEPHANIA TETRANDRA ROOT EXTRACT
C0070122|T121|32937|RXNORM|PAROXETINE|PAROXETINE
C3538346|T121|1372577|RXNORM|EVENING PRIMROSE OIL / LINOLEATE|EVENING PRIMROSE OIL / LINOLEATE
C0982325|T121|1363621|RXNORM|PEG-8 DIOLEATE|PEG-8 DIOLEATE
C2929507|T121|1008607|RXNORM|ECHINACEA ANGUSTIFOLIA ROOT EXTRACT / GOLDEN SEAL ROOT|ECHINACEA ANGUSTIFOLIA ROOT EXTRACT / GOLDEN SEAL ROOT
C2740867|T129|899906|RXNORM|RASPBERRY ALLERGENIC EXTRACT|RUBUS IDAEUS ALLERGENIC EXTRACT
C3256599|T109|1307154|RXNORM|C20-40 PARETH-10|C20-40 PARETH-10
C3474160|T121|1307155|RXNORM|GLYCOL PALMITATE|GLYCOL PALMITATE
C3256344|T109|1307156|RXNORM|BUTYLPHENYL METHYLPROPIONAL|BUTYLPHENYL METHYLPROPIONAL
C3255930|T109|1307157|RXNORM|DI-PPG-3 MYRISTYL ETHER ADIPATE|DI-PPG-3 MYRISTYL ETHER ADIPATE
C3256793|T109|1307150|RXNORM|OOLONG TEA LEAF EXTRACT|OOLONG TEA LEAF EXTRACT
C3255704|T121|1307151|RXNORM|NELUMBO NUCIFERA FLOWER WAX|NELUMBO NUCIFERA FLOWER WAX
C1881892|T121|1307152|RXNORM|GLYCERYL CAPRYLATE|GLYCERYL MONOCAPRYLATE
C3256769|T121|1307153|RXNORM|GLUCOSYL STEVIOL|GLUCOSYL STEVIOL
C0165603|T121|60212|RXNORM|ATOVAQUONE|ATOVAQUONE
C3488916|T121|1309467|RXNORM|HOTTONIA PALUSTRIS FLOWER EXTRACT|HOTTONIA PALUSTRIS FLOWER EXTRACT
C3256044|T109|1309464|RXNORM|FAGUS SYLVATICA FLOWER BUD EXTRACT|FAGUS SYLVATICA FLOWER BUD EXTRACT
C0085424|T129|1309465|RXNORM|INTERLEUKIN-9|INTERLEUKIN-9
C3256725|T121|1309462|RXNORM|SAPONARIA OFFICINALIS ROOT EXTRACT|SAPONARIA OFFICINALIS ROOT EXTRACT
C3256727|T109|1309463|RXNORM|SAUSSUREA COSTUS ROOT EXTRACT|AUCKLANDIA COSTUS ROOT EXTRACT
C3256719|T109|1309460|RXNORM|SALVIA HISPANICA SEED EXTRACT|CHIA SEED EXTRACT
C3488969|T121|1309461|RXNORM|SAMBUCUS NIGRA SUBSP. CANADENSIS FLOWERING TOP EXTRACT|SAMBUCUS NIGRA SUBSP. CANADENSIS FLOWERING TOP EXTRACT
C1875796|T121|705067|RXNORM|SULFUR / ZINC OXIDE|SULFUR / ZINC OXIDE
C3488447|T121|1426419|RXNORM|LAMIUM ALBUM EXTRACT|WHITE NETTLE EXTRACT
C3255735|T121|1426418|RXNORM|HYDROGENATED SOYBEAN LECITHIN|HYDROGENATED SOYBEAN LECITHIN
C3488970|T121|1309468|RXNORM|SCHINUS MOLLE BARK EXTRACT|SCHINUS MOLLE BARK EXTRACT
C3255842|T109|1309469|RXNORM|HOUTTUYNIA CORDATA FLOWERING TOP EXTRACT|HOUTTUYNIA CORDATA FLOWERING TOP EXTRACT
C0301459|T129|89854|RXNORM|MUMPS SKIN TEST ANTIGEN|MUMPS SKIN TEST ANTIGEN
C0061202|T123|25696|RXNORM|GENISTEIN|GENISTEIN
C2756418|T129|968130|RXNORM|STEMPHYLIUM SARCINIFORME EXTRACT|STEMPHYLIUM SARCINIFORME EXTRACT
C0981816|T130|314301|RXNORM|ALBUMIN,IODINATED I-131 SERUM|ALBUMIN,IODINATED I-131 SERUM
C2741291|T129|900764|RXNORM|SCOTCH PINE POLLEN EXTRACT|PINUS SYLVESTRIS POLLEN EXTRACT
C3651724|T121|1430251|RXNORM|PHYLLOSTACHYS NIGRA SAP EXTRACT|PHYLLOSTACHYS NIGRA SAP EXTRACT
C0622984|T120|1430252|RXNORM|1-PHENYLAZO-2-NAPHTHYLAMINE|1-PHENYLAZO-2-NAPHTHYLAMINE
C0717756|T121|214553|RXNORM|ESTRADIOL / TESTOSTERONE|ESTRADIOL / TESTOSTERONE
C0718030|T121|214807|RXNORM|PSEUDOEPHEDRINE / TRIPROLIDINE|PSEUDOEPHEDRINE / TRIPROLIDINE
C0718029|T121|214806|RXNORM|PSEUDOEPHEDRINE / TERFENADINE|PSEUDOEPHEDRINE / TERFENADINE
C0717760|T121|214557|RXNORM|ETHINYL ESTRADIOL / ETHYNODIOL|ETHINYL ESTRADIOL / ETHYNODIOL
C0717758|T121|214555|RXNORM|ETANERCEPT|ETANERCEPT
C0982111|T127|314583|RXNORM|D-BIOTIN|D-BIOTIN
C0717762|T121|214559|RXNORM|ETHINYL ESTRADIOL / NORGESTIMATE|ETHINYL ESTRADIOL / NORGESTIMATE
C0717761|T121|214558|RXNORM|ETHINYL ESTRADIOL / LEVONORGESTREL|ETHINYL ESTRADIOL / LEVONORGESTREL
C3488475|T121|1341385|RXNORM|TEUCRIUM MARUM EXTRACT|TEUCRIUM MARUM EXTRACT
C3488471|T121|1341384|RXNORM|ARTEMISIA VULGARIS ROOT EXTRACT|ARTEMISIA VULGARIS ROOT EXTRACT
C3486632|T121|1309791|RXNORM|EUTROCHIUM PURPUREUM ROOT|EUTROCHIUM PURPUREUM ROOT
C3255598|T121|1309793|RXNORM|HAWTHORN LEAF WITH FLOWER EXTRACT|HAWTHORN LEAF WITH FLOWER EXTRACT
C3486599|T121|1309794|RXNORM|CERATOSTIGMA WILLMOTTIANUM FLOWER EXTRACT|CERATOSTIGMA WILLMOTTIANUM FLOWER EXTRACT
C3255599|T121|1309795|RXNORM|HEDERA HELIX LEAF EXTRACT|HEDERA HELIX LEAF EXTRACT
C3488180|T121|1309796|RXNORM|TABEBUIA HETEROPHYLLA BARK EXTRACT|TABEBUIA HETEROPHYLLA BARK EXTRACT
C3488183|T121|1309798|RXNORM|QUEBRACHO BARK EXTRACT|QUEBRACHO BARK EXTRACT
C0001041|T123|194|RXNORM|ACETYLCHOLINE|ACETYLCHOLINE
C0001047|T121|197|RXNORM|ACETYLCYSTEINE|ACETYLCYSTEINE
C0001047|T121|197|RXNORM|ACETYLCYSTEINE|ACETYLCYSTEINE
C0001047|T121|197|RXNORM|ACETYLCYSTEINE|ACETYLCYSTEINE
C0001040|T127|193|RXNORM|ACETYLCARNITINE|ACETYLCARNITINE
C0040933|T004|328140|RXNORM|TRICOPHYTON PREPARATION|TRICHOPHYTON (FUNGUS)
C1122975|T121|328141|RXNORM|ANGELICA SINENSIS PREPARATION|ANGELICA SINENSIS PREPARATION
C0056783|T121|21993|RXNORM|CYCLONIUM|CYCLONIUM
C0056780|T121|21990|RXNORM|CYCLOMETHYCAINE|CYCLOMETHYCAINE
C2756786|T121|1370435|RXNORM|GLYCYRRHIZA GLABRA EXTRACT|GLYCYRRHIZA GLABRA EXTRACT
C0085237|T121|42359|RXNORM|TOCAINIDE|TOCAINIDE
C2955472|T116|1370439|RXNORM|ALBUMIN MICROSPHERES, HUMAN|ALBUMIN MICROSPHERES, HUMAN
C2937472|T121|1009219|RXNORM|ALISKIREN / AMLODIPINE|ALISKIREN / AMLODIPINE
C0085228|T121|42355|RXNORM|FLUVOXAMINE|FLUVOXAMINE
C0538727|T121|140480|RXNORM|ICODEXTRIN|ICODEXTRIN
C0085217|T197|42351|RXNORM|LITHIUM CARBONATE|LITHIUM CARBONATE
C0051162|T121|17311|RXNORM|ALIZAPRIDE|ALIZAPRIDE
C1578240|T121|477364|RXNORM|SOLFENACIN|SOLFENACIN
C2698759|T121|1312715|RXNORM|PENTADECALACTONE|PENTADECALACTONE
C2929818|T121|1008921|RXNORM|CALCIUM CARBONATE / MAGNESIUM TRISILICATE|CALCIUM CARBONATE / MAGNESIUM TRISILICATE
C2929817|T121|1008920|RXNORM|ALUMINUM STEARATE / GUAIAZULENE / PENTOSAN POLYSULFATE|ALUMINUM STEARATE / GUAIAZULENE / PENTOSAN POLYSULFATE
C2929820|T121|1008923|RXNORM|INOSITOL / VITAMIN B6|INOSITOL / VITAMIN B6
C2929819|T121|1008922|RXNORM|BENDROFLUMETHIAZIDE / SPIRONOLACTONE|BENDROFLUMETHIAZIDE / SPIRONOLACTONE
C2929822|T121|1008925|RXNORM|GLUTAMATE / ZINC CHLORIDE|GLUTAMATE / ZINC CHLORIDE
C0039350|T123|10337|RXNORM|TAURINE|TAURINE
C2929824|T121|1008927|RXNORM|NIACIN / VITAMIN B6|NIACIN / VITAMIN B6
C2929823|T121|1008926|RXNORM|DEXTROMETHORPHAN / GUAIACOLSULFONATE|DEXTROMETHORPHAN / GUAIACOLSULFONATE
C2929826|T121|1008929|RXNORM|ALANINE / ARGININE / ASPARTATE / CALCIUM CHLORIDE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / ASPARTATE / CALCIUM CHLORIDE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C0028158|T196|7456|RXNORM|CHLOPHENIRAMINE|NITROGEN
C0030438|T121|7909|RXNORM|PARALDEHYDE|PARALDEHYDE
C1099045|T121|321650|RXNORM|IODINE / POTASSIUM IODIDE|IODINE / POTASSIUM IODIDE
C1099045|T121|321650|RXNORM|IODINE / POTASSIUM IODIDE|IODINE / POTASSIUM IODIDE
C0393080|T121|121243|RXNORM|VORICONAZOLE|VORICONAZOLE
C0030415|T122|7906|RXNORM|PARAFFIN|PARAFFIN
C2356014|T121|802546|RXNORM|CODEINE / DEXCHLORPHENIRAMINE / PHENYLEPHRINE|CODEINE / DEXCHLORPHENIRAMINE / PHENYLEPHRINE
C3530902|T121|1365710|RXNORM|CETEARETH-22|CETEARETH-22
C0771521|T121|236265|RXNORM|ISOMYRTOL|ISOMYRTOL
C3834235|T121|1543765|RXNORM|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-BRISBANE-60-2008 STRAIN|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-BRISBANE-60-2008 STRAIN
C0771526|T121|236268|RXNORM|BICLOTYMOL|BICLOTYMOL
C3531205|T109|1366320|RXNORM|ANGELICA BISERRATA ROOT EXTRACT|ANGELICA BISERRATA ROOT EXTRACT
C2364541|T129|805541|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-FLORIDA-4-2006 STRAIN|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-FLORIDA-4-2006 STRAIN
C0055402|T121|20823|RXNORM|CHLOROCRESOL|CHLOROCRESOL
C3486601|T121|1306351|RXNORM|CETRARIA ISLANDICA SUBSP. ISLANDICA EXTRACT|CETRARIA ISLANDICA SUBSP. ISLANDICA EXTRACT
C1509365|T121|1368901|RXNORM|ISOSTEARYL PALMITATE|ISOSTEARYL PALMITATE
C2723780|T129|867369|RXNORM|COMMON COCKLEBURR POLLEN EXTRACT|COMMON COCKLEBURR POLLEN EXTRACT
C2701360|T129|852158|RXNORM|RUSSIAN THISTLE POLLEN EXTRACT|SALSOLA KALI POLLEN EXTRACT
C3857951|T109|1552172|RXNORM|GUIZOTIA ABYSSINICA SEED OIL|GUIZOTIA ABYSSINICA SEED OIL
C3818775|T121|1492182|RXNORM|AGROPYRON FRAGILE WHOLE EXTRACT|AGROPYRON FRAGILE WHOLE EXTRACT
C0044487|T121|1425941|RXNORM|1-MYRISTYLPICOLINIUM|MIRIPIRIUM CHLORIDE
C1291212|T121|618278|RXNORM|AZELATE|AZELATE
C0392426|T121|121069|RXNORM|DIMETHOXANATE|DIMETHOXANATE
C1702726|T121|618272|RXNORM|FLUFENAMATE|FLUFENAMATE
C0772446|T121|237108|RXNORM|SODIUM ACETATE TRIHYDRATE|SODIUM ACETATE TRIHYDRATE
C0075632|T121|37418|RXNORM|SUMATRIPTAN|SUMATRIPTAN
C0873066|T121|259404|RXNORM|BARBERRY EXTRACT|BARBERRY EXTRACT
C0012403|T121|3455|RXNORM|DIMETHYL SULFOXIDE|DIMETHYL SULFOXIDE
C3486817|T121|1337635|RXNORM|OXALIS MONTANA LEAF EXTRACT|OXALIS MONTANA LEAF EXTRACT
C0057920|T121|22971|RXNORM|DIETHANOLAMINE FUSIDATE|DIETHANOLAMINE FUSIDATE
C2710464|T121|1426385|RXNORM|C18-36 ACID TRIGLYCERIDE|C18-36 ACID TRIGLYCERIDE
C3864825|T109|1597295|RXNORM|N,N-BIS(2-HYDROXYETHYL)LACTAMIDE|N,N-BIS(2-HYDROXYETHYL)LACTAMIDE
C0084528|T121|41996|RXNORM|SERTINDOLE|SERTINDOLE
C0062686|T121|26879|RXNORM|HEXYLCAINE|HEXYLCAINE
C3857949|T109|1552357|RXNORM|POLYGLYCERYL-3 DIOLEATE|POLYGLYCERYL-3 DIOLEATE
C2747700|T129|966979|RXNORM|PAECILOMYCES VARIOTII EXTRACT|PAECILOMYCES VARIOTII EXTRACT
C1258950|T109|1552358|RXNORM|HESPERADIN|HESPERADIN
C2920800|T129|999457|RXNORM|FUSARIUM COMPACTUM EXTRACT|FUSARIUM COMPACTUM EXTRACT
C3853725|T121|1597291|RXNORM|MYRTUS COMMUNIS WHOLE EXTRACT|MYRTUS COMMUNIS WHOLE EXTRACT
C2929579|T121|1008679|RXNORM|CAFFEINE / CARZENIDE / PROPYPHENAZONE|CAFFEINE / CARZENIDE / PROPYPHENAZONE
C2929578|T121|1008678|RXNORM|HEPTAMINOL / INOSITOL / RUTIN|HEPTAMINOL / INOSITOL / RUTIN
C0772206|T121|236881|RXNORM|BUTOXYCAINE|BUTOXYCAINE
C0772205|T121|236880|RXNORM|ETHYL HEXYL SALICYLATE|ETHYL HEXYL SALICYLATE
C3486564|T121|1310036|RXNORM|TSUGA CANADENSIS BARK EXTRACT|TSUGA CANADENSIS BARK EXTRACT
C2929571|T121|1008671|RXNORM|ANTIPYRINE / MEPROBAMATE / PAPAVERINE|ANTIPYRINE / MEPROBAMATE / PAPAVERINE
C2929570|T121|1008670|RXNORM|LAURETH-9 / UREA|POLIDOCANOL / UREA
C2929573|T121|1008673|RXNORM|ASCORBIC ACID / CALCIUM CITRATE / SILICON DIOXIDE|ASCORBIC ACID / CALCIUM CITRATE / SILICON DIOXIDE
C2929572|T121|1008672|RXNORM|DIBUCAINE / POLICRESULEN|DIBUCAINE / POLICRESULEN
C2929575|T121|1008675|RXNORM|CALCIUM PHOSPHATE / PICOLINIC ACID|CALCIUM PHOSPHATE / PICOLINIC ACID
C2929574|T121|1008674|RXNORM|CLIMBAZOLE / PIROCTONE OLAMINE|CLIMBAZOLE / PIROCTONE OLAMINE
C2929577|T121|1008677|RXNORM|LOPERAMIDE / PHTHALYLSULFACETAMIDE / PHTHALYLSULFATHIAZOLE|LOPERAMIDE / PHTHALYLSULFACETAMIDE / PHTHALYLSULFATHIAZOLE
C2929576|T121|1008676|RXNORM|ASCORBIC ACID / ZINC CITRATE|ASCORBIC ACID / ZINC CITRATE
C2194013|T121|818018|RXNORM|ATROPINE / EPINEPHRINE|ATROPINE / EPINEPHRINE
C0939900|T121|285246|RXNORM|PLANTAIN PREPARATION|PLANTAIN PREPARATION
C3834047|T109|1543742|RXNORM|BEEF TONGUE PREPARATION|BEEF TONGUE PREPARATION
C2168864|T121|818014|RXNORM|GUAIFENESIN / PYRILAMINE|GUAIFENESIN / PYRILAMINE
C1509274|T121|1311623|RXNORM|CETEARETH-30|CETEARETH-30
C0019134|T123|5224|RXNORM|HEPARIN|HEPARIN
C3256460|T109|1309480|RXNORM|TUSSILAGO FARFARA FLOWER EXTRACT|TUSSILAGO FARFARA FLOWER EXTRACT
C3256354|T109|1311622|RXNORM|CETEARETH-25|CETEARETH-25
C0772316|T121|236982|RXNORM|GREATER CELANDINE|GREATER CELANDINE
C1572598|T121|1311624|RXNORM|CETEARETH-6|CETEARETH-6
C2929486|T121|1008583|RXNORM|DANTHRON / POLOXAMER 188|DANTHRON / POLOXAMER 188
C2929485|T121|1008582|RXNORM|BETAINE / GLUTAMATE / OX BILE EXTRACT|BETAINE / GLUTAMATE / OX BILE EXTRACT
C2929483|T121|1008580|RXNORM|NALIDIXATE / PHENAZOPYRIDINE|NALIDIXATE / PHENAZOPYRIDINE
C2701174|T129|851934|RXNORM|WESTERN WATERHEMP POLLEN EXTRACT|AMARANTHUS TUBERCULATUS POLLEN EXTRACT
C2929489|T121|1008586|RXNORM|ANTHRALIN / SALICYLIC ACID|ANTHRALIN / SALICYLIC ACID
C2929488|T121|1008585|RXNORM|FERROUS FUMARATE / FOLIC ACID / POLYSACCHARIDE IRON COMPLEX|FERROUS FUMARATE / FOLIC ACID / POLYSACCHARIDE IRON COMPLEX
C2929487|T121|1008584|RXNORM|MELATONIN / VITAMIN B6|MELATONIN / VITAMIN B6
C0981880|T130|851938|RXNORM|FALSE RAGWEED POLLEN EXTRACT|AMBROSIA ACANTHICARPA POLLEN EXTRACT
C2929492|T121|1008589|RXNORM|OXELADIN / PROMETHAZINE|OXELADIN / PROMETHAZINE
C2929491|T121|1008588|RXNORM|CHROMOUS CHLORIDE / COPPER SULFATE / MANGANESE CHLORIDE / SELENIOUS ACID / SODIUM IODIDE / ZINC SULFATE|CHROMOUS CHLORIDE / COPPER SULFATE / MANGANESE CHLORIDE / SELENIOUS ACID / SODIUM IODIDE / ZINC SULFATE
C0051919|T121|17941|RXNORM|ANISINDIONE|ANISINDIONE
C3486725|T197|1311628|RXNORM|CUPRIC ARSENITE|CUPRIC ARSENITE
C0071304|T121|33910|RXNORM|ISRADIPINE|ISRADIPINE
C0052416|T197|18330|RXNORM|ARSENIC TRIOXIDE|ARSENIC TRIOXIDE
C3256495|T121|1372011|RXNORM|ACER SACCHARUM SAP EXTRACT|ACER SACCHARUM SAP EXTRACT
C3256206|T121|1372010|RXNORM|CRITHMUM MARITIMUM EXTRACT|CRITHMUM MARITIMUM EXTRACT
C3256685|T121|1372013|RXNORM|GELIDIELLA ACEROSA EXTRACT|GELIDIELLA ACEROSA EXTRACT
C3818783|T109|1491867|RXNORM|PIGMENT ORANGE 2|PIGMENT ORANGE 2
C3255700|T121|1307976|RXNORM|NOTOPTERYGIUM INCISUM ROOT EXTRACT|NOTOPTERYGIUM INCISUM ROOT EXTRACT
C3256788|T121|1307977|RXNORM|NELUMBO NUCIFERA LEAF EXTRACT|NELUMBO NUCIFERA LEAF EXTRACT
C3488926|T121|1307974|RXNORM|CNIDIUM OFFICINALE ROOT EXTRACT|CNIDIUM OFFICINALE ROOT EXTRACT
C3256994|T121|1307975|RXNORM|PAEONIA SUFFRUTICOSA ROOT EXTRACT|PAEONIA SUFFRUTICOSA ROOT EXTRACT
C3256196|T121|1307972|RXNORM|KALMIA LATIFOLIA LEAF|KALMIA LATIFOLIA LEAF
C1881920|T121|1307970|RXNORM|VERBASCUM DENSIFLORUM LEAF EXTRACT|MULLEIN LEAF EXTRACT
C3255879|T121|1307971|RXNORM|STEVIA REBAUDIUNA LEAF EXTRACT|STEVIA REBAUDIUNA LEAF EXTRACT
C3162437|T121|1114112|RXNORM|AZFICEL-T|AZFICEL-T
C3486865|T121|1310203|RXNORM|LEDUM PALUSTRE TWIG EXTRACT|RHODODENDRON TOMENTOSUM LEAFY TWIG EXTRACT
C3464705|T109|1313733|RXNORM|4-HYDROXY-2,5-DIMETHYLFURAN-2(3H)-ONE|DIMETHYLHYDROXY FURANONE
C3496033|T121|1311257|RXNORM|SUS SCROFA SPINAL CORD PREPARATION|PORCINE SPINAL CORD PREPARATION
C0732784|T121|226976|RXNORM|LIDOCAINE / PHENYLEPHRINE|LIDOCAINE / PHENYLEPHRINE
C3500636|T121|1314926|RXNORM|LYCOPERDON UTRIFORME FRUITING BODY EXTRACT|LYCOPERDON UTRIFORME FRUITING BODY EXTRACT
C1095878|T121|319799|RXNORM|ERYSIMUM PREPARATION|ERYSIMUM PREPARATION
C0002374|T197|615|RXNORM|ALUMINUM OXIDE|ALUMINIUM OXIDE
C3666442|T121|1436959|RXNORM|ISOSTEARIC DIETHANOLAMIDE|ISOSTEARIC DIETHANOLAMIDE
C2727177|T129|886638|RXNORM|CAT FLEA ALLERGENIC EXTRACT|CTENOCEPHALIDES FELIS ALLERGENIC EXTRACT
C3651697|T121|1428848|RXNORM|ADANSONIA DIGITATA LEAF EXTRACT|ADANSONIA DIGITATA LEAF EXTRACT
C3651767|T121|1428849|RXNORM|ADANSONIA DIGITATA SEED EXTRACT|ADANSONIA DIGITATA SEED EXTRACT
C3651771|T121|1428844|RXNORM|DIANTHUS CARYOPHYLLUS FLOWER EXTRACT|DIANTHUS CARYOPHYLLUS FLOWER EXTRACT
C3651770|T121|1428845|RXNORM|FICUS CARICA FLOWER EXTRACT|FICUS CARICA FLOWER EXTRACT
C3651769|T121|1428846|RXNORM|GARDEN SNAIL MUCIN PREPARATION|GARDEN SNAIL MUCIN PREPARATION
C3651768|T121|1428847|RXNORM|CUCUMIS MELO EXTRACT|CUCUMIS MELO EXTRACT
C1445375|T121|1428840|RXNORM|PSIDIUM GUAJAVA EXTRACT|PSIDIUM GUAJAVA EXTRACT
C3651773|T121|1428841|RXNORM|MORUS AUSTRALIS WOOD EXTRACT|MORUS AUSTRALIS WOOD EXTRACT
C3651772|T121|1428842|RXNORM|VIGNA RADIATA EXTRACT|VIGNA RADIATA EXTRACT
C1445784|T121|1428843|RXNORM|IRIS GERMANICA EXTRACT|IRIS GERMANICA EXTRACT
C2723725|T129|867311|RXNORM|LIVE OAK POLLEN EXTRACT|QUERCUS VIRGINIANA POLLEN EXTRACT
C2723729|T129|867315|RXNORM|RABBIT SKIN EXTRACT|RABBIT SKIN EXTRACT
C2186923|T121|815765|RXNORM|CLOPAMIDE / DIHYDROERGOCRISTINE / RESERPINE|CLOPAMIDE / DIHYDROERGOCRISTINE / RESERPINE
C2193892|T121|812260|RXNORM|ETHINYL ESTRADIOL / LYNESTRENOL|ETHINYL ESTRADIOL / LYNESTRENOL
C1329999|T121|404794|RXNORM|DIHYDROCODEINE / GUAIFENESIN / PSEUDOEPHEDRINE|DIHYDROCODEINE / GUAIFENESIN / PSEUDOEPHEDRINE
C2080566|T121|815946|RXNORM|ASCORBIC ACID / PHENYLPROPANOLAMINE|ASCORBIC ACID / PHENYLPROPANOLAMINE
C3856075|T121|1549545|RXNORM|DIHYDROSTREPTOMYCIN / PENICILLIN G|DIHYDROSTREPTOMYCIN / PENICILLIN G
C2701078|T129|851744|RXNORM|RED MAPLE POLLEN EXTRACT|RED MAPLE POLLEN EXTRACT
C0262967|T195|1549540|RXNORM|DIHYDROSTREPTOMYCIN|DIHYDROSTREPTOMYCIN
C2928394|T121|1007472|RXNORM|ASPIRIN / CHLORMEZANONE|ASPIRIN / CHLORMEZANONE
C2928395|T121|1007473|RXNORM|ESTRIOL / THYMOL / UREA|ESTRIOL / THYMOL / UREA
C2928392|T121|1007470|RXNORM|DI-ISOPROPYLAMMONIUM / OROTIC ACID|DI-ISOPROPYLAMMONIUM / OROTIC ACID
C2928393|T121|1007471|RXNORM|ALUMINUM HYDROXIDE / SIMETHICONE|ALUMINUM HYDROXIDE / SIMETHICONE
C2928398|T121|1007476|RXNORM|PENTAERYTHRITOL / PROPRANOLOL|PENTAERYTHRITOL / PROPRANOLOL
C2928399|T121|1007477|RXNORM|CODEINE / ETHYLMORPHINE|CODEINE / ETHYLMORPHINE
C2928396|T121|1007474|RXNORM|ETHINYL ESTRADIOL / NORGESTRIENONE|ETHINYL ESTRADIOL / NORGESTRIENONE
C2928397|T121|1007475|RXNORM|BENZALKONIUM / BENZOCAINE / HEXYLRESORCINOL|BENZALKONIUM / BENZOCAINE / HEXYLRESORCINOL
C3255874|T109|1367149|RXNORM|STEAROXYTRIMETHYLSILANE|STEAROXYTRIMETHYLSILANE
C2946981|T121|1040053|RXNORM|DEXTROMETHORPHAN / QUINIDINE|DEXTROMETHORPHAN / QUINIDINE
C2928401|T121|1007479|RXNORM|ACETIC ACID / BENZOCAINE|ACETIC ACID / BENZOCAINE
C3709926|T121|1488577|RXNORM|BIOTIN / PANTHENOL|BIOTIN / PANTHENOL
C0126000|T121|52106|RXNORM|LITHIUM GLUCONATE|LITHIUM GLUCONATE
C1875087|T121|691072|RXNORM|DYPHYLLINE / EPHEDRINE / GUAIFENESIN / PHENOBARBITAL|DYPHYLLINE / EPHEDRINE / GUAIFENESIN / PHENOBARBITAL
C0055468|T121|20881|RXNORM|CHLORPHENOXAMINE|CHLORPHENOXAMINE
C0024027|T121|6472|RXNORM|LOVASTATIN|LOVASTATIN
C0075061|T121|1546393|RXNORM|FOSINOPRILAT|FOSINOPRILAT
C0024002|T121|6470|RXNORM|LORAZEPAM|LORAZEPAM
C0024056|T121|6475|RXNORM|LOXAPINE|LOXAPINE
C0888195|T197|267798|RXNORM|DISODIUM PYROPHOSPHATE|DISODIUM PYROPHOSPHATE
C0773826|T121|237929|RXNORM|SENNA LEAVES|SENNA LEAVES
C2929529|T121|1008629|RXNORM|CARBINOXAMINE MALEATE / CARBINOXAMINE TANNATE|CARBINOXAMINE MALEATE / CARBINOXAMINE TANNATE
C0070072|T121|32894|RXNORM|PARAMETHADIONE|PARAMETHADIONE
C3848542|T196|1546392|RXNORM|CHLORITE ION|CHLORITE ION
C0053777|T122|19464|RXNORM|BISDEQUALINIUM|BISDEQUALINIUM
C0053774|T121|19461|RXNORM|BISABOLOL|BISABOLOL
C1828179|T121|687103|RXNORM|BENZOCAINE / CETYLPYRIDINIUM|BENZOCAINE / CETYLPYRIDINIUM
C0031937|T121|8332|RXNORM|PINDOLOL|PINDOLOL
C0031938|T121|8333|RXNORM|PINE TAR|PINE TAR
C0031935|T121|8331|RXNORM|PIMOZIDE|PIMOZIDE
C0025241|T121|6718|RXNORM|MELPHALAN|MELPHALAN
C0025242|T121|6719|RXNORM|MEMANTINE|MEMANTINE
C0031954|T121|8338|RXNORM|PIPERACETAZINE|PIPERACETAZINE
C0031955|T195|8339|RXNORM|PIPERACILLIN|PIPERACILLIN
C0043458|T123|1314423|RXNORM|ZEIN|ZEIN
C0304987|T197|91540|RXNORM|IODOHIPPURATE I131 SODIUM|IODOHIPPURATE I131 SODIUM
C0025219|T125|6711|RXNORM|MELATONIN|MELATONIN
C0317591|T007|100272|RXNORM|LACTOBACILLUS BULGARICUS|LACTOBACILLUS BULGARICUS
C1276887|T121|389179|RXNORM|FELODIPINE / RAMIPRIL|FELODIPINE / RAMIPRIL
C0302928|T197|1546391|RXNORM|CHLORIC ACID|CHLORIC ACID
C0317597|T007|100278|RXNORM|LACTOBACILLUS CASEI RHAMNOSUS|LACTOBACILLUS CASEI RHAMNOSUS
C0059703|T121|24464|RXNORM|ETHAVERINE|ETHAVERINE
C3645121|T121|1426628|RXNORM|METHYLESCULETIN ACETATE|METHYLESCULETIN ACETATE
C3535844|T121|1370649|RXNORM|LAURYL SULFOSUCCINATE|LAURYL SULFOSUCCINATE
C0059699|T121|24460|RXNORM|ETHANOLAMINE OLEATE|ETHANOLAMINE OLEATE
C0036774|T123|1426381|RXNORM|SERUM ALBUMIN, BOVINE|SERUM ALBUMIN, BOVINE
C3255976|T109|1426622|RXNORM|PROPYLENE GLYCOL DICAPRYLATE-DICAPRATE|PROPYLENE GLYCOL DICAPRYLATE-DICAPRATE
C3645117|T121|1426623|RXNORM|ISOPROPYL MALEATE|ISOPROPYL MALEATE
C3255977|T109|1426620|RXNORM|PROPYLENE GLYCOL DIETHYLHEXANOATE|PROPYLENE GLYCOL DIETHYLHEXANOATE
C0294713|T109|1426621|RXNORM|HYDROXYISOHEXYL 3-CYCLOHEXENE CARBOXALDEHYDE|HYDROXYISOHEXYL 3-CYCLOHEXENE CARBOXALDEHYDE
C3645119|T121|1426626|RXNORM|PALM KERNEL ACID|PALM KERNEL ACID
C0059708|T121|24468|RXNORM|ETHENZAMIDE|ETHENZAMIDE
C3645118|T121|1426624|RXNORM|PALM ACID|PALM ACID
C3256225|T109|1426625|RXNORM|DIMETHYLOCTADECYL(3-(TRIMETHOXYSILYL)PROPYL)AMMONIUM CHLORIDE|DIMETHYLOCTADECYL(3-(TRIMETHOXYSILYL)PROPYL)AMMONIUM CHLORIDE
C3265177|T121|1307741|RXNORM|RAPESEED STEROL EXTRACT|RAPESEED STEROL EXTRACT
C3255674|T121|1307740|RXNORM|HELIANTHUS ANNUUS SEED WAX EXTRACT|HELIANTHUS ANNUUS SEED WAX EXTRACT
C3255981|T121|1307743|RXNORM|SYZYGIUM JAMBOS LEAF EXTRACT|SYZYGIUM JAMBOS LEAF EXTRACT
C3256214|T121|1307742|RXNORM|CUSCUTA JAPONICA SEED EXTRACT|CUSCUTA JAPONICA SEED EXTRACT
C3255701|T121|1307745|RXNORM|NYMPHAEA ALBA FLOWER EXTRACT|NYMPHAEA ALBA FLOWER EXTRACT
C3473990|T109|1307744|RXNORM|ROSA GALLICA FLOWER OIL|ROSA GALLICA FLOWER OIL
C3257505|T121|1307747|RXNORM|HIBISCUS ROSA-SINENSIS LEAF EXTRACT|HIBISCUS ROSA-SINENSIS LEAF EXTRACT
C3255693|T121|1307746|RXNORM|LIPPIA CITRIODORA FLOWER EXTRACT|LIPPIA CITRIODORA FLOWER EXTRACT
C2349151|T121|1307749|RXNORM|SALIX ALBA BARK EXTRACT|WHITE WILLOW BARK EXTRACT
C3256269|T109|1307748|RXNORM|RICE OIL|RICE OIL
C0001002|T121|178|RXNORM|ACETONE|ACETONE
C2973446|T129|1147320|RXNORM|BRENTUXIMAB VEDOTIN|BRENTUXIMAB VEDOTIN
C0717307|T121|214128|RXNORM|ACETAMINOPHEN / BROMPHENIRAMINE / PHENYLPROPANOLAMINE|ACETAMINOPHEN / BROMPHENIRAMINE / PHENYLPROPANOLAMINE
C2057739|T121|813683|RXNORM|DEXAMETHASONE / THEOPHYLLINE|DEXAMETHASONE / THEOPHYLLINE
C0072540|T121|34930|RXNORM|PSEUDOISOCYTIDINE|PSEUDOISOCYTIDINE
C2047354|T121|813131|RXNORM|HYDROCHLOROTHIAZIDE / POTASSIUM CHLORIDE|HYDROCHLOROTHIAZIDE / POTASSIUM CHLORIDE
C3651745|T121|1429392|RXNORM|LIQUIDAMBAR FORMOSANA RESIN|LIQUIDAMBAR FORMOSANA RESIN
C3255642|T109|1306168|RXNORM|BALSAM FIR LEEFY TWIG EXTRACT|BALSAM FIR LEEFY TWIG EXTRACT
C3255643|T109|1306169|RXNORM|BAMBUSA ARUNDINACEA STEM EXTRACT|BAMBUSA ARUNDINACEA STEM EXTRACT
C0014758|T121|4040|RXNORM|ERYTHRITYL TETRANITRATE|ERITRITYL TETRANITRATE
C2189302|T121|816810|RXNORM|BROMAZEPAM / VERALIPRIDE|BROMAZEPAM / VERALIPRIDE
C0719098|T121|215831|RXNORM|CALCIUM CITRATE / VITAMIN D|CALCIUM CITRATE / VITAMIN D
C0719097|T121|215830|RXNORM|CALCIUM CARBONATE / VITAMIN D|CALCIUM CARBONATE / VITAMIN D
C1879986|T168|1306162|RXNORM|CAMELLIA OIL|CAMELLIA OIL
C3256753|T109|1306163|RXNORM|CAMPHOR LEAF OIL|CAMPHOR LEAF OIL
C3256665|T109|1306160|RXNORM|CALOPHYLLUM TACAMAHACA SEED OIL|CALOPHYLLUM TACAMAHACA SEED OIL
C3256669|T109|1306161|RXNORM|CAMELLIA JAPONICA SEED OIL|CAMELLIA JAPONICA SEED OIL
C2948039|T121|1306166|RXNORM|ARNICA MONTANA FLOWER EXTRACT|ARNICA MONTANA FLOWER EXTRACT
C2949322|T121|1306167|RXNORM|ANGELICA DAHURICA ROOT EXTRACT|ANGELICA DAHURICA ROOT EXTRACT
C3256827|T109|1306164|RXNORM|CARAPA GUIANENSIS SEED OIL|CARAPA GUIANENSIS SEED OIL
C2938850|T121|1306165|RXNORM|ALTHAEA OFFICINALIS ROOT EXTRACT|ALTHAEA OFFICINALIS ROOT EXTRACT
C3500510|T121|1314678|RXNORM|COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENATE / POLYSACCHARIDE IRON COMPLEX / PYRIDOXINE / RIBOFLAVIN / SODIUM ASCORBATE / THIAMINE / VITAMIN B 12 / ZINC SULFATE|COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENATE / POLYSACCHARIDE IRON COMPLEX / PYRIDOXINE / RIBOFLAVIN / SODIUM ASCORBATE / THIAMINE / VITAMIN B 12 / ZINC SULFATE
C3695933|T121|1485045|RXNORM|HYDROXYPROPYL CELLULOSE (TYPE J)|HYDROXYPROPYL CELLULOSE (TYPE J)
C1442898|T129|465062|RXNORM|TRICHOPHYTON MENTAGROPHYTES ANTIGEN|TRICHOPHYTON MENTAGROPHYTES ANTIGEN
C0060132|T121|24809|RXNORM|FEBUPROL|FEBUPROL
C1337387|T129|408134|RXNORM|BOTULISM ANTITOXIN TRIV A,B&E|BOTULISM ANTITOXIN TRIV A,B&E
C0056593|T197|21833|RXNORM|CUPRIC CHLORIDE|CUPRIC CHLORIDE
C0060130|T121|24807|RXNORM|FEBARBAMATE|FEBARBAMATE
C0066274|T130|1551460|RXNORM|METHYL ORANGE|METHYL ORANGE
C0056598|T197|21837|RXNORM|CUPRIC OXIDE|CUPRIC OXIDE
C0981868|T129|852355|RXNORM|FREMONT COTTONWOOD POLLEN EXTRACT|POPULUS FREMONTII POLLEN EXTRACT
C2939943|T130|1014340|RXNORM|ITALIAN RYE GRASS POLLEN EXTRACT|LOLIUM PERENNE SSP. MULTIFLORUM POLLEN EXTRACT
C0953467|T121|291204|RXNORM|TACALCITOL|TACALCITOL
C2701534|T129|852359|RXNORM|PALO VERDE POLLEN EXTRACT|PARKINSONIA FLORIDA POLLEN EXTRACT
C1176329|T121|358274|RXNORM|AMBRISENTAN|AMBRISENTAN
C0892648|T196|1546395|RXNORM|MOLYBDATE ION|MOLYBDATE ION
C1875038|T121|690855|RXNORM|DISOFENIN / STANNOUS CHLORIDE|DISOFENIN / STANNOUS CHLORIDE
C3528961|T109|1363831|RXNORM|PISTACIA LENTISCUS SEED OIL|PISTACIA LENTISCUS SEED OIL
C3530901|T121|1365709|RXNORM|ASARUM HETEROTROPOIDES VAR. MANDSHURICUM ROOT EXTRACT|ASARUM HETEROTROPOIDES VAR. MANDSHURICUM ROOT EXTRACT
C0008929|T121|2578|RXNORM|CLEMASTINE|CLEMASTINE
C0212021|T121|68730|RXNORM|MILBEMYCIN OXIME|MILBEMYCIN OXIME
C2348018|T109|1335893|RXNORM|CURCUMA ZEDORIA ROOT EXTRACT|CURCUMA ZEDORIA ROOT EXTRACT
C0596235|T196|1316581|RXNORM|CALCIUM ION|CA 2+
C0033059|T121|8674|RXNORM|PRENYLAMINE|PRENYLAMINE
C0043572|T121|11454|RXNORM|GLUCOMANNAN|GLUCOMANNAN
C1337158|T121|407906|RXNORM|CHROMIUM CITRATE|CHROMIUM CITRATE
C0303029|T196|1546394|RXNORM|IODINE I-131|IODINE I-131
C0770546|T123|235473|RXNORM|HEPARIN, PORCINE|HEPARIN, PORCINE
C3496118|T121|1368706|RXNORM|STEARATE|STEARATE
C2961510|T121|1053102|RXNORM|ASPIRIN / DEXTROMETHORPHAN / PHENYLEPHRINE|ASPIRIN / DEXTROMETHORPHAN / PHENYLEPHRINE
C0937891|T121|1368704|RXNORM|MICROCRYSTALLINE WAX|MICROCRYSTALLINE WAX
C0077100|T109|1368702|RXNORM|TRIETHYLENE GLYCOL|TRIETHYLENE GLYCOL
C0083072|T109|1368703|RXNORM|ISOPENTANE|ISOPENTANE
C0058460|T197|1368701|RXNORM|DISILVER OXIDE|DISILVER OXIDE
C0018318|T121|5036|RXNORM|GUANETHIDINE|GUANETHIDINE
C1615664|T121|578315|RXNORM|HOODIA GORDONII EXTRACT|HOODIA GORDONII EXTRACT
C0018305|T121|5032|RXNORM|GUAIFENESIN|GUAIFENESIN
C0018312|T121|5033|RXNORM|GUANABENZ|GUANABENZ
C3255957|T121|1368708|RXNORM|MARITIME PINE EXTRACT|MARITIME PINE EXTRACT
C0018304|T121|5031|RXNORM|GUAIACOL|GUAIACOL
C0050940|T121|17128|RXNORM|LANSOPRAZOLE|LANSOPRAZOLE
C0050940|T121|17128|RXNORM|LANSOPRAZOLE|LANSOPRAZOLE
C0050940|T121|17128|RXNORM|LANSOPRAZOLE|LANSOPRAZOLE
C1166176|T121|350465|RXNORM|1-ALPHA-VITAMIN D|1-ALPHA-VITAMIN D
C1445198|T129|894783|RXNORM|GOOSE FEATHER EXTRACT|ANSER ANSER FEATHER EXTRACT
C3818768|T109|1492339|RXNORM|POLYGONUM CUSPIDATUM LEAF EXTRACT|POLYGONUM CUSPIDATUM LEAF EXTRACT
C3818769|T121|1492338|RXNORM|GLYCERETH-6|GLYCERETH-6
C0003371|T129|973|RXNORM|ANTILYMPHOCYTE IMMUNOGLOBULIN|ANTILYMPHOCYTE IMMUNOGLOBULIN
C0000956|T121|154|RXNORM|9-OCTADECENYL ACETATE, (9Z)-|ACENOCOUMAROL
C0002333|T121|596|RXNORM|ALPRAZOLAM|ALPRAZOLAM
C1875133|T121|692988|RXNORM|ESTRONE / TESTOSTERONE|ESTRONE / TESTOSTERONE
C0770121|T121|235219|RXNORM|DIGITALIS LEAF EXTRACT|DIGITALIS LEAVES
C3651718|T122|1430440|RXNORM|PEG-80 SORBITAN PALMITATE|PEG-80 SORBITAN PALMITATE
C2194287|T121|822959|RXNORM|BROMHEXINE / FENOTEROL|BROMHEXINE / FENOTEROL
C1516487|T121|494309|RXNORM|ACETAMINOPHEN / CHLORZOXAZONE|ACETAMINOPHEN / CHLORZOXAZONE
C3531630|T121|1367391|RXNORM|RHAMNUS CATHARTICA FRUIT EXTRACT|RHAMNUS CATHARTICA FRUIT EXTRACT
C0646029|T197|1423457|RXNORM|ALUMINUM HYDROXYPHOSPHATE|ALUMINUM HYDROXYPHOSPHATE
C0939798|T121|1367399|RXNORM|SYMPHYTUM UPLANDICUM LEAF EXTRACT|SYMPHYTUM UPLANDICUM LEAF EXTRACT
C0055936|T125|21285|RXNORM|CLOPREDNOL|CLOPREDNOL
C0178695|T121|62372|RXNORM|HYALURONATE|HYALURONATE
C0178695|T121|62372|RXNORM|HYALURONATE|HYALURONATE
C0178695|T121|62372|RXNORM|HYALURONATE|HYALURONATE
C0350881|T121|102792|RXNORM|CALCIUM SULFALOXATE|CALCIUM SULFALOXATE
C0071099|T121|33740|RXNORM|PIPAZETHATE|PIPAZETATE
C0031237|T129|8080|RXNORM|PERTUSSIS VACCINE|PERTUSSIS VACCINE
C0873038|T121|485858|RXNORM|BOSWELLIA PREPARATION|BOSWELLIA PREPARATION
C3714522|T121|1535478|RXNORM|EQUISETUM ARVENSE WHOLE EXTRACT|EQUISETUM ARVENSE WHOLE EXTRACT
C3818716|T121|1535479|RXNORM|EUCOMMIA ULMOIDES WHOLE EXTRACT|EUCOMMIA ULMOIDES WHOLE EXTRACT
C0672188|T130|194098|RXNORM|S-BENZOYLMERCAPTOACETYLTRIGLYCINE|S-BENZOYLMERCAPTOACETYLTRIGLYCINE
C2241979|T129|762595|RXNORM|TYPHOID VACCINE LIVE TY21A|SALMONELLA TYPHI TY21A LIVE ANTIGEN
C0387288|T121|118886|RXNORM|VERTEPORFIN|VERTEPORFIN
C3818720|T121|1535473|RXNORM|AMOMUM VILLOSUM VAR. XANTHIOIDES WHOLE EXTRACT|AMOMUM VILLOSUM VAR. XANTHIOIDES WHOLE EXTRACT
C3818719|T121|1535474|RXNORM|BROUSSONETIA KAZINOKI WHOLE EXTRACT|BROUSSONETIA KAZINOKI WHOLE EXTRACT
C3818718|T121|1535475|RXNORM|BROUSSONETIA PAPYRIFERA WHOLE EXTRACT|BROUSSONETIA PAPYRIFERA WHOLE EXTRACT
C0536004|T121|139233|RXNORM|MAGNESIUM OROTATE|MAGNESIUM OROTATE
C2930049|T121|1009156|RXNORM|CHLORPHENIRAMINE / METHSCOPOLAMINE / PHENYLEPHRINE|CHLORPHENIRAMINE / METHSCOPOLAMINE / PHENYLEPHRINE
C2930049|T121|1009156|RXNORM|CHLORPHENIRAMINE / METHSCOPOLAMINE / PHENYLEPHRINE|CHLORPHENIRAMINE / METHSCOPOLAMINE / PHENYLEPHRINE
C2930048|T121|1009155|RXNORM|CHYMOTRYPSIN / TRYPSIN|CHYMOTRYPSIN / TRYPSIN
C2930047|T121|1009154|RXNORM|POTASSIUM CITRATE / POTASSIUM GLUCONATE|POTASSIUM CITRATE / POTASSIUM GLUCONATE
C2930046|T121|1009153|RXNORM|POTASSIUM BICARBONATE / POTASSIUM CITRATE|POTASSIUM BICARBONATE / POTASSIUM CITRATE
C2930045|T121|1009152|RXNORM|POTASSIUM CHLORIDE / POTASSIUM GLUCONATE|POTASSIUM CHLORIDE / POTASSIUM GLUCONATE
C2930044|T121|1009151|RXNORM|CORTICOTROPIN / ZINC HYDROXIDE|CORTICOTROPIN / ZINC HYDROXIDE
C1099456|T121|321988|RXNORM|ESCITALOPRAM|ESCITALOPRAM
C0991832|T125|317235|RXNORM|NPH INSULIN, BEEF|INSULIN BEEF, ISOPHANE
C0164613|T129|59744|RXNORM|INTERFERON ALFACON-1|INTERFERON ALFACON-1
C0063908|T130|27863|RXNORM|ISO-SULFAN BLUE|ISO-SULFAN BLUE
C2928041|T121|1007119|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE|ACETAMINOPHEN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE
C2928040|T121|1007118|RXNORM|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE / PYRILAMINE|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE / PYRILAMINE
C0072858|T121|1546359|RXNORM|QUINAPRILAT|QUINAPRILAT
C0164608|T121|59743|RXNORM|QUINETHAZONE|QUINETHAZONE
C2928037|T121|1007115|RXNORM|POLYMYXIN B / TRIAMCINOLONE|POLYMYXIN B / TRIAMCINOLONE
C2928036|T121|1007114|RXNORM|CYNARA PREPARATION / DEHYDROCHOLATE|CYNARA PREPARATION / DEHYDROCHOLATE
C2928039|T121|1007117|RXNORM|CHLORPHENIRAMINE / PHENYLTOLOXAMINE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / PHENYLTOLOXAMINE / PSEUDOEPHEDRINE
C2928038|T121|1007116|RXNORM|FLUOROMETHOLONE / TETRAHYDROZOLINE|FLUOROMETHOLONE / TETRAHYDROZOLINE
C2826087|T121|1546353|RXNORM|2-ETHYLHEXYL 4-PHENYLBENZOPHENONE-2'-CARBOXYLATE|2-ETHYLHEXYL 4-PHENYLBENZOPHENONE-2'-CARBOXYLATE
C2928032|T121|1007110|RXNORM|BROMHEXINE / PENICILLIN V|BROMHEXINE / PENICILLIN V
C2928035|T121|1007113|RXNORM|ALLOIN / PHENOLPHTHALEIN|ALLOIN / PHENOLPHTHALEIN
C2928034|T121|1007112|RXNORM|ASPIRIN / PYRIDINOLCARBAMATE|ASPIRIN / PYRIDINOLCARBAMATE
C1875664|T121|689944|RXNORM|PETROLEUM DISTILLATE / PIPERONYL BUTOXIDE / PYRETHRINS|PETROLEUM DISTILLATE / PIPERONYL BUTOXIDE / PYRETHRINS
C0991843|T109|1309249|RXNORM|LANOLIN OIL|LANOLIN OIL
C0039865|T121|10471|RXNORM|THIETHYLPERAZINE|THIETHYLPERAZINE
C2073839|T121|816818|RXNORM|ASPIRIN / CHLORPHENIRAMINE|ASPIRIN / CHLORPHENIRAMINE
C0039871|T131|10473|RXNORM|THIOTEPA|THIOTEPA
C0039867|T121|10472|RXNORM|THIMEROSAL|THIMEROSAL
C3488334|T129|1309242|RXNORM|SOLIDAGO VIRGAUREA POLLEN EXTRACT|SOLIDAGO VIRGAUREA POLLEN EXTRACT
C0010198|T168|1309243|RXNORM|COTTONSEED OIL|COTTONSEED OIL
C0632804|T109|1309240|RXNORM|JASMINE OIL|JASMINE OIL
C0304103|T109|1309241|RXNORM|CORIANDER OIL|CORIANDER OIL
C1509729|T109|1309246|RXNORM|POLYOXYL 35 CASTOR OIL|POLYOXYL 35 CASTOR OIL
C0036845|T168|1309247|RXNORM|SESAME OIL|SESAME OIL
C0758616|T109|1309245|RXNORM|JUNIPER BERRY OIL|JUNIPER BERRY OIL
C3645243|T121|1427026|RXNORM|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-BRISBANE-60-2008-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-BRISBANE-60-2008-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS
C3645239|T129|1427022|RXNORM|INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS|INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS
C3645237|T129|1427020|RXNORM|INFLUENZA B VIRUS VACCINE, B-BRISBANE-60-2008-LIKE VIRUS|INFLUENZA B VIRUS VACCINE, B-BRISBANE-60-2008-LIKE VIRUS
C1873633|T121|700810|RXNORM|LISDEXAMFETAMINE|LISDEXAMFETAMINE
C2193931|T121|820748|RXNORM|DIPHENHYDRAMINE / NAPHAZOLINE|DIPHENHYDRAMINE / NAPHAZOLINE
C1445387|T121|1428417|RXNORM|CYNODON DACTYLON EXTRACT|CYNODON DACTYLON EXTRACT
C0065656|T121|29275|RXNORM|MANIDIPINE|MANIDIPINE
C3848536|T121|1546402|RXNORM|SULFONATED OLEIC ACID|SULFONATED OLEIC ACID
C0071103|T121|33743|RXNORM|PIPENZOLATE|PIPENZOLATE
C0064226|T123|28116|RXNORM|KAMALA EXTRACT|KAMALA EXTRACT
C0149368|T121|58295|RXNORM|ZINC ACETATE|ZINC ACETATE
C0149368|T121|58295|RXNORM|ZINC ACETATE|ZINC ACETATE
C0071129|T121|33767|RXNORM|PIRBUTEROL|PIRBUTEROL
C0071126|T195|33764|RXNORM|PIRARUBICIN|PIRARUBICIN
C0772046|T197|236741|RXNORM|MAGNESIUM SULFATE HEPTAHYDRATE|MAGNESIUM SULFATE HEPTAHYDRATE
C0070426|T121|1546400|RXNORM|PERINDOPRILAT|PERINDOPRILAT
C0033979|T123|8928|RXNORM|PSYLLIUM|PSYLLIUM
C2928724|T121|1007809|RXNORM|MAGNESIUM SULFATE / POTASSIUM SULFATE / SODIUM SULFATE|MAGNESIUM SULFATE / POTASSIUM SULFATE / SODIUM SULFATE
C2928723|T121|1007808|RXNORM|IVERMECTIN / PYRANTEL|IVERMECTIN / PYRANTEL
C2586798|T129|830457|RXNORM|RABIES VIRUS VACCINE FLURY-LEP STRAIN|RABIES VIRUS VACCINE FLURY-LEP STRAIN
C2928718|T121|1007803|RXNORM|METHENAMINE / SALICYLIC ACID|METHENAMINE / SALICYLIC ACID
C2928718|T121|1007803|RXNORM|METHENAMINE / SALICYLIC ACID|METHENAMINE / SALICYLIC ACID
C2928717|T121|1007802|RXNORM|DEXTRAN 70 / GLYCERIN / HYPROMELLOSE|DEXTRAN 70 / GLYCERIN / HYPROMELLOSE
C2928716|T121|1007801|RXNORM|BILBERRY EXTRACT / BLACK PEPPER PREPARATION|BILBERRY EXTRACT / BLACK PEPPER PREPARATION
C2928715|T121|1007800|RXNORM|BUTABARBITAL / HOMATROPINE|BUTABARBITAL / HOMATROPINE
C2928722|T121|1007807|RXNORM|ASCORBIC ACID / FOLIC ACID / IRON CARBONYL / VITAMIN B 12|ASCORBIC ACID / FOLIC ACID / IRON CARBONYL / VITAMIN B 12
C2928721|T121|1007806|RXNORM|GUAIACOLSULFONIC ACID / PHENYLEPHRINE / PROMETHAZINE|GUAIACOLSULFONIC ACID / PHENYLEPHRINE / PROMETHAZINE
C2928720|T121|1007805|RXNORM|MINERAL OIL / PRAMOXINE / ZINC OXIDE|MINERAL OIL / PRAMOXINE / ZINC OXIDE
C0298067|T121|1592254|RXNORM|PIRFENIDONE|PIRFENIDONE
C0370067|T121|113931|RXNORM|CLAVULANATE / TICARCILLIN|CLAVULANATE / TICARCILLIN
C0049477|T121|15978|RXNORM|ACEXAMIC ACID|ACEXAMIC ACID
C0068673|T121|31722|RXNORM|NIAPRAZINE|NIAPRAZINE
C2726176|T129|1010879|RXNORM|BAY LEAF ALLERGENIC EXTRACT|LAURUS NOBILIS ALLERGENIC EXTRACT
C3256707|T109|1314208|RXNORM|OCTYLDODECYL STEARATE|OCTYLDODECYL STEARATE
C3486690|T121|1309992|RXNORM|FUMARIA OFFICINALIS FLOWERING TOP EXTRACT|FUMARIA OFFICINALIS FLOWERING TOP EXTRACT
C0052993|T197|18789|RXNORM|BASIC ALUMINUM CARBONATE GEL|BASIC ALUMINUM CARBONATE GEL
C0590796|T121|151221|RXNORM|CYCLOPENTHIAZIDE / OXPRENOLOL|CYCLOPENTHIAZIDE / OXPRENOLOL
C3256339|T109|1305639|RXNORM|AMYRIS BALSAMIFERA OIL|AMYRIS BALSAMIFERA OIL
C0102271|T168|1305638|RXNORM|ALMOND OIL|ALMOND OIL
C3256062|T168|1305636|RXNORM|MENTHA ARVENSIS FLOWER OIL|MENTHA ARVENSIS FLOWER OIL
C1635037|T121|607999|RXNORM|METFORMIN / PIOGLITAZONE|METFORMIN / PIOGLITAZONE
C1721512|T109|1305634|RXNORM|CINNAMON OIL, BARK|CINNAMON OIL, BARK
C3255743|T109|1305633|RXNORM|CHAMAECYPARIS OBTUSA WOOD OIL|CHAMAECYPARIS OBTUSA WOOD OIL
C3256627|T121|1314205|RXNORM|POLYGLYCERIN-10|POLYGLYCERIN-10
C3474157|T168|1305631|RXNORM|CAMELINA SATIVA SEED OIL|CAMELINA SATIVA SEED OIL
C2927366|T129|1005909|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-CALIFORNIA-7-2009 (H1N1) STRAIN|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-CALIFORNIA-7-2009 (H1N1) STRAIN
C3651785|T121|1428414|RXNORM|AGROSTEMMA GITHAGO SEED EXTRACT|AGROSTEMMA GITHAGO SEED EXTRACT
C0648444|T121|1491978|RXNORM|BORNYL ACETATE|BORNYL ACETATE
C1881356|T196|1546443|RXNORM|LANTHANUM CATION (3+)|LANTHANUM CATION (3+)
C0359084|T121|107013|RXNORM|NEOMYCIN / TRIAMCINOLONE|NEOMYCIN / TRIAMCINOLONE
C0359083|T121|107012|RXNORM|ECONAZOLE / TRIAMCINOLONE|ECONAZOLE / TRIAMCINOLONE
C0359082|T121|107011|RXNORM|NYSTATIN / TRIAMCINOLONE|NYSTATIN / TRIAMCINOLONE
C0359081|T121|107010|RXNORM|CHLORTETRACYCLINE / TRIAMCINOLONE|CHLORTETRACYCLINE / TRIAMCINOLONE
C2142857|T121|814483|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / CODEINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / CHLORPHENIRAMINE / CODEINE / PSEUDOEPHEDRINE
C2722033|T129|867202|RXNORM|CLADOSPORIUM SPHAEROSPERMUM ALLERGENIC EXTRACT|CLADOSPORIUM SPHAEROSPERMUM ALLERGENIC EXTRACT
C3191261|T121|1145801|RXNORM|EMTRICITABINE / RILPIVIRINE / TENOFOVIR DISOPROXIL|EMTRICITABINE / RILPIVIRINE / TENOFOVIR DISOPROXIL
C1874520|T121|690269|RXNORM|BENZOCAINE / LICORICE / MENTHOL|BENZOCAINE / LICORICE / MENTHOL
C3282452|T121|1352501|RXNORM|EVERNIA PRUNASTRI EXTRACT|EVERNIA PRUNASTRI EXTRACT
C2701564|T129|852398|RXNORM|COCHLIOBOLUS SATIVUS EXTRACT|COCHLIOBOLUS SATIVUS EXTRACT
C2929352|T121|1008448|RXNORM|MAGNESIUM GLUCONATE / MAGNESIUM OXIDE|MAGNESIUM GLUCONATE / MAGNESIUM OXIDE
C2929353|T121|1008449|RXNORM|CALCIUM CHLORIDE, DIHYDRATION / LACTATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CHLORIDE, DIHYDRATION / LACTATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C2929350|T121|1008446|RXNORM|MAGNESIUM OXIDE / SODIUM BICARBONATE|MAGNESIUM OXIDE / SODIUM BICARBONATE
C2929351|T121|1008447|RXNORM|DAPSONE / FERROUS OXALATE|DAPSONE / FERROUS OXALATE
C2929348|T121|1008444|RXNORM|ESTRADIOL / FLUPREDNIDENE|ESTRADIOL / FLUPREDNIDENE
C2929349|T121|1008445|RXNORM|ALUMINUM HYDROXIDE / THEOPHYLLINE|ALUMINUM HYDROXIDE / THEOPHYLLINE
C2929346|T121|1008442|RXNORM|BISMUTH SUBGALLATE / MEPENZOLATE / PHTHALYLSULFATHIAZOLE|BISMUTH SUBGALLATE / MEPENZOLATE / PHTHALYLSULFATHIAZOLE
C2928313|T121|1007391|RXNORM|BISMUTH SUBGALLATE / HYDROCORTISONE|BISMUTH SUBGALLATE / HYDROCORTISONE
C2929344|T121|1008440|RXNORM|IBUPROFEN / SCOPOLAMINE|IBUPROFEN / SCOPOLAMINE
C2929345|T121|1008441|RXNORM|ORPHENADRINE / PROPYPHENAZONE|ORPHENADRINE / PROPYPHENAZONE
C3848520|T196|1546442|RXNORM|IODATE ION|IODATE ION
C2928319|T121|1007397|RXNORM|GLUCOSAMINE HYDROCHLORIDE / GLUCOSAMINE SULFATE|GLUCOSAMINE HYDROCHLORIDE / GLUCOSAMINE SULFATE
C1874011|T121|690205|RXNORM|ACETIC ACID / SALICYLIC ACID|ACETIC ACID / SALICYLIC ACID
C3247243|T129|1191668|RXNORM|GONADOTROPIN RELEASING FACTOR ANALOG-DIPHTHERIA TOXOID CONJUGATE|GONADOTROPIN RELEASING FACTOR ANALOG-DIPHTHERIA TOXOID CONJUGATE
C1874008|T121|690201|RXNORM|ACETIC ACID / DESONIDE|ACETIC ACID / DESONIDE
C2928318|T121|1007396|RXNORM|COLLOIDAL OATMEAL / SALICYLIC ACID|COLLOIDAL OATMEAL / SALICYLIC ACID
C1165938|T121|350262|RXNORM|CINCHONA OFFICINALIS PREPARATION|CINCHONA OFFICINALIS PREPARATION
C0771999|T197|1433888|RXNORM|GOLD TRIBROMIDE|GOLD TRIBROMIDE
C3663845|T122|1433886|RXNORM|HYDROXYPROPYL CELLULOSE (TYPE M)|HYDROXYPROPYL CELLULOSE (TYPE M)
C2928316|T121|1007394|RXNORM|METHYLPARABEN / PROPYLPARABEN|METHYLPARABEN / PROPYLPARABEN
C2194159|T121|813961|RXNORM|ASCORBIC ACID / ASPIRIN|ASCORBIC ACID / ASPIRIN
C0994438|T121|317825|RXNORM|HORSE CHESTNUT PREPARATION|HORSE CHESTNUT PREPARATION
C0994437|T109|317824|RXNORM|CEPHAELIS IPECACUANHA PREPARATION|CEPHAELIS IPECACUANHA PREPARATION
C2928321|T121|1007399|RXNORM|AMYLASES / LIPASE|AMYLASES / LIPASE
C0301370|T121|89781|RXNORM|BELLADONNA EXTRACT, USP|ATROPA BELLADONA EXTRACT
C0301369|T121|89780|RXNORM|ANISOTROPINE|ANISOTROPINE
C0301371|T121|89782|RXNORM|DIPHEMANIL|DIPHEMANIL
C0301374|T121|89785|RXNORM|METHSCOPOLAMINE|METHYLSCOPOLAMINE
C0301373|T121|89784|RXNORM|ISOPROPAMIDE|ISOPROPAMIDE
C0005070|T121|1406|RXNORM|BENZOIN|BENZOIN RESIN
C0246415|T121|72962|RXNORM|DOCETAXEL|DOCETAXEL
C2702357|T129|892543|RXNORM|CODFISH ALLERGENIC EXTRACT|CODFISH ALLERGENIC EXTRACT
C0246421|T121|72965|RXNORM|LETROZOLE|LETROZOLE
C1095785|T007|487252|RXNORM|SPIRULINA|SPIRULINA
C0305055|T129|91601|RXNORM|LYMPHOCYTE IMMUNE GLOBULIN|LYMPHOCYTE IMMUNE GLOBULIN
C0305058|T129|91603|RXNORM|TETANUS IMMUNE GLOBULIN, HUMAN|TETANUS IMMUNE GLOBULIN, HUMAN
C0305057|T129|91602|RXNORM|EQUINE DIPHTHERIA ANTITOXIN|EQUINE DIPHTHERIA ANTITOXIN
C3555483|T109|1376500|RXNORM|PANAX PSEUDOGINSENG ROOT EXTRACT|PANAX PSEUDOGINSENG ROOT EXTRACT
C0073047|T121|35350|RXNORM|REMOXIPRIDE|REMOXIPRIDE
C2701305|T129|852102|RXNORM|PULLULARIA EXTRACT|AUREOBASIDIUM PULLULANS VAR. PULLUTANS EXTRACT
C3282853|T121|1313260|RXNORM|OCTYLDODECYL LACTATE|OCTYLDODECYL LACTATE
C0068986|T121|31988|RXNORM|NORFENEFRINE|NORFENEFRINE
C2701309|T129|852106|RXNORM|ALKALI BLITE POLLEN EXTRACT|SUAEDA NIGRA POLLEN EXTRACT
C0042674|T121|11201|RXNORM|VINCAMINE|VINCAMINE
C0042679|T121|11202|RXNORM|VINCRISTINE|VINCRISTINE
C2928970|T121|1008059|RXNORM|BROMPHENIRAMINE / CODEINE / GUAIFENESIN|BROMPHENIRAMINE / CODEINE / GUAIFENESIN
C2928969|T121|1008058|RXNORM|BUTAFOSFAN / VITAMIN B 12|BUTAFOSFAN / VITAMIN B 12
C2928966|T121|1008055|RXNORM|PREDNISOLONE / TRIMEPRAZINE|PREDNISOLONE / TRIMEPRAZINE
C2928965|T121|1008054|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007, IVR-148 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-URUGUAY-716-2007, NYMC X-175C (H3N2) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007, IVR-148 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-URUGUAY-716-2007, NYMC X-175C (H3N2) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN
C2928968|T121|1008057|RXNORM|FRUCTOSE / GLUCOSE / SODIUM CITRATE|FRUCTOSE / GLUCOSE / SODIUM CITRATE
C2928967|T121|1008056|RXNORM|CALCIUM CARBONATE / MAGNESIUM OXIDE / VALERIAN ROOT EXTRACT / VALINE|CALCIUM CARBONATE / MAGNESIUM OXIDE / VALERIAN ROOT EXTRACT / VALINE
C2928962|T121|1008051|RXNORM|CAFFEINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN B6|CAFFEINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN B6
C2928961|T121|1008050|RXNORM|MENTHOL / METHYL SALICYLATE / TOURMALINE|MENTHOL / METHYL SALICYLATE / TOURMALINE
C2928964|T121|1008053|RXNORM|CHLOROXYLENOL / COPPER SULFATE|CHLOROXYLENOL / COPPER SULFATE
C2928963|T121|1008052|RXNORM|AMYLOCAINE / TRICHLOROACETALDEHYDE|AMYLOCAINE / TRICHLOROACETALDEHYDE
C3667870|T109|1440231|RXNORM|MYRISTAMIDOPROPYL PG-DIMONIUM CHLORIDE PHOSPHATE|MYRISTAMIDOPROPYL PG-DIMONIUM CHLORIDE PHOSPHATE
C0070139|T130|32950|RXNORM|PATENT BLUE VIOLET|PATENT BLUE VIOLET
C2701442|T129|852244|RXNORM|CANIS LUPUS FAMILIARIS EXTRACT|CANIS LUPUS FAMILIARIS EXTRACT
C3667872|T109|1440235|RXNORM|PEG-8 GLYCERYL ISOSTEARATE|PEG-8 GLYCERYL ISOSTEARATE
C2741441|T129|901199|RXNORM|SESAME SEED ALLERGENIC EXTRACT|SESAMUM INDICUM SEED ALLERGENIC EXTRACT
C3667873|T109|1440237|RXNORM|PEG-80 SORBITAN LAURATE|PEG-80 SORBITAN LAURATE
C0053323|T121|19075|RXNORM|BENZYLPARABEN|BENZYLPARABEN
C3667874|T121|1440239|RXNORM|PPG-12-SMDI COPOLYMER|PPG-12-SMDI COPOLYMER
C0163641|T121|1116238|RXNORM|TOLU BALSAM|TOLU BALSAM
C0053327|T195|19079|RXNORM|BENZYLPENICILLOYL POLYLYSINE|BENZYLPENICILLOYL POLYLYSINE
C2604635|T121|1367839|RXNORM|MIPOMERSEN|MIPOMERSEN
C3486808|T121|1351787|RXNORM|SCHOENOCAULON OFFICINALE SEED EXTRACT|SCHOENOCAULON OFFICINALE SEED EXTRACT
C0254824|T121|76273|RXNORM|PROPINOX|PROPINOX
C0297269|T121|87866|RXNORM|ARDEPARIN|ARDEPARIN
C3255682|T109|1426383|RXNORM|HIMANTHALIA ELONGATA EXTRACT|HIMANTHALIA ELONGATA EXTRACT
C0600615|T130|155156|RXNORM|POLOXAMER|POLOXAMER
C0600611|T121|155152|RXNORM|POLOXAMER 188|POLOXAMER 188
C3484911|T129|1303855|RXNORM|INFLUENZA B VIRUS VACCINE, B-WISCONSIN-1-2010-LIKE VIRUS|INFLUENZA B VIRUS VACCINE, B-WISCONSIN-1-2010-LIKE VIRUS
C3256591|T109|1309401|RXNORM|AFRAMOMUM ANGUSTIFOLIUM SEED EXTRACT|AFRAMOMUM ANGUSTIFOLIUM SEED EXTRACT
C3256411|T109|1309403|RXNORM|ANOGEISSUS LEIOCARPUS BARK EXTRACT|ANOGEISSUS LEIOCARPUS BARK EXTRACT
C3484909|T129|1303851|RXNORM|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS
C2929913|T121|1009018|RXNORM|AMPRENAVIR / VITAMIN E|AMPRENAVIR / VITAMIN E
C3256494|T109|1309406|RXNORM|ACER SACCHARUM BARK-SAP EXTRACT|ACER SACCHARUM BARK-SAP EXTRACT
C3256018|T109|1309407|RXNORM|BETULA PLATYPHYLLA VAR. JAPONICA BARK EXTRACT|BETULA PLATYPHYLLA VAR. JAPONICA BARK EXTRACT
C2193908|T121|817139|RXNORM|FENOFIBRATE / PANTETHINE|FENOFIBRATE / PANTETHINE
C3644976|T130|1426161|RXNORM|PIGMENT RED 48|PIGMENT RED 48
C3644975|T122|1426160|RXNORM|PEG-175 DIISOSTEARATE|PEG-175 DIISOSTEARATE
C3644978|T109|1426163|RXNORM|ETHYL LAUROYL ARGINATE|ETHYL LAUROYL ARGINATE
C2929911|T121|1009016|RXNORM|HOPS EXTRACT / VALERIAN ROOT EXTRACT|HOPS EXTRACT / VALERIAN ROOT EXTRACT
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, BEECH|PRASTERONE
C0058415|T121|23410|RXNORM|DIPIVEFRIN|DIPIVEFRINE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, BEE|PRASTERONE
C0003438|T121|1009|RXNORM|GLUCOSE / MILRINONE|ANTITHROMBIN III
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, BIRCH|PRASTERONE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, BERMUDA GRASS|PRASTERONE
C0058425|T121|23419|RXNORM|DIPROPIZINE|DROPROPIZINE
C2929909|T121|1009014|RXNORM|2-PHENYLPHENOL / CHLOROCRESOL / CLOROPHENE|2-PHENYLPHENOL / CHLOROCRESOL / CLOROPHENE
C0025942|T121|6932|RXNORM|MICONAZOLE|MICONAZOLE
C0025942|T121|6932|RXNORM|MICONAZOLE|MICONAZOLE
C0025942|T121|6932|RXNORM|MICONAZOLE|MICONAZOLE
C0025942|T121|6932|RXNORM|MICONAZOLE|MICONAZOLE
C0025942|T121|6932|RXNORM|MICONAZOLE|MICONAZOLE
C2721771|T121|877015|RXNORM|LEVOLEUCOVORIN|LEVOLEUCOVORIN
C2927826|T121|1006902|RXNORM|BETAINE / GLUTAMATE / PEPSIN A|BETAINE / GLUTAMATE / PEPSIN A
C1257880|T121|382272|RXNORM|LINOLEIC ACIDS, CONJUGATED|LINOLEIC ACIDS, CONJUGATED
C2927829|T121|1006905|RXNORM|CARBETAPENTANE / GUAIACOLSULFONATE / PHENYLEPHRINE|CARBETAPENTANE / GUAIACOLSULFONATE / PHENYLEPHRINE
C1170011|T125|352385|RXNORM|INSULIN, ASPART PROTAMINE, HUMAN|INSULIN, ASPART PROTAMINE, HUMAN
C3833355|T109|1541236|RXNORM|C12-17 ALKANE|C12-17 ALKANE
C2929908|T121|1009013|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE / PYRILAMINE|DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE / PYRILAMINE
C0994408|T121|317808|RXNORM|ELDER EXTRACT|ELDER EXTRACT
C2929905|T121|1009010|RXNORM|PREDNISOLONE / SALICYLIC ACID|PREDNISOLONE / SALICYLIC ACID
C0718057|T121|214829|RXNORM|SODIUM BICARBONATE / SODIUM CITRATE|SODIUM BICARBONATE / SODIUM CITRATE
C2929906|T121|1009011|RXNORM|CALCIUM PHOSPHATE / DEHYDROEPIANDROSTERONE|CALCIUM PHOSPHATE / PRASTERONE
C0298130|T121|88249|RXNORM|MONTELUKAST|MONTELUKAST
C2242160|T129|763100|RXNORM|POLIOVIRUS VACCINE INACTIVATED, TYPE 3 (SAUKETT)|POLIOVIRUS VACCINE INACTIVATED, TYPE 3 (SAUKETT)
C3860108|T121|1594579|RXNORM|CLEMATIS HEXAPETALA WHOLE EXTRACT|CLEMATIS HEXAPETALA WHOLE EXTRACT
C2746955|T129|904498|RXNORM|CAROB ALLERGENIC EXTRACT|CERATONIA SILIQUA ALLERGENIC EXTRACT
C0937649|T121|283587|RXNORM|YUCCA ROOT|YUCCA ROOT
C0007955|T196|2296|RXNORM|CHARCOAL|CHARCOAL
C0057950|T109|1538383|RXNORM|DIETHYLENE GLYCOL MONOMETHYL ETHER|DIETHYLENE GLYCOL MONOMETHYL ETHER
C2730186|T129|892526|RXNORM|CASHEW NUT ALLERGENIC EXTRACT|ANACARDIUM OCCIDENTALE ALLERGENIC EXTRACT
C1302054|T126|392509|RXNORM|LARONIDASE|LARONIDASE
C1302053|T121|392508|RXNORM|ERYTHROMYCIN / TRETINOIN|ERYTHROMYCIN / TRETINOIN
C3643658|T121|1422085|RXNORM|ATORVASTATIN / EZETIMIBE|ATORVASTATIN / EZETIMIBE
C1412008|T121|453012|RXNORM|PROTAMONE|PROTAMONE
C0282386|T195|82122|RXNORM|LEVOFLOXACIN|LEVOFLOXACIN
C0282386|T195|82122|RXNORM|LEVOFLOXACIN|LEVOFLOXACIN
C1302047|T121|392503|RXNORM|MEQUINOL / TRETINOIN|MEQUINOL / TRETINOIN
C2929647|T121|1008748|RXNORM|HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE / TETANUS TOXOID VACCINE, INACTIVATED|HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE / TETANUS TOXOID VACCINE, INACTIVATED
C1533426|T109|1314848|RXNORM|ISOSTEARYL NEOPENTANOATE|ISOSTEARYL NEOPENTANOATE
C0982317|T109|1314849|RXNORM|PEG-40 STEARATE|PEG-40 STEARATE
C0074536|T197|1314846|RXNORM|SILVER CHLORIDE|SILVER CHLORIDE
C0033148|T121|8691|RXNORM|PRIMIDONE|PRIMIDONE
C3256147|T121|1314844|RXNORM|CORALLINA OFFICINALIS EXTRACT|CORALLINA OFFICINALIS EXTRACT
C0000986|T109|1370450|RXNORM|ACETIC ANHYDRIDE|ACETIC ANHYDRIDE
C3500585|T109|1314842|RXNORM|BEHENETH-20|BEHENETH-20
C0041009|T121|10811|RXNORM|TRIHEXYPHENIDYL|TRIHEXYPHENIDYL
C0085379|T129|42405|RXNORM|MUROMONAB-CD3|MUROMONAB-CD3
C0981943|T129|895919|RXNORM|SPINY PIGWEED POLLEN EXTRACT|AMARANTHUS SPINOSUS POLLEN EXTRACT
C0041345|T121|10917|RXNORM|TUBOCURARINE|TUBOCURARINE
C3538671|T121|1373248|RXNORM|CALAMINE / MENTHOL / ZINC OXIDE|CALAMINE / MENTHOL / ZINC OXIDE
C0031379|T121|8120|RXNORM|PHENAZOPYRIDINE|PHENAZOPYRIDINE
C0045549|T121|1482535|RXNORM|2,5-DIAMINOTOLUENE|2,5-DIAMINOTOLUENE
C0039245|T121|10318|RXNORM|TACRINE|TACRINE
C2929846|T121|1008949|RXNORM|CAFFEINE / PHENOBARBITAL|CAFFEINE / PHENOBARBITAL
C2929845|T121|1008948|RXNORM|SODIUM BICARBONATE / SODIUM FLUORIDE|SODIUM BICARBONATE / SODIUM FLUORIDE
C2929840|T121|1008943|RXNORM|LANOLIN / SILICONES|LANOLIN / SILICONES
C0027603|T195|7299|RXNORM|NEOMYCIN|NEOMYCIN
C0027603|T195|7299|RXNORM|NEOMYCIN|NEOMYCIN
C2929838|T121|1008941|RXNORM|CHOLINE / PROCAINE|CHOLINE / PROCAINE
C2929837|T121|1008940|RXNORM|ASCORBIC ACID / SODIUM FLUORIDE / VITAMIN A / VITAMIN D|ASCORBIC ACID / SODIUM FLUORIDE / VITAMIN A / VITAMIN D
C2929844|T121|1008947|RXNORM|CAFFEINE / DIMENHYDRINATE|CAFFEINE / DIMENHYDRINATE
C2929843|T121|1008946|RXNORM|MURAMIDASE / VITAMIN B6|MURAMIDASE / VITAMIN B6
C2929842|T121|1008945|RXNORM|ETOFENAMATE / NIACIN|ETOFENAMATE / NIACIN
C2929841|T121|1008944|RXNORM|ETHANOL / RESORCINOL / SULFUR|ETHANOL / RESORCINOL / SULFUR
C2929991|T121|1009096|RXNORM|LYCOPENE / VITAMIN E|LYCOPENE / VITAMIN E
C2929992|T121|1009097|RXNORM|ASCORBIC ACID / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D|ASCORBIC ACID / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D
C2929989|T121|1009094|RXNORM|AMILORIDE / FUROSEMIDE / INDAPAMIDE|AMILORIDE / FUROSEMIDE / INDAPAMIDE
C2929990|T121|1009095|RXNORM|BACITRACIN / TIXOCORTOL|BACITRACIN / TIXOCORTOL
C2929987|T121|1009092|RXNORM|ESTRADIOL / TYROTHRICIN|ESTRADIOL / TYROTHRICIN
C2929988|T121|1009093|RXNORM|LIDOCAINE / RUSCOGENIN|LIDOCAINE / RUSCOGENIN
C2929985|T121|1009090|RXNORM|BENZALKONIUM / BENZOCAINE / ZINC CHLORIDE|BENZALKONIUM / BENZOCAINE / ZINC CHLORIDE
C2929986|T121|1009091|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE
C2183097|T121|819146|RXNORM|DEXTROMETHORPHAN / POTASSIUM IODIDE|DEXTROMETHORPHAN / POTASSIUM IODIDE
C2701757|T129|852716|RXNORM|YELLOW PINE POLLEN EXTRACT|PINUS PONDEROSA POLLEN EXTRACT
C3555523|T121|1374402|RXNORM|MANSOA ALLIACEA LEAF EXTRACT|MANSOA ALLIACEA LEAF EXTRACT
C2929993|T121|1009098|RXNORM|BICLOTYMOL / CHLORPHENIRAMINE / PHENYLEPHRINE|BICLOTYMOL / CHLORPHENIRAMINE / PHENYLEPHRINE
C2929994|T121|1009099|RXNORM|ASCORBIC ACID / VITAMIN A|ASCORBIC ACID / VITAMIN A
C1719942|T121|645245|RXNORM|DEXTROMETHORPHAN / TRIPROLIDINE|DEXTROMETHORPHAN / TRIPROLIDINE
C3832921|T130|1539907|RXNORM|D&C RED NO. 6 BARIUM LAKE|D&C RED NO. 6 BARIUM LAKE
C0771503|T121|236249|RXNORM|PARETHOXYCAINE|PARETHOXYCAINE
C0771502|T121|236248|RXNORM|AMYLMETACRESOL|AMYLMETACRESOL
C0937916|T121|283809|RXNORM|TRAVOPROST|TRAVOPROST
C1174893|T121|356887|RXNORM|LEVOCETIRIZINE|LEVOCETIRIZINE
C0937912|T121|283805|RXNORM|BEAN POD EXTRACT|BEAN POD EXTRACT
C2193980|T121|819537|RXNORM|EPHEDRINE / GUAIFENESIN / NOSCAPINE|EPHEDRINE / GUAIFENESIN / NOSCAPINE
C0771815|T121|236531|RXNORM|BUCHU|BUCHU
C1874570|T121|690448|RXNORM|BISACODYL / TANNIC ACID|BISACODYL / TANNIC ACID
C2080637|T121|821472|RXNORM|PHLOROGLUCINOL / TRIMETHOXYBENZENE|PHLOROGLUCINOL / TRIMETHOXYBENZENE
C0216660|T121|69722|RXNORM|ZANAMIVIR|ZANAMIVIR
C2183736|T121|817502|RXNORM|DIPHENHYDRAMINE / RESORCINOL|DIPHENHYDRAMINE / RESORCINOL
C0030040|T121|7801|RXNORM|OXPRENOLOL|OXPRENOLOL
C0392214|T109|121047|RXNORM|PROPIONATE|PROPIONATE
C3256620|T121|1311591|RXNORM|FRITILLARIA PRZEWALSKII BULB EXTRACT|FRITILLARIA PRZEWALSKII BULB EXTRACT
C3695970|T109|1483728|RXNORM|AMODIMETHICONE (3500 CST)|AMODIMETHICONE (3500 CST)
C3695969|T121|1483729|RXNORM|ASPARAGUS ADSCENDENS ROOT EXTRACT|ASPARAGUS ADSCENDENS ROOT EXTRACT
C1268566|T196|1483727|RXNORM|SODIUM NA-22|SODIUM NA-22
C3651947|T122|1431306|RXNORM|TAURATE|TAURATE
C2825462|T121|1025342|RXNORM|LEVOMEFOLIC ACID|LEVOMEFOLIC ACID
C0360192|T121|107784|RXNORM|COLFOSCERIL|COLFOSCERIL
C0105750|T121|46967|RXNORM|BERACTANT|BERACTANT
C0055964|T121|21311|RXNORM|CLOXAZOLAM|CLOXAZOLAM
C2701372|T129|852170|RXNORM|ARROYO WILLOW POLLEN EXTRACT|SALIX LASIOLEPIS POLLEN EXTRACT
C2939991|T121|1014404|RXNORM|ASCORBIC ACID / FOLIC ACID / POLYSACCHARIDE IRON COMPLEX|ASCORBIC ACID / FOLIC ACID / POLYSACCHARIDE IRON COMPLEX
C0012322|T122|3430|RXNORM|DIHYDROXYACETONE|DIHYDROXYACETONE
C0051500|T121|17599|RXNORM|ALTHIAZIDE|ALTHIAZIDE
C0770962|T127|235788|RXNORM|NICOBOXIL|NICOBOXIL
C0003166|T121|873|RXNORM|ANTHRALIN|ANTHRALIN
C3531181|T109|1366231|RXNORM|PEG PPG116-66 COPOLYMER|PEG PPG116-66 COPOLYMER
C0007018|T197|2037|RXNORM|CARBON MONOXIDE|CARBON MONOXIDE
C0770959|T121|235787|RXNORM|CAPSICUM OLEORESIN|CAPSICUM OLEORESIN
C0007012|T197|2034|RXNORM|CARBON DIOXIDE|CARBON DIOXIDE
C3531182|T109|1366232|RXNORM|DIMETHICONOL (2000 CST)|DIMETHICONOL (2000 CST)
C0770958|T121|235786|RXNORM|CALCIUM OROTATE|CALCIUM OROTATE
C0017718|T121|4845|RXNORM|GLUCOSAMINE|GLUCOSAMINE
C2929513|T121|1008613|RXNORM|PHENOBARBITAL / PIPENZOLATE|PHENOBARBITAL / PIPENZOLATE
C2929512|T121|1008612|RXNORM|BENZOCAINE / METHYLBENZETHONIUM|BENZOCAINE / METHYLBENZETHONIUM
C2929511|T121|1008611|RXNORM|GARLIC PREPARATION / SOY LECITHIN|GARLIC PREPARATION / SOYBEAN LECITHIN
C2929510|T121|1008610|RXNORM|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PHENYLEPHRINE / PSEUDOEPHEDRINE / SCOPOLAMINE|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PHENYLEPHRINE / PSEUDOEPHEDRINE / SCOPOLAMINE
C2929517|T121|1008617|RXNORM|PANCREATIN / POTASSIUM BICARBONATE / SODIUM BICARBONATE|PANCREATIN / POTASSIUM BICARBONATE / SODIUM BICARBONATE
C2929516|T121|1008616|RXNORM|AMMONIUM CHLORIDE / GUAIACOLSULFONIC ACID|AMMONIUM CHLORIDE / GUAIACOLSULFONIC ACID
C2929515|T121|1008615|RXNORM|DICALCIUM PHOSPHATE / VITAMIN B 12|DICALCIUM PHOSPHATE / VITAMIN B 12
C2080573|T121|820128|RXNORM|BROMPHENIRAMINE / GUAIFENESIN / PHENYLPROPANOLAMINE|BROMPHENIRAMINE / GUAIFENESIN / PHENYLPROPANOLAMINE
C2929519|T121|1008619|RXNORM|BELLADONNA ALKALOIDS / CAFFEINE / ERGOTAMINE / PHENOBARBITAL|BELLADONNA ALKALOIDS / CAFFEINE / ERGOTAMINE / PHENOBARBITAL
C2929518|T121|1008618|RXNORM|ANTAZOLINE / TETRAHYDROZOLINE|ANTAZOLINE / TETRAHYDROZOLINE
C3257689|T121|1363437|RXNORM|LIME PEEL EXTRACT|LIME PEEL EXTRACT
C0246249|T197|72901|RXNORM|FERUMOXIDES|FERUMOXIDES
C1874470|T121|690057|RXNORM|BENDROFLUMETHIAZIDE / POTASSIUM CHLORIDE|BENDROFLUMETHIAZIDE / POTASSIUM CHLORIDE
C1874469|T121|690054|RXNORM|BENACTYZINE / MEPROBAMATE|BENACTYZINE / MEPROBAMATE
C3474581|T109|1363431|RXNORM|CAPRYLYL TRISILOXANE|CAPRYLYL TRISILOXANE
C3535620|T121|1370827|RXNORM|POLYETHYLENE GLYCOL 8000000|POLYETHYLENE GLYCOL 8000000
C2756541|T129|968492|RXNORM|BARLEY SMUT EXTRACT|USTILAGO NUDA EXTRACT
C0939224|T121|284628|RXNORM|CANDESARTAN / HYDROCHLOROTHIAZIDE|CANDESARTAN / HYDROCHLOROTHIAZIDE
C3538039|T121|1371911|RXNORM|PASSIFLORA INCARNATA SEED EXTRACT|PASSIFLORA INCARNATA SEED EXTRACT
C3535924|T121|1368916|RXNORM|GAMMA-AMINOBUTYRATE / MELATONIN / VALERIAN ROOT EXTRACT|GAMMA-AMINOBUTYRATE / MELATONIN / VALERIAN ROOT EXTRACT
C3538040|T122|1371912|RXNORM|TRIDECETH-5|TRIDECETH-5
C0043971|T121|1363030|RXNORM|1,3-PROPANEDIOL|1,3-PROPANEDIOL
C0772450|T121|237112|RXNORM|MYCOPHENOLATE MOFETIL HYDROCHLORIDE|MYCOPHENOLATE MOFETIL HYDROCHLORIDE
C0772453|T121|237115|RXNORM|GRAPE SEED|GRAPE SEED
C0772454|T121|237116|RXNORM|GRAPE SEED EXTRACT|GRAPE SEED EXTRACT
C0075478|T130|37296|RXNORM|SUCROSE OCTAACETATE|SUCROSE OCTAACETATE
C0073076|T121|35373|RXNORM|REPROTEROL|REPROTEROL
C0042646|T121|11194|RXNORM|VIDARABINE|VIDARABINE
C0042646|T121|11194|RXNORM|VIDARABINE|VIDARABINE
C3486798|T121|1311249|RXNORM|SUS SCROFA FRONTAL LOBE PREPARATION|PORCINE FRONTAL LOBE PREPARATION
C0042665|T121|11196|RXNORM|VILOXAZINE|VILOXAZINE
C3496026|T121|1311247|RXNORM|SUS SCROFA ANKLE JOINT PREPARATION|PORCINE ANKLE JOINT PREPARATION
C0042670|T123|11198|RXNORM|VINBLASTINE|VINBLASTINE
C3497927|T121|1311245|RXNORM|SUS SCROFA NERVE PREPARATION|PORCINE NERVE PREPARATION
C3497926|T121|1311244|RXNORM|SUS SCROFA LIMBIC SYSTEM PREPARATION|PORCINE LIMBIC SYSTEM PREPARATION
C3484424|T121|1311242|RXNORM|SUS SCROFA STOMACH PREPARATION|PORCINE STOMACH PREPARATION
C3487985|T121|1311241|RXNORM|SUS SCROFA PITUITARY GLAND PREPARATION|PORCINE PITUITARY GLAND PREPARATION
C3487984|T121|1311240|RXNORM|SUS SCROFA HYPOTHALAMUS PREPARATION|PORCINE HYPOTHALAMUS PREPARATION
C0873002|T121|259342|RXNORM|CAYENNE|CAYENNE EXTRACT
C0058156|T121|1362922|RXNORM|DIISOPROPANOLAMINE|DIISOPROPANOLAMINE
C0010711|T121|3041|RXNORM|CYTARABINE|CYTARABINE
C2701376|T129|852174|RXNORM|PUSSY WILLOW POLLEN EXTRACT|SALIX DISCOLOR POLLEN EXTRACT
C2194080|T121|819464|RXNORM|METOCLOPRAMIDE / SIMETHICONE|METOCLOPRAMIDE / SIMETHICONE
C0055630|T197|1539810|RXNORM|CHROMIUM TRIOXIDE|CHROMIUM TRIOXIDE
C1815835|T129|805486|RXNORM|VARICELLA VIRUS VACCINE LIVE (OKA-MERCK) STRAIN|VARICELLA VIRUS VACCINE LIVE (OKA-MERCK) STRAIN
C0028040|T131|7407|RXNORM|NICOTINE|NICOTINE
C0982199|T121|314666|RXNORM|HYDRASTIS PREPARATION|HYDRASTIS PREPARATION
C0078849|T121|40003|RXNORM|ZOTEPINE|ZOTEPINE
C3486790|T121|1310229|RXNORM|ECBALLIUM ELATERIUM FRUIT EXTRACT|ECBALLIUM ELATERIUM FRUIT EXTRACT
C3486770|T121|1310227|RXNORM|PIPER CUBEBA FRUIT EXTRACT|PIPER CUBEBA FRUIT EXTRACT
C0939870|T121|1310220|RXNORM|ACONITUM NAPELLUS EXTRACT|ACONITUM NAPELLUS EXTRACT
C3668773|T121|1441400|RXNORM|VITEX AGNUS-CASTUS WHOLE EXTRACT|VITEX AGNUS-CASTUS WHOLE EXTRACT
C3486584|T121|1311069|RXNORM|PORK BRAIN PREPARATION|PORK BRAIN PREPARATION
C0003765|T123|1091|RXNORM|ARGININE|ARGININE
C0003765|T123|1091|RXNORM|ARGININE|ARGININE
C2917638|T121|1311063|RXNORM|GIANT PUFFBALL EXTRACT|GIANT PUFFBALL EXTRACT
C3484411|T197|1311062|RXNORM|OYSTER SHELL CALCIUM CARBONATE PREPARATION|OYSTER SHELL CALCIUM CARBONATE PREPARATION
C0001699|T007|1311061|RXNORM|KLEBSIELLA PNEUMONIAE|KLEBSIELLA PNEUMONIAE
C3484410|T121|1311060|RXNORM|MUCUNA PRURIENS FRUIT TRICHOME EXTRACT|MUCUNA PRURIENS FRUIT TRICHOME EXTRACT
C0003779|T125|1098|RXNORM|ARGIPRESSIN|ARGIPRESSIN
C3489014|T121|1311066|RXNORM|SPONGIA OFFICINALIS SKELETON EXTRACT|SPONGIA OFFICINALIS SKELETON EXTRACT
C0052972|T197|1311065|RXNORM|BARIUM CHLORIDE|BARIUM CHLORIDE
C1721343|T121|662263|RXNORM|DORZOLAMIDE / TIMOLOL|DORZOLAMIDE / TIMOLOL
C3542442|T121|1428866|RXNORM|CARROT EXTRACT|DAUCUS CAROTA SUBSP. SATIVUS EXTRACT
C2699766|T121|1428867|RXNORM|DIETHADIONE|DIETHADIONE
C3651756|T109|1428864|RXNORM|CAPRYLYL TRIMETHICONE|CAPRYLYL TRIMETHICONE
C3651755|T122|1428865|RXNORM|CETETH-7|CETETH-7
C1619629|T121|614373|RXNORM|DEFERASIROX|DEFERASIROX
C3651757|T109|1428863|RXNORM|C10-36 OLEFIN|C10-36 OLEFIN
C3651759|T109|1428860|RXNORM|AZELAMIDE MONOETHANOLAMINE|AZELAMIDE MONOETHANOLAMINE
C1875437|T121|700826|RXNORM|LEVONORDEFRIN / MEPIVACAINE|LEVONORDEFRIN / MEPIVACAINE
C0304600|T121|91299|RXNORM|PIPERONYL BUTOXIDE / PYRETHRINS|PIPERONYL BUTOXIDE / PYRETHRINS
C3848580|T129|1546168|RXNORM|PEGINTERFERON BETA-1A|PEGINTERFERON BETA-1A
C3651754|T130|1428868|RXNORM|DISODIUM HEDTA|DISODIUM HEDTA
C0057936|T131|1428869|RXNORM|DIETHYL SULFATE|DIETHYL SULFATE
C3488643|T121|1309989|RXNORM|CELERY SEED EXTRACT|CELERY SEED EXTRACT
C3465264|T121|1309988|RXNORM|MORUS ALBA LEAF EXTRACT|MORUS ALBA LEAF EXTRACT
C3488234|T121|1309985|RXNORM|TARAXACUM PALUSTRE ROOT EXTRACT|TARAXACUM PALUSTRE ROOT EXTRACT
C3489041|T121|1309987|RXNORM|EUPATORIUM CANNABINUM EXTRACT|EUPATORIUM CANNABINUM FLOWERING TOP EXTRACT
C3488252|T121|1309986|RXNORM|FRAXINUS EXCELSIOR LEAF EXTRACT|FRAXINUS EXCELSIOR LEAF EXTRACT
C0772003|T121|1309981|RXNORM|RUBUS IDAEUS LEAF EXTRACT|RUBUS IDAEUS LEAF EXTRACT
C3465042|T109|1309980|RXNORM|SOYBEAN SEED OIL|SOYBEAN SEED OIL
C3484403|T121|1309983|RXNORM|SYMPLOCARPUS FOETIDUS ROOT EXTRACT|SYMPLOCARPUS FOETIDUS ROOT EXTRACT
C3486819|T121|1310112|RXNORM|SEMPERVIVUM TECTORUM LEAF EXTRACT|SEMPERVIVUM TECTORUM LEAF EXTRACT
C0065961|T121|29518|RXNORM|MEPINDOLOL|MEPINDOLOL
C3834071|T122|1541745|RXNORM|DIPENTAERYTHRITYL HEXASTEARATE|DIPENTAERYTHRITYL HEXASTEARATE
C3834072|T122|1541744|RXNORM|CHOLESTERYL ISOSTEARATE|CHOLESTERYL ISOSTEARATE
C0065374|T121|29046|RXNORM|LISINOPRIL|LISINOPRIL
C0162947|T109|1541746|RXNORM|METHYL RICINOLEATE|METHYL RICINOLEATE
C3834075|T122|1541741|RXNORM|HYDROXYPROPYL BISSTEARAMIDE MONOETHANOLAMIDE|HYDROXYPROPYL BISSTEARAMIDE MONOETHANOLAMIDE
C3714982|T122|1541740|RXNORM|TARAXACUM MONGOLICUM EXTRACT|TARAXACUM MONGOLICUM EXTRACT
C3834073|T122|1541743|RXNORM|TREHALOSE ISOSTEARATE ESTERS|TREHALOSE ISOSTEARATE ESTERS
C0305007|T197|91559|RXNORM|SODIUM PHOSPHATE P32|SODIUM PHOSPHATE (32P)
C0004718|T121|1321|RXNORM|BAMETHAN|BAMETHAN
C0004743|T121|1325|RXNORM|BARBITAL|BARBITAL
C2146623|T121|812243|RXNORM|ACETAMINOPHEN / CAFFEINE / MAGNESIUM SALICYLATE|ACETAMINOPHEN / CAFFEINE / MAGNESIUM SALICYLATE
C2194017|T121|812242|RXNORM|BETAMETHASONE / CHLORPHENIRAMINE|BETAMETHASONE / CHLORPHENIRAMINE
C0876880|T121|262231|RXNORM|HYOSCYAMINE / METHENAMINE|HYOSCYAMINE / METHENAMINE
C0529793|T121|136411|RXNORM|SILDENAFIL|SILDENAFIL
C0529793|T121|136411|RXNORM|SILDENAFIL|SILDENAFIL
C0025826|T125|6904|RXNORM|METHYLTESTOSTERONE|METHYLTESTOSTERONE
C0033124|T121|8686|RXNORM|PRILOCAINE|PRILOCAINE
C0033126|T121|8687|RXNORM|PRIMAQUINE|PRIMAQUINE
C0025810|T121|6901|RXNORM|METHYLPHENIDATE|METHYLPHENIDATE
C0023899|T121|6459|RXNORM|LIVER EXTRACT|LIVER EXTRACT
C2928417|T121|1007495|RXNORM|RED CLOVER PREPARATION / SOYBEAN PREPARATION / VITAMIN E|RED CLOVER PREPARATION / SOYBEAN PREPARATION / VITAMIN E
C2928418|T121|1007496|RXNORM|APPLE PECTIN / LACTOBACILLUS ACIDOPHILUS|APPLE PECTIN / LACTOBACILLUS ACIDOPHILUS
C2928419|T121|1007497|RXNORM|GARLIC PREPARATION / GINKGO BILOBA EXTRACT / GINSENG PREPARATION|GARLIC PREPARATION / GINKGO BILOBA EXTRACT / GINSENG PREPARATION
C2928412|T121|1007490|RXNORM|ALUM, POTASSIUM / LIDOCAINE|ALUM, POTASSIUM / LIDOCAINE
C3152842|T129|1098200|RXNORM|NEUROSPORA SITOPHILA EXTRACT|NEUROSPORA SITOPHILA EXTRACT
C2928414|T121|1007492|RXNORM|BENZYDAMINE / BROMHEXINE|BENZYDAMINE / BROMHEXINE
C0031411|T121|8133|RXNORM|PHENMETRAZINE|PHENMETRAZINE
C0216278|T121|69646|RXNORM|TINZAPARIN|TINZAPARIN
C3486694|T121|1346618|RXNORM|GALPHIMIA GLAUCA FLOWERING TOP EXTRACT|GALPHIMIA GLAUCA FLOWERING TOP EXTRACT
C3486704|T121|1346619|RXNORM|GERANIUM MACULATUM ROOT EXTRACT|GERANIUM MACULATUM ROOT EXTRACT
C3667111|T121|1438637|RXNORM|OCTYL SULFATE|OCTYL SULFATE
C3486663|T121|1346616|RXNORM|CALTHA PALUSTRIS EXTRACT|CALTHA PALUSTRIS EXTRACT
C3486682|T121|1346617|RXNORM|BLATTA ORIENTALIS PREPARATION|ORIENTAL COCKROACH PREPARATION
C3256019|T121|1307567|RXNORM|BETULA PLATYPHYLLA VAR JAPONICA RESIN|BETULA PLATYPHYLLA VAR JAPONICA RESIN
C2702400|T129|867198|RXNORM|CLADOSPORIUM CLADOSPORIOIDES EXTRACT|CLADOSPORIUM CLADOSPORIOIDES EXTRACT
C2928144|T121|1007222|RXNORM|FORMALDEHYDE / GLUTARAL / GLYOXAL|FORMALDEHYDE / GLUTARAL / GLYOXAL
C0939819|T121|285168|RXNORM|VERATRUM ALBUM PREPARATION|VERATRUM ALBUM PREPARATION
C0060245|T197|24912|RXNORM|FERRIC SUBSULFATE SOLUTION|MONSEL'S SOLUTION
C0031962|T131|8345|RXNORM|PIPERONYL BUTOXIDE|PIPERONYL BUTOXIDE
C3256218|T109|1307560|RXNORM|CYDONIA OBLONGA SEED EXTRACT|CYDONIA OBLONGA SEED EXTRACT
C0873010|T121|259350|RXNORM|MIRANOL 2MHT MODIFIED|MIRANOL 2MHT MODIFIED
C3666982|T121|1438109|RXNORM|LYCOPODIUM COMPLANATUM WHOLE EXTRACT|LYCOPODIUM COMPLANATUM WHOLE EXTRACT
C0873018|T121|259357|RXNORM|BORON GLUCONATE|BORON GLUCONATE
C1445380|T129|892539|RXNORM|CLAM ALLERGENIC EXTRACT|CLAM ALLERGENIC EXTRACT
C0353697|T121|103990|RXNORM|CARBIDOPA / LEVODOPA|CARBIDOPA / LEVODOPA
C0047231|T121|1435285|RXNORM|3-AMINOPHENOL|M-AMINOPHENOL
C0016913|T007|1592903|RXNORM|ANAEROCOCCUS TETRADIUS|ANAEROCOCCUS TETRADIUS
C0031978|T121|8352|RXNORM|PIRENZEPINE|PIRENZEPINE
C0031979|T121|8353|RXNORM|PIRIBEDIL|PIRIBEDIL
C0031982|T121|8354|RXNORM|PIRINITRAMIDE|PIRINITRAMIDE
C0031990|T121|8356|RXNORM|PIROXICAM|PIROXICAM
C1874354|T121|689498|RXNORM|ASCORBIC ACID / NIACIN|ASCORBIC ACID / NIACIN
C3651786|T121|1428413|RXNORM|CALCIUM HYDRIDE|CALCIUM HYDRIDE
C0072973|T121|35296|RXNORM|RAMIPRIL|RAMIPRIL
C3859428|T007|1592901|RXNORM|MORAXELLA CATARRHALIS SUBSP. CATARRHALIS|MORAXELLA CATARRHALIS SUBSP. CATARRHALIS
C0057908|T109|1593447|RXNORM|DIDODECYL PHOSPHATE|DIDODECYL PHOSPHATE
C3256849|T109|1427202|RXNORM|LAURYL PCA|LAURYL PIDOLATE
C3859630|T121|1593448|RXNORM|2,5-DI-TERT-PENTYLHYDROQUINONE|2,5-DI-TERT-PENTYLHYDROQUINONE
C3859427|T121|1592900|RXNORM|POLYGONATUM CYRTONEMA ROOT EXTRACT|POLYGONATUM CYRTONEMA ROOT EXTRACT
C1874350|T121|689494|RXNORM|ASCORBIC ACID / HESPERIDIN|ASCORBIC ACID / HESPERIDIN
C3489069|T121|1355185|RXNORM|FOMITOPSIS PINICOLA FRUITING BODY EXTRACT|FOMITOPSIS PINICOLA FRUITING BODY EXTRACT
C2079567|T121|814600|RXNORM|NORTRIPTYLINE / PERPHENAZINE|NORTRIPTYLINE / PERPHENAZINE
C0059678|T121|24441|RXNORM|ETIFOXINE|ETIFOXINE
C0358712|T121|106732|RXNORM|CLEMASTINE / PHENYLPROPANOLAMINE|CLEMASTINE / PHENYLPROPANOLAMINE
C3465352|T122|1427207|RXNORM|SYNTHETIC WAX (1900 MW)|SYNTHETIC WAX (1900 MW)
C0117953|T130|50110|RXNORM|DICHLORODIFLUOROMETHANE|DICHLORODIFLUOROMETHANE
C2740876|T129|899916|RXNORM|SCALLOP ALLERGENIC EXTRACT|SCALLOP ALLERGENIC EXTRACT
C3282116|T121|1307729|RXNORM|PAEONIA SUFFRUTICOSA ROOT BARK EXTRACT|PAEONIA SUFFRUTICOSA ROOT BARK EXTRACT
C3651953|T121|1428137|RXNORM|CHLOPHEDIANOL / THONZYLAMINE|CHLOPHEDIANOL / THONZYLAMINE
C0717652|T121|214452|RXNORM|COLCHICINE / PROBENECID|COLCHICINE / PROBENECID
C0717650|T121|214450|RXNORM|CODEINE / PHENYLEPHRINE / PYRILAMINE|CODEINE / PHENYLEPHRINE / PYRILAMINE
C0717651|T121|214451|RXNORM|CODEINE / PSEUDOEPHEDRINE / TRIPROLIDINE|CODEINE / PSEUDOEPHEDRINE / TRIPROLIDINE
C3257189|T168|1307723|RXNORM|RASPBERRY JUICE|RUBUS IDAEUS JUICE
C3255784|T109|1307722|RXNORM|OAT KERNEL OIL|OAT KERNEL OIL
C0772361|T121|1307721|RXNORM|WHITE MULBERRY EXTRACT|WHITE MULBERRY EXTRACT
C3256537|T121|1307720|RXNORM|FERULA ASSA-FOETIDA ROOT EXTRACT|FERULA ASSA-FOETIDA ROOT EXTRACT
C3256754|T121|1307727|RXNORM|CANNA INDICA ROOT EXTRACT|CANNA INDICA ROOT EXTRACT
C3255858|T121|1307726|RXNORM|PANAX GINSENG FLOWER EXTRACT|PANAX GINSENG FLOWER EXTRACT
C3281945|T121|1307724|RXNORM|MYRCIARIA DUBIA SEED EXTRACT|MYRCIARIA DUBIA SEED EXTRACT
C2939834|T121|1014182|RXNORM|CALCIUM CITRATE / ERGOCALCIFEROL / MAGNESIUM OXIDE|CALCIUM CITRATE / ERGOCALCIFEROL / MAGNESIUM OXIDE
C3714904|T121|1546352|RXNORM|2,3-DIMERCAPTO-1-PROPANESULFONIC ACID|2,3-DIMERCAPTO-1-PROPANESULFONIC ACID
C2701673|T129|852597|RXNORM|UTAH JUNIPER POLLEN EXTRACT|JUNIPERUS OSTEOSPERMA POLLEN EXTRACT
C2342892|T121|794809|RXNORM|MENTHOL / ZINC OXIDE|MENTHOL / ZINC OXIDE
C3848625|T121|1544131|RXNORM|PLECTRANTHUS BARBATUS WHOLE EXTRACT|PLECTRANTHUS BARBATUS WHOLE EXTRACT
C3667887|T109|1440254|RXNORM|ETHYL PALMATE|ETHYL PALMATE
C3848624|T109|1544135|RXNORM|VINYLPYRROLIDONE-EICOSENE COPOLYMER|VINYLPYRROLIDONE-EICOSENE COPOLYMER
C3857947|T121|1552448|RXNORM|BOS TAURUS ESOPHAGUS PREPARATION|BOS TAURUS ESOPHAGUS PREPARATION
C3848622|T121|1544137|RXNORM|BOS TAURUS LYMPH VESSEL PREPARATION|BOS TAURUS LYMPH VESSEL PREPARATION
C3848623|T121|1544136|RXNORM|BOS TAURUS CONJUNCTIVA PREPARATION|BOS TAURUS CONJUNCTIVA PREPARATION
C2194234|T121|819156|RXNORM|SALICYLIC ACID / TRICLOSAN|SALICYLIC ACID / TRICLOSAN
C3818685|T109|1537759|RXNORM|TRIMETHYLSILYL TREATED DIIMETHICONOL-TRIMETHYLSILOXYSILICATE CROSSPOLYMER (40-60 WW)|TRIMETHYLSILYL TREATED DIIMETHICONOL-TRIMETHYLSILOXYSILICATE CROSSPOLYMER (40-60 WW)
C3818686|T109|1537758|RXNORM|COMMIPHORA AFRICANA RESIN|COMMIPHORA AFRICANA RESIN
C0055151|T121|20614|RXNORM|CETRIMONIUM|CETRIMONIUM
C0995182|T121|318340|RXNORM|ALOE VERA PREPARATION|ALOE VERA PREPARATION
C3815858|T121|1537753|RXNORM|VALERIANA OFFICINALIS WHOLE EXTRACT|VALERIANA OFFICINALIS WHOLE EXTRACT
C0719127|T121|215858|RXNORM|CAMPHOR / PHENOL|CAMPHOR / PHENOL
C3818689|T121|1537751|RXNORM|WOOD TAR HYDROCARBON DISTILLATE|WOOD TAR HYDROCARBON DISTILLATE
C0051721|T197|17789|RXNORM|AMMONIUM MOLYBDATE|AMMONIUM MOLYBDATE
C3818687|T121|1537757|RXNORM|GLECHOMA LONGITUBA WHOLE EXTRACT|GLECHOMA LONGITUBA WHOLE EXTRACT
C3814375|T121|1537756|RXNORM|ARGEMONE MEXICANA EXTRACT|ARGEMONE MEXICANA EXTRACT
C0074027|T121|1537755|RXNORM|SANGUINARINE|SANGUINARINE
C0021252|T121|5784|RXNORM|INDORAMIN|INDORAMIN
C0021246|T121|5781|RXNORM|INDOMETHACIN|INDOMETHACIN
C0021246|T121|5781|RXNORM|INDOMETHACIN|INDOMETHACIN
C0876715|T121|262099|RXNORM|PHENAZOPYRIDINE / SULFAMETHOXAZOLE|PHENAZOPYRIDINE / SULFAMETHOXAZOLE
C1445822|T121|466588|RXNORM|ALUMINUM HYDROXIDE / MAGNESIUM HYDROXIDE / SIMETHICONE|ALUMINUM HYDROXIDE / MAGNESIUM HYDROXIDE / SIMETHICONE
C1176308|T121|358257|RXNORM|TOLVAPTAN|TOLVAPTAN
C1176306|T121|358255|RXNORM|APREPITANT|APREPITANT
C1337367|T121|408114|RXNORM|GOLDEN SEAL EXTRACT|GOLDEN SEAL EXTRACT
C3709740|T121|1488226|RXNORM|GALIUM BOREALE LEAF EXTRACT|GALIUM BOREALE LEAF EXTRACT
C1445815|T121|466581|RXNORM|ACETAMINOPHEN / CAFFEINE / SALICYLAMIDE|ACETAMINOPHEN / CAFFEINE / SALICYLAMIDE
C1176309|T121|358258|RXNORM|BORTEZOMIB|BORTEZOMIB
C0617623|T121|166283|RXNORM|LIDOCAINE / PRILOCAINE|LIDOCAINE / PRILOCAINE
C0617623|T121|166283|RXNORM|LIDOCAINE / PRILOCAINE|LIDOCAINE / PRILOCAINE
C1445818|T121|466584|RXNORM|ACETAMINOPHEN / ASPIRIN / CAFFEINE|ACETAMINOPHEN / ASPIRIN / CAFFEINE
C2929598|T121|1008698|RXNORM|ATROPINE / CARZENIDE / DIPYRONE|ATROPINE / CARZENIDE / DIPYRONE
C3848521|T196|1546440|RXNORM|HYPOPHOSPHITE ION|HYPOPHOSPHITE ION
C2701549|T129|852376|RXNORM|BLACK COTTONWOOD POLLEN EXTRACT|POPULUS TRICHOCARPA POLLEN EXTRACT
C3668709|T121|1441297|RXNORM|AGARICUS CAMPESTRIS VAR. CAMPESTRIS WHOLE EXTRACT|AGARICUS CAMPESTRIS VAR. CAMPESTRIS WHOLE EXTRACT
C2939957|T129|1014360|RXNORM|LONGLEAF PINE POLLEN EXTRACT|PINUS PALUSTRIS POLLEN EXTRACT
C0034272|T127|684879|RXNORM|PYRIDOXINE|PYRIDOXINE
C2920812|T129|999487|RXNORM|WHEAT STEM RUST EXTRACT|PUCCINIA GRAMINIS EXTRACT
C0303208|T197|90402|RXNORM|CHROMIC SULFATE|CHROMIC SULFATE
C1330007|T121|404802|RXNORM|GUAIFENESIN / PHENYLEPHRINE / PYRILAMINE|GUAIFENESIN / PHENYLEPHRINE / PYRILAMINE
C0538927|T121|140587|RXNORM|CELECOXIB|CELECOXIB
C2194146|T121|816628|RXNORM|MAZINDOL / TIRATRICOL|MAZINDOL / TIRATRICOL
C0043501|T130|11431|RXNORM|ZINC-DTPA|ZINC-DTPA
C3256425|T121|1307738|RXNORM|PHRAGMITES AUSTRALIS ROOT EXTRACT|PHRAGMITES AUSTRALIS ROOT EXTRACT
C3256740|T121|1307739|RXNORM|VACCINIUM ANGUSTIFOLIUM LEAF EXTRACT|VACCINIUM ANGUSTIFOLIUM LEAF EXTRACT
C2364553|T129|805553|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED B-FLORIDA-4-2006 STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED B-FLORIDA-4-2006 STRAIN
C2961528|T121|1053120|RXNORM|ASPIRIN / DEXTROMETHORPHAN / DOXYLAMINE / PHENYLEPHRINE|ASPIRIN / DEXTROMETHORPHAN / DOXYLAMINE / PHENYLEPHRINE
C0016282|T121|4453|RXNORM|FLUFENAMIC ACID|FLUFENAMIC ACID
C0016280|T125|4452|RXNORM|FLUDROCORTISONE|FLUDROCORTISONE
C0016278|T121|4451|RXNORM|FLUCYTOSINE|FLUCYTOSINE
C0016277|T121|4450|RXNORM|FLUCONAZOLE|FLUCONAZOLE
C0016293|T121|4457|RXNORM|FLUMAZENIL|FLUMAZENIL
C2827104|T122|1305738|RXNORM|CARBOMER HOMOPOLYMER TYPE C|CARBOMER 980
C0016295|T121|4459|RXNORM|FLUNARIZINE|FLUNARIZINE
C2827146|T121|1305739|RXNORM|ETHYLCELLULOSE (100 MPA S)|ETHYLCELLULOSE (100 MPA S)
C0071123|T121|33761|RXNORM|PIPROZOLINE|PIPROZOLINE
C0048207|T121|1485787|RXNORM|4-COUMARIC ACID|4-COUMARIC ACID
C1620322|T109|1356761|RXNORM|ASCORBYL TETRAISOPALMITATE|ASCORBYL TETRAISOPALMITATE
C3504850|T109|1356760|RXNORM|SUCROSE TETRAISOSTEARATE|SUCROSE TETRAISOSTEARATE
C3464654|T121|1356763|RXNORM|SILK, ACID HYDROLYZED (1000 MW)|SILK, ACID HYDROLYZED (1000 MW)
C0058623|T121|37534|RXNORM|TADENAN|TADENAN
C1451182|T109|1356765|RXNORM|DIOCTYL MALEATE|DIOCTYL MALEATE
C3504851|T109|1356764|RXNORM|POLYACRYLAMIDE (1300000 MW)|POLYACRYLAMIDE (1300000 MW)
C3256629|T109|1356767|RXNORM|POLYGLYCERYL-10 OLEATE|POLYGLYCERYL-10 OLEATE
C3504852|T109|1356766|RXNORM|PEG-PPG-14-7 DIMETHYL ETHER|PEG-PPG-14-7 DIMETHYL ETHER
C0074758|T197|36710|RXNORM|TRIBASIC SODIUM PHOSPHATE|TRIBASIC SODIUM PHOSPHATE
C3504853|T109|1356768|RXNORM|SODIUM METHYL STEAROYL TAURATE|SODIUM METHYL STEAROYL TAURATE
C0250480|T121|74169|RXNORM|PIPERACILLIN / TAZOBACTAM|PIPERACILLIN / TAZOBACTAM
C0074765|T197|36717|RXNORM|SODIUM SELENATE|SODIUM SELENATE
C0060187|T121|24860|RXNORM|FENOZOLONE|FENOZOLONE
C0060194|T121|24867|RXNORM|FENPROPOREX|FENPROPOREX
C2741022|T129|900131|RXNORM|TAMARACK POLLEN EXTRACT|LARIX OCCIDENTALIS POLLEN EXTRACT
C0055860|T195|21216|RXNORM|CLAVULANIC ACID|CLAVULANIC ACID
C1630394|T121|608868|RXNORM|ETHINYL ESTRADIOL / GESTODENE|ETHINYL ESTRADIOL / GESTODENE
C0002083|T121|508|RXNORM|ALLANTOIN|ALLANTOIN
C0066805|T121|30227|RXNORM|MOROXYDINE|MOROXYDINE
C3848577|T197|1546210|RXNORM|GOLD MONOSULFIDE|GOLD MONOSULFIDE
C2146624|T121|820463|RXNORM|ACETAMINOPHEN / MELATONIN|ACETAMINOPHEN / MELATONIN
C3256603|T121|1423924|RXNORM|CORN GRAIN EXTRACT|CORN MEAL EXTRACT
C0077666|T126|1423925|RXNORM|UBIQUINONE Q2|UBIQUINONE Q2
C0056037|T197|1423923|RXNORM|COBALTOUS NITRATE|COBALTOUS NITRATE
C3643348|T121|1423921|RXNORM|ESCHSCHOLZIA CALIFORNICA FLOWERING TOP EXTRACT|CALIFORNIA POPPY FLOWERING TOP EXTRACT
C3818722|T109|1535452|RXNORM|AESCULUS HIPPOCASTANUM SEED OIL|AESCULUS HIPPOCASTANUM SEED OIL
C3818721|T121|1535457|RXNORM|CERITINIB|CERITINIB
C1723401|T129|1092437|RXNORM|BELIMUMAB|BELIMUMAB
C3833035|T121|1540240|RXNORM|VACCINIUM ANGUSTIFOLIUM WHOLE EXTRACT|VACCINIUM ANGUSTIFOLIUM WHOLE EXTRACT
C0771436|T121|236186|RXNORM|TENONITROZOLE|TENONITROZOLE
C0044548|T121|12166|RXNORM|1-OCTACOSANOL|1-OCTACOSANOL
C0537147|T121|139778|RXNORM|TEGASEROD|TEGASEROD
C0022181|T131|6027|RXNORM|SACCHAROMYCES BOULARDII LYO|ISOFLUROPHATE
C0771438|T121|236188|RXNORM|TIEMONIUM|TIEMONIUM
C0537670|T129|139994|RXNORM|OPRELVEKIN|OPRELVEKIN
C0165477|T121|1546379|RXNORM|TRANDOLAPRILAT|TRANDOLAPRILAT
C3848548|T130|1546378|RXNORM|ROSE BENGAL AT|ROSE BENGAL AT
C3848551|T196|1546370|RXNORM|THALLOUS CATION TL-201|THALLOUS CATION TL-201
C0303225|T196|1546372|RXNORM|GALLIUM-67|GALLIUM-67
C3848549|T196|1546374|RXNORM|GOLD CATION (3+)|GOLD CATION (3+)
C0072970|T121|1546377|RXNORM|RAMIPRILAT|RAMIPRILAT
C0083236|T197|1546376|RXNORM|LITHIUM HYDROXIDE|LITHIUM HYDROXIDE
C0039832|T121|10450|RXNORM|THIABENDAZOLE|THIABENDAZOLE
C0038425|T195|10109|RXNORM|STREPTOMYCIN|STREPTOMYCIN
C0036720|T123|9671|RXNORM|SERINE|SERINE
C0039840|T127|10454|RXNORM|THIAMINE|THIAMINE (VIT B1)
C0038416|T121|10105|RXNORM|STREPTODORNASE / STREPTOKINASE|STREPTODORNASE / STREPTOKINASE
C0038415|T126|10104|RXNORM|STREPTODORNASE|STREPTODORNASE
C0038418|T126|10106|RXNORM|STREPTOKINASE|STREPTOKINASE
C0056519|T121|21766|RXNORM|CROTAMITON|CROTAMITON
C2740585|T129|899355|RXNORM|BASIL ALLERGENIC EXTRACT|OCIMUM BASILICUM ALLERGENIC EXTRACT
C3256859|T121|1427009|RXNORM|PROPYLENE GLYCOL DICAPRATE|PROPYLENE GLYCOL DICAPRATE
C0981976|T129|899359|RXNORM|SUGAR BEET ALLERGENIC EXTRACT|BETA VULGARIS ALLERGENIC EXTRACT
C2741458|T129|901265|RXNORM|WHITE FISH ALLERGENIC EXTRACT|WHITE FISH ALLERGENIC EXTRACT
C0772323|T109|236988|RXNORM|WHITE BRYONY EXTRACT|WHITE BRYONY EXTRACT
C0772078|T121|236768|RXNORM|SULFATED MUCOPOLYSACCHARIDES|SULFATED MUCOPOLYSACCHARIDES
C0090306|T121|43611|RXNORM|LATANOPROST|LATANOPROST ACID
C0071102|T121|33742|RXNORM|PIPECURONIUM|PIPECURONIUM
C0772321|T130|236987|RXNORM|MANGAFODIPIR|MANGAFODIPIR
C0939895|T121|285241|RXNORM|GINGER EXTRACT|GINGER EXTRACT
C0939894|T121|285240|RXNORM|VERATRUM VIRIDE PREPARATION|VERATRUM VIRIDE PREPARATION
C0939897|T121|285243|RXNORM|ALFALFA PREPARATION|ALFALFA PREPARATION
C0071108|T125|33747|RXNORM|ESTROPIPATE|ESTROPIPATE
C0071108|T125|33747|RXNORM|ESTROPIPATE|ESTROPIPATE
C2344304|T129|798279|RXNORM|HAEMOPHILUS INFLUENZAE TYPE B, CAPSULAR POLYSACCHARIDE INACTIVATED TETANUS TOXOID CONJUGATE VACCINE|HAEMOPHILUS INFLUENZAE TYPE B, CAPSULAR POLYSACCHARIDE INACTIVATED TETANUS TOXOID CONJUGATE VACCINE
C0066795|T121|30218|RXNORM|MORAZONE|MORAZONE
C3692449|T121|1442093|RXNORM|AFOXOLANER|AFOXOLANER
C0163082|T121|59094|RXNORM|CYCLOPENTAMINE|CYCLOPENTAMINE
C0105583|T130|1313278|RXNORM|BENZENESULFONATE|BENZENESULFONATE
C2726174|T129|891637|RXNORM|KIDNEY BEAN ALLERGENIC EXTRACT|KIDNEY BEAN ALLERGENIC EXTRACT
C0004954|T123|1359|RXNORM|LINALOOL, (-)-|BELLADONNA ALKALOIDS
C2702332|T129|891633|RXNORM|HAZELNUT ALLERGENIC EXTRACT|HAZELNUT ALLERGENIC EXTRACT
C3505681|T121|1359088|RXNORM|PINUS LAMBERTIANA RESIN|PINUS LAMBERTIANA RESIN
C3498012|T121|1314222|RXNORM|TAXUS BACCATA FRUIT EXTRACT|TAXUS BACCATA FRUIT EXTRACT
C3498009|T109|1314223|RXNORM|METHYL SORBATE|METHYL SORBATE
C0144544|T121|1314221|RXNORM|TARTRATE|TARTRATE
C3474308|T121|1314226|RXNORM|SYRINGA VULGARIS WHOLE EXTRACT|SYRINGA VULGARIS WHOLE EXTRACT
C0243264|T121|1314227|RXNORM|HYDROXYTYROSOL|HYDROXYTYROSOL
C3497919|T121|1314224|RXNORM|SANTALUM ALBUM SEED EXTRACT|SANTALUM ALBUM SEED EXTRACT
C3282691|T121|1314225|RXNORM|TETRADECENE|TETRADECENE
C3496662|T121|1314228|RXNORM|MUSA BASJOO WHOLE EXTRACT|MUSA BASJOO WHOLE EXTRACT
C3282785|T121|1314229|RXNORM|TETRAPROPYL ORTHOSILICATE|TETRAPROPYL ORTHOSILICATE
C3831982|T121|1538287|RXNORM|CALCIUM CARBONATE / POTASSIUM BICARBONATE / SODIUM BICARBONATE|CALCIUM CARBONATE / POTASSIUM BICARBONATE / SODIUM BICARBONATE
C0119860|T121|1085955|RXNORM|POLYSULFATED GLYCOSAMINOGLYCAN|POLYSULFATED GLYCOSAMINOGLYCAN
C3505677|T121|1359084|RXNORM|BIS-HYDROXYETHOXYPROPYL DIMETHICONE (50 CST)|BIS-HYDROXYETHOXYPROPYL DIMETHICONE (50 CST)
C1445191|T129|892851|RXNORM|DUCK FEATHER EXTRACT|ANAS PLATYRHYNCHOS FEATHER EXTRACT
C2702377|T129|892584|RXNORM|SALMON ALLERGENIC EXTRACT|SALMON ALLERGENIC EXTRACT
C3505680|T109|1359087|RXNORM|PEG-55 HYDROGENATED CASTOR OIL|PEG-55 HYDROGENATED CASTOR OIL
C3528000|T121|1546446|RXNORM|OMACETAXINE|OMACETAXINE
C2723711|T129|867297|RXNORM|PLAINS COTTONWOOD POLLEN EXTRACT|POPULUS DELTOIDES SUBSP. MONILIFERA POLLEN EXTRACT
C0002328|T121|595|RXNORM|ALGESTONE|ALGESTONE
C0002327|T121|594|RXNORM|ALPHAPRODINE|ALPHAPRODINE
C0002334|T121|597|RXNORM|ALPRENOLOL|ALPRENOLOL
C1722260|T121|1114326|RXNORM|INDACATEROL|INDACATEROL
C0002340|T123|599|RXNORM|ALSEROXYLON|ALSEROXYLON
C0002335|T121|598|RXNORM|ALPROSTADIL|ALPROSTADIL
C2241685|T121|761364|RXNORM|DIHYDROCODEINE / PHENYLEPHRINE|DIHYDROCODEINE / PHENYLEPHRINE
C0059471|T121|24274|RXNORM|EPROZINOL|EPROZINOL
C0059469|T121|24272|RXNORM|EPRAZINONE|EPRAZINONE
C0532699|T121|137732|RXNORM|CHROMIUM NICOTINIC ACID COMPLEX|CHROMIUM NICOTINIC ACID COMPLEX
C2929332|T121|1008428|RXNORM|CHLORHEXIDINE / PHENYLEPHRINE|CHLORHEXIDINE / PHENYLEPHRINE
C2929333|T121|1008429|RXNORM|BUZEPIDE METIODIDE / HALOPERIDOL|BUZEPIDE METIODIDE / HALOPERIDOL
C0012191|T121|3384|RXNORM|DIETHYLCARBAMAZINE|DIETHYLCARBAMAZINE
C0064113|T121|28031|RXNORM|ITRACONAZOLE|ITRACONAZOLE
C2929324|T121|1008420|RXNORM|ASCORBIC ACID / CALCIUM PHOSPHATE|ASCORBIC ACID / CALCIUM PHOSPHATE
C2929325|T121|1008421|RXNORM|ALLANTOIN / COAL TAR / LACTATE|ALLANTOIN / COAL TAR / LACTATE
C2929326|T121|1008422|RXNORM|ASCORBIC ACID / BIOTIN|ASCORBIC ACID / BIOTIN
C2929327|T121|1008423|RXNORM|BUTETAMATE / HELICIN|BUTETAMATE / HELICIN
C2929328|T121|1008424|RXNORM|CETRIMONIUM / LIDOCAINE / TYROTHRICIN|CETRIMONIUM / LIDOCAINE / TYROTHRICIN
C2929329|T121|1008425|RXNORM|HYDROCORTISONE / HYDROQUINONE / TRETINOIN|HYDROCORTISONE / HYDROQUINONE / TRETINOIN
C2929330|T121|1008426|RXNORM|LIDOCAINE / METHYL SALICYLATE / ZINC OXIDE|LIDOCAINE / METHYL SALICYLATE / ZINC OXIDE
C2929331|T121|1008427|RXNORM|ACEXAMIC ACID / NEOMYCIN|ACEXAMIC ACID / NEOMYCIN
C2928315|T121|1007393|RXNORM|BISMUTH SUBGALLATE / PHTHALYLSULFATHIAZOLE|BISMUTH SUBGALLATE / PHTHALYLSULFATHIAZOLE
C2928314|T121|1007392|RXNORM|SQUALENE / VITAMIN E|SQUALENE / VITAMIN E
C2928742|T121|1007827|RXNORM|ACETAMINOPHEN / PAMABROM / VITAMIN E|ACETAMINOPHEN / PAMABROM / VITAMIN E
C2928312|T121|1007390|RXNORM|SODIUM FLUORIDE / STANNOUS FLUORIDE|SODIUM FLUORIDE / STANNOUS FLUORIDE
C2928736|T121|1007821|RXNORM|CYCLOMETHYCAINE / DIPHENHYDRAMINE|CYCLOMETHYCAINE / DIPHENHYDRAMINE
C2928735|T121|1007820|RXNORM|AMYLASES / ENDOPEPTIDASES / LIPASE|AMYLASES / ENDOPEPTIDASES / LIPASE
C2928738|T121|1007823|RXNORM|CYCLONIUM / IBUPROFEN|CYCLONIUM / IBUPROFEN
C1874514|T121|690261|RXNORM|BENZOCAINE / CHLOROXYLENOL / ZINC OXIDE|BENZOCAINE / CHLOROXYLENOL / ZINC OXIDE
C1874516|T121|690263|RXNORM|BENZOCAINE / CLOVE OIL|BENZOCAINE / CLOVE OIL
C2928320|T121|1007398|RXNORM|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / INTRINSIC FACTOR|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / INTRINSIC FACTOR
C2928744|T121|1007829|RXNORM|ECHINACEA PURPUREA EXTRACT / GOLDEN SEAL EXTRACT|ECHINACEA PURPUREA EXTRACT / GOLDEN SEAL EXTRACT
C2928743|T121|1007828|RXNORM|BENZOCAINE / ZINC CHLORIDE|BENZOCAINE / ZINC CHLORIDE
C1874518|T121|690267|RXNORM|BENZOCAINE / ICHTHAMMOL|BENZOCAINE / ICHTHAMMOL
C3852512|T121|1597381|RXNORM|DASABUVIR|DASABUVIR
C0087064|T123|1364853|RXNORM|TAURINE DEOXYCHOLATE|TAURINE DEOXYCHOLATE
C1120386|T195|325887|RXNORM|MICAFUNGIN|MICAFUNGIN
C0065992|T197|1311475|RXNORM|MERCURIC SULFATE|MERCURIC SULFATE
C0006223|T196|1311476|RXNORM|BROMINE|BROMINE
C3256412|T121|1311477|RXNORM|CHONDRUS CRISPUS EXTRACT|CHONDRUS CRISPUS EXTRACT
C2012248|T121|821174|RXNORM|ASCORBIC ACID / GLUCOSE|ASCORBIC ACID / GLUCOSE
C0007016|T197|1311478|RXNORM|CARBON DISULFIDE|CARBON DISULFIDE
C3256678|T121|1311479|RXNORM|FRANKINCENSE EXTRACT|FRANKINCENSE EXTRACT
C1109213|T121|324007|RXNORM|DICRESULENE POLYMER|DICRESULENE POLYMER
C1445383|T121|1319268|RXNORM|ANTHOXANTHUM ODORATUM EXTRACT|ANTHOXANTHUM ODORATUM EXTRACT
C2203711|T121|813863|RXNORM|ASCORBIC ACID / ZINC SULFATE|ASCORBIC ACID / ZINC SULFATE
C0066621|T121|30077|RXNORM|MIVACURIUM|MIVACURIUM
C0939216|T121|284620|RXNORM|ABACAVIR / LAMIVUDINE / ZIDOVUDINE|ABACAVIR / LAMIVUDINE / ZIDOVUDINE
C0939218|T121|284622|RXNORM|ARTICAINE / EPINEPHRINE|ARTICAINE / EPINEPHRINE
C0939219|T121|284623|RXNORM|ATOVAQUONE / PROGUANIL|ATOVAQUONE / PROGUANIL
C0359015|T121|106960|RXNORM|CHLORAMPHENICOL / HYDROCORTISONE|CHLORAMPHENICOL / HYDROCORTISONE
C3247503|T121|1192515|RXNORM|BENZETHONIUM / BENZOCAINE / MENTHOL|BENZETHONIUM / BENZOCAINE / MENTHOL
C0076660|T121|38260|RXNORM|TIBOLONE|TIBOLONE
C0359018|T121|106963|RXNORM|HYDROCORTISONE / NEOMYCIN|HYDROCORTISONE / NEOMYCIN
C0359018|T121|106963|RXNORM|HYDROCORTISONE / NEOMYCIN|HYDROCORTISONE / NEOMYCIN
C0359019|T121|106964|RXNORM|HYDROCORTISONE / LIDOCAINE|HYDROCORTISONE / LIDOCAINE
C0359019|T121|106964|RXNORM|HYDROCORTISONE / LIDOCAINE|HYDROCORTISONE / LIDOCAINE
C0939225|T121|284629|RXNORM|CARBETAPENTANE / GUAIFENESIN / PHENYLEPHRINE|CARBETAPENTANE / GUAIFENESIN / PHENYLEPHRINE
C2701411|T129|852213|RXNORM|SHEEP SORREL POLLEN EXTRACT|RUMEX ACETOSELLA POLLEN EXTRACT
C0359025|T121|106967|RXNORM|HYDROCORTISONE / MICONAZOLE|HYDROCORTISONE / MICONAZOLE
C3489267|T121|1313308|RXNORM|ALLIUM CEPA WHOLE EXTRACT|ALLIUM CEPA WHOLE EXTRACT
C0051710|T197|1313309|RXNORM|AMMONIUM BROMIDE|AMMONIUM BROMIDE
C3486547|T126|1313304|RXNORM|3-PHYTASE B (ASPERGILLUS NIGER)|3-PHYTASE B (ASPERGILLUS NIGER)
C1880230|T123|1313305|RXNORM|5-HYDROXYTRYPTOPHAN, DL-|5-HYDROXYTRYPTOPHAN, DL-
C0771793|T197|1313302|RXNORM|MANGANESE PHOSPHATE|MANGANESE PHOSPHATE
C3489249|T121|1313303|RXNORM|2,5-PIPERAZINEDIONE|2,5-PIPERAZINEDIONE
C2348752|T121|1372247|RXNORM|GERANIUM EXTRACT|GERANIUM EXTRACT
C2928518|T121|1007600|RXNORM|FOLIC ACID / POLYSACCHARIDE IRON COMPLEX / VITAMIN B 12|FOLIC ACID / POLYSACCHARIDE IRON COMPLEX / VITAMIN B 12
C2928458|T121|1007537|RXNORM|CHONDROITIN SULFATES / GLUCOSAMINE / METHYLSULFONYLMETHANE|CHONDROITIN SULFATES / GLUCOSAMINE / METHYLSULFONYLMETHANE
C2928457|T121|1007536|RXNORM|CRANBERRY PREPARATION / EVENING PRIMROSE OIL|CRANBERRY PREPARATION / EVENING PRIMROSE OIL
C2928456|T121|1007535|RXNORM|HYALURONATE / UREA|HYALURONATE / UREA
C2928455|T121|1007534|RXNORM|MEASLES VIRUS VACCINE LIVE, ENDERS' ATTENUATED EDMONSTON STRAIN / MUMPS VIRUS VACCINE LIVE, JERYL LYNN STRAIN / RUBELLA VIRUS VACCINE LIVE (WISTAR RA 27-3 STRAIN)|MEASLES VIRUS VACCINE LIVE, ENDERS' ATTENUATED EDMONSTON STRAIN / MUMPS VIRUS VACCINE LIVE, JERYL LYNN STRAIN / RUBELLA VIRUS VACCINE LIVE (WISTAR RA 27-3 STRAIN)
C2928454|T121|1007533|RXNORM|ALANINE / ARGININE / CALCIUM CHLORIDE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / SODIUM ACETATE TRIHYDRATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / CALCIUM CHLORIDE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / SODIUM ACETATE TRIHYDRATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2928453|T121|1007532|RXNORM|PETROLATUM / RESORCINOL|PETROLATUM / RESORCINOL
C2928452|T121|1007531|RXNORM|CANNABINOL / TETRAHYDROCANNABINOL|CANNABINOL / TETRAHYDROCANNABINOL
C2006132|T121|1007530|RXNORM|CALCIUM CHLORIDE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM CITRATE|CALCIUM CHLORIDE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM CITRATE
C3667885|T109|1440252|RXNORM|HYDROGENATED AVOCADO OIL|HYDROGENATED AVOCADO OIL
C0353716|T121|103999|RXNORM|METHYLTESTOSTERONE / PEMOLINE / YOHIMBINE|METHYLTESTOSTERONE / PEMOLINE / YOHIMBINE
C3667889|T121|1440257|RXNORM|BENZYL NICOTINAMIDE|BENZYL NICOTINAMIDE
C0071758|T197|34303|RXNORM|POTASSIUM CHROMATE(VI)|POTASSIUM CHROMATE(VI)
C2928460|T121|1007539|RXNORM|BELLADONNA EXTRACT, USP / EPHEDRINE|BELLADONNA EXTRACT, USP / EPHEDRINE
C2928459|T121|1007538|RXNORM|CALCIUM CHLORIDE / GLUCOSE / LACTATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CHLORIDE / GLUCOSE / LACTATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C0995188|T129|318341|RXNORM|CETUXIMAB|CETUXIMAB
C1875485|T121|691137|RXNORM|METHACHOLINE / METHYL SALICYLATE|METHACHOLINE / METHYL SALICYLATE
C0770555|T121|235479|RXNORM|THYROID, PORCINE|THYROID, PORCINE
C0048678|T130|1362740|RXNORM|4-PHENYLENEDIAMINE|4-PHENYLENEDIAMINE
C3859811|T109|1593853|RXNORM|HUMAN SKIN PREPARATION|HUMAN SKIN PREPARATION
C1875487|T121|691138|RXNORM|METHENAMINE / POTASSIUM PHOSPHATE|METHENAMINE / POTASSIUM PHOSPHATE
C1703334|T195|642274|RXNORM|RETAPAMULIN|RETAPAMULIN
C3191910|T121|1146773|RXNORM|MENTHOL / PETROLATUM|MENTHOL / PETROLATUM
C3255840|T109|1309429|RXNORM|WASABI ROOT EXTRACT|WASABI ROOT EXTRACT
C1702615|T121|616546|RXNORM|WHITE KIDNEY BEAN EXTRACT|WHITE KIDNEY BEAN EXTRACT
C0056026|T197|1362742|RXNORM|COBALT SULFATE|COBALT SULFATE
C1095802|T121|319779|RXNORM|ASAFETIDA EXTRACT|FERULA ASSAFOETIDA RESIN EXTRACT
C3256219|T109|1309422|RXNORM|CYMBOPOGON SCHOENANTHUS LEAF EXTRACT|CYMBOPOGON SCHOENANTHUS LEAF EXTRACT
C3256227|T109|1309423|RXNORM|DIOSPYROS KAKI LEAF EXTRACT|DIOSPYROS KAKI LEAF EXTRACT
C3256212|T109|1309420|RXNORM|CUPRESSUS SEMPERVIRENS SEED EXTRACT|CUPRESSUS SEMPERVIRENS SEED EXTRACT
C3256837|T109|1309421|RXNORM|DRYNARIA FORTUNEI ROOT EXTRACT|DRYNARIA FORTUNEI ROOT EXTRACT
C3256684|T121|1309426|RXNORM|GARDENIA TAITENSIS FLOWER EXTRACT|GARDENIA TAITENSIS FLOWER EXTRACT
C3256687|T109|1309427|RXNORM|GENTIANA MACROPHYLLA ROOT EXTRACT|GENTIANA MACROPHYLLA ROOT EXTRACT
C3256619|T109|1309424|RXNORM|FRANKINCENSE OIL|FRANKINCENSE OIL
C3255668|T109|1309425|RXNORM|EPILOBIUM ANGUSTIFOLIUM LEAF EXTRACT|EPILOBIUM ANGUSTIFOLIUM LEAF EXTRACT
C0031406|T121|8130|RXNORM|PHENINDIONE|PHENINDIONE
C2928509|T121|1007591|RXNORM|CHROMIUM PICOLINATE / VITAMIN B6|CHROMIUM PICOLINATE / VITAMIN B6
C0058445|T195|23437|RXNORM|DIRITHROMYCIN|DIRITHROMYCIN
C1601799|T196|486961|RXNORM|PHOSPHATE ION|PHOSPHATE ION
C0982437|T121|314875|RXNORM|TOCOPHERYL ACID SUCCINATE,D-ALPHA|TOCOPHERYL ACID SUCCINATE,D-ALPHA
C1725516|T121|1423272|RXNORM|AMMONIUM XYLENESULFONATE|AMMONIUM XYLENESULFONATE
C0717802|T121|214597|RXNORM|GUAIFENESIN / PHENYLEPHRINE|GUAIFENESIN / PHENYLEPHRINE
C0717801|T121|214596|RXNORM|GUAIFENESIN / OXTRIPHYLLINE|GUAIFENESIN / OXTRIPHYLLINE
C0717799|T121|214594|RXNORM|GUAIFENESIN / HYDROCODONE|GUAIFENESIN / HYDROCODONE
C0304888|T121|91472|RXNORM|SHARK LIVER OIL|SHARK LIVER OIL
C0717804|T121|214599|RXNORM|GUAIFENESIN / PSEUDOEPHEDRINE|GUAIFENESIN / PSEUDOEPHEDRINE
C0717803|T121|214598|RXNORM|GUAIFENESIN / PHENYLPROPANOLAMINE|GUAIFENESIN / PHENYLPROPANOLAMINE
C2701364|T129|852162|RXNORM|BLACK WILLOW POLLEN EXTRACT|BLACK WILLOW POLLEN EXTRACT
C0074754|T197|1366983|RXNORM|SODIUM PEROXIDE|SODIUM PEROXIDE
C1873980|T121|689777|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLPROPANOLAMINE|ACETAMINOPHEN / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLPROPANOLAMINE
C1873979|T121|689776|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE|ACETAMINOPHEN / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE
C2701368|T129|852166|RXNORM|WATER BIRCH POLLEN EXTRACT|BETULA OCCIDENTALIS POLLEN EXTRACT
C3255600|T121|1311601|RXNORM|HEDERA HELIX TOP EXTRACT|HEDERA HELIX TOP EXTRACT
C0056784|T121|1366989|RXNORM|GAMMA-CYCLODEXTRIN|GAMMA-CYCLODEXTRIN
C1873982|T121|689779|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / PHENYLEPHRINE / PYRILAMINE|ACETAMINOPHEN / DEXTROMETHORPHAN / PHENYLEPHRINE / PYRILAMINE
C1873981|T121|689778|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE|ACETAMINOPHEN / DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE
C1955474|T129|733003|RXNORM|PLERIXAFOR|PLERIXAFOR
C0032153|T204|1432989|RXNORM|PLASMODIUM MALARIAE|PLASMODIUM MALARIAE
C1302069|T121|392520|RXNORM|METRONIDAZOLE / NYSTATIN|METRONIDAZOLE / NYSTATIN
C2928511|T121|1007593|RXNORM|DEHYDROCHOLATE / PAPAVERINE|DEHYDROCHOLATE / PAPAVERINE
C0085542|T121|42463|RXNORM|PRAVASTATIN|PRAVASTATIN
C1337310|T109|1370470|RXNORM|CLARY SAGE EXTRACT|CLARY SAGE EXTRACT
C1302104|T121|687315|RXNORM|DOMIPHEN / LIDOCAINE|DOMIPHEN / LIDOCAINE
C3643654|T121|1422066|RXNORM|N-ALKYL ETHYLBENZYL DIMETHYL AMMONIUM (C12-C14)|N-ALKYL ETHYLBENZYL DIMETHYL AMMONIUM (C12-C14)
C0022499|T197|6102|RXNORM|KAOLIN|KAOLIN
C3864823|T109|1597389|RXNORM|QUATERNIUM-33|QUATERNIUM-33
C0041411|T130|10938|RXNORM|TURPENTINE|TURPENTINE
C0139007|T121|55244|RXNORM|PROTHIPENDYL|PROTHIPENDYL
C3832941|T121|1539965|RXNORM|ANGELICA DAHURICA VAR. FORMOSANA WHOLE EXTRACT|ANGELICA DAHURICA VAR. FORMOSANA WHOLE EXTRACT
C2928513|T121|1007595|RXNORM|LANOLIN / PETROLATUM / ZINC OXIDE|LANOLIN / PETROLATUM / ZINC OXIDE
C2929895|T121|1009000|RXNORM|TRETINOIN / UREA|TRETINOIN / UREA
C3464190|T121|1291430|RXNORM|DOCOSAENOIC ACID / EICOSAPENTAENOATE|DOCOSAENOIC ACID / EICOSAPENTAENOATE
C0771958|T129|236658|RXNORM|BOTULISM ANTITOXIN A|BOTULISM ANTITOXIN A
C0637887|T197|1337969|RXNORM|ANTIMONY PENTASULFIDE|ANTIMONY PENTASULFIDE
C0771792|T121|236512|RXNORM|AMINOHYDROXYBUTYRIC ACID|AMINOHYDROXYBUTYRIC ACID
C0937932|T126|283821|RXNORM|RASBURICASE|RASBURICASE
C2730227|T129|892616|RXNORM|EGG WHITE (CHICKEN) ALLERGENIC EXTRACT|EGG WHITE (CHICKEN) ALLERGENIC EXTRACT
C0937941|T121|283829|RXNORM|CIDER VINEGAR|CIDER VINEGAR
C2075280|T121|818449|RXNORM|CISAPRIDE / SIMETHICONE|CISAPRIDE / SIMETHICONE
C1874973|T121|690467|RXNORM|DEXCHLORPHENIRAMINE / GUAIFENESIN / PSEUDOEPHEDRINE|DEXCHLORPHENIRAMINE / GUAIFENESIN / PSEUDOEPHEDRINE
C1874972|T121|690466|RXNORM|DEXCHLORPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|DEXCHLORPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C0357131|T121|105695|RXNORM|EPOETIN BETA|EPOETIN BETA
C0357126|T121|105694|RXNORM|EPOETIN ALFA|EPOETIN ALFA
C0772197|T121|236872|RXNORM|CHLOROTHEOPHYLLINE|CHLOROTHEOPHYLLINE
C0718909|T121|215648|RXNORM|COMPOUND BENZOIN TINCTURE (USP)|COMPOUND BENZOIN TINCTURE (USP)
C0116569|T121|49737|RXNORM|ESMOLOL|ESMOLOL
C2350948|T121|1300701|RXNORM|LORCASERIN|LORCASERIN
C0038481|T131|1310185|RXNORM|STRYCHNINE NITRATE|STRYCHNINE NITRATE
C0012289|T121|3416|RXNORM|DIHYDROERGOCRISTINE|DIHYDROERGOCRISTINE
C0012290|T121|3417|RXNORM|DIHYDROERGOCRYPTINE|DIHYDROERGOCRYPTINE
C0012288|T121|3415|RXNORM|DIHYDROERGOCORNINE|DIHYDROERGOCORNINE
C0056039|T127|21373|RXNORM|COBAMAMIDE|COBAMAMIDE
C3666922|T121|1437983|RXNORM|HYPROMELLOSE 2910 (10000 MPA.S)|HYPROMELLOSE 2910 (10000 MPA.S)
C3666924|T121|1437985|RXNORM|CITRUS SINENSIS WHOLE EXTRACT|CITRUS SINENSIS WHOLE EXTRACT
C3666923|T121|1437984|RXNORM|BENZORESORCINOL|BENZORESORCINOL
C0012291|T121|3418|RXNORM|DIHYDROERGOTAMINE|DIHYDROERGOTAMINE
C2348063|T130|1437986|RXNORM|D&C RED NO. 34|D&C RED NO. 34
C1530072|T121|1086769|RXNORM|VILAZODONE|VILAZODONE
C2940008|T121|1014426|RXNORM|ALANINE / ARGININE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / PROLINE / SERINE / SODIUM BISULFITE / THREONINE / TRYPTOPHAN / VALINE|ALANINE / ARGININE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / PROLINE / SERINE / SODIUM BISULFITE / THREONINE / TRYPTOPHAN / VALINE
C3160115|T121|1112496|RXNORM|SAW PALMETTO EXTRACT / ZINC PICOLINATE|SAW PALMETTO EXTRACT / ZINC PICOLINATE
C2929861|T121|1008965|RXNORM|ATROPINE / BENZOATE / HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / PHENYL SALICYLATE|ATROPINE / BENZOATE / HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / PHENYL SALICYLATE
C2929860|T121|1008964|RXNORM|KAVA PREPARATION / PASSION FLOWER EXTRACT / VALERIAN ROOT EXTRACT|KAVA PREPARATION / PASSION FLOWER EXTRACT / VALERIAN ROOT EXTRACT
C2929863|T121|1008967|RXNORM|DIPTHERIA PROTEIN / HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE|DIPTHERIA PROTEIN / HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE
C2929862|T121|1008966|RXNORM|BENZOYL PEROXIDE / COLLOID SULFUR|BENZOYL PEROXIDE / COLLOID SULFUR
C2929857|T121|1008961|RXNORM|BACITRACIN / LIDOCAINE / NEOMYCIN|BACITRACIN / LIDOCAINE / NEOMYCIN
C2929856|T121|1008960|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / SCOPOLAMINE|CHLORPHENIRAMINE / DEXTROMETHORPHAN / SCOPOLAMINE
C2929859|T121|1008963|RXNORM|ASCORBIC ACID / POLYSACCHARIDE IRON COMPLEX|ASCORBIC ACID / POLYSACCHARIDE IRON COMPLEX
C2929858|T121|1008962|RXNORM|ISOTHIPENDYL / PIPAZETHATE|ISOTHIPENDYL / PIPAZETHATE
C0006976|T195|2015|RXNORM|CARBENICILLIN|CARBENICILLIN
C3859935|T109|1594338|RXNORM|PIPERAZINE, 1-(4'-METHOXY(1,1'-BIPHENYL)-2-YL)-|PIPERAZINE, 1-(4'-METHOXY(1,1'-BIPHENYL)-2-YL)-
C2929865|T121|1008969|RXNORM|ALGINIC ACID / ALUMINUM HYDROXIDE / MAGNESIUM CARBONATE|ALGINIC ACID / ALUMINUM HYDROXIDE / MAGNESIUM CARBONATE
C2929864|T121|1008968|RXNORM|BENZETHONIUM / DYCLONINE|BENZETHONIUM / DYCLONINE
C3488450|T121|1313973|RXNORM|VISCUM ALBUM WHOLE EXTRACT|VISCUM ALBUM WHOLE EXTRACT
C3497931|T121|1311367|RXNORM|SUS SCROFA KNEE JOINT PREPARATION|PORCINE KNEE JOINT PREPARATION
C2929539|T121|1008639|RXNORM|NAPHAZOLINE / POLYETHYLENE GLYCOL 300|NAPHAZOLINE / POLYETHYLENE GLYCOL 300
C3486673|T129|1313972|RXNORM|MUCOR RACEMOSUS IMMUNOSERUM RABBIT|MUCOR RACEMOSUS IMMUNOSERUM RABBIT
C2929535|T121|1008635|RXNORM|DEXTROMETHORPHAN / DOXYLAMINE / PHENYLEPHRINE|DEXTROMETHORPHAN / DOXYLAMINE / PHENYLEPHRINE
C2929534|T121|1008634|RXNORM|LUTEIN / ZEAXANTHIN|LUTEIN / ZEAXANTHIN
C2929537|T121|1008637|RXNORM|PHOSPHOLIPIDS / PROTEINS|PHOSPHOLIPIDS / PROTEINS
C2929536|T121|1008636|RXNORM|FOLIC ACID / PYRIDOXINE / VITAMIN B 12|FOLIC ACID / PYRIDOXINE / VITAMIN B 12
C2929531|T121|1008631|RXNORM|ASCORBIC ACID / CALCIUM CARBONATE / FERROUS FUMARATE / FOLIC ACID|ASCORBIC ACID / CALCIUM CARBONATE / FERROUS FUMARATE / FOLIC ACID
C2929530|T121|1008630|RXNORM|EUCALYPTOL / GUAIACOL ETHYLGLYCOLATE|EUCALYPTOL / GUAIACOL ETHYLGLYCOLATE
C1714033|T121|637366|RXNORM|WHEAT DEXTRIN|WHEAT DEXTRIN
C3834057|T109|1543079|RXNORM|ETHYL 10-UNDECENOATE|ETHYL 10-UNDECENOATE
C3834058|T109|1543078|RXNORM|METHYL UNDECYLENATE|METHYL UNDECYLENATE
C0075209|T121|1313977|RXNORM|STEARAMINE|STEARAMINE
C3834059|T121|1543077|RXNORM|EUPHORBIA HIRTA FLOWERING TOP EXTRACT|EUPHORBIA HIRTA FLOWERING TOP EXTRACT
C0305062|T129|798306|RXNORM|TETANUS TOXOID VACCINE, INACTIVATED|CLOSTRIDIUM TETANI TOXOID ANTIGEN, INACTIVATED
C0071545|T121|1363053|RXNORM|POLYDEXTROSE|POLYDEXTROSE
C0067912|T109|1363052|RXNORM|N-DECYL ALCOHOL|1-DECANOL
C0066776|T121|1363051|RXNORM|MONOPHOSPHORYL LIPID A|MONOPHOSPHORYL LIPID A
C0065601|T121|1363050|RXNORM|MALTODEXTRIN|MALTODEXTRIN
C0074915|T121|1363057|RXNORM|SORBITAN MONOSTEARATE|SORBITAN MONOSTEARATE
C0074913|T122|1363056|RXNORM|SORBITAN MONOOLEATE|SORBITAN MONOOLEATE
C0074912|T121|1363055|RXNORM|SORBITAN MONOLAURATE|SORBITAN MONOLAURATE
C0073970|T109|1363054|RXNORM|SALICYL ALCOHOL|SALICYL ALCOHOL
C0075159|T197|1363059|RXNORM|STANNIC OXIDE|STANNIC OXIDE
C0074916|T121|1363058|RXNORM|SORBITAN SESQUIOLEATE|SORBITAN SESQUIOLEATE
C0039419|T197|1423270|RXNORM|TECHNETIUM TC 99M SULFUR COLLOID|TECHNETIUM (99MTC) SULFUR COLLOID
C0040193|T195|10591|RXNORM|TICARCILLIN|TICARCILLIN
C0040219|T121|10597|RXNORM|TILIDINE|TILIDINE
C0040207|T121|10594|RXNORM|TICLOPIDINE|TICLOPIDINE
C3486596|T121|1310024|RXNORM|COMOCLADIA DENTATA BARK-LEAF EXTRACT|COMOCLADIA DENTATA BARK-LEAF EXTRACT
C3489345|T121|1310025|RXNORM|CASTANEA SATIVE LEAF EXTRACT|CASTANEA SATIVE LEAF EXTRACT
C3538038|T122|1371910|RXNORM|IPOMOEA PURPUREA SEED EXTRACT|IPOMOEA PURPUREA SEED EXTRACT
C3267301|T121|1310021|RXNORM|CRATAEGUS MONOGYNA FLOWER EXTRACT|CRATAEGUS MONOGYNA FLOWER EXTRACT
C3473231|T121|1310022|RXNORM|STYPHNOLOBIUM JAPONICUM ROOT EXTRACT|STYPHNOLOBIUM JAPONICUM ROOT EXTRACT
C3489112|T121|1310023|RXNORM|CYNANCHUM VINCETOXICUM LEAF EXTRACT|CYNANCHUM VINCETOXICUM LEAF EXTRACT
C3488090|T121|1311269|RXNORM|SUS SCROFA RENAL PELVIS PREPARATION|PORCINE RENAL PELVIS PREPARATION
C3486563|T121|1311268|RXNORM|SUS SCROFA COLON PREPARATION|PORCINE COLON PREPARATION
C3255875|T109|1313978|RXNORM|STEARYL BEHENATE|STEARYL BEHENATE
C2722042|T129|973274|RXNORM|OYSTER ALLERGENIC EXTRACT|OYSTER ALLERGENIC EXTRACT
C0024658|T121|1311261|RXNORM|MALTOSE|MALTOSE
C2928416|T121|1007494|RXNORM|COBALAMINS / VITAMIN B 12|COBALAMINS / VITAMIN B 12
C3486842|T121|1311262|RXNORM|SUS SCROFA TENDON PREPARATION|PORCINE TENDON PREPARATION
C2608748|T121|1311265|RXNORM|LYTTA VESICATORIA PREPARATION|CANTHARIS PREPARATION
C3496034|T121|1311264|RXNORM|SUS SCROFA TONSIL PREPARATION|PORCINE TONSIL PREPARATION
C3486549|T121|1311266|RXNORM|SUS SCROFA VAGUS NERVE PREPARATION|PORCINE VAGUS NERVE PREPARATION
C0054840|T121|20355|RXNORM|CARZENIDE|CARZENIDE
C2746264|T129|902215|RXNORM|COMMON COCKLEBUR POLLEN EXTRACT|XANTHIUM STRUMARIUM VAR. CANADENSE POLLEN EXTRACT
C0054836|T121|20352|RXNORM|CARVEDILOL|CARVEDILOL
C0076448|T121|38077|RXNORM|THIOBUTABARBITAL|THIOBUTABARBITAL
C3255958|T121|1424909|RXNORM|MARRUBIUM VULGARE EXTRACT|COMMON HOREHOUND EXTRACT
C3473402|T109|1307939|RXNORM|LITSEA OIL|LITSEA OIL
C0063384|T121|27438|RXNORM|IMIDAZOLE-2-HYDROXYBENZOATE|IMIDAZOLE SALICYLATE
C1814271|T130|1306061|RXNORM|TETRAKIS(1-ISOCYANO-2-METHOXY-2-METHYL-PROPANE)-COPPER(I) TETRAFLUOROBORATE|TETRAKIS(1-ISOCYANO-2-METHOXY-2-METHYL-PROPANE)-COPPER(I) TETRAFLUOROBORATE
C0072511|T121|34906|RXNORM|PROXYPHYLLINE|PROXYPHYLLINE
C0072510|T121|34905|RXNORM|PROPARACAINE|PROPARACAINE
C3484416|T121|1310248|RXNORM|BERBERIS VULGARIS FRUIT EXTRACT|BERBERIS VULGARIS FRUIT EXTRACT
C3488934|T121|1310249|RXNORM|BOS TAURUS BILE PREPARATION|BOVINE BILE PREPARATION
C1689936|T121|608362|RXNORM|ICHTHAMMOL / ZINC OXIDE|ICHTHAMMOL / ZINC OXIDE
C3190778|T121|1145109|RXNORM|AZELATE / CUPRIC OXIDE / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / ZINC OXIDE|AZELATE / CUPRIC OXIDE / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / ZINC OXIDE
C0078956|T126|40028|RXNORM|ANISTREPLASE|ANISTREPLASE
C3486683|T121|1310244|RXNORM|BOS TAURUS ADRENAL GLAND PREPARATION|BOVINE ADRENAL GLAND PREPARATION
C0145106|T195|57021|RXNORM|TEICOPLANIN|TEICOPLANIN
C3495980|T121|1310246|RXNORM|BOS TAURUS ANKLE JOINT PREPARATION|BOVINE ANKLE JOINT PREPARATION
C1876822|T121|700809|RXNORM|DEXBROMPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE|DEXBROMPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE
C3152932|T121|1098361|RXNORM|NAPHAZOLINE / POLYSORBATE 80|NAPHAZOLINE / POLYSORBATE 80
C2700605|T196|1546418|RXNORM|CHROMIC CATION|CHROMIC CATION
C2928625|T121|1007709|RXNORM|BENZOCAINE / CHLORHEXIDINE|BENZOCAINE / CHLORHEXIDINE
C2928620|T121|1007704|RXNORM|ACETAMINOPHEN / SALICYLIC ACID|ACETAMINOPHEN / SALICYLIC ACID
C2928621|T121|1007705|RXNORM|ALUMINUM MAGNESIUM SILICATE / CALCIUM CARBONATE|ALUMINUM MAGNESIUM SILICATE / CALCIUM CARBONATE
C2928622|T121|1007706|RXNORM|ACETAMINOPHEN / DIHYDROERGOTAMINE|ACETAMINOPHEN / DIHYDROERGOTAMINE
C2928623|T121|1007707|RXNORM|ACONITE / LACTOSE|ACONITE / LACTOSE
C2928616|T121|1007700|RXNORM|FLUOCORTOLONE / LIDOCAINE|FLUOCORTOLONE / LIDOCAINE
C3205070|T121|1150100|RXNORM|BIFIDOBACTERIUM LACTIS / BIFIDOBACTERIUM LONGUM / LACTOBACILLUS ACIDOPHILUS|BIFIDOBACTERIUM LACTIS / BIFIDOBACTERIUM LONGUM / LACTOBACILLUS ACIDOPHILUS
C2928618|T121|1007702|RXNORM|ACEPROMETAZINE / MEPROBAMATE|ACEPROMETAZINE / MEPROBAMATE
C2928619|T121|1007703|RXNORM|CLONIXIN / PROPINOX|CLONIXIN / PROPINOX
C0719818|T121|216524|RXNORM|DEXAMETHASONE / NEOMYCIN|DEXAMETHASONE / NEOMYCIN
C0719818|T121|216524|RXNORM|DEXAMETHASONE / NEOMYCIN|DEXAMETHASONE / NEOMYCIN
C0719819|T121|216525|RXNORM|DEXAMETHASONE / NEOMYCIN / POLYMYXIN B|DEXAMETHASONE / NEOMYCIN / POLYMYXIN B
C1874210|T121|691307|RXNORM|AMMONIUM CHLORIDE / IPECAC|AMMONIUM CHLORIDE / IPECAC
C0064044|T109|1364275|RXNORM|ISOPRENE|ISOPRENE
C1739462|T126|644101|RXNORM|IDURSULFASE|IDURSULFASE
C0937772|T121|283680|RXNORM|GOLDEN SEAL ROOT EXTRACT|GOLDEN SEAL ROOT EXTRACT
C0304096|T109|1426919|RXNORM|BAY OIL (PIMENTA RACEMOSA)|BAY OIL (PIMENTA RACEMOSA)
C0065605|T121|1362894|RXNORM|MALTOL|MALTOL
C0065654|T123|1362895|RXNORM|MANGIFERIN|MANGIFERIN
C0066503|T197|1362896|RXNORM|MICA|MICA
C0067074|T121|1362897|RXNORM|MYRISTYL ALCOHOL|MYRISTYL ALCOHOL
C0055809|T121|1362890|RXNORM|CITRAL|CITRAL
C2728186|T129|1010932|RXNORM|LEEK ALLERGENIC EXTRACT|LEEK ALLERGENIC EXTRACT
C0059788|T121|1362892|RXNORM|ETHYL-P-HYDROXYBENZOATE|ETHYL-P-HYDROXYBENZOATE
C0063124|T109|1362893|RXNORM|HYDROXYCITRONELLAL|HYDROXYCITRONELLAL
C0071639|T121|1362898|RXNORM|POLYOXYETHYLENE-24-CHOLESTERYL ETHER|POLYOXYETHYLENE-24-CHOLESTERYL ETHER
C0071771|T197|1362899|RXNORM|POTASSIUM METABISULFITE|POTASSIUM METABISULFITE
C3710066|T109|1488998|RXNORM|ACACIA DEALBATA FLOWER EXTRACT|ACACIA DEALBATA FLOWER EXTRACT
C3710067|T109|1488999|RXNORM|BOERHAVIA DIFFUSA ROOT EXTRACT|BOERHAVIA DIFFUSA ROOT EXTRACT
C3709488|T121|1487529|RXNORM|CETYL BEHENATE|CETYL BEHENATE
C0004886|T129|1344|RXNORM|BCG VACCINE|BCG VACCINE
C0004905|T125|1347|RXNORM|BECLOMETHASONE|BECLOMETHASONE
C0004905|T125|1347|RXNORM|BECLOMETHASONE|BECLOMETHASONE
C3556191|T121|1373721|RXNORM|3-O-ETHYL ASCORBATE|3-O-ETHYL ASCORBATE
C3555532|T121|1373722|RXNORM|CITRUS SINENSIS FLOWER EXTRACT|CITRUS SINENSIS FLOWER EXTRACT
C3555531|T121|1373723|RXNORM|GOSSYPIUM HERBACEUM WHOLE EXTRACT|GOSSYPIUM HERBACEUM WHOLE EXTRACT
C3555530|T121|1373724|RXNORM|METHYL 3-HYDROXYBENZOATE|METHYL 3-HYDROXYBENZOATE
C3555529|T121|1373725|RXNORM|PEG-PPG-17-18 DIMETHICONE|PEG-PPG-17-18 DIMETHICONE
C3555528|T121|1373726|RXNORM|POLYGLYCERYL-3 RICINOLEATE|POLYGLYCERYL-3 RICINOLEATE
C2354879|T121|1373727|RXNORM|RETINYL RETINOATE|RETINYL RETINOATE
C3555527|T121|1373728|RXNORM|ROSA CANINA SEED EXTRACT|ROSA CANINA SEED EXTRACT
C0031364|T131|8113|RXNORM|PHENACETIN|PHENACETIN
C0025893|T195|6927|RXNORM|MEZLOCILLIN|MEZLOCILLIN
C0025887|T121|6926|RXNORM|MEXILETINE|MEXILETINE
C0025869|T130|6920|RXNORM|METRIZAMIDE|METRIZAMIDE
C0025876|T125|6923|RXNORM|METYRAPONE|METYRAPONE
C0025872|T121|6922|RXNORM|METRONIDAZOLE|METRONIDAZOLE
C0025872|T121|6922|RXNORM|METRONIDAZOLE|METRONIDAZOLE
C0025872|T121|6922|RXNORM|METRONIDAZOLE|METRONIDAZOLE
C0025872|T121|6922|RXNORM|METRONIDAZOLE|METRONIDAZOLE
C0025872|T121|6922|RXNORM|METRONIDAZOLE|METRONIDAZOLE
C0062525|T129|26744|RXNORM|HEPATITIS B IMMUNE GLOBULIN|HEPATITIS B IMMUNOGLOBIN
C0029300|T123|7712|RXNORM|OROTIC ACID|OROTIC ACID
C0029309|T121|7715|RXNORM|ORPHENADRINE|ORPHENADRINE
C3247810|T121|1193036|RXNORM|CHOLECALCIFEROL / FOLIC ACID / OMEGA-3 ACID ETHYL ESTERS (USP) / PHYTOSTEROLS / PYRIDOXINE / VITAMIN B 12|CHOLECALCIFEROL / FOLIC ACID / OMEGA-3 ACID ETHYL ESTERS (USP) / PHYTOSTEROLS / PYRIDOXINE / VITAMIN B 12
C0982338|T121|314784|RXNORM|YELLOW PHENOLPHTHALEIN|YELLOW PHENOLPHTHALEIN
C3819168|T121|1492302|RXNORM|HYDROXYPROPYL BIS-HYDROXYETHYLDIMONIUM|HYDROXYPROPYL BIS-HYDROXYETHYLDIMONIUM
C1434556|T121|1421444|RXNORM|ETILEVODOPA|ETILEVODOPA
C2356037|T130|802624|RXNORM|GADOXETATE|GADOXETATE
C3484548|T121|1311044|RXNORM|EPIMEDIUM GRANDIFLORUM TOP EXTRACT|EPIMEDIUM GRANDIFLORUM TOP EXTRACT
C3489192|T121|1311047|RXNORM|IMMATURE JUGLANS REGIA FRUIT RIND EXTRACT|IMMATURE JUGLANS REGIA FRUIT RIND EXTRACT
C3484575|T121|1311041|RXNORM|CALVATIA GIGANTEA EXTRACT|CALVATIA GIGANTEA EXTRACT
C3484401|T121|1311040|RXNORM|BROWN RICE PREPARATION|BROWN RICE PREPARATION
C3256914|T109|1426645|RXNORM|GUAVA EXTRACT|GUAVA EXTRACT
C2917628|T121|992917|RXNORM|BAPTISIA TINCTORIA EXTRACT|BAPTISIA TINCTORIA EXTRACT
C3256806|T109|1426646|RXNORM|SILICA DIMETHYL SILYLATE|SILICA DIMETHYL SILYLATE
C3486219|T121|1312537|RXNORM|ALPHA-AMYLCINNAMYL ALCOHOL|ALPHA-AMYLCINNAMYL ALCOHOL
C0717904|T121|214691|RXNORM|MANNITOL / SORBITOL|MANNITOL / SORBITOL
C3488920|T109|1309351|RXNORM|MAGNOLIA OFFICINALIS FLOWER EXTRACT|MAGNOLIA OFFICINALIS FLOWER EXTRACT
C0005642|T196|1599|RXNORM|BISMUTH|BISMUTH
C0053508|T121|1312538|RXNORM|BETA-THUJAPLICIN|BETA-THUJAPLICIN
C0717912|T121|214699|RXNORM|MEPERIDINE / PROMETHAZINE|MEPERIDINE / PROMETHAZINE
C0873033|T121|259372|RXNORM|FRUCTOOLIGOSACCHARIDE|FRUCTOOLIGOSACCHARIDE
C3256879|T121|1425403|RXNORM|YUCCA SCHIDIGERA EXTRACT|YUCCA SCHIDIGERA EXTRACT
C1703327|T121|1425406|RXNORM|MYRISTYL NICOTINATE|MYRISTYL NICOTINATE
C0633017|T121|1425405|RXNORM|N-VALYLTRYPTOPHAN|N-VALYLTRYPTOPHAN
C3256812|T121|1425404|RXNORM|VERBENA OFFICINALIS EXTRACT|VERBENA OFFICINALIS EXTRACT
C2587184|T121|831503|RXNORM|FIBRINOGEN CONCENTRATE (HUMAN)|FIBRINOGEN CONCENTRATE (HUMAN)
C3710065|T109|1488997|RXNORM|LAWSONIA INERMIS FLOWERING TOP EXTRACT|LAWSONIA INERMIS FLOWERING TOP EXTRACT
C1276807|T121|389132|RXNORM|BUDESONIDE / FORMOTEROL|BUDESONIDE / FORMOTEROL
C2731877|T129|896213|RXNORM|COMMON WORMWOOD POLLEN EXTRACT|ARTEMISIA ANNUA POLLEN EXTRACT
C0118092|T121|50138|RXNORM|FONAZINE|DIMETOTIAZINE
C3695962|T121|1484280|RXNORM|ZEA MAYS SUBSP. MAYS WHOLE EXTRACT|ZEA MAYS SUBSP. MAYS WHOLE EXTRACT
C1210517|T007|1544936|RXNORM|BARTONELLA WASHOENSIS|BARTONELLA WASHOENSIS
C3695961|T122|1484281|RXNORM|ISOPROPYLPHTHALIMIDE|ISOPROPYLPHTHALIMIDE
C3535913|T121|1368646|RXNORM|FOSCOLATE|FOSCOLATE
C3500587|T109|1314847|RXNORM|TOXICODENDRON VERNICIFLUUM FRUIT RIND WAX|TOXICODENDRON VERNICIFLUUM FRUIT RIND WAX
C3644625|T109|1425356|RXNORM|SALVIA SCLAREA SEED OIL|SALVIA SCLAREA SEED OIL
C0717670|T121|214470|RXNORM|DENILEUKIN DIFTITOX|DENILEUKIN DIFTITOX
C0717671|T121|214471|RXNORM|DESERPIDINE / HYDROCHLOROTHIAZIDE|DESERPIDINE / HYDROCHLOROTHIAZIDE
C0717672|T121|214472|RXNORM|DESERPIDINE / METHYCLOTHIAZIDE|DESERPIDINE / METHYCLOTHIAZIDE
C0717678|T121|214478|RXNORM|DEXAMETHASONE / LIDOCAINE|DEXAMETHASONE / LIDOCAINE
C1565750|T121|593411|RXNORM|SITAGLIPTIN|SITAGLIPTIN
C0028277|T121|7500|RXNORM|NOMIFENSINE|NOMIFENSINE
C0073083|T131|35380|RXNORM|RESMETHRIN|RESMETHRIN
C0304977|T197|91531|RXNORM|SODIUM IODIDE I123|SODIUM IODIDE (123I)
C2701653|T129|852577|RXNORM|ENGLISH WALNUT POLLEN EXTRACT|JUGLANS REGIA POLLEN EXTRACT
C2929296|T121|1008392|RXNORM|CARBON DIOXIDE / NITROGEN / OXYGEN|CARBON DIOXIDE / NITROGEN / OXYGEN
C2929297|T121|1008393|RXNORM|DEXCHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE|DEXCHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE
C2929294|T121|1008390|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED, A-H1N1 (A-BRISBANE-59-2007) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED, A-H3N2 (A-URUGUAY-716-2007) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED, INFLUENZA B (B-FLORIDA-4-2006) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED, A-H1N1 (A-BRISBANE-59-2007) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED, A-H3N2 (A-URUGUAY-716-2007) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED, INFLUENZA B (B-FLORIDA-4-2006) STRAIN
C2929295|T121|1008391|RXNORM|CARBON MONOXIDE / NEON / NITROGEN / OXYGEN|CARBON MONOXIDE / NEON / NITROGEN / OXYGEN
C2929301|T121|1008397|RXNORM|CHROMIUM CITRATE / MANGANESE CITRATE / VANADIUM|CHROMIUM CITRATE / MANGANESE CITRATE / VANADIUM
C2929299|T121|1008395|RXNORM|MENINGOCOCCAL GROUP A POLYSACCHARIDE / MENINGOCOCCAL GROUP C POLYSACCHARIDE / MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP W-135 / MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP Y|MENINGOCOCCAL GROUP A POLYSACCHARIDE / MENINGOCOCCAL GROUP C POLYSACCHARIDE / MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP W-135 / MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP Y
C2929302|T121|1008398|RXNORM|MECHLORETHAMINE / TERPIN HYDRATE|MECHLORETHAMINE / TERPIN HYDRATE
C2929303|T121|1008399|RXNORM|CLOTRIMAZOLE / HEXAMIDINE|CLOTRIMAZOLE / HEXAMIDINE
C0046519|T121|13714|RXNORM|ENSULIZOLE|PHENYLBENZIMIDAZOLE SULFONIC ACID
C0546173|T127|142407|RXNORM|CALCIUM ASCORBATE|CALCIUM ASCORBATE
C0057258|T121|22396|RXNORM|DEFLAZACORT|DEFLAZACORT
C0009185|T130|2660|RXNORM|FLOR DE PIEDRA|COCCIDIOIDIN
C0024321|T125|6529|RXNORM|LYNESTRENOL|LYNESTRENOL
C0013030|T123|3628|RXNORM|DOPAMINE|DOPAMINE
C1875441|T121|690895|RXNORM|LIDOCAINE / SODIUM CHLORIDE|LIDOCAINE / SODIUM CHLORIDE
C1875440|T121|690893|RXNORM|LIDOCAINE / POVIDONE-IODINE|LIDOCAINE / POVIDONE-IODINE
C0013015|T121|3626|RXNORM|DOMPERIDONE|DOMPERIDONE
C3644996|T109|1426261|RXNORM|JASMINE LACTONE|JASMINE LACTONE
C2701494|T129|852311|RXNORM|WHEAT RUST EXTRACT|PUCCINIA STRIIFORMIS VAR. STRIIFORMIS EXTRACT
C3474159|T121|1307679|RXNORM|CHILEAN HAZELNUT OIL|CHILEAN HAZELNUT OIL
C2701498|T129|852315|RXNORM|KAPOK TREE FIBER EXTRACT|CEIBA PENTANDRA FIBER EXTRACT
C3256346|T121|1307678|RXNORM|BAMBUSA VULGARIS WHOLE EXTRACT|BAMBUSA VULGARIS WHOLE EXTRACT
C3848566|T196|1546281|RXNORM|INDIUM CATION IN-111|INDIUM CATION IN-111
C2940372|T121|1020419|RXNORM|CAPSAICIN / LIDOCAINE / MENTHOL / METHYL SALICYLATE|CAPSAICIN / LIDOCAINE / MENTHOL / METHYL SALICYLATE
C0043474|T121|11413|RXNORM|ZIDOVUDINE|ZIDOVUDINE
C1533391|T116|477454|RXNORM|COLLAGEN, HYDROLYZED|COLLAGEN, HYDROLYZED
C0795589|T196|253158|RXNORM|UREA [14C]|UREA [14C]
C0043481|T196|11416|RXNORM|ZINC|ZINC
C0795592|T121|253159|RXNORM|CHROMIUM ASPARTATE|CHROMIUM ASPARTATE
C3472713|T109|1307705|RXNORM|PELARGONIUM GRAVEOLENS FLOWER OIL|PELARGONIUM GRAVEOLENS FLOWER OIL
C3256050|T121|1307704|RXNORM|HYPERICUM PERFORATUM LEAF EXTRACT|HYPERICUM PERFORATUM LEAF EXTRACT
C3256677|T121|1307707|RXNORM|FLICKINGERIA FIMBRIATA STEM EXTRACT|FLICKINGERIA FIMBRIATA STEM EXTRACT
C3255610|T121|1307706|RXNORM|PUNICA GRANATUM FLOWER EXTRACT|PUNICA GRANATUM FLOWER EXTRACT
C3257421|T121|1307701|RXNORM|YUCCA SCHIDIGERA ROOT EXTRACT|YUCCA SCHIDIGERA ROOT EXTRACT
C3255963|T121|1307700|RXNORM|PEG-10 RAPESEED STEROL|PEG-10 RAPESEED STEROL
C3475282|T109|1307703|RXNORM|PERILLA FRUTESCENS SEED OIL|PERILLA FRUTESCENS SEED OIL
C3256587|T121|1307674|RXNORM|ACTINIDIA POLYGAMA FRUIT EXTRACT|ACTINIDIA POLYGAMA FRUIT EXTRACT
C2726218|T129|968506|RXNORM|SYNCEPHALASTRUM RACEMOSUM ALLERGENIC EXTRACT|SYNCEPHALASTRUM RACEMOSUM ALLERGENIC EXTRACT
C0081609|T197|1316091|RXNORM|ANTIMONY TRISULFIDE|ANTIMONY TRISULFIDE
C3256516|T121|1307709|RXNORM|DIPTERYX ODORATA SEED EXTRACT|DIPTERYX ODORATA SEED EXTRACT
C3256183|T168|1307708|RXNORM|RICE GERM OIL|RICE GERM OIL
C3848564|T196|1546284|RXNORM|BISMUTH CATION|BISMUTH CATION
C3256430|T121|1307671|RXNORM|PINUS TABULIFORMIS BARK EXTRACT|PINUS TABULIFORMIS BARK EXTRACT
C0752345|T122|1424910|RXNORM|HIGH-DENSITY POLYETHYLENE|HIGH-DENSITY POLYETHYLENE
C3467876|T121|1424911|RXNORM|DABRAFENIB|DABRAFENIB
C0077410|T127|38893|RXNORM|TROXERUTIN|TROXERUTIN
C3256247|T121|1307670|RXNORM|PERSICARIA TINCTORIA LEAF EXTRACT|PERSICARIA TINCTORIA LEAF EXTRACT
C0046100|T121|13369|RXNORM|OCTINOXATE|OCTINOXATE
C0579233|T007|1363918|RXNORM|STREPTOCOCCUS AGALACTIAE|STREPTOCOCCUS AGALACTIAE
C0318157|T007|1363919|RXNORM|STREPTOCOCCUS VIRIDANS GROUP|STREPTOCOCCUS VIRIDANS GROUP
C0010467|T130|2955|RXNORM|CURCUMIN|CURCUMIN
C0006464|T121|477631|RXNORM|BUTABARBITAL|BUTABARBITAL
C3503768|T121|1363916|RXNORM|CARMOISINE|CARMOISINE
C0038410|T007|1363917|RXNORM|STREPTOCOCCUS PNEUMONIAE|STREPTOCOCCUS PNEUMONIAE
C0000294|T121|44|RXNORM|FLUORIDES|MESNA
C3529010|T121|1363915|RXNORM|BIS-ETHOXYDIGLYCOL SUCCINATE|BIS-ETHOXYDIGLYCOL SUCCINATE
C2741010|T129|900113|RXNORM|REDBERRY JUNIPER POLLEN EXTRACT|JUNIPERUS PINCHOTII POLLEN
C3504820|T121|1356709|RXNORM|LYSINE THIAZOLIDINE CARBOXYLATE|LYSINE THIAZOLIDINE CARBOXYLATE
C3504819|T121|1356708|RXNORM|LEUCOJUM AESTIVUM BULB EXTRACT|LEUCOJUM AESTIVUM BULB EXTRACT
C3555524|T121|1374401|RXNORM|MANSOA ALLIACEA BARK EXTRACT|MANSOA ALLIACEA BARK EXTRACT
C3818724|T109|1535215|RXNORM|DI-C12-13 ALKYL TARTRATE|DI-C12-13 ALKYL TARTRATE
C3504815|T121|1356703|RXNORM|PROPYLENE GLYCOL MYRISTYL ETHER ACETATE|PROPYLENE GLYCOL MYRISTYL ETHER ACETATE
C1509675|T121|1356702|RXNORM|PPG-10 CETYL ETHER|PPG-10 CETYL ETHER
C3504814|T121|1356701|RXNORM|HYDROXYLATED LANOLIN|HYDROXYLATED LANOLIN
C3504813|T121|1356700|RXNORM|CUCUMIS MELO VAR. CANTALUPENSIS WHOLE EXTRACT|CUCUMIS MELO VAR. CANTALUPENSIS WHOLE EXTRACT
C3504818|T109|1356707|RXNORM|PEG-7 HYDROGENATED CASTOR OIL|PEG-7 HYDROGENATED CASTOR OIL
C3504817|T121|1356706|RXNORM|SILANEDIOL SALICYLATE|SILANEDIOL SALICYLATE
C3504816|T121|1356705|RXNORM|TABEBUIA IMPETIGINOSA WHOLE EXTRACT|TABEBUIA IMPETIGINOSA WHOLE EXTRACT
C3503277|T121|1356704|RXNORM|SAUSSUREA GOSSIPIPHORA EXTRACT|SAUSSUREA GOSSIPIPHORA EXTRACT
C0060173|T121|24846|RXNORM|FENIPENTOL|FENIPENTOL
C0060167|T121|24840|RXNORM|FENETHYLLINE|FENETYLLINE
C1165377|T121|349753|RXNORM|SODIUM PHOSPHATE, MONOBASIC, ANHYDROUS|SODIUM PHOSPHATE, MONOBASIC, ANHYDROUS
C0981934|T129|349978|RXNORM|OAT SMUT ALLERGENIC EXTRACT|USTILAGO AVENAE ALLERGENIC EXTRACT
C3488181|T121|1426898|RXNORM|QUININE ARSENITE|QUININE ARSENITE
C0525005|T121|134527|RXNORM|NELFINAVIR|NELFINAVIR
C1874166|T121|705056|RXNORM|ALUMINUM HYDROXIDE / CALCIUM CARBONATE / MAGNESIUM HYDROXIDE|ALUMINUM HYDROXIDE / CALCIUM CARBONATE / MAGNESIUM HYDROXIDE
C2369985|T121|827116|RXNORM|CARBETAPENTANE / PSEUDOEPHEDRINE / PYRILAMINE|CARBETAPENTANE / PSEUDOEPHEDRINE / PYRILAMINE
C3256401|T121|1310495|RXNORM|BETA-CITRONELLOL, (R)-|BETA-CITRONELLOL, (R)-
C2080551|T121|817497|RXNORM|GUAIFENESIN / HYDROCODONE / PHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE|GUAIFENESIN / HYDROCODONE / PHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C1330008|T121|817496|RXNORM|HYDROCHLOROTHIAZIDE / OLMESARTAN|HYDROCHLOROTHIAZIDE / OLMESARTAN
C2742502|T129|1535922|RXNORM|RAMUCIRUMAB|RAMUCIRUMAB
C2827078|T121|1305896|RXNORM|ALUMINUM ZIRCONIUM TETRACHLOROHYDREX GLY|ALUMINUM ZIRCONIUM TETRACHLOROHYDREX GLY
C3818702|T109|1535931|RXNORM|PYROLIGNEOUS ACID|PYROLIGNEOUS ACID
C1828054|T121|802591|RXNORM|BENZOCAINE / TYROTHRICIN|BENZOCAINE / TYROTHRICIN
C0146196|T121|1535930|RXNORM|TOLTRAZURIL|TOLTRAZURIL
C3853832|T121|1591950|RXNORM|CINCHONA OFFICINALIS WHOLE EXTRACT|CINCHONA OFFICINALIS WHOLE EXTRACT
C0023413|T127|6313|RXNORM|LEUCOVORIN|LEUCOVORIN
C2930014|T121|1009119|RXNORM|MANNITOL / MECOBALAMIN|MANNITOL / MECOBALAMIN
C2930013|T121|1009118|RXNORM|FLUOCINONIDE / NEOMYCIN|FLUOCINONIDE / NEOMYCIN
C0033371|T125|1426890|RXNORM|PROLACTIN|PROLACTIN
C2930008|T121|1009113|RXNORM|POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC|POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC
C2930007|T121|1009112|RXNORM|DEXTROMETHORPHAN / THEOPHYLLINE|DEXTROMETHORPHAN / THEOPHYLLINE
C2930006|T121|1009111|RXNORM|ALANINE / ARGININE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM ACETATE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TYROSINE / VALI|ALANINE / ARGININE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM ACETATE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TYROSINE / VALINE
C2930005|T121|1009110|RXNORM|CHLORHEXIDINE / ETHANOL|CHLORHEXIDINE / ETHANOL
C2930012|T121|1009117|RXNORM|AJMALICINE / ALMITRINE|AJMALICINE / ALMITRINE
C2930011|T121|1009116|RXNORM|LOPERAMIDE / NEOMYCIN|LOPERAMIDE / NEOMYCIN
C2930010|T121|1009115|RXNORM|GINSENG PREPARATION / VITAMIN B 12|GINSENG PREPARATION / VITAMIN B 12
C2930009|T121|1009114|RXNORM|DIAZEPAM / OCTYLONIUM|DIAZEPAM / OCTYLONIUM
C0525678|T121|134748|RXNORM|RASAGILINE|RASAGILINE
C3645207|T121|1426892|RXNORM|POLIDRONIUM|POLIDRONIUM
C1533695|T197|1426894|RXNORM|POTASSIUM ARSENITE|POTASSIUM ARSENITE
C0064624|T121|1546426|RXNORM|LAIDLOMYCIN|LAIDLOMYCIN
C0039771|T121|10438|RXNORM|THEOPHYLLINE|THEOPHYLLINE
C3495132|T121|1351898|RXNORM|ASCARIS LUMBRICOIDES PREPARATION|ASCARIS LUMBRICOIDES PREPARATION
C2731567|T129|895588|RXNORM|RED DELICIOUS APPLE ALLERGENIC EXTRACT|RED DELICIOUS APPLE ALLERGENIC EXTRACT
C0038467|T196|10122|RXNORM|STRONTIUM|STRONTIUM
C0039736|T131|10432|RXNORM|THALIDOMIDE|THALIDOMIDE
C3495100|T121|1351897|RXNORM|PARIETARIA OFFICINALIS EXTRACT|PARIETARIA OFFICINALIS EXTRACT
C0039763|T121|10437|RXNORM|THEOBROMINE|THEOBROMINE
C0946377|T121|1427069|RXNORM|SEBACATE|SEBACATE
C3645256|T121|1427063|RXNORM|STAPHYLOCOCCUS AUREUS IMMUNOSERUM|STAPHYLOCOCCUS AUREUS IMMUNOSERUM
C0771424|T121|236174|RXNORM|PRIFINIUM|PRIFINIUM
C3497913|T121|1427060|RXNORM|PROPYLENE GLYCOL HEPTANOATE|PROPYLENE GLYCOL HEPTANOATE
C0220926|T197|1427067|RXNORM|THIOCYANATE|THIOCYANATE
C3159524|T121|1427065|RXNORM|METHYL UNDECENOYL LEUCINATE|METHYL UNDECENOYL LEUCINATE
C3475215|T121|1427064|RXNORM|ACETYLATED SUCROSE DISTEARATE|ACETYLATED SUCROSE DISTEARATE
C3486721|T121|1336265|RXNORM|BRYONIA DIOICA ROOT EXTRACT|BRYONIA DIOICA ROOT EXTRACT
C3666925|T121|1437987|RXNORM|TRIMETHYLPENTANEDIYL DIBENZOATE|TRIMETHYLPENTANEDIYL DIBENZOATE
C0360068|T121|619354|RXNORM|HYDROTALCITE / SIMETHICONE|HYDROTALCITE / SIMETHICONE
C3474935|T121|1421890|RXNORM|POLYGLYCERYL-6 DISTEARATE|POLYGLYCERYL-6 DISTEARATE
C3536941|T121|1430254|RXNORM|LINALOOL, (+)-|LINALOOL, (+)-
C2351315|T109|1421892|RXNORM|HEXYL SALICYLATE|HEXYL SALICYLATE
C0012294|T121|3419|RXNORM|DIHYDROERGOTOXINE|DIHYDROERGOTOXINE
C2740250|T129|898324|RXNORM|LODGEPOLE PINE POLLEN EXTRACT|PINUS CONTORTA POLLEN EXTRACT
C3181682|T121|1363268|RXNORM|CABOZANTINIB|CABOZANTINIB
C2702419|T129|891658|RXNORM|PEANUT ALLERGENIC EXTRACT|PEANUT ALLERGENIC EXTRACT
C2356374|T129|804187|RXNORM|YELLOW-FEVER VIRUS VACCINE, 17D-204 STRAIN|YELLOW-FEVER VIRUS VACCINE, 17D-204 STRAIN
C3857950|T121|1552276|RXNORM|BOS TAURUS PARASYMPATHETIC NERVE PREPARATION|BOS TAURUS PARASYMPATHETIC NERVE PREPARATION
C2726186|T129|891652|RXNORM|NUTMEG ALLERGENIC EXTRACT|NUTMEG ALLERGENIC EXTRACT
C0939803|T121|1372255|RXNORM|GOLDENSEAL EXTRACT|HYDRASTIS CANADENSIS EXTRACT
C0304112|T121|1305670|RXNORM|PINE NEEDLE OIL (PINUS SYLVESTRIS)|PINE NEEDLE OIL (PINUS SYLVESTRIS)
C3486625|T121|1372253|RXNORM|MELILOTUS EXTRACT|MELILOTUS INDICUS SEED EXTRACT
C3256845|T121|1372251|RXNORM|GREATER GALANGAL EXTRACT|THAI GALANGAL EXTRACT
C3255837|T121|1372250|RXNORM|ACHILLEA MILLEFOLIUM EXTRACT|ACHILLEA MELLEFOLIUM EXTRACT
C0600489|T130|155122|RXNORM|PHENOLPHTHALEIN|PHENOLPHTHALEIN
C3163233|T121|1115926|RXNORM|BURWEED MARSHELDER POLLEN EXTRACT / ROUGH MARSHELDER POLLEN EXTRACT|BURWEED MARSHELDER POLLEN EXTRACT / ROUGH MARSHELDER POLLEN EXTRACT
C3473193|T121|1298292|RXNORM|ASCORBIC ACID / BETA CAROTENE / ERGOCALCIFEROL / FOLIC ACID / NIACIN / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E|ASCORBIC ACID / BETA CAROTENE / ERGOCALCIFEROL / FOLIC ACID / NIACIN / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E
C0051654|T121|1006397|RXNORM|AMINOPENTAMIDE|AMINOPENTAMIDE
C2702352|T129|891514|RXNORM|BRAZIL NUT ALLERGENIC EXTRACT|BRAZIL NUT ALLERGENIC EXTRACT
C1874196|T121|690790|RXNORM|AMINOPHYLLINE / EPHEDRINE / PHENOBARBITAL / POTASSIUM IODIDE|AMINOPHYLLINE / EPHEDRINE / PHENOBARBITAL / POTASSIUM IODIDE
C1874198|T121|690793|RXNORM|AMINOPHYLLINE / POTASSIUM IODIDE|AMINOPHYLLINE / POTASSIUM IODIDE
C1874197|T121||RXNORM|AMINOPHYLLINE / PHENOBARBITAL
C0065932|T127|29491|RXNORM|MENADIOL|MENADIOL
C0065936|T127|29495|RXNORM|MENATETRENONE|MENATETRENONE
C2722022|T129|867274|RXNORM|NEUROSPORA INTERMEDIA ALLERGENIC EXTRACT|NEUROSPORA INTERMEDIA ALLERGENIC EXTRACT
C0054147|T130|1114345|RXNORM|BRONOPOL|BRONOPOL
C2929306|T121|1008402|RXNORM|ALUMINUM CHLORIDE / POTASSIUM CHLORATE|ALUMINUM CHLORIDE / POTASSIUM CHLORATE
C2929307|T121|1008403|RXNORM|NITROFURANTOIN / SULFADIAZINE|NITROFURANTOIN / SULFADIAZINE
C2929304|T121|1008400|RXNORM|CAFFEINE / GUARANA PREPARATION|CAFFEINE / GUARANA PREPARATION
C2929305|T121|1008401|RXNORM|CODEINE / GUAIFENESIN / PHENYLTOLOXAMINE|CODEINE / GUAIFENESIN / PHENYLTOLOXAMINE
C2929310|T121|1008406|RXNORM|ALBUTEROL / AMBROXOL|ALBUTEROL / AMBROXOL
C2929311|T121|1008407|RXNORM|LAURETH-9 / MEPIVACAINE|MEPIVACAINE / POLIDOCANOL
C2929308|T121|1008404|RXNORM|ANTIPYRINE / CALCIUM CHLORIDE|ANTIPYRINE / CALCIUM CHLORIDE
C2929309|T121|1008405|RXNORM|DIHYDROERGOTAMINE / ETILEFRINE|DIHYDROERGOTAMINE / ETILEFRINE
C2057529|T121|819395|RXNORM|ETHYLMORPHINE / TERPIN HYDRATE|ETHYLMORPHINE / TERPIN HYDRATE
C2740799|T129|899742|RXNORM|DATE ALLERGENIC EXTRACT|DATE ALLERGENIC EXTRACT
C2929312|T121|1008408|RXNORM|DIPYRONE / TIEMONIUM|DIPYRONE / TIEMONIUM
C2929313|T121|1008409|RXNORM|NORFENEFRINE / PHOLEDRINE|NORFENEFRINE / PHOLEDRINE
C2740802|T129|899746|RXNORM|FLOUNDER ALLERGENIC EXTRACT|FLOUNDER ALLERGENIC EXTRACT
C0005096|T121|1422|RXNORM|BENZPHETAMINE|BENZPHETAMINE
C1874500|T121|690247|RXNORM|BENZOCAINE / BUTAMBEN / TETRACAINE|BENZOCAINE / BUTAMBEN / TETRACAINE
C1874499|T121|690246|RXNORM|BENZOCAINE / BORIC ACID|BENZOCAINE / BORIC ACID
C1874498|T121|690245|RXNORM|BENZOCAINE / BISMUTH SUBNITRATE / CERIUM OXALATE|BENZOCAINE / BISMUTH SUBNITRATE / CERIUM OXALATE
C0005100|T121|1426|RXNORM|BENZYL ALCOHOL|BENZYL ALCOHOL
C0005100|T121|1426|RXNORM|BENZYL ALCOHOL|BENZYL ALCOHOL
C0012133|T121|3364|RXNORM|DIDANOSINE|DIDANOSINE
C0064088|T121|28012|RXNORM|ISOTHIPENDYL|ISOTHIPENDYL
C3864968|T121|1597118|RXNORM|CHONDROITIN SULFATES / GLUCOSAMINE / IBUPROFEN|CHONDROITIN SULFATES / GLUCOSAMINE / IBUPROFEN
C0012125|T121|3361|RXNORM|DICYCLOMINE|DICYCLOVERINE
C0768182|T129|234449|RXNORM|IODINE-131-TOSITUMOMAB|TOSITUMOMAB/IODINE (131I) TOSITUMOMAB
C0012132|T121|3363|RXNORM|ZALCITABINE|ZALCITABINE
C2194208|T121|818806|RXNORM|FERROUS FUMARATE / THIAMINE|FERROUS FUMARATE / THIAMINE
C0006982|T121|2019|RXNORM|CARBIDOPA|CARBIDOPA
C3859185|T121|1592295|RXNORM|FORMALDEHYDE SULFOXYLATE|FORMALDEHYDE SULFOXYLATE
C0304139|T109|1362137|RXNORM|HYSSOP OIL|HYSSOP OIL
C0382876|T109|1362136|RXNORM|TETRAHYDRODIFERULOYLMETHANE|TETRAHYDRODIFERULOYLMETHANE
C0015528|T126|4271|RXNORM|FACTOR XIII|FACTOR XIII
C3528223|T109|1362134|RXNORM|ARABICA COFFEE OIL|ARABICA COFFEE OIL
C3700903|T116|1486022|RXNORM|PALMITOYLLYSYLVALYLDIAMINOBUTYROYLTHREONINE|PALMITOYLLYSYLVALYLDIAMINOBUTYROYLTHREONINE
C0015620|T121|4278|RXNORM|FAMOTIDINE|FAMOTIDINE
C0243879|T109|1486028|RXNORM|2-HYDROXYDECANOATE|2-HYDROXYDECANOATE
C3528225|T109|1362138|RXNORM|JOJOBA BUTTER|JOJOBA BUTTER
C0020411|T130|5556|RXNORM|HYMECROMONE|HYMECROMONE
C0020404|T121|5553|RXNORM|HYDROXYZINE|HYDROXYZINE
C0020402|T121|5552|RXNORM|HYDROXYUREA|HYDROXYUREA
C2079566|T121|812477|RXNORM|AMITRIPTYLINE / DIAZEPAM / PERPHENAZINE|AMITRIPTYLINE / DIAZEPAM / PERPHENAZINE
C0006979|T121|2017|RXNORM|CARBENOXOLONE|CARBENOXOLONE
C3257280|T121|1311584|RXNORM|CYMBOPOGON SCHOENANTHUS TOP EXTRACT|CYMBOPOGON SCHOENANTHUS TOP EXTRACT
C0771555|T121|1592259|RXNORM|POTASSIUM ASCORBATE|POTASSIUM ASCORBATE
C0304612|T121|91311|RXNORM|DIFLORASONE|DIFLORASONE
C0025856|T121|1311585|RXNORM|METOMIDATE|METOMIDATE
C0076648|T121|38248|RXNORM|TIADENOL|TIADENOL
C0771339|T121|1424676|RXNORM|CALTERIDOL|CALTERIDOL
C3256281|T109|1424674|RXNORM|C20-22 ALKYL PHOSPHATE|C20-22 ALKYL PHOSPHATE
C3255718|T121|1311586|RXNORM|PINUS MASSONIANA RESIN|PINUS MASSONIANA RESIN
C0771601|T197|1424671|RXNORM|CALCIUM HYPOPHOSPHITE|CALCIUM HYPOPHOSPHITE
C3256337|T109|1309394|RXNORM|AMPELOPSIS JAPONICA ROOT EXTRACT|AMPELOPSIS JAPONICA ROOT EXTRACT
C0032821|T196|8588|RXNORM|POTASSIUM|KALIUM
C0077192|T131|1426813|RXNORM|TRIMETHYLOLPROPANE TRIACRYLATE|TRIMETHYLOLPROPANE TRIACRYLATE
C3256340|T109|1309397|RXNORM|ANACYCLUS PYRETHRUM ROOT EXTRACT|ANACYCLUS PYRETHRUM ROOT EXTRACT
C1952586|T121|1309390|RXNORM|SAFFLOWER EXTRACT|SAFFLOWER EXTRACT
C3257532|T121|1309391|RXNORM|SUNFLOWER SEED EXTRACT|SUNFLOWER SEED EXTRACT
C3256015|T109|1309392|RXNORM|ALPINIA ZERUMBET LEAF EXTRACT|ALPINIA ZERUMBET LEAF EXTRACT
C1509305|T121|1426816|RXNORM|DEXTRATES|DEXTRATES
C3485005|T121|1311580|RXNORM|CULLEN CORYLIFOLIUM FRUIT EXTRACT|CULLEN CORYLIFOLIUM FRUIT EXTRACT
C3256590|T121|1309398|RXNORM|AESCULUS HIPPOCASTANUM BARK EXTRACT|AESCULUS HIPPOCASTANUM BARK EXTRACT
C3255625|T121|1311581|RXNORM|ZANTHOXYLUM PIPERITUM FRUIT PULP EXTRACT|ZANTHOXYLUM PIPERITUM FRUIT PULP EXTRACT
C0663378|T121|1311582|RXNORM|NIFURPIPONE|NIFURPIPONE
C1095912|T121|1362688|RXNORM|SHIITAKE MUSHROOM PREPARATION|SHIITAKE MUSHROOM PREPARATION
C1633985|T121|622157|RXNORM|BENZALKONIUM / CETRIMIDE|BENZALKONIUM / CETRIMIDE
C2699757|T121|1303098|RXNORM|ACLIDINIUM|ACLIDINIUM
C3663397|T121|1432979|RXNORM|ONCORHYNCHUS MASOU SPERM DNA|ONCORHYNCHUS MASOU SPERM DNA
C0028004|T121|1311583|RXNORM|NICARBAZIN|NICARBAZIN
C0014047|T005|1439114|RXNORM|JAPANESE ENCEPHALITIS VIRUS|JAPANESE ENCEPHALITIS VIRUS
C0021741|T129|5882|RXNORM|INTERFERON GAMMA-1B|INTERFERON GAMMA-1B
C0021735|T129|5880|RXNORM|INTERFERON ALFA-2B|INTERFERON ALFA-2B
C0021735|T129|5880|RXNORM|INTERFERON ALFA-2B|INTERFERON ALFA-2B
C2346747|T121|1440271|RXNORM|AMOPROXAN|AMOPROXAN
C0051733|T121|1440270|RXNORM|AMONAFIDE|AMONAFIDE
C3848705|T121|1545149|RXNORM|CANAGLIFLOZIN / METFORMIN|CANAGLIFLOZIN / METFORMIN
C2928508|T121|1007590|RXNORM|FERROUS GLYCINE SULFATE / FOLIC ACID|FERROUS GLYCINE SULFATE / FOLIC ACID
C0016911|T196|1310171|RXNORM|GADOLINIUM|GADOLINIUM
C2929175|T121|1008268|RXNORM|BLACK PEPPER PREPARATION / ECHINACEA PREPARATION|BLACK PEPPER PREPARATION / ECHINACEA PREPARATION
C2928433|T121|1007511|RXNORM|CALCIUM CARBONATE / ERGOCALCIFEROL / SOYBEAN PREPARATION|CALCIUM CARBONATE / ERGOCALCIFEROL / SOYBEAN PREPARATION
C2928432|T121|1007510|RXNORM|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / CUPRIC OXIDE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM OXIDE / NIACIN / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / CUPRIC OXIDE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM OXIDE / NIACIN / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC OXIDE
C2928435|T121|1007513|RXNORM|MAGNESIUM SULFATE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC|MAGNESIUM SULFATE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC
C2928510|T121|1007592|RXNORM|CHLORZOXAZONE / FLUFENAMATE|CHLORZOXAZONE / FLUFENAMATE
C2928437|T121|1007515|RXNORM|SODIUM PHOSPHATE, DIBASIC / UREA|SODIUM PHOSPHATE, DIBASIC / UREA
C2928436|T121|1007514|RXNORM|CALCIUM CARBONATE / ERGOCALCIFEROL / VITAMIN K 1|CALCIUM CARBONATE / ERGOCALCIFEROL / VITAMIN K 1
C2928439|T121|1007517|RXNORM|BENZETHONIUM / DIMETHICONE|BENZETHONIUM / DIMETHICONE
C2928438|T121|1007516|RXNORM|CALCIUM PHOSPHATE / ERGOCALCIFEROL|CALCIUM PHOSPHATE / ERGOCALCIFEROL
C2928441|T121|1007519|RXNORM|CALCIUM ASCORBATE / FERROUS ASPARTO GLYCINATE / POLYSACCHARIDE IRON COMPLEX / SUCCINIC ACID|CALCIUM ASCORBATE / FERROUS ASPARTO GLYCINATE / POLYSACCHARIDE IRON COMPLEX / SUCCINIC ACID
C2928440|T121|1007518|RXNORM|HEPARINOIDS / LAURETH-4|HEPARINOIDS / LAURETH-4
C2918506|T121|995720|RXNORM|CLADOSOPRIUM CLADOSPORIOIDES ALLERGENIC EXTRACT|CLADOSOPRIUM CLADOSPORIOIDES ALLERGENIC EXTRACT
C2928512|T121|1007594|RXNORM|BUTACAINE / OLEATE|BUTACAINE / OLEATE
C0076079|T195|37775|RXNORM|TEMOCILLIN|TEMOCILLIN
C2928187|T121|1007265|RXNORM|NITRIC OXIDE / NITROGEN|NITRIC OXIDE / NITROGEN
C2928514|T121|1007596|RXNORM|GONADORELIN / THYROTROPIN-RELEASING HORMONE|GONADORELIN / THYROTROPIN-RELEASING HORMONE
C0245109|T121|72435|RXNORM|ANAKINRA|ANAKINRA
C2756450|T129|968197|RXNORM|TRICHODERMA HARZIANUM EXTRACT|TRICHODERMA HARZIANUM EXTRACT
C3855916|T129|1549330|RXNORM|COCCIDIODIDES IMMITIS SPHERULE PREPARATION|COCCIDIOIDES IMMITIS SPHERULE
C3855917|T109|1549331|RXNORM|ROSIN PARTIALLY DIMERIZED GLYCEROL ESTER|ROSIN PARTIALLY DIMERIZED GLYCEROL ESTER
C0074289|T123|1549332|RXNORM|SELENOCYSTEINE|SELENOCYSTEINE
C1276898|T121|389190|RXNORM|FIBRINOGEN / THROMBIN|FIBRINOGEN / THROMBIN
C0043040|T131|11291|RXNORM|WASP VENOMS|WASP VENOMS
C0718096|T121|214866|RXNORM|TRANDOLAPRIL / VERAPAMIL|TRANDOLAPRIL / VERAPAMIL
C4281713|T121|27291|RXNORM|HYDROXYPROPYLCELLULOSE|HYDROXYPROPYL CELLULOSE
C0065832|T121|29410|RXNORM|MEBEVERINE|MEBEVERINE
C3818815|T109|1489759|RXNORM|AMMONIUM LAUROYL SARCOSINATE|AMMONIUM LAUROYL SARCOSINATE
C0037521|T197|9884|RXNORM|SODIUM IODIDE|SODIUM IODIDE
C1456409|T121|475969|RXNORM|ETRAVIRINE|ETRAVIRINE
C1456408|T125|475968|RXNORM|LIRAGLUTIDE|LIRAGLUTIDE
C1875661|T121|689759|RXNORM|PHOSPHORIC ACID / SODIUM FLUORIDE|PHOSPHORIC ACID / SODIUM FLUORIDE
C3486597|T121|1313321|RXNORM|CUPRIC CARBONATE BASIC|CUPRIC CARBONATE BASIC
C1875660|T121|689757|RXNORM|PHENYLEPHRINE / ZINC SULFATE|PHENYLEPHRINE / ZINC SULFATE
C1875659|T121|689756|RXNORM|PHENYLEPHRINE / SULFACETAMIDE|PHENYLEPHRINE / SULFACETAMIDE
C1875658|T121|689755|RXNORM|PHENYLEPHRINE / SCOPOLAMINE|PHENYLEPHRINE / SCOPOLAMINE
C3538555|T109|1373037|RXNORM|TURMERIC OIL|TURMERIC OIL
C2701343|T129|852140|RXNORM|PEPPER TREE POLLEN EXTRACT|SCHINUS MOLLE POLLEN EXTRACT
C1875657|T121|689752|RXNORM|PHENYLEPHRINE / PREDNISOLONE / SULFACETAMIDE|PHENYLEPHRINE / PREDNISOLONE / SULFACETAMIDE
C1875655|T121|689750|RXNORM|PHENYLEPHRINE / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE|PHENYLEPHRINE / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE
C1828124|T121|687333|RXNORM|ESTRADIOL / LEVONORGESTREL|ESTRADIOL / LEVONORGESTREL
C0029193|T121|7688|RXNORM|METAPROTERENOL|METAPROTERENOL
C0029193|T121|7688|RXNORM|METAPROTERENOL|METAPROTERENOL
C1831905|T121|711942|RXNORM|ELTROMBOPAG|ELTROMBOPAG
C1654726|T121|978673|RXNORM|HEME IRON POLYPEPTIDE|HEME IRON POLYPEPTIDE
C0384228|T121|117466|RXNORM|TENOFOVIR|TENOFOVIR
C3700877|T121|1487085|RXNORM|CRAMBE MARITIMA WHOLE EXTRACT|CRAMBE MARITIMA WHOLE EXTRACT
C0772481|T121|237141|RXNORM|TIBEZONIUM IODIDE|TIBEZONIUM IODIDE
C0290883|T121|84857|RXNORM|ANASTROZOLE|ANASTROZOLE
C1874489|T121|690077|RXNORM|BENZALKONIUM / LIDOCAINE|BENZALKONIUM / LIDOCAINE
C0733758|T125|227518|RXNORM|FOLLICLE STIMULATING HORMONE|FOLLICLE STIMULATING HORMONE
C2928073|T121|1007151|RXNORM|CINNARIZINE / DOBESILIC ACID|CINNARIZINE / DOBESILIC ACID
C1443660|T121|465366|RXNORM|BUPIVACAINE / LIDOCAINE|BUPIVACAINE / LIDOCAINE
C0041479|T123|10958|RXNORM|TYRAMINE|TYRAMINE
C2073800|T121|819896|RXNORM|BROMHEXINE / CHLOPHEDIANOL|BROMHEXINE / CHLOPHEDIANOL
C3651729|T168|1429968|RXNORM|WINE GRAPE JUICE|WINE GRAPE JUICE
C0598436|T121|154643|RXNORM|MESTRANOL / NORETHINDRONE|MESTRANOL / NORETHINDRONE
C0937627|T121|283567|RXNORM|GREEN TEA LEAF EXTRACT|GREEN TEA LEAF EXTRACT
C2702407|T129|995699|RXNORM|COCHLIOBOLUS SPICIFER ALLERGENIC EXTRACT|COCHLIOBOLUS SPICIFER ALLERGENIC EXTRACT
C0055804|T121|21171|RXNORM|CITIOLONE|CITIOLONE
C0717511|T121|214317|RXNORM|BISOPROLOL / HYDROCHLOROTHIAZIDE|BISOPROLOL / HYDROCHLOROTHIAZIDE
C3496088|T121|1315116|RXNORM|EGGPLANT EXTRACT|EGGPLANT EXTRACT
C2194020|T121|814034|RXNORM|BETAMETHASONE / TERFENADINE|BETAMETHASONE / TERFENADINE
C1508746|T121|1315115|RXNORM|EGG EXTRACT|EGG EXTRACT
C3179549|T121|1551291|RXNORM|DULAGLUTIDE|DULAGLUTIDE
C0007558|T195|2190|RXNORM|CEFSULODIN|CEFSULODIN
C0937629|T121|283569|RXNORM|GYMNEMA SYLVESTRE PREPARATION|GYMNEMA SYLVESTRE PREPARATION
C1704256|T123|1426465|RXNORM|TRANSFORMING GROWTH FACTOR BETA 1|TRANSFORMING GROWTH FACTOR BETA 1
C0218501|T131|1433761|RXNORM|FIPRONIL|FIPRONIL
C3496085|T129|1315113|RXNORM|COTTON FIBER EXTRACT|COTTON FIBER EXTRACT
C2142852|T121|818422|RXNORM|BROMPHENIRAMINE / CODEINE / PSEUDOEPHEDRINE|BROMPHENIRAMINE / CODEINE / PSEUDOEPHEDRINE
C3256613|T109|1426466|RXNORM|DUNALIELLA SALINA EXTRACT|DUNALIELLA SALINA EXTRACT
C3500693|T121|1315112|RXNORM|CASEIN, LACTOCOCCUS LACTIS CULTURED, PENICILLIUM CAMEMBERTI CULTURED, AGED|CASEIN, LACTOCOCCUS LACTIS CULTURED, PENICILLIUM CAMEMBERTI CULTURED, AGED
C2929094|T121|1008187|RXNORM|BISMUTH SUBNITRATE / LAURETH-9 / ZINC OXIDE|BISMUTH SUBNITRATE / POLIDOCANOL / ZINC OXIDE
C2929093|T121|1008186|RXNORM|BENZOCAINE / HEXYLRESORCINOL|BENZOCAINE / HEXYLRESORCINOL
C2929092|T121|1008185|RXNORM|CETRIMIDE / LIDOCAINE|CETRIMIDE / LIDOCAINE
C2929091|T121|1008184|RXNORM|DIAZEPAM / SCOPOLAMINE|DIAZEPAM / SCOPOLAMINE
C2929090|T121|1008183|RXNORM|LIDOCAINE / NEOMYCIN|LIDOCAINE / NEOMYCIN
C2929089|T121|1008182|RXNORM|DIPHENHYDRAMINE / LIDOCAINE|DIPHENHYDRAMINE / LIDOCAINE
C2929088|T121|1008181|RXNORM|THIAMINE / VITAMIN E|THIAMINE / VITAMIN E
C2929087|T121|1008180|RXNORM|IODOQUINOL / PAPAVERINE / SUCCINYLSULFATHIAZOLE|IODOQUINOL / PAPAVERINE / SUCCINYLSULFATHIAZOLE
C0016967|T121|4637|RXNORM|GALANTAMINE|GALANTAMINE
C3500691|T121|1315110|RXNORM|CASEIN, LACTOCOCCUS LACTIS CULTURED|CASEIN, LACTOCOCCUS LACTIS CULTURED
C3505775|T109|1359283|RXNORM|TETRASILANE|TETRASILANE
C2929096|T121|1008189|RXNORM|EUCALYPTUS EXTRACT / METHYL SALICYLATE|EUCALYPTUS EXTRACT / METHYL SALICYLATE
C2929095|T121|1008188|RXNORM|BENPHOTHIAMINE / VITAMIN B6|BENPHOTHIAMINE / VITAMIN B6
C2709772|T129|854968|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 7F VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 7F VACCINE
C0370086|T121|618564|RXNORM|TRICHLOROACETATE|TRICHLOROACETATE
C3535919|T121|1368487|RXNORM|HYDROXYPROPYL BISSTEARYLDIMONIUM|HYDROXYPROPYL BISSTEARYLDIMONIUM
C0056601|T197|1423796|RXNORM|CUPROUS CHLORIDE|CUPROUS CHLORIDE
C3643350|T121|1423791|RXNORM|SUCROSE TETRASTEARATE TRIACETATE|SUCROSE TETRASTEARATE TRIACETATE
C3643349|T121|1423793|RXNORM|SODIUM LAURYL GLYCOL CARBOXYLATE|SODIUM LAURYL GLYCOL CARBOXYLATE
C0630395|T109|1423792|RXNORM|TILIROSIDE|TILIROSIDE
C0873078|T121|259415|RXNORM|ECHINACEA ANGUSTIFOLIA ROOT EXTRACT|ECHINACEA ANGUSTIFOLIA ROOT EXTRACT
C0074718|T197|1364794|RXNORM|SODIUM ARSENATE|SODIUM ARSENATE
C0076836|T121|38409|RXNORM|TOREMIFENE|TOREMIFENE
C1166253|T121|350528|RXNORM|SUMBUL|SUMBUL
C0076823|T121|38400|RXNORM|ATOMOXETINE|ATOMOXETINE
C2940023|T129|1014447|RXNORM|YELLOW SWEET CLOVER POLLEN EXTRACT|MELILOTUS OFFICINALIS POLLEN EXTRACT
C0772335|T121|236999|RXNORM|HELICIN|HELICIN
C0076829|T121|38404|RXNORM|TOPIRAMATE|TOPIRAMATE
C0770338|T121|235376|RXNORM|IRON BILE SALTS|IRON BILE SALTS
C0040238|T196|10603|RXNORM|TIN|TIN
C0040233|T121|10600|RXNORM|TIMOLOL|TIMOLOL
C0040233|T121|10600|RXNORM|TIMOLOL|TIMOLOL
C0770337|T121|235375|RXNORM|MALT EXTRACT|MALT EXTRACT
C2929884|T121|1008989|RXNORM|NICOBOXIL / VANILLYL-N-NONYLAMIDE|NICOBOXIL / VANILLYL-N-NONYLAMIDE
C2929883|T121|1008988|RXNORM|ASPIRIN / NAFRONYL|ASPIRIN / NAFRONYL
C2929882|T121|1008987|RXNORM|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM ACETATE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / POTASSIUM ACETATE / PROLINE / SERINE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM ACETATE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / POTASSIUM ACETATE / PROLINE / SERINE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929881|T121|1008986|RXNORM|BETAINE / GLUTAMATE / METHYLCELLULOSE|BETAINE / GLUTAMATE / METHYLCELLULOSE
C2929880|T121|1008985|RXNORM|OXYGEN / XENON-133|OXYGEN / XENON-133
C2929879|T121|1008984|RXNORM|DEXTROMETHORPHAN / GUAIACOLSULFONATE / GUAIFENESIN / PYRILAMINE|DEXTROMETHORPHAN / GUAIACOLSULFONATE / GUAIFENESIN / PYRILAMINE
C2929877|T121|1008982|RXNORM|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929877|T121|1008982|RXNORM|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929876|T121|1008981|RXNORM|MEFRUSIDE / METHYLDOPA|MEFRUSIDE / METHYLDOPA
C2930441|T121|1008980|RXNORM|ACEBUTOLOL / NIFEDIPINE|ACEBUTOLOL / NIFEDIPINE
C0771662|T121|236395|RXNORM|METHYL DIACETYLCYSTEINATE|METHYL DIACETYLCYSTEINATE
C3282530|T121|1251581|RXNORM|IMIDACLOPRID / MOXIDECTIN|IMIDACLOPRID / MOXIDECTIN
C0771660|T121|236393|RXNORM|MIRISTALKONIUM|MIRISTALKONIUM
C0052585|T195|18469|RXNORM|SPARFLOXACIN|SPARFLOXACIN
C3488038|T025|1345682|RXNORM|HUMAN BREAST TUMOR CELL|HUMAN BREAST TUMOR CELL
C3486753|T121|1345680|RXNORM|LILIUM LANCIFOLIUM BULB EXTRACT|LILIUM LANCIFOLIUM BULB EXTRACT
C3487969|T121|1345681|RXNORM|JACOBAEA MARITIMA EXTRACT|JACOBAEA MARITIMA EXTRACT
C0064056|T121|27985|RXNORM|ISOPROPYL MYRISTATE|ISOPROPYL MYRISTATE
C0068314|T195|31435|RXNORM|ALLERGENIC EXTRACT, COTTONWOOD FREMONT|VALRUBICIN
C3486710|T121|1310006|RXNORM|BROMUS RAMOSUS FLOWER EXTRACT|BROMUS RAMOSUS FLOWER EXTRACT
C3484460|T121|1310007|RXNORM|ARALIA HISPIDA ROOT EXTRACT|ARALIA HISPIDA ROOT EXTRACT
C3472771|T121|1310004|RXNORM|PRUNUS PERSICA SEED EXTRACT|PRUNUS PERSICA SEED EXTRACT
C3257270|T121|1310005|RXNORM|PLANTAGO MAJOR LEAF EXTRACT|PLANTAGO MAJOR LEAF EXTRACT
C3486703|T121|1310002|RXNORM|HIPPOMANE MANCINELLA FRUITING LEAFY TWIG EXTRACT|HIPPOMANE MANCINELLA FRUITING LEAFY TWIG EXTRACT
C0772501|T121|237159|RXNORM|LEVALBUTEROL|LEVOSALBUTAMOL
C3465331|T121|1310000|RXNORM|PICEA ABIES FLOWER BUD EXTRACT|PICEA ABIES FLOWER BUD EXTRACT
C3486702|T121|1310001|RXNORM|HIERACIUM PILOSELLA FLOWERING TOP|HIERACIUM PILOSELLA FLOWERING TOP
C0872917|T121|259283|RXNORM|YUCCA EXTRACT|YUCCA EXTRACT
C3257279|T121|1310008|RXNORM|HIBISCUS ROSA-SINENSIS FLOWERING TOP EXTRACT|HIBISCUS ROSA-SINENSIS FLOWERING TOP EXTRACT
C3489004|T121|1310009|RXNORM|PRUNUS PERSICA FLOWER EXTRACT|PRUNUS PERSICA FLOWER EXTRACT
C0037134|T121|9793|RXNORM|SILVER SULFADIAZINE|SILVER SULFADIAZINE
C0081816|T197|40762|RXNORM|BISMUTH ALUMINATE|BISMUTH ALUMINATE
C0037138|T122|9796|RXNORM|SIMETHICONE|SIMETHICONE
C0037135|T121|9794|RXNORM|SILYMARIN|SILYMARIN
C2370726|T121|828682|RXNORM|FOSPROPOFOL|FOSPROPOFOL
C2730270|T129|892734|RXNORM|CALIFORNIA MUGWORT POLLEN EXTRACT|ARTEMISIA DOUGLASIANA POLLEN EXTRACT
C2975314|T195|1113697|RXNORM|GAMITHROMYCIN|GAMITHROMYCIN
C3665003|T122|1435110|RXNORM|POLYGLYCERYL-2 MONOISOSTEARATE|POLYGLYCERYL-2 MONOISOSTEARATE
C0052772|T195|18609|RXNORM|AZIDOCILLIN|AZIDOCILLIN
C0052762|T121|18603|RXNORM|AZELASTINE|AZELASTINE
C0052762|T121|18603|RXNORM|AZELASTINE|AZELASTINE
C0052759|T121|18600|RXNORM|AZATADINE|AZATADINE
C3538280|T121|1372481|RXNORM|POLYQUATERNIUM-37 (3000 MPA.S)|POLYQUATERNIUM-37 (3000 MPA.S)
C0939669|T121|285036|RXNORM|ACETAMINOPHEN / DOXYLAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / DOXYLAMINE / PSEUDOEPHEDRINE
C0771150|T121|1305554|RXNORM|ALCLOXA|ALCLOXA
C0002937|T121|820|RXNORM|INORGANIC PHOSPHATE|ANETHOLE TRITHIONE
C0907349|T121|274771|RXNORM|NELARABINE|NELARABINE
C3497614|T121|1310262|RXNORM|BOS TAURUS KNEE JOINT PREPARATION|BOVINE KNEE JOINT PREPARATION
C3497615|T121|1310263|RXNORM|BOS TAURUS LIMBIC SYSTEM PREPARATION|BOVINE LIMBIC SYSTEM PREPARATION
C3495984|T121|1310260|RXNORM|BOS TAURUS HIPPOCAMPUS PREPARATION|BOVINE HIPPOCAMPUS PREPARATION
C0032143|T126|8410|RXNORM|ALTEPLASE|ALTEPLASE
C2938201|T121|1310266|RXNORM|ANEMONE NEMOROSA EXTRACT|ANEMONE NEMOROSA EXTRACT
C3497618|T121|1310267|RXNORM|BOS TAURUS NERVE PREPARATION|BOVINE NERVE PREPARATION
C3497616|T121|1310264|RXNORM|BOS TAURUS LYMPH PREPARATION|BOVINE LYMPH PREPARATION
C3497617|T121|1310265|RXNORM|BOS TAURUS MESENCHYME PREPARATION|BOVINE MESENCHYME PREPARATION
C0039738|T196|1311633|RXNORM|THALLIUM|THALLIUM
C0621910|T121|168651|RXNORM|PREDNAZOLINE|PREDNAZOLINE
C3255773|T121|1311630|RXNORM|LOWBUSH BLUEBERRY EXTRACT|LOWBUSH BLUEBERRY EXTRACT
C0066779|T121|30206|RXNORM|MONOSULFIRAM|SULFIRAM
C1098510|T121|321208|RXNORM|FONDAPARINUX|FONDAPARINUX
C3486845|T121|1311263|RXNORM|SUS SCROFA THYMUS PREPARATION|PORCINE THYMUS PREPARATION
C2928641|T121|1007726|RXNORM|BISDEQUALINIUM / PREDNISOLONE|BISDEQUALINIUM / PREDNISOLONE
C2928642|T121|1007727|RXNORM|GLUCONOLACTONE / MAGNESIUM CARBONATE|GLUCONOLACTONE / MAGNESIUM CARBONATE
C2928639|T121|1007724|RXNORM|DEHYDROEPIANDROSTERONE / ESTRADIOL|ESTRADIOL / PRASTERONE
C2928640|T121|1007725|RXNORM|IDOXURIDINE / PREDNISOLONE|IDOXURIDINE / PREDNISOLONE
C2928637|T121|1007722|RXNORM|POVIDONE / TETRACYCLINE|POVIDONE / TETRACYCLINE
C2928638|T121|1007723|RXNORM|PODOPHYLLIN / SALICYLIC ACID|PODOPHYLLIN / SALICYLIC ACID
C2928636|T121|1007720|RXNORM|ALANINE / ARGININE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2928636|T121|1007720|RXNORM|ALANINE / ARGININE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C0600296|T121|155046|RXNORM|PENTOSAN POLYSULFATE|PENTOSAN POLYSULFATE
C0073629|T121|35825|RXNORM|GANIRELIX|GANIRELIX
C2928643|T121|1007728|RXNORM|ASCORBIC ACID / D-BIOTIN / FOLIC ACID / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|ASCORBIC ACID / D-BIOTIN / FOLIC ACID / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C3848522|T196|1546439|RXNORM|GERMANIUM CATION (4+)|GERMANIUM CATION (4+)
C3555535|T121|1373445|RXNORM|ISOSTEARYL HYDROXYSTEARATE|ISOSTEARYL HYDROXYSTEARATE
C3555536|T109|1373444|RXNORM|TAMANU OIL|TAMANU OIL
C3555534|T109|1373446|RXNORM|POLYQUATERNIUM-6 (15000 MW)|POLYQUATERNIUM-6 (15000 MW)
C0049065|T121|15657|RXNORM|DECITABINE|DECITABINE
C0039416|T130|1488818|RXNORM|TECHNETIUM TC 99M MEDRONATE|TECHNETIUM TC 99M MEDRONATE
C0065329|T121|29006|RXNORM|LYAPOLATE|LYAPOLATE
C0065331|T123|29008|RXNORM|LYCOPENE|LYCOPENE
C3531130|T121|1366142|RXNORM|CHOLECALCIFEROL / VITAMIN E|CHOLECALCIFEROL / VITAMIN E
C0076275|T121|37925|RXNORM|ORLISTAT|ORLISTAT
C0304348|T121|91101|RXNORM|ACETYL SALICYLATE|ACETYL SALICYLATE
C2728194|T129|1010915|RXNORM|CHOCOLATE ALLERGENIC EXTRACT|CHOCOLATE ALLERGENIC EXTRACT
C2701217|T129|851998|RXNORM|GIANT RAGWEED POLLEN EXTRACT|AMBROSIA TRIFIDA POLLEN EXTRACT
C0037209|T195|9806|RXNORM|SISOMICIN|SISOMICIN
C0981982|T130|851994|RXNORM|TIMOTHY GRASS POLLEN EXTRACT|TIMOTHY GRASS POLLEN EXTRACT
C2701211|T129|851990|RXNORM|SLENDER RAGWEED POLLEN EXTRACT|AMBROSIA TENUIFOLIA POLLEN EXTRACT
C3710013|T109|1488816|RXNORM|SAPONARIA OFFICINALIS LEAF EXTRACT|SAPONARIA OFFICINALIS LEAF EXTRACT
C0031495|T121|8175|RXNORM|PHENYLPROPANOLAMINE|PHENYLPROPANOLAMINE
C3709472|T121|1487507|RXNORM|PRUNUS ARMENIACA LEAF EXTRACT|PRUNUS ARMENIACA LEAF EXTRACT
C3709471|T109|1487505|RXNORM|GERANIUM MACULATUM ROOT OIL|GERANIUM MACULATUM ROOT OIL
C0319878|T004|1310914|RXNORM|CANDIDA PARAPSILOSIS|CANDIDA PARAPSILOSIS
C0033477|T007|1310910|RXNORM|PROPIONIBACTERIUM ACNES|PROPIONIBACTERIUM ACNES
C0033809|T007|1310913|RXNORM|PSEUDOMONAS AERUGINOSA|PSEUDOMONAS AERUGINOSA
C2193903|T121|822432|RXNORM|BUTHIAZIDE / METIPRANOLOL|BUTHIAZIDE / METIPRANOLOL
C3818785|T109|1491859|RXNORM|PINUS SYLVESTRIS BARK EXTRACT|PINUS SYLVESTRIS BARK EXTRACT
C3818786|T109|1491858|RXNORM|JOJOBA OIL, RANDOMIZED|JOJOBA OIL, RANDOMIZED
C0378091|T121|114817|RXNORM|ROXATIDINE|ROXATIDINE
C1720023|T121|644563|RXNORM|LAUROMACROGOLS / UREA|LAUROMACROGOLS / UREA
C3832873|T121|1539815|RXNORM|IMMATURE CITRUS SINENSIS FRUIT EXTRACT|IMMATURE CITRUS SINENSIS FRUIT EXTRACT
C2740662|T129|899480|RXNORM|HOPS ALLERGENIC EXTRACT|HOPS ALLERGENIC EXTRACT
C3159389|T121|1111064|RXNORM|BROMPHENIRAMINE / CHLOPHEDIANOL / PHENYLEPHRINE|BROMPHENIRAMINE / CHLOPHEDIANOL / PHENYLEPHRINE
C0851287|T196|258478|RXNORM|PHOSPHORUS 32|PHOSPHORUS 32
C0066774|T121|30202|RXNORM|MOFEBUTAZONE|MOFEBUTAZONE
C0521890|T195|1314589|RXNORM|TIAMULIN FUMARATE|TIAMULIN FUMARATE
C3255939|T121|1314588|RXNORM|HYDROGENATED POLYDECENE (550 MW)|HYDROGENATED POLYDECENE (550 MW)
C0993602|T121|1314587|RXNORM|CARDAMOM EXTRACT|CARDAMOM EXTRACT
C3500456|T121|1314586|RXNORM|CARTHAMUS TINCTORIUS SEEDCAKE EXTRACT|CARTHAMUS TINCTORIUS SEEDCAKE EXTRACT
C3500455|T121|1314585|RXNORM|POLYETHYLENE GLYCOL 11000|POLYETHYLENE GLYCOL 11000
C3500454|T121|1314584|RXNORM|UNCARIA SINENSIS WHOLE PREPARATION|UNCARIA SINENSIS WHOLE PREPARATION
C3500453|T121|1314583|RXNORM|HYDRASTIS CANADENSIS WHOLE PREPARATION|HYDRASTIS CANADENSIS WHOLE PREPARATION
C0107994|T121|47579|RXNORM|CABERGOLINE|CABERGOLINE
C0002607|T197|1299884|RXNORM|AMMONIA|AMMONIA
C0304110|T121|1314580|RXNORM|BITTER ORANGE OIL|BITTER ORANGE OIL
C3695977|T109|1483422|RXNORM|CUCUMBER SEED OIL|CUCUMBER SEED OIL
C3486676|T121|1353884|RXNORM|RHUS AROMATICA ROOT BARK EXTRACT|RHUS AROMATICA ROOT BARK EXTRACT
C0075770|T123|594680|RXNORM|DOCOSANOL|DOCOSANOL
C0717880|T121|214671|RXNORM|LAMIVUDINE / ZIDOVUDINE|LAMIVUDINE / ZIDOVUDINE
C3864827|T109|1597186|RXNORM|COMBRETUM MICRANTHUM LEAF EXTRACT|COMBRETUM MICRANTHUM LEAF EXTRACT
C2080485|T121|814664|RXNORM|ASPIRIN / PHENYLEPHRINE|ASPIRIN / PHENYLEPHRINE
C0939860|T121|285208|RXNORM|ARNICA MONTANA EXTRACT|ARNICA MONTANA EXTRACT
C2929124|T121|1008217|RXNORM|CLEMASTINE / DEXAMETHASONE|CLEMASTINE / DEXAMETHASONE
C2929123|T121|1008216|RXNORM|CLONIDINE / CYCLOTHIAZIDE|CLONIDINE / CYCLOTHIAZIDE
C2929122|T121|1008215|RXNORM|ASCORBIC ACID / DEQUALINIUM / TYROTHRICIN|ASCORBIC ACID / DEQUALINIUM / TYROTHRICIN
C2929121|T121|1008214|RXNORM|CHOLECALCIFEROL / SODIUM FLUORIDE|CHOLECALCIFEROL / SODIUM FLUORIDE
C2929120|T121|1008213|RXNORM|TETRACAINE / TRICARBAURINIUM|TETRACAINE / TRICARBAURINIUM
C2929119|T121|1008212|RXNORM|CINNARIZINE / DIHYDROERGOTAMINE|CINNARIZINE / DIHYDROERGOTAMINE
C2929118|T121|1008211|RXNORM|CAFFEINE / CHLORPHENOXAMINE|CAFFEINE / CHLORPHENOXAMINE
C2929117|T121|1008210|RXNORM|ESTRIOL / LACTOBACILLUS ACIDOPHILUS|ESTRIOL / LACTOBACILLUS ACIDOPHILUS
C2929126|T121|1008219|RXNORM|BENZOCAINE / ZINC OXIDE|BENZOCAINE / ZINC OXIDE
C2929125|T121|1008218|RXNORM|PHLOROGLUCINOL / TRIMETHOBENZAMIDE|PHLOROGLUCINOL / TRIMETHOBENZAMIDE
C3833229|T109|1540870|RXNORM|ETHYL METHICONE (8 MPA.S)|ETHYL METHICONE (8 MPA.S)
C0004969|T121|1367|RXNORM|BENCYCLANE|BENCYCLANE
C3833231|T109|1540872|RXNORM|EUCALYPTUS RADIATA FLOWER TOP OIL|EUCALYPTUS RADIATA FLOWER TOP OIL
C3833232|T109|1540873|RXNORM|MEADOWFOAM SEED OIL FATTY ACIDS|MEADOWFOAM SEED OIL FATTY ACIDS
C3833233|T109|1540874|RXNORM|CENTIPEDA MINIMA WHOLE EXTRACT|CENTIPEDA MINIMA WHOLE EXTRACT
C3714575|T109|1540875|RXNORM|PERFLUOROPERHYDROPHENANTHRENE|PERFLUOROPERHYDROPHENANTHRENE
C3833234|T121|1540876|RXNORM|POLYGLYCERYL-4 OLEATE|POLYGLYCERYL-4 OLEATE
C0004962|T121|1361|RXNORM|BENACTYZINE|BENACTYZINE
C3833236|T109|1540878|RXNORM|OCTYLDODECYL BEHENATE|OCTYLDODECYL BEHENATE
C3833237|T109|1540879|RXNORM|UNDECYL ETHYLENEGLYCOL MONOETHER|UNDECYL ETHYLENEGLYCOL MONOETHER
C1095887|T121|319808|RXNORM|BROCCOLI PREPARATION|BROCCOLI PREPARATION
C0004975|T121|1369|RXNORM|BENDROFLUMETHIAZIDE|BENDROFLUMETHIAZIDE
C3709741|T121|1488227|RXNORM|EQUUS CABALLUS LEG CALLOUS PREPARATION|EQUUS CABALLUS LEG CALLOUS PREPARATION
C0717615|T121|214418|RXNORM|CHLORTHALIDONE / CLONIDINE|CHLORTHALIDONE / CLONIDINE
C0717616|T121|214419|RXNORM|CHLORTHALIDONE / RESERPINE|CHLORTHALIDONE / RESERPINE
C3488922|T109|1309336|RXNORM|MANIHOT ESCULENTA ROOT EXTRACT|CASSAVA
C2701641|T129|852551|RXNORM|BURWEED MARSHELDER POLLEN EXTRACT|IVA XANTHIFOLIA POLLEN EXTRACT
C0046547|T109|1358473|RXNORM|2-PYRROLIDONE|2-PYRROLIDONE
C0717608|T121|214411|RXNORM|CHLORPHENIRAMINE / METHSCOPOLAMINE / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / METHSCOPOLAMINE / PHENYLPROPANOLAMINE
C0717613|T121|214416|RXNORM|CHLORPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE|CHLORPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE
C3505482|T121|1358476|RXNORM|CHERRY PLUM EXTRACT|CHERRY PLUM EXTRACT
C3505481|T121|1358475|RXNORM|CEANOTHUS AMERICANUS WHOLE EXTRACT|CEANOTHUS AMERICANUS WHOLE EXTRACT
C3505480|T121|1358474|RXNORM|BERBERIS VULGARIS WHOLE EXTRACT|BERBERIS VULGARIS WHOLE EXTRACT
C0014708|T121|4024|RXNORM|ERGOLOID MESYLATES, USP|ERGOLOID MESYLATES, USP
C0014710|T121|4025|RXNORM|ERGOTAMINE|ERGOTAMINE
C0014707|T123|4023|RXNORM|ERGOT ALKALOIDS|ERGOT ALKALOIDS
C0073571|T121|35780|RXNORM|ROPIVACAINE|ROPIVACAINE
C0014704|T121|4021|RXNORM|ERGONOVINE|ERGONOVINE
C3257224|T121|1241795|RXNORM|CUPRIC OXIDE / FOLIC ACID / NIACINAMIDE / ZINC OXIDE|CUPRIC OXIDE / FOLIC ACID / NIACINAMIDE / ZINC OXIDE
C2701290|T129|852087|RXNORM|SHAD SCALE POLLEN EXTRACT|ATRIPLEX CONFERTIFOLIA POLLEN EXTRACT
C1956630|T121|1432796|RXNORM|PARTHENIUM HYSTEROPHORUS EXTRACT|PARTHENIUM HYSTEROPHORUS EXTRACT
C2929283|T121|1008378|RXNORM|CETYLPYRIDINIUM / DYCLONINE|CETYLPYRIDINIUM / DYCLONINE
C2929284|T121|1008379|RXNORM|LECITHIN / PHOSPHATIDYLETHANOLAMINES / PHOSPHATIDYLINOSITOLS|LECITHIN / PHOSPHATIDYLETHANOLAMINES / PHOSPHATIDYLINOSITOLS
C2929279|T121|1008374|RXNORM|CATALASE / SUPEROXIDE DISMUTASE|CATALASE / SUPEROXIDE DISMUTASE
C2929280|T121|1008375|RXNORM|BENZETHONIUM / LIDOCAINE|BENZETHONIUM / LIDOCAINE
C2929281|T121|1008376|RXNORM|CAMPHOR / PETROLATUM|CAMPHOR / PETROLATUM
C0078221|T129|807219|RXNORM|TYPHOID VI POLYSACCHARIDE VACCINE, S TYPHI TY2 STRAIN|TYPHOID VI POLYSACCHARIDE VACCINE, S TYPHI TY2 STRAIN
C2929275|T121|1008370|RXNORM|AMOXICILLIN / DICLOFENAC|AMOXICILLIN / DICLOFENAC
C2929276|T121|1008371|RXNORM|ATROPINE / SCOPOLAMINE / SIMETHICONE|ATROPINE / SCOPOLAMINE / SIMETHICONE
C2929277|T121|1008372|RXNORM|CITIOLONE / SILYMARIN|CITIOLONE / SILYMARIN
C2929278|T121|1008373|RXNORM|ALUMINUM ACETATE / BORIC ACID|ALUMINUM ACETATE / BORIC ACID
C3256333|T109|1307094|RXNORM|AMNONIUM ACRYLOYLDIMETHYLTAURATE - VP COPOLYMER|AMNONIUM ACRYLOYLDIMETHYLTAURATE - VP COPOLYMER
C0077096|T131|1307097|RXNORM|TRIETHYLAMINE|TRIETHYLAMINE
C3255967|T121|1307096|RXNORM|PEG-12 GLYCERYL DIMYRISTATE|PEG-12 GLYCERYL DIMYRISTATE
C3473405|T121|1307091|RXNORM|HEPTYL UNDECYLENATE|HEPTYL UNDECYLENATE
C3473399|T121|1307090|RXNORM|PENTAERYTHRITYL TETRASTEARATE|PENTAERYTHRITYL TETRASTEARATE
C3255869|T109|1307093|RXNORM|STEARAMIDOPROPYL PG-DIMONIUM CHLORIDE PHOSPHATE|STEARAMIDOPROPYL PROPYLENE GLYCOL-DIMONIUM CHLORIDE PHOSPHATE
C3256543|T109|1307092|RXNORM|ISODECYL NEOPENTANOATE|ISODECYL NEOPENTANOATE
C0069638|T121|32526|RXNORM|ORGOTEIN|ORGOTEIN
C0014582|T121|3995|RXNORM|EPIRUBICIN|EPIRUBICIN
C3256323|T121|1307099|RXNORM|ACETYL TETRAPEPTIDE-9|ACETYL TETRAPEPTIDE-9
C0014563|T125|3992|RXNORM|EPINEPHRINE|EPINEPHRINE
C0014563|T125|3992|RXNORM|EPINEPHRINE|EPINEPHRINE
C0014563|T125|3992|RXNORM|EPINEPHRINE|EPINEPHRINE
C0014563|T125|3992|RXNORM|EPINEPHRINE|EPINEPHRINE
C0014563|T125|3992|RXNORM|EPINEPHRINE|EPINEPHRINE
C0014563|T125|3992|RXNORM|EPINEPHRINE|EPINEPHRINE
C3538274|T121|1372474|RXNORM|AMYLASES / BETAINE / OX BILE EXTRACT / PANCREATIN / PAPAIN / PEPSIN A|AMYLASES / BETAINE / OX BILE EXTRACT / PANCREATIN / PAPAIN / PEPSIN A
C2947386|T121|1041523|RXNORM|ACETIC ACID / ANTIPYRINE / BENZOCAINE / POLICOSANOL|ACETIC ACID / ANTIPYRINE / BENZOCAINE / POLICOSANOL
C3486295|T121|1426702|RXNORM|POLYETHYLENE GLYCOL 300000|POLYETHYLENE GLYCOL 300000
C2727836|T129|999450|RXNORM|EUROTIUM HERBARIORUM EXTRACT|EUROTIUM HERBARIORUM ALLERGENIC EXTRACT
C2701518|T129|852339|RXNORM|ASPEN POLLEN EXTRACT|POPULUS TREMULA POLLEN EXTRACT
C0982180|T121|314647|RXNORM|GLYCERYL MONOLAURATE|GLYCERYL MONOLAURATE
C3499937|T121|1313179|RXNORM|PPG-17|POLYOXYPROPYLENE (17)
C1121677|T121|1313178|RXNORM|PPG-15 STEARYL ETHER|PPG-15 STEARYL ETHER
C3499933|T121|1313173|RXNORM|N,N-DIMETHYLGLYCINE|N,N-DIMETHYLGLYCINE
C3499931|T121|1313171|RXNORM|NONOXYNOL-8|NONOXYNOL-8
C3499936|T121|1313177|RXNORM|PEG-5 GLYCERYL STEARATE|PEG-5 GLYCERYL STEARATE
C0768280|T197|1313176|RXNORM|NICKEL ACETATE|NICKEL ACETATE
C3848535|T196|1546409|RXNORM|TRIPOLYPHOSPHATE ION|TRIPOLYPHOSPHATE ION
C3651721|T130|1430394|RXNORM|BENZILIC ACID|BENZILIC ACID
C3651720|T121|1430397|RXNORM|ACETYLMANDELIC ACID, (+)-|ACETYLMANDELIC ACID, (+)-
C3651722|T109|1430391|RXNORM|ULKENIA DHA OIL|ULKENIA DHA OIL
C2698944|T121|1430390|RXNORM|RACEMENTHOL|RACEMENTHOL
C2079534|T121|815872|RXNORM|BENZYL BENZOATE / PERMETHRIN|BENZYL BENZOATE / PERMETHRIN
C3504704|T121|1356492|RXNORM|SAPINDUS MUKOROSSI FRUIT RIND EXTRACT|SAPINDUS MUKOROSSI FRUIT RIND EXTRACT
C3504703|T121|1356491|RXNORM|PIPERIDINEPROPIONIC ACID|PIPERIDINEPROPIONIC ACID
C3504702|T121|1356490|RXNORM|PEG-60 GLYCERYL ISOSTEARATE|PEG-60 GLYCERYL ISOSTEARATE
C2701435|T129|852237|RXNORM|LAMBS QUARTERS POLLEN EXTRACT|CHENOPODIUM ALBUM POLLEN EXTRACT
C0209210|T121|68091|RXNORM|DOLASETRON|DOLASETRON
C3848553|T196|1546368|RXNORM|CESIUM CATION|CESIUM CATION
C0001443|T123|296|RXNORM|ADENOSINE|ADENOSINE
C0001443|T123|296|RXNORM|ADENOSINE|ADENOSINE
C0772319|T125|1546408|RXNORM|UNOPROSTONE|UNOPROSTONE
C0069937|T121|32786|RXNORM|PADIMATE-O|PADIMATE-O
C0001407|T123|290|RXNORM|ADENINE|ADENINE
C0282340|T130|82097|RXNORM|ROSE BENGAL SODIUM I 131|ROSE BENGAL SODIUM I 131
C3267656|T121|1306058|RXNORM|TRIBULUS TERRESTRIS ROOT EXTRACT|TRIBULUS TERRESTRIS ROOT EXTRACT
C3464669|T195|1306059|RXNORM|TILDIPIROSIN|TILDIPIROSIN
C3474474|T109|1306057|RXNORM|WHITE PINE OIL|WHITE PINE OIL
C0351000|T121|102848|RXNORM|GLYMIDINE|GLYMIDINE
C1719877|T121|645364|RXNORM|ALUMINUM HYDROXIDE / DIMETHICONE|ALUMINUM HYDROXIDE / DIMETHICONE
C0654934|T121|1426854|RXNORM|AMILOXATE|AMILOXATE
C0060493|T121|25112|RXNORM|FLUMEQUINE|FLUMEQUINE
C0350998|T121|102846|RXNORM|GLIBORNURIDE|GLIBORNURIDE
C3163347|T121|1116106|RXNORM|CHLORHEXIDINE / MICONAZOLE|CHLORHEXIDINE / MICONAZOLE
C2702425|T129|867284|RXNORM|PHOMA EXIGUA VAR. EXIGUA EXTRACT|PHOMA EXIGUA VAR. EXIGUA EXTRACT
C0116832|T121|1546423|RXNORM|ETHYL SALICYLATE|ETHYL SALICYLATE
C0085994|T123|42588|RXNORM|CHENODEOXYCHOLATE|CHENODEOXYCHOLATE
C3154678|T121|1102195|RXNORM|ASCORBIC ACID / BIOTIN / FERROUS BISGLYCINATE / FOLIC ACID / FORMIC ACID / IRON-DEXTRAN COMPLEX / NIACIN / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|ASCORBIC ACID / BIOTIN / FERROUS BISGLYCINATE / FOLIC ACID / FORMIC ACID / IRON-DEXTRAN COMPLEX / NIACIN / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C3813541|T121|1535496|RXNORM|POLYGONUM ARENASTRUM WHOLE EXTRACT|POLYGONUM ARENASTRUM WHOLE EXTRACT
C3818707|T121|1535497|RXNORM|STEMONA SESSILIFOLIA ROOT EXTRACT|STEMONA SESSILIFOLIA ROOT EXTRACT
C3818709|T109|1535494|RXNORM|LOTUS CORNICULATUS FLOWER VOLATILE OIL|LOTUS CORNICULATUS FLOWER VOLATILE OIL
C3818708|T121|1535495|RXNORM|PEUCEDANUM PRAERUPTORUM ROOT EXTRACT|PEUCEDANUM PRAERUPTORUM ROOT EXTRACT
C3474073|T121|1358899|RXNORM|HOUTTUYNIA CORDATA WHOLE EXTRACT|HOUTTUYNIA CORDATA WHOLE EXTRACT
C0008402|T121|2447|RXNORM|CHOLESTYRAMINE RESIN|CHOLESTYRAMINE RESIN
C3818713|T121|1535490|RXNORM|GLYCYRRHIZA GLABRA WHOLE EXTRACT|GLYCYRRHIZA GLABRA WHOLE EXTRACT
C3818712|T121|1535491|RXNORM|GLYCYRRHIZA URALENSIS WHOLE EXTRACT|GLYCYRRHIZA URALENSIS WHOLE EXTRACT
C3474071|T121|1358895|RXNORM|DIANTHUS CHINENSIS WHOLE EXTRACT|DIANTHUS CHINENSIS WHOLE EXTRACT
C3256843|T109|1358897|RXNORM|GRAPEFRUIT PEEL EXTRACT|GRAPEFRUIT PEEL EXTRACT
C0008405|T123|2449|RXNORM|CHOLINE|CHOLINE
C0008405|T123|2449|RXNORM|CHOLINE|CHOLINE
C3489061|T121|1358891|RXNORM|THUJA OCCIDENTALIS WHOLE EXTRACT|THUJA OCCIDENTALIS WHOLE EXTRACT
C3257275|T121|1241895|RXNORM|NIACIN / PANTOTHENIC ACID / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN B6|NIACIN / PANTOTHENIC ACID / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN B6
C3488680|T121|1358893|RXNORM|SOLANUM NIGRUM WHOLE EXTRACT|SOLANUM NIGRUM WHOLE EXTRACT
C3485018|T121|1358892|RXNORM|SYZYGIUM AROMATICUM WHOLE EXTRACT|SYZYGIUM AROMATICUM WHOLE EXTRACT
C0004599|T195|1291|RXNORM|ASCORBIC ACID / CRANBERRY PREPARATION / LACTOBACILLUS SPOROGENES|BACITRACIN
C0041455|T123|1426856|RXNORM|COLLAGEN TYPE I|COLLAGEN TYPE I
C3818700|T121|1535944|RXNORM|COAGULATION FACTOR IX RECOMBINANT IMMUNOGLOBULIN G1 FUSION PROTEIN|EFTRENONACOG ALFA
C2930030|T121|1009135|RXNORM|PENBUTOLOL / PIRETANIDE|PENBUTOLOL / PIRETANIDE
C0050559|T121|16818|RXNORM|ACITRETIN|ACITRETIN
C2930032|T121|1009137|RXNORM|AMILORIDE / BENDROFLUMETHIAZIDE|AMILORIDE / BENDROFLUMETHIAZIDE
C2930031|T121|1009136|RXNORM|PAPAIN / PAPAYA PREPARATION|PAPAIN / PAPAYA PREPARATION
C2930026|T121|1009131|RXNORM|ATROPINE / ICTASOL|ATROPINE / ICTASOL
C2930025|T121|1009130|RXNORM|BEE POLLEN / ROYAL JELLY|BEE POLLEN / ROYAL JELLY
C2930028|T121|1009133|RXNORM|PHENYLEPHRINE / SULFATED MUCOPOLYSACCHARIDES|PHENYLEPHRINE / SULFATED MUCOPOLYSACCHARIDES
C2929318|T121|1008414|RXNORM|CHLOROCRESOL / CLOROPHENE|CHLOROCRESOL / CLOROPHENE
C3505487|T121|1358481|RXNORM|VITIS VINIFERA WHOLE EXTRACT|VITIS VINIFERA WHOLE EXTRACT
C2930034|T121|1009139|RXNORM|HYDRALAZINE / HYDROCHLOROTHIAZIDE / METOPROLOL|HYDRALAZINE / HYDROCHLOROTHIAZIDE / METOPROLOL
C2930033|T121|1009138|RXNORM|HYALURONATE / PILOCARPINE|HYALURONATE / PILOCARPINE
C0050558|T121|16817|RXNORM|ACIPIMOX|ACIPIMOX
C0023586|T121|6378|RXNORM|LEVORPHANOL|LEVORPHANOL
C0771395|T121|236149|RXNORM|AMYL SALICYLATE|AMYL SALICYLATE
C0023554|T121|6370|RXNORM|LEVALLORPHAN|LEVALLORPHAN
C0023556|T121|6371|RXNORM|LEVAMISOLE|LEVAMISOLE
C0771387|T121|236142|RXNORM|ZINC ASPARTATE|ZINC ASPARTATE
C0023566|T125|6373|RXNORM|LEVONORGESTREL|LEVONORGESTREL
C0023570|T123|6375|RXNORM|LEVODOPA|LEVODOPA
C2347816|T196|1546419|RXNORM|COBALTOUS CATION|COBALTOUS CATION
C1875264|T121|689920|RXNORM|HYDROCORTISONE / POLYMYXIN B|HYDROCORTISONE / POLYMYXIN B
C0009975|T121|2839|RXNORM|COPPER GLUCONATE|COPPER GLUCONATE
C1875265|T121|689922|RXNORM|HYDROCORTISONE / SALICYLIC ACID / SULFUR|HYDROCORTISONE / SALICYLIC ACID / SULFUR
C1875266|T121|689923|RXNORM|HYDROCORTISONE / SULFUR / ZINC OXIDE|HYDROCORTISONE / SULFUR / ZINC OXIDE
C1874791|T121|689299|RXNORM|CHLOROPHYLL / PAPAIN / UREA|CHLOROPHYLL / PAPAIN / UREA
C1875270|T121|689929|RXNORM|HYDROGEN PEROXIDE / POVIDONE-IODINE|HYDROGEN PEROXIDE / POVIDONE-IODINE
C2741531|T129|901365|RXNORM|CUMIN ALLERGENIC EXTRACT|CUMINUM CYMINUM ALLERGENIC EXTRACT
C3256822|T109|1427045|RXNORM|ETHYLENE-VINYL ACETATE COPOLYMER (9% VINYL ACETATE)|ETHYLENE-VINYL ACETATE COPOLYMER (9% VINYL ACETATE)
C0036579|T121|9639|RXNORM|SELEGILINE|SELEGILINE
C0036579|T121|9639|RXNORM|SELEGILINE|SELEGILINE
C3257534|T109|1427046|RXNORM|WHEAT BRAN EXTRACT|TRITICUM VULGARE EXTRACT
C0112317|T195|1358488|RXNORM|DANOFLOXACIN|DANOFLOXACIN
C3475125|T121|1427043|RXNORM|PEG-PPG-36-41 DIMETHYL ETHER|PEG-PPG-36-41 DIMETHYL ETHER
C3484813|T121|1427042|RXNORM|SUCROSE STEARATE-PALMITATE ESTER (75% MONO ESTER)|SUCROSE STEARATE-PALMITATE ESTER (75% MONO ESTER)
C0058291|T109|1427048|RXNORM|DIMYRISTOYLPHOSPHATIDYLGLYCEROL|DIMYRISTOYLPHOSPHATIDYLGLYCEROL
C3535627|T121|1370729|RXNORM|ANGELICA SINENSIS WHOLE EXTRACT|ANGELICA SINENSIS WHOLE EXTRACT
C2744711|T109|1370728|RXNORM|SUCROSE COCOATE|SUCROSE COCOATE
C1445691|T121|466457|RXNORM|FLUORESCEIN / PROPARACAINE|FLUORESCEIN / PROPARACAINE
C2827132|T121|1546417|RXNORM|DENATONIUM|DENATONIUM
C0001134|T197|236|RXNORM|NA PHOSPHATE,DIBASIC DIHYDRATE|ACIDULATED PHOSPHATE FLUORIDE
C1445687|T121|466453|RXNORM|BROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE|BROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE
C0034131|T130|8948|RXNORM|PURIFIED PROTEIN DERIVATIVE OF TUBERCULIN|PURIFIED PROTEIN DERIVATIVE OF TUBERCULIN
C1445693|T121|466459|RXNORM|GLUCOSAMINE / METHYLSULFONYLMETHANE|GLUCOSAMINE / METHYLSULFONYLMETHANE
C1654082|T121|1486501|RXNORM|BARIUM ACETATE|BARIUM ACETATE
C2928617|T121|1007701|RXNORM|CHYMOSIN / LACTASE|CHYMOSIN / LACTASE
C3848533|T121|1546412|RXNORM|MORINDA OFFICIANALIS ROOT EXTRACT|MORINDA OFFICIANALIS ROOT EXTRACT
C3848532|T121|1546413|RXNORM|METHYLHOMATROPINE|METHYLHOMATROPINE
C0005116|T121|1436|RXNORM|BEPRIDIL|BEPRIDIL
C2702406|T129|891676|RXNORM|STRING BEAN ALLERGENIC EXTRACT|STRING BEAN ALLERGENIC EXTRACT
C0005117|T121|1437|RXNORM|BERBERINE|BERBERINE
C0961965|T121|1491625|RXNORM|METRELEPTIN|METRELEPTIN
C0000956|T121|154|RXNORM|STRONTIUM CATION SR-89|ACENOCOUMAROL
C0287262|T131|83586|RXNORM|LUFENURON|LUFENURON
C3538155|T121|1372271|RXNORM|CHINESE CHESTNUT EXTRACT|CHINESE CHESTNUT EXTRACT
C0005740|T195|1622|RXNORM|BLEOMYCIN|BLEOMYCIN
C0006931|T121|1992|RXNORM|CAPSAICIN|CAPSAICIN
C0006931|T121|1992|RXNORM|CAPSAICIN|CAPSAICIN
C3256649|T109|1305659|RXNORM|SALIX ALBA BARK VOLATILE OIL|SALIX ALBA BARK VOLATILE OIL
C2348197|T109|1305658|RXNORM|SHEANUT OIL|SHEANUT OIL
C2979418|T121|1090831|RXNORM|ASCORBIC ACID / BETA CAROTENE / COPPER SULFATE / LUTEIN / SELENITE / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / BETA CAROTENE / COPPER SULFATE / LUTEIN / SELENITE / VITAMIN E / ZINC OXIDE
C0006945|T121|1999|RXNORM|CARBACHOL|CARBACHOL
C0006938|T121|1998|RXNORM|CAPTOPRIL|CAPTOPRIL
C0260069|T109|1305657|RXNORM|SPEARMINT OIL|SPEARMINT OIL
C3486324|T109|1305656|RXNORM|STAR ANISE OIL|STAR ANISE OIL
C0105754|T109|1305651|RXNORM|BERGAMOT OIL|BERGAMOT OIL
C3265531|T109|1305650|RXNORM|BAY LEAF OIL|BAY LEAF OIL
C1572635|T109|1305653|RXNORM|WORMWOOD OIL|WORMWOOD OIL
C3256128|T109|1305652|RXNORM|BOSWELLIA SERRATA RESIN OIL|BOSWELLIA SERRATA RESIN OIL
C0982275|T129|314724|RXNORM|MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP W-135|MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP W-135
C3500835|T109|1356135|RXNORM|GINKO BILOBA LEAF OIL|GINKO BILOBA LEAF OIL
C3700898|T121|1486502|RXNORM|ILEX AQUIFOLIUM FRUITING TOP EXTRACT|ILEX AQUIFOLIUM FRUITING TOP EXTRACT
C0066477|T121|29961|RXNORM|METYLPERON|MELPERONE
C0064567|T121|28381|RXNORM|AMINO ACIDS 20%|LACHESINE
C3256202|T121|1356138|RXNORM|LAURAMIDOPROPYLAMINE OXIDE|LAURAMIDOPROPYLAMINE OXIDE
C0031479|T121|8167|RXNORM|PHENYLHYDRAZINE|PHENYLHYDRAZINE
C2356380|T121|804304|RXNORM|CALAMINE / PRAMOXINE|CALAMINE / PRAMOXINE
C2928747|T121|1007832|RXNORM|DEXCHLORPHENIRAMINE / METHSCOPOLAMINE / PSEUDOEPHEDRINE|DEXCHLORPHENIRAMINE / METHSCOPOLAMINE / PSEUDOEPHEDRINE
C2928748|T121|1007833|RXNORM|RIBOFLAVIN / VITAMIN B6|RIBOFLAVIN / VITAMIN B6
C0004057|T121|1191|RXNORM|ASPIRIN|ASPIRIN
C0004057|T121|1191|RXNORM|ASPIRIN|ASPIRIN
C0004057|T121|1191|RXNORM|ASPIRIN|ASPIRIN
C0004057|T121|1191|RXNORM|ASPIRIN|ASPIRIN
C0770624|T122|235535|RXNORM|CARBOMER|CARBOMER
C0012066|T121|3347|RXNORM|DICHLOROACETATE|DICHLOROACETATE
C3256690|T121|1307879|RXNORM|JASMINUM OFFICINALE FLOWER EXTRACT|JASMINUM OFFICINALE FLOWER EXTRACT
C2928746|T121|1007831|RXNORM|ASCORBIC ACID / FERROUS GLUCONATE / FOLIC ACID|ASCORBIC ACID / FERROUS GLUCONATE / FOLIC ACID
C0066837|T121|30257|RXNORM|MOXONIDINE|MOXONIDINE
C2928306|T121|1007384|RXNORM|PIROXICAM / VITAMIN B 12|PIROXICAM / VITAMIN B 12
C2241628|T121|802519|RXNORM|ALISKIREN / HYDROCHLOROTHIAZIDE|ALISKIREN / HYDROCHLOROTHIAZIDE
C0059726|T109|1362891|RXNORM|ETHOHEXADIOL|ETHOHEXADIOL
C2365117|T130|1367088|RXNORM|OFTASCEINE|OFTASCEINE
C3859161|T109|1592264|RXNORM|SODIUM LAURETH-4 PHOSPHATE|SODIUM LAURETH-4 PHOSPHATE
C2983890|T121|1336135|RXNORM|SACCHAROMYCES CEREVISIAE RNA|SACCHAROMYCES CEREVISIAE RNA
C3535893|T121|1370587|RXNORM|MYRISTALKONIUM|MYRISTALKONIUM
C0015506|T123|4257|RXNORM|FACTOR VIII|FACTOR VIII
C0015506|T123|4257|RXNORM|FACTOR VIII|FACTOR VIII
C0015505|T126|4256|RXNORM|FACTOR VIIA|FACTOR VIIA
C0015505|T126|4256|RXNORM|FACTOR VIIA|FACTOR VIIA
C3538371|T121|1372641|RXNORM|CHINESE YAM EXTRACT|CHINESE YAM EXTRACT
C0020352|T121|5531|RXNORM|HETASTARCH|HYDROXYETHYLSTARCH
C3535894|T121|1370586|RXNORM|GLYCYRRHIZATE|GLYCYRRHIZATE
C0962603|T121|299635|RXNORM|ALEFACEPT|ALEFACEPT
C0063779|T121|27748|RXNORM|IODOFORM|IODOFORM
C3535899|T121|1370581|RXNORM|2-SULFOLAURATE|2-SULFOLAURATE
C1302124|T121|392564|RXNORM|ACEBUTOLOL / HYDROCHLOROTHIAZIDE|ACEBUTOLOL / HYDROCHLOROTHIAZIDE
C3535900|T121|1370580|RXNORM|LAUROYL ASPARTATE|LAUROYL ASPARTATE
C3488952|T129|1313274|RXNORM|INFLUENZA B VIRUS, B PANAMA-45-90 HEMMAGGLUTININ ANTIGEN, INACTIVATED|INFLUENZA B VIRUS, B PANAMA-45-90 HEMMAGGLUTININ ANTIGEN, INACTIVATED
C3700896|T109|1486507|RXNORM|CALOPHYLLUM TACAMAHACA WHOLE EXTRACT|CALOPHYLLUM TACAMAHACA WHOLE EXTRACT
C2928754|T121|1007839|RXNORM|CHLOROBUTANOL / TANNIC ACID|CHLOROBUTANOL / TANNIC ACID
C0358975|T121|106928|RXNORM|BETAMETHASONE / CLOTRIMAZOLE|BETAMETHASONE / CLOTRIMAZOLE
C2983955|T129|1318050|RXNORM|INTERLEUKIN-12, HUMAN|INTERLEUKIN-12, HUMAN
C3256512|T109|1426384|RXNORM|C12-20 ALKYL BENZOATE|C12-20 ALKYL BENZOATE
C3256402|T109|1424651|RXNORM|BETA-D-GALACTOPYRANOSE|BETA-D-GALACTOPYRANOSE
C3256400|T109|1424650|RXNORM|BETA-CITRONELLOL, (+-)-|BETA-CITRONELLOL, (+-)-
C3535898|T121|1370582|RXNORM|P-CHLORO-M-CRESOL|P-CHLORO-M-CRESOL
C1679366|T109|1424655|RXNORM|1,2-DIMYRISTOYL-SN-GLYCERO-3-(PHOSPHO-RAC-(1-GLYCEROL))|1,2-DIMYRISTOYL-SN-GLYCERO-3-(PHOSPHO-RAC-(1-GLYCEROL))
C3256405|T109|1424656|RXNORM|1,2-DIOLEOYL-SN-GLYCERO-3-PHOSPHOCHOLINE|1,2-DIOLEOYL-SN-GLYCERO-3-PHOSPHOCHOLINE
C1872109|T129|709271|RXNORM|CERTOLIZUMAB PEGOL|CERTOLIZUMAB PEGOL
C3486609|T121|1309808|RXNORM|FERULA SUMBUL ROOT EXTRACT|FERULA SUMBUL ROOT EXTRACT
C3488357|T121|1309809|RXNORM|MALUS DOMESTICA FLOWER EXTRACT|MALUS DOMESTICA FLOWER EXTRACT
C3486686|T121|1426873|RXNORM|HEKLA LAVA|HEKLA LAVA
C3486608|T121|1309805|RXNORM|ASCLEPIAS TUBEROSA FLOWERING TOP EXTRACT|ASCLEPIAS TUBEROSA FLOWERING TOP EXTRACT
C3255602|T121|1309806|RXNORM|LIGUSTICUM TENUISSIMUM LEAF EXTRACT|LIGUSTICUM TENUISSIMUM LEAF EXTRACT
C3488342|T121|1309807|RXNORM|CYNANCHUM VINCETOXICUM ROOT EXTRACT|VINCETOXICUM HIRUNDINARIA ROOT EXTRACT
C3486603|T121|1309800|RXNORM|ARUNDO PLINIANA ROOT EXTRACT|ARUNDO PLINIANA ROOT EXTRACT
C0050408|T121|1426875|RXNORM|ACEMANNAN|ACEMANNAN
C3255601|T121|1309803|RXNORM|LIGUSTICUM SINENSE SUBSP. CHUANXIONG ROOT EXTRACT|LIGUSTICUM SINENSE SUBSP. CHUANXIONG ROOT EXTRACT
C3819183|T121|1490716|RXNORM|COENZYME Q10 / GLYCINE / ISOLEUCINE|COENZYME Q10 / GLYCINE / ISOLEUCINE
C0301408|T121|89811|RXNORM|VINBARBITAL|VINBARBITAL
C0301407|T121|89810|RXNORM|TALBUTAL|TALBUTAL
C0301409|T121|89812|RXNORM|CAPTODIAMINE|CAPTODIAME
C1996229|T121|834773|RXNORM|BROMPHENIRAMINE / DIPHENHYDRAMINE|BROMPHENIRAMINE / DIPHENHYDRAMINE
C0301418|T121|89818|RXNORM|STYRAMATE|STYRAMATE
C1136535|T129|338036|RXNORM|PEGFILGRASTIM|PEGFILGRASTIM
C2001856|T121|1302966|RXNORM|CARFILZOMIB|CARFILZOMIB
C0123859|T121|51471|RXNORM|IODOXAMID|IODOXAMID
C2739885|T129|897316|RXNORM|SALTBUSH POLLEN EXTRACT|ATRIPLEX WRIGHTII POLLEN EXTRACT
C0123865|T130|51474|RXNORM|IOTROLAN|IOTROLAN
C1952576|T121|729717|RXNORM|METFORMIN / SITAGLIPTIN|METFORMIN / SITAGLIPTIN
C0107103|T123|47324|RXNORM|BRAIN-DERIVED NEUROTROPHIC FACTOR|BRAIN-DERIVED NEUROTROPHIC FACTOR
C3848597|T109|1545167|RXNORM|N-TERT-OCTYLACRYLAMIDE|N-TERT-OCTYLACRYLAMIDE
C0072828|T121|35185|RXNORM|QUAZEPAM|QUAZEPAM
C0024452|T195|6572|RXNORM|MAFENIDE|MAFENIDE
C2928499|T121|1007579|RXNORM|CALCIUM ASCORBATE / POTASSIUM|CALCIUM ASCORBATE / POTASSIUM
C2928498|T121|1007578|RXNORM|BENZOCAINE / ZIRCONIUM OXIDE|BENZOCAINE / ZIRCONIUM OXIDE
C0024467|T196|6574|RXNORM|MAGNESIUM|MAGNESIUM
C2928493|T121|1007573|RXNORM|FOLIC ACID / VITAMIN B 12|FOLIC ACID / VITAMIN B 12
C2928493|T121|1007573|RXNORM|FOLIC ACID / VITAMIN B 12|FOLIC ACID / VITAMIN B 12
C2928492|T121|1007572|RXNORM|ACETAMINOPHEN / CODEINE / GUAIFENESIN / PSEUDOEPHEDRINE|ACETAMINOPHEN / CODEINE / GUAIFENESIN / PSEUDOEPHEDRINE
C2928491|T121|1007571|RXNORM|CALCIUM PHOSPHATE / CHOLECALCIFEROL / SOYBEAN PREPARATION|CALCIUM PHOSPHATE / CHOLECALCIFEROL / SOYBEAN PREPARATION
C0024472|T197|6579|RXNORM|MAGNESIUM CHLORIDE|MAGNESIUM CHLORIDE
C1608841|T129|847083|RXNORM|USTEKINUMAB|USTEKINUMAB
C2928496|T121|1007576|RXNORM|LIDOCAINE / POLYMYXIN B|LIDOCAINE / POLYMYXIN B
C2928495|T121|1007575|RXNORM|DOMPERIDONE / RANITIDINE|DOMPERIDONE / RANITIDINE
C2928494|T121|1007574|RXNORM|THIAMINE / VITAMIN B 12|THIAMINE / VITAMIN B 12
C0249959|T121|73891|RXNORM|BLACK CURRANT OIL|BLACK CURRANT OIL
C1874687|T121|691178|RXNORM|CAMPHOR / EUCALYPTUS OIL / MENTHOL|CAMPHOR / EUCALYPTUS OIL / MENTHOL
C0771875|T121|236583|RXNORM|MITE EXTRACT|MITE EXTRACT
C2730258|T129|892674|RXNORM|BAKER'S YEAST ALLERGENIC EXTRACT|BAKER'S YEAST ALLERGENIC EXTRACT
C0982390|T121|314832|RXNORM|SODIUM LAURYL SULFOACETATE|SODIUM LAURYL SULFOACETATE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, HICKORY|PRASTERONE
C2698764|T121|1356552|RXNORM|PERAMPANEL|PERAMPANEL
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, HORMODENDRUM HORDEI|PRASTERONE
C0982396|T197|314838|RXNORM|SODIUM PHOSPHATE, DIBASIC, ANHYDROUS|SODIUM PHOSPHATE, DIBASIC, ANHYDROUS
C0145184|T121|57047|RXNORM|TERIZIDONE|TERIZIDONE
C2701613|T129|852509|RXNORM|SUNFLOWER POLLEN EXTRACT|HELIANTHUS ANNUUS POLLEN EXTRACT
C1165931|T121|350255|RXNORM|HEPATITIS NOSODES|HEPATITIS NOSODES
C3555540|T197|1373351|RXNORM|SILODRATE|SILODRATE
C3535891|T121|1370590|RXNORM|DIHYDROXYPROPYLTRIMONIUM|DIHYDROXYPROPYLTRIMONIUM
C2605143|T121|1366947|RXNORM|2-NAPHTHALENESULFONATE|2-NAPHTHALENESULFONATE
C0813171|T121|258326|RXNORM|ST. JOHN'S WORT EXTRACT|HYPERICI HERBA
C0220795|T121|70589|RXNORM|BENZOATE|BENZOATE
C3538575|T121|1373114|RXNORM|IODOFORM / ZINC OXIDE|IODOFORM / ZINC OXIDE
C0104238|T197|1375924|RXNORM|ARSENATE|ARESENATE ION
C3486691|T121|1313342|RXNORM|FAGUS SYLVATICA NUT EXTRACT|FAGUS SYLVATICA NUT EXTRACT
C0060515|T197|1313343|RXNORM|FLUORAPATITE|FLUORAPATITE
C0058217|T131|1313349|RXNORM|DIMETHYL ETHER|DIMETHYL ETHER
C1875645|T121|689737|RXNORM|PHENAZOPYRIDINE / SULFAMETHIZOLE|PHENAZOPYRIDINE / SULFAMETHIZOLE
C0001655|T125|376|RXNORM|CORTICOTROPIN|CORTICOTROPIN
C1875160|T121|687351|RXNORM|FLUOCINOLONE / NEOMYCIN|FLUOCINOLONE / NEOMYCIN
C0069370|T121|32311|RXNORM|OCTYLONIUM|OCTYLONIUM
C0069772|T121|32645|RXNORM|OXIRACETAM|OXIRACETAM
C0164398|T121|59639|RXNORM|ATOSIBAN|ATOSIBAN
C3709739|T121|1488225|RXNORM|SUS SCROFA FALLOPIAN TUBE PREPARATION|SUS SCROFA FALLOPIAN TUBE PREPARATION
C0053116|T127|18891|RXNORM|BENPHOTHIAMINE|BENPHOTHIAMINE
C0069776|T121|32649|RXNORM|OXITROPIUM|OXITROPIUM
C3651758|T109|1428862|RXNORM|BUTYLENE GLYCOL DICAPRATE|BUTYLENE GLYCOL DICAPRATE
C0022635|T121|6142|RXNORM|KETOPROFEN|KETOPROFEN
C0772233|T197|236907|RXNORM|POTASSIUM SULFIDE|POTASSIUM SULFIDE
C0022643|T121|6147|RXNORM|KHELLIN|KHELLIN
C0022642|T121|6146|RXNORM|KETOTIFEN|KETOTIFEN
C0044052|T130|1428547|RXNORM|1,6-HEXAMETHYLENE DIISOCYANATE|1,6-HEXAMETHYLENE DIISOCYANATE
C1453642|T195|473837|RXNORM|TELAVANCIN|TELAVANCIN
C0137996|T121|54993|RXNORM|POTASSIUM CITRATE|POTASSIUM CITRATE
C0050505|T130|1425216|RXNORM|ACETYLCELLULOSE|CELLULOSE ACETATE
C0041536|T123|10975|RXNORM|UBIQUINONE|UBIQUINONE
C3162427|T121|1425214|RXNORM|CAVIAR PREPARATION|CAVIAR PREPARATION
C0055049|T122|1425215|RXNORM|CELLULOSE ACETATE PHTHALATE|CELLACEFATE
C0145185|T125|57048|RXNORM|TERLIPRESSIN|TERLIPRESSIN
C0971350|T121|1425218|RXNORM|CETEARYL ALCOHOL|CETEARYL ALCOHOL
C2717318|T109|1425219|RXNORM|CETEARYL GLUCOSIDE|CETEARYL GLUCOSIDE
C2194188|T121|816394|RXNORM|ASCORBIC ACID / CALCIUM ASCORBATE|ASCORBIC ACID / CALCIUM ASCORBATE
C3651732|T121|1429948|RXNORM|POLYGALA TENUIFOLIA ROOT EXTRACT|POLYGALA TENUIFOLIA ROOT EXTRACT
C3834048|T109|1543741|RXNORM|PEG-90 STEARATE|PEG-90 STEARATE
C3651733|T121|1429943|RXNORM|METHACRYLATE-METHOXY PEG-10 MALEATE-STYRENE COPOLYMER|METHACRYLATE-METHOXY PEG-10 MALEATE-STYRENE COPOLYMER
C0055735|T130|21113|RXNORM|CINAMETIC ACID|CINAMETIC ACID
C1566826|T121|1102270|RXNORM|RILPIVIRINE|RILPIVIRINE
C0022940|T007|1592255|RXNORM|LACTOBACILLUS CASEI|LACTOBACILLUS CASEI
C0772234|T121|236908|RXNORM|METHYL BUTETISALICYLATE|METHYL BUTETISALICYLATE
C3257788|T121|1242956|RXNORM|BURWEED MARSHELDER POLLEN EXTRACT / POVERTY WEED POLLEN EXTRACT / ROUGH MARSHELDER POLLEN EXTRACT|BURWEED MARSHELDER POLLEN EXTRACT / POVERTY WEED POLLEN EXTRACT / ROUGH MARSHELDER POLLEN EXTRACT
C1629853|T121|608571|RXNORM|LIDOCAINE / ZINC OXIDE|LIDOCAINE / ZINC OXIDE
C0057610|T127|22701|RXNORM|DEXPANTHENOL|(+)-PANTHENOL
C0057610|T127|22701|RXNORM|DEXPANTHENOL|(+)-PANTHENOL
C1445834|T121|466600|RXNORM|CAMPHOR / MENTHOL|CAMPHOR / MENTHOL
C1445834|T121|466600|RXNORM|CAMPHOR / MENTHOL|CAMPHOR / MENTHOL
C0717531|T121|214336|RXNORM|CAFFEINE / ERGOTAMINE|CAFFEINE / ERGOTAMINE
C0057621|T121|22708|RXNORM|DEXTRANOMER|DEXTRANOMER
C0057621|T121|22708|RXNORM|DEXTRANOMER|DEXTRANOMER
C0061751|T121|26143|RXNORM|GLYCYRRHIZIC ACID|GLYCYRRHIZIC ACID
C1874812|T121|689389|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE|CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE
C3864971|T121|1596423|RXNORM|IODINE / ISOPROPYL ALCOHOL / SODIUM IODIDE|IODINE / ISOPROPYL ALCOHOL / SODIUM IODIDE
C1170397|T121|352767|RXNORM|METHSCOPOLAMINE / PSEUDOEPHEDRINE|METHSCOPOLAMINE / PSEUDOEPHEDRINE
C0216784|T121|69749|RXNORM|VALSARTAN|VALSARTAN
C3538361|T121|1372631|RXNORM|PIGMENT RED 5|PIGMENT RED 5
C2725260|T121|1482502|RXNORM|ESLICARBAZEPINE|ESLICARBAZEPINE
C1329988|T121|404783|RXNORM|CARBETAPENTANE / PSEUDOEPHEDRINE|CARBETAPENTANE / PSEUDOEPHEDRINE
C3255838|T109|1306197|RXNORM|ACORUS GRAMINEUS ROOT EXTRACT|ACORUS GRAMINEUS ROOT EXTRACT
C0051601|T121|46276|RXNORM|AMINAPHTHONE|AMINAPHTHONE
C2981355|T109|1426435|RXNORM|POLYOXYL 50 HYDROGENATED CASTOR OIL|PEG-50 HYDROGENATED CASTOR OIL
C3669357|T121|1482787|RXNORM|HYSSOPUS OFFICINALIS WHOLE EXTRACT|HYSSOPUS OFFICINALIS WHOLE EXTRACT
C3695989|T121|1482786|RXNORM|PPG-2 HYDROXYETHYL STEARAMIDE|PPG-2 HYDROXYETHYL STEARAMIDE
C2744563|T195|1368469|RXNORM|TYLVALOSIN|TYLVALOSIN
C1874807|T121|689381|RXNORM|CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C3695987|T121|1482789|RXNORM|CORDIA SEBESTENA FLOWER EXTRACT|CORDIA SEBESTENA FLOWER EXTRACT
C3695988|T121|1482788|RXNORM|CISTUS INCANUS FLOWERING TOP EXTRACT|CISTUS INCANUS FLOWERING TOP EXTRACT
C0007047|T121|2051|RXNORM|CARBOPROST|CARBOPROST
C0039943|T121|10502|RXNORM|THIORIDAZINE|THIORIDAZINE
C3485471|T121|1368159|RXNORM|ISOCETYL ETHYLHEXANOATE|ISOCETYL ETHYLHEXANOATE
C3474293|T121|1368158|RXNORM|QUATERNIUM-91|QUATERNIUM-91
C0016564|T131|4530|RXNORM|FORMALDEHYDE|FORMALDEHYDE
C0016564|T131|4530|RXNORM|FORMALDEHYDE|FORMALDEHYDE
C0017642|T121|4821|RXNORM|GLIPIZIDE|GLIPIZIDE
C0030827|T195|7980|RXNORM|PENICILLIN G|PENICILLIN G
C0353942|T168|104125|RXNORM|BRAN|BRAN
C0030840|T195|7984|RXNORM|PENICILLIN V|PENICILLIN V
C3848543|T196|1546390|RXNORM|CHLORATE ION|CHLORATE ION
C2741586|T129|901507|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP C OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|NEISSERIA MENINGITIDIS SEROGROUP C OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C0040341|T195|10627|RXNORM|TOBRAMYCIN|TOBRAMYCIN
C0040341|T195|10627|RXNORM|TOBRAMYCIN|TOBRAMYCIN
C0040341|T195|10627|RXNORM|TOBRAMYCIN|TOBRAMYCIN
C0070455|T131|33199|RXNORM|PERMETHRIN|PERMETHRIN
C3696419|T121|1484782|RXNORM|MICONAZOLE / SALICYLIC ACID|MICONAZOLE / SALICYLIC ACID
C0772125|T121|236809|RXNORM|GINKGO BILOBA EXTRACT|GINKGO BILOBA EXTRACT
C2702362|T129|892665|RXNORM|COW MILK ALLERGENIC EXTRACT|COW MILK ALLERGENIC EXTRACT
C0772117|T121|236801|RXNORM|YOHIMBE BARK PREPARATION|YOHIMBE BARK PREPARATION
C0772118|T121|236802|RXNORM|DAMIANA EXTRACT|DAMIANA EXTRACT
C0026408|T195|1368208|RXNORM|MONENSIN|MONENSIN
C3535693|T121|1368151|RXNORM|CHELIDONIUM MAJUS ROOT EXTRACT|CHELIDONIUM MAJUS ROOT EXTRACT
C0440463|T121|124431|RXNORM|YELLOW HORNET VENOM|YELLOW HORNET VENOM
C0106916|T121|1368202|RXNORM|BORNEOL|BORNEOL
C0057874|T121|1368201|RXNORM|DICLAZURIL|DICLAZURIL
C3255839|T109|1306198|RXNORM|AMMONIO METHACRYLATE COPOLYMER TYPE B|AMMONIO METHACRYLATE COPOLYMER TYPE B
C2827258|T121|1368207|RXNORM|MENTHYL SALICYLATE|MENTHYL SALICYLATE
C3472792|T121|1368206|RXNORM|LENTINULA EDODES MYCELIUM EXTRACT|LENTINULA EDODES MYCELIUM EXTRACT
C3485560|T121|1368205|RXNORM|BETA VULGARIS EXTRACT|BETA VULGARIS EXTRACT
C3535921|T123|1368204|RXNORM|BEHENATE|BEHENATE
C3692999|T121|1442993|RXNORM|HYOSCYAMUS NIGER WHOLE EXTRACT|HYOSCYAMUS NIGER WHOLE EXTRACT
C3485069|T121|1310063|RXNORM|FRANGULA ALNUS BARK EXTRACT|FRANGULA ALNUS BARK EXTRACT
C3475109|T109|1310064|RXNORM|CITRUS SINENSIS FRUIT OIL|CITRUS SINENSIS FRUIT OIL
C3484475|T121|1310065|RXNORM|RHEUM OFFICINALE ROOT EXTRACT|RHEUM OFFICINALE ROOT EXTRACT
C3475151|T121|1310066|RXNORM|MATRICARIA RECUTITA LEAF EXTRACT|MATRICARIA CHAMOMILLA LEAF EXTRACT
C3255611|T121|1310067|RXNORM|PUNICA GRANATUM SEED EXTRACT|PUNICA GRANATUM SEED EXTRACT
C3255616|T121|1310068|RXNORM|TRICHOSANTHES CUCUMERINA SEED EXTRACT|TRICHOSANTHES CUCUMERINA SEED EXTRACT
C3475323|T121|1310069|RXNORM|HYPOXIS HEMEROCALLIDEA ROOT EXTRACT|HYPOXIS HEMEROCALLIDEA ROOT EXTRACT
C3693002|T121|1442998|RXNORM|CETYL DIMETHICONE 150|CETYL DIMETHICONE 150
C0304632|T121|91327|RXNORM|OCTISALATE|OCTISALATE
C0304629|T109|91324|RXNORM|MERADIMATE|MERADIMATE
C0056478|T109|1362910|RXNORM|CREOSOL|CREOSOL
C2080601|T121|820369|RXNORM|GUAIFENESIN / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE|GUAIFENESIN / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE
C2741584|T129|901505|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP A OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|NEISSERIA MENINGITIDIS SEROGROUP A OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C0304137|T109|1309388|RXNORM|OIL OF GINGER|GINGER ROOT OIL
C3528818|T121|1363429|RXNORM|ALPHA-ARBUTIN|ALPHA-ARBUTIN
C2731464|T121|895365|RXNORM|SYDNEY GOLDEN WATTLE POLLEN EXTRACT|ACACIA LONGIFOLIA POLLEN EXTRACT
C2183062|T121|823322|RXNORM|CHLORPHENIRAMINE / DEXAMETHASONE|CHLORPHENIRAMINE / DEXAMETHASONE
C1696465|T122|8375|RXNORM|PLACEBO|PLACEBO
C3153172|T121|1098639|RXNORM|HYPROMELLOSE / TETRAHYDROZOLINE / ZINC SULFATE|HYPROMELLOSE / TETRAHYDROZOLINE / ZINC SULFATE
C0032032|T195|8372|RXNORM|PIVAMPICILLIN|PIVAMPICILLIN
C0032036|T121|8373|RXNORM|PIZOTYLINE|PIZOTYLINE
C0982134|T121|314605|RXNORM|EGG YOLK PHOSPHOLIPIDS|EGG YOLK PHOSPHOLIPIDS
C3555490|T121|1376215|RXNORM|SAMBUCUS CANADENSIS FLOWER EXTRACT|SAMBUCUS CANADENSIS FLOWER EXTRACT
C3555491|T121|1376214|RXNORM|CORYDALIS AMBIGUA TUBER EXTRACT|CORYDALIS AMBIGUA TUBER EXTRACT
C3255661|T121|1310288|RXNORM|CHAENOMELES SPECIOSA FRUIT|CHAENOMELES SPECIOSA FRUIT
C3486220|T121|1310289|RXNORM|BOS TAURUS PARATHYROID GLAND PREPARATION|BOVINE PARATHYROID GLAND PREPARATION
C3555494|T121|1376211|RXNORM|COPTIS CHINENSIS ROOT EXTRACT|COPTIS CHINENSIS ROOT EXTRACT
C3692541|T121|1442192|RXNORM|ARISTOLOCHIA SERPENTARIA ROOT EXTRACT|ARISTOLOCHIA SERPENTARIA ROOT EXTRACT
C3488554|T121|1310285|RXNORM|GAULTHERIA PROCUMBENS TOP EXTRACT|GAULTHERIA PROCUMBENS TOP EXTRACT
C0969589|T121|304962|RXNORM|ARFORMOTEROL|ARFORMOTEROL
C3254761|T109|1310287|RXNORM|LUFFA ACUTANGULA FRUIT EXTRACT|LUFFA EXTRACT
C3488416|T121|1310280|RXNORM|ACORUS CALAMUS EXTRACT|ACORUS CALAMUS EXTRACT
C3488419|T121|1310281|RXNORM|SCOMBEROMORUS CAVALLA EXTRACT|SCOMBEROMORUS CAVALLA EXTRACT
C3488449|T121|1310282|RXNORM|TRILLIUM ERECTUM EXTRACT|TRILLIUM ERECTUM EXTRACT
C1739768|T121|1114195|RXNORM|RIVAROXABAN|RIVAROXABAN
C0305040|T197|91588|RXNORM|THALLOUS CHLORIDE TL201|THALLOUS CHLORIDE TL201
C3257523|T109|1305719|RXNORM|CUCUMBER EXTRACT|CUCUMBER EXTRACT
C3819179|T121|1492051|RXNORM|DEXTROMETHORPHAN / PHENYLEPHRINE / TRIPROLIDINE|DEXTROMETHORPHAN / PHENYLEPHRINE / TRIPROLIDINE
C0939230|T121|636632|RXNORM|ESTRADIOL / MEDROXYPROGESTERONE|ESTRADIOL / MEDROXYPROGESTERONE
C2928655|T121|1007740|RXNORM|LACTOBACILLUS ACIDOPHILUS / PECTIN|LACTOBACILLUS ACIDOPHILUS / PECTIN
C2928656|T121|1007741|RXNORM|HALOMETASONE / TRICLOSAN|HALOMETASONE / TRICLOSAN
C2928657|T121|1007742|RXNORM|BROMHEXINE / BUTETAMATE|BROMHEXINE / BUTETAMATE
C2928658|T121|1007743|RXNORM|ACETONE / ETHANOL|ACETONE / ETHANOL
C2928659|T121|1007744|RXNORM|CARBOCYSTEINE / SOBREROL|CARBOCYSTEINE / SOBREROL
C2928660|T121|1007745|RXNORM|BROMHEXINE / GUAIFENESIN|BROMHEXINE / GUAIFENESIN
C2928661|T121|1007746|RXNORM|AMMONIUM CHLORIDE / ISOAMINILE|AMMONIUM CHLORIDE / ISOAMINILE
C2928662|T121|1007747|RXNORM|DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / SODIUM ACETATE / SODIUM CHLORIDE|DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / SODIUM ACETATE / SODIUM CHLORIDE
C2928663|T121|1007748|RXNORM|MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE / SODIUM PHOSPHATE, DIBASIC|MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE / SODIUM PHOSPHATE, DIBASIC
C2928664|T121|1007749|RXNORM|DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE|DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE
C2980841|T129|1426665|RXNORM|TRICHOSPORON CUTANEUM ALLERGENIC EXTRACT|TRICHOSPORON CUTANEUM ALLERGENIC EXTRACT
C2928881|T121|1007968|RXNORM|DEMELVERIN / TRIHEXYPHENIDYL|DEMELVERIN / TRIHEXYPHENIDYL
C2928882|T121|1007969|RXNORM|CALCIUM PHOSPHATE / SODIUM FLUORIDE|CALCIUM PHOSPHATE / SODIUM FLUORIDE
C3475221|T121|1312539|RXNORM|ALOE VERA WHOLE EXTRACT|ALOE VERA WHOLE EXTRACT
C1329993|T121|404788|RXNORM|CHLORPHENIRAMINE / DIHYDROCODEINE / PHENYLEPHRINE|CHLORPHENIRAMINE / DIHYDROCODEINE / PHENYLEPHRINE
C0072315|T121|34769|RXNORM|PROGLUMETACIN|PROGLUMETACIN
C1874725|T121|691347|RXNORM|CARBOXYMETHYLCELLULOSE / DOCUSATE|CARBOXYMETHYLCELLULOSE / DOCUSATE
C1874724|T121|691346|RXNORM|CARBOXYMETHYLCELLULOSE / CASANTHRANOL / DOCUSATE|CARBOXYMETHYLCELLULOSE / CASANTHRANOL / DOCUSATE
C1874726|T121|691348|RXNORM|CARBOXYMETHYLCELLULOSE / DOCUSATE / PHENOLPHTHALEIN|CARBOXYMETHYLCELLULOSE / DOCUSATE / PHENOLPHTHALEIN
C2938411|T129|1012190|RXNORM|NAVY KIDNEY BEAN ALLERGENIC EXTRACT|NAVY KIDNEY BEAN ALLERGENIC EXTRACT
C1178459|T121|360262|RXNORM|APPLE CIDER VINEGAR|APPLE CIDER VINEGAR
C0026651|T195|7069|RXNORM|MOXALACTAM|MOXALACTAM
C0939921|T121|285265|RXNORM|BITTER APPLE PREPARATION|BITTER APPLE PREPARATION
C3486004|T109|1426662|RXNORM|TRIISOSTEARIN|TRIISOSTEARIN
C0031635|T121|8226|RXNORM|PHOSPHOCYSTEAMINE|PHOSPHOCYSTEAMINE
C2109244|T121|814091|RXNORM|JUNIPER TAR / ZINC PYRITHIONE|JUNIPER TAR / ZINC PYRITHIONE
C0054323|T121|19943|RXNORM|BUZEPIDE METIODIDE|BUZEPIDE METIODIDE
C0077046|T109|1439115|RXNORM|TRICHLOROSUCROSE|SUCRALOSE
C3489114|T121|1311229|RXNORM|SUS SCROFA ILEUM PREPARATION|PORCINE ILEUM PREPARATION
C0315276|T007|1311228|RXNORM|MORGANELLA MORGANII|MORGANELLA MORGANII
C0021757|T129|1311225|RXNORM|INTERLEUKIN-3|INTERLEUKIN-3
C0021236|T121|1311224|RXNORM|INDOLE|INDOLE
C2937963|T129|1010971|RXNORM|PEPPERMINT ALLERGENIC EXTRACT|PEPPERMINT ALLERGENIC EXTRACT
C3489113|T121|1311226|RXNORM|SUS SCROFA BILE DUCT PREPARATION|PORCINE BILE DUCT PREPARATION
C0102819|T121|1314612|RXNORM|ALTRENOGEST|ALTRENOGEST
C3488294|T121|1311223|RXNORM|SUS SCROFA THALAMUS LATERAL GENICULATE NUCLEUS PREPARATION|PORCINE THALAMUS LATERAL GENICULATE NUCLEUS PREPARATION
C3700904|T109|1485786|RXNORM|MUCUNA PRURIENS SEED EXTRACT|MUCUNA PRURIENS SEED EXTRACT
C0026056|T121|6960|RXNORM|MIDAZOLAM|MIDAZOLAM
C0026078|T121|6963|RXNORM|MIDODRINE|MIDODRINE
C3700905|T109|1485785|RXNORM|APPLE FRUIT OIL|APPLE FRUIT OIL
C0032911|T121|8628|RXNORM|PRAZIQUANTEL|PRAZIQUANTEL
C0032912|T121|8629|RXNORM|PRAZOSIN|PRAZOSIN
C3463996|T109|1426663|RXNORM|LIQUID PETROLEUM|LIQUID PETROLEUM
C0031453|T123|8156|RXNORM|PHENYLALANINE|PHENYLALANINE
C0032910|T121|8627|RXNORM|PRAZEPAM|PRAZEPAM
C0031447|T121|8152|RXNORM|PHENTERMINE|PHENTERMINE
C0031448|T121|8153|RXNORM|PHENTOLAMINE|PHENTOLAMINE
C0031444|T121|8150|RXNORM|PHENPROCOUMON|PHENPROCOUMON
C0023861|T007|1491871|RXNORM|LISTERIA MONOCYTOGENES|LISTERIA MONOCYTOGENES
C0023238|T007|1491870|RXNORM|LEGIONELLA PNEUMOPHILA|LEGIONELLA PNEUMOPHILA
C0036960|T007|1491872|RXNORM|SHIGELLA SONNEI|SHIGELLA SONNEI
C0081876|T121|40790|RXNORM|PANTOPRAZOLE|PANTOPRAZOLE
C3474472|T121|1423273|RXNORM|PPG-26-BUTETH-26|PPG-26-BUTETH-26
C0982395|T197|314837|RXNORM|SODIUM PHOSPHATE DIHYDRATE|SODIUM PHOSPHATE DIHYDRATE
C2057753|T121|812199|RXNORM|NOSCAPINE / THEOPHYLLINE|NOSCAPINE / THEOPHYLLINE
C3256595|T121|1307572|RXNORM|ALBIZIA JULIBRISSIN BARK EXTRACT|ALBIZIA JULIBRISSIN BARK EXTRACT
C2740652|T129|899466|RXNORM|ONION ALLERGENIC EXTRACT|ONION ALLERGENIC EXTRACT
C3667115|T121|1438641|RXNORM|COLLOIDAL OATMEAL / MENTHOL|COLLOIDAL OATMEAL / MENTHOL
C1875699|T121|690166|RXNORM|PROMETHAZINE / PSEUDOEPHEDRINE|PROMETHAZINE / PSEUDOEPHEDRINE
C3540829|T121|1435397|RXNORM|PUERARIA MONTANA VAR. LOBATA WHOLE EXTRACT|PUERARIA MONTANA VAR. LOBATA WHOLE EXTRACT
C0318366|T005|1435394|RXNORM|HUMAN COXSACKIEVIRUS A2|HUMAN COXSACKIEVIRUS A2
C0318371|T005|1435395|RXNORM|HUMAN COXSACKIEVIRUS A7|HUMAN COXSACKIEVIRUS A7
C2607479|T123|1534763|RXNORM|ALBIGLUTIDE|ALBIGLUTIDE
C3665154|T121|1435393|RXNORM|FRASERA CAROLINIENSIS ROOT EXTRACT|FRASERA CAROLINIENSIS ROOT EXTRACT
C3665152|T121|1435390|RXNORM|ETHYL JOJOBATE|ETHYL JOJOBATE
C1875694|T121|690161|RXNORM|PREDNISOLONE / SULFACETAMIDE|PREDNISOLONE / SULFACETAMIDE
C0527076|T197|1311081|RXNORM|CADMIUM IODIDE|CADMIUM IODIDE
C1950072|T121|1311080|RXNORM|WOOD ANT PREPARATION|FORMICA RUFA PREPARATION
C3486674|T121|1311083|RXNORM|RANCID BEEF PREPARATION|RANCID BEEF PREPARATION
C0043314|T123|1311085|RXNORM|XANTHINE|XANTHINE
C3486618|T121|1311084|RXNORM|CHOLINE HYDROXIDE|CHOLINE HYDROXIDE
C0039994|T196|1534769|RXNORM|THORIUM|THORIUM
C0035973|T196|1534768|RXNORM|RUTHENIUM|RUTHENIUM
C3473404|T121|1312579|RXNORM|FILIPENDULA ULMARIA WHOLE EXTRACT|FILIPENDULA ULMARIA WHOLE EXTRACT
C3256739|T121|1426661|RXNORM|USNEA BARBATA EXTRACT|USNEA BARBATA EXTRACT
C3663611|T122|1433497|RXNORM|SOYETHYL MORPHOLINIUM ETHOSULFATE|SOYETHYL MORPHOLINIUM ETHOSULFATE
C3663610|T122|1433496|RXNORM|POLY(METHYL METHACRYLATE; 450000 MW)|POLY(METHYL METHACRYLATE; 450000 MW)
C3663609|T122|1433495|RXNORM|ETHYL ACRYLATE-METHACRYLIC ACID-STEARETH-20 METHACRYLATE COPOLYMER|ETHYL ACRYLATE-METHACRYLIC ACID-STEARETH-20 METHACRYLATE COPOLYMER
C0032611|T122|1358182|RXNORM|POLYTETRAFLUOROETHYLENE|POLYTETRAFLUOROETHYLENE
C0717858|T121|214652|RXNORM|IBUPROFEN / PSEUDOEPHEDRINE|IBUPROFEN / PSEUDOEPHEDRINE
C3255754|T122|1312573|RXNORM|ETHYL ACRYLATE AND METHYL METHACRYLATE COPOLYMER (2:1; 600000 MW)|ETHYL ACRYLATE AND METHYL METHACRYLATE COPOLYMER (2:1; 600000 MW)
C3255759|T109|1312574|RXNORM|ETHYL VALERATE|ETHYL VALERATE
C2827148|T121|1312575|RXNORM|ETHYLCELLULOSE (7 MPA.S)|ETHYLCELLULOSE (7 MPA.S)
C3255765|T121|1312576|RXNORM|ETHYLENE-VINYL ACETATE COPOLYMER (19% VINYLACETATE)|ETHYLENE-VINYL ACETATE COPOLYMER (19% VINYLACETATE)
C3255767|T109|1312577|RXNORM|ETHYLENE-VINYL ACETATE COPOLYMER (40% VINYL ACETATE)|ETHYLENE-VINYL ACETATE COPOLYMER (40% VINYL ACETATE)
C1620942|T121|580117|RXNORM|AFRICAN PYGEUM EXTRACT|AFRICAN PYGEUM EXTRACT
C0724570|T197|221090|RXNORM|DIBASIC SODIUM PHOSPHATE HEPTAHYDRATE|DIBASIC SODIUM PHOSPHATE HEPTAHYDRATE
C0724573|T121|221091|RXNORM|DIPTHERIA PROTEIN|DIPTHERIA PROTEIN
C0008260|T123|2388|RXNORM|CHLOROPHYLL|CHLOROPHYLL
C1166032|T121|350344|RXNORM|CONIUM PREPARATION|CONIUM PREPARATION
C2349150|T121|1319902|RXNORM|WHITE OAK BARK EXTRACT|QUERCUS ALBA BARK EXTRACT
C1618310|T121|580119|RXNORM|STINGING NETTLE EXTRACT|STINGING NETTLE EXTRACT
C2929138|T121|1008231|RXNORM|ANTIPYRINE / BENZOCAINE / ZINC ACETATE|ANTIPYRINE / BENZOCAINE / ZINC ACETATE
C2929137|T121|1008230|RXNORM|ALANINE / ARGININE / ASPARTATE / CYSTEINE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / TAURINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / ASPARTATE / CYSTEINE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / TAURINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929140|T121|1008233|RXNORM|GUARANA PREPARATION / LEVOCARNITINE|GUARANA PREPARATION / LEVOCARNITINE
C2929139|T121|1008232|RXNORM|SALICYLAMIDE / VITAMIN B 12|SALICYLAMIDE / VITAMIN B 12
C2929142|T121|1008235|RXNORM|ASCORBIC ACID / D-BIOTIN / FOLIC ACID / NIACINAMIDE / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|ASCORBIC ACID / D-BIOTIN / FOLIC ACID / NIACINAMIDE / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C2929141|T121|1008234|RXNORM|PHOLCODINE / PSEUDOEPHEDRINE|PHOLCODINE / PSEUDOEPHEDRINE
C2929144|T121|1008237|RXNORM|CALCIUM CARBONATE / DEHYDROEPIANDROSTERONE|CALCIUM CARBONATE / PRASTERONE
C2929143|T121|1008236|RXNORM|CHLORAMPHENICOL / PREDNISOLONE|CHLORAMPHENICOL / PREDNISOLONE
C2929145|T121|1008238|RXNORM|COLCHICINE / PODOPHYLLIN|COLCHICINE / PODOPHYLLIN
C3700990|T121|1486780|RXNORM|FORMALDEHYDE / METHANOL|FORMALDEHYDE / METHANOL
C0245561|T121|72625|RXNORM|DULOXETINE|DULOXETINE
C0005038|T131|1388|RXNORM|LINDANE|LINDANE
C3536832|T197|411|RXNORM|AIR|MEDICAL AIR
C1095908|T121|319829|RXNORM|LEGUME PREPARATION|LEGUME PREPARATION
C3667875|T121|1440241|RXNORM|SAFFLOWER SEED EXTRACT|SAFFLOWER SEED EXTRACT
C0005035|T121|1385|RXNORM|BENZBROMARONE|BENZBROMARONE
C1095903|T121|319824|RXNORM|GENTIAN PREPARATION|GENTIAN PREPARATION
C1095902|T121|319823|RXNORM|THYME PREPARATION|THYME PREPARATION
C2111789|T121|815276|RXNORM|POLYETHYLENE GLYCOL 3350 / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE / SODIUM SULFATE|POLYETHYLENE GLYCOL 3350 / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE / SODIUM SULFATE
C2701629|T129|852532|RXNORM|ROUGH MARSHELDER POLLEN EXTRACT|IVA ANNUA POLLEN EXTRACT
C2709738|T129|854934|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 11A VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 11A VACCINE
C0149389|T121|58301|RXNORM|ZINC PICOLINATE|ZINC PICOLINATE
C2701633|T129|852539|RXNORM|POVERTY WEED POLLEN EXTRACT|IVA AXILLARIS POLLEN EXTRACT
C1648605|T121|606096|RXNORM|ACETAMINOPHEN / GUAIFENESIN|ACETAMINOPHEN / GUAIFENESIN
C2929261|T121|1008356|RXNORM|CHLOROXYLENOL / LIDOCAINE|CHLOROXYLENOL / LIDOCAINE
C2069095|T121|1008357|RXNORM|FOLIC ACID / POLYSACCHARIDE IRON COMPLEX|FOLIC ACID / POLYSACCHARIDE IRON COMPLEX
C2929259|T121|1008354|RXNORM|COAL TAR / MERCURY, AMMONIATED / METHENAMINE|COAL TAR / MERCURY, AMMONIATED / METHENAMINE
C2929260|T121|1008355|RXNORM|FORMALDEHYDE / SALICYLIC ACID|FORMALDEHYDE / SALICYLIC ACID
C2929257|T121|1008352|RXNORM|TESTOSTERONE 17-PHENYLPROPIONATE / TESTOSTERONE ISOCAPROATE / TESTOSTERONE PROPIONATE|TESTOSTERONE 17-PHENYLPROPIONATE / TESTOSTERONE ISOCAPROATE / TESTOSTERONE PROPIONATE
C3700986|T109|1486522|RXNORM|2-SULFOPALMITATE|2-SULFOPALMITATE
C2929255|T121|1008350|RXNORM|MELATONIN / PYRIDOXINE|MELATONIN / PYRIDOXINE
C0066275|T109|1486520|RXNORM|METHYL PALMITATE|METHYL PALMITATE
C2194326|T121|818306|RXNORM|ACETAMINOPHEN / MEPHENESIN|ACETAMINOPHEN / MEPHENESIN
C1166079|T121|350386|RXNORM|MANDRAGORA OFFICINARUM PREPARATION|MANDRAGORA OFFICINARUM PREPARATION
C2929263|T121|1008358|RXNORM|CHROMOUS CHLORIDE / COPPER SULFATE / MANGANESE CHLORIDE / ZINC CHLORIDE|CHROMOUS CHLORIDE / COPPER SULFATE / MANGANESE CHLORIDE / ZINC CHLORIDE
C2929264|T121|1008359|RXNORM|ESTRADIOL / ETHINYL ESTRADIOL / LEVONORGESTREL|ESTRADIOL / ETHINYL ESTRADIOL / LEVONORGESTREL
C1445179|T129|894961|RXNORM|CANARY FEATHER EXTRACT|SERINUS CANARIA FEATHER EXTRACT
C0043339|T196|11363|RXNORM|XENON|XENON
C0205758|T121|66887|RXNORM|RACEPINEPHRINE|RACEPINEPHRINE
C0600416|T121|155097|RXNORM|HAWTHORN PREPARATION|HAWTHORN PREPARATION
C2827266|T121|1307079|RXNORM|METHYL BENZOIN|METHYL BENZOIN
C3256110|T121|1305743|RXNORM|ILEX PARAGUARIENSIS LEAF EXTRACT|ILEX PARAGUARIENSIS LEAF EXTRACT
C2940158|T129|1014690|RXNORM|JACK PINE POLLEN EXTRACT|PINUS BANKSIANA POLLEN EXTRACT
C2709746|T129|854942|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 17F VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 17F VACCINE
C1706292|T109|1309228|RXNORM|HYPERICUM EXTRACT|HYPERICUM EXTRACT
C0935916|T121|282357|RXNORM|FULVESTRANT|FULVESTRANT
C0038689|T195|10180|RXNORM|SULFAMETHOXAZOLE|SULFAMETHOXAZOLE
C0014644|T005|1316054|RXNORM|EPSTEIN-BARR VIRUS|EPSTEIN-BARR VIRUS
C0014323|T204|1316053|RXNORM|ENTAMOEBA HISTOLYTICA|ENTAMOEBA HISTOLYTICA
C2193953|T121|815852|RXNORM|CODEINE / EPHEDRINE|CODEINE / EPHEDRINE
C3643345|T121|1424359|RXNORM|PERSICARIA TINCTORIA TOP EXTRACT|PERSICARIA TINCTORIA TOP EXTRACT
C0282328|T123|82089|RXNORM|ISPAGHULA EXTRACT|ISPAGHULA EXTRACT
C0282327|T121|82088|RXNORM|PLANTAGO SEED|PLANTAGO SEED
C0253029|T121|1305749|RXNORM|GLYCERYL BEHENATE|GLYCERYL BEHENATE
C3255853|T109|1424357|RXNORM|PADINA PAVONICA EXTRACT|PADINA PAVONICA EXTRACT
C2080474|T121|813172|RXNORM|LIDOCAINE / PHENYLBUTAZONE|LIDOCAINE / PHENYLBUTAZONE
C3255634|T109|1305748|RXNORM|GLYCERETH-2 COCOATE|GLYCERETH-2 COCOATE
C3645000|T121|1426267|RXNORM|ACRIFLAVINE / GENTIAN VIOLET / SODIUM PROPIONATE|ACRIFLAVINE / GENTIAN VIOLET / SODIUM PROPIONATE
C3834062|T121|1542900|RXNORM|CAULOSIDE D|CAULOSIDE D
C3834061|T121|1542901|RXNORM|PROPYLENE GLYCOL 1-(2-METHYLBUTYRATE)|PROPYLENE GLYCOL 1-(2-METHYLBUTYRATE)
C2955629|T121|1050797|RXNORM|ALISKIREN / AMLODIPINE / HYDROCHLOROTHIAZIDE|ALISKIREN / AMLODIPINE / HYDROCHLOROTHIAZIDE
C3853907|T121|1595298|RXNORM|COCAMIDOPROPYL PROPYLENE GLYCOL-DIMONIUM CHLORIDE|COCAMIDOPROPYL PROPYLENE GLYCOL-DIMONIUM CHLORIDE
C0060520|T130|25138|RXNORM|FLUORESCEIN|FLUORESCEIN
C0109265|T109|1309221|RXNORM|CHAMOMILE FLOWER OIL|CHAMOMILE FLOWER OIL
C3854119|T121|1549107|RXNORM|LYSIMACHIA NUMMULARIA EXTRACT|LYSIMACHIA NUMMULARIA EXTRACT
C1435444|T121|460132|RXNORM|DARUNAVIR|DARUNAVIR
C0064723|T197|1549104|RXNORM|LEAD SULFIDE|LEAD SULFIDE
C3855804|T121|1549103|RXNORM|HYACINTHUS ORIENTALIS WHOLE EXTRACT|HYACINTHUS ORIENTALIS WHOLE EXTRACT
C3855803|T121|1549102|RXNORM|BOS TAURUS ARTERY PREPARATION|BOS TAURUS ARTERY PREPARATION
C2741520|T129|901346|RXNORM|TAPIOCA STARCH ALLERGENIC EXTRACT|TAPIOCA STARCH ALLERGENIC EXTRACT
C0074127|T130|36224|RXNORM|SCARLET RED|SCARLET RED
C1259855|T197|1549109|RXNORM|PLATINIC CHLORIDE|PLATINIC CHLORIDE
C3855807|T121|1549108|RXNORM|PICEA ABIES LEAF EXTRACT|PICEA ABIES LEAF EXTRACT
C3651790|T121|1428044|RXNORM|EGG SHELL MEMBRANE|EGG SHELL MEMBRANE
C0872895|T121|259265|RXNORM|GINKGO BILOBA LEAF EXTRACT|GINKGO BILOBA LEAF EXTRACT
C0872893|T121|259263|RXNORM|ESTROGENIC SUBSTANCES|ESTROGENIC SUBSTANCES
C0872887|T121|259260|RXNORM|BUTTON MUSHROOM EXTRACT|BUTTON MUSHROOM EXTRACT
C0872889|T121|259261|RXNORM|CHASTE BERRY EXTRACT|CHASTE BERRY EXTRACT
C2347037|T121|1319885|RXNORM|BLACK WALNUT LEAVES EXTRACT|JUGLANS NIGRA LEAF EXTRACT
C0021225|T130|259268|RXNORM|PENTETATE INDIUM DISODIUM,IN-111|INDIUM IN-111 PENTETATE DISODIUM
C0082646|T130|41144|RXNORM|GADODIAMIDE|GADODIAMIDE
C0025051|T121|6680|RXNORM|MEDAZEPAM|MEDAZEPAM
C3860003|T109|1594416|RXNORM|BUTYL ETHER|BUTYL ETHER
C2929722|T121|1008824|RXNORM|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / VITAMIN B 12|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / VITAMIN B 12
C2929723|T121|1008825|RXNORM|CINNARIZINE / HEPTAMINOL|CINNARIZINE / HEPTAMINOL
C2929724|T121|1008826|RXNORM|AMOXICILLIN / CARBOCYSTEINE|AMOXICILLIN / CARBOCYSTEINE
C2929725|T121|1008827|RXNORM|CETRIMIDE / LIDOCAINE / MENTHOL|CETRIMIDE / LIDOCAINE / MENTHOL
C2193831|T121|1008820|RXNORM|AMPICILLIN / DICLOXACILLIN|AMPICILLIN / DICLOXACILLIN
C2929719|T121|1008821|RXNORM|CASTOR OIL / PERUVIAN BALSAM|CASTOR OIL / PERUVIAN BALSAM
C2929720|T121|1008822|RXNORM|SWEETLEAF PREPARATION / ZINC CHLORIDE|SWEETLEAF PREPARATION / ZINC CHLORIDE
C2929721|T121|1008823|RXNORM|GINKGO BILOBA EXTRACT / HEPTAMINOL / TROXERUTIN|GINKGO BILOBA EXTRACT / HEPTAMINOL / TROXERUTIN
C0008328|T125|2420|RXNORM|CHOLECYSTOKININ|CHOLECYSTOKININ, HUMAN
C2929726|T121|1008828|RXNORM|CAFFEINE / PROPYPHENAZONE|CAFFEINE / PROPYPHENAZONE
C2929727|T121|1008829|RXNORM|HYDROCORTISONE / ICTASOL|HYDROCORTISONE / ICTASOL
C0008359|T129|2427|RXNORM|CHOLERA VACCINE|CHOLERA VACCINE
C3833028|T121|1540229|RXNORM|KETOROLAC / PHENYLEPHRINE|KETOROLAC / PHENYLEPHRINE
C0982027|T121|314506|RXNORM|APIOLE|APIOLE
C3848575|T196|1546269|RXNORM|URANIUM CATION (6+)|URANIUM CATION (6+)
C2939575|T121|1013615|RXNORM|CHLORCYCLIZINE / CODEINE / PHENYLEPHRINE|CHLORCYCLIZINE / CODEINE / PHENYLEPHRINE
C0059836|T121|236122|RXNORM|ETHYLNICOTINATE|ETHYLNICOTINATE
C0771364|T121|236121|RXNORM|ECHINACEA ANGUSTIFOLIA EXTRACT|ECHINACEA ANGUSTIFOLIA EXTRACT
C3255717|T109|1426421|RXNORM|PIMPINELLA ANISUM EXTRACT|PIMPINELLA ANISUM EXTRACT
C0009053|T126|898492|RXNORM|COLLAGENASE CLOSTRIDIUM HISTOLYTICUM|COLLAGENASE CLOSTRIDIUM HISTOLYTICUM
C0058895|T121|23796|RXNORM|EBASTINE|EBASTINE
C3474374|T121|1300887|RXNORM|CAMPHOR / PHENOL / TANNIC ACID / ZINC OXIDE|CAMPHOR / PHENOL / TANNIC ACID / ZINC OXIDE
C2702423|T129|1294634|RXNORM|RED PAPER WASP VENOM PROTEIN|POLISTES ANNULARIS VENOM
C0035525|T121|9344|RXNORM|RIBAVIRIN|RIBAVIRIN
C0038670|T121|10169|RXNORM|SULFACETAMIDE|SULFACETAMIDE
C0038670|T121|10169|RXNORM|SULFACETAMIDE|SULFACETAMIDE
C0038666|T195|10168|RXNORM|SULBENICILLIN|SULBENICILLIN
C0038665|T195|10167|RXNORM|SULBACTAM|SULBACTAM
C0218986|T129|70223|RXNORM|ALDESLEUKIN|ALDESLEUKIN
C3531215|T109|1366331|RXNORM|TAGETES MINUTA FLOWER OIL|TAGETES MINUTA FLOWER OIL
C3531214|T109|1366330|RXNORM|PINUS PALUSTRIS LEAF EXTRACT|PINUS PALUSTRIS LEAF EXTRACT
C0146224|T121|57308|RXNORM|TOPOTECAN|TOPOTECAN
C0055906|T121|21255|RXNORM|CLOFEXAMIDE|CLOFEXAMIDE
C0055904|T121|21254|RXNORM|CHLOPHEDIANOL|CHLOPHEDIANOL
C1365461|T109|436163|RXNORM|TEA TREE EXTRACT|TEA TREE EXTRACT
C0300990|T197|1552051|RXNORM|COPPER ARSENATE|COPPER ARSENATE
C3859186|T109|1592296|RXNORM|KALE EXTRACT|KALE EXTRACT
C0006400|T121|1815|RXNORM|BUPIVACAINE|BUPIVACAINE
C0006403|T121|1817|RXNORM|BUPRANOLOL|BUPRANOLOL
C1445713|T121|466479|RXNORM|NEOMYCIN / POLYMYXIN B / PRAMOXINE|NEOMYCIN / POLYMYXIN B / PRAMOXINE
C1445712|T121|466478|RXNORM|LIDOCAINE / NEOMYCIN / POLYMYXIN B|LIDOCAINE / NEOMYCIN / POLYMYXIN B
C0939876|T121|285223|RXNORM|CAT'S CLAW PREPARATION|CAT'S CLAW PREPARATION
C0939875|T121|285222|RXNORM|CALENDULA OFFICINALIS EXTRACT|CALENDULA OFFICINALIS EXTRACT
C0939872|T121|285220|RXNORM|CHELIDONIUM MAJUS PREPARATION|CHELIDONIUM MAJUS EXTRACT
C0006405|T121|1819|RXNORM|BUPRENORPHINE|BUPRENORPHINE
C2825635|T195|1437806|RXNORM|TULATHROMYCIN A|TULATHROMYCIN A
C1445704|T121|466470|RXNORM|IODINE / METHYL SALICYLATE|IODINE / METHYL SALICYLATE
C0525133|T197|134568|RXNORM|BENTOQUATAM|BENTOQUATAM
C3651714|T168|1431150|RXNORM|NIGELLA SATIVA SEED OIL|CARAWAY BLACK OIL
C3651948|T197|1431152|RXNORM|FLUOROSILICATE|FLUOROSILICATE
C3651712|T121|1431153|RXNORM|MYRISTAMINE OXIDE|MYRISTAMINE OXIDE
C0079856|T121|40169|RXNORM|MORICIZINE|MORICIZINE
C2347036|T129|891695|RXNORM|BLACK WALNUT ALLERGENIC EXTRACT|WALLIA NIGRA ALLERGENIC EXTRACT
C3255676|T109|1314281|RXNORM|HEXAMETHYLINDANOPYRAN|HEXAMETHYLINDANOPYRAN
C3255802|T121|1314282|RXNORM|POLYACRYLIC ACID (450000 MW)|POLYACRYLIC ACID (450000 MW)
C3255813|T196|1314283|RXNORM|STANNOUS CATION|STANNOUS CATION
C3255857|T121|1314284|RXNORM|PALMITOYL TRIPEPTIDE-5|PALMITOYL TRIPEPTIDE-5
C3255873|T109|1314285|RXNORM|STEARIC DIETHANOLAMIDE|STEARIC DIETHANOLAMIDE
C3255878|T121|1314286|RXNORM|STEARYL MYRISTATE|STEARYL MYRISTATE
C3255937|T109|1314287|RXNORM|HYDROGENATED POLYBUTENE (1300 MW)|HYDROGENATED POLYBUTENE (1300 MW)
C3255964|T121|1314288|RXNORM|PEG-10 SOY STEROL|PEG-10 SOY STEROL
C3256087|T109|1314289|RXNORM|QUATERNIUM-15 CIS-FORM|QUATERNIUM-15 CIS-FORM
C3855256|T109|1547621|RXNORM|PSEUDOLARIX AMABILIS BARK EXTRACT|PSEUDOLARIX AMABILIS BARK EXTRACT
C3855257|T109|1547622|RXNORM|PEG-32 HYDROGENATED PALM GLYCERIDES|PEG-32 HYDROGENATED PALM GLYCERIDES
C3855258|T109|1547623|RXNORM|CHRYSANTHEMIN EXTRACT|CHRYSANTHEMIN EXTRACT
C2079440|T121|1355936|RXNORM|CYCLOPENTAMINE / ISOPROTERENOL|CYCLOPENTAMINE / ISOPROTERENOL
C3530627|T121|1364986|RXNORM|ACONITUM KUSNEZOFFI ROOT EXTRACT|ACONITUM KUSNEZOFFI ROOT EXTRACT
C0055458|T197|1543755|RXNORM|CHLOROUS ACID|CHLOROUS ACID
C0011588|T121|3226|RXNORM|DEQUALINIUM|DEQUALINIUM
C3665327|T109|1435890|RXNORM|BUCKMINSTERFULLERENE|BUCKMINSTERFULLERENE
C0303403|T196|90540|RXNORM|INDIUM-111|INDIUM-111
C0164814|T121|59838|RXNORM|HALAZONE|HALAZONE
C0164815|T121|59839|RXNORM|PENCICLOVIR|PENCICLOVIR
C1509794|T121|477189|RXNORM|SAW PALMETTO FRUIT EXTRACT|SAW PALMETTO FRUIT EXTRACT
C3505683|T121|1359090|RXNORM|POLYQUATERNIUM-51 (2-METHACRYLOYLOXYETHYL PHOSPHORYLCHOLINE:N-BUTYL METHACRYLATE; 3:7)|POLYQUATERNIUM-51 (2-METHACRYLOYLOXYETHYL PHOSPHORYLCHOLINE:N-BUTYL METHACRYLATE; 3:7)
C0993551|T130|317675|RXNORM|SAMARIUM SM 153 LEXIDRONAM PENTASODIUM|SAMARIUM SM 153 LEXIDRONAM PENTASODIUM
C0259507|T121|78484|RXNORM|DANAPAROID|DANAPAROID
C3505684|T127|1359091|RXNORM|TOCOPHERYL NICOTINATE, D-.ALPHA.|TOCOPHERYL NICOTINATE, D-.ALPHA.
C1874533|T121|690286|RXNORM|BENZOXIQUINE / ICHTHAMMOL|BENZOXIQUINE / ICHTHAMMOL
C0012010|T121|3322|RXNORM|DIAZEPAM|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM|DIAZEPAM
C0149381|T121|58300|RXNORM|ZINC GLUCONATE|ZINC GLUCONATE
C0020223|T121|5470|RXNORM|HYDRALAZINE|HYDRALAZINE
C0012022|T121|3327|RXNORM|DIAZOXIDE|DIAZOXIDE
C0012022|T121|3327|RXNORM|DIAZOXIDE|DIAZOXIDE
C0643520|T109|1426427|RXNORM|OLEYL OLEATE|OLEYL OLEATE
C3855118|T121|1547444|RXNORM|CALCIUM ACETATE / MAGNESIUM ACETATE / POTASSIUM ACETATE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM GLUCONATE|CALCIUM ACETATE / MAGNESIUM ACETATE / POTASSIUM ACETATE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM GLUCONATE
C0612804|T109|1308067|RXNORM|ORIGANUM OIL|ORIGANUM OIL
C2928797|T121|1007883|RXNORM|HYDROCORTISONE / SALICYLIC ACID / SODIUM THIOSULFATE|HYDROCORTISONE / SALICYLIC ACID / SODIUM THIOSULFATE
C2928796|T121|1007882|RXNORM|NICARDIPINE / PYRITHIOXIN|NICARDIPINE / PYRITHIOXIN
C2928795|T121|1007881|RXNORM|GINSENG ROOT / SIBERIAN GINSENG ROOT|GINSENG ROOT / SIBERIAN GINSENG ROOT
C0360564|T121|108118|RXNORM|MOMETASONE|MOMETASONE
C0360564|T121|108118|RXNORM|MOMETASONE|MOMETASONE
C0360564|T121|108118|RXNORM|MOMETASONE|MOMETASONE
C2928801|T121|1007887|RXNORM|ASAFETIDA EXTRACT / CAPSICUM EXTRACT / CASCARA SAGRADA / GINGER EXTRACT / NUX VOMICA EXTRACT|ASAFETIDA EXTRACT / CAPSICUM EXTRACT / CASCARA SAGRADA / GINGER EXTRACT / NUX VOMICA EXTRACT
C3256326|T121|1307854|RXNORM|ACHYRANTHES BIDENTATA ROOT EXTRACT|ACHYRANTHES BIDENTATA ROOT EXTRACT
C2928799|T121|1007885|RXNORM|CETYLPYRIDINIUM / DOMIPHEN|CETYLPYRIDINIUM / DOMIPHEN
C2928798|T121|1007884|RXNORM|AMYLASES / ENDOPEPTIDASES / LIPASE / PANCREATIN|AMYLASES / ENDOPEPTIDASES / LIPASE / PANCREATIN
C3465033|T121|1307858|RXNORM|MORINDA CITRIFOLIA LEAF EXTRACT|MORINDA CITRIFOLIA LEAF EXTRACT
C2928803|T121|1007889|RXNORM|PUMPKIN SEED OIL / SAW PALMETTO EXTRACT / ZINC GLUCONATE|PUMPKIN SEED OIL / SAW PALMETTO EXTRACT / ZINC GLUCONATE
C2928802|T121|1007888|RXNORM|CALCIUM CARBONATE / NUX VOMICA EXTRACT / PHENOBARBITAL|CALCIUM CARBONATE / NUX VOMICA EXTRACT / PHENOBARBITAL
C0056058|T109|1367422|RXNORM|COCO-BETAINE|COCO-BETAINE
C3531638|T121|1367423|RXNORM|DIPHENYLTRICHLOROETHANE|DIPHENYLTRICHLOROETHANE
C3859423|T121|1592894|RXNORM|CETYL GLYCOL|CETYL GLYCOL
C0772228|T121|1310546|RXNORM|ACESULFAME|ACESULFAME
C0045818|T121|1310544|RXNORM|2-AMINO-2-METHYL-1-PROPANOL|2-AMINO-2-METHYL-1-PROPANOL
C0043940|T121|1310543|RXNORM|1,3-DIMETHYLOL-5,5-DIMETHYLHYDANTOIN|1,3-DIMETHYLOL-5,5-DIMETHYLHYDANTOIN
C0043904|T121|1310542|RXNORM|1,3-BUTYLENE GLYCOL|1,3-BUTYLENE GLYCOL
C2348061|T130|1310541|RXNORM|D&C RED NO. 21|D&C RED NO. 21
C3859425|T121|1592896|RXNORM|ETHYLHEXYLGLYCERYL BEHENATE|ETHYLHEXYLGLYCERYL BEHENATE
C1509527|T121|1310548|RXNORM|ALKYL (C12-15) BENZOATE|ALKYL (C12-15) BENZOATE
C3486868|T168|1311144|RXNORM|SEPIA OFFICINALIS JUICE EXTRACT|SEPIA OFFICINALIS JUICE
C0071112|T121|1311146|RXNORM|PIPERINE|PIPERINE
C0054673|T130|1311147|RXNORM|DIETHYLENE GLYCOL MONOETHYL ETHER|DIETHYLENE GLYCOL MONOETHYL ETHER
C1533168|T121|1311140|RXNORM|SORBATE|SORBATE
C1875650|T121|689746|RXNORM|PHENOBARBITAL / SODIUM NITRITE|PHENOBARBITAL / SODIUM NITRITE
C3484472|T121|1311143|RXNORM|AJI PEPPER EXTRACT|AJI PEPPER EXTRACT
C3464624|T121|1292776|RXNORM|ASCORBIC ACID / CHOLECALCIFEROL / VITAMIN A|ASCORBIC ACID / CHOLECALCIFEROL / VITAMIN A
C2937462|T121|1311148|RXNORM|LYCOPUS VIRGINICUS EXTRACT|LYCOPUS VIRGINICUS EXTRACT
C0027375|T121|1311149|RXNORM|NAPHTHALENE|NAPHTHALENE
C2726150|T129|974527|RXNORM|THYME ALLERGENIC EXTRACT|THYMUS VULGARIS ALLERGENIC EXTRACT
C0048047|T109|1435279|RXNORM|4-AMINOPHENOL|4-AMINOPHENOL
C0020316|T127|5514|RXNORM|HYDROXOCOBALAMIN|HYDROXOCOBALAMIN
C0020316|T127|5514|RXNORM|HYDROXOCOBALAMIN|HYDROXOCOBALAMIN
C2183076|T121|815449|RXNORM|DEXBROMPHENIRAMINE / PHENYLEPHRINE|DEXBROMPHENIRAMINE / PHENYLEPHRINE
C3486624|T121|1309826|RXNORM|MEDICAGO SATIVA LEAF EXTRACT|MEDICAGO SATIVA LEAF EXTRACT
C3489254|T121|1309827|RXNORM|MORELLA CERIFERA ROOT BARK EXTRACT|MORELLA CERIFERA ROOT BARK EXTRACT
C2928011|T121|1007088|RXNORM|BETAMETHASONE DIPROPIONATE / BETAMETHASONE SODIUM PHOSPHATE|BETAMETHASONE DIPROPIONATE / BETAMETHASONE SODIUM PHOSPHATE
C3486621|T121|1309822|RXNORM|CICHORIUM INTYBUS FLOWER EXTRACT|CICHORIUM INTYBUS FLOWER EXTRACT
C0296800|T121|87636|RXNORM|FEXOFENADINE|FEXOFENADINE
C3488609|T121|1309820|RXNORM|VIBURNUM OPULUS ROOT|VIBURNUM OPULUS ROOT
C2928006|T121|1007083|RXNORM|DILTIAZEM / HYDROCHLOROTHIAZIDE|DILTIAZEM / HYDROCHLOROTHIAZIDE
C2928005|T121|1007082|RXNORM|DIMETHICONE / GLYCERIN|DIMETHICONE / GLYCERIN
C0296806|T130|87639|RXNORM|IOBITRIDOL|IOBITRIDOL
C2928003|T121|1007080|RXNORM|ASCORBIC ACID / CALCIUM CARBONATE / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM OXIDE / NIACINAMIDE / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D / VITAMIN E / ZINC SULFATE|ASCORBIC ACID / CALCIUM CARBONATE / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM OXIDE / NIACINAMIDE / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D / VITAMIN E / ZINC SULFATE
C2928010|T121|1007087|RXNORM|ASCORBIC ACID / BETA CAROTENE / CUPROUS OXIDE / LUTEIN / SODIUM SELENATE / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / BETA CAROTENE / CUPROUS OXIDE / LUTEIN / SODIUM SELENATE / VITAMIN E / ZINC OXIDE
C2928009|T121|1007086|RXNORM|ASCORBIC ACID / FOLIC ACID / NIACIN / PYRIDOXINE / RIBOFLAVIN / SODIUM FLUORIDE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D / VITAMIN E|ASCORBIC ACID / FOLIC ACID / NIACIN / PYRIDOXINE / RIBOFLAVIN / SODIUM FLUORIDE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D / VITAMIN E
C2928008|T121|1007085|RXNORM|ACETAMINOPHEN / CLEMASTINE / PHENYLPROPANOLAMINE|ACETAMINOPHEN / CLEMASTINE / PHENYLPROPANOLAMINE
C2928007|T121|1007084|RXNORM|CHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE / PSEUDOEPHEDRINE / PYRILAMINE|CHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE / PSEUDOEPHEDRINE / PYRILAMINE
C2723651|T129|867232|RXNORM|HELMINTHOSPORIUM SOLANI ALLERGENIC EXTRACT|HELMINTHOSPORIUM SOLANI ALLERGENIC EXTRACT
C0066412|T121|29900|RXNORM|METHYLNICOTINATE|METHYLNICOTINATE
C0002191|T123|535|RXNORM|ALPHA 1-ANTITRYPSIN|ALFA1 ANTITRYPSIN
C0056396|T121|21660|RXNORM|CORTIVAZOL|CORTIVAZOL
C3834237|T121|1543728|RXNORM|AMYLASES / BACILLUS COAGULANS / ENDOPEPTIDASES / LIPASE|AMYLASES / BACILLUS COAGULANS / ENDOPEPTIDASES / LIPASE
C0301434|T121|89831|RXNORM|ZINC PHENOLSULFONATE|ZINC PHENOLSULFONATE
C0058753|T121|23678|RXNORM|DROMOSTANOLONE|DROMOSTANOLONE
C2928476|T121|1007555|RXNORM|ASCORBIC ACID / CHOLECALCIFEROL / SODIUM FLUORIDE / VITAMIN A|ASCORBIC ACID / CHOLECALCIFEROL / SODIUM FLUORIDE / VITAMIN A
C2928148|T121|1007226|RXNORM|CITRIC ACID / TARTARIC ACID|CITRIC ACID / TARTARIC ACID
C2928147|T121|1007225|RXNORM|TRIAMTERENE / XIPAMIDE|TRIAMTERENE / XIPAMIDE
C2928477|T121|1007556|RXNORM|HAEMOPHILUS INFLUENZAE B (ROSS STRAIN) CAPSULAR POLYSACCHARIDE MENINGOCOCCAL PROTEIN CONJUGATE VACCINE / HEPATITIS B SURFACE ANTIGEN VACCINE|HAEMOPHILUS INFLUENZAE B (ROSS STRAIN) CAPSULAR POLYSACCHARIDE MENINGOCOCCAL PROTEIN CONJUGATE VACCINE / HEPATITIS B SURFACE ANTIGEN VACCINE
C2928145|T121|1007223|RXNORM|ACETAMINOPHEN / ADIPHENINE|ACETAMINOPHEN / ADIPHENINE
C2928471|T121|1007550|RXNORM|SALICYLIC ACID / TRICHLOROACETALDEHYDE|SALICYLIC ACID / TRICHLOROACETALDEHYDE
C2928474|T121|1007553|RXNORM|BENZOCAINE / CALAMINE / CAMPHOR|BENZOCAINE / CALAMINE / CAMPHOR
C2928142|T121|1007220|RXNORM|DODECYL SULFATE / LANOLIN|DODECYL SULFATE / LANOLIN
C2918538|T129|995768|RXNORM|CLADOSPORIUM CLADOSPORIOIDES ALLERGENIC EXTRACT|CLADOSPORIUM CLADOSPORIOIDES ALLERGENIC EXTRACT
C2057674|T121|1007559|RXNORM|CHLORTETRACYCLINE / DEMECLOCYCLINE / TETRACYCLINE|CHLORTETRACYCLINE / DEMECLOCYCLINE / TETRACYCLINE
C2928479|T121|1007558|RXNORM|GINGER EXTRACT / PYRIDOXINE|GINGER EXTRACT / PYRIDOXINE
C2928151|T121|1007229|RXNORM|FENBUTRAZATE / PHENMETRAZINE|FENBUTRAZATE / PHENMETRAZINE
C2928150|T121|1007228|RXNORM|ALUMINUM HYDROXIDE / SILICON DIOXIDE|ALUMINUM HYDROXIDE / SILICON DIOXIDE
C0071768|T197|34312|RXNORM|POTASSIUM IODATE|POTASSIUM IODATE
C0163657|T121|59308|RXNORM|CHROMIUM PICOLINATE|CHROMIUM PICOLINATE
C1655488|T121|606797|RXNORM|ACETAMINOPHEN / CAFFEINE / PHENYLTOLOXAMINE / SALICYLAMIDE|ACETAMINOPHEN / CAFFEINE / PHENYLTOLOXAMINE / SALICYLAMIDE
C0033223|T121|8702|RXNORM|PROCARBAZINE|PROCARBAZINE
C0011817|T121|3290|RXNORM|DEXTROMORAMIDE|DEXTROMORAMIDE
C0024200|T195|6513|RXNORM|LYMECYCLINE|LYMECYCLINE
C2701572|T129|852412|RXNORM|JUTE FIBER EXTRACT|CORCORUS CAPSULARIS FIBER EXTRACT
C0048250|T121|15027|RXNORM|4-DIMETHYLAMINOPHENOL|4-DIMETHYLAMINOPHENOL
C0071767|T197|34311|RXNORM|POTASSIUM HYDROXIDE|POTASSIUM HYDROXIDE
C3535678|T196|1368379|RXNORM|SULFIDE ION|SULFIDE ION
C0071701|T131|1541597|RXNORM|POLYVINYL ACETATE|POLYVINYL ACETATE
C3535679|T109|1368378|RXNORM|TERMINALIA BELLIRICA FRUIT EXTRACT|TERMINALIA BELLIRICA FRUIT EXTRACT
C2701600|T129|852491|RXNORM|GREEN ASH POLLEN EXTRACT|FRAXINUS PENNSYLVANICA POLLEN EXTRACT
C0013954|T121|3816|RXNORM|EMEPRONIUM|EMEPRONIUM
C3503280|T121|1370109|RXNORM|VACCINIUM MYRTILLUS WHOLE EXTRACT|VACCINIUM MYRTILLUS WHOLE EXTRACT
C3535647|T109|1370108|RXNORM|DIBUTYL LAUROYL GLUTAMIDE|DIBUTYL LAUROYL GLUTAMIDE
C0072151|T125|34625|RXNORM|PROMESTRIENE|PROMESTRIENE
C0937846|T121|283742|RXNORM|ESOMEPRAZOLE|ESOMEPRAZOLE
C0937844|T121|283740|RXNORM|SWEETLEAF PREPARATION|SWEETLEAF PREPARATION
C3489018|T121|1310131|RXNORM|VISCUM ALBUM FRUIT EXTRACT|VISCUM ALBUM FRUIT EXTRACT
C3535649|T121|1370105|RXNORM|WALTHERIA INDICA LEAF EXTRACT|WALTHERIA INDICA LEAF EXTRACT
C3535650|T121|1370104|RXNORM|FREESIA ALBA FLOWER EXTRACT|FREESIA ALBA FLOWER EXTRACT
C0873118|T121|259453|RXNORM|LEVOBUPIVACAINE|LEVOBUPIVACAINE
C0601355|T121|1366920|RXNORM|CETYL SULFATE|CETYL SULFATE
C0244223|T197|1366921|RXNORM|SODIUM CHLORATE|SODIUM CHLORATE
C0055565|T121|1366924|RXNORM|CHOLESTERYL SULFATE|CHOLESTERYL SULFATE
C1875259|T121|689716|RXNORM|HYDROCHLOROTHIAZIDE / LABETALOL|HYDROCHLOROTHIAZIDE / LABETALOL
C1875258|T121|689714|RXNORM|HYDRALAZINE / RESERPINE|HYDRALAZINE / RESERPINE
C0772051|T130|177906|RXNORM|SAMARIUM SM 153 LEXIDRONAM|SAMARIUM (153SM) LEXDRONAM
C1720478|T121|712584|RXNORM|ALDIOXA / CHLOROXYLENOL|ALDIOXA / CHLOROXYLENOL
C0058702|T121|23638|RXNORM|DOPEXAMINE|DOPEXAMINE
C0028476|T121|7543|RXNORM|NOXYTHIOLIN|NOXYTHIOLIN
C2701384|T130|905276|RXNORM|GERMAN COCKROACH ALLERGENIC EXTRACT|BLATTELLA GERMANICA ALLERGENIC EXTRACT
C3474466|T109|1307684|RXNORM|EUCALYPTUS POLYBRACTEA LEAF OIL|EUCALYPTUS POLYBRACTEA LEAF OIL
C0376261|T121|114202|RXNORM|LACTATE|LACTATE
C0376261|T121|114202|RXNORM|LACTATE|LACTATE
C0376261|T121|114202|RXNORM|LACTATE|LACTATE
C0376261|T121|114202|RXNORM|LACTATE|LACTATE
C3465254|T109|1307686|RXNORM|CEDRUS DEODARA WOOD OIL|CEDRUS DEODARA WOOD OIL
C3255608|T121|1307687|RXNORM|PUERARIA MONTANA VAR. CHINENSIS ROOT EXTRACT|PUERARIA MONTANA VAR. CHINENSIS ROOT EXTRACT
C3256330|T109|1307680|RXNORM|AMINOMETHYL PROPANEDIOL|AMINOMETHYL PROPANEDIOL
C3255955|T109|1307681|RXNORM|MANGO SEED OIL|MANGO SEED OIL
C3256680|T109|1307682|RXNORM|GALANGAL OIL|GALANGAL OIL
C3255733|T109|1307683|RXNORM|HYDROGENATED COCONUT OIL|HYDROGENATED COCONUT OIL
C3535632|T121|1370465|RXNORM|BOS TAURUS NASAL MUCOSA PREPARATION|BOVINE NASAL MUCOSA PREPARATION
C2827497|T109|1307688|RXNORM|POLYOXYL 60 HYDROGENATED CASTOR OIL|PEG-60 HYDROGENATED CASTOR OIL
C3255961|T109|1307689|RXNORM|PAPRIKA OIL|PAPRIKA OIL
C0053947|T121|19610|RXNORM|BORNAPRINE|BORNAPRINE
C1874158|T121|690990|RXNORM|ALUMINUM ACETATE / ZINC OXIDE|ALUMINUM ACETATE / ZINC OXIDE
C3192263|T121|1147220|RXNORM|VEMURAFENIB|VEMURAFENIB
C1874164|T121|690996|RXNORM|ALUMINUM HYDROXIDE / ASPIRIN / CODEINE / MAGNESIUM HYDROXIDE|ALUMINUM HYDROXIDE / ASPIRIN / CODEINE / MAGNESIUM HYDROXIDE
C0030946|T126|8031|RXNORM|ENDOPEPTIDASES|ENDOPEPTIDASES
C1328025|T129|1298944|RXNORM|PERTUZUMAB|PERTUZUMAB
C1321284|T121|687323|RXNORM|EPINEPHRINE / GUANETHIDINE|EPINEPHRINE / GUANETHIDINE
C3859661|T121|1593610|RXNORM|SPINACIA OLERACEA ROOT EXTRACT|SPINACIA OLERACEA ROOT EXTRACT
C3859662|T121|1593611|RXNORM|ARGANIA SPINOSA LEAF EXTRACT|ARGANIA SPINOSA LEAF EXTRACT
C3555459|T121|1421149|RXNORM|BOS TAURUS PROSTATE GLAND PREPARATION|BOVINE PROSTATE GLAND PREPARATION
C0041928|T196|10999|RXNORM|URANIUM|URANIUM
C0041920|T121|10996|RXNORM|URACIL MUSTARD|URACIL MUSTARD
C0041917|T123|10995|RXNORM|URACIL|URACIL
C3859664|T121|1593618|RXNORM|ACETAMINOPHEN / CHLOPHEDIANOL / PYRILAMINE|ACETAMINOPHEN / CHLOPHEDIANOL / PYRILAMINE
C0168273|T121|60819|RXNORM|BIVALIRUDIN|BIVALIRUDIN
C0041738|T121|10991|RXNORM|UNITHIOL|UNITHIOL
C0057946|T109|1429928|RXNORM|DIETHYLENE GLYCOL|DIETHYLENE GLYCOL
C1170748|T121|353110|RXNORM|FIBRINOLYSIS INHIBITOR|FIBRINOLYSIS INHIBITOR
C0059871|T121|24611|RXNORM|ETOFYLLINE|ETOFYLLINE
C3651740|T121|1429926|RXNORM|CANNABIS SATIVA SEED EXTRACT|CANNABIS SATIVA SEED EXTRACT
C3651739|T121|1429927|RXNORM|CHAMAECYPARIS OBTUSA WHOLE EXTRACT|CHAMAECYPARIS OBTUSA WHOLE EXTRACT
C3465034|T121|1307539|RXNORM|MORUS NIGRA ROOT EXTRACT|MORUS NIGRA ROOT EXTRACT
C0055752|T121|21130|RXNORM|CINNAMEDRINE|CINNAMEDRINE
C0060282|T197|24947|RXNORM|FERROUS SULFATE|FERROUS SULFATE
C0060277|T121|24942|RXNORM|FERROUS GLUCONATE|FERROUS GLUCONATE
C0060275|T197|24940|RXNORM|FERROUS CHLORIDE|FERROUS CHLORIDE
C0060276|T121|24941|RXNORM|FERROUS FUMARATE|FERROUS FUMARATE
C2701470|T129|852276|RXNORM|GAMBELS OAK POLLEN EXTRACT|QUERCUS GAMBELII POLLEN EXTRACT
C0717555|T121|214358|RXNORM|CARAMIPHEN / PHENYLPROPANOLAMINE|CARAMIPHEN / PHENYLPROPANOLAMINE
C0981937|T129|852272|RXNORM|PECAN POLLEN EXTRACT|PECAN POLLEN EXTRACT
C0771946|T125|236646|RXNORM|INSULIN, PROTAMINE ZINC, HUMAN|INSULIN, PROTAMINE ZINC, HUMAN
C0077539|T121|38998|RXNORM|TYLOXAPOL|TYLOXAPOL
C0717546|T121|214350|RXNORM|CALCIUM GLYCEROPHOSPHATE / CALCIUM LACTATE|CALCIUM GLYCEROPHOSPHATE / CALCIUM LACTATE
C0717551|T129|214355|RXNORM|CANDIDA ALBICANS EXTRACT|YEAST EXTRACT
C0717550|T121|214354|RXNORM|CANDESARTAN|CANDESARTAN
C0717554|T121|214357|RXNORM|CAPTOPRIL / HYDROCHLOROTHIAZIDE|CAPTOPRIL / HYDROCHLOROTHIAZIDE
C1831808|T121|1364430|RXNORM|APIXABAN|APIXABAN
C0772192|T121|236867|RXNORM|OCTODRINE|OCTODRINE
C0007641|T126|2219|RXNORM|CELLULASE|CELLULASE
C0068788|T121|31819|RXNORM|NITAZOXANIDE|NITAZOXANIDE
C0771939|T121|236641|RXNORM|CAPSELLA BURSA-PASTORIS EXTRACT|CAPSELLA BURSA-PASTORIS EXTRACT
C2730220|T129|892604|RXNORM|CASEIN (COW MILK) ALLERGENIC EXTRACT|CASEIN (COW MILK) ALLERGENIC EXTRACT
C0022616|T121|6131|RXNORM|KETANSERIN|KETANSERIN
C0663733|T121|190548|RXNORM|TIPRANAVIR|TIPRANAVIR
C0058961|T121|23852|RXNORM|EFLOXATE|EFLOXATE
C0527038|T121|135313|RXNORM|ISOPROPYL UNOPROSTONE|ISOPROPYL UNOPROSTONE
C0054417|T197|1368199|RXNORM|CADMIUM SULFIDE|CADMIUM SULFIDE
C0043773|T121|1368198|RXNORM|1,2-BENZISOTHIAZOLINE-3-ONE|1,2-BENZISOTHIAZOLINE-3-ONE
C3256842|T109|1368193|RXNORM|GLYCERYL LINOLEATE|GLYCERYL LINOLEATE
C3486815|T121|1328310|RXNORM|ORNITHOGALUM UMBELLATUM EXTRACT|ORNITHOGALUM UMBELLATUM EXTRACT
C3488312|T121|1328313|RXNORM|THYMUS SERPYLLUM EXTRACT|THYMUS SERPYLLUM EXTRACT
C3487991|T121|1328312|RXNORM|CONIUM MACULATUM FLOWERING TOP EXTRACT|CONIUM MACULATUM FLOWERING TOP EXTRACT
C3488964|T109|1328315|RXNORM|PORPHYRIDIUM PURPUREUM EXTRACT|PORPHYRIDIUM PURPUREUM EXTRACT
C2961423|T121|1368196|RXNORM|HARD FAT|HARD FAT
C3267547|T121|1368195|RXNORM|DIETHYLHEXYL SYRINGYLIDENEMALONATE|DIETHYLHEXYL SYRINGYLIDENEMALONATE
C3257700|T109|1368194|RXNORM|1-ETHYL-2-PYRROLECARBOXALDEHYDE|1-ETHYL-2-PYRROLECARBOXALDEHYDE
C1321946|T121|402527|RXNORM|CHLORPHENINDIONE|CHLORPHENINDIONE
C0060477|T121|25096|RXNORM|FLUBENDAZOLE|FLUBENDAZOLE
C2344291|T129|798262|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 11 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 11 VACCINE
C0610988|T121|162592|RXNORM|DIETHYLAMINE SALICYLATE|DIETHYLAMINE SALICYLATE
C0016410|T127|4511|RXNORM|FOLIC ACID|FOLIC ACID
C2980923|T129|1094193|RXNORM|BROOMWEED POLLEN EXTRACT|AMPHIACHYRIS DRACUNCULOIDES POLLEN EXTRACT
C3256278|T109|1424672|RXNORM|C12-20 ALKYL GLUCOSIDE|C12-20 ALKYL GLUCOSIDE
C0043832|T121|11645|RXNORM|DEFERIPRONE|DEFERIPRONE
C3695981|T109|1483231|RXNORM|KARUM SEED OIL|KARUM SEED OIL
C3695980|T109|1483232|RXNORM|OCTYLDODECYL OLEATE|OCTYLDODECYL OLEATE
C3714887|T121|1492183|RXNORM|HYDROXYETHYL CELLULOSE (280 MPA.S AT 2%)|HYDROXYETHYL CELLULOSE (280 MPA.S AT 2%)
C0019392|T127|5281|RXNORM|HESPERIDIN|HESPERIDIN
C3281529|T121|1307702|RXNORM|MUSA X PARADISIACA LEAF EXTRACT|MUSA X PARADISIACA LEAF EXTRACT
C0012004|T130|3319|RXNORM|DIATRIZOATE|DIATRIZOATE
C0076793|T121|38372|RXNORM|TOLCICLATE|TOLCICLATE
C0128513|T121|52769|RXNORM|MILRINONE|MILRINONE
C3486846|T121|1311354|RXNORM|SUS SCROFA TOOTH PREPARATION|PORCINE TOOTH PREPARATION
C3813564|T121|1539684|RXNORM|LEONTOPODIUM ALPINUM EXTRACT|LEONTOPODIUM NIVALE SUBSP. ALPINUM WHOLE FLOWERING EXTRACT
C0064007|T121|27946|RXNORM|ISOMETHEPTENE|ISOMETHEPTENE
C1531015|T121|498509|RXNORM|PEGAPTANIB|PEGAPTANIB
C3537762|T121|1371443|RXNORM|2,2,2-TRIFLUOROACETOPHENONE|2,2,2-TRIFLUOROACETOPHENONE
C3474470|T121|1310048|RXNORM|HELICHRYSUM ITALICUM FLOWER EXTRACT|HELICHRYSUM ITALICUM FLOWER EXTRACT
C2351132|T121|817579|RXNORM|ACETAMINOPHEN / CODEINE|ACETAMINOPHEN / CODEINE
C2718773|T129|853491|RXNORM|CANAKINUMAB|CANAKINUMAB
C1166208|T121|350488|RXNORM|SERENOA PREPARATION|SERENOA PREPARATION
C0074554|T121|36567|RXNORM|SIMVASTATIN|SIMVASTATIN
C3486573|T121|1310043|RXNORM|CICUTA VIROSA ROOT EXTRACT|CICUTA VIROSA ROOT EXTRACT
C0937879|T121|1310040|RXNORM|MILLET EXTRACT|MILLET EXTRACT
C3162669|T121|1114601|RXNORM|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / CHOLINE / FERROUS FUMARATE / FOLIC ACID / NIACIN / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / CHOLINE / FERROUS FUMARATE / FOLIC ACID / NIACIN / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN E / ZINC OXIDE
C3495652|T121|1310046|RXNORM|SESAME SEED EXTRACT|SESAME SEED EXTRACT
C3474163|T109|1310047|RXNORM|NELUMBO NUCIFERA FLOWER OIL|NELUMBO NUCIFERA FLOWER OIL
C3474158|T168|1310044|RXNORM|CASHEW OIL|CASHEW OIL
C3486727|T121|1310045|RXNORM|LARIX DECIDUA FLOWERING TOP EXTRACT|LARIX DECIDUA FLOWERING TOP EXTRACT
C3500189|T109|1313968|RXNORM|POLYQUATERNIUM-51 (2-METHACRYLOYLOXYETHYL PHOSPHORYLCHOLINE-N-BUTYL METHACRYLATE; 4:1)|POLYQUATERNIUM-51 (2-METHACRYLOYLOXYETHYL PHOSPHORYLCHOLINE-N-BUTYL METHACRYLATE; 4:1)
C0087163|T127|42955|RXNORM|LEVOCARNITINE|LEVOCARNITINE
C0087162|T127|42954|RXNORM|VITAMIN B6|VITAMIN B6
C3537766|T121|1371447|RXNORM|DIMETHICONE PEG-10 PHOSPHATE|DIMETHICONE PEG-10 PHOSPHATE
C3537765|T121|1371446|RXNORM|GLYCERETH-7 TRIMETHYL ETHER|GLYCERETH-7 TRIMETHYL ETHER
C1629836|T007|602811|RXNORM|LACTOBACILLUS RHAMNOSUS GG|LACTOBACILLUS RHAMNOSUS GG
C0063449|T121|27492|RXNORM|INDANAZOLINE|INDANAZOLINE
C3531674|T109|1367499|RXNORM|STEARYL TRIETHOXYSILANE|STEARYL TRIETHOXYSILANE
C3531673|T109|1367498|RXNORM|POLYGLYCERYL-3 DISTEARATE|POLYGLYCERYL-3 DISTEARATE
C0533545|T195|138099|RXNORM|GEMIFLOXACIN|GEMIFLOXACIN
C0035891|T195|9478|RXNORM|ROXITHROMYCIN|ROXITHROMYCIN
C2702401|T129|1098619|RXNORM|TRICHOPHYTON TONSURANS ALLERGENIC EXTRACT|TRICHOPHYTON TONSURANS ALLERGENIC EXTRACT
C3864855|T121|1594930|RXNORM|PORTULACA GRANDIFLORA WHOLE EXTRACT|PORTULACA GRANDIFLORA WHOLE EXTRACT
C3864854|T121|1594931|RXNORM|PORTULACA GRANDIFLORA SEED EXTRACT|PORTULACA GRANDIFLORA SEED EXTRACT
C3853574|T121|1594933|RXNORM|MENTHA SPICATA EXTRACT|MENTHA SPICATA EXTRACT
C3488949|T121|1322552|RXNORM|ANGOSTURA BARK EXTRACT|ANGOSTURA BARK EXTRACT
C3531671|T109|1367495|RXNORM|PEG-7 METHYL ETHER|PEG-7 METHYL ETHER
C1871004|T121|715869|RXNORM|MAROPITANT|MAROPITANT
C3531670|T109|1367494|RXNORM|OCTADECENE|OCTADECENE
C2194290|T121|820299|RXNORM|CITRIC ACID / SODIUM BICARBONATE|CITRIC ACID / SODIUM BICARBONATE
C0034295|T121|9020|RXNORM|PYRITHIOXIN|PYRITHIOXIN
C3256848|T109|1426922|RXNORM|LAURYL LAURATE|LAURYL LAURATE
C0034303|T130|9022|RXNORM|PYROGALLOL|PYROGALLOL
C3255887|T197|1305556|RXNORM|ALUMINUM HYDRATE|ALUMINUM HYDRATE
C2344347|T129|798372|RXNORM|MUMPS VIRUS VACCINE LIVE, JERYL LYNN STRAIN|MUMPS VIRUS VACCINE LIVE, JERYL LYNN STRAIN
C2928684|T121|1007769|RXNORM|BISMUTH SUBCITRATE / METRONIDAZOLE / TETRACYCLINE|BISMUTH SUBCITRATE / METRONIDAZOLE / TETRACYCLINE
C2928861|T121|1007948|RXNORM|CLIOQUINOL / PHTHALYLSULFATHIAZOLE|CLIOQUINOL / PHTHALYLSULFATHIAZOLE
C2928862|T121|1007949|RXNORM|CINAMETIC ACID / METOCLOPRAMIDE / SIMETHICONE|CINAMETIC ACID / METOCLOPRAMIDE / SIMETHICONE
C2928677|T121|1007762|RXNORM|HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / THREONINE / TRYPTOPHAN / VALINE|HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / THREONINE / TRYPTOPHAN / VALINE
C2928678|T121|1007763|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL / SOYBEAN PREPARATION|CALCIUM CARBONATE / CHOLECALCIFEROL / SOYBEAN PREPARATION
C2928675|T121|1007760|RXNORM|COENZYME Q10 / FOLIC ACID / VITAMIN B 12 / VITAMIN B6|COENZYME Q10 / FOLIC ACID / VITAMIN B 12 / VITAMIN B6
C2928676|T121|1007761|RXNORM|EFAVIRENZ / EMTRICITABINE / TENOFOVIR DISOPROXIL|EFAVIRENZ / EMTRICITABINE / TENOFOVIR DISOPROXIL
C2928681|T121|1007766|RXNORM|CHLORPHENIRAMINE / DIPYRONE|CHLORPHENIRAMINE / DIPYRONE
C2928682|T121|1007767|RXNORM|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PSEUDOEPHEDRINE / SCOPOLAMINE|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PSEUDOEPHEDRINE / SCOPOLAMINE
C2928679|T121|1007764|RXNORM|CHROMIUM PICOLINATE / NIACIN|CHROMIUM PICOLINATE / NIACIN
C2928680|T121|1007765|RXNORM|CHLORPHENIRAMINE / EPHEDRINE / OXOLAMINE|CHLORPHENIRAMINE / EPHEDRINE / OXOLAMINE
C0038744|T121|10206|RXNORM|SULFISOMIDINE|SULFISOMIDINE
C0038745|T121|10207|RXNORM|SULFISOXAZOLE|SULFISOXAZOLE
C0038745|T121|10207|RXNORM|SULFISOXAZOLE|SULFISOXAZOLE
C0038742|T121|10205|RXNORM|SULFINPYRAZONE|SULFINPYRAZONE
C3281528|T121|1426928|RXNORM|GLYCERYL PALMITATE|GLYCERYL PALMITATE
C1874741|T121|691366|RXNORM|CASTOR OIL / PERUVIAN BALSAM / TRYPSIN|CASTOR OIL / PERUVIAN BALSAM / TRYPSIN
C3256588|T109|1305553|RXNORM|ADENOPHORA STRICTA ROOT EXTRACT|ADENOPHORA STRICTA ROOT EXTRACT
C2728191|T129|1010954|RXNORM|LICORICE ALLERGENIC EXTRACT|LICORICE ALLERGENIC EXTRACT
C0644503|T121|180806|RXNORM|BUTALAMINE|BUTALAMINE
C0359958|T121|107610|RXNORM|COCAINE / HOMATROPINE|COCAINE / HOMATROPINE
C0937908|T121|1364288|RXNORM|ECHINACEA PALLIDA PREPARATION|ECHINACEA PALLIDA PREPARATION
C2981254|T004|1329940|RXNORM|ASPERGILLUS FLAVUS VAR. ORYZAE|ASPERGILLUS FLAVUS VAR. ORYZAE
C0982067|T109|1425217|RXNORM|CERESIN|CERESIN
C3484454|T121|1353217|RXNORM|NUTMEG EXTRACT|NUTMEG EXTRACT
C0076040|T121|37744|RXNORM|TEFERROL|IRON POLYMALTOSE
C1313616|T121|1370971|RXNORM|OSPEMIFENE|OSPEMIFENE
C3695963|T121|1484279|RXNORM|CUCUMIS SATIVUS WHOLE EXTRACT|CUCUMIS SATIVUS WHOLE EXTRACT
C0040829|T121|1484278|RXNORM|TRENBOLONE|TRENBOLONE
C3488473|T121|1426870|RXNORM|MOSCHUS MOSCHIFERUS MUSK SAC RESIN|MOSCHUS MOSCHIFERUS MUSK SAC RESIN
C0937596|T121|283538|RXNORM|ANTHRAQUINONE GLYCOSIDE|ANTHRAQUINONE GLYCOSIDE
C3486304|T121|1426678|RXNORM|C12-14 PARETH-3|C12-14 PARETH-3
C0032836|T121|8602|RXNORM|POTASSIUM OROTATE|POTASSIUM OROTATE
C0937595|T121|283537|RXNORM|ANAMU PREPARATION|ANAMU PREPARATION
C0058978|T121|1304974|RXNORM|ICOSAPENT ETHYL|ICOSAPENT ETHYL
C0032841|T121|8606|RXNORM|POTASSIUM SORBATE|POTASSIUM SORBATE
C0032838|T197|8604|RXNORM|POTASSIUM PERMANGANATE|POTASSIUM PERMANGANATE
C0026187|T195|6980|RXNORM|MINOCYCLINE|MINOCYCLINE
C0026187|T195|6980|RXNORM|MINOCYCLINE|MINOCYCLINE
C3159366|T129|1111024|RXNORM|VALLEY OAK POLLEN EXTRACT|QUERCUS LOBATA POLLEN EXTRACT
C2723639|T129|867218|RXNORM|DOGFENNEL POLLEN EXTRACT|EUPATORIUM CAPILLIFOLIUM POLLEN EXTRACT
C3864843|T121|1595884|RXNORM|SODIUM PROPOXYHYDROXYPROPYL THIOSULFATE SILICA|SODIUM PROPOXYHYDROXYPROPYL THIOSULFATE SILICA
C0078023|T197|39364|RXNORM|VANADYL SULFATE|VANADYL SULFATE
C2929680|T121|1008781|RXNORM|5-HYDROXYTRYPTOPHAN / VITAMIN B6|5-HYDROXYTRYPTOPHAN / VITAMIN B6
C2929679|T121|1008780|RXNORM|CHONDROITIN SULFATES / PAPAIN|CHONDROITIN SULFATES / PAPAIN
C2929682|T121|1008783|RXNORM|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / POLYSACCHARIDE IRON COMPLEX|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / POLYSACCHARIDE IRON COMPLEX
C2929681|T121|1008782|RXNORM|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC / THREONINE / TRYPTOPH|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929684|T121|1008785|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 1 VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 10A VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 11A VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 12F VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHAR|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 1 VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 10A VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 11A VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 12F VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 14 VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 15B VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 17F VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 18C VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 19A VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 19F VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 2 VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 20 VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 22F VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 23F VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 3 VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 33F VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 4 VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 5 VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 6B VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 7F VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 8 VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 9N VACCINE / PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 9V VACCINE
C2929683|T121|1008784|RXNORM|MAGNESIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE|MAGNESIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE
C2929686|T121|1008787|RXNORM|BENZOCAINE / CAPSAICIN / MENTHOL / METHYL SALICYLATE|BENZOCAINE / CAPSAICIN / MENTHOL / METHYL SALICYLATE
C2929685|T121|1008786|RXNORM|DIPYRONE / PROPOXYPHENE|DIPYRONE / PROPOXYPHENE
C2929688|T121|1008789|RXNORM|EFAVIRENZ / LAMIVUDINE / TENOFOVIR DISOPROXIL|EFAVIRENZ / LAMIVUDINE / TENOFOVIR DISOPROXIL
C2929687|T121|1008788|RXNORM|BENZOATE / HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / PHENYL SALICYLATE|BENZOATE / HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / PHENYL SALICYLATE
C3651782|T121|1428418|RXNORM|FRAXINUS AMERICANA BARK EXTRACT|FRAXINUS AMERICANA BARK EXTRACT
C0047828|T121|14699|RXNORM|DIHYDROXYBUTYL ETHER|DIHYDROXYBUTYL ETHER
C3281701|T109|1426671|RXNORM|UNDECYLENOYL GLYCINE|UNDECYLENOYL GLYCINE
C3488255|T121|1426670|RXNORM|VESPA CRABRO PREPARATION|VESPA CRABRO PREPARATION
C0034245|T131|8991|RXNORM|PYRETHRINS|PYRETHRINS
C0003442|T129|1011|RXNORM|LYMPHOCYTE IMMUNE GLOBULIN, ANTI-THYMOCYTE GLOBULIN|LYMPHOCYTE IMMUNE GLOBULIN, ANTI-THYMOCYTE GLOBULIN
C3530628|T121|1364987|RXNORM|CARICA PAPAYA WHOLE EXTRACT|CARICA PAPAYA WHOLE EXTRACT
C2727825|T129|889548|RXNORM|COTTON ALLERGENIC EXTRACT|GOSSYPIUM HIRSUTUM ALLERGENIC EXTRACT
C3496736|T109|1426675|RXNORM|SYNTHETIC WAX (1800 MW)|SYNTHETIC WAX (1800 MW)
C3539943|T121|1428412|RXNORM|ALTHAEA OFFICINALIS WHOLE EXTRACT|ALTHAEA OFFICINALIS WHOLE EXTRACT
C1871020|T121|1313706|RXNORM|HEXYL DECANOATE|HEXYL DECANOATE
C2726192|T129|966995|RXNORM|PHOMA DESTRUCTIVA ALLERGENIC EXTRACT|PHOMA DESTRUCTIVA ALLERGENIC EXTRACT
C2981326|T168|1310511|RXNORM|HIGH FRUCTOSE CORN SYRUP|HIGH FRUCTOSE CORN SYRUP
C3497847|T197|1426676|RXNORM|TRIMETHYLSILOXYSILICATE (M-Q 0.8-1.0)|TRIMETHYLSILOXYSILICATE (M-Q 0.8-1.0)
C3495099|T121|1342649|RXNORM|ADONIS VERNALIS EXTRACT|ADONIS VERNALIS EXTRACT
C0041942|T123|11002|RXNORM|UREA|UREA
C0041942|T123|11002|RXNORM|UREA|UREA
C0041942|T123|11002|RXNORM|UREA|UREA
C2929166|T121|1008259|RXNORM|CYSTINE / VITAMIN B6|CYSTINE / VITAMIN B6
C3255811|T122|1310513|RXNORM|SORBITAN ISOSTEARATE|SORBITAN ISOSTEARATE
C2981012|T121|1094349|RXNORM|DEXTROMETHORPHAN / DOXYLAMINE / PSEUDOEPHEDRINE|DEXTROMETHORPHAN / DOXYLAMINE / PSEUDOEPHEDRINE
C3833238|T109|1540880|RXNORM|CISTUS LADANIFER RESIN|CISTUS LADANIFER RESIN
C2929159|T121|1008252|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / DIPHENHYDRAMINE|ACETAMINOPHEN / DEXTROMETHORPHAN / DIPHENHYDRAMINE
C2929158|T121|1008251|RXNORM|BETAINE / IODINE / PAPAIN / PEPSIN A|BETAINE / IODINE / PAPAIN / PEPSIN A
C2929157|T121|1008250|RXNORM|ASCORBIC ACID / QUERCETIN|ASCORBIC ACID / QUERCETIN
C2929164|T121|1008257|RXNORM|AMINOPHYLLINE / EPHEDRINE / POTASSIUM IODIDE|AMINOPHYLLINE / EPHEDRINE / POTASSIUM IODIDE
C2929163|T121|1008256|RXNORM|BROMPHENIRAMINE / DIHYDROCODEINE / PSEUDOEPHEDRINE|BROMPHENIRAMINE / DIHYDROCODEINE / PSEUDOEPHEDRINE
C2929162|T121|1008255|RXNORM|BROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE|BROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE
C2929161|T121|1008254|RXNORM|ALANINE / ARGININE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929161|T121|1008254|RXNORM|ALANINE / ARGININE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2949213|T121|1046220|RXNORM|BENZALKONIUM / MENTHOL / PETROLATUM|BENZALKONIUM / MENTHOL / PETROLATUM
C3864830|T129|1596932|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 45 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 45 VACCINE
C0001927|T121|435|RXNORM|ALBUTEROL|ALBUTEROL
C0001927|T121|435|RXNORM|ALBUTEROL|ALBUTEROL
C3834051|T121|1543411|RXNORM|FRITILLARIA DELAVAYI BULB EXTRACT|FRITILLARIA DELAVAYI BULB EXTRACT
C0001911|T121|430|RXNORM|ALBENDAZOLE|ALBENDAZOLE
C2194161|T121|819659|RXNORM|ASPIRIN / PAPAIN|ASPIRIN / PAPAIN
C0981911|T129|852519|RXNORM|HOUSE DUST EXTRACT|HOUSE DUST EXTRACT
C2193905|T121|818431|RXNORM|MERSALYL / THEOPHYLLINE|MERSALYL / THEOPHYLLINE
C2701257|T129|852046|RXNORM|NETTLE POLLEN EXTRACT|URTICA DIOICA POLLEN EXTRACT
C2701617|T129|852514|RXNORM|VELVET GRASS POLLEN EXTRACT|HOLCUS LANATUS POLLEN EXTRACT
C2929235|T121|1008330|RXNORM|NORMETHADONE / OXILOFRINE|NORMETHADONE / OXILOFRINE
C2929236|T121|1008331|RXNORM|DIPHENHYDRAMINE / METHAQUALONE|DIPHENHYDRAMINE / METHAQUALONE
C2929237|T121|1008332|RXNORM|SULFADIAZINE / TETROXOPRIM|SULFADIAZINE / TETROXOPRIM
C2929238|T121|1008333|RXNORM|ASCORBIC ACID / FOLIC ACID|ASCORBIC ACID / FOLIC ACID
C2929239|T121|1008334|RXNORM|BENZOCAINE / SULFUR|BENZOCAINE / SULFUR
C2929240|T121|1008335|RXNORM|BENZOCAINE / TANNIC ACID|BENZOCAINE / TANNIC ACID
C2929241|T121|1008336|RXNORM|MEPHENESIN / PHENYLBUTAZONE|MEPHENESIN / PHENYLBUTAZONE
C2929243|T121|1008338|RXNORM|CAPSAICIN / LIDOCAINE|CAPSAICIN / LIDOCAINE
C2929244|T121|1008339|RXNORM|GLUCOSAMINE / S-ADENOSYLMETHIONINE|GLUCOSAMINE / S-ADENOSYLMETHIONINE
C0633482|T121|174965|RXNORM|MYRTOL|MYRTOL
C0019497|T121|5321|RXNORM|HEXYLRESORCINOL|HEXYLRESORCINOL
C3255843|T121|1311608|RXNORM|HOVENIA DULCIS FRUIT EXTRACT|HOVENIA DULCIS FRUIT EXTRACT
C3700987|T109|1486024|RXNORM|HYDROXYCAPRYLATE|HYDROXYCAPRYLATE
C3665206|T121|1435518|RXNORM|7-BEHENOYLSTEARATE|7-BEHENOYLSTEARATE
C3665207|T121|1435519|RXNORM|DIMETHYLMETHOXY CHROMANYL PALMITATE|DIMETHYLMETHOXY CHROMANYL PALMITATE
C0717839|T121|214633|RXNORM|HYDROCODONE / PHENYLEPHRINE / PYRILAMINE|HYDROCODONE / PHENYLEPHRINE / PYRILAMINE
C0717837|T121|214631|RXNORM|HYDROCODONE / PSEUDOEPHEDRINE|HYDROCODONE / PSEUDOEPHEDRINE
C3464710|T121|1312556|RXNORM|DIMETHOXY DI-P-CRESOL|DIMETHOXY DI-P-CRESOL
C3282036|T121|1312557|RXNORM|DIPALMITOYLETHYL HYDROXYETHYLMONIUM METHOSULFATE|DIPALMITOYLETHYL HYDROXYETHYLMONIUM METHOSULFATE
C3256171|T109|1307050|RXNORM|METHYL DIHYDROJASMONATE|METHYL DIHYDROJASMONATE
C3496831|T121|1312558|RXNORM|DIPHENYLSILOXY PHENYL TRIMETHICONE|DIPHENYLSILOXY PHENYL TRIMETHICONE
C3256834|T121|1312559|RXNORM|DIPROPYLENE GLYCOL CAPRATE-CAPRYLATE DIESTER|DIPROPYLENE GLYCOL CAPRATE-CAPRYLATE DIESTER
C2093620|T129|904554|RXNORM|KARAYA GUM ALLERGENIC EXTRACT|KARAYA GUM ALLERGENIC EXTRACT
C2724975|T121|880446|RXNORM|CODEINE / PSEUDOEPHEDRINE / PYRILAMINE|CODEINE / PSEUDOEPHEDRINE / PYRILAMINE
C3651747|T122|1429043|RXNORM|BIS-HYDROXYETHOXYPROPYL DIMETHICONE (37 CST)|BIS-HYDROXYETHOXYPROPYL DIMETHICONE (37 CST)
C3257425|T121|1307668|RXNORM|FILIPENDULA ULMARIA LEAF EXTRACT|FILIPENDULA ULMARIA LEAF EXTRACT
C2920773|T129|999408|RXNORM|ASPERGILLUS TERREUS EXTRACT|ASPERGILLUS TERREUS EXTRACT
C3864831|T129|1596931|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 33 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 33 VACCINE
C3256501|T121|1307669|RXNORM|ARISAEMA ERUBESCENS ROOT EXTRACT|ARISAEMA ERUBESCENS ROOT EXTRACT
C0065152|T121|28863|RXNORM|LOFEXIDINE|LOFEXIDINE
C1134467|T121|337068|RXNORM|METHYL 5-AMINOLEVULINATE|METHYL AMINOLEVULINATE
C0033702|T007|1316073|RXNORM|PROTEUS VULGARIS|PROTEUS VULGARIS
C1615680|T121|581550|RXNORM|CITRUS PECTIN EXTRACT|CITRUS PECTIN EXTRACT
C0538777|T123|140502|RXNORM|ANCESTIM|ANCESTIM
C0036956|T007|1316076|RXNORM|SHIGELLA DYSENTERIAE|SHIGELLA DYSENTERIAE
C0717374|T121|214188|RXNORM|ACETAMINOPHEN / SALICYLAMIDE|ACETAMINOPHEN / SALICYLAMIDE
C2037256|T121|813667|RXNORM|CLORAZEPATE / SULPIRIDE|CLORAZEPATE / SULPIRIDE
C3256428|T121|1307663|RXNORM|PINELLIA TERNATA ROOT EXTRACT|PINELLIA TERNATA ROOT EXTRACT
C0717369|T121|214184|RXNORM|ACETAMINOPHEN / PAMABROM|ACETAMINOPHEN / PAMABROM
C0717370|T121|214185|RXNORM|ACETAMINOPHEN / PENTAZOCINE|ACETAMINOPHEN / PENTAZOCINE
C0717371|T121|214186|RXNORM|ACETAMINOPHEN / PHENYLEPHRINE|ACETAMINOPHEN / PHENYLEPHRINE
C0717373|T121|214187|RXNORM|ACETAMINOPHEN / PSEUDOEPHEDRINE|ACETAMINOPHEN / PSEUDOEPHEDRINE
C0717365|T121|214180|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN|ACETAMINOPHEN / DEXTROMETHORPHAN
C0717366|T121|214181|RXNORM|ACETAMINOPHEN / DIPHENHYDRAMINE|ACETAMINOPHEN / DIPHENHYDRAMINE
C0717367|T121|214182|RXNORM|ACETAMINOPHEN / HYDROCODONE|ACETAMINOPHEN / HYDROCODONE
C0717368|T121|214183|RXNORM|ACETAMINOPHEN / OXYCODONE|ACETAMINOPHEN / OXYCODONE
C3465006|T121|1307661|RXNORM|AZADIRACHTA INDICA BARK EXTRACT|AZADIRACHTA INDICA BARK EXTRACT
C3487958|T121|1309699|RXNORM|LACTUCA VIROSA LEAF EXTRACT|LACTUCA VIROSA LEAF EXTRACT
C1663809|T109|1426289|RXNORM|TRIDECYL TRIMELLITATE|TRIDECYL TRIMELLITATE
C3486860|T121|1309695|RXNORM|GELSEMIUM SEMPERVIRENS ROOT EXTRACT|GELSEMIUM SEMPERVIRENS ROOT EXTRACT
C3488689|T121|1309694|RXNORM|SELENICEREUS GRANDIFLORUS STEM EXTRACT|SELENICEREUS GRANDIFLORUS STEM EXTRACT
C3489213|T121|1309697|RXNORM|HAMAMELIS VIRGINIANA ROOT BARK-STEM BARK EXTRACT|HAMAMELIS VIRGINIANA ROOT BARK-STEM BARK EXTRACT
C2718418|T129|857953|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-BRISBANE-60-2008 STRAIN|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-BRISBANE-60-2008 STRAIN
C2604029|T197|1309691|RXNORM|ARSENIC TRIIODIDE|ARSENIC TRIIODIDE
C2947577|T121|1309690|RXNORM|DIOSCOREA VILLOSA TUBER EXTRACT|DIOSCOREA VILLOSA TUBER EXTRACT
C3484471|T121|1309692|RXNORM|STRYCHNOS IGNATII SEED EXTRACT|STRYCHNOS IGNATII SEED EXTRACT
C2702015|T121|853142|RXNORM|TOURMALINE|TOURMALINE
C1874173|T121|705058|RXNORM|ALUMINUM SULFATE / CALCIUM ACETATE|ALUMINUM SULFATE / CALCIUM ACETATE
C3464493|T121|1344626|RXNORM|LUPINUS ALBUS SEED EXTRACT|LUPINUS ALBUS SEED EXTRACT
C3667050|T121|1438291|RXNORM|ROSA CANINA LEAF EXTRACT|ROSA CANINA LEAF EXTRACT
C0102139|T126|46049|RXNORM|ALGLUCERASE|ALGLUCERASE
C0085857|T121|42547|RXNORM|AUROTHIOMALATE|AUROTHIOMALATE
C3864828|T129|1596934|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 58 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 58 VACCINE
C3496144|T109|1370373|RXNORM|BRINE SHRIMP EXTRACT|BRINE SHRIMP EXTRACT
C0102118|T121|46041|RXNORM|ALENDRONATE|ALENDRONATE
C0041056|T121|10834|RXNORM|TRIMIPRAMINE|TRIMIPRAMINE
C0041044|T121|10831|RXNORM|SULFAMETHOXAZOLE / TRIMETHOPRIM|SULFAMETHOXAZOLE / TRIMETHOPRIM
C0000589|T121|1426888|RXNORM|5-METHOXYTRYPTAMINE|5-METHOXYTRYPTAMINE
C3693115|T121|1482550|RXNORM|WHEAT SPROUT EXTRACT|WHEAT SPROUT EXTRACT
C0050133|T195|1482551|RXNORM|9,10-ANTHRAQUINONE|9,10-ANTHRAQUINONE
C0021218|T120|1426889|RXNORM|INDIGO|INDIGO
C1874360|T121|689509|RXNORM|ASPIRIN / CAFFEINE / CHLORPHENIRAMINE|ASPIRIN / CAFFEINE / CHLORPHENIRAMINE
C2929707|T121|1008808|RXNORM|CASCARA SAGRADA / SENNOSIDES, USP|CASCARA SAGRADA / SENNOSIDES, USP
C2929708|T121|1008809|RXNORM|BUTABARBITAL / MEPROBAMATE|BUTABARBITAL / MEPROBAMATE
C2929705|T121|1008806|RXNORM|LODGEPOLE PINE POLLEN EXTRACT / YELLOW PINE POLLEN EXTRACT|LODGEPOLE PINE POLLEN EXTRACT / YELLOW PINE POLLEN EXTRACT
C2929706|T121|1008807|RXNORM|EMODEPSIDE / PRAZIQUANTEL|EMODEPSIDE / PRAZIQUANTEL
C2929703|T121|1008804|RXNORM|GREEN ASH POLLEN EXTRACT / WHITE ASH POLLEN EXTRACT|GREEN ASH POLLEN EXTRACT / WHITE ASH POLLEN EXTRACT
C2929701|T121|1008802|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / DIPHENHYDRAMINE / PHENYLEPHRINE|ACETAMINOPHEN / DEXTROMETHORPHAN / DIPHENHYDRAMINE / PHENYLEPHRINE
C2929699|T121|1008800|RXNORM|CALCIUM CARBONATE / CALCIUM GLUCONATE / CHOLECALCIFEROL|CALCIUM CARBONATE / CALCIUM GLUCONATE / CHOLECALCIFEROL
C2929700|T121|1008801|RXNORM|AMLODIPINE / HYDROCHLOROTHIAZIDE / OLMESARTAN|AMLODIPINE / HYDROCHLOROTHIAZIDE / OLMESARTAN
C1874665|T121|691028|RXNORM|CALCIUM GLUCONATE / NIACINAMIDE / PHENOBARBITAL|CALCIUM GLUCONATE / NIACINAMIDE / PHENOBARBITAL
C0055716|T121|21095|RXNORM|CICLOXILIC ACID|CICLOXILIC ACID
C3475017|T121|1302463|RXNORM|INULIN / LACTOBACILLUS RHAMNOSUS GG|INULIN / LACTOBACILLUS RHAMNOSUS GG
C0055711|T121|21090|RXNORM|CICLOPIROX|CICLOPIROX
C2722053|T129|892338|RXNORM|KHUSKIA ORYZAE ALLERGENIC EXTRACT|KHUSKIA ORYZAE ALLERGENIC EXTRACT
C0030092|T195|7821|RXNORM|OXYTETRACYCLINE|OXYTETRACYCLINE
C0055720|T121|21099|RXNORM|CIFENLINE|CIBENZOLINE
C0030095|T125|7824|RXNORM|OXYTOCIN|OXYTOCIN
C2193907|T121|816562|RXNORM|BUMETANIDE / POTASSIUM CHLORIDE|BUMETANIDE / POTASSIUM CHLORIDE
C1874909|T121|690102|RXNORM|CODEINE / TERPIN HYDRATE|CODEINE / TERPIN HYDRATE
C2365098|T121|1426448|RXNORM|CERAMIDE 2|CERAMIDE 2
C0173083|T121|61805|RXNORM|NITISINONE|NITISINONE
C0771343|T121|236106|RXNORM|POISON IVY EXTRACT|POISON IVY EXTRACT
C0771726|T121|236452|RXNORM|DI-ISOPROPYLAMMONIUM|DI-ISOPROPYLAMMONIUM
C3256681|T121|1312593|RXNORM|GARDEN CRESS SPROUT EXTRACT|GARDEN CRESS SPROUT EXTRACT
C2684346|T129|852819|RXNORM|PERENNIAL RYE GRASS POLLEN EXTRACT|LOLIUM PERENNE POLLEN EXTRACT
C3853726|T109|1552036|RXNORM|ARISTOLOCHIA CLEMATITIS WHOLE EXTRACT|ARISTOLOCHIA CLEMATITIS WHOLE EXTRACT
C0770991|T121|235812|RXNORM|HEXYLNICOTINATE|HEXYLNICOTINATE
C1451502|T121|1244607|RXNORM|TAFLUPROST|TAFLUPROST
C0034235|T121|8984|RXNORM|PYRANTEL|PYRANTEL
C0034239|T121|8987|RXNORM|PYRAZINAMIDE|PYRAZINAMIDE
C1171081|T168|1370769|RXNORM|RASPBERRY EXTRACT|RASPBERRY EXTRACT
C3256876|T109|1427080|RXNORM|WHEAT MIDDLINGS EXTRACT|WHEAT MIDDLINGS EXTRACT
C0058645|T122|1427083|RXNORM|LAURTRIMONIUM|LAURTRIMONIUM
C1533312|T121|1370766|RXNORM|BARLEY EXTRACT|BARLEY EXTRACT
C1122970|T121|1370761|RXNORM|QUINCE EXTRACT|QUINCE EXTRACT
C3486607|T121|1348451|RXNORM|ASCLEPIAS CURASSAVICA EXTRACT|ASCLEPIAS CURASSAVICA EXTRACT
C0302923|T197|1427087|RXNORM|PHOSPHONIC ACID|PHOSPHOROUS ACID
C3179443|T121|1427086|RXNORM|AVOTERMIN|AVOTERMIN
C2928490|T121|1007570|RXNORM|DIMETHICONE / MICONAZOLE / ZINC OXIDE|DIMETHICONE / MICONAZOLE / ZINC OXIDE
C3692236|T121|1441543|RXNORM|ALNUS GLUTINOSA BARK EXTRACT|BLACK ALDER BARK EXTRACT
C3692237|T121|1441544|RXNORM|ALSTONIA CONSTRICTA BARK EXTRACT|ALSTONIA CONSTRICTA BARK EXTRACT
C2827079|T121|1441545|RXNORM|AMMONIUM VALERATE|AMMONIUM VALERATE
C0003036|T131|1441546|RXNORM|ANILINE|ANILINE
C3535909|T121|1369685|RXNORM|LINOLEAMIDOPROPYL PG-DIMONIUM|LINOLEAMIDOPROPYL PG-DIMONIUM
C1302004|T121|392466|RXNORM|CHLORTHALIDONE / TRIAMTERENE|CHLORTHALIDONE / TRIAMTERENE
C0008290|T121|2406|RXNORM|CHLORPROTHIXENE|CHLORPROTHIXENE
C0018033|T121|4980|RXNORM|AUROTHIOGLUCOSE|AUROTHIOGLUCOSE
C0008287|T121|2404|RXNORM|CHLORPROPAMIDE|CHLORPROPAMIDE
C3486759|T121|1353887|RXNORM|DIEFFENBACHIA SEGUINE EXTRACT|DIEFFENBACHIA SEGUINE EXTRACT
C0008286|T121|2403|RXNORM|CHLORPROMAZINE|CHLORPROMAZINE
C0008281|T121|2400|RXNORM|CHLORPHENIRAMINE|CHLORPHENIRAMINE
C0008281|T121|2400|RXNORM|CHLORPHENIRAMINE|CHLORPHENIRAMINE
C0018062|T125|4986|RXNORM|CHORIONIC GONADOTROPIN|CHORIONIC GONADOTROPIN
C3486761|T121|1353888|RXNORM|LOBARIA PULMONARIA EXTRACT|LOBARIA PULMONARIA EXTRACT
C0525079|T121|134547|RXNORM|BENDAMUSTINE|BENDAMUSTINE
C0008293|T195|2408|RXNORM|CHLORTETRACYCLINE|CHLORTETRACYCLINE
C0008293|T195|2408|RXNORM|CHLORTETRACYCLINE|CHLORTETRACYCLINE
C0008294|T121|2409|RXNORM|CHLORTHALIDONE|CHLORTHALIDONE
C1444903|T121|465680|RXNORM|FLUOCINOLONE / HYDROQUINONE / TRETINOIN|FLUOCINOLONE / HYDROQUINONE / TRETINOIN
C2701136|T129|851890|RXNORM|TREE OF HEAVEN POLLEN EXTRACT|AILANTHUS ALTISSIMA POLLEN EXTRACT
C2927584|T129|1006371|RXNORM|MANGO BLOSSOM POLLEN EXTRACT|MANGIFERA INDICA POLLEN EXTRACT
C1961041|T121|820887|RXNORM|CHLORHEXIDINE / NEOMYCIN|CHLORHEXIDINE / NEOMYCIN
C3854066|T121|1547608|RXNORM|EUPHORBIA AMYGDALOIDES EXTRACT|EUPHORBIA AMYGDALOIDES EXTRACT
C0006796|T121|1951|RXNORM|CAMBENDAZOLE|CAMBENDAZOLE
C1693169|T121|631158|RXNORM|ACETAMINOPHEN / GUAIFENESIN / PHENYLEPHRINE|ACETAMINOPHEN / GUAIFENESIN / PHENYLEPHRINE
C1874171|T121|690771|RXNORM|ALUMINUM HYDROXIDE / MAGNESIUM TRISILICATE / PHENYLBUTAZONE|ALUMINUM HYDROXIDE / MAGNESIUM TRISILICATE / PHENYLBUTAZONE
C0006809|T121|1952|RXNORM|CAMPHOR|CAMPHOR
C0011689|T121|3248|RXNORM|DESLANOSIDE|DESLANOSIDE
C3486562|T129|1367198|RXNORM|REPTOCOCCUS VIRIDANS GROUP IMMUNOSERUM RABBIT|REPTOCOCCUS VIRIDANS GROUP IMMUNOSERUM RABBIT
C3486567|T129|1367199|RXNORM|MALARIAL PLASMODIUM GROUP IMMUNOSERUM RABBIT|MALARIAL PLASMODIUM GROUP IMMUNOSERUM RABBIT
C3486560|T129|1367196|RXNORM|MYCOBACTERIUM MICROTI IMMUNOSERUM RABBIT|MYCOBACTERIUM MICROTI IMMUNOSERUM RABBIT
C3486561|T129|1367197|RXNORM|STREPTOCOCCUS PYOGENES IMMUNOSERUM RABBIT|STREPTOCOCCUS PYOGENES IMMUNOSERUM RABBIT
C3486558|T129|1367194|RXNORM|STREPTOCOCCUS PNEUMONIAE IMMUNOSERUM RABBIT|STREPTOCOCCUS PNEUMONIAE IMMUNOSERUM RABBIT
C3486559|T129|1367195|RXNORM|MYCOBACTERIUM BOVIS IMMUNOSERUM RABBIT|MYCOBACTERIUM BOVIS IMMUNOSERUM RABBIT
C0011685|T121|3247|RXNORM|DESIPRAMINE|DESIPRAMINE
C3486556|T129|1367193|RXNORM|LACTOCOCCUS LACTIS IMMUNOSERUM RABBIT|LACTOCOCCUS LACTIS IMMUNOSERUM RABBIT
C3475126|T121|1367190|RXNORM|PENTYLAMINE|PENTYLAMINE
C0043801|T131|1367191|RXNORM|1,2-DIBROMO-3-CHLOROPROPANE|1,2-DIBROMO-3-CHLOROPROPANE
C0303762|T121|90737|RXNORM|PETROLEUM DISTILLATE|PETROLEUM DISTILLATE
C3528936|T121|1363758|RXNORM|EUCALYPTOL / MENTHOL / SODIUM FLUORIDE / THYMOL|EUCALYPTOL / MENTHOL / SODIUM FLUORIDE / THYMOL
C3528063|T121|1361667|RXNORM|HEPATITIS A VACCINE (INACTIVATED) STRAIN HM175 / TYPHOID VI POLYSACCHARIDE VACCINE, S TYPHI TY2 STRAIN|HEPATITIS A VACCINE (INACTIVATED) STRAIN HM175 / TYPHOID VI POLYSACCHARIDE VACCINE, S TYPHI TY2 STRAIN
C0083031|T129|1311380|RXNORM|INTERLEUKIN-11|INTERLEUKIN-11
C0040383|T109|1311381|RXNORM|TOLUENE|TOLUENE
C0037248|T123|1311386|RXNORM|SKATOLE|SKATOLE
C0008240|T123|1311387|RXNORM|CHLOROGENIC ACID|CHLOROGENIC ACID
C0039462|T196|1311384|RXNORM|TELLURIUM|TELLURIUM
C3486841|T121|1311385|RXNORM|SINUSITISINUM|SINUSITISINUM
C0019846|T196|1311388|RXNORM|HOLMIUM|HOLMIUM
C0016979|T130|1311389|RXNORM|GALLIC ACID|GALLIC ACID
C0020281|T197|5499|RXNORM|HYDROGEN PEROXIDE|HYDROGEN PEROXIDE
C0020281|T197|5499|RXNORM|HYDROGEN PEROXIDE|HYDROGEN PEROXIDE
C0020273|T121|5495|RXNORM|HYDROFLUMETHIAZIDE|HYDROFLUMETHIAZIDE
C2828287|T109|1426442|RXNORM|FERRIC AMMONIUM FERROCYANIDE|FERRIC AMMONIUM FERROCYANIDE
C3531468|T129|1366997|RXNORM|INFLUENZA A VIRUS ANTIGEN, PANAMA 2007-99 (H3N2)|INFLUENZA A VIRUS ANTIGEN, PANAMA 2007-99 (H3N2)
C0020268|T125|5492|RXNORM|HYDROCORTISONE|HYDROCORTISONE
C0020268|T125|5492|RXNORM|HYDROCORTISONE|HYDROCORTISONE
C0020268|T125|5492|RXNORM|HYDROCORTISONE|HYDROCORTISONE
C0020268|T125|5492|RXNORM|HYDROCORTISONE|HYDROCORTISONE
C0020268|T125|5492|RXNORM|HYDROCORTISONE|HYDROCORTISONE
C0020268|T125|5492|RXNORM|HYDROCORTISONE|HYDROCORTISONE
C0020268|T125|5492|RXNORM|HYDROCORTISONE|HYDROCORTISONE
C3854019|T195|1596450|RXNORM|GENTAMICIN|GENTAMICIN
C0007080|T121|2068|RXNORM|CARBUTAMIDE|CARBUTAMIDE
C3256513|T121|1307839|RXNORM|CLEMATIS VITALBA LEAF EXTRACT|CLEMATIS VITALBA LEAF EXTRACT
C3256592|T121|1307838|RXNORM|AGAVE AMERICANA LEAF EXTRACT|CENTURY PLANT LEAF EXTRACT
C3488538|T121|1353222|RXNORM|AMMI VISNAGA FRUIT EXTRACT|VISNAGA DAUCOIDES FRUIT EXTRACT
C3486824|T121|1353221|RXNORM|EPIFAGUS VIRGINIANA EXTRACT|EPIFAGUS VIRGINIANA EXTRACT
C3486711|T121|1353220|RXNORM|ATROPA BELLADONNA ROOT EXTRACT|ATROPA BELLADONNA ROOT EXTRACT
C0054803|T122|1307833|RXNORM|CARNAUBA WAX|CARNAUBA WAX
C3256014|T121|1307832|RXNORM|ALPINIA OFFICINARUM LEAF EXTRACT|ALPINIA OFFICINARUM LEAF EXTRACT
C3256138|T121|1307831|RXNORM|COIX LACRYMA-JOBI SEED EXTRACT|COIX LACRYMA-JOBI SEED EXTRACT
C0108407|T122|1307830|RXNORM|CARBOMER-934|CARBOMER HOMOPOLYMER TYPE B (ALLYL SUCROSE CROSSLINKED)
C3256915|T121|1307837|RXNORM|GUAZUMA ULMIFOLIA LEAF EXTRACT|GUAZUMA ULMIFOLIA LEAF EXTRACT
C0086079|T121|42618|RXNORM|CRYPTENAMINE|CRYPTENAMINE
C3255901|T109|1307835|RXNORM|MYRTLE LEAF OIL|MYRTLE LEAF OIL
C3464953|T121|1307834|RXNORM|MORINGA OLEIFERA LEAF EXTRACT|MORINGA OLEIFERA LEAF EXTRACT
C3256215|T109|1363578|RXNORM|CYCLOMETHICONE 4|CYCLOMETHICONE 4
C3256223|T109|1363579|RXNORM|DIMETHICONOL (41 MPA.S)|DIMETHICONOL (41 MPA.S)
C0982105|T130|1310563|RXNORM|D & C RED # 30 ALUMINUM LAKE|D & C RED # 30 ALUMINUM LAKE
C0040263|T121|10612|RXNORM|TINIDAZOLE|TINIDAZOLE
C0059756|T121|1310565|RXNORM|ETHYL CELLULOSE|ETHYL CELLULOSE
C1509304|T120|1310564|RXNORM|D&C RED NO. 7|D&C RED NO. 7
C0851342|T197|1310566|RXNORM|MAGNESIUM SILICATE|MAGNESIUM SILICATE
C1699573|T121|1363570|RXNORM|PEG-30 DIPOLYHYDROXYSTEARATE|PEG-30-DIPOLYHYDROXYSTEARATE
C0001963|T131|1310568|RXNORM|METHANOL|METHANOL
C1952498|T121|1363572|RXNORM|METHYL GLUCETH-20|METHYL GLUCETH-20
C2608247|T121|1363573|RXNORM|LAURETH-10|LAURETH-10
C2342361|T109|1363574|RXNORM|METHYL STEARATE|METHYL STEARATE
C2607173|T109|1363575|RXNORM|HEXYLDECANOL|HEXYLDECANOL
C2603860|T131|1363576|RXNORM|COCAMIDOPROPYLAMINE OXIDE|COCAMIDOPROPYLAMINE OXIDE
C3256203|T109|1363577|RXNORM|LAURETH-12|LAURETH-12
C0040557|T204|1432991|RXNORM|TOXOPLASMA GONDII|TOXOPLASMA GONDII
C2730119|T129|892360|RXNORM|GRAIN MOTH EXTRACT|SITOTROGA CEREALELLA EXTRACT
C0301311|T121|89729|RXNORM|ACRISORCIN|ACRISORCIN
C2608095|T121|1314409|RXNORM|DL-LACTIC ACID|DL-LACTIC ACID
C3486757|T121|1311167|RXNORM|PORK KIDNEY PREPARATION|PORK KIDNEY PREPARATION
C1871062|T122|1311164|RXNORM|CARBOPOL 981|CARBOMER HOMOPOLYMER TYPE A (ALLYL PENTAERYTHRITOL CROSSLINKED)
C1589331|T129|544488|RXNORM|BOTULISM IMMUNE GLOBULIN IV HUMAN|BOTULISM IMMUNE GLOBULIN IV HUMAN
C0301304|T121|89722|RXNORM|PHENYLMERCURIC NITRATE|PHENYLMERCURIC NITRATE
C0301303|T121|89721|RXNORM|NITROMERSOL|NITROMERSOL
C0086073|T121|42612|RXNORM|CROMOLYN|CROMOLYN
C0086073|T121|42612|RXNORM|CROMOLYN|CROMOLYN
C0086073|T121|42612|RXNORM|CROMOLYN|CROMOLYN
C0086073|T121|42612|RXNORM|CROMOLYN|CROMOLYN
C0042629|T007|1432992|RXNORM|VIBRIO CHOLERAE|VIBRIO CHOLERAE
C0014824|T130|4061|RXNORM|ERYTHROSINE|ERYTHROSINE
C3832914|T121|1539899|RXNORM|CHLOROXYLENOL / SALICYLIC ACID / SODIUM THIOSULFATE|CHLOROXYLENOL / SALICYLIC ACID / SODIUM THIOSULFATE
C0053114|T121|18889|RXNORM|BENOXINATE|OXYBUPROCAINE
C0007068|T121|2062|RXNORM|CARBOXYMETHYLCELLULOSE|CARBOXYMETHYLCELLULOSE
C2182926|T121|817999|RXNORM|CHLORDIAZEPOXIDE / DESIPRAMINE|CHLORDIAZEPOXIDE / DESIPRAMINE
C1703661|T121|618060|RXNORM|THIOCTATE|THIOCTATE
C0082491|T121|41078|RXNORM|ETHOXAZENE|ETHOXAZENE
C0002144|T121|519|RXNORM|ALLOPURINOL|ALLOPURINOL
C0065865|T121|29439|RXNORM|MEDRYSONE|MEDRYSONE
C0065858|T121|29434|RXNORM|MEDIFOXAMINE|MEDIFOXAMINE
C0002119|T131|513|RXNORM|ALLETHRIN|ALLETHRIN
C0939813|T121|285163|RXNORM|BITTERSWEET EXTRACT|BITTERSWEET EXTRACT
C0002132|T121|516|RXNORM|ALLOBARBITAL|ALLOBARBITAL
C0004320|T121|1227|RXNORM|AURANOFIN|AURANOFIN
C0301464|T121|89858|RXNORM|ALUMINUM CARBONATE|ALUMINUM CARBONATE
C1328051|T121|729750|RXNORM|COENZYME Q10 / VITAMIN E|COENZYME Q10 / VITAMIN E
C0002403|T121|620|RXNORM|AMANTADINE|AMANTADINE
C0004259|T121|1223|RXNORM|ATROPINE|ATROPINE
C0004259|T121|1223|RXNORM|ATROPINE|ATROPINE
C0004259|T121|1223|RXNORM|ATROPINE|ATROPINE
C0002435|T195|626|RXNORM|AMDINOCILLIN|AMDINOCILLIN
C0002421|T121|625|RXNORM|AMBROXOL|AMBROXOL
C2928944|T121|1008033|RXNORM|HYDROCORTISONE / KETOCONAZOLE|HYDROCORTISONE / KETOCONAZOLE
C3856017|T121|1549461|RXNORM|ESTRADIOL / TRENBOLONE|ESTRADIOL / TRENBOLONE
C0058716|T121|23651|RXNORM|DOXACURIUM|DOXACURIUM
C0024337|T123|6536|RXNORM|LYSINE|LYSINE
C2928122|T121|1007200|RXNORM|HYDROXYZINE / MECLIZINE|HYDROXYZINE / MECLIZINE
C2928125|T121|1007203|RXNORM|DEQUALINIUM / HEXETIDINE|DEQUALINIUM / HEXETIDINE
C2928124|T121|1007202|RXNORM|CETRIMIDE / DIPHENHYDRAMINE / MOROXYDINE|CETRIMIDE / DIPHENHYDRAMINE / MOROXYDINE
C2928127|T121|1007205|RXNORM|CALCIUM GLUCONATE / CALCIUM SACCHARATE|CALCIUM GLUCONATE / CALCIUM SACCHARATE
C2928126|T121|1007204|RXNORM|CODEINE / PROPYPHENAZONE|CODEINE / PROPYPHENAZONE
C2928129|T121|1007207|RXNORM|SODIUM BICARBONATE / SODIUM PHOSPHATE, MONOBASIC|SODIUM BICARBONATE / SODIUM PHOSPHATE, MONOBASIC
C0024328|T125|6531|RXNORM|LYPRESSIN|LYPRESSIN
C2928131|T121|1007209|RXNORM|GOLDENSEAL EXTRACT / PAPAIN|GOLDENSEAL EXTRACT / PAPAIN
C2928130|T121|1007208|RXNORM|DEXPANTHENOL / ZINC OXIDE|DEXPANTHENOL / ZINC OXIDE
C2918527|T129|995747|RXNORM|BALD CYPRESS POLLEN EXTRACT|TAXODIUM DISTICHUM POLLEN EXTRACT
C0063750|T121|27723|RXNORM|IODINATED GLYCEROL|IODINATED GLYCEROL
C0063750|T121|27723|RXNORM|IODINATED GLYCEROL|IODINATED GLYCEROL
C0033508|T121|8792|RXNORM|PROPYLHEXEDRINE|PROPYLHEXEDRINE
C2918524|T129|995743|RXNORM|CANADA GOLDENROD POLLEN EXTRACT|SOLIDAGO CANADENSIS POLLEN EXTRACT
C0602896|T121|156762|RXNORM|BUTETHAMATE CITRATE|BUTETHAMATE CITRATE
C2928195|T121|1007273|RXNORM|ACTIVATED CHARCOAL / CALCIUM CARBONATE|ACTIVATED CHARCOAL / CALCIUM CARBONATE
C3531389|T109|1366710|RXNORM|SILK, ENZYME HYDROLYZED (1000 MW)|SILK, ENZYME HYDROLYZED (1000 MW)
C0033511|T121|8794|RXNORM|PROPYLTHIOURACIL|PROPYLTHIOURACIL
C0677942|T196|196342|RXNORM|SAMARIUM SM153|SAMARIUM SM153
C3700899|T121|1486392|RXNORM|MORINDA OFFICINALIS WHOLE EXTRACT|MORINDA OFFICINALIS WHOLE EXTRACT
C0033513|T123|8795|RXNORM|PROSCILLARIDIN|PROSCILLARIDIN
C0052593|T121|18475|RXNORM|ATIPAMEZOLE|ATIPAMEZOLE
C0771858|T129|798444|RXNORM|HAEMOPHILUS INFLUENZAE B (ROSS STRAIN) CAPSULAR POLYSACCHARIDE MENINGOCOCCAL PROTEIN CONJUGATE VACCINE|HAEMOPHILUS INFLUENZAE B (ROSS STRAIN) CAPSULAR POLYSACCHARIDE MENINGOCOCCAL PROTEIN CONJUGATE VACCINE
C2018744|T121|814684|RXNORM|BUTHIAZIDE / SPIRONOLACTONE|BUTHIAZIDE / SPIRONOLACTONE
C0939815|T121|285165|RXNORM|STRYCHNOS IGNATII PREPARATION|STRYCHNOS IGNATII PREPARATION
C1874696|T121|691188|RXNORM|CAMPHOR / MENTHOL / METHYL SALICYLATE|CAMPHOR / MENTHOL / METHYL SALICYLATE
C2183762|T121|814681|RXNORM|CHLORMEZANONE / DIPYRONE|CHLORMEZANONE / DIPYRONE
C0248572|T121|73455|RXNORM|DORAMECTIN|DORAMECTIN
C2756324|T129|967960|RXNORM|PENICILLIUM ITALICUM EXTRACT|PENICILLIUM ITALICUM EXTRACT
C0873140|T121|259473|RXNORM|AMERICAN GINSENG ROOT|AMERICAN GINSENG ROOT
C0873139|T121|259472|RXNORM|SIBERIAN GINSENG ROOT EXTRACT|SIBERIAN GINSENG ROOT EXTRACT
C0873138|T121|259471|RXNORM|KOREAN GINSENG ROOT EXTRACT|KOREAN GINSENG ROOT EXTRACT
C0873137|T121|259470|RXNORM|KOREAN GINSENG PREPARATION|KOREAN GINSENG PREPARATION
C3538611|T121|1373153|RXNORM|HYDROXYETHYL BEHENAMIDOPROPYL DIMONIUM CHLORIDE|HYDROXYETHYL BEHENAMIDOPROPYL DIMONIUM CHLORIDE
C3538610|T121|1373152|RXNORM|ETHYLBISIMINOMETHYLGUAIACOL MANGANESE CHLORIDE|ETHYLBISIMINOMETHYLGUAIACOL MANGANESE CHLORIDE
C0018302|T130|1373150|RXNORM|GUAIAC|GUAIAC
C3538615|T121|1373157|RXNORM|POLYGONATUM BIFLORUM ROOT ETXRACT|POLYGONATUM BIFLORUM ROOT ETXRACT
C3538614|T121|1373156|RXNORM|NELUMBO NUCIFERA WHOLE EXTRACT|NELUMBO NUCIFERA WHOLE EXTRACT
C3538613|T121|1373155|RXNORM|NELUMBO NUCIFERA ROOT EXTRACT|NELUMBO NUCIFERA ROOT EXTRACT
C3538612|T121|1373154|RXNORM|LAURYL PEG-9 POLYDIMETHYLSILOXYETHYL DIMETHICONE|LAURYL PEG-9 POLYDIMETHYLSILOXYETHYL DIMETHICONE
C0072127|T121|34604|RXNORM|PROLINTANE|PROLINTANE
C3538617|T121|1373159|RXNORM|PRUNUS ARMENIACA WHOLE EXTRACT|PRUNUS ARMENIACA WHOLE EXTRACT
C3538616|T121|1373158|RXNORM|POLYGONATUM ODORATUM WHOLE EXTRACT|POLYGONATUM ODORATUM WHOLE EXTRACT
C0031676|T123|8246|RXNORM|PHOSPHOLIPIDS|PHOSPHOLIPIDS
C2709744|T129|854940|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 15B VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 15B VACCINE
C0163557|T121|1047072|RXNORM|MOXIDECTIN|MOXIDECTIN
C3500118|T121|1313834|RXNORM|ASCORBIC ACID / BACILLUS COAGULANS / CRANBERRY PREPARATION|ASCORBIC ACID / BACILLUS COAGULANS / CRANBERRY PREPARATION
C3531377|T109|1366670|RXNORM|ISOPROPYLBENZYL SALICYLATE|ISOPROPYLBENZYL SALICYLATE
C3531378|T109|1366671|RXNORM|ISOCETYL STEAROYL STEARATE|ISOCETYL STEAROYL STEARATE
C0073603|T121|35805|RXNORM|ROYAL JELLY|ROYAL JELLY
C1529800|T121|498193|RXNORM|BOSENTAN MONOHYDRATE|BOSENTAN MONOHYDRATE
C2961881|T121|1053719|RXNORM|CHLOPHEDIANOL / GUAIFENESIN|CHLOPHEDIANOL / GUAIFENESIN
C1119918|T121|325526|RXNORM|GINSENG PREPARATION|GINSENG PREPARATION
C0297985|T197|88188|RXNORM|ZINC BROMIDE|ZINC BROMIDE
C0057143|T121|22298|RXNORM|DAPIPRAZOLE|DAPIPRAZOLE
C0057144|T195|22299|RXNORM|DAPTOMYCIN|DAPTOMYCIN
C0057135|T121|22293|RXNORM|DANTHRON|DANTRON
C0015109|T121|4166|RXNORM|ETHYLMORPHINE|ETHYLMORPHINE
C0719248|T121|215976|RXNORM|MAGNESIUM, CHELATED|MAGNESIUM, CHELATED
C0015099|T125|4162|RXNORM|ETHYLESTRENOL|ETHYLESTRENOL
C0937630|T121|283570|RXNORM|HAWTHORN BERRY|HAWTHORN BERRY
C0015116|T121|4169|RXNORM|ETILEFRINE|ETILEFRINE
C2980906|T121|1094155|RXNORM|REDROOT PIGWEED POLLEN EXTRACT / SPINY PIGWEED POLLEN EXTRACT|REDROOT PIGWEED POLLEN EXTRACT / SPINY PIGWEED POLLEN EXTRACT
C0068660|T130|1364276|RXNORM|NEW COCCINE|NEW COCCINE
C3486524|T121|1314323|RXNORM|BUDDLEJA DAVIDII WHOLE EXTRACT|BUDDLEJA DAVIDII WHOLE EXTRACT
C2981043|T121|1094405|RXNORM|CHLOPHEDIANOL / TRIPROLIDINE|CHLOPHEDIANOL / TRIPROLIDINE
C2073834|T121|1303250|RXNORM|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE
C3484865|T121|1314322|RXNORM|KJELLMANIELLA GYRATA PREPARATION|KJELLMANIELLA GYRATA PREPARATION
C3256331|T109|1307558|RXNORM|AMINOPROPYL ASCORBYL PHOSPHATE|AMINOPROPYL ASCORBYL PHOSPHATE
C3464667|T121|1307559|RXNORM|MATRICARIA CHAMOMILLA WHOLE EXTRACT|MATRICARIA CHAMOMILLA WHOLE EXTRACT
C2347826|T121|1339883|RXNORM|COLLINSONIA EXTRACT|COLLINSONIA EXTRACT
C2347823|T121|1314321|RXNORM|CAULOPHYLLUM ROBUSTUM ROOT EXTRACT|CAULOPHYLLUM ROBUSTUM ROOT EXTRACT
C3256631|T121|1307550|RXNORM|POLYGONATUM ODORATUM ROOT EXTRACT|POLYGONATUM ODORATUM ROOT EXTRACT
C0050461|T121|16738|RXNORM|RACECADOTRIL|RACECADOTRIL
C3256615|T121|1307553|RXNORM|FILIPENDULA ULMARIA FLOWER EXTRACT|FILIPENDULA ULMARIA FLOWER EXTRACT
C3474824|T121|1307554|RXNORM|ARTEMISIA CAPILLARIS FLOWER EXTRACT|ARTEMISIA CAPILLARIS FLOWER EXTRACT
C3256479|T121|1307555|RXNORM|1-(4-(4-CHLOROPHENYL)-3-PHENYL-2-BUTENYL)-PYRROLIDINE 1,5-NAPHTHALENEDISULFONATE|PYRROBUTAMINE NAPHTHALENE DISULFONATE
C3256149|T109|1307556|RXNORM|CORNUS OFFICINALIS FRUIT EXTRACT|CORNUS OFFICINALIS FRUIT EXTRACT
C3486307|T121|1307557|RXNORM|MENTHA X ROTUNDIFOLIA LEAF EXTRACT|MENTHA X ROTUNDIFOLIA LEAF EXTRACT
C0875914|T121|261408|RXNORM|CARBETAPENTANE / CHLORPHENIRAMINE / PHENYLEPHRINE|CARBETAPENTANE / CHLORPHENIRAMINE / PHENYLEPHRINE
C2701447|T129|852252|RXNORM|DOMESTIC GOAT SKIN EXTRACT|CAPRA HIRCUS SKIN EXTRACT
C0772505|T121|237162|RXNORM|DEXKETOPROFEN|DEXKETOPROFEN
C3643369|T109|1421434|RXNORM|COCO DIISOPROPANOLAMIDE|COCO DIISOPROPANOLAMIDE
C0071538|T121|1364277|RXNORM|POLYDATIN|POLYDATIN
C2701451|T129|852256|RXNORM|DOMESTIC COW SKIN EXTRACT|DOMESTIC COW SKIN EXTRACT
C2701753|T129|852709|RXNORM|SHORTLEAF PINE POLLEN EXTRACT|PINUS ECHINATA POLLEN EXTRACT
C1112096|T121|324044|RXNORM|DESOGESTREL / ETHINYL ESTRADIOL|DESOGESTREL / ETHINYL ESTRADIOL
C2701749|T129|852704|RXNORM|DATE PALM POLLEN EXTRACT|PHOENIX DACTYLIFERA POLLEN EXTRACT
C1110663|T121|324040|RXNORM|PODOPHYLLUM PREPARATION|PODOPHYLLUM PREPARATION
C2727011|T129|1014711|RXNORM|SUGARCANE ALLERGENIC EXTRACT|SUGARCANE ALLERGENIC EXTRACT
C1112082|T121||RXNORM|HYDROCHLOROTHIAZIDE / SPIRONOLACTONE
C0007738|T195|2239|RXNORM|CEPHRADINE|CEPHRADINE
C0007737|T195|2238|RXNORM|CEPHAPIRIN|CEPHAPIRIN
C3500688|T121|1315107|RXNORM|ARGERATINA AROMATICA ROOT EXTRACT|ARGERATINA AROMATICA ROOT EXTRACT
C2016765|T121|817886|RXNORM|SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC|SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC
C2016765|T121|817886|RXNORM|SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC|SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC
C2016765|T121|817886|RXNORM|SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC|SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC
C3555512|T109|1375415|RXNORM|CASTOR FIBER SCENT GLAND SECRETION|CASTOR FIBER SCENT GLAND SECRETION
C0007550|T195|2182|RXNORM|CEFMETAZOLE|CEFMETAZOLE
C0007716|T195|2231|RXNORM|CEPHALEXIN|CEPHALEXIN
C0007727|T195|2233|RXNORM|CEPHALORIDINE|CEPHALORIDINE
C3530454|T121|1364410|RXNORM|IOXAPINE|IOXAPINE
C0007735|T195|2236|RXNORM|CEPHALOTHIN|CEPHALOTHIN
C0021971|T130|5936|RXNORM|IODIPAMIDE|ADIPIODONE
C3256623|T109|1426452|RXNORM|ISOSTEARAMIDOPROPYL MORPHOLINE LACTATE|ISOSTEARAMIDOPROPYL MORPHOLINE LACTATE
C0021968|T196|5933|RXNORM|IODINE|MOLECULAR IODINE
C3256135|T109|1426455|RXNORM|COCO-GLYCERIDES|COCO-GLYCERIDES
C0020835|T129|1426454|RXNORM|IMMUNOGLOBULIN A|IMMUNOGLOBULIN A
C0012522|T121|3498|RXNORM|DIPHENHYDRAMINE|DIPHENHYDRAMINE
C0012522|T121|3498|RXNORM|DIPHENHYDRAMINE|DIPHENHYDRAMINE
C0600319|T130|155060|RXNORM|PYROGLUTAMATE|PIDOLATE
C3255766|T109|1426456|RXNORM|ETHYLENE-VINYL ACETATE COPOLYMER (28% VINYL ACETATE)|ETHYLENE-VINYL ACETATE COPOLYMER (28% VINYL ACETATE)
C0125901|T123|595958|RXNORM|LINOLENATE|LINOLENATE
C0016745|T121|4570|RXNORM|FRUCTOSE|FRUCTOSE
C2726996|T129|973447|RXNORM|CRICKET ALLERGENIC EXTRACT|ACHETA DOMESTICUS ALLERGENIC EXTRACT
C1654825|T121|605496|RXNORM|CARBETAPENTANE / GUAIFENESIN|CARBETAPENTANE / GUAIFENESIN
C0007557|T195|2189|RXNORM|CEFOXITIN|CEFOXITIN
C3696422|T121|1483211|RXNORM|CHLOROXYLENOL / ETHANOL|CHLOROXYLENOL / ETHANOL
C2183745|T121|817082|RXNORM|DIPHENYLPYRALINE / PHENYLEPHRINE|DIPHENYLPYRALINE / PHENYLEPHRINE
C0304095|T168|90926|RXNORM|ANISE OIL|ANISE OIL
C2756506|T129|968437|RXNORM|WHEAT LOOSE SMUT EXTRACT|WHEAT LOOSE SMUT ALLERGENIC EXTRACT
C2698280|T121|1291301|RXNORM|AVANAFIL|AVANAFIL
C0031398|T121|8126|RXNORM|PHENYLETHYL ALCOHOL|PHENYLETHYL ALCOHOL
C3255921|T109|1306207|RXNORM|CITRUS MAXIMA FRUIT RIND EXTRACT|CITRUS MAXIMA FRUIT RIND EXTRACT
C3255917|T109|1306206|RXNORM|CITRUS AURANTIUM FRUIT RIND EXTRACT|CITRUS AURANTIUM FRUIT RIND EXTRACT
C3255914|T109|1306205|RXNORM|CITRUS AURANTIUM FLOWER EXTRACT|CITRUS AURANTIUM FLOWER EXTRACT
C3255911|T109|1306204|RXNORM|CHRYSANTHEMUM X MORIFOLIUM FLOWER EXTRACT|CHRYSANTHEMUM X MORIFOLIUM FLOWER EXTRACT
C3255910|T109|1306203|RXNORM|CHYSANTHELLUM INDICUM TOP EXTRACT|CHYSANTHELLUM INDICUM TOP EXTRACT
C3255908|T109|1306201|RXNORM|CHOLETH-20|CHOLETH-20
C3255907|T109|1306200|RXNORM|CHOLESTERYL STEARATE|CHOLESTERYL STEARATE
C0055146|T121|20609|RXNORM|CETIEDIL|CETIEDIL
C3255924|T109|1306209|RXNORM|CITRUS MAXIMA SEED EXTRACT|CITRUS MAXIMA SEED EXTRACT
C3255923|T109|1306208|RXNORM|CITRUS MAXIMA LEAF EXTRACT|CITRUS MAXIMA LEAF EXTRACT
C3663106|T168|1432476|RXNORM|OPUNTIA FICUS-INDICA FRUIT JUICE EXTRACT|OPUNTIA FICUS-INDICA FRUIT JUICE
C3663107|T121|1432477|RXNORM|TILIA CORDATA, WHOLE EXTRACT|TILIA CORDATA, WHOLE EXTRACT
C3663104|T121|1432474|RXNORM|WHOLE MELIA AZEDERACH EXTRACT|WHOLE MELIA AZEDERACH EXTRACT
C3663105|T121|1432475|RXNORM|WHOLE ERIODICTYON CALIFORNICUM EXTRACT|WHOLE ERIODICTYON CALIFORNICUM EXTRACT
C3663103|T121|1432472|RXNORM|CODONOPSIS LANCEOLATA ROOT EXTRACT|CODONOPSIS LANCEOLATA ROOT EXTRACT
C3542474|T121|1432473|RXNORM|LARICIFOMES OFFICINALIS WHOLE EXTRACT|LARICIFOMES OFFICINALIS WHOLE EXTRACT
C3831878|T109|1538052|RXNORM|LAURETH-30|LAURETH-30
C3484463|T121|1310013|RXNORM|DALBERGIA PINNATA ROOT EXTRACT|DALBERGIA PINNATA ROOT EXTRACT
C3663108|T121|1432478|RXNORM|PUNICA GRANATUM WHOLE EXTRACT|PUNICA GRANATUM WHOLE EXTRACT
C3663109|T121|1432479|RXNORM|DIETHOXYETHYL SUCCINATE|DIETHOXYETHYL SUCCINATE
C1302013|T121|392475|RXNORM|ATENOLOL / NIFEDIPINE|ATENOLOL / NIFEDIPINE
C1302012|T121|392474|RXNORM|NYSTATIN / TOLNAFTATE|NYSTATIN / TOLNAFTATE
C1302016|T121|392477|RXNORM|ASCORBIC ACID / CLIOQUINOL|ASCORBIC ACID / CLIOQUINOL
C2983812|T121|1300786|RXNORM|MIRABEGRON|MIRABEGRON
C1302010|T121|392472|RXNORM|EPHEDRINE / THEOPHYLLINE|EPHEDRINE / THEOPHYLLINE
C3643372|T109|1421431|RXNORM|TRIDECYL SALICYLATE|TRIDECYL SALICYLATE
C0965129|T121|301542|RXNORM|ROSUVASTATIN|ROSUVASTATIN
C3696417|T121|1483778|RXNORM|ACETAMIDOPROPYL TRIMONIUM|ACETAMIDOPROPYL TRIMONIUM
C0102834|T121|46239|RXNORM|ALUMINUM ACETOTARTRATE|ALUMINIUM ACETOTARTRATE
C1707080|T121|657797|RXNORM|TEMSIROLIMUS|TEMSIROLIMUS
C3695946|T121|1484857|RXNORM|POLYACRYLIC ACID (8000 MW)|POLYACRYLIC ACID (8000 MW)
C3496185|T121|1368650|RXNORM|CINNAMATE|CINNAMATE
C1682316|T121|619676|RXNORM|ACETAMINOPHEN / METHIONINE|ACETAMINOPHEN / METHIONINE
C1874873|T121|689865|RXNORM|CLIOQUINOL / COAL TAR / HYDROCORTISONE|CLIOQUINOL / COAL TAR / HYDROCORTISONE
C1874874|T121|689867|RXNORM|CLIOQUINOL / HYDROCORTISONE / PRAMOXINE|CLIOQUINOL / HYDROCORTISONE / PRAMOXINE
C1099675|T121|322165|RXNORM|THIOSALICYLIC ACID|THIOSALICYLIC ACID
C1268876|T121|386938|RXNORM|FOLLITROPIN ALFA|FOLLITROPIN ALFA
C3256449|T109|1311640|RXNORM|TALLOW ACID, BEEF|TALLOW ACID, BEEF
C3664998|T121|1435105|RXNORM|TRAMETES VERSICOLOR WHOLE EXTRACT|TRAMETES VERSICOLOR WHOLE EXTRACT
C3465009|T109|1427142|RXNORM|BENZYLIDENE DIMETHOXYDIMETHYLINDANONE|BENZYLIDENE DIMETHOXYDIMETHYLINDANONE
C3256756|T109|1427143|RXNORM|CAPROOYL TETRAPEPTIDE-3|CAPROOYL TETRAPEPTIDE-3
C1509676|T121|1427148|RXNORM|PPG-3 MYRISTYL ETHER|PPG-3 MYRISTYL ETHER
C0054690|T121|1427149|RXNORM|CARBOCYSTEINE-LYSINE|CARBOCYSTEINE-LYSINE
C0771967|T121|236665|RXNORM|BLACK COHOSH EXTRACT|BLACK COHOSH EXTRACT
C0771966|T121|236664|RXNORM|CHASTE TREE PREPARATION|CHASTE TREE PREPARATION
C0771960|T129|236660|RXNORM|BOTULISM ANTITOXIN E|BOTULISM ANTITOXIN E
C0070709|T121|33408|RXNORM|PHENYLTOLOXAMINE|PHENYLTOLOXAMINE
C2702371|T129|892628|RXNORM|PORK ALLERGENIC EXTRACT|PORK ALLERGENIC EXTRACT
C0052506|T121|18405|RXNORM|ASIATICOSIDE|ASIATICOSIDE
C2928842|T121|1007928|RXNORM|PANTOTHENATE / VITAMIN B6|PANTOTHENATE / VITAMIN B6
C2928843|T121|1007929|RXNORM|HYDROCHLOROTHIAZIDE / TRIAMTERENE / VERAPAMIL|HYDROCHLOROTHIAZIDE / TRIAMTERENE / VERAPAMIL
C0070557|T195|33277|RXNORM|PHENETHICILLIN|PHENETICILLIN
C2928834|T121|1007920|RXNORM|DANTHRON / PANTOTHENIC ACID|DANTHRON / PANTOTHENIC ACID
C2928835|T121|1007921|RXNORM|GUAIAZULENE / PENTOSAN POLYSULFATE|GUAIAZULENE / PENTOSAN POLYSULFATE
C2928836|T121|1007922|RXNORM|GREATER CELANDINE / SILYMARIN|GREATER CELANDINE / SILYMARIN
C2928837|T121|1007923|RXNORM|DEANOL / HEPTAMINOL|DEANOL / HEPTAMINOL
C2928838|T121|1007924|RXNORM|CAPSAICIN / METHYLNICOTINATE|CAPSAICIN / METHYLNICOTINATE
C2928839|T121|1007925|RXNORM|LEVOCARNITINE / PICOLINIC ACID|LEVOCARNITINE / PICOLINIC ACID
C2928840|T121|1007926|RXNORM|ASCORBIC ACID / CALCIUM LACTATE|ASCORBIC ACID / CALCIUM LACTATE
C2928841|T121|1007927|RXNORM|BENZYLPARABEN / PROPYLPARABEN|BENZYLPARABEN / PROPYLPARABEN
C0026400|T121|7023|RXNORM|MOLSIDOMINE|MOLSIDOMINE
C1453538|T109|1489548|RXNORM|MONOMENTHYL GLUTARATE|MONOMENTHYL GLUTARATE
C0076286|T121|37935|RXNORM|TETRAHYDROZOLINE|TETRYZOLINE
C0076286|T121|37935|RXNORM|TETRAHYDROZOLINE|TETRYZOLINE
C0034261|T121|9000|RXNORM|PYRIDOSTIGMINE|PYRIDOSTIGMINE
C3818822|T121|1489544|RXNORM|CHINESE RHUBARB ROOT EXRACT|CHINESE RHUBARB ROOT EXRACT
C3256618|T109|1312592|RXNORM|FOSVESET|FOSVESET
C3818820|T121|1489546|RXNORM|COMMIPHORA MYRRHA TOP EXTRACT|COMMIPHORA MYRRHA TOP EXTRACT
C3818819|T121|1489547|RXNORM|GERANIUM WILFORDII TOP EXTRACT|GERANIUM WILFORDII TOP EXTRACT
C0034282|T121|9009|RXNORM|PYRILAMINE|PYRILAMINE
C0038774|T196|10223|RXNORM|SULFUR|SULFUR
C0038774|T196|10223|RXNORM|SULFUR|SULFUR
C3500490|T121|1314653|RXNORM|COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / SODIUM ASCORBATE / THIAMINE / VITAMIN B 12 / ZINC SULFATE|COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / SODIUM ASCORBATE / THIAMINE / VITAMIN B 12 / ZINC SULFATE
C0060549|T130|25161|RXNORM|FLUOREXON STAIN|FLUOREXON STAIN
C1144109|T109|1314657|RXNORM|ETHYLHEXYL TRIAZONE|OCTYL TRIAZONE
C1113645|T129|1314656|RXNORM|RADISH EXTRACT|RADISH EXTRACT
C0065525|T197|1362814|RXNORM|MAGNESIUM NITRATE|MAGNESIUM NITRATE
C2983889|T121|1329960|RXNORM|HUMAN PLACENTA HYDROLYSATE|HUMAN PLACENTA HYDROLYSATE
C3528650|T121|1362811|RXNORM|BETAINE / BROMELAINS / PANCREATIN / PAPAIN / PEPSIN A|BETAINE / BROMELAINS / PANCREATIN / PAPAIN / PEPSIN A
C3256493|T121|1362813|RXNORM|ACACIA DECURRENS EXTRACT|ACACIA DECURRENS EXTRACT
C0039329|T120|1305578|RXNORM|TARTRAZINE|TARTRAZINE
C0064970|T130|1305579|RXNORM|LIGHT GREEN SF YELLOWISH|LIGHT GREEN SF YELLOWISH
C0060120|T130|1305574|RXNORM|FD&C YELLOW NO. 6|FD&C YELLOW NO. 6
C0066052|T130|1305576|RXNORM|METANIL YELLOW|METANIL YELLOW
C0443770|T121|991260|RXNORM|HEPTANOIC ACID|HEPTANOIC ACID
C0028735|T121|7595|RXNORM|NYLIDRIN|NYLIDRIN
C0046079|T121|1433902|RXNORM|2-DIETHYLAMINOETHANOL|2-DIETHYLAMINOETHANOL
C0030031|T195|7798|RXNORM|OXOLINIC ACID|OXOLINIC ACID
C2740621|T129|899420|RXNORM|GINGER ALLERGENIC EXTRACT|ZINGIBER OFFICINALE ALLERGENIC EXTRACT
C3857943|T121|1552576|RXNORM|TRIETHANOLAMINE 2-CYCLOHEXYL-4,6-DINITROPHENOLATE|TRIETHANOLAMINE 2-CYCLOHEXYL-4,6-DINITROPHENOLATE
C3857944|T121|1552574|RXNORM|AINSLIAEA FRAGRANS TOP EXTRACT|AINSLIAEA FRAGRANS TOP EXTRACT
C0054274|T121|1552575|RXNORM|DIETHYLENE GLYCOL MONOBUTYL ETHER|DIETHYLENE GLYCOL MONOBUTYL ETHER
C0000959|T121|155|RXNORM|ACEPROMAZINE|ACEPROMAZINE
C2740627|T129|899428|RXNORM|HADDOCK ALLERGENIC EXTRACT|MELANOGRAMMUS AEGLEFINUS ALLERGENIC EXTRACT
C0049690|T127|1088438|RXNORM|6-O-PALMITOYLASCORBIC ACID|6-O-PALMITOYLASCORBIC ACID
C3257508|T109|1426782|RXNORM|ULVA COMPRESSA EXTRACT|ULVA COMPRESSA EXTRACT
C0051809|T121|596724|RXNORM|ANAGRELIDE|ANAGRELIDE
C3859497|T121|1593134|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP B RECOMBINANT LP2086 A05 PROTEIN VARIANT ANTIGEN / NEISSERIA MENINGITIDIS SEROGROUP B RECOMBINANT LP2086 B01 PROTEIN VARIANT ANTIGEN|NEISSERIA MENINGITIDIS SEROGROUP B RECOMBINANT LP2086 A05 PROTEIN VARIANT ANTIGEN / NEISSERIA MENINGITIDIS SEROGROUP B RECOMBINANT LP2086 B01 PROTEIN VARIANT ANTIGEN
C1961852|T121|236901|RXNORM|SOMATORELIN|SOMATORELIN
C0939844|T121|285193|RXNORM|RED CLOVER PREPARATION|RED CLOVER PREPARATION
C2929182|T121|1008275|RXNORM|DIPROPIZINE / GUAIFENESIN|DIPROPIZINE / GUAIFENESIN
C2929181|T121|1008274|RXNORM|ISOPROPYL ALCOHOL / POVIDONE-IODINE|ISOPROPYL ALCOHOL / POVIDONE-IODINE
C2929184|T121|1008277|RXNORM|BENZALKONIUM / PRAMOXINE|BENZALKONIUM / PRAMOXINE
C2929178|T121|1008271|RXNORM|DIBUNATE / GUAIACOLSULFONATE|DIBUNATE / GUAIACOLSULFONATE
C2929180|T121|1008273|RXNORM|ALANINE / ARGININE / ASPARTATE / CYSTEINE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM METABISULFITE / TAURINE / THREONINE / TRYPTOPHAN / TYRO|ALANINE / ARGININE / ASPARTATE / CYSTEINE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM METABISULFITE / TAURINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929179|T121|1008272|RXNORM|DIPHTHERIA TOXOID VACCINE, INACTIVATED / HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE|DIPHTHERIA TOXOID VACCINE, INACTIVATED / HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE
C2929186|T121|1008279|RXNORM|COBAMAMIDE / VITAMIN B 12|COBAMAMIDE / VITAMIN B 12
C2929185|T121|1008278|RXNORM|CAMPHOR / MENTHOL / PHENOL / SALICYLIC ACID|CAMPHOR / MENTHOL / PHENOL / SALICYLIC ACID
C3463997|T121|1311598|RXNORM|HAMAMELIS VIRGINIANA TOP WATER EXTRACT|HAMAMELIS VIRGINIANA TOP WATER EXTRACT
C1096768|T121|319866|RXNORM|MEGLUMINE ANTIMONIATE|MEGLUMINE ANTIMONIATE
C1096766|T121|319864|RXNORM|CISATRACURIUM|CISATRACURIUM
C1096793|T121|319868|RXNORM|1,4-BENZOQUINONE|1,4-BENZOQUINONE
C0982278|T121|1367118|RXNORM|METHYL GLUCETH-10|METHYL GLUCETH-10
C3255965|T109|1312710|RXNORM|PEG-12 DILAURATE|PEG-12 DILAURATE
C3256070|T109|1312711|RXNORM|PEG-3 ALPHA-LINOLENAMIDE|PEG-3 ALPHA-LINOLENAMIDE
C3256073|T121|1312712|RXNORM|PEG-4 STEARATE|PEG-4 STEARATE
C3256172|T121|1312714|RXNORM|METHYL DIISOPROPYL PROPIONAMIDE|METHYL DIISOPROPYL PROPIONAMIDE
C0304346|T121|91099|RXNORM|THIOSALICYLATE|THIOSALICYLATE
C3256176|T109|1312716|RXNORM|PENTAERYTHRITYL DISTEARATE|PENTAERYTHRITYL DISTEARATE
C3256248|T121|1312717|RXNORM|PHELLINUS LINTEUS MYCELIUM EXTRACT|PHELLINUS LINTEUS MYCELIUM EXTRACT
C3256254|T121|1312719|RXNORM|4-((4,6-BIS(OCTYLTHIO)-1,3,5-TRIAZIN-2-YL)AMINO)-2,6-BIS(1,1-DIMETHYLETHYL)-PHENOL|4-((4,6-BIS(OCTYLTHIO)-1,3,5-TRIAZIN-2-YL)AMINO)-2,6-BIS(1,1-DIMETHYLETHYL)-PHENOL
C2186922|T121|812468|RXNORM|DIHYDRALAZINE / HYDROCHLOROTHIAZIDE / RESERPINE|DIHYDRALAZINE / HYDROCHLOROTHIAZIDE / RESERPINE
C0981931|T129|314415|RXNORM|MUCOR PLUMBEUS ALLERGENIC EXTRACT|MUCOR PLUMBEUS ALLERGENIC EXTRACT
C0068333|T121|31447|RXNORM|NABILONE|NABILONE
C0014912|T125|4083|RXNORM|ESTRADIOL|ESTRADIOL
C0014912|T125|4083|RXNORM|ESTRADIOL|ESTRADIOL
C0014921|T121|4089|RXNORM|ESTRAMUSTINE|ESTRAMUSTINE
C0257343|T121|77492|RXNORM|TAMSULOSIN|TAMSULOSIN
C2080580|T121|817377|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / GUAIFENESIN / PHENYLPROPANOLAMINE|ACETAMINOPHEN / CHLORPHENIRAMINE / GUAIFENESIN / PHENYLPROPANOLAMINE
C0247025|T121|73137|RXNORM|TIROFIBAN|TIROFIBAN
C0068334|T121|31448|RXNORM|NABUMETONE|NABUMETONE
C3864826|T130|1597292|RXNORM|SOLVENT RED 4|SOLVENT RED 4
C3853718|T121|1597293|RXNORM|ORIGANUM VULGARE SUBSP. HIRTUM WHOLE EXTRACT|ORIGANUM VULGARE SUBSP. HIRTUM WHOLE EXTRACT
C1509273|T121|1311621|RXNORM|CETEARETH-15|CETEARETH-15
C1533387|T109|1311620|RXNORM|CETEARETH-12|CETEARETH-12
C2929225|T121|1008318|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-CALIFORNIA-07-2009 X-179A (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-VICTORIA-210-2009 X-187 (H3N2) (A-PERTH-16-2009) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-CALIFORNIA-07-2009 X-179A (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-VICTORIA-210-2009 X-187 (H3N2) (A-PERTH-16-2009) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN
C2929226|T121|1008319|RXNORM|CAFFEINE / CODEINE / PHENIRAMINE / PHENYLEPHRINE / SALICYLIC ACID|CAFFEINE / CODEINE / PHENIRAMINE / PHENYLEPHRINE / SALICYLIC ACID
C0043155|T121|11327|RXNORM|WHITE WAX|WHITE WAX
C3497971|T121|1311627|RXNORM|LIMONIUM VULGARE FLOWERING TOP EXTRACT|LIMONIUM VULGARE FLOWERING TOP EXTRACT
C0028013|T196|1311629|RXNORM|NICKEL|NICKEL
C2929220|T121|1008313|RXNORM|PLANTAGO SEED / SENNOSIDES, USP|PLANTAGO SEED / SENNOSIDES, USP
C2929218|T121|1008311|RXNORM|PRUNE PREPARATION / SENNOSIDES, USP|PRUNE PREPARATION / SENNOSIDES, USP
C2929223|T121|1008316|RXNORM|HYDROGEN PEROXIDE / LACTATE|HYDROGEN PEROXIDE / LACTATE
C2929224|T121|1008317|RXNORM|CAMPHOR / MENTHOL / METHYL SALICYLATE / THYMOL|CAMPHOR / MENTHOL / METHYL SALICYLATE / THYMOL
C2929221|T121|1008314|RXNORM|CALCIUM POLYCARBOPHIL / SENNOSIDES, USP|CALCIUM POLYCARBOPHIL / SENNOSIDES, USP
C2929222|T121|1008315|RXNORM|CODEINE / GUAIFENESIN / PROMETHAZINE|CODEINE / GUAIFENESIN / PROMETHAZINE
C3710016|T109|1488820|RXNORM|PINUS KORAIENSIS SEED OIL|PINUS KORAIENSIS SEED OIL
C3710017|T109|1488821|RXNORM|PINUS MUGO SUBSP. MUGO BARK EXTRACT|PINUS MUGO SUBSP. MUGO BARK EXTRACT
C2348650|T109|1488822|RXNORM|TANSY OIL|TANSY OIL
C3710018|T109|1488823|RXNORM|SUS SCROFA VENTRICLE PREPARATION|PORCINE VENTRICLE PREPARATION
C3255677|T109|1307037|RXNORM|HEXANEDIOL|HEXANEDIOL
C3257443|T121|1307035|RXNORM|LENS CULINARIS FRUIT EXTRACT|LENS CULINARIS FRUIT EXTRACT
C3474583|T121|1307039|RXNORM|METHYLBENZYL METHYLBENZIMIDAZOLE PIPERIDINYLMETHANONE|METHYLBENZYL METHYLBENZIMIDAZOLE PIPERIDINYLMETHANONE
C3256614|T109|1307038|RXNORM|DECYL OLEATE|DECYL OLEATE
C1141002|T121|340262|RXNORM|PRUNE PREPARATION|PRUNE PREPARATION
C0717824|T121|214618|RXNORM|HYDROCHLOROTHIAZIDE / LISINOPRIL|HYDROCHLOROTHIAZIDE / LISINOPRIL
C0717825|T121|214619|RXNORM|HYDROCHLOROTHIAZIDE / LOSARTAN|HYDROCHLOROTHIAZIDE / LOSARTAN
C3695944|T109|1484859|RXNORM|SOY ACID|SOY ACID
C0717820|T121|214614|RXNORM|HOMATROPINE / HYDROCODONE|HOMATROPINE / HYDROCODONE
C0717821|T121|214615|RXNORM|HYDRALAZINE / HYDROCHLOROTHIAZIDE|HYDRALAZINE / HYDROCHLOROTHIAZIDE
C0717822|T121|214616|RXNORM|HYDRALAZINE / HYDROCHLOROTHIAZIDE / RESERPINE|HYDRALAZINE / HYDROCHLOROTHIAZIDE / RESERPINE
C0717823|T121|214617|RXNORM|HYDROCHLOROTHIAZIDE / IRBESARTAN|HYDROCHLOROTHIAZIDE / IRBESARTAN
C3474471|T121|1313199|RXNORM|PENTAERYTHRITYL TETRACAPRYLATE-TETRACAPRATE|PENTAERYTHRITYL TETRACAPRYLATE-TETRACAPRATE
C2726151|T129|999463|RXNORM|GEOTRICHUM CANDIDUM ALLERGENIC EXTRACT|GEOTRICHUM CANDIDUM ALLERGENIC EXTRACT
C3504692|T109|1356479|RXNORM|ABIES BALSAMEA LEAF OIL|ABIES BALSAMEA LEAF OIL
C3695945|T109|1484858|RXNORM|ISOPROPYL LINOLEATE|ISOPROPYL LINOLEATE
C0058344|T121|23350|RXNORM|DIOXYBENZONE|DIOXYBENZONE
C0106291|T121|47111|RXNORM|BIFEMELANE|BIFEMELANE
C3152335|T121|1094890|RXNORM|LIDOCAINE / MENTHOL / METHYL SALICYLATE|LIDOCAINE / MENTHOL / METHYL SALICYLATE
C0251516|T130|74671|RXNORM|CORTICORELIN OVINE|CORTICORELIN OVINE
C3473991|T121|1307789|RXNORM|SAURURUS CHINENSIS FLOWER EXTRACT|SAURURUS CHINENSIS FLOWER EXTRACT
C3256813|T109|1307788|RXNORM|VETIVER OIL|VETIVER OIL
C3256896|T121|1307784|RXNORM|CARTHAMUS TINCTORIUS (SAFFLOWER) OLEOSOMES EXTRACT|CARTHAMUS TINCTORIUS (SAFFLOWER) OLEOSOMES EXTRACT
C3488909|T121|1307787|RXNORM|BANCHA TEA, LEAF, TWIG PREPARATION|BANCHA TEA, LEAF, TWIG PREPARATION
C3256404|T121|1307781|RXNORM|1,2-DIARACHIDOYL-SN-GLYCERO-3-PHOSPHOCHOLINE|1,2-DIARACHIDOYL-SN-GLYCERO-3-PHOSPHOCHOLINE
C3256280|T121|1307780|RXNORM|C20-22 ALCOHOLS|C20-22 ALCOHOLS
C3256901|T109|1307783|RXNORM|CETEARETH-33|CETEARETH-33
C3486532|T121|1307782|RXNORM|SYRINGA VULGARIS FLOWER EXTRACT|SYRINGA VULGARIS FLOWER EXTRACT
C2701271|T129|852062|RXNORM|TOBACCO LEAF EXTRACT|TOBACCO LEAF EXTRACT
C3503436|T121|1358491|RXNORM|SUGARCANE EXTRACT|SUGARCANE EXTRACT
C1655908|T121|1358490|RXNORM|POLYETHYLENE GLYCOL 4500|POLYETHYLENE GLYCOL 4500
C0982258|T121|314711|RXNORM|LICORICE EXTRACT|LICORICE EXTRACT
C2347236|T121|819929|RXNORM|BUTAFOSFAN|BUTAFOSFAN
C0054152|T121|19791|RXNORM|BROVANEXINE|BROVANEXINE
C0054151|T121|19790|RXNORM|BROTIZOLAM|BROTIZOLAM
C0536495|T195|139462|RXNORM|MOXIFLOXACIN|MOXIFLOXACIN
C0536495|T195|139462|RXNORM|MOXIFLOXACIN|MOXIFLOXACIN
C3855821|T109|1549143|RXNORM|POLIXETONIUM|POLIXETONIUM
C2037257|T121|814917|RXNORM|DIAZEPAM / SULPIRIDE|DIAZEPAM / SULPIRIDE
C1433763|T129|458451|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18
C0024778|T121|6646|RXNORM|MAPROTILINE|MAPROTILINE
C0085154|T121|42319|RXNORM|NIZATIDINE|NIZATIDINE
C3811626|T116|1536616|RXNORM|FLATHEAD SOLE PREPARATION|FLATHEAD SOLE PREPARATION
C1874370|T121|689522|RXNORM|ASPIRIN / CARISOPRODOL / CODEINE|ASPIRIN / CARISOPRODOL / CODEINE
C1807658|T121|689524|RXNORM|ASPIRIN / CITRIC ACID / SODIUM BICARBONATE|ASPIRIN / CITRIC ACID / SODIUM BICARBONATE
C2939977|T129|1014385|RXNORM|BERMUDA GRASS SMUT EXTRACT|USTILAGO CYNODONTIS EXTRACT
C3669022|T121|1482536|RXNORM|ERYNGIUM MARITIMUM EXTRACT|ERYNGIUM MARITIMUM EXTRACT
C0041014|T125|10814|RXNORM|TRIIODOTHYRONINE|LIOTHYRONINE
C3555525|T121|1374400|RXNORM|HIMATANTHUS LANCIFOLIUS BARK EXTRACT|HIMATANTHUS LANCIFOLIUS BARK EXTRACT
C1874374|T121|689529|RXNORM|ASPIRIN / ETHOHEPTAZINE / MEPROBAMATE|ASPIRIN / ETHOHEPTAZINE / MEPROBAMATE
C0041023|T121|10819|RXNORM|TRIMEBUTINE|TRIMEBUTINE
C3555522|T121|1374403|RXNORM|MINQUARTIA GUIANENSIS BARK EXTRACT|MINQUARTIA GUIANENSIS BARK EXTRACT
C3555521|T121|1374404|RXNORM|PHYLLANTHUS NIRURI WHOLE EXTRACT|PHYLLANTHUS NIRURI WHOLE EXTRACT
C3555520|T121|1374405|RXNORM|PIPER ADUNCUM LEAF EXTRACT|PIPER ADUNCUM LEAF EXTRACT
C3555519|T109|1374406|RXNORM|SORBITAN DIOLEATE|SORBITAN DIOLEATE
C2929766|T121|1008868|RXNORM|CODEINE / GUAIACOLSULFONATE|CODEINE / GUAIACOLSULFONATE
C2929767|T121|1008869|RXNORM|BILBERRY EXTRACT / CALCIUM CITRATE / MAGNESIUM GLYCINATE / POTASSIUM CITRATE / VITAMIN E|BILBERRY EXTRACT / CALCIUM CITRATE / MAGNESIUM GLYCINATE / POTASSIUM CITRATE / VITAMIN E
C0030053|T121|7805|RXNORM|OXYFEDRINE|OXYFEDRINE
C0030049|T121|7804|RXNORM|OXYCODONE|OXYCODONE
C0030054|T196|7806|RXNORM|OXYGEN|OXYGEN
C2929758|T121|1008860|RXNORM|AMPHETAMINE / PHENOBARBITAL|AMPHETAMINE / PHENOBARBITAL
C2929759|T121|1008861|RXNORM|ASCORBIC ACID / INOSITOL|ASCORBIC ACID / INOSITOL
C2929760|T121|1008862|RXNORM|ASCORBIC ACID / RUTIN / VINCAMINE|ASCORBIC ACID / RUTIN / VINCAMINE
C2929761|T121|1008863|RXNORM|DEXPANTHENOL / PREDNISOLONE / SALICYLIC ACID|DEXPANTHENOL / PREDNISOLONE / SALICYLIC ACID
C2929762|T121|1008864|RXNORM|LAURETH-9 / PREDNISOLONE / PROMETHAZINE|POLIDOCANOL / PREDNISOLONE / PROMETHAZINE
C2929764|T121|1008866|RXNORM|ACETAMINOPHEN / PAMABROM / VITAMIN B6|ACETAMINOPHEN / PAMABROM / VITAMIN B6
C2929765|T121|1008867|RXNORM|LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS BIFIDUS|LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS BIFIDUS
C0054235|T121|19861|RXNORM|BUTAMBEN|BUTAMBEN
C0054234|T121|19860|RXNORM|BUTALBITAL|BUTALBITAL
C0054236|T121|19862|RXNORM|BUTAMIRATE|BUTAMIRATE
C3848527|T196|1546429|RXNORM|GADOLINIUM CATION (3+)|GADOLINIUM CATION (3+)
C0023726|T195|6398|RXNORM|LINCOMYCIN|LINCOMYCIN
C0540209|T121|1426467|RXNORM|3-IODO-2-PROPYNYLBUTYLCARBAMATE|IODOPROPYNYL BUTYLCARBAMATE
C0023665|T121|6390|RXNORM|LIDOFLAZINE|LIDOFLAZINE
C0008273|T121|2396|RXNORM|CHLOROTHIAZIDE|CHLOROTHIAZIDE
C0008275|T125|2397|RXNORM|CHLOROTRIANISENE|CHLOROTRIANISENE
C3818763|T196|1492441|RXNORM|IODINE I-120|IODINE I-120
C0008269|T121|2393|RXNORM|CHLOROQUINE|CHLOROQUINE
C0521934|T121|1492443|RXNORM|TRICAINE METHANESULFONATE|TRICAINE METHANESULFONATE
C3818762|T109|1492442|RXNORM|ORCHIS MASCULA TUBER EXTRACT|ORCHIS MASCULA TUBER EXTRACT
C0008280|T121|2399|RXNORM|CHLORPHENESIN|CHLORPHENESIN
C0888714|T130|1426460|RXNORM|D&C BLUE NO. 4|D&C BLUE NO. 4
C1703862|T121|618442|RXNORM|TIAPROFENATE|TIAPROFENATE
C0772093|T004|236782|RXNORM|SACCHAROMYCES BOULARDII|SACCHAROMYCES BOULARDII
C0060236|T197|1428835|RXNORM|FERRIC HYDROXIDE|FERRIC HYDROXIDE
C1445663|T121|466431|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C3255877|T109|1313979|RXNORM|STEARYL GLUCOSIDE|STEARYL GLUCOSIDE
C0772095|T121|236784|RXNORM|DETAJMIUM BITARTRATE|DETAJMIUM BITARTRATE
C0055856|T195|21212|RXNORM|CLARITHROMYCIN|CLARITHROMYCIN
C0055856|T195|21212|RXNORM|CLARITHROMYCIN|CLARITHROMYCIN
C3651776|T121|1428837|RXNORM|MELIA AZEDARACH BARK EXTRACT|MELIA AZEDARACH BARK EXTRACT
C3473111|T121|1298165|RXNORM|CALCIUM CARBONATE / VITAMIN B 12|CALCIUM CARBONATE / VITAMIN B 12
C3714499|T121|1546422|RXNORM|EPICRIPTINE|EPICRIPTINE
C2935436|T129|1371041|RXNORM|TRASTUZUMAB-DM1 CONJUGATE|ADO-TRASTUZUMAB EMTANSINE
C2106235|T121|815532|RXNORM|COAL TAR / HYDROCORTISONE|COAL TAR / HYDROCORTISONE
C3848529|T197|1546424|RXNORM|NITRITE ION|NITRITE ION
C0007537|T195|2176|RXNORM|CEFACLOR|CEFACLOR
C0007538|T195|2177|RXNORM|CEFADROXIL|CEFADROXIL
C0017992|T121|4967|RXNORM|GLYOXAL|GLYOXAL
C0007541|T195|2178|RXNORM|CEFAMANDOLE|CEFAMANDOLE
C3651778|T109|1428832|RXNORM|2-(L-MENTHOXY)ETHANOL|2-(L-MENTHOXY)ETHANOL
C2726136|T129|1006310|RXNORM|ASPERGILLUS REPENS ALLERGENIC EXTRACT|ASPERGILLUS REPENS ALLERGENIC EXTRACT
C1165729|T129|851878|RXNORM|ORCHARD GRASS POLLEN EXTRACT|ORCHARD GRASS POLLEN EXTRACT
C2701126|T129|851874|RXNORM|HARD MAPLE POLLEN EXTRACT|ACER SACCHARUM POLLEN EXTRACT
C0981893|T129|851870|RXNORM|REDTOP GRASS POLLEN EXTRACT|AGROSTIS GIGANTEA POLLEN EXTRACT
C1875415|T121|690713|RXNORM|KAOLIN / PAREGORIC / PECTIN|KAOLIN / PAREGORIC / PECTIN
C0011777|T121|3264|RXNORM|DEXAMETHASONE|DEXAMETHASONE
C0011777|T121|3264|RXNORM|DEXAMETHASONE|DEXAMETHASONE
C0011777|T121|3264|RXNORM|DEXAMETHASONE|DEXAMETHASONE
C0011777|T121|3264|RXNORM|DEXAMETHASONE|DEXAMETHASONE
C0011777|T121|3264|RXNORM|DEXAMETHASONE|DEXAMETHASONE
C0011777|T121|3264|RXNORM|DEXAMETHASONE|DEXAMETHASONE
C0011777|T121|3264|RXNORM|DEXAMETHASONE|DEXAMETHASONE
C0011785|T121|3267|RXNORM|DEXETIMIDE|DEXETIMIDE
C0011786|T121|3268|RXNORM|DEXFENFLURAMINE|DEXFENFLURAMINE
C0005098|T121|1424|RXNORM|BENZTROPINE|BENZTROPINE
C1874721|T121|692971|RXNORM|CARBON MONOXIDE / HELIUM / NITROGEN / OXYGEN|CARBON MONOXIDE / HELIUM / NITROGEN / OXYGEN
C1874720|T121|692970|RXNORM|CARBON DIOXIDE / OXYGEN|CARBON DIOXIDE / OXYGEN
C1875125|T121|692979|RXNORM|ESTRADIOL / HYDROXYPROGESTERONE|17-ALPHA-HYDROXYPROGESTERONE / ESTRADIOL
C3833114|T197|1540524|RXNORM|ALUMINUM HYDRIDE|ALUMINUM HYDRIDE
C2954513|T121|1048074|RXNORM|CHLOPHEDIANOL / GUAIFENESIN / PHENYLEPHRINE|CHLOPHEDIANOL / GUAIFENESIN / PHENYLEPHRINE
C0303739|T196|90719|RXNORM|169 YTTERBIUM|169 YTTERBIUM
C3486634|T121|1310367|RXNORM|EUPHORBIA RESINIFERA RESIN EXTRACT|EUPHORBIA RESINIFERA RESIN
C0369246|T195|113608|RXNORM|FUSIDATE|FUSIDATE
C2929392|T121|1008488|RXNORM|ADENINE / GLUCOSE|ADENINE / GLUCOSE
C2929393|T121|1008489|RXNORM|GUAIACOLSULFONIC ACID / PHENYLEPHRINE|GUAIACOLSULFONIC ACID / PHENYLEPHRINE
C3488573|T121|1311368|RXNORM|PLANTAGO MAJOR EXTRACT|PLANTAGO MAJOR EXTRACT
C2929386|T121|1008482|RXNORM|DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE / PYRILAMINE|DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE / PYRILAMINE
C2929387|T121|1008483|RXNORM|ALUMINUM POTASSIUM SULFATE / PHENOL|ALUMINUM POTASSIUM SULFATE / PHENOL
C3497930|T121|1311366|RXNORM|SUS SCROFA ACHILLES TENDON PREPARATION|PORCINE ACHILLES TENDON PREPARATION
C2929385|T121|1008481|RXNORM|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE / PYRILAMINE|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE / PYRILAMINE
C2929390|T121|1008486|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-SOUTH DAKOTA-6-2007 (H1N1) (A-BRISBANE-59-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-URUGUAY -716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-FLORIDA-4-2006 STRAIN|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-SOUTH DAKOTA-6-2007 (H1N1) (A-BRISBANE-59-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-URUGUAY -716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-FLORIDA-4-2006 STRAIN
C2929391|T121|1008487|RXNORM|CITRUS PECTIN EXTRACT / LACTOBACILLUS ACIDOPHILUS|CITRUS PECTIN EXTRACT / LACTOBACILLUS ACIDOPHILUS
C2929388|T121|1008484|RXNORM|GINKGO BILOBA EXTRACT / GINKGO BILOBA LEAF EXTRACT|GINKGO BILOBA EXTRACT / GINKGO BILOBA LEAF EXTRACT
C2929389|T121|1008485|RXNORM|ACETAMINOPHEN / PHENYLEPHRINE / PHENYLTOLOXAMINE|ACETAMINOPHEN / PHENYLEPHRINE / PHENYLTOLOXAMINE
C0078596|T121|1307815|RXNORM|XANTHAN GUM|XANTHAN GUM
C3472815|T121|1307814|RXNORM|PERILLA FRUTESCENS SEED EXTRACT|PERILLA FRUTESCENS SEED EXTRACT
C3256659|T121|1307817|RXNORM|ASARUM SIEBOLDII ROOT EXTRACT|ASARUM SIEBOLDII ROOT EXTRACT
C3267745|T121|1307816|RXNORM|MAGNOLIA ACUMINATA FLOWER EXTRACT|MAGNOLIA ACUMINATA FLOWER EXTRACT
C0043892|T121|38716|RXNORM|TRIMETHYLPHLOROGLUCINOL|TRIMETHYLPHLOROGLUCINOL
C3474082|T121|1307810|RXNORM|QUERCUS SUBER BARK EXTRACT|QUERCUS SUBER BARK EXTRACT
C3256437|T121|1307812|RXNORM|PLUMERIA RUBRA FLOWER EXTRACT|PLUMERIA RUBRA FLOWER EXTRACT
C0076959|T121|38508|RXNORM|TREOSULFAN|TREOSULFAN
C3255596|T121|1307819|RXNORM|HAMAMELIS VIRGINIANA LEAF WATER EXTRACT|HAMAMELIS VIRGINIANA LEAF WATER EXTRACT
C3256671|T121|1307818|RXNORM|CAMELLIA SINENSIS ROOT EXTRACT|CAMELLIA SINENSIS ROOT EXTRACT
C3489043|T121|1358961|RXNORM|ONONIS REPENS WHOLE EXTRACT|ONONIS REPENS WHOLE EXTRACT
C3496117|T121|1358960|RXNORM|CUPRESSUS SEMPERVIRENS LEAF EXTRACT|CUPRESSUS SEMPERVIRENS LEAF EXTRACT
C3474042|T121|1358963|RXNORM|NARDOSTACHYS CHINENSIS WHOLE EXTRACT|NARDOSTACHYS CHINENSIS WHOLE EXTRACT
C3475120|T121|1358962|RXNORM|MACLURA TRICUSPIDATA WHOLE EXTRACT|MACLURA TRICUSPIDATA WHOLE EXTRACT
C0452454|T168|1358965|RXNORM|APPLE JUICE|APPLE JUICE
C3256421|T168|1358964|RXNORM|MANGO JUICE|MANGO JUICE
C0781149|T109|1358967|RXNORM|NEATSFOOT OIL|NEATSFOOT OIL
C0452458|T168|1358966|RXNORM|ORANGE JUICE|ORANGE JUICE
C0054435|T121|20032|RXNORM|BENZOATE / CAFFEINE|BENZOATE / CAFFEINE
C3662998|T121|1432296|RXNORM|CITRUS PARADISI, WHOLE EXTRACT|CITRUS PARADISI, WHOLE EXTRACT
C0762662|T121|232158|RXNORM|ROFECOXIB|ROFECOXIB
C0937641|T121|283580|RXNORM|MILK THISTLE SEED|MILK THISTLE SEED
C3486780|T121|1311274|RXNORM|SUS SCROFA BONE PREPARATION|PORCINE BONE PREPARATION
C2962856|T121|1087280|RXNORM|BORON / CALCIUM CARBONATE / CHOLECALCIFEROL / FOLIC ACID / MAGNESIUM OXIDE / PYRIDOXINE / VITAMIN B 12|BORON / CALCIUM CARBONATE / CHOLECALCIFEROL / FOLIC ACID / MAGNESIUM OXIDE / PYRIDOXINE / VITAMIN B 12
C0521965|T125|133070|RXNORM|PAROXYPROPIONE|PAROXYPROPIONE
C0046099|T109|1432294|RXNORM|2-ETHYLHEXYL ACRYLATE|2-ETHYLHEXYL ACRYLATE
C3497707|T121|1310502|RXNORM|CHLORPHENIRAMINE / IBUPROFEN / PHENYLEPHRINE|CHLORPHENIRAMINE / IBUPROFEN / PHENYLEPHRINE
C3497901|T121|1311109|RXNORM|SPONGIA OFFICINALIS PREPARATION|SPONGIA OFFICINALIS PREPARATION
C3535888|T123|1370593|RXNORM|CARNOSINE HYDROCHLORIDE|CARNOSINE HYDROCHLORIDE
C3485577|T121|1311100|RXNORM|SYMPHORICARPOS ALBUS FRUIT EXTRACT|SYMPHORICARPOS ALBUS FRUIT EXTRACT
C3485576|T121|1311101|RXNORM|SANICULA EUROPAEA EXTRACT|SANICULA EUROPAEA EXTRACT
C3486669|T121|1311102|RXNORM|CANIS LUPUS FAMILIARIS MILK PREPARATION|CANIS LUPUS FAMILIARIS MILK PREPARATION
C3497900|T197|1311103|RXNORM|YTTERBIUM OXIDE|YTTERBIUM OXIDE
C0907967|T197|1311105|RXNORM|SAMARIUM OXIDE|SAMARIUM OXIDE
C1623336|T197|1311107|RXNORM|NEODYMIUM OXIDE|NEODYMIUM OXIDE
C3152977|T121|1098425|RXNORM|NIACINAMIDE / PANTHENOL / ZINC PYRITHIONE|NIACINAMIDE / PANTHENOL / ZINC PYRITHIONE
C3848567|T196|1546280|RXNORM|NICKEL CATION|NICKEL CATION
C3848565|T196|1546283|RXNORM|ANTIMONY CATION (5+)|ANTIMONY CATION (5+)
C2948028|T121|1309199|RXNORM|ALOE VERA FLOWER EXTRACT|ALOE VERA FLOWER EXTRACT
C0025760|T121|6883|RXNORM|METHYLERGONOVINE|METHYLERGONOVINE
C2927972|T121|1007049|RXNORM|IODOPHORS / ISOPROPYL ALCOHOL|IODOPHORS / ISOPROPYL ALCOHOL
C2927971|T121|1007048|RXNORM|POVIDONE / TETRAHYDROZOLINE|POVIDONE / TETRAHYDROZOLINE
C2927970|T121|1007047|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-URUGUAY-716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-FLORIDA-4-2006 STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-URUGUAY-716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-FLORIDA-4-2006 STRAIN
C2927969|T121|1007046|RXNORM|CALCIUM CHLORIDE / GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CHLORIDE / GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / SODIUM CHLORIDE
C2927968|T121|1007045|RXNORM|DICHLORODIFLUOROMETHANE / ETHYL CHLORIDE|DICHLORODIFLUOROMETHANE / ETHYL CHLORIDE
C2927967|T121|1007044|RXNORM|POLOXAMER 407 / SIMETHICONE|POLOXAMER 407 / SIMETHICONE
C2927966|T121|1007043|RXNORM|GREEN TEA LEAF EXTRACT / THEAFLAVIN|GREEN TEA LEAF EXTRACT / THEAFLAVIN
C2927965|T121|1007042|RXNORM|GARLIC PREPARATION / LECITHIN|GARLIC PREPARATION / LECITHIN
C3282782|T121|1313241|RXNORM|ISOEICOSANE|ISOEICOSANE
C3502969|T123|1370594|RXNORM|LAURATE|LAURATE
C1875534|T121|691448|RXNORM|NIACIN / PHENIRAMINE|NIACIN / PHENIRAMINE
C3256134|T121|1426393|RXNORM|COCO MONOETHANOLAMIDE|COCO MONOETHANOLAMIDE
C1451406|T195|1309314|RXNORM|TULATHROMYCIN|TULATHROMYCIN
C1875533|T121|691447|RXNORM|NIACIN / PENTYLENETETRAZOLE|NIACIN / PENTYLENETETRAZOLE
C1875530|T121|691444|RXNORM|NIACIN / NIACINAMIDE / PHENOBARBITAL|NIACIN / NIACINAMIDE / PHENOBARBITAL
C3535887|T109|1370595|RXNORM|STARCH GLYCOLATE TYPE A CORN|STARCH GLYCOLATE TYPE A CORN
C3488975|T109|1309310|RXNORM|OREGANO FLOWERING TOP EXTRACT|OREGANO FLOWERING TOP EXTRACT
C0074751|T197|1364915|RXNORM|SODIUM PERCARBONATE|SODIUM PERCARBONATE
C0757571|T121|1426897|RXNORM|QUATERNIUM-22|QUATERNIUM-22
C0164505|T121|59695|RXNORM|CHLOROTHEN|CHLOROTHEN
C3488331|T121|1336266|RXNORM|ANAGALLIS ARVENSIS EXTRACT|ANAGALLIS ARVENSIS EXTRACT
C3488470|T121|1336267|RXNORM|ARTEMISIA ABROTANUM FLOWERING TOP EXTRACT|ARTEMISIA ABROTANUM FLOWERING TOP EXTRACT
C3484461|T121|1336264|RXNORM|CHIMAPHILA MACULATA EXTRACT|CHIMAPHILA MACULATA EXTRACT
C0065841|T195|29418|RXNORM|MECLOCYCLINE|MECLOCYCLINE
C3488422|T121|1426396|RXNORM|SEA SCALLOP PREPARATION|SEA SCALLOP PREPARATION
C0065834|T121|29411|RXNORM|MEBHYDROLINE|MEBHYDROLIN
C3834238|T121|1541621|RXNORM|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-TEXAS-50-2012 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-BRISBANE-60-2008-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-TEXAS-50-2012 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-BRISBANE-60-2008-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS
C3489124|T121|1336269|RXNORM|GRATIOLA OFFICINALIS EXTRACT|GRATIOLA OFFICINALIS EXTRACT
C0108111|T121|47618|RXNORM|CALCIUM GLUCEPTATE|CALCIUM GLUCOHEPTONATE
C3535883|T121|1370599|RXNORM|RICINOLEIC MONOETHANOLAMIDE SULFOSUCCINATE|RICINOLEIC MONOETHANOLAMIDE SULFOSUCCINATE
C3256642|T109|1426394|RXNORM|POLYQUATERNIUM-7 (70-30 ACRYLAMIDE-DADMAC; 1600 KD)|POLYQUATERNIUM-7 (70-30 ACRYLAMIDE-DADMAC 1600000 MW)
C0108092|T122|47610|RXNORM|CALCIUM ALGINATE|CALCIUM ALGINATE
C0108101|T121|47613|RXNORM|CALCIUM CITRATE|CALCIUM CITRATE
C3256705|T109|1426395|RXNORM|OCTOXYNOL-40|OCTOXYNOL-40
C0108108|T121|47617|RXNORM|CALCIUM GALACTOGLUCONATE BROMIDE|CALCIUM GALACTOGLUCONATE BROMIDE
C0004147|T121|1202|RXNORM|ATENOLOL|ATENOLOL
C2928517|T121|1007599|RXNORM|HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / PHENYL SALICYLATE|HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / PHENYL SALICYLATE
C2928516|T121|1007598|RXNORM|ECHINACEA PREPARATION / GOLDENSEAL EXTRACT|ECHINACEA PREPARATION / GOLDENSEAL EXTRACT
C2928191|T121|1007269|RXNORM|ACETAMINOPHEN / GUAIFENESIN / PSEUDOEPHEDRINE|ACETAMINOPHEN / GUAIFENESIN / PSEUDOEPHEDRINE
C2928190|T121|1007268|RXNORM|FENUGREEK SEED PREPARATION / LEGUME PREPARATION|FENUGREEK SEED PREPARATION / LEGUME PREPARATION
C2928185|T121|1007263|RXNORM|ESTRADIOL / PREDNISOLONE|ESTRADIOL / PREDNISOLONE
C2928184|T121|1007262|RXNORM|BISACODYL / DOCUSATE|BISACODYL / DOCUSATE
C2928183|T121|1007261|RXNORM|PREDNISOLONE / RIFAMYCINS|PREDNISOLONE / RIFAMYCINS
C2928182|T121|1007260|RXNORM|OXYTETRACYCLINE / PREDNISOLONE|OXYTETRACYCLINE / PREDNISOLONE
C2928189|T121|1007267|RXNORM|PRAMOXINE / ZINC SULFATE|PRAMOXINE / ZINC SULFATE
C2928188|T121|1007266|RXNORM|LACTATE / PRAMOXINE|LACTATE / PRAMOXINE
C2928515|T121|1007597|RXNORM|FERROUS PHOSPHATE / POTASSIUM CHLORIDE|FERROUS PHOSPHATE / POTASSIUM CHLORIDE
C2928186|T121|1007264|RXNORM|OXYQUINOLINE / PREDNISOLONE|OXYQUINOLINE / PREDNISOLONE
C0040899|T121|10772|RXNORM|TRICHLORMETHIAZIDE|TRICHLORMETHIAZIDE
C3531402|T109|1366737|RXNORM|LIMONIUM GERBERI FLOWERING TOP EXTRACT|LIMONIUM GERBERI FLOWERING TOP EXTRACT
C3531403|T109|1366739|RXNORM|DECAMETHYLTETRASILOXANE|DECAMETHYLTETRASILOXANE
C2701423|T129|852225|RXNORM|CHEAT GRASS POLLEN EXTRACT|BROMUS SECALINUS POLLEN EXTRACT
C1874699|T121|691192|RXNORM|CAMPHOR / PARACHLOROPHENOL|CAMPHOR / PARACHLOROPHENOL
C0009185|T130|2660|RXNORM|COCCIDIOIDIN|COCCIDIOIDIN
C0244821|T121|72302|RXNORM|ROPINIROLE|ROPINIROLE
C0873075|T121|259412|RXNORM|GRIFFONIA PREPARATION|GRIFFONIA PREPARATION
C3848588|T121|1545791|RXNORM|POPULUS TREMULA WHOLE EXTRACT|POPULUS TREMULA WHOLE EXTRACT
C3499588|T121|1312458|RXNORM|PETROLATUM / VITAMIN E|PETROLATUM / VITAMIN E
C2746119|T129|901636|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 7F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 7F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C2919267|T126|901805|RXNORM|VELAGLUCERASE ALFA|VELAGLUCERASE ALFA
C0896320|T121|273888|RXNORM|CALCIUM THREONATE|CALCIUM THREONATE
C0073631|T121|35827|RXNORM|KETOROLAC|KETOROLAC
C0073631|T121|35827|RXNORM|KETOROLAC|KETOROLAC
C3661282|T121|1455099|RXNORM|VORTIOXETINE|VORTIOXETINE
C2929968|T121|1009073|RXNORM|MERADIMATE / TITANIUM DIOXIDE|MERADIMATE / TITANIUM DIOXIDE
C0037215|T121|9808|RXNORM|SITOSTEROLS|SITOSTEROLS
C0673966|T121|194881|RXNORM|BRINZOLAMIDE|BRINZOLAMIDE
C0073633|T121|35829|RXNORM|RANOLAZINE|RANOLAZINE
C0037167|T125|9800|RXNORM|SINCALIDE|SINCALIDE
C0813211|T121||RXNORM|HYDROCHLOROTHIAZIDE / TRIAMTERENE
C0874047|T121|260020|RXNORM|HORSE CHESTNUT SEED|HORSE CHESTNUT SEED
C0301478|T121|89870|RXNORM|OX BILE EXTRACT|OX BILE EXTRACT
C0171302|T121|61455|RXNORM|MIZOLASTINE|MIZOLASTINE
C0724516|T121|221053|RXNORM|ADIASTATIC BARLEY MALT EXTRACT|ADIASTATIC BARLEY MALT EXTRACT
C0772239|T121|236911|RXNORM|ZINC CITRATE|ZINC CITRATE
C0302211|T197|90120|RXNORM|MAGNESIUM SALT|MAGNESIUM SALT
C2722029|T129|862453|RXNORM|BARLEY ALLERGENIC EXTRACT|BARLEY ALLERGENIC EXTRACT
C0982183|T121|1367188|RXNORM|GLYCOL DISTEARATE|GLYCOL DISTEARATE
C1095905|T121|319826|RXNORM|BEETS PREPARATION|BEET JUICE
C0175162|T121|1360721|RXNORM|THONZYLAMINE|THONZYLAMINE
C1577357|T121|486456|RXNORM|METHYLFOLIC ACID|METHYLFOLIC ACID
C3644809|T109|1425900|RXNORM|ROSA CANINA FLOWER OIL|ROSA CANINA FLOWER OIL
C0015058|T121|4141|RXNORM|ETHYL CHLORIDE|ETHYL CHLORIDE
C3488281|T121|1351789|RXNORM|CASTORBEAN SEED EXTRACT|CASTORBEAN SEED EXTRACT
C2116317|T121|812786|RXNORM|AMILORIDE / HYDROCHLOROTHIAZIDE / TIMOLOL|AMILORIDE / HYDROCHLOROTHIAZIDE / TIMOLOL
C0982459|T121|314896|RXNORM|WHEAT GERM PREPARATION|WHEAT GERM PREPARATION
C3486736|T121|1351786|RXNORM|BETULA PENDULA LEAF EXTRACT|BETULA PENDULA LEAF EXTRACT
C3267239|T121|1245705|RXNORM|CHLOPHEDIANOL / CHLORPHENIRAMINE / PHENYLEPHRINE|CHLOPHEDIANOL / CHLORPHENIRAMINE / PHENYLEPHRINE
C0717592|T121|214395|RXNORM|CHLORPHENIRAMINE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / PSEUDOEPHEDRINE
C0717591|T121|214394|RXNORM|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE
C0717587|T121|214390|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN|CHLORPHENIRAMINE / DEXTROMETHORPHAN
C0717590|T121|214393|RXNORM|CHLORPHENIRAMINE / PHENYLEPHRINE|CHLORPHENIRAMINE / PHENYLEPHRINE
C0717589|T121|214392|RXNORM|CHLORPHENIRAMINE / HYDROCODONE|CHLORPHENIRAMINE / HYDROCODONE
C2940189|T129|1014739|RXNORM|BITTER DOCK POLLEN EXTRACT|RUMEX OBTUSIFOLIUS POLLEN EXTRACT
C3486696|T121|1313275|RXNORM|ACONITIC ACID, (Z)-|ACONITIC ACID, (Z)-
C2700070|T121|1426386|RXNORM|TRIBEHENIN|TRIBEHENIN
C3473019|T122|1313270|RXNORM|POLYACRYLAMIDE (CROSSLINKED; 0.01-0.2 MOLE PERCENT BISACRYLAMIDE)|POLYACRYLAMIDE (CROSSLINKED; 0.01-0.2 MOLE PERCENT BISACRYLAMIDE)
C3473023|T109|1313271|RXNORM|RIMETHYLOLPROPANE TRICAPRYLATE-TRICAPRATE|RIMETHYLOLPROPANE TRICAPRYLATE-TRICAPRATE
C3255595|T109|1426382|RXNORM|HAEMATOCOCCUS PLUVIALIS EXTRACT|HAEMATOCOCCUS PLUVIALIS EXTRACT
C2940183|T129|1014731|RXNORM|CANADIAN BLUEGRASS POLLEN EXTRACT|POA COMPRESSA POLLEN EXTRACT
C2701431|T129|852233|RXNORM|BOTTLEBRUSH POLLEN EXTRACT|MELALEUCA CITRINA POLLEN EXTRACT
C1571583|T121|1037042|RXNORM|DABIGATRAN ETEXILATE|DABIGATRAN ETEXILATE
C2940186|T129|1014735|RXNORM|WHITE SWEET CLOVER POLLEN EXTRACT|MELILOTUS ALBUS POLLEN EXTRACT
C3489391|T121|1313279|RXNORM|URANYL NITRATE HEXAHYDRATE|URANYL NITRATE HEXAHYDRATE
C1106203|T121|323994|RXNORM|ALFALFA OIL|ALFALFA OIL
C2827241|T121|1364479|RXNORM|LOMITAPIDE|LOMITAPIDE
C3256282|T109|1424679|RXNORM|CANDELILLA WAX POWDER|CANDELILLA WAX POWDER
C2929017|T121|1008109|RXNORM|BAMETHAN / TROXERUTIN|BAMETHAN / TROXERUTIN
C2929016|T121|1008108|RXNORM|ALGESTONE / ESTRADIOL|ALGESTONE / ESTRADIOL
C2929015|T121|1008107|RXNORM|CETRIMONIUM / CHLORHEXIDINE|CETRIMONIUM / CHLORHEXIDINE
C2929014|T121|1008106|RXNORM|BORIC ACID / PHENOL|BORIC ACID / PHENOL
C2929013|T121|1008105|RXNORM|TOLNAFTATE / TRIACETIN|TOLNAFTATE / TRIACETIN
C2929012|T121|1008104|RXNORM|ALLANTOIN / DYCLONINE|ALLANTOIN / DYCLONINE
C2929011|T121|1008103|RXNORM|BETAXOLOL / PILOCARPINE|BETAXOLOL / PILOCARPINE
C2929009|T121|1008101|RXNORM|P-HYDROXYAMPHETAMINE / TROPICAMIDE|P-HYDROXYAMPHETAMINE / TROPICAMIDE
C2929008|T121|1008100|RXNORM|ASCORBIC ACID / VITAMIN E|ASCORBIC ACID / VITAMIN E
C0069751|T121|32624|RXNORM|OXCARBAZEPINE|OXCARBAZEPINE
C0069753|T121|32626|RXNORM|OXELADIN|OXELADIN
C0076649|T121|38249|RXNORM|TIADILON|TIADILON
C2725893|T129|974129|RXNORM|SARDINE ALLERGENIC EXTRACT|EUROPEAN PILCHARD ALLERGENIC EXTRACT
C0037114|T122|9778|RXNORM|SILICONES|SILICONES
C0357929|T121|106212|RXNORM|CALAMINE|CALAMINE
C3255747|T109|1306195|RXNORM|CHENOPODIUM QUINOA SEED EXTRACT|CHENOPODIUM QUINOA SEED EXTRACT
C3255745|T109|1306194|RXNORM|CHAMAEMELUM NOBILE FLOWER EXTRACT|CHAMAEMELUM NOBILE FLOWER EXTRACT
C3255742|T109|1306193|RXNORM|BELLIS PERENNIS FLOWER EXTRACT|BELLIS PERENNIS FLOWER EXTRACT
C3255741|T109|1306192|RXNORM|BEHENYL PHOSPHATE|BEHENYL PHOSPHATE
C3255740|T109|1306191|RXNORM|BEACH STRAWBERRY EXTRACT|BEACH STRAWBERRY EXTRACT
C3255739|T109|1306190|RXNORM|BATILOL|BATILOL
C3257291|T109|1368157|RXNORM|PEG-10 DIMETHICONE (600 CST)|PEG-10 DIMETHICONE (600 CST)
C3245080|T121|1368156|RXNORM|PEG-150 STEARATE|PEG-150 STEARATE
C3535618|T109|1368155|RXNORM|PEG-30 STEARATE|PEG-30 STEARATE
C0015087|T131|1368154|RXNORM|ETHYLENE OXIDE|ETHYLENE OXIDE
C0055754|T121|1368153|RXNORM|CINNAMIC ALDEHYDE|CINNAMALDEHYDE
C3473981|T121|1368152|RXNORM|CHITOSAN MEDIUM MOLECULAR WEIGHT (200-800 MPA.S)|CHITOSAN MEDIUM MOLECULAR WEIGHT (200-800 MPA.S)
C3255905|T109|1306199|RXNORM|ALFALFA SEED EXTRACT|ALFALFA SEED EXTRACT
C3535925|T121|1368402|RXNORM|ALOGLIPTIN / PIOGLITAZONE|ALOGLIPTIN / PIOGLITAZONE
C0031705|T196|8263|RXNORM|PHOSPHORUS|PHOSPHORUS
C0304114|T121|90945|RXNORM|ROSEMARY OIL|ROSEMARY OIL
C1722685|T121|658708|RXNORM|ECALLANTIDE|ECALLANTIDE
C0016673|T195|4556|RXNORM|FRAMYCETIN|FRAMYCETIN
C0054838|T121|1368148|RXNORM|CARYOPHYLLENE|CARYOPHYLLENE
C0016610|T195|4550|RXNORM|FOSFOMYCIN|FOSFOMYCIN
C3472714|T121|1368149|RXNORM|CENTAURIUM ERYTHRAEA PREPARATION|CENTAURIUM ERYTHRAEA PREPARATION
C0032823|T123|8589|RXNORM|POTASSIUM ASPARTATE|POTASSIUM ASPARTATE
C3832971|T109|1540025|RXNORM|EUCALYPTUS CAMALDULENSIS LEAF OIL|EUCALYPTUS CAMALDULENSIS LEAF OIL
C3162761|T121|1114858|RXNORM|MELATONIN / VITAMIN B 12|MELATONIN / VITAMIN B 12
C1815866|T121|670544|RXNORM|SANGUINARIA CANADENSIS ROOT EXTRACT|SANGUINARIA CANADENSIS ROOT EXTRACT
C3256496|T121|1309395|RXNORM|ACORUS CALAMUS ROOT EXTRACT|ACORUS CALAMUS ROOT EXTRACT
C2344269|T129|798224|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 19F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 19F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C3162754|T121|1114850|RXNORM|CHLOROPHYLL / GARLIC PREPARATION / PARSLEY EXTRACT|CHLOROPHYLL / GARLIC PREPARATION / PARSLEY EXTRACT
C0291772|T121|85248|RXNORM|ALOSETRON|ALOSETRON
C0060234|T197|24902|RXNORM|PRUSSIAN BLUE|PRUSSIAN BLUE
C3485004|T121|1307573|RXNORM|ANGELICA PUBESCENS ROOT EXTRACT|ANGELICA PUBESCENS ROOT EXTRACT
C3256539|T121|1307570|RXNORM|IRVINGIA GABONENSIS SEED EXTRACT|IRVINGIA GABONENSIS SEED EXTRACT
C2827072|T130|1307571|RXNORM|1,4-SORBITAN|1,4-SORBITAN
C3256656|T121|1307576|RXNORM|ALCEA ROSEA FLOWER EXTRACT|ALCEA ROSEA FLOWER EXTRACT
C3256146|T121|1307577|RXNORM|COPTIS JAPONICA ROOT EXTRACT|COPTIS JAPONICA ROOT EXTRACT
C3464709|T121|1307574|RXNORM|CHENOPODIUM ALBUM FLOWER EXTRACT|CHENOPODIUM ALBUM FLOWER EXTRACT
C3256721|T121|1307575|RXNORM|SANGUISORBA MINOR ROOT EXTRACT|SANGUISORBA MINOR ROOT EXTRACT
C3256710|T121|1307578|RXNORM|OENOTHERA BIENNIS LEAF EXTRACT|OENOTHERA BIENNIS LEAF EXTRACT
C0060241|T121|24909|RXNORM|FERRIC OXIDE, SACCHARATED|IRON SACCHARATE
C0302236|T129|979384|RXNORM|NORTH AMERICAN CORAL SNAKE ANTIVENIN|NORTH AMERICAN CORAL SNAKE ANTIVENIN
C0020275|T196|5497|RXNORM|HYDROGEN|HYDROGEN
C0440280|T121|124323|RXNORM|GRAPEFRUIT EXTRACT|GRAPEFRUIT EXTRACT
C3256293|T109|1368140|RXNORM|BUTYL ESTER OF METHYL VINYL ETHER-MALEIC ANHYDRIDE COPOLYMER (125 KD)|BUTYL ESTER OF METHYL VINYL ETHER/MALEIC ANHYDRIDE COPOLYMER (125000 MW)
C0063953|T121|27901|RXNORM|ISOCONAZOLE|ISOCONAZOLE
C3257292|T109|1368141|RXNORM|BUTYLENE GLYCOL DICAPRYLATE-DICAPRATE|BUTYLENE GLYCOL DICAPRYLATE-DICAPRATE
C2746961|T129|904507|RXNORM|EGG (CHICKEN) ALLERGENIC EXTRACT|EGG (CHICKEN) ALLERGENIC EXTRACT
C0060629|T121|25231|RXNORM|FOMOCAIN|FOMOCAIN
C0015843|T121|4335|RXNORM|FENSPIRIDE|FENSPIRIDE
C3488448|T121|1310133|RXNORM|ONOSMODIUM VIRGINIANUM WHOLE EXTRACT|ONOSMODIUM VIRGINIANUM WHOLE EXTRACT
C2726970|T129|885750|RXNORM|SOUTHERN RAGWEED POLLEN EXTRACT|AMBROSIA BIDENTATA POLLEN EXTRACT
C2344267|T129|798222|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 18C CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 18C CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C1301996|T121|392458|RXNORM|DAPSONE / PYRIMETHAMINE|DAPSONE / PYRIMETHAMINE
C1301995|T121|392457|RXNORM|PHYSOSTIGMINE / PILOCARPINE|PHYSOSTIGMINE / PILOCARPINE
C1301992|T121|392454|RXNORM|BENZOYL PEROXIDE / HYDROCORTISONE|BENZOYL PEROXIDE / HYDROCORTISONE
C2740303|T121|898430|RXNORM|DIHYDROCODEINE / PHENYLEPHRINE / PYRILAMINE|DIHYDROCODEINE / PHENYLEPHRINE / PYRILAMINE
C0060274|T197|473387|RXNORM|FERUMOXYTOL|FERUMOXYTOL
C0086444|T121|42736|RXNORM|DEXRAZOXANE|DEXRAZOXANE
C2719767|T129|860189|RXNORM|ONABOTULINUMTOXINA|ONABOTULINUMTOXINA
C2719767|T129|860189|RXNORM|ONABOTULINUMTOXINA|ONABOTULINUMTOXINA
C0055011|T195|20489|RXNORM|CEFPODOXIME|CEFPODOXIME
C2927830|T121|1006906|RXNORM|SODIUM BICARBONATE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC|SODIUM BICARBONATE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC
C0055004|T195|20482|RXNORM|CEFETAMET|CEFETAMET
C0055003|T195|20481|RXNORM|CEFEPIME|CEFEPIME
C1958588|T121|1592684|RXNORM|DIRLOTAPIDE|DIRLOTAPIDE
C0055008|T195|20486|RXNORM|CEFORANIDE|CEFORANIDE
C0055007|T195|20485|RXNORM|CEFODIZIME|CEFODIZIME
C0040976|T130|10798|RXNORM|TRIENTINE|TRIENTINE
C0040958|T121|10795|RXNORM|TRICLOSAN|TRICLOSAN
C0040958|T121|10795|RXNORM|TRICLOSAN|TRICLOSAN
C1874860|T121|689842|RXNORM|CITRIC ACID / SIMETHICONE / SODIUM BICARBONATE|CITRIC ACID / SIMETHICONE / SODIUM BICARBONATE
C1874859|T121|689841|RXNORM|CITRIC ACID / POTASSIUM CITRATE / SODIUM CITRATE|CITRIC ACID / POTASSIUM CITRATE / SODIUM CITRATE
C3663395|T121|1432976|RXNORM|CYBERLINDNERA JADINII RNA|CYBERLINDNERA JADINII RNA
C3663394|T121|1432975|RXNORM|CAPRIC DIETHANOLAMIDE|CAPRIC DIETHANOLAMIDE
C3486754|T109|1427168|RXNORM|LING PREPARATION|LING PREPARATION
C3818739|T121|1495206|RXNORM|VERBASCUM DENSIFLORUM FLOWER EXTRACT|VERBASCUM DENSIFLORUM FLOWER EXTRACT
C3500831|T121|1356131|RXNORM|SUS SCROFA DANDER PREPARATION|SUS SCROFA DANDER PREPARATION
C2194082|T121|812838|RXNORM|BROMAZEPAM / DOMPERIDONE / SIMETHICONE|BROMAZEPAM / DOMPERIDONE / SIMETHICONE
C0771949|T121|236649|RXNORM|PROCYANIDOLIC OLIGOMER|PROCYANIDOLIC OLIGOMER
C2741542|T129|901382|RXNORM|LEMON ALLERGENIC EXTRACT|CITRUS LIMON ALLERGENIC EXTRACT
C0771575|T121|236315|RXNORM|GUAIETOLIN|GUAIETOLIN
C0771574|T121|236314|RXNORM|GUAIACOL ETHYLGLYCOLATE|GUAIACOL ETHYLGLYCOLATE
C0982419|T121|1426355|RXNORM|STEARYL HEPTANOATE|STEARYL HEPTANOATE
C3488925|T121|1320410|RXNORM|CENTAUREA BENEDICTA EXTRACT|CENTAUREA BENEDICTA EXTRACT
C3489145|T121|1320411|RXNORM|AQUILEGIA VULGARIS EXTRACT|AQUILEGIA VULGARIS EXTRACT
C2938403|T130|1012179|RXNORM|WHITE KIDNEY BEAN ALLERGENIC EXTRACT|PHASEOLUS VULGARIS ALLERGENIC EXTRACT
C3663396|T121|1432978|RXNORM|DEHYDROABIETATE|DEHYDROABIETATE
C0051711|T121|1310190|RXNORM|AMMONIUM CARBONATE|AMMONIUM CARBONATE
C3486858|T121|1310193|RXNORM|MERCURIUS SOLUBILIS PREPARATION|MERCURIUS SOLUBILIS PREPARATION
C3700993|T121|1485894|RXNORM|PANTHENOL / ZINC PYRITHIONE|PANTHENOL / ZINC PYRITHIONE
C0038807|T121|10240|RXNORM|SULTHIAME|SULTIAME
C2702351|T129|891771|RXNORM|APPLE ALLERGENIC EXTRACT|APPLE ALLERGENIC EXTRACT
C0026259|T121|7005|RXNORM|MITOXANTRONE|MITOXANTRONE
C0026256|T121|7004|RXNORM|MITOTANE|MITOTANE
C0038838|T126|10245|RXNORM|SUPEROXIDE DISMUTASE|SUPEROXIDE DISMUTASE
C2937983|T129|1010999|RXNORM|NECTARINE ALLERGENIC EXTRACT|NECTARINE ALLERGENIC EXTRACT
C0027608|T196|7301|RXNORM|NEON|NEON
C0070563|T121|33283|RXNORM|PHENINDAMINE|PHENINDAMINE
C3256119|T121|1305555|RXNORM|ALUMINUM DIMYRISTATE|ALUMINUM DIMYRISTATE
C0044438|T131|1305552|RXNORM|1-METHYL-2-PYRROLIDINONE|METHYL PYRROLIDONE
C0052865|T195|18687|RXNORM|BACAMPICILLIN|BACAMPICILLIN
C3256294|T109|1305550|RXNORM|CANNABIS SATIVA SEED OIL|CANNABIS SATIVA SEED OIL
C3152269|T129|1305551|RXNORM|CARYA LACINIOSA POLLEN EXTRACT|CARYA LACINIOSA POLLEN EXTRACT
C1144149|T121|342369|RXNORM|LENALIDOMIDE|LENALIDOMIDE
C3864845|T129|1595881|RXNORM|COTTONMOUTH VENOM|AGKISTRODON PISCIVORUS VENOM
C0580776|T131|1595880|RXNORM|GILA MONSTER VENOM|HELODERMA SUSPECTUM VENOM
C1998431|T130|1305558|RXNORM|AMMONIA N-13|AMMONIA N-13
C3465351|T109|1305559|RXNORM|AMMONIUM ACRYLODIMETHYLTAURATE|AMMONIUM ACRYLODIMETHYLTAURATE
C1631068|T121|608566|RXNORM|CETYLPYRIDINIUM / LIDOCAINE|CETYLPYRIDINIUM / LIDOCAINE
C1628498|T121|608568|RXNORM|LIDOCAINE / TETRACAINE|LIDOCAINE / TETRACAINE
C0002711|T121|742|RXNORM|AMYL NITRITE|AMYL NITRITE
C0002711|T121|742|RXNORM|AMYL NITRITE|AMYL NITRITE
C0002712|T126|743|RXNORM|AMYLASES|AMYLASES
C0021745|T129|5885|RXNORM|INTERFERON TYPE II|INTERFERON TYPE II
C0066485|T121|1442202|RXNORM|MEVALONOLACTONE|MEVALONOLACTONE
C0997449|T004|1442200|RXNORM|MONASCUS PURPUREUS|RED YEAST
C2927655|T129|1006506|RXNORM|TALL OAT GRASS POLLEN EXTRACT|ARRHENATHERUM ELATIUS POLLEN EXTRACT
C0937851|T121|283746|RXNORM|TASONERMIN|TASONERMIN
C1874913|T121|690105|RXNORM|COLISTIN / HYDROCORTISONE / NEOMYCIN / THONZONIUM|COLISTIN / HYDROCORTISONE / NEOMYCIN / THONZONIUM
C0003639|T121|1054|RXNORM|APRINDINE|APRINDINE
C1874908|T121|690101|RXNORM|CODEINE / PYRILAMINE|CODEINE / PYRILAMINE
C0003641|T123|1056|RXNORM|APROTININ|APROTININ
C1509720|T121|1368184|RXNORM|NONOXYNOL-4|NONOXYNOL-4
C2731457|T129|895353|RXNORM|COOTAMUNDRA WATTLE POLLEN EXTRACT|COOTAMUNDRA WATTLE POLLEN EXTRACT
C3667898|T121|1440278|RXNORM|PLATANUS OCCIDENTALIS WHOLE EXTRACT|PLATANUS OCCIDENTALIS WHOLE EXTRACT
C2928816|T121|1007902|RXNORM|CORNSTARCH / KAOLIN / ZINC OXIDE|CORNSTARCH / KAOLIN / ZINC OXIDE
C2928817|T121|1007903|RXNORM|BUTAMBEN / NITROMERSOL|BUTAMBEN / NITROMERSOL
C2928814|T121|1007900|RXNORM|BENZYL ALCOHOL / PRAMOXINE|BENZYL ALCOHOL / PRAMOXINE
C2928815|T121|1007901|RXNORM|GUAIFENESIN / PHENYLEPHRINE / POTASSIUM CITRATE|GUAIFENESIN / PHENYLEPHRINE / POTASSIUM CITRATE
C2928820|T121|1007906|RXNORM|CIDER VINEGAR / KELP PREPARATION / LECITHIN / VITAMIN B6|CIDER VINEGAR / KELP PREPARATION / LECITHIN / VITAMIN B6
C2928821|T121|1007907|RXNORM|FRAMYCETIN / HYDROCORTISONE|FRAMYCETIN / HYDROCORTISONE
C2928818|T121|1007904|RXNORM|DEXTROMETHORPHAN / PHENYLEPHRINE / SODIUM CITRATE|DEXTROMETHORPHAN / PHENYLEPHRINE / SODIUM CITRATE
C2928819|T121|1007905|RXNORM|SULFONATED PHENOL / SULFURIC ACID|SULFONATED PHENOL / SULFURIC ACID
C2826347|T196|1334548|RXNORM|BARIUM CATION|BARIUM CATION
C2928822|T121|1007908|RXNORM|CHOLINE / CYSTEINE|CHOLINE / CYSTEINE
C2928823|T121|1007909|RXNORM|NALOXONE / TILIDINE|NALOXONE / TILIDINE
C3645180|T122|1426830|RXNORM|COCOAMPHOACETATE|COCOAMPHOACETATE
C0015772|T121|4316|RXNORM|FELODIPINE|FELODIPINE
C0015777|T121|4319|RXNORM|FELYPRESSIN|FELYPRESSIN
C0026926|T007|1492936|RXNORM|MYCOBACTERIUM TUBERCULOSIS|MYCOBACTERIUM TUBERCULOSIS
C0526399|T121|135056|RXNORM|LERCANIDIPINE|LERCANIDIPINE
C2928434|T121|1007512|RXNORM|CALCIUM CITRATE / ERGOCALCIFEROL|CALCIUM CITRATE / ERGOCALCIFEROL
C2929206|T121|1008299|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 16 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 16 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18 VACCINE
C2929205|T121|1008298|RXNORM|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE
C2929204|T121|1008297|RXNORM|CLORSULON / IVERMECTIN|CLORSULON / IVERMECTIN
C2929203|T121|1008296|RXNORM|PALM OIL / SOYBEAN OIL|PALM OIL / SOYBEAN OIL
C2929202|T121|1008295|RXNORM|ACETAMINOPHEN / CLEMASTINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / CLEMASTINE / PSEUDOEPHEDRINE
C2929201|T121|1008294|RXNORM|MICONAZOLE / POLYMYXIN B / PREDNISOLONE|MICONAZOLE / POLYMYXIN B / PREDNISOLONE
C2929200|T121|1008293|RXNORM|CUPROUS OXIDE / FOLIC ACID / NIACINAMIDE / ZINC OXIDE|CUPROUS OXIDE / FOLIC ACID / NIACINAMIDE / ZINC OXIDE
C2929199|T121|1008292|RXNORM|BERBERINE / CHOLECALCIFEROL / HOPS EXTRACT / VITAMIN K|BERBERINE / CHOLECALCIFEROL / HOPS EXTRACT / VITAMIN K
C2929198|T121|1008291|RXNORM|PHYTOSTEROLS / SAW PALMETTO EXTRACT|PHYTOSTEROLS / SAW PALMETTO EXTRACT
C2929197|T121|1008290|RXNORM|GLUCOSAMINE / HYALURONATE / METHYLSULFONYLMETHANE|GLUCOSAMINE / HYALURONATE / METHYLSULFONYLMETHANE
C0358859|T121|106846|RXNORM|AMPICILLIN / CLOXACILLIN|AMPICILLIN / CLOXACILLIN
C0011082|T121|3118|RXNORM|DEBRISOQUIN|DEBRISOQUIN
C0011064|T121|3116|RXNORM|DEANOL|DEANOL
C2073874|T121|815781|RXNORM|CHLORPHENIRAMINE / PHENYLEPHRINE / SCOPOLAMINE|CHLORPHENIRAMINE / PHENYLEPHRINE / SCOPOLAMINE
C0937631|T121|283571|RXNORM|HAWTHORN BERRY EXTRACT|HAWTHORN BERRY EXTRACT
C3832869|T121|1539809|RXNORM|CETEARYL NONANOATE|CETEARYL NONANOATE
C3464714|T121|1312738|RXNORM|POLYETHYLENE GLYCOL 400000|POLYETHYLENE GLYCOL 400000
C0076130|T109|1312739|RXNORM|TERPINYL ACETATE|TERPINYL ACETATE
C3500689|T121|1315108|RXNORM|ARCHED SWIMMING CRAB, COOKED PREPARATION|ARCHED SWIMMING CRAB, COOKED PREPARATION
C3500690|T121|1315109|RXNORM|CASEIN, EMMENTAL CULTURED|CASEIN, EMMENTAL CULTURED
C0937638|T121|283577|RXNORM|LYCOPODIUM CLAVATUM PREPARATION|LYCOPODIUM CLAVATUM PREPARATION
C2726183|T129|995727|RXNORM|MYCOCLADUS CORYMBIFERUS EXTRACT|MYCOCLADUS CORYMBIFERUS EXTRACT
C3496664|T121|1312732|RXNORM|TORREYA NUCIFERA WHOLE EXTRACT|TORREYA NUCIFERA WHOLE EXTRACT
C0937639|T121|283578|RXNORM|MAGNESIUM MALATE|MAGNESIUM MALATE
C3265135|T121|1312730|RXNORM|QUATERNIUM-14|QUATERNIUM-14
C3265585|T121|1312731|RXNORM|POLYETHYLENE GLYCOL 7000000|POLYETHYLENE GLYCOL 7000000
C3281531|T121|1312736|RXNORM|POLYISOBUTYLENE (2300 MW)|POLYISOBUTYLENE (2300 MW)
C0032952|T125|8640|RXNORM|PREDNISONE|PREDNISONE
C3465316|T109|1427228|RXNORM|POLY(METHYL ACRYLATE-CO-METHYL METHACRYLATE-CO-METHACRYLIC ACID 7:3:1; 280000 MW)|POLY(METHYL ACRYLATE-CO-METHYL METHACRYLATE-CO-METHACRYLIC ACID 7:3:1; 280000 MW)
C0068353|T121|31462|RXNORM|NADOXOLOL|NADOXOLOL
C0754820|T130|228833|RXNORM|GADOVERSETAMIDE|GADOVERSETAMIDE
C3700880|T121|1486818|RXNORM|4,5-DICHLORO-2-OCTYL-3-ISOTHIAZOLONE|4,5-DICHLORO-2-OCTYL-3-ISOTHIAZOLONE
C0205704|T121|66869|RXNORM|CASCARA SAGRADA|CASCARA SAGRADA
C0205704|T121|66869|RXNORM|CASCARA SAGRADA|CASCARA SAGRADA
C3257690|T121|1311648|RXNORM|PANAX GINSENG FRUIT EXTRACT|PANAX GINSENG FRUIT EXTRACT
C1646261|T121|607162|RXNORM|BROMPHENIRAMINE / CARBETAPENTANE / PHENYLEPHRINE|BROMPHENIRAMINE / CARBETAPENTANE / PHENYLEPHRINE
C1656846|T121|607163|RXNORM|BROMPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE|BROMPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE
C3256371|T121|1311643|RXNORM|MORUS NIGRA FRUIT EXTRACT|MORUS NIGRA FRUIT EXTRACT
C3256364|T168|1311642|RXNORM|MORINDA CITRIFOLIA FRUIT JUICE|NONI FRUIT JUICE
C2980817|T109|1311641|RXNORM|MORINDA CITRIFOLIA FRUIT EXTRACT|NONI FRUIT EXTRACT
C1099677|T121|322167|RXNORM|SOLIFENACIN|SOLIFENACIN
C3256991|T121|1311647|RXNORM|ORANGE PEEL WAX|ORANGE PEEL WAX
C3256785|T121|1311646|RXNORM|NARCISSUS TAZETTA BULB EXTRACT|NARCISSUS TAZETTA BULB EXTRACT
C3256374|T121|1311645|RXNORM|MYRCIARIA DUBIA FRUIT EXTRACT|MYRCIARIA DUBIA FRUIT EXTRACT
C2928590|T121|1007674|RXNORM|AMPHOTERICIN B / TRIAMCINOLONE|AMPHOTERICIN B / TRIAMCINOLONE
C2928591|T121|1007675|RXNORM|POTASSIUM TARTRATE / SODIUM BICARBONATE|POTASSIUM TARTRATE / SODIUM BICARBONATE
C2928592|T121|1007676|RXNORM|BARBITAL / PYRILAMINE|BARBITAL / PYRILAMINE
C2928593|T121|1007677|RXNORM|BISMUTH / NAPHAZOLINE|BISMUTH / NAPHAZOLINE
C2928586|T121|1007670|RXNORM|BENZOCAINE / ETHACRIDINE|BENZOCAINE / ETHACRIDINE
C2928587|T121|1007671|RXNORM|CHLORAMPHENICOL / IDOXURIDINE|CHLORAMPHENICOL / IDOXURIDINE
C2928588|T121|1007672|RXNORM|MENTHOL / TROLAMINE SALICYLATE|MENTHOL / TROLAMINE SALICYLATE
C2928589|T121|1007673|RXNORM|LIDOCAINE / MAGNESIUM SULFATE|LIDOCAINE / MAGNESIUM SULFATE
C3643655|T121|1424007|RXNORM|BENZOYL PEROXIDE / SALICYLIC ACID / SULFUR|BENZOYL PEROXIDE / SALICYLIC ACID / SULFUR
C2928594|T121|1007678|RXNORM|DEXPANTHENOL / DIPHENHYDRAMINE / LIDOCAINE|DEXPANTHENOL / DIPHENHYDRAMINE / LIDOCAINE
C2928595|T121|1007679|RXNORM|CAFFEINE / DIPYRONE|CAFFEINE / DIPYRONE
C3256168|T121|1312598|RXNORM|HEXYLDECYL LAURATE|HEXYLDECYL LAURATE
C3486289|T109|1312599|RXNORM|HEXYLDECYL STEARATE|HEXYLDECYL STEARATE
C3505261|T121|1358169|RXNORM|CHROMIUM, CHELATED / MANGANESE GLUCONATE / ZINC CITRATE|CHROMIUM, CHELATED / MANGANESE GLUCONATE / ZINC CITRATE
C0078703|T121|39879|RXNORM|MEPIRODIPINE|BARNIDIPINE
C3666392|T121|1436556|RXNORM|CAFFEINE / CHOLINE|CAFFEINE / CHOLINE
C2080572|T121|820044|RXNORM|BROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLPROPANOLAMINE|BROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLPROPANOLAMINE
C0001157|T131|242|RXNORM|ACONITE|ACONITE
C2194304|T121|812314|RXNORM|FLUNARIZINE / NICERGOLINE|FLUNARIZINE / NICERGOLINE
C0058371|T121|23370|RXNORM|DIPHENIDOL|DIPHENIDOL
C0717693|T121|214492|RXNORM|DEXTROMETHORPHAN / PSEUDOEPHEDRINE|DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C0717692|T121|214491|RXNORM|DEXTROMETHORPHAN / PROMETHAZINE|DEXTROMETHORPHAN / PROMETHAZINE
C0717697|T121|214496|RXNORM|DEXTROMETHORPHAN / PHENYLEPHRINE / PYRILAMINE|DEXTROMETHORPHAN / PHENYLEPHRINE / PYRILAMINE
C0717695|T121|214494|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE|DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE
C0717696|T121|214495|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE|DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE
C0717696|T121|214495|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE|DEXTROMETHORPHAN / GUAIFENESIN / PSEUDOEPHEDRINE
C1874320|T121|689242|RXNORM|ANTIPYRINE / PHENYLEPHRINE|ANTIPYRINE / PHENYLEPHRINE
C3152798|T129|1098130|RXNORM|NARROWLEAF MARSHELDER POLLEN EXTRACT|IVA ANGUSIFOLIA POLLEN EXTRACT
C0084110|T121|1314381|RXNORM|POLYAMINOPROPYL BIGUANIDE|POLYAMINOPROPYL BIGUANIDE
C2947555|T121|1041833|RXNORM|CALCIUM CARBONATE / WHEAT DEXTRIN|CALCIUM CARBONATE / WHEAT DEXTRIN
C2701223|T129|852007|RXNORM|WORMWOOD SAGE POLLEN EXTRACT|ARTEMISIA ABSINTHIUM POLLEN EXTRACT
C3700872|T109|1487142|RXNORM|PEG-60 SORBITAN STEARATE|PEG-60 SORBITAN STEARATE
C3700873|T109|1487140|RXNORM|SALVIA OFFICINALIS ROOT EXTRACT|SALVIA OFFICINALIS ROOT EXTRACT
C3249499|T129|1232604|RXNORM|PALE DOCK POLLEN EXTRACT|RUMEX ALTISSIMUS POLLEN EXTRACT
C0066415|T121|29903|RXNORM|METHYLPARABEN|METHYLPARABEN
C0025010|T129|6669|RXNORM|MEASLES VACCINE|MEASLES VACCINE
C2746114|T129|901631|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 5 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 5 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C2746116|T129|901633|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 6A CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 6A CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C3848573|T196|1546271|RXNORM|NITRATE ION|NITRATE ION
C0110681|T131|1373349|RXNORM|COPPER NAPHTHENATE|COPPER NAPHTHENATE
C0285387|T130|1362135|RXNORM|BASIL OIL|BASIL OIL
C0024977|T121|6664|RXNORM|MAZINDOL|MAZINDOL
C0041213|T130|10878|RXNORM|TRYPAN BLUE|TRYPAN BLUE
C0724635|T197|221125|RXNORM|SODIUM PHOSPHATE,MONOBASIC,MONOHYDRATE|SODIUM PHOSPHATE,MONOBASIC,MONOHYDRATE
C3247831|T121|1193101|RXNORM|FOLIC ACID / OMEGA-3 ACID ETHYL ESTERS (USP) / PHYTOSTEROLS / PYRIDOXINE / VITAMIN B 12|FOLIC ACID / OMEGA-3 ACID ETHYL ESTERS (USP) / PHYTOSTEROLS / PYRIDOXINE / VITAMIN B 12
C0059764|T121|52882|RXNORM|MONOETHYL FUMARATE|MONOETHYL FUMARATE
C0049301|T121|15850|RXNORM|5-METHYL-8-HYDROXYQUINOLINE|5-METHYL-8-HYDROXYQUINOLINE
C1874378|T121|689540|RXNORM|ASPIRIN / PROMETHAZINE / PSEUDOEPHEDRINE|ASPIRIN / PROMETHAZINE / PSEUDOEPHEDRINE
C1874379|T121|689541|RXNORM|ASPIRIN / PROPOXYPHENE|ASPIRIN / PROPOXYPHENE
C0128922|T197|52885|RXNORM|MONOFLUOROPHOSPHATE|MONOFLUOROPHOSPHATE
C0054219|T121|19847|RXNORM|BUMADIZONE|BUMADIZONE
C3848569|T196|1546276|RXNORM|CADMIUM CATION|CADMIUM CATION
C0973231|T197|1546277|RXNORM|BICARBONATE ION|BICARBONATE ION
C1873940|T121|687078|RXNORM|ACETAMINOPHEN / ASPIRIN|ACETAMINOPHEN / ASPIRIN
C0717427|T197|214236|RXNORM|ANHYDROUS CALCIUM IODIDE|ANHYDROUS CALCIUM IODIDE
C0717428|T121|214237|RXNORM|ANHYDROUS CALCIUM IODIDE / CODEINE|ANHYDROUS CALCIUM IODIDE / CODEINE
C0771682|T121|236410|RXNORM|PALMITOYL COLLAGEN ACID|PALMITOYL COLLAGEN ACID
C0717424|T121|214233|RXNORM|AMPICILLIN / PROBENECID|AMPICILLIN / PROBENECID
C0717418|T121|214230|RXNORM|AMOBARBITAL / SECOBARBITAL|AMOBARBITAL / SECOBARBITAL
C3818821|T121|1489545|RXNORM|CINNAMOMUM AROMATICUM WHOLE EXTRACT|CINNAMOMUM AROMATICUM WHOLE EXTRACT
C3474995|T121|1302427|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / GUAIFENESIN|ACETAMINOPHEN / CHLORPHENIRAMINE / GUAIFENESIN
C3486708|T121|1347559|RXNORM|BOWFIN PREPARATION|BOWFIN PREPARATION
C1174995|T129|356988|RXNORM|EFALIZUMAB|EFALIZUMAB
C3818761|T121|1492933|RXNORM|SOPHORA TONKINENSIS WHOLE EXTRACT|SOPHORA TONKINENSIS WHOLE EXTRACT
C3813117|T121|1492935|RXNORM|PARIS QUADRIFOLIA EXTRACT|PARIS QUADRIFOLIA EXTRACT
C3818760|T121|1492934|RXNORM|SALIX ALBA FLOWER EXTRACT|SALIX ALBA FLOWER EXTRACT
C3818759|T121|1492937|RXNORM|LONICERA CONFUSA FLOWER EXTRACT|LONICERA CONFUSA FLOWER EXTRACT
C0443384|T121|124848|RXNORM|DICHLOROTETRAFLUOROETHANE|DICHLOROTETRAFLUOROETHANE
C3812145|T121|1492939|RXNORM|GRINDELIA HIRSUTULA WHOLE EXTRACT|GRINDELIA HIRSUTULA WHOLE EXTRACT
C3818758|T121|1492938|RXNORM|IRIS DOMESTICA WHOLE EXTRACT|IRIS DOMESTICA WHOLE EXTRACT
C0061851|T121|26225|RXNORM|ONDANSETRON|ONDANSETRON
C1443048|T129|465118|RXNORM|TRICHOPHYTON ANTIGEN|TRICHOPHYTON ANTIGEN
C0008221|T121|2372|RXNORM|CHLORMETHIAZOLE|CHLORMETHIAZOLE
C0008223|T121|2373|RXNORM|CHLORMEZANONE|CHLORMEZANONE
C0056727|T121|21945|RXNORM|CYCLOADIPHENINE|CYCLOADIPHENINE
C2701649|T129|852569|RXNORM|BLACK WALNUT POLLEN EXTRACT|JUGLANS NIGRA POLLEN EXTRACT
C3484407|T121|1347557|RXNORM|AMBROSIA ARTEMISIIFOLIA EXTRACT|AMBROSIA ARTEMISIIFOLIA EXTRACT
C2740612|T129|899398|RXNORM|CABBAGE ALLERGENIC EXTRACT|CABBAGE ALLERGENIC EXTRACT
C0055877|T121|21232|RXNORM|CLIDINIUM|CLIDINIUM
C2740609|T129|899394|RXNORM|BUCKWHEAT ALLERGENIC EXTRACT|BUCKWHEAT ALLERGENIC EXTRACT
C0056732|T121|21949|RXNORM|CYCLOBENZAPRINE|CYCLOBENZAPRINE
C2194327|T121|820045|RXNORM|ACETAMINOPHEN / MEPROBAMATE|ACETAMINOPHEN / MEPROBAMATE
C2740796|T129|899738|RXNORM|CUCUMBER ALLERGENIC EXTRACT|CUCUMIS SATIVUS ALLERGENIC EXTRACT
C3254782|T121|1235388|RXNORM|ASCORBIC ACID / FOLIC ACID / NIACIN / RIBOFLAVIN / SODIUM FLUORIDE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN D / VITAMIN E|ASCORBIC ACID / FOLIC ACID / NIACIN / RIBOFLAVIN / SODIUM FLUORIDE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN D / VITAMIN E
C0795616|T121|253171|RXNORM|GOLDEN SEAL ROOT|GOLDEN SEAL ROOT
C1739459|T121|646818|RXNORM|PANGAMATE|PANGAMATE
C2929740|T121|1008842|RXNORM|GLYCERIN / HYPROMELLOSE|GLYCERIN / HYPROMELLOSE
C2929738|T121|1008840|RXNORM|CHROMIUM POLYNICOTINATE / THIOCTATE|CHROMIUM POLYNICOTINATE / THIOCTATE
C1329978|T121|404773|RXNORM|AMLODIPINE / ATORVASTATIN|AMLODIPINE / ATORVASTATIN
C2929744|T121|1008846|RXNORM|DEXTROMETHORPHAN / GUAIACOL|DEXTROMETHORPHAN / GUAIACOL
C2929745|T121|1008847|RXNORM|ARACHIS OIL / CHLOROBUTANOL / DICHLOROBENZENE|CHLOROBUTANOL / DICHLOROBENZENE / PEANUT OIL
C2929742|T121|1008844|RXNORM|RED MULBERRY POLLEN EXTRACT / WHITE MULBERRY POLLEN EXTRACT|RED MULBERRY POLLEN EXTRACT / WHITE MULBERRY POLLEN EXTRACT
C2929743|T121|1008845|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-CALIFORNIA-07-2009 X-181 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-VICTORIA-210-2009 X-187 (H3N2) (A-PERTH-16-2009) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-CALIFORNIA-07-2009 X-181 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-VICTORIA-210-2009 X-187 (H3N2) (A-PERTH-16-2009) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN
C3860186|T109|1594765|RXNORM|PPG-2 HYDROXYETHYL COCAMIDE/ISOSTEARAMIDE|PPG-2 HYDROXYETHYL COCAMIDE/ISOSTEARAMIDE
C3860185|T121|1594764|RXNORM|PAEONIA LACTIFLORA FLOWER EXTRACT|PAEONIA LACTIFLORA FLOWER EXTRACT
C2929746|T121|1008848|RXNORM|CAPSAICIN / MENTHOL / METHYL SALICYLATE|CAPSAICIN / MENTHOL / METHYL SALICYLATE
C2929747|T121|1008849|RXNORM|SALICYLIC ACID / UREA|SALICYLIC ACID / UREA
C3834089|T122|1541725|RXNORM|GARDENIA RESINIFERA RESIN|GARDENIA RESINIFERA RESIN
C0007299|T121|2116|RXNORM|CARTEOLOL|CARTEOLOL
C0007299|T121|2116|RXNORM|CARTEOLOL|CARTEOLOL
C2927921|T121|1006998|RXNORM|ACETAMINOPHEN / ASTEMIZOLE / PHENYLEPHRINE|ACETAMINOPHEN / ASTEMIZOLE / PHENYLEPHRINE
C2927922|T121|1006999|RXNORM|DODECYL SULFATE / ZINC PYRITHIONE|DODECYL SULFATE / ZINC PYRITHIONE
C2927919|T121|1006996|RXNORM|ESTROGENS, CONJUGATED (USP) / MEDROGESTONE|ESTROGENS, CONJUGATED (USP) / MEDROGESTONE
C2927920|T121|1006997|RXNORM|BENZOCAINE / SALICYLIC ACID|BENZOCAINE / SALICYLIC ACID
C2927917|T121|1006994|RXNORM|PIRETANIDE / RAMIPRIL|PIRETANIDE / RAMIPRIL
C2927918|T121|1006995|RXNORM|ALUMINUM HYDROXIDE / ASPIRIN / CAFFEINE|ALUMINUM HYDROXIDE / ASPIRIN / CAFFEINE
C2927915|T121|1006992|RXNORM|MERBROMIN / PENICILLIN G|MERBROMIN / PENICILLIN G
C2927916|T121|1006993|RXNORM|NIACINAMIDE / QUININE / THIAMINE|NIACINAMIDE / QUININE / THIAMINE
C2927913|T121|1006990|RXNORM|BENZALKONIUM / PANTOTHENIC ACID|BENZALKONIUM / PANTOTHENIC ACID
C2927914|T121|1006991|RXNORM|HYDROCORTISONE / NATAMYCIN / NEOMYCIN|HYDROCORTISONE / NATAMYCIN / NEOMYCIN
C0006711|T197|1919|RXNORM|CALCIUM PHOSPHATE|CALCIUM PHOSPHATE
C1012255|T204|1368365|RXNORM|TRICHINELLA BRITOVI|TRICHINELLA BRITOVI
C3489040|T121|1368361|RXNORM|SOLANUM LYCOPERSICUM EXTRACT|SOLANUM LYCOPERSICUM EXTRACT
C0011816|T121|3289|RXNORM|DEXTROMETHORPHAN|DEXTROMETHORPHAN
C0011812|T121|3288|RXNORM|DEXTROAMPHETAMINE|DEXTROAMPHETAMINE
C1875427|T121|690733|RXNORM|LANOLIN / MINERAL OIL|LANOLIN / MINERAL OIL
C0006701|T197|1910|RXNORM|CALCIUM HYDROXIDE|CALCIUM HYDROXIDE
C3247211|T121|1191504|RXNORM|BUPIVACAINE LIPOSOME|BUPIVACAINE LIPOSOME
C3714579|T121|1541720|RXNORM|LAURUS NOBILIS WHOLE EXTRACT|LAURUS NOBILIS WHOLE EXTRACT
C0081913|T121|158660|RXNORM|PROXIGERMANIUM|PROXIGERMANIUM
C3488429|T109|1309747|RXNORM|CERVUS ELAPHUS HORN OIL|CERVUS ELAPHUS HORN OIL
C3488275|T121|1309746|RXNORM|THUJA PLICATA LEAF EXTRACT|THUJA PLICATA LEAF EXTRACT
C3488274|T121|1309745|RXNORM|ROSA CANINA FLOWER EXTRACT|ROSA CANINA FLOWER EXTRACT
C0076313|T109|1363713|RXNORM|TETRAMETHYLTHIURAM MONOSULFIDE|TETRAMETHYLTHIURAM MONOSULFIDE
C3488273|T121|1309743|RXNORM|MALUS SYLVESTRIS FLOWER EXTRACT|MALUS SYLVESTRIS FLOWER EXTRACT
C0117000|T109|1363715|RXNORM|EUTANOL G|EUTANOL G
C0070559|T121|1309741|RXNORM|PHENETHYLAMINE|PHENETHYLAMINE
C0283192|T109|1363717|RXNORM|ISOMALT|ISOMALT
C0052884|T195|1363718|RXNORM|BACITRACIN METHYLENE DISALICYLATE|BACITRACIN METHYLENE DISALICYLATE
C0521891|T195|1363719|RXNORM|TYLOSIN PHOSPHATE|TYLOSIN PHOSPHATE
C1875136|T121|692993|RXNORM|ETHINYL ESTRADIOL / FLUOXYMESTERONE|ETHINYL ESTRADIOL / FLUOXYMESTERONE
C3488290|T121|1309748|RXNORM|CLEMATIS VITALBA TOP EXTRACT|CLEMATIS VITALBA PRE-FLOWERING TOP EXTRACT
C0076341|T121|37985|RXNORM|TETRAZEPAM|TETRAZEPAM
C3854003|T121|1594763|RXNORM|FERULA COMMUNIS SUBSP. GLAUCA EXTRACT|FERULA COMMUNIS SUBSP. GLAUCA EXTRACT
C0039936|T121|10498|RXNORM|THIOPROPERAZINE|THIOPROPERAZINE
C0039925|T121|10493|RXNORM|THIOPENTAL|THIOPENTAL
C3256373|T126|1314198|RXNORM|MUTANASE SCHIZOSACCHAROMYCES POMBE|MUTANASE SCHIZOSACCHAROMYCES POMBE
C3256431|T109|1314199|RXNORM|PIPER METHYSTICUM WHOLE EXTRACT|PIPER METHYSTICUM WHOLE EXTRACT
C3527637|T121|1360623|RXNORM|PLATYCLADUS ORIENTALIS POLLEN EXTRACT|PLATYCLADUS ORIENTALIS POLLEN EXTRACT
C3527636|T121|1360622|RXNORM|ECLIPTA PROSTRATA WHOLE EXTRACT|ECLIPTA PROSTRATA WHOLE EXTRACT
C3527639|T121|1360625|RXNORM|TRIPTERYGIUM WILFORDII ROOT EXTRACT|TRIPTERYGIUM WILFORDII ROOT EXTRACT
C3527638|T121|1360624|RXNORM|SANGUISORBA OFFICINALIS LEAF EXTRACT|SANGUISORBA OFFICINALIS LEAF EXTRACT
C3527641|T109|1360627|RXNORM|PINE NEEDLE OIL (PINUS MUGO)|PINE NEEDLE OIL (PINUS MUGO)
C3527640|T121|1360626|RXNORM|(ALL-Z)-4,7,10,13,16-DOCOSAPENTAENOIC ACID,|(ALL-Z)-4,7,10,13,16-DOCOSAPENTAENOIC ACID,
C3256066|T121|1314190|RXNORM|PEG-20 SOY STEROL|PEG-20 SOY STEROL
C3256068|T121|1314191|RXNORM|PEG-200 DILAURATE|PEG-200 DILAURATE
C3256069|T121|1314192|RXNORM|PEG-25 PROPYLENE GLYCOL STEARATE|PEG-25 PROPYLENE GLYCOL STEARATE
C3256076|T121|1314193|RXNORM|PEG-6 METHYL ETHER|PEG-6 METHYL ETHER
C3256080|T121|1314194|RXNORM|PEG-8 DIMETHICONE|PEG-8 DIMETHICONE
C2825348|T129|1314195|RXNORM|IMMUNOGLOBULIN M, HUMAN|IMMUNOGLOBULIN M, HUMAN
C3256179|T121|1314196|RXNORM|PENTAERYTHRITYL TETRAOLEATE|PENTAERYTHRITYL TETRAOLEATE
C3256249|T121|1314197|RXNORM|PHELLINUS LINTEUS WHOLE EXTRACT|PHELLINUS LINTEUS WHOLE EXTRACT
C3651952|T121|1428952|RXNORM|ALPHA HYDROXY ACIDS / UREA|ALPHA HYDROXY ACIDS / UREA
C0054409|T123|20012|RXNORM|CADEXOMER IODINE|CADEXOMER IODINE
C2146627|T121|814486|RXNORM|ACETAMINOPHEN / PROMETHAZINE|ACETAMINOPHEN / PROMETHAZINE
C3667076|T121|1438492|RXNORM|HEXADECANOLACTONE|HEXADECANOLACTONE
C2726211|T129|974687|RXNORM|RADISH ALLERGENIC EXTRACT|RAPHANUS SATIVUS EXTRACT
C0874041|T121|260014|RXNORM|WATERMELON PREPARATION|WATERMELON PREPARATION
C2927178|T121|1002293|RXNORM|FORMOTEROL / MOMETASONE|FORMOTEROL / MOMETASONE
C1718383|T121|1310520|RXNORM|TERIFLUNOMIDE|TERIFLUNOMIDE
C0874039|T121|260012|RXNORM|SALICIN EXTRACT|SALICIN EXTRACT
C0982246|T121|1364294|RXNORM|ACETYLATED LANOLIN ALCOHOLS|ACETYLATED LANOLIN ALCOHOLS
C1095904|T121|1364295|RXNORM|CLOVE PREPARATION|CLOVE PREPARATION
C3257525|T121|1358901|RXNORM|KIWI FRUIT EXTRACT|KIWI FRUIT EXTRACT
C3256646|T121|1358900|RXNORM|PONCIRUS TRIFOLIATA FRUIT EXTRACT|PONCIRUS TRIFOLIATA FRUIT EXTRACT
C1698893|T130|1364290|RXNORM|GADOFOSVESET|GADOFOSVESET
C0939864|T168|1364291|RXNORM|LEMON EXTRACT|LEMON EXTRACT
C0939919|T121|1364292|RXNORM|LOBELIA INFLATA PREPARATION|LOBELIA INFLATA PREPARATION
C0982088|T121|1364293|RXNORM|COCO-CAPRYLATE|COCO-CAPRYLATE
C0292819|T121|85763|RXNORM|FOMIVIRSEN|FOMIVIRSEN
C0292818|T121|85762|RXNORM|RITONAVIR|RITONAVIR
C0092801|T121|44157|RXNORM|CLADRIBINE|CLADRIBINE
C3190695|T121|1145020|RXNORM|ALLANTOIN / CHLOROXYLENOL|ALLANTOIN / CHLOROXYLENOL
C0092777|T121|44151|RXNORM|CLOFARABINE|CLOFARABINE
C2073836|T121|1144260|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / SALICYLAMIDE|ACETAMINOPHEN / CHLORPHENIRAMINE / SALICYLAMIDE
C0037517|T197|9880|RXNORM|SODIUM HYDROXIDE|SODIUM HYDROXIDE
C3163606|T121|1116741|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-CHRISTCHURCH-16-2010 NIB-74 (H1N1) (A-CALIFORNIA-7-2009) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-VICTORIA-210-2009 X-187 (H3N2) (A-PERTH-16-2009) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-CHRISTCHURCH-16-2010 NIB-74 (H1N1) (A-CALIFORNIA-7-2009) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-VICTORIA-210-2009 X-187 (H3N2) (A-PERTH-16-2009) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN
C2927992|T121|1007069|RXNORM|DIBUNATE / GUAIFENESIN|DIBUNATE / GUAIFENESIN
C2927991|T121|1007068|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL / MAGNESIUM OXIDE|CALCIUM CARBONATE / CHOLECALCIFEROL / MAGNESIUM OXIDE
C0056244|T121|1309334|RXNORM|CONIFERYL ALCOHOL|CONIFERYL ALCOHOL
C3488608|T109|1309332|RXNORM|MATRICARIA CHAMOMILLA FLOWERING TOP OIL|MATRICARIA CHAMOMILLA FLOWERING TOP OIL
C3488929|T121|1309330|RXNORM|MELALEUCA ALTERNIFOLIA LEAF EXTRACT|MELALEUCA ALTERNIFOLIA LEAF EXTRACT
C3488963|T109|1309331|RXNORM|CUPRESSUS SEMPERVIRENS LEAF OIL|CUPRESSUS SEMPERVIRENS LEAF OIL
C2927984|T121|1007061|RXNORM|DIMETHICONE / METHYLNICOTINATE|DIMETHICONE / METHYLNICOTINATE
C2927983|T121|1007060|RXNORM|BUCLIZINE / HYDROXYZINE / NIACIN|BUCLIZINE / HYDROXYZINE / NIACIN
C2927986|T121|1007063|RXNORM|CALCIUM ASPARTATE / MAGNESIUM SALT / POTASSIUM ASPARTATE|CALCIUM ASPARTATE / MAGNESIUM SALT / POTASSIUM ASPARTATE
C2927985|T121|1007062|RXNORM|GINKGO BILOBA EXTRACT / GLUTAMINE|GINKGO BILOBA EXTRACT / GLUTAMINE
C0025696|T121|6860|RXNORM|METHYCLOTHIAZIDE|METHYCLOTHIAZIDE
C2927987|T121|1007064|RXNORM|GLYCERIN / HYPROMELLOSE / POLYETHYLENE GLYCOL 400|GLYCERIN / HYPROMELLOSE / POLYETHYLENE GLYCOL 400
C2927990|T121|1007067|RXNORM|CRANBERRY PREPARATION / OLIVE LEAF EXTRACT|CRANBERRY PREPARATION / OLIVE LEAF EXTRACT
C1874793|T121|689301|RXNORM|CHLOROPHYLLIN COPPER COMPLEX / SODIUM CHLORIDE|CHLOROPHYLLIN COPPER COMPLEX / SODIUM CHLORIDE
C1874794|T121|689302|RXNORM|CHLOROPHYLLIN COPPER COMPLEX / SODIUM PROPIONATE|CHLOROPHYLLIN COPPER COMPLEX / SODIUM PROPIONATE
C1874795|T121|689303|RXNORM|CHLOROQUINE / PRIMAQUINE|CHLOROQUINE / PRIMAQUINE
C1875164|T121|689304|RXNORM|FLUOROMETHOLONE / SULFACETAMIDE|FLUOROMETHOLONE / SULFACETAMIDE
C0360172|T121|107770|RXNORM|MEPENZOLATE|MEPENZOLATE
C0360174|T121|107771|RXNORM|DEMECARIUM|DEMECARIUM
C3204554|T129|1119986|RXNORM|CENTRUROIDES (SCORPION) IMMUNE F(AB')2 (EQUINE)|CENTRUROIDES (SCORPION) IMMUNE F(AB')2 (EQUINE)
C1321984|T121|402565|RXNORM|DIBUNATE|DIBUNATE
C3486832|T121|1311346|RXNORM|SUS SCROFA SUPERIOR GASTRIC PLEXUS PREPARATION|PORCINE SUPERIOR GASTRIC PLEXUS PREPARATION
C3486831|T121|1311344|RXNORM|SUS SCROFA SPLEEN PREPARATION|PORCINE SPLEEN PREPARATION
C1714166|T121|636827|RXNORM|GUAIACOLSULFONATE|GUAIACOLSULFONATE
C3486830|T121|1311343|RXNORM|SUS SCROFA RECTUM PREPARATION|PORCINE RECTUM PREPARATION
C3486828|T121|1311340|RXNORM|SUS SCROFA PROSTATE PREPARATION|PORCINE PROSTATE PREPARATION
C3486829|T121|1311341|RXNORM|SUS SCROFA PYLORUS PREPARATION|PORCINE PYLORUS PREPARATION
C0981971|T129|314455|RXNORM|SILK ALLERGENIC EXTRACT|BOMBYX MORI FIBER ALLERGENIC EXTRACT
C3486843|T121|1311349|RXNORM|SUS SCROFA TESTICLE PREPARATION|PORCINE TESTICLE PREPARATION
C2928166|T121|1007244|RXNORM|TALC / ZINC OXIDE|TALC / ZINC OXIDE
C2928169|T121|1007247|RXNORM|CHLOROXYLENOL / UNDECYLENATE|CHLOROXYLENOL / UNDECYLENATE
C2928169|T121|1007247|RXNORM|CHLOROXYLENOL / UNDECYLENATE|CHLOROXYLENOL / UNDECYLENATE
C2928168|T121|1007246|RXNORM|COBAMAMIDE / FOLIC ACID|COBAMAMIDE / FOLIC ACID
C2928163|T121|1007241|RXNORM|ACEXAMIC ACID / CETRIMONIUM|ACEXAMIC ACID / CETRIMONIUM
C2928162|T121|1007240|RXNORM|ACETIAMINE / ASPIRIN|ACETIAMINE / ASPIRIN
C2928164|T121|1007242|RXNORM|COBAMAMIDE / CYPROHEPTADINE|COBAMAMIDE / CYPROHEPTADINE
C3256850|T109|1368363|RXNORM|LAURYL PYRROLIDONE|LAURYL PYRROLIDONE
C2928171|T121|1007249|RXNORM|FRUCTOOLIGOSACCHARIDE / LACTOBACILLUS ACIDOPHILUS|FRUCTOOLIGOSACCHARIDE / LACTOBACILLUS ACIDOPHILUS
C0004499|T195|1266|RXNORM|AZLOCILLIN|AZLOCILLIN
C0244404|T121|72143|RXNORM|RALOXIFENE|RALOXIFENE
C0255289|T129|76469|RXNORM|BCG, LIVE, CONNAUGHT STRAIN|BCG, LIVE, CONNAUGHT STRAIN
C0033488|T123|8783|RXNORM|PROPOLIS|PROPOLIS
C0033487|T121|8782|RXNORM|PROPOFOL|PROPOFOL
C0033497|T121|8787|RXNORM|PROPRANOLOL|PROPRANOLOL
C0033493|T121|8785|RXNORM|PROPOXYPHENE|PROPOXYPHENE
C0030840|T195|7984|RXNORM|HEPATITIS B SURFACE ANTIGEN (AUSTRALIA ANTIGEN) MSD, VACCINE|PENICILLIN V
C1117793|T121|325518|RXNORM|TRIMETHOXYBENZENE|TRIMETHOXYBENZENE
C1117888|T121|325519|RXNORM|POTASSIUM ESTRONE|POTASSIUM ESTRONE
C0078168|T121|39468|RXNORM|VERALIPRIDE|VERALIPRIDE
C1875431|T121|690737|RXNORM|LANOLIN / MINERAL OIL / PETROLATUM|LANOLIN / MINERAL OIL / PETROLATUM
C0028833|T125|7617|RXNORM|OCTREOTIDE|OCTREOTIDE
C1116570|T121|325514|RXNORM|INDIGOTINDISULFONATE|INDIGOTINDISULFONATE
C3255688|T121|1311551|RXNORM|LILIUM CANDIDUM BULB EXTRACT|LILIUM CANDIDUM BULB EXTRACT
C0011707|T125|3255|RXNORM|PETROLATUM DISTILLATES|DESOXIMETASONE
C1117748|T121|325517|RXNORM|PHENYLEHRINE|PHENYLEHRINE
C3488644|T121|1311122|RXNORM|TRITICUM AESTIVUM EXTRACT|TRITICUM AESTIVUM EXTRACT
C0378482|T121|114979|RXNORM|RABEPRAZOLE|RABEPRAZOLE
C3267232|T121|1314336|RXNORM|C13-15 ALKANE|C13-15 ALKANE
C3486719|T121|1311121|RXNORM|PSEUDOGNAPHALIUM OBTUSIFOLIUM EXTRACT|PSEUDOGNAPHALIUM OBTUSIFOLIUM EXTRACT
C0001455|T123|1314330|RXNORM|CYCLIC AMP|CYCLIC AMP
C3256096|T121|1311127|RXNORM|ASCOPHYLLUM NODOSUM EXTRACT|ASCOPHYLLUM NODOSUM EXTRACT
C3256345|T109|1314332|RXNORM|BAMBUSA VULGARIS TOP EXTRACT|BAMBUSA VULGARIS TOP EXTRACT
C3489052|T121|1311125|RXNORM|MYRTUS COMMUNIS TOP EXTRACT|MYRTUS COMMUNIS TOP EXTRACT
C0378466|T121|114970|RXNORM|ZAFIRLUKAST|ZAFIRLUKAST
C0132768|T109|1314253|RXNORM|NONANAL|NONANAL
C3489053|T121|1311128|RXNORM|CITHARACANTHUS SPINICRUS PREPARATION|CITHARACANTHUS SPINICRUS PREPARATION
C3489117|T204|1311129|RXNORM|YEAST MANNAN PREPARATION|YEAST MANNAN PREPARATION
C0006947|T131|1314339|RXNORM|CARBADOX|CARBADOX
C3709596|T121|1487829|RXNORM|CINNAMOMUM CAMPHORA WHOLE EXTRACT|CINNAMOMUM CAMPHORA WHOLE EXTRACT
C0068065|T121|1363710|RXNORM|N-ISOPROPYL-N-PHENYL-4-PHENYLENEDIAMINE|N-ISOPROPYL-N-PHENYL-4-PHENYLENEDIAMINE
C0071568|T126|34132|RXNORM|PEGASPARGASE|PEGASPARGASE
C3472777|T121|1314251|RXNORM|POVIDONE K15|POVIDONE K15
C0938417|T121|284110|RXNORM|FE HEME POLYPEPTIDE|FE HEME POLYPEPTIDE
C0068253|T131|1363711|RXNORM|N-OXYDIETHYLENE-2-BENZOTHIAZOLE SULFENAMIDE|N-OXYDIETHYLENE-2-BENZOTHIAZOLE SULFENAMIDE
C0072176|T195|34649|RXNORM|PROPICILLIN|PROPICILLIN
C3256454|T121|1314250|RXNORM|TRIMETHYLSILANE|TRIMETHYLSILANE
C0069936|T121|1363712|RXNORM|PADIMATE A|PADIMATE A
C3709594|T121|1487827|RXNORM|CANARIUM LUZONICUM WHOLE EXTRACT|CANARIUM LUZONICUM WHOLE EXTRACT
C0044551|T109|1487826|RXNORM|1-OCTANOL|1-OCTANOL
C1276848|T121|883815|RXNORM|DEXAMETHASONE / TOBRAMYCIN|DEXAMETHASONE / TOBRAMYCIN
C0033382|T123|8737|RXNORM|PROLINE|PROLINE
C0083735|T123|1363714|RXNORM|NEUROTROPHIN 3|NEUROTROPHIN 3
C3692372|T121|1441830|RXNORM|DOXYLAMINE / PHENYLEPHRINE|DOXYLAMINE / PHENYLEPHRINE
C1719977|T121|729578|RXNORM|ISOPROPYL MYRISTATE / MINERAL OIL|ISOPROPYL MYRISTATE / MINERAL OIL
C0162753|T130|1363716|RXNORM|SAFFRON STAIN|SAFFRON STAIN
C0620168|T130|1552361|RXNORM|2,6-DIMETHYL-5-HEPTENAL|2,6-DIMETHYL-5-HEPTENAL
C0071780|T197|34323|RXNORM|POTASSIUM SULFATE|POTASSIUM SULFATE
C0961649|T121|298983|RXNORM|PONAZURIL|PONAZURIL
C2700232|T196|1546282|RXNORM|GALLIUM CATION|GALLIUM CATION
C0301704|T109|89959|RXNORM|PHOSPHATIDYLSERINE|PHOSPHATIDYLSERINE
C0058133|T121|23161|RXNORM|ALDIOXA|ALDIOXA
C0058135|T121|23163|RXNORM|DIHYDROXYALUMINUM SODIUM CARBONATE|DIHYDROXYALUMINUM SODIUM CARBONATE
C1519169|T121|496653|RXNORM|SALICYLIC ACID / SULFUR|SALICYLIC ACID / SULFUR
C1519169|T121|496653|RXNORM|SALICYLIC ACID / SULFUR|SALICYLIC ACID / SULFUR
C0108143|T122|47633|RXNORM|CALCIUM STEARATE|CALCIUM STEARATE
C0108139|T121|47630|RXNORM|CALCIUM POLYSTYRENE SULFONATE PRODUCT|CALCIUM POLYSTYRENE SULFONATE PRODUCT
C3818793|T121|1490797|RXNORM|FERROUS CYSTEINE GLYCINATE|FERROUS CYSTEINE GLYCINATE
C0001026|T123|1490796|RXNORM|ACETYL COENZYME A|ACETYL COENZYME A
C0301508|T129|89890|RXNORM|YELLOW FEVER VACCINE|YELLOW FEVER, LIVE ATTENUATED
C3819182|T121|1490790|RXNORM|CAMPHOR / LEVOMENTHOL|CAMPHOR / LEVOMENTHOL
C0032483|T122|8516|RXNORM|POLYETHYLENE GLYCOLS|POLYETHYLENE GLYCOLS
C2106233|T121|813232|RXNORM|CHLOROXYLENOL / COAL TAR|CHLOROXYLENOL / COAL TAR
C3857948|T121|1552360|RXNORM|PEG-200 HYDROGENATED GLYCERYL PALMATE|PEG-200 HYDROGENATED GLYCERYL PALMATE
C0054668|T121|20217|RXNORM|CARBETAPENTANE|PENTOXYVERINE
C0030969|T121|8042|RXNORM|PERAZINE|PERAZINE
C0062092|T121|26412|RXNORM|HALAZEPAM|HALAZEPAM
C2731409|T109|895223|RXNORM|ACACIA BAILEYANA POLLEN EXTRACT|ACACIA BAILEYANA POLLEN EXTRACT
C0062097|T121|26416|RXNORM|HALOMETASONE|HALOMETASONE
C3488311|T121|1309749|RXNORM|CALLUNA VULGARIS FLOWERING TOP EXTRACT|CALLUNA VULGARIS FLOWERING TOP EXTRACT
C2974521|T121|1537034|RXNORM|VORAPAXAR|VORAPAXAR
C2980882|T121|1094114|RXNORM|ECHINACEA ANGUSTIFOLIA ROOT EXTRACT / ECHINACEA PURPUREA ROOT EXTRACT|ECHINACEA ANGUSTIFOLIA ROOT EXTRACT / ECHINACEA PURPUREA ROOT EXTRACT
C0015025|T125|4129|RXNORM|ETHISTERONE|ETHISTERONE
C0376637|T121|114289|RXNORM|INDINAVIR|INDINAVIR
C1145579|T121|342940|RXNORM|PAU D'ARCO PREPARATION|PAU D'ARCO PREPARATION
C0015021|T121|4127|RXNORM|ETHIONAMIDE|ETHIONAMIDE
C0015020|T121|4126|RXNORM|AMIFOSTINE|AMIFOSTINE
C0015018|T130|4125|RXNORM|ETHIODIZED OIL|ETHIODIZED OIL
C0015011|T125|4124|RXNORM|ETHINYL ESTRADIOL|ETHINYL ESTRADIOL
C2183094|T121|815192|RXNORM|CITRIC ACID / DEXTROMETHORPHAN / GUAIFENESIN / POTASSIUM CITRATE|CITRIC ACID / DEXTROMETHORPHAN / GUAIFENESIN / POTASSIUM CITRATE
C2701770|T129|852742|RXNORM|ENGLISH PLANTAIN POLLEN EXTRACT|PLANTAGO LANCEOLATA POLLEN EXTRACT
C1108725|T121|324003|RXNORM|BISMUTH DIPROPYLACETATE|BISMUTH DIPROPYLACETATE
C2701415|T129|852217|RXNORM|SMOOTH BROME POLLEN EXTRACT|BROMUS INERMIX POLLEN EXTRACT
C1109120|T121|324005|RXNORM|D-TRANSALLETHRIN|D-TRANSALLETHRIN
C2940200|T129|1014755|RXNORM|WESTERN BLACK WILLOW POLLEN EXTRACT|SALIX LUCIDA SSP. LASIANDRA POLLEN EXTRACT
C0728888|T007|1544929|RXNORM|ENTEROBACTER AEROGENES|ENTEROBACTER AEROGENES
C0254119|T129|75917|RXNORM|INTERFERON BETA-1A|INTERFERON BETA-1A
C2073897|T121|818485|RXNORM|CHLORPHENIRAMINE / GUAIFENESIN / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PYRILAMINE|CHLORPHENIRAMINE / GUAIFENESIN / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PYRILAMINE
C3256082|T121|1313258|RXNORM|PEG-8 RICINOLEATE|PEG-8 RICINOLEATE
C0628659|T109|1313259|RXNORM|TOCOPHERYL RETINOATE|TOCOPHERYL RETINOATE
C3255968|T121|1313256|RXNORM|PEG-12 LAURATE|PEG-12 LAURATE
C3255969|T121|1313257|RXNORM|PEG-12 STEARATE|PEG-12 STEARATE
C3256382|T109|1426365|RXNORM|TRIDECETH-6|TRIDECETH-6
C3257533|T109|1426364|RXNORM|TANGERINE EXTRACT|TANGERINE EXTRACT
C2603645|T109|1426360|RXNORM|STEARYL STEARATE|STEARYL STEARATE
C2929036|T121|1008129|RXNORM|DIAZEPAM / HYOSCYAMINE|DIAZEPAM / HYOSCYAMINE
C2929035|T121|1008128|RXNORM|ATROPINE / HYOSCYAMINE / METHENAMINE / PHENYL SALICYLATE|ATROPINE / HYOSCYAMINE / METHENAMINE / PHENYL SALICYLATE
C2194256|T121|815995|RXNORM|ETHINYL ESTRADIOL / METHYLTESTOSTERONE|ETHINYL ESTRADIOL / METHYLTESTOSTERONE
C2075682|T121|815990|RXNORM|BROMAZEPAM / CLEBOPRIDE / SIMETHICONE|BROMAZEPAM / CLEBOPRIDE / SIMETHICONE
C2929028|T121|1008121|RXNORM|DIFLUCORTOLONE / ISOCONAZOLE|DIFLUCORTOLONE / ISOCONAZOLE
C2929027|T121|1008120|RXNORM|PYRIDOXAL / TYROSINE|PYRIDOXAL / TYROSINE
C2929030|T121|1008123|RXNORM|BORIC ACID / PHENYLEPHRINE|BORIC ACID / PHENYLEPHRINE
C0043668|T127|11516|RXNORM|DOXERCALCIFEROL|DOXERCALCIFEROL
C2929032|T121|1008125|RXNORM|DIPYRONE / HOMATROPINE|DIPYRONE / HOMATROPINE
C2929031|T121|1008124|RXNORM|ACETAMINOPHEN / CALCIUM CARBONATE / MAGNESIUM CARBONATE / MAGNESIUM OXIDE|ACETAMINOPHEN / CALCIUM CARBONATE / MAGNESIUM CARBONATE / MAGNESIUM OXIDE
C2929034|T121|1008127|RXNORM|CETRIMIDES / CHLORHEXIDINE|CETRIMIDES / CHLORHEXIDINE
C0022057|T121|5979|RXNORM|IPRINDOLE|IPRINDOLE
C0022038|T130|5973|RXNORM|IOXAGLATE|IOXAGLATE
C2726167|T129|968426|RXNORM|TRICHOTHECIUM ROSEUM EXTRACT|TRICHOTHECIUM ROSEUM EXTRACT
C0022049|T130|5976|RXNORM|IPODATE|IPODATE
C0022046|T121|5975|RXNORM|IPECAC|IPECACUANHA
C2726166|T129|968422|RXNORM|TRICHOPHYTON SCHOENLEINII ALLERGENIC EXTRACT|TRICHOPHYTON SCHOENLEINII ALLERGENIC EXTRACT
C3255929|T109|1368179|RXNORM|DI-C12-15 ALKYL FUMARATE|DI-C12-15 ALKYL FUMARATE
C0026941|T007|1360621|RXNORM|MYCOPLASMA PNEUMONIAE|MYCOPLASMA PNEUMONIAE
C0058470|T130|1368171|RXNORM|DISPERSE BLUE 106|DISPERSE BLUE 106
C0058383|T109|1368170|RXNORM|DIPHENYLGUANIDINE|DIPHENYLGUANIDINE
C0068450|T121|1368173|RXNORM|NARINGENIN|NARINGENIN
C0063914|T130|1368172|RXNORM|ISOAMYL ACETATE|ISOAMYL ACETATE
C0072229|T109|1368175|RXNORM|PROPYLENE OXIDE|PROPYLENE OXIDE
C0070686|T121|1368174|RXNORM|PHENYLISOTHIOCYANATE|PHENYLISOTHIOCYANATE
C0078260|T130|1368177|RXNORM|VINYL ACETATE|VINYL ACETATE
C0078032|T121|1368176|RXNORM|VANILLIN|VANILLIN
C0293969|T125|1492039|RXNORM|PRALMORELIN|PRALMORELIN
C0060405|T195|25037|RXNORM|CEFDINIR|CEFDINIR
C3818779|T109|1492035|RXNORM|CAPRYLOYL SALICYLIC ACID|CAPRYLOYL SALICYLIC ACID
C0060400|T195|25033|RXNORM|CEFIXIME|CEFIXIME
C3818777|T109|1492037|RXNORM|GENIPA AMERICANA FRUIT EXTRACT|GENIPA AMERICANA FRUIT EXTRACT
C1875139|T121|693000|RXNORM|ETHYNODIOL / MESTRANOL|ETHYNODIOL / MESTRANOL
C0217385|T130|69893|RXNORM|PENTETREOTIDE|PENTETREOTIDE
C1617275|T121|579893|RXNORM|CORNSILK|CORNSILK
C3527643|T121|1360629|RXNORM|ZANTHOXYLUM BUNGEANUM FRUIT EXTRACT|ZANTHOXYLUM BUNGEANUM FRUIT EXTRACT
C2701762|T129|905258|RXNORM|AMERICAN COCKROACH ALLERGENIC EXTRACT|PERIPLANETA AMERICANA ALLERGENIC EXTRACT
C3464315|T121|1307598|RXNORM|GLYCYRRHIZA INFLATA ROOT EXTRACT|GLYCYRRHIZA INFLATA ROOT EXTRACT
C3256173|T121|1307599|RXNORM|PELARGONIUM GRAVEOLENS FLOWERING TOP EXTRACT|PELARGONIUM GRAVEOLENS FLOWERING TOP EXTRACT
C3527642|T121|1360628|RXNORM|RUMEX CRISPUS WHOLE EXTRACT|RUMEX CRISPUS WHOLE EXTRACT
C3256350|T121|1307594|RXNORM|CEDRUS ATLANTICA BARK EXTRACT|CEDRUS ATLANTICA BARK EXTRACT
C3257766|T121|1307595|RXNORM|COLA ACUMINATA SEED EXTRACT|COLA ACUMINATA SEED EXTRACT
C2348464|T121|1307596|RXNORM|EQUISETUM ARVENSE BRANCH EXTRACT|EQUISETUM ARVENSE BRANCH EXTRACT
C3256733|T121|1307597|RXNORM|SELENICEREUS GRANDIFLORUS FLOWER EXTRACT|SELENICEREUS GRANDIFLORUS FLOWER EXTRACT
C3256755|T121|1307590|RXNORM|CAPER BERRY EXTRACT|CAPER BERRY EXTRACT
C3255696|T121|1307591|RXNORM|LONICERA DASYSTYLA FLOWER BUD EXTRACT|LONICERA DASYSTYLA FLOWER BUD EXTRACT
C3256594|T109|1307592|RXNORM|AJUGA TURKESTANICA TOP EXTRACT|AJUGA TURKESTANICA TOP EXTRACT
C2699491|T121|1307593|RXNORM|SOPHORA FLAVESCENS ROOT EXTRACT|SOPHORA FLAVESCENS ROOT EXTRACT
C0213771|T121|69120|RXNORM|TIOTROPIUM|TIOTROPIUM
C0008947|T195|2582|RXNORM|CLINDAMYCIN|CLINDAMYCIN
C0008947|T195|2582|RXNORM|CLINDAMYCIN|CLINDAMYCIN
C0008947|T195|2582|RXNORM|CLINDAMYCIN|CLINDAMYCIN
C0008932|T121|2580|RXNORM|CLENBUTEROL|CLENBUTEROL
C3486602|T121|1322548|RXNORM|CHAMAELIRIUM LUTEUM ROOT EXTRACT|CHAMAELIRIUM LUTEUM ROOT EXTRACT
C0043125|T005|1316080|RXNORM|WEST NILE VIRUS|WEST NILE VIRUS
C3486653|T129|1322549|RXNORM|BACILLUS ANTHRACIS IMMUNOSERUM RABBIT|BACILLUS ANTHRACIS IMMUNOSERUM RABBIT
C0052300|T168|18235|RXNORM|ARACHIS OIL|GROUNDNUT OIL
C0060657|T121|25255|RXNORM|FORMOTEROL|FORMOTEROL
C2742797|T129|1538097|RXNORM|VEDOLIZUMAB|VEDOLIZUMAB
C2928696|T121|1007781|RXNORM|DOCOSAHEXAENOATE / PHOSPHOLIPIDS|DOCOSAHEXAENOATE / PHOSPHOLIPIDS
C2728172|T129|972689|RXNORM|BEEF LIVER ALLERGENIC EXTRACT|BEEF LIVER ALLERGENIC EXTRACT
C0963398|T121|300195|RXNORM|TENOFOVIR DISOPROXIL|TENOFOVIR DISOPROXIL
C3486791|T121|1347560|RXNORM|MAHONIA AQUIFOLIUM ROOT BARK EXTRACT|BERBERIS AQUIFOLIUM ROOT BARK EXTRACT
C3487959|T121|1347563|RXNORM|MELILOTUS OFFICINALIS TOP EXTRACT|MELILOTUS OFFICINALIS TOP EXTRACT
C2183735|T121|820457|RXNORM|DIPHENHYDRAMINE / PYRILAMINE|DIPHENHYDRAMINE / PYRILAMINE
C0079488|T007|1318501|RXNORM|HELICOBACTER PYLORI|HELICOBACTER PYLORI
C3651728|T121|1429969|RXNORM|LONICERA CAPRIFOLIUM FLOWERING TOP EXTRACT|LONICERA CAPRIFOLIUM FLOWERING TOP EXTRACT
C0022252|T121|6058|RXNORM|ISOSORBIDE DINITRATE|ISOSORBIDE DINITRATE
C0022245|T121|6054|RXNORM|ISOPROTERENOL|ISOPROTERENOL
C0022245|T121|6054|RXNORM|ISOPROTERENOL|ISOPROTERENOL
C0022251|T121|6057|RXNORM|ISOSORBIDE|ISOSORBIDE
C0022251|T121|6057|RXNORM|ISOSORBIDE|ISOSORBIDE
C2364498|T129|805469|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED, A-H3N2 (A-URUGUAY-716-2007) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED, A-H3N2 (A-URUGUAY-716-2007) STRAIN
C1876564|T121|700888|RXNORM|CHROMIUM POLYNICOTINATE|CHROMIUM POLYNICOTINATE
C2057679|T121|1006923|RXNORM|NOVOBIOCIN / TETRACYCLINE|NOVOBIOCIN / TETRACYCLINE
C3864975|T121|1594955|RXNORM|CAPSAICIN / LIDOCAINE / MENTHOL|CAPSAICIN / LIDOCAINE / MENTHOL
C0009137|T121|2635|RXNORM|COAL TAR|COAL TAR
C0063371|T131|1442172|RXNORM|ENILCONAZOLE|ENILCONAZOLE
C3486391|T121|1322547|RXNORM|CYNARA SCOLYMUS LEAF EXTRACT|CYNARA SCOLYMUS LEAF EXTRACT
C0982221|T125|314684|RXNORM|INSULIN, PROTAMINE LISPRO, HUMAN|INSULIN, PROTAMINE LISPRO, HUMAN
C0982224|T125|314685|RXNORM|INSULIN, PROTAMINE ZINC, BEEF-PORK|INSULIN, PROTAMINE ZINC, BEEF-PORK
C0982226|T121|314686|RXNORM|INSULIN, REGULAR, BEEF|INSULIN, REGULAR, BEEF
C2682879|T121|845639|RXNORM|DIMETHICONE / ZINC OXIDE|DIMETHICONE / ZINC OXIDE
C0982217|T125|314682|RXNORM|LENTE INSULIN, BEEF-PORK|LENTE INSULIN, BEEF-PORK
C0982219|T125|314683|RXNORM|INSULIN, ZINC, HUMAN|INSULIN, ZINC, HUMAN
C3535859|T121|1370628|RXNORM|CETOSTEARYL SULFATE|CETOSTEARYL SULFATE
C2828272|T197|1370629|RXNORM|MANGANESE ACETATE|MANGANESE ACETATE
C1445804|T168|466570|RXNORM|PUMPKIN SEED OIL|PUMPKIN SEED OIL
C3535862|T121|1370624|RXNORM|STARCH GLYCOLATE TYPE B POTATO|STARCH GLYCOLATE TYPE B POTATO
C3535861|T121|1370625|RXNORM|STEAROYL GLUTAMATE|STEAROYL GLUTAMATE
C3535860|T121|1370626|RXNORM|STEARYL FUMARATE|STEARYL FUMARATE
C3503279|T130|1370627|RXNORM|THIOGLYCOLATE|THIOGLYCOLATE
C3535865|T121|1370620|RXNORM|PALM KERNELATE|PALM KERNELATE
C3503116|T109|1370621|RXNORM|PALMITATE|PALMITATE
C3535864|T109|1370622|RXNORM|PALMITOYL PROLINE|PALMITOYL PROLINE
C3535863|T121|1370623|RXNORM|PYRROLIDONE CARBOXYLATE|PYRROLIDONE CARBOXYLATE
C2722056|T129|904606|RXNORM|PISTACHIO NUT ALLERGENIC EXTRACT|PISTACIA VERA ALLERGENIC EXTRACT
C0937909|T121|969119|RXNORM|ECHINACEA PALLIDA ROOT EXTRACT|ECHINACEA PALLIDA ROOT EXTRACT
C0369845|T195|113831|RXNORM|PIPEMIDATE|PIPEMIDATE
C2729782|T129|891752|RXNORM|AMERICAN CHESTNUT ALLERGENIC EXTRACT|CASTANEA DENTATA ALLERGENIC EXTRACT
C2927539|T129|1006297|RXNORM|ASPERGILLUS NIGER VAR. NIGER ALLERGENIC EXTRACT|ASPERGILLUS NIGER VAR. NIGER ALLERGENIC EXTRACT
C3537535|T109|1370992|RXNORM|BARBASCO EXTRACT|BARBASCO EXTRACT
C3537533|T109|1370990|RXNORM|PLANATUS OCCIDENTALIS BARK EXTRACT|PLANATUS OCCIDENTALIS BARK EXTRACT
C3537534|T109|1370991|RXNORM|BILBERRY SEED EXTRACT|BILBERRY SEED EXTRACT
C3257375|T121|1242095|RXNORM|ETHANOL / ISOPROPYL ALCOHOL / POVIDONE-IODINE|ETHANOL / ISOPROPYL ALCOHOL / POVIDONE-IODINE
C3256960|T109|1305532|RXNORM|TANGERINE PEEL EXTRACT|TANGERINE PEEL EXTRACT
C1875027|T121|690690|RXNORM|DIPHENHYDRAMINE / GUAIFENESIN / MENTHOL / SODIUM CITRATE|DIPHENHYDRAMINE / GUAIFENESIN / MENTHOL / SODIUM CITRATE
C0012702|T121|3541|RXNORM|DISOPYRAMIDE|DISOPYRAMIDE
C1875029|T121|690692|RXNORM|DIPHENHYDRAMINE / PHENOL|DIPHENHYDRAMINE / PHENOL
C1330000|T121|690693|RXNORM|DIPHENHYDRAMINE / PHENYLEPHRINE|DIPHENHYDRAMINE / PHENYLEPHRINE
C0771864|T121|236573|RXNORM|LITHIUM HYDROGEN ASPARTATE|LITHIUM HYDROGEN ASPARTATE
C0055578|T121|20976|RXNORM|OXTRIPHYLLINE|CHOLINE THEOPHYLLINATE
C1143123|T121|341379|RXNORM|NITENPYRAM|NITENPYRAM
C1875269|T121|692832|RXNORM|HYDROFLUORIC ACID / SODIUM FLUORIDE / STANNOUS FLUORIDE|HYDROFLUORIC ACID / SODIUM FLUORIDE / STANNOUS FLUORIDE
C1166210|T121|350490|RXNORM|URTICA DIOICA PREPARATION|URTICA DIOICA PREPARATION
C1875267|T121|692830|RXNORM|HYDROFLUORIC ACID / PHOSPHORIC ACID / SODIUM FLUORIDE|HYDROFLUORIC ACID / PHOSPHORIC ACID / SODIUM FLUORIDE
C1875268|T121|692831|RXNORM|HYDROFLUORIC ACID / SODIUM FLUORIDE|HYDROFLUORIC ACID / SODIUM FLUORIDE
C0031700|T197|8259|RXNORM|PHOSPHORIC ACID|PHOSPHORIC ACID
C0053800|T131|1433347|RXNORM|BISPHENOL A|BISPHENOL A
C1174115|T109|1364296|RXNORM|ISOBUTYLPARABEN|ISOBUTYLPARABEN
C2194278|T121|814818|RXNORM|DEXTROMETHORPHAN / METHOXYPHENAMINE|DEXTROMETHORPHAN / METHOXYPHENAMINE
C3536724|T121|1433760|RXNORM|ERODIUM CICUTARIUM EXTRACT|ERODIUM CICUTARIUM EXTRACT
C0010524|T131|2969|RXNORM|CYCLAMATE|CYCLAMATE
C0010523|T195|2968|RXNORM|CYCLACILLIN|CYCLACILLIN
C2025629|T121|814761|RXNORM|CELLULASE / DIAZEPAM / FENIPENTOL / PANCREATIN|CELLULASE / DIAZEPAM / FENIPENTOL / PANCREATIN
C2928858|T121|1007945|RXNORM|ADIPIC ACID / AMMONIUM|ADIPIC ACID / AMMONIUM
C2929628|T121|1008729|RXNORM|DIMETHICONE / TITANIUM DIOXIDE|DIMETHICONE / TITANIUM DIOXIDE
C2929627|T121|1008728|RXNORM|ALLANTOIN / BENZOCAINE / CAMPHOR / DIMETHICONE / PETROLATUM|ALLANTOIN / BENZOCAINE / CAMPHOR / DIMETHICONE / PETROLATUM
C2929625|T121|1008726|RXNORM|MECLIZINE / NIACIN|MECLIZINE / NIACIN
C3163163|T121|1115799|RXNORM|MAGNESIUM CITRATE / MAGNESIUM OXIDE / POTASSIUM CITRATE / PYRIDOXINE|MAGNESIUM CITRATE / MAGNESIUM OXIDE / POTASSIUM CITRATE / PYRIDOXINE
C2929623|T121|1008724|RXNORM|NIACIN / RIBOFLAVIN|NIACIN / RIBOFLAVIN
C2929622|T121|1008723|RXNORM|ASCORBIC ACID / FLUORIDE ION / FOLIC ACID / NIACIN / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D / VITAMIN E|ASCORBIC ACID / FLUORIDE ION / FOLIC ACID / NIACIN / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D / VITAMIN E
C2929621|T121|1008722|RXNORM|BORAGE OIL / GAMMA-LINOLENATE / LINOLEATE|BORAGE OIL / GAMMA-LINOLENATE / LINOLEATE
C2929620|T121|1008721|RXNORM|ACETAMINOPHEN / MAGNESIUM SALICYLATE / PAMABROM|ACETAMINOPHEN / MAGNESIUM SALICYLATE / PAMABROM
C2929619|T121|1008720|RXNORM|AMMONIUM CHLORIDE / EPHEDRINE|AMMONIUM CHLORIDE / EPHEDRINE
C2727802|T129|974741|RXNORM|MOSQUITO ALLERGENIC EXTRACT|AEDES TAENIORHYNCHUS ALLERGENIC EXTRACT
C3256767|T109|1309431|RXNORM|GLEHNIA LITTORALIS ROOT EXTRACT|GLEHNIA LITTORALIS ROOT EXTRACT
C2193878|T121|818109|RXNORM|METRONIDAZOLE / SPIRAMYCIN|METRONIDAZOLE / SPIRAMYCIN
C2047874|T121|818102|RXNORM|ACETAMINOPHEN / IBUPROFEN|ACETAMINOPHEN / IBUPROFEN
C3643343|T121|1424459|RXNORM|PALMITOYL LYSYLDIOXYMETHIONYLLYSINE|PALMITOYL LYSYLDIOXYMETHIONYLLYSINE
C3643344|T121|1424458|RXNORM|C9-11 PARETH-8|C9-11 PARETH-8
C2938369|T121|1012111|RXNORM|CHLORCYCLIZINE / CODEINE|CHLORCYCLIZINE / CODEINE
C0066685|T121|30131|RXNORM|MOEXIPRIL|MOEXIPRIL
C0030817|T121|7975|RXNORM|EDTMP|PENICILLAMINE
C0027752|T123|7327|RXNORM|NERVE GROWTH FACTOR|NERVE GROWTH FACTOR
C3855134|T109|1547466|RXNORM|AGRIMONIA PILOSA WHOLE EXTRACT|AGRIMONIA PILOSA WHOLE EXTRACT
C0015846|T121|4337|RXNORM|FENTANYL|FENTANYL
C0057948|T130|1486708|RXNORM|DIETHYLENE GLYCOL DISTEARATE|DIETHYLENE GLYCOL DISTEARATE
C0015840|T121|4333|RXNORM|FENOTEROL|FENOTEROL
C2928856|T121|1007943|RXNORM|OLEANDOMYCIN / TETRACYCLINE|OLEANDOMYCIN / TETRACYCLINE
C0015837|T121|4331|RXNORM|FENOPROFEN|FENOPROFEN
C0011145|T130|3131|RXNORM|DEFEROXAMINE|DEFEROXAMINE
C0047683|T125|14584|RXNORM|ETONOGESTREL|ETONOGESTREL
C3496090|T121|1315126|RXNORM|BLUE CRAB PREPARATION|BLUE CRAB PREPARATION
C3496181|T121|1315124|RXNORM|WHITE RICE EXTRACT|WHITE RICE EXTRACT
C0616779|T121|1315125|RXNORM|BENZOPHENONE-2|BENZOPHENONE-2
C3500696|T121|1315122|RXNORM|SERRATED SWIMMING CRAB, COOKED PREPARATION|SERRATED SWIMMING CRAB, COOKED PREPARATION
C2949233|T121|1046247|RXNORM|ALPHA TOCOPHEROL / LEVOMENTHOL|ALPHA TOCOPHEROL / LEVOMENTHOL
C3496086|T121|1315120|RXNORM|LAMB PREPARATION|LAMB PREPARATION
C3500695|T129|1315121|RXNORM|OYSTER, UNSPECIFIED PREPARATION|OYSTER, UNSPECIFIED PREPARATION
C0521943|T197|133050|RXNORM|ACTIVATED ATTAPULGITE|ACTIVATED ATTAPULGITE
C3488938|T109|1309291|RXNORM|RASPBERRY SEED OIL|RASPBERRY SEED OIL
C3488944|T109|1309290|RXNORM|ROSA RUBIGINOSA SEED OIL|ROSA RUBIGINOSA SEED OIL
C3488988|T109|1309293|RXNORM|CARROT SEED OIL|CARROT SEED OIL
C1138839|T121|1309292|RXNORM|ANISE SEED EXTRACT|ANISE SEED EXTRACT
C3488918|T109|1309295|RXNORM|CITRUS AURANTIIFOLIA LEAF OIL|CITRUS AURANTIIFOLIA LEAF OIL
C3488984|T109|1309294|RXNORM|PRUNELLA VULGARIS FLOWERING TOP EXTRACT|PRUNELLA VULGARIS FLOWERING TOP EXTRACT
C3488956|T109|1309296|RXNORM|PISCIDIA PISCIPULA ROOT BARK EXTRACT|PISCIDIA PISCIPULA ROOT BARK EXTRACT
C0937612|T121|283553|RXNORM|COLA EXTRACT|COLA EXTRACT
C0937610|T121|283551|RXNORM|CINCHONA PUBESCENS PREPARATION|CINCHONA PUBESCENS PREPARATION
C0057834|T131|22895|RXNORM|DICLORAN|DICLORAN
C0937617|T121|283557|RXNORM|DROSERA ROTUNDIFOLIA EXTRACT|DROSERA ROTUNDIFOLIA FLOWERING TOP EXTRACT
C0937615|T121|283556|RXNORM|DELPHINIUM STAPHISAGRIA PREPARATION|DELPHINIUM STAPHISAGRIA PREPARATION
C0937614|T121|283555|RXNORM|CUTTLE FISH INK|CUTTLE FISH INK
C0937613|T121|283554|RXNORM|CORDYCEPS SINENSIS PREPARATION|CORDYCEPS SINENSIS PREPARATION
C3256129|T121|1311665|RXNORM|BRASSICA RAPA VAR. RAPA EXTRACT|BRASSICA RAPA VAR. RAPA EXTRACT
C3256867|T121|1311664|RXNORM|PRUNUS SEROTINA FRUIT EXTRACT|PRUNUS SEROTINA FRUIT EXTRACT
C3256260|T121|1311667|RXNORM|ROSA MULTIFLORA FRUIT EXTRACT|ROSA MULTIFLORA FRUIT EXTRACT
C3464715|T121|1311666|RXNORM|PYRACANTHA FORTUNEANA FRUIT EXTRACT|PYRACANTHA FORTUNEANA FRUIT EXTRACT
C3256866|T121|1311663|RXNORM|PRUNUS MUME FRUIT EXTRACT|PRUNUS MUME FRUIT EXTRACT
C2928855|T121|1007941|RXNORM|ESTRADIOL / ESTRIOL / NORETHINDRONE|ESTRADIOL / ESTRIOL / NORETHINDRONE
C3256261|T121|1311668|RXNORM|ROSA ROXBURGHII FRUIT EXTRACT|ROSA ROXBURGHII FRUIT EXTRACT
C2979049|T121|1090007|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / FOLIC ACID / PHYTOSTEROLS / POLICOSANOL / VITAMIN B 12 / VITAMIN B6|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / FOLIC ACID / PHYTOSTEROLS / POLICOSANOL / VITAMIN B 12 / VITAMIN B6
C0137822|T197|1364922|RXNORM|POLYMETAPHOSPHATE|POLYMETAPHOSPHATE
C0021186|T121|5764|RXNORM|INDAPAMIDE|INDAPAMIDE
C2745274|T121|1545063|RXNORM|TAFAMIDIS|TAFAMIDIS
C0163025|T121|59064|RXNORM|PIPERIDOLATE|PIPERIDOLATE
C2928574|T121|1007658|RXNORM|ACETYLENE / NITROGEN / OXYGEN|ACETYLENE / NITROGEN / OXYGEN
C2928575|T121|1007659|RXNORM|CARBON DIOXIDE / CARBON MONOXIDE / NITROGEN / OXYGEN|CARBON DIOXIDE / CARBON MONOXIDE / NITROGEN / OXYGEN
C2928572|T121|1007656|RXNORM|CARBON DIOXIDE / HYDROGEN / NITROGEN|CARBON DIOXIDE / HYDROGEN / NITROGEN
C2928573|T121|1007657|RXNORM|GINKGO BILOBA EXTRACT / VINCAMINE|GINKGO BILOBA EXTRACT / VINCAMINE
C2928570|T121|1007654|RXNORM|ACETAMINOPHEN / MAGNESIUM SALICYLATE|ACETAMINOPHEN / MAGNESIUM SALICYLATE
C2928571|T121|1007655|RXNORM|GINSENG PREPARATION / GUARANA PREPARATION|GINSENG PREPARATION / GUARANA PREPARATION
C2928568|T121|1007652|RXNORM|MENTHOL / PEPPERMINT OIL|MENTHOL / PEPPERMINT OIL
C2928569|T121|1007653|RXNORM|CHLOROBUTANOL / POSTERIOR PITUITARY HORMONES|CHLOROBUTANOL / POSTERIOR PITUITARY HORMONES
C2928566|T121|1007650|RXNORM|GUAIACOLSULFONATE / MORPHINE|GUAIACOLSULFONATE / MORPHINE
C2928567|T121|1007651|RXNORM|ESTROGENS, CONJUGATED (USP) / ESTRONE|ESTROGENS, CONJUGATED (USP) / ESTRONE
C0061347|T121|25806|RXNORM|CALCIUM GLUBIONATE|CALCIUM GLUBIONATE
C3265058|T121|1244007|RXNORM|ASCORBIC ACID / CHOLECALCIFEROL / FERROUS SULFATE / SODIUM FLUORIDE / VITAMIN A|ASCORBIC ACID / CHOLECALCIFEROL / FERROUS SULFATE / SODIUM FLUORIDE / VITAMIN A
C0718043|T126|214817|RXNORM|SACROSIDASE|SACROSIDASE
C1875122|T121|691251|RXNORM|ERGOTAMINE / HYOSCYAMINE / PHENOBARBITAL|ERGOTAMINE / HYOSCYAMINE / PHENOBARBITAL
C2741444|T129|901203|RXNORM|SUNFLOWER SEED ALLERGENIC EXTRACT|HELIANTHUS ANNUUS SEED ALLERGENIC EXTRACT
C1001866|T007|1550045|RXNORM|BIFIDOBACTERIUM ANIMALIS|BIFIDOBACTERIUM ANIMALIS
C2073864|T121|812621|RXNORM|ACETAMINOPHEN / ASCORBIC ACID / CAFFEINE / CHLORPHENIRAMINE / PHENYLEPHRINE|ACETAMINOPHEN / ASCORBIC ACID / CAFFEINE / CHLORPHENIRAMINE / PHENYLEPHRINE
C3693001|T125|1442996|RXNORM|THYROID, OVINE|THYROID, OVINE
C3496793|T121|1307298|RXNORM|ENZALUTAMIDE|ENZALUTAMIDE
C3152793|T129|1098118|RXNORM|CULTIVATED BARLEY POLLEN EXTRACT|HORDEUM VULGARE POLLEN EXTRACT
C0163391|T197|59203|RXNORM|POTASSIUM CHLORATE|POTASSIUM CHLORATE
C3265918|T168|1309337|RXNORM|CHINESE CINNAMON OIL|CHINESE CINNAMON OIL
C1692318|T121|82003|RXNORM|DOCUSATE|DOCUSATE
C1692318|T121|82003|RXNORM|DOCUSATE|DOCUSATE
C0000956|T121|154|RXNORM|ROTAVIRUS VACCINES|ACENOCOUMAROL
C0010552|T121|2978|RXNORM|CYCLOBARBITAL|CYCLOBARBITAL
C0028095|T121|7427|RXNORM|NIMORAZOLE|NIMORAZOLE
C0121902|T121|50975|RXNORM|HISTRELIN|HISTRELIN
C2701243|T129|852029|RXNORM|MUGWORT SAGE POLLEN EXTRACT|ARTEMISIA VULGARIS POLLEN EXTRACT
C0028089|T121|7424|RXNORM|NIKETHAMIDE|NIKETHAMIDE
C0028073|T121|7421|RXNORM|NIFURTIMOX|NIFURTIMOX
C0247194|T121|73178|RXNORM|ILOPERIDONE|ILOPERIDONE
C2731191|T129|894750|RXNORM|PARA GRASS POLLEN EXTRACT|UROCHLOA MUTICA POLLEN EXTRACT
C0981863|T129|852020|RXNORM|COMMON SAGEBRUSH POLLEN EXTRACT|ARTEMISIA TRIDENTATA POLLEN EXTRACT
C0795617|T121|253172|RXNORM|GRAPE EXTRACT|GRAPE EXTRACT
C2701239|T129|852025|RXNORM|COCKLEBUR POLLEN EXTRACT|XANTHIUM STRUMARIUM POLLEN EXTRACT
C0050175|T121|16521|RXNORM|ADEFOVIR|ADEFOVIR
C3538278|T121|1372478|RXNORM|ASARUM HETEROTROPOIDES EXTRACT|ASARUM HETEROTROPOIDES EXTRACT
C0070203|T121|32987|RXNORM|PECTIN|PECTIN
C2928357|T121|1007435|RXNORM|METOCLOPRAMIDE / PAPAIN / SIMETHICONE|METOCLOPRAMIDE / PAPAIN / SIMETHICONE
C2928354|T121|1007432|RXNORM|NITROFURANTOIN / PHENAZOPYRIDINE / SULFADIAZINE|NITROFURANTOIN / PHENAZOPYRIDINE / SULFADIAZINE
C3486742|T121|1330088|RXNORM|SPONGILLA LACUSTRIS EXTRACT|SPONGILLA LACUSTRIS EXTRACT
C3486765|T121|1330089|RXNORM|OKOUBAKA AUBREVILLEI BARK EXTRACT|OKOUBAKA AUBREVILLEI BARK EXTRACT
C0024547|T131|6606|RXNORM|MALATHION|MALATHION
C0060440|T109|1536070|RXNORM|FLAVONE|FLAVONE
C3484530|T129|1330085|RXNORM|BEEF LIVER PREPARATION|BEEF LIVER PREPARATION
C0044923|T121|12449|RXNORM|GEMEPROST|GEMEPROST
C0383765|T197|1366982|RXNORM|SODIUM OXIDE|SODIUM OXIDE
C0085795|T195|42527|RXNORM|AMPHOTERICIN|AMPHOTERICIN
C1873953|T121|689566|RXNORM|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE
C1873954|T121|689567|RXNORM|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE
C1873949|T121|689561|RXNORM|ACETAMINOPHEN / BUTALBITAL / CAFFEINE / CODEINE|ACETAMINOPHEN / BUTALBITAL / CAFFEINE / CODEINE
C1873950|T121|689562|RXNORM|ACETAMINOPHEN / BUTALBITAL / CAFFEINE / HYDROCODONE|ACETAMINOPHEN / BUTALBITAL / CAFFEINE / HYDROCODONE
C1873951|T121|689563|RXNORM|ACETAMINOPHEN / BUTALBITAL / CODEINE|ACETAMINOPHEN / BUTALBITAL / CODEINE
C2927988|T121|1007065|RXNORM|CARBETAPENTANE CITRATE / CARBETAPENTANE TANNATE / PHENYLEPHRINE HYDROCHLORIDE / PHENYLEPHRINE TANNATE|CARBETAPENTANE CITRATE / CARBETAPENTANE TANNATE / PHENYLEPHRINE HYDROCHLORIDE / PHENYLEPHRINE TANNATE
C0291140|T126|84959|RXNORM|IMIGLUCERASE|IMIGLUCERASE
C1873955|T121|689568|RXNORM|ACETAMINOPHEN / CAFFEINE / CODEINE / SALICYLAMIDE|ACETAMINOPHEN / CAFFEINE / CODEINE / SALICYLAMIDE
C1873956|T121|689569|RXNORM|ACETAMINOPHEN / CAFFEINE / DIHYDROCODEINE|ACETAMINOPHEN / CAFFEINE / DIHYDROCODEINE
C0601126|T121|1426773|RXNORM|DIPENTAMETHYLENETHIURAM DISULFIDE|DIPENTAMETHYLENETHIURAM DISULFIDE
C3488915|T109|1309338|RXNORM|EAST INDIAN LEMONGRASS OIL|EAST INDIAN LEMONGRASS OIL
C0969943|T121|1426777|RXNORM|LIMONENE, (-)-|LIMONENE, (-)-
C0724600|T125|221108|RXNORM|NPH INSULIN, PORK|INSULIN PORK, ISOPHANE
C0724601|T125|221109|RXNORM|INSULIN, REGULAR, PORK|INSULIN, REGULAR, PORK
C0076370|T196|1309339|RXNORM|THALLIUM SULFATE|THALLIUM SULFATE
C3856083|T121|1549554|RXNORM|ALISMA PLANTAGO-AQUATICA WHOLE EXTRACT|ALISMA PLANTAGO-AQUATICA WHOLE EXTRACT
C0055645|T197|21032|RXNORM|CHROMOUS CHLORIDE|CHROMOUS CHLORIDE
C0069388|T130|1495079|RXNORM|SOLVENT RED 27|SOLVENT RED 27
C3818742|T109|1495078|RXNORM|PPG-12-PEG-50 LANOLIN|PPG-12-PEG-50 LANOLIN
C3666710|T121|1437550|RXNORM|C10-16 PARETH-1|C10-16 PARETH-1
C3666711|T121|1437551|RXNORM|C9-11 PARETH-3|C9-11 PARETH-3
C3818743|T109|1495075|RXNORM|ISOTHIAZOLE|ISOTHIAZOLE
C0066562|T121|1495077|RXNORM|MINAXOLONE|MINAXOLONE
C3464111|T121|1291283|RXNORM|BENZALKONIUM / UREA|BENZALKONIUM / UREA
C3818744|T109|1495073|RXNORM|ISODECYL ISONONANOATE|ISODECYL ISONONANOATE
C0717400|T121|214212|RXNORM|AMILORIDE / HYDROCHLOROTHIAZIDE|AMILORIDE / HYDROCHLOROTHIAZIDE
C3663719|T121|1433642|RXNORM|DIMETHYL SEBACATE|DIMETHYL SEBACATE
C1714089|T109|1433643|RXNORM|PEG-5 SOY STEROL|PEG-5 SOY STEROL
C0717404|T121|214216|RXNORM|AMINOPHYLLINE / GUAIFENESIN|AMINOPHYLLINE / GUAIFENESIN
C3663718|T121|1433641|RXNORM|DAEMONOROPS DRACO WHOLE EXTRACT|DAEMONOROPS DRACO WHOLE EXTRACT
C2078991|T121|816868|RXNORM|IODINE / VITAMIN A|IODINE / VITAMIN A
C1875165|T121|689306|RXNORM|FLURANDRENOLIDE / NEOMYCIN|FLURANDRENOLIDE / NEOMYCIN
C0000608|T121|99|RXNORM|DIPHENHYDRAMINE / LIDOCAINE / NYSTATIN|6-AMINOCAPROIC ACID
C1311893|T122|1425088|RXNORM|3-(TRIETHOXYSILYL)PROPYLAMINE|3-(TRIETHOXYSILYL)PROPYLAMINE
C1706570|T109|1425087|RXNORM|SANDALWOOD EXTRACT|SANDALWOOD EXTRACT
C1874669|T121|691033|RXNORM|CALCIUM IODIDE / ISOPROTERENOL|CALCIUM IODIDE / ISOPROTERENOL
C3642395|T121|1423797|RXNORM|MAHONIA AQUIFOLIUM WHOLE EXTRACT|MAHONIA AQUIFOLIUM WHOLE EXTRACT
C2701733|T129|852680|RXNORM|RED MULBERRY POLLEN EXTRACT|MORUS RUBRA POLLEN EXTRACT
C2725037|T121|880688|RXNORM|DIHYDROCODEINE / GUAIFENESIN / PHENYLEPHRINE|DIHYDROCODEINE / GUAIFENESIN / PHENYLEPHRINE
C0008196|T121|2358|RXNORM|CHLORHEXIDINE|CHLORHEXIDINE
C0008196|T121|2358|RXNORM|CHLORHEXIDINE|CHLORHEXIDINE
C3153766|T121|1100065|RXNORM|FAMOTIDINE / IBUPROFEN|FAMOTIDINE / IBUPROFEN
C0008174|T121|2353|RXNORM|CLORAZEPATE|CLORAZEPATE
C1874666|T121|691030|RXNORM|CALCIUM GLYCEROPHOSPHATE / CALCIUM LEVULINATE|CALCIUM GLYCEROPHOSPHATE / CALCIUM LEVULINATE
C0008188|T121|2356|RXNORM|CHLORDIAZEPOXIDE|CHLORDIAZEPOXIDE
C0008183|T121|2354|RXNORM|CHLORCYCLIZINE|CHLORCYCLIZINE
C1527027|T195|877510|RXNORM|ROMIDEPSIN|ROMIDEPSIN
C3667092|T121|1438509|RXNORM|PEARL (HYRIOPSIS CUMINGII) EXTRACT|PEARL (HYRIOPSIS CUMINGII) EXTRACT
C2194018|T121|813869|RXNORM|BETAMETHASONE / DEXCHLORPHENIRAMINE|BETAMETHASONE / DEXCHLORPHENIRAMINE
C0006674|T127|1894|RXNORM|CALCITRIOL|CALCITRIOL
C0006674|T127|1894|RXNORM|CALCITRIOL|CALCITRIOL
C0006675|T196|1895|RXNORM|CALCIUM|CALCIUM
C0006681|T197|1897|RXNORM|CALCIUM CARBONATE|CALCIUM CARBONATE
C0006681|T197|1897|RXNORM|CALCIUM CARBONATE|CALCIUM CARBONATE
C0006681|T197|1897|RXNORM|CALCIUM CARBONATE|CALCIUM CARBONATE
C3256329|T121|1311153|RXNORM|AMINO METHACRYLATE COPOLYMER|DIMETHYLAMINOETHYL METHACRYLATE - BUTYL METHACRYLATE - METHYL METHACRYLATE COPOLYMER
C2741474|T129|901283|RXNORM|SWORDFISH ALLERGENIC EXTRACT|XIPHIAS GLADIUS ALLERGENIC EXTRACT
C0303458|T196|90574|RXNORM|99 MOLYBDENUM|99 MOLYBDENUM
C0066673|T121|30121|RXNORM|MOCLOBEMIDE|MOCLOBEMIDE
C1313386|T125|400008|RXNORM|INSULIN, GLULISINE, HUMAN|INSULIN, GLULISINE, HUMAN
C0007367|T126|2133|RXNORM|CATALASE|CATALASE
C2747602|T129|966692|RXNORM|ALGAL FUNGI ALLERGENIC EXTRACT|PHYCOMYCES BLAKESLEEANUS ALLERGENIC EXTRACT
C3486834|T121|1311347|RXNORM|SUS SCROFA TEMPORAL LOBE PREPARATION|PORCINE TEMPORAL LOBE PREPARATION
C0017135|T123|4698|RXNORM|GASTRIC MUCINS|GASTRIC MUCINS
C3695973|T121|1483620|RXNORM|ROSA RUGOSA FLOWER BUD EXTRACT|ROSA RUGOSA FLOWER BUD EXTRACT
C2702372|T129|892632|RXNORM|POTATO ALLERGENIC EXTRACT|POTATO ALLERGENIC EXTRACT
C3538502|T121|1372927|RXNORM|GYNOSTEMMA PENTAPHYLLUM TOP EXTRACT|GYNOSTEMMA PENTAPHYLLUM TOP EXTRACT
C3255933|T109|1372926|RXNORM|DICAPRYLYL CARBONATE|DICAPRYLYL CARBONATE
C3695960|T122|1484396|RXNORM|PEG-80 STEARATE|PEG-80 STEARATE
C3538504|T121|1372929|RXNORM|DISTEARDIMONIUM HECTORITE|DISTEARDIMONIUM HECTORITE
C3538503|T121|1372928|RXNORM|HETEROTHECA INULOIDES FLOWER EXTRACT|HETEROTHECA INULOIDES FLOWER EXTRACT
C0357080|T121|105669|RXNORM|POLYSACCHARIDE IRON COMPLEX|POLYSACCHARIDE IRON COMPLEX
C3848528|T121|1546427|RXNORM|ETHYLMERCURITHIOSALICYLIC ACID|ETHYLMERCURITHIOSALICYLIC ACID
C2342354|T109|1367138|RXNORM|DICAPRYLYL ETHER|DICAPRYLYL ETHER
C2356501|T121|1367139|RXNORM|ETHYLHEXYL ISONONANOATE|ETHYLHEXYL ISONONANOATE
C1613432|T121|1367134|RXNORM|ETHYLHEXYLGLYCERIN|ETHYLHEXYLGLYCERIN
C1655177|T197|1367135|RXNORM|STANNOUS OXIDE|STANNOUS OXIDE
C1814776|T121|1367136|RXNORM|NEOPENTYL GLYCOL DIISOSTEARATE|NEOPENTYL GLYCOL DIISOSTEARATE
C0301185|T122|1367137|RXNORM|DIBUTYL ADIPATE|DIBUTYL ADIPATE
C1509712|T121|1367130|RXNORM|POLYGLYCERYL-4 ISOSTEARATE|POLYGLYCERYL-4 ISOSTEARATE
C1509774|T109|1367131|RXNORM|STEARETH-100|STEARETH-100
C1533418|T122|1367133|RXNORM|POLYOXYL 8 STEARATE|POLYETHYLENE GLYCOL 400 MONOSTEARATE
C3486577|T131|1309761|RXNORM|TOXICODENDRON VERNIX LEAFY TWIG EXTRACT|TOXICODENDRON VERNIX LEAFY TWIG EXTRACT
C3488686|T121|1309763|RXNORM|SOLIDAGO VIRGAUREA FLOWERING TOP EXTRACT|SOLIDAGO VIRGAUREA FLOWERING TOP EXTRACT
C3486583|T121|1309762|RXNORM|NUPHAR LUTEUM ROOT EXTRACT|NUPHAR LUTEUM ROOT EXTRACT
C3487976|T121|1309764|RXNORM|KRAMERIA LAPPACEA ROOT EXTRACT|KRAMERIA LAPPACEA ROOT EXTRACT
C3486586|T121|1309767|RXNORM|PTERIDIUM AQUILINUM ROOT EXTRACT|PTERIDIUM AQUILINUM ROOT EXTRACT
C3488687|T121|1309766|RXNORM|BERBERIS VULGARIS ROOT BARK EXTRACT|BERBERIS VULGARIS ROOT BARK EXTRACT
C1872203|T121|1364105|RXNORM|PASIREOTIDE|PASIREOTIDE
C3528920|T121|1363730|RXNORM|SAMBUCUS NIGRA WHOLE EXTRACT|SAMBUCUS NIGRA WHOLE EXTRACT
C3486835|T121|1311348|RXNORM|SUS SCROFA PARATHYROID GLAND PREPARATION|PORCINE PARATHYROID GLAND PREPARATION
C0795585|T121|253157|RXNORM|BEE POLLEN|BEE POLLEN
C0770612|T121|235524|RXNORM|LICORICE ROOT EXTRACT|LICORICE ROOT EXTRACT
C1533519|T121|477531|RXNORM|ECHINACEA PURPUREA AERIAL PARTS EXTRACT|ECHINACEA PURPUREA AERIAL PARTS EXTRACT
C1166245|T121|350520|RXNORM|CARDUUS MARIANUS PREPARATION|CARDUUS MARIANUS PREPARATION
C3256031|T121|1363596|RXNORM|DIETHYLHEXYL 2,6-NAPHTHALATE|DIETHYLHEXYL 2,6-NAPHTHALATE
C0982120|T121|1363597|RXNORM|DIGLYCOL STEARATE|DIGLYCOL STEARATE
C3256028|T109|1363594|RXNORM|DIETHANOLAMINE BIS(C8-C18 PERFLUOROALKYLETHYL)PHOSPHATE|DIETHANOLAMINE BIS(C8-C18 PERFLUOROALKYLETHYL)PHOSPHATE
C3256029|T121|1363595|RXNORM|DIETHANOLAMINE CETYL PHOSPHATE|DIETHANOLAMINE CETYL PHOSPHATE
C0915913|T109|1363593|RXNORM|COCAMIDOPROPYL HYDROXYSULTAINE|COCAMIDOPROPYL HYDROXYSULTAINE
C3256013|T121|1363590|RXNORM|HYPROMELLOSE 2910 50CP|HYPROMELLOSE 2910 50CP
C3644402|T121|1424840|RXNORM|ASCORBIC ACID / CHOLECALCIFEROL|ASCORBIC ACID / CHOLECALCIFEROL
C3153223|T121|1098755|RXNORM|CHLOPHEDIANOL / PSEUDOEPHEDRINE / TRIPROLIDINE|CHLOPHEDIANOL / PSEUDOEPHEDRINE / TRIPROLIDINE
C3256038|T109|1363598|RXNORM|DIHYDROXYETHYL COCAMINE OXIDE|DIHYDROXYETHYL COCAMINE OXIDE
C3256040|T121|1363599|RXNORM|DIISOBUTYL ADIPATE|DIISOBUTYL ADIPATE
C0874066|T121|260039|RXNORM|SANGRE DE GRADO|SANGRE DE GRADO
C0874065|T121|260038|RXNORM|KOREAN GINSENG ROOT|KOREAN GINSENG ROOT
C0074714|T121|36669|RXNORM|SOBREROL|SOBREROL
C3538276|T121|1372476|RXNORM|RHUS CHINENSIS WHOLE EXTRACT|RHUS CHINENSIS WHOLE EXTRACT
C0009213|T168|2669|RXNORM|P-AMINOSALICYLIC ACID MONOSODIUM SALT|COD LIVER OIL
C0908935|T121|275635|RXNORM|DESLORATADINE|DESLORATADINE
C0023401|T123|6308|RXNORM|LEUCINE|LEUCINE
C2927926|T121|1007003|RXNORM|ACEBUTOLOL / MEFRUSIDE|ACEBUTOLOL / MEFRUSIDE
C2927925|T121|1007002|RXNORM|PENTOSAN POLYSULFATE / TROXERUTIN / XANTHINOL|PENTOSAN POLYSULFATE / TROXERUTIN / XANTHINOL
C1639214|T121|608716|RXNORM|DIBUCAINE / HYDROCORTISONE|DIBUCAINE / HYDROCORTISONE
C1639214|T121|608716|RXNORM|DIBUCAINE / HYDROCORTISONE|DIBUCAINE / HYDROCORTISONE
C2927923|T121|1007000|RXNORM|COLISTIN / FURAZOLIDONE|COLISTIN / FURAZOLIDONE
C2927930|T121|1007007|RXNORM|LORATADINE / POVIDONE|LORATADINE / POVIDONE
C2927929|T121|1007006|RXNORM|ACTIVATED CHARCOAL / SALICYLIC ACID / SULFUR|ACTIVATED CHARCOAL / SALICYLIC ACID / SULFUR
C2927928|T121|1007005|RXNORM|ASPIRIN / QUININE|ASPIRIN / QUININE
C2927927|T121|1007004|RXNORM|CHLOROTHEOPHYLLINE / DIPHENHYDRAMINE|CHLOROTHEOPHYLLINE / DIPHENHYDRAMINE
C2057737|T121|818865|RXNORM|ALBUTEROL / KETOTIFEN / THEOPHYLLINE|ALBUTEROL / KETOTIFEN / THEOPHYLLINE
C2927932|T121|1007009|RXNORM|IODOQUINOL / PAPAVERINE / PHTHALYLSULFATHIAZOLE|IODOQUINOL / PAPAVERINE / PHTHALYLSULFATHIAZOLE
C2927931|T121|1007008|RXNORM|ALGINIC ACID / CARBOXYMETHYLCELLULOSE|ALGINIC ACID / CARBOXYMETHYLCELLULOSE
C3538556|T121|1373038|RXNORM|VITIS VINIFERA LEAF EXTRACT|VITIS VINIFERA LEAF EXTRACT
C0010029|T168|2854|RXNORM|CORN OIL|CORN OIL
C2928170|T121|1007248|RXNORM|CALCIUM PHOSPHATE / PHOSPHORUS|CALCIUM PHOSPHATE / PHOSPHORUS
C3488921|T109|1309350|RXNORM|MALVA SYLVESTRIS FLOWER EXTRACT|HIGH MALLOW FLOWER EXTRACT
C1122087|T129|327361|RXNORM|ADALIMUMAB|ADALIMUMAB
C3488919|T121|1309352|RXNORM|MAGNOLIA GRANDIFLORA FLOWER EXTRACT|MAGNOLIA GRANDIFLORA FLOWER EXTRACT
C3488907|T109|1309353|RXNORM|LIGUSTICUM SINENSE ROOT EXTRACT|LIGUSTICUM SINENSE ROOT EXTRACT
C3265864|T109|1309354|RXNORM|HELICHRYSUM ITALICUM FLOWER OIL|HELICHRYSUM ITALICUM FLOWER OIL
C3818705|T109|1535606|RXNORM|PEG-14 DIMETHICONE|PEG-14 DIMETHICONE
C3265488|T121|1244924|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL / VITAMIN K|CALCIUM CARBONATE / CHOLECALCIFEROL / VITAMIN K
C3488912|T109|1309358|RXNORM|HELICHRYSUM ITALICUM FLOWERING TOP EXTRACT|HELICHRYSUM ITALICUM FLOWERING TOP EXTRACT
C3488913|T109|1309359|RXNORM|HIPPOPHAE RHAMNOIDES SEED OIL|HIPPOPHAE RHAMNOIDES SEED OIL
C2343925|T121|797431|RXNORM|MENTHOL / PETROLATUM / PRAMOXINE|MENTHOL / PETROLATUM / PRAMOXINE
C0025668|T121|6847|RXNORM|METHOHEXITAL|METHOHEXITAL
C0025659|T121|6845|RXNORM|METHOCARBAMOL|METHOCARBAMOL
C0068333|T121|31447|RXNORM|ALLERGENIC EXTRACT, WEED, WEST MIX|NABILONE
C0068333|T121|31447|RXNORM|ALLERGENIC EXTRACT, WASP|NABILONE
C0981986|T130|314470|RXNORM|ALLERGENIC EXTRACT, WALNUT|WALNUT ALLERGENIC EXTRACT
C0016677|T007|1432988|RXNORM|FRANCISELLA TULARENSIS|FRANCISELLA TULARENSIS
C0065888|T130|29459|RXNORM|MEGLUMINE IOXITHALAMATE|MEGLUMINE IOXITHALAMATE
C0068333|T121|31447|RXNORM|ALLERGENIC EXTRACT, WESTERN RAGWEED|NABILONE
C0533153|T121|137939|RXNORM|SILVER ACETATE|SILVER ACETATE
C0068333|T121|31447|RXNORM|ALLERGENIC EXTRACT,YELLOW JACKET|NABILONE
C1874796|T121|689367|RXNORM|CHLOROTHEN / METHAPYRILENE / PYRILAMINE|CHLOROTHEN / METHAPYRILENE / PYRILAMINE
C3486787|T121|1311320|RXNORM|SUS SCROFA CONJUNCTIVA PREPARATION|PORCINE CONJUNCTIVA PREPARATION
C3486788|T121|1311321|RXNORM|SUS SCROFA CORPUS LUTEUM PREPARATION|PORCINE CORPUS LUTEUM PREPARATION
C3486789|T121|1311322|RXNORM|SUS SCROFA BRONCHUS PREPARATION|PORCINE BRONCHUS PREPARATION
C0076166|T121|37840|RXNORM|TERTATOLOL|TERTATOLOL
C3486794|T121|1311324|RXNORM|SUS SCROFA DIENCEPHALON PREPARATION|PORCINE DIENCEPHALON PREPARATION
C3486795|T121|1311325|RXNORM|SUS SCROFA DUODENUM PREPARATION|PORCINE DUODENUM PREPARATION
C0070975|T121|33632|RXNORM|PHTHALYLSULFATHIAZOLE|PHTHALYLSULFATHIAZOLE
C3486796|T121|1311327|RXNORM|SUS SCROFA EMBRYO PREPARATION|PORCINE EMBRYO PREPARATION
C3486797|T121|1311328|RXNORM|SUS SCROFA ESOPHAGUS PREPARATION|PORCINE ESOPHAGUS PREPARATION
C3486800|T121|1311329|RXNORM|SUS SCROFA JEJUNUM PREPARATION|PORCINE JEJUNUM PREPARATION
C0770343|T126|235379|RXNORM|PANCRELIPASE|PANCRELIPASE
C2350866|T121|1045453|RXNORM|ERIBULIN|ERIBULIN
C2929196|T121|1008289|RXNORM|GLYCERIN / PETROLATUM|GLYCERIN / PETROLATUM
C3663403|T121|1432985|RXNORM|CHOLECALCIFEROL / INULIN|CHOLECALCIFEROL / INULIN
C0306604|T125|93108|RXNORM|INSULIN, ZINC, PORK|INSULIN, ZINC, PORK
C0137988|T197|54989|RXNORM|ALUMINUM POTASSIUM SULFATE|ALUM
C3256481|T121|1426374|RXNORM|1-GLYCERYL MONOOLEATE|GLYCERYL 1-OLEATE
C3695931|T109|1485119|RXNORM|PEG-6 SORBITAN OLEATE|PEG-6 SORBITAN OLEATE
C0026782|T129|763656|RXNORM|MUMPS VACCINE|MUMPS VACCINE
C0997436|T004|1426666|RXNORM|PENICILLIUM BREVICOMPACTUM|PENICILLIUM BREVICOMPACTUM
C0074710|T121|746741|RXNORM|PRAMIPEXOLE|PRAMIPEXOLE
C3496039|T121|1426667|RXNORM|AVICULARIA AVICULARIA PREPARATION|AVICULARIA AVICULARIA PREPARATION
C0378335|T130|114918|RXNORM|TECHNETIUM TC 99M BICISATE|TECHNETIUM (99MTC) BICISATE
C3475150|T109|1426664|RXNORM|DIMETHICONE 200|DIMETHICONE 200
C0043431|T196|1311498|RXNORM|YTTERBIUM|YTTERBIUM
C0938430|T168|1311499|RXNORM|SEA SALT|SEA SALT
C3496038|T121|1314318|RXNORM|SELAGINELLA TAMARISCINA EXTRACT|SELAGINELLA TAMARISCINA EXTRACT
C0066227|T121|1314316|RXNORM|METHYL BENZOATE|METHYL BENZOATE
C3496735|T121|1314317|RXNORM|PPG-14 PALMETH-60 HEXYL DICARBAMATE|PPG-14 PALMETH-60 HEXYL DICARBAMATE
C0039297|T196|1311490|RXNORM|TANTALUM|TANTALUM
C3475128|T121|1314315|RXNORM|DIMETHYL BENZYL CARBINYL ACETATE|DIMETHYL BENZYL CARBINYL ACETATE
C0040066|T196|1311496|RXNORM|THULIUM|THULIUM
C3256424|T121|1311497|RXNORM|MELISSA OFFICINALIS EXTRACT|MELISSA OFFICINALIS EXTRACT
C0242865|T109|1311494|RXNORM|AMBERGRIS|AMBERGRIS
C3474041|T121|1314311|RXNORM|HALIMEDA OPUNTIA EXTRACT|HALIMEDA OPUNTIA EXTRACT
C3485639|T121|1304496|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / CHOLECALCIFEROL / FOLIC ACID / IRON CARBONYL / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|ALPHA TOCOPHEROL / ASCORBIC ACID / CHOLECALCIFEROL / FOLIC ACID / IRON CARBONYL / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C3486678|T121|1309971|RXNORM|ROBINIA PSEUDOACACIA BARK EXTRACT|ROBINIA PSEUDOACACIA BARK EXTRACT
C3465040|T109|1309972|RXNORM|POLYOXYL 60 CASTOR OIL|POLYOXYL 60 CASTOR OIL
C0993202|T129|901845|RXNORM|ALTERNARIA ALTERNATA ALLERGENIC EXTRACT|ALTERNARIA ALTERNATA ALLERGENIC EXTRACT
C3485672|T121|1313732|RXNORM|2-ETHYLHEXYL BENZOATE|2-ETHYLHEXYL BENZOATE
C2919980|T121|1309979|RXNORM|PASSIFLORA INCARNATA FLOWERING TOP EXTRACT|PASSIFLORA INCARNATA FLOWERING TOP EXTRACT
C0359665|T121|107360|RXNORM|HYPROMELLOSE / PHENYLEPHRINE|HYPROMELLOSE / PHENYLEPHRINE
C1873992|T121|689799|RXNORM|ACETAMINOPHEN / PHENYLTOLOXAMINE / SALICYLAMIDE|ACETAMINOPHEN / PHENYLTOLOXAMINE / SALICYLAMIDE
C1614004|T121|1425503|RXNORM|COCO GLUCOSIDE|COCO GLUCOSIDE
C0110382|T130|1425501|RXNORM|COCHINEAL|COCHINEAL STAIN
C1873991|T121|689797|RXNORM|ACETAMINOPHEN / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE|ACETAMINOPHEN / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE
C1873990|T121|689796|RXNORM|ACETAMINOPHEN / PHENYLPROPANOLAMINE|ACETAMINOPHEN / PHENYLPROPANOLAMINE
C2978509|T121|1089032|RXNORM|BENZOCAINE / CETYLPYRIDINIUM / MENTHOL / TANNIC ACID|BENZOCAINE / CETYLPYRIDINIUM / MENTHOL / TANNIC ACID
C1873989|T121|689794|RXNORM|ACETAMINOPHEN / PHENOBARBITAL|ACETAMINOPHEN / PHENOBARBITAL
C2929457|T121|1008554|RXNORM|ACETAMINOPHEN / CODEINE / MAGNESIUM SALICYLATE / PHENYLTOLOXAMINE|ACETAMINOPHEN / CODEINE / MAGNESIUM SALICYLATE / PHENYLTOLOXAMINE
C2929458|T121|1008555|RXNORM|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / VITAMIN E|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / VITAMIN E
C2929459|T121|1008556|RXNORM|CALCIUM CARBONATE / MAGNESIUM OXIDE / VITAMIN D|CALCIUM CARBONATE / MAGNESIUM OXIDE / VITAMIN D
C2929460|T121|1008557|RXNORM|CHLORPHENIRAMINE / PARAMETHASONE|CHLORPHENIRAMINE / PARAMETHASONE
C2929453|T121|1008550|RXNORM|BROMPHENIRAMINE / CHLOPHEDIANOL / PSEUDOEPHEDRINE|BROMPHENIRAMINE / CHLOPHEDIANOL / PSEUDOEPHEDRINE
C2929454|T121|1008551|RXNORM|DEHYDROCHOLATE / DOCUSATE|DEHYDROCHOLATE / DOCUSATE
C2929455|T121|1008552|RXNORM|ESTROGENS, CONJUGATED (USP) / ESTROGENS, ESTERIFIED (USP) / MEDROXYPROGESTERONE|ESTROGENS, CONJUGATED (USP) / ESTROGENS, ESTERIFIED (USP) / MEDROXYPROGESTERONE
C2731839|T130|896135|RXNORM|SHORT RAGWEED POLLEN EXTRACT|AMBROSIA ARTEMISIIFOLIA POLLEN EXTRACT
C3484795|T121|1303726|RXNORM|BACITRACIN / PRAMOXINE|BACITRACIN / PRAMOXINE
C2929461|T121|1008558|RXNORM|AMPICILLIN / DICLOFENAC|AMPICILLIN / DICLOFENAC
C0717767|T121|1008559|RXNORM|FERROUS FUMARATE / FOLIC ACID|FERROUS FUMARATE / FOLIC ACID
C0142853|T121|56476|RXNORM|SODIUM GLUCONATE|SODIUM GLUCONATE
C0002499|T195|641|RXNORM|AMIKACIN|AMIKACIN
C1874950|T121|690316|RXNORM|DANTHRON / DOCUSATE|DANTHRON / DOCUSATE
C0002502|T121|644|RXNORM|AMILORIDE|AMILORIDE
C1874947|T121|690313|RXNORM|CYCLOPHOSPHAMIDE / MANNITOL|CYCLOPHOSPHAMIDE / MANNITOL
C1874946|T121|690312|RXNORM|CYCLOPENTOLATE / PHENYLEPHRINE|CYCLOPENTOLATE / PHENYLEPHRINE
C0010927|T121|3098|RXNORM|DACARBAZINE|DACARBAZINE
C3257602|T121|1242519|RXNORM|ALLANTOIN / BENZETHONIUM|ALLANTOIN / BENZETHONIUM
C2142879|T121|816996|RXNORM|GUAIFENESIN / PSEUDOEPHEDRINE / TRIPROLIDINE|GUAIFENESIN / PSEUDOEPHEDRINE / TRIPROLIDINE
C3857935|T121|1591920|RXNORM|1-(C14-C18 ESTEROYL)-2-DOCOSAHEXANOYL-SN-GLYCERO-3-PHOSPHOCHOLINE|1-(C14-C18 ESTEROYL)-2-DOCOSAHEXANOYL-SN-GLYCERO-3-PHOSPHOCHOLINE
C3857934|T121|1591921|RXNORM|1-(C14-C18 ESTEROYL)-2-DOCOSAHEXANOYL-SN-GLYCERO-3-PHOSPHOETHANOLAMINE|1-(C14-C18 ESTEROYL)-2-DOCOSAHEXANOYL-SN-GLYCERO-3-PHOSPHOETHANOLAMINE
C3848604|T121|1544634|RXNORM|CUCURBITA PEPO FLOWER EXTRACT|CUCURBITA PEPO FLOWER EXTRACT
C0014939|T125|4100|RXNORM|ESTROGENS|ESTROGENS
C0014942|T125|4103|RXNORM|ESTRONE|ESTRONE
C3864967|T121|1597378|RXNORM|OMBITASVIR / PARITAPREVIR / RITONAVIR|OMBITASVIR / PARITAPREVIR / RITONAVIR
C2701553|T129|852382|RXNORM|WHITE POPLAR POLLEN EXTRACT|POPULUS ALBA POLLEN EXTRACT
C0293359|T125|86009|RXNORM|INSULIN LISPRO|INSULIN LISPRO
C0014960|T121|4106|RXNORM|ETHACRIDINE|ETHACRIDINE
C3159605|T121|1111555|RXNORM|FERROUS BISGLYCINATE / POLYSACCHARIDE IRON COMPLEX|FERROUS BISGLYCINATE / POLYSACCHARIDE IRON COMPLEX
C3852670|T121|1597371|RXNORM|OMBITASVIR|OMBITASVIR
C0358951|T121|1000711|RXNORM|BETAMETHASONE / SALICYLIC ACID|BETAMETHASONE / SALICYLIC ACID
C0005023|T130|1314334|RXNORM|BENZALDEHYDE|BENZALDEHYDE
C0059985|T121|24698|RXNORM|FLUDARABINE|FLUDARABINE
C3257694|T109|1314335|RXNORM|C12-14 ISOPARAFFIN|C12-14 ISOPARAFFIN
C3266878|T121|1333213|RXNORM|IRIS VERSICOLOR ROOT EXTRACT|IRIS VERSICOLOR ROOT EXTRACT
C0036580|T197|9640|RXNORM|SELENITE|SELENITE
C0051511|T197|17610|RXNORM|ALUMINUM CHLORHYDRATE|ALUMINIUM CHLOROHYDRATE
C3267233|T121|1314337|RXNORM|C13-16 ISOPARAFFIN|C13-16 ISOPARAFFIN
C2911925|T121|978140|RXNORM|DIMETHICONE / MENTHOL|DIMETHICONE / MENTHOL
C0064263|T121|28144|RXNORM|EMEDASTINE|EMEDASTINE
C0075160|T197|37032|RXNORM|STANNOUS CHLORIDE|STANNOUS CHLORIDE
C1110602|T121|324028|RXNORM|PETROLEUM PREPARATION|PETROLEUM PREPARATION
C0125339|T121|393540|RXNORM|LAURETH-4|LAURETH-4
C2940212|T130|1014774|RXNORM|CULTIVATED RYE GRASS POLLEN EXTRACT|SECALE CEREALE POLLEN EXTRACT
C1533314|T121|1314333|RXNORM|BEHENTRIMONIUM METHOSULFATE|BEHENTRIMONIUM METHOSULFATE
C2929050|T121|1008143|RXNORM|ASCORBIC ACID / BEE POLLEN|ASCORBIC ACID / BEE POLLEN
C2929049|T121|1008142|RXNORM|ACETAMINOPHEN / ASCORBIC ACID / EUCALYPTOL|ACETAMINOPHEN / ASCORBIC ACID / EUCALYPTOL
C1874348|T121|1008141|RXNORM|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID
C2929047|T121|1008140|RXNORM|CALCIUM POLYSTYRENE SULFONATE PRODUCT / METHYLCELLULOSE|CALCIUM POLYSTYRENE SULFONATE PRODUCT / METHYLCELLULOSE
C2929054|T121|1008147|RXNORM|GINSENG PREPARATION / ST. JOHN'S WORT EXTRACT|GINSENG PREPARATION / ST. JOHN'S WORT EXTRACT
C2929053|T121|1008146|RXNORM|GARLIC PREPARATION / INOSITOL / POLICOSANOL|GARLIC PREPARATION / INOSITOL / POLICOSANOL
C2929052|T121|1008145|RXNORM|EMTRICITABINE / TENOFOVIR DISOPROXIL|EMTRICITABINE / TENOFOVIR DISOPROXIL
C2929051|T121|1008144|RXNORM|LIVER,DESICCATED / PHENOBARBITAL|LIVER,DESICCATED / PHENOBARBITAL
C3488936|T109|1313230|RXNORM|CORYDALIS YANHUSUO TUBER EXTRACT|CORYDALIS YANHUSUO TUBER EXTRACT
C0005018|T197|1375|RXNORM|EPINEPHRINE / LIDOCAINE / TETRACAINE|BENTONITE
C2929056|T121|1008149|RXNORM|DIAZEPAM / FENPROPOREX|DIAZEPAM / FENPROPOREX
C2929055|T121|1008148|RXNORM|CARBON DIOXIDE / HELIUM|CARBON DIOXIDE / HELIUM
C2604598|T109|1313234|RXNORM|TRIHEPTANOIN|TRIHEPTANOIN
C3265134|T109|1313236|RXNORM|PISTACIA LENTISCUS RESIN|PISTACIA LENTISCUS RESIN
C3484432|T121|1310003|RXNORM|VISCUM ALBUM LEAF EXTRACT|VISCUM ALBUM LEAF EXTRACT
C1743856|T109|1426373|RXNORM|OCTADECYLTRIMETHYLAMMONIUM|OCTADECYLTRIMETHYLAMMONIUM
C3853936|T121|1594966|RXNORM|SOLANUM TUBEROSUM EXTRACT|SOLANUM TUBEROSUM EXTRACT
C2726165|T130|968401|RXNORM|TRICHODERMA VIRIDE ALLERGENIC EXTRACT|TRICHODERMA VIRIDE ALLERGENIC EXTRACT
C0022005|T130|5956|RXNORM|IOHEXOL|IOHEXOL
C3555476|T121|1420963|RXNORM|FERULA ASSA-FOETIDA WHOLE EXTRACT|FERULA ASSA-FOETIDA WHOLE EXTRACT
C3555477|T121|1420962|RXNORM|DENDROBIUM NOBILE STEM EXTRACT|DENDROBIUM NOBILE STEM EXTRACT
C3555478|T121|1420961|RXNORM|DAEMONODROPS DRACO RESIN EXTRACT|DAEMONODROPS DRACO RESIN
C2928740|T121|1007825|RXNORM|BELLADONNA ALKALOIDS / CHLORPHENIRAMINE / PSEUDOEPHEDRINE|BELLADONNA ALKALOIDS / CHLORPHENIRAMINE / PSEUDOEPHEDRINE
C3555474|T109|1420965|RXNORM|HYDNOCARPUS KURZII SEED OIL|HYDNOCARPUS KURZII SEED OIL
C0061182|T121|1420964|RXNORM|GELLAN GUM (LOW ACYL)|GELLAN GUM (LOW ACYL)
C1509381|T121|1427070|RXNORM|LAURAMIDE|LAURAMIDE
C3256910|T121|1307609|RXNORM|DENDRANTHEMA INDICUM FLOWER EXTRACT|CHRYSANTHEMUM INDICUM FLOWER EXTRACT
C3255951|T121|1307604|RXNORM|MALPIGHIA EMARGINATA SEED EXTRACT|MALPIGHIA EMARGINATA SEED EXTRACT
C0169964|T125|61148|RXNORM|SOMATROPIN|SOMATROPIN
C3256752|T121|1307606|RXNORM|AVENA SATIVA LEAF EXTRACT|AVENA SATIVA LEAF EXTRACT
C3255945|T121|1307607|RXNORM|MAGNOLIA BIONDII BARK EXTRACT|MAGNOLIA BIONDII BARK EXTRACT
C3282108|T121|1307600|RXNORM|IPOMOEA NIL SEED EXTRACT|IPOMOEA NIL SEED EXTRACT
C3256197|T121|1307601|RXNORM|KHAYA SENEGALENSIS BARK EXTRACT|KHAYA SENEGALENSIS BARK EXTRACT
C3256370|T121|1307602|RXNORM|MORUS AUSTRALIS ROOT EXTRACT|MORUS AUSTRALIS ROOT EXTRACT
C3473228|T121|1307603|RXNORM|MORINGA OLEIFERA BARK EXTRACT|MORINGA OLEIFERA BARK EXTRACT
C0017735|T126|1427073|RXNORM|GLUCOSE OXIDASE|GLUCOSE OXIDASE
C3486821|T121|1309513|RXNORM|SHARK PREPARATION|SHARK PREPARATION
C3485055|T121|1309510|RXNORM|ARTEMISIA CINA FLOWER EXTRACT|ARTEMISIA CINA FLOWER EXTRACT
C2928739|T121|1007824|RXNORM|PSEUDOEPHEDRINE / PYRILAMINE|PSEUDOEPHEDRINE / PYRILAMINE
C0167117|T121|60548|RXNORM|EXENATIDE|EXENATIDE
C3256694|T109|1426449|RXNORM|MICROCOCCUS LUTEUS PREPARATION|MICROCOCCUS LUTEUS PREPARATION
C0054837|T109|1427075|RXNORM|CARVONE|CARVONE
C3499861|T121|1313043|RXNORM|CAPRYLIC-CAPRIC-LAURIC TRIGLYCERIDE|CAPRYLIC-CAPRIC-LAURIC TRIGLYCERIDE
C0025042|T121|6678|RXNORM|MECLOFENAMIC ACID|MECLOFENAMIC ACID
C1318649|T121|401713|RXNORM|CARGLUMIC ACID|CARGLUMIC ACID
C3256632|T109|1309456|RXNORM|POLYGONUM BISTORTA ROOT EXTRACT|POLYGONUM BISTORTA ROOT EXTRACT
C3643361|T109|1421634|RXNORM|DIOCTYLDODECYL DODECANEDIOATE|DIOCTYLDODECYL DODECANEDIOATE
C0056504|T121|21753|RXNORM|CROCONAZOLE|CROCONAZOLE
C2106251|T121|817189|RXNORM|COAL TAR / SULFUR|COAL TAR / SULFUR
C3859818|T129|1594964|RXNORM|PHEASANT FEATHER EXTRACT|PHASIANUS COLCHICUS FEATHER EXTRACT
C1875769|T121|693069|RXNORM|SODIUM CHLORIDE / SODIUM SULFITE / SODIUM THIOSULFATE|SODIUM CHLORIDE / SODIUM SULFITE / SODIUM THIOSULFATE
C0056608|T121|1313047|RXNORM|CURDLAN|CURDLAN
C3499863|T121|1313046|RXNORM|ACETYL OCTAPEPTIDE-3|ACETYL OCTAPEPTIDE-3
C1101838|T121|861634|RXNORM|PITAVASTATIN|PITAVASTATIN
C3818741|T109|1495154|RXNORM|CARTHAMUS TINCTORIUS FLOWER OIL|CARTHAMUS TINCTORIUS FLOWER OIL
C3499862|T121|1313045|RXNORM|GLYCYRRHIZA GLABRA LEAF EXTRACT|GLYCYRRHIZA GLABRA LEAF EXTRACT
C0063252|T121|27340|RXNORM|DESFLURANE|DESFLURANE
C3255664|T109|1426441|RXNORM|ELEMI EXTRACT|CANARIUM LUZONICUM EXTRACT
C0873093|T121|259430|RXNORM|SOY GERM|SOY GERM
C0031618|T123|8215|RXNORM|NAPHAZOLINE / PYRILAMINE|PHOSPHATIDYLETHANOLAMINES
C2073924|T121|821036|RXNORM|CHLORZOXAZONE / IBUPROFEN|CHLORZOXAZONE / IBUPROFEN
C2075857|T121|821034|RXNORM|AMBROXOL / CLOBUTINOL|AMBROXOL / CLOBUTINOL
C3818740|T121|1495155|RXNORM|EUCALYPTUS PIPERITA LEAF EXTRACT|EUCALYPTUS PIPERITA LEAF EXTRACT
C1959892|T121|729517|RXNORM|CODEINE / KAOLIN|CODEINE / KAOLIN
C0873097|T121|259434|RXNORM|SLIPPERY ELM BARK|SLIPPERY ELM BARK
C3245206|T121|1190579|RXNORM|CODEINE / DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE|CODEINE / DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE
C0527189|T121|135391|RXNORM|OLOPATADINE|OLOPATADINE
C0527189|T121|135391|RXNORM|OLOPATADINE|OLOPATADINE
C3643355|T109|1422193|RXNORM|POLOXAMER 403|POLOXAMER 403
C0074742|T197|1422194|RXNORM|SODIUM IODATE|SODIUM IODATE
C0022209|T121|6038|RXNORM|ISONIAZID|ISONIAZID
C0022192|T123|6033|RXNORM|ISOLEUCINE|ISOLEUCINE
C1873993|T121|689802|RXNORM|ACETAMINOPHEN / PSEUDOEPHEDRINE / TRIPROLIDINE|ACETAMINOPHEN / PSEUDOEPHEDRINE / TRIPROLIDINE
C0771161|T197|235954|RXNORM|BISMUTH HYDROXIDE|BISMUTH HYDROXIDE
C0220892|T195|70618|RXNORM|PENICILLIN|PENICILLIN
C0009170|T131|2653|RXNORM|COCAINE|COCAINE
C0220873|T130|70612|RXNORM|MALATE|MALATE
C0220871|T123|70611|RXNORM|LINOLEATE|LINOLEATE
C0369188|T121|113588|RXNORM|ERYTHROMYCIN / SULFISOXAZOLE|ERYTHROMYCIN / SULFISOXAZOLE
C0220884|T123|70616|RXNORM|OLEATE|OLEATE
C3535877|T122|1370606|RXNORM|C12-15 PARETH-3 SULFATE|C12-15 PARETH-3 SULFATE
C3535876|T121|1370607|RXNORM|DIETHYL OXALACETATE|DIETHYL OXALACETATE
C3535879|T121|1370604|RXNORM|SULFOSALICYLATE|SULFOSALICYLATE
C3535878|T121|1370605|RXNORM|ASCORBYL PHOSPHATE|ASCORBYL PHOSPHATE
C3535881|T121|1370602|RXNORM|CAPROAMPHODIPROPIONATE|CAPROAMPHODIPROPIONATE
C3535880|T122|1370603|RXNORM|ETHYLENE DICOCAMIDE PEG-15 DISULFATE|ETHYLENE DICOCAMIDE PEG-15 DISULFATE
C0178627|T130|1370600|RXNORM|ETHYLENEDIAMINETETRAACETATE|ETHYLENEDIAMINETETRAACETATE
C3535882|T121|1370601|RXNORM|XYLENESULFONATE|XYLENESULFONATE
C3535875|T121|1370608|RXNORM|LAUROYL ISETHIONATE|LAUROYL ISETHIONATE
C3535874|T121|1370609|RXNORM|METHYL 2-SULFOLAURATE|METHYL 2-SULFOLAURATE
C1445787|T121|466553|RXNORM|PENICILLIN G BENZATHINE / PENICILLIN G PROCAINE|PENICILLIN G BENZATHINE / PENICILLIN G PROCAINE
C1445789|T121|466555|RXNORM|GUAIFENESIN / PHENYLEPHRINE / PHENYLPROPANOLAMINE|GUAIFENESIN / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C1445790|T121|466556|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN / PHENYLPROPANOLAMINE|DEXTROMETHORPHAN / GUAIFENESIN / PHENYLPROPANOLAMINE
C0017535|T204|1439028|RXNORM|GIARDIA LAMBLIA|GIARDIA LAMBLIA
C3696420|T121|1484769|RXNORM|CHLORHEXIDINE / KETOCONAZOLE / SALICYLOYL PHYTOSPHINGOSINE|CHLORHEXIDINE / KETOCONAZOLE / SALICYLOYL PHYTOSPHINGOSINE
C1337283|T121|969139|RXNORM|HAWTHORN FLOWER EXTRACT|CRATAEGUS LAEVIGATA FLOWER EXTRACT
C0034403|T121|9061|RXNORM|QUINACRINE|QUINACRINE
C3505267|T121|1358176|RXNORM|GENTIANA URNULA FLOWER EXTRACT|GENTIANA URNULA FLOWER EXTRACT
C0072595|T109|1425878|RXNORM|PULLULAN|PULLULAN
C0600190|T122|1425879|RXNORM|NITROCELLULOSE|NITROCELLULOSE
C2016117|T121|820923|RXNORM|ACETAMINOPHEN / AMBROXOL / OXATOMIDE|ACETAMINOPHEN / AMBROXOL / OXATOMIDE
C0039086|T121|10288|RXNORM|SYNEPHRINE|SYNEPHRINE
C0034410|T125|9066|RXNORM|QUINESTROL|QUINESTROL
C0034414|T121|9068|RXNORM|QUINIDINE|QUINIDINE
C3668959|T121|1442792|RXNORM|STACHYS OFFICINALIS EXTRACT|STACHYS OFFICINALIS EXTRACT
C2701182|T129|851942|RXNORM|CANYON RAGWEED POLLEN EXTRACT|AMBROSIA AMBROSIOIDES POLLEN EXTRACT
C0038515|T131|1362878|RXNORM|STYRENE|STYRENE
C0038777|T197|1362879|RXNORM|SULFUR DIOXIDE|SULFUR DIOXIDE
C3855221|T109|1547569|RXNORM|BRASSICA JUNCEA SEED OIL|BRASSICA JUNCEA SEED OIL
C3855220|T109|1547568|RXNORM|BORAGO OFFICINIALIS WHOLE EXTRACT|BORAGO OFFICINIALIS WHOLE EXTRACT
C0001964|T121|1362872|RXNORM|1-PROPANOL|1-PROPANOL
C0056301|T197|21579|RXNORM|COPPER SULFATE|COPPER SULFATE
C0001056|T121|1362871|RXNORM|ACETYLGLUCOSAMINE|N-ACETYLGLUCOSAMINE
C0024574|T130|1362876|RXNORM|MALEIC ANHYDRIDE|MALEIC ANHYDRIDE
C0033434|T109|1362877|RXNORM|PROPANE|PROPANE
C0022683|T197|1362874|RXNORM|DIATOMACEOUS EARTH|DIATOMACEOUS EARTH
C3505265|T121|1358173|RXNORM|GALANTHUS NIVALIS SEED EXTRACT|GALANTHUS NIVALIS SEED EXTRACT
C3282505|T121|1328285|RXNORM|AHNFELTIOPSIS CONCINNA EXTRACT|AHNFELTIOPSIS CONCINNA EXTRACT
C1675326|T121|619693|RXNORM|PERAMIVIR|PERAMIVIR
C1875019|T121|690679|RXNORM|DICYCLOMINE / PHENOBARBITAL|DICYCLOMINE / PHENOBARBITAL
C1875018|T121|690677|RXNORM|DICHLOROTETRAFLUOROETHANE / ETHYL CHLORIDE|DICHLOROTETRAFLUOROETHANE / ETHYL CHLORIDE
C3505263|T197|1358171|RXNORM|CALCIUM ALUMINUM BOROSILICATE|CALCIUM ALUMINUM BOROSILICATE
C0043920|T131|1305516|RXNORM|1,3-DICHLORO-2-PROPANOL|1,3-DICHLORO-2-PROPANOL
C0046095|T109|1305517|RXNORM|2-ETHYLHEXANOIC ACID|2-ETHYLHEXANOIC ACID
C0636819|T121|1305515|RXNORM|1,1-DIFLUOROETHANE|1,1-DIFLUOROETHANE
C0074767|T197|1363697|RXNORM|SODIUM SILICATE|SODIUM SILICATE
C0072222|T121|1363696|RXNORM|PROPYLENE CARBONATE|PROPYLENE CARBONATE
C1655464|T121|605569|RXNORM|CARBINOXAMINE / PHENYLEPHRINE|CARBINOXAMINE / PHENYLEPHRINE
C0016343|T121|4488|RXNORM|FLOXURIDINE|FLOXURIDINE
C0102860|T109|1363698|RXNORM|ALUMINUM TRISTEARATE|ALUMINUM TRISTEARATE
C0010286|T123|2907|RXNORM|CREATINE|CREATINE
C0002611|T197|709|RXNORM|AMMONIUM|AMMONIUM
C0002600|T121|704|RXNORM|AMITRIPTYLINE|AMITRIPTYLINE
C2146620|T121|814290|RXNORM|ACETAMINOPHEN / DOXYLAMINE|ACETAMINOPHEN / DOXYLAMINE
C0002598|T121|703|RXNORM|AMIODARONE|AMIODARONE
C2929607|T121|1008708|RXNORM|PUMPKIN SEED OIL / SAW PALMETTO EXTRACT|PUMPKIN SEED OIL / SAW PALMETTO EXTRACT
C2929600|T121|1008701|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / DOXYLAMINE / PHENYLEPHRINE|ACETAMINOPHEN / DEXTROMETHORPHAN / DOXYLAMINE / PHENYLEPHRINE
C2929602|T121|1008703|RXNORM|MAGNESIUM ACETATE / POTASSIUM ACETATE / SODIUM CHLORIDE|MAGNESIUM ACETATE / POTASSIUM ACETATE / SODIUM CHLORIDE
C2929601|T121|1008702|RXNORM|PYRIDOXINE / VITAMIN B 12|PYRIDOXINE / VITAMIN B 12
C2929604|T121|1008705|RXNORM|DIPHENHYDRAMINE / PRAMOXINE|DIPHENHYDRAMINE / PRAMOXINE
C2929603|T121|1008704|RXNORM|DOCUSATE / SENNOSIDE B|DOCUSATE / SENNOSIDE B
C2929606|T121|1008707|RXNORM|BISMUTH CHLORIDE OXIDE / PREDNISOLONE / ZINC OXIDE|BISMUTH CHLORIDE OXIDE / PREDNISOLONE / ZINC OXIDE
C2929605|T121|1008706|RXNORM|ACETAMINOPHEN / DEXCHLORPHENIRAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / DEXCHLORPHENIRAMINE / PSEUDOEPHEDRINE
C3264621|T121|1243041|RXNORM|IVACAFTOR|IVACAFTOR
C0054635|T121|20191|RXNORM|CARAMIPHEN|CARAMIPHEN
C0054636|T121|20192|RXNORM|CARAZOLOL|CARAZOLOL
C2193983|T121|812410|RXNORM|BROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN|BROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN
C1445298|T121|1352033|RXNORM|FAGOPYRUM ESCULENTUM EXTRACT|FAGOPYRUM ESCULENTUM EXTRACT
C0058134|T121|23162|RXNORM|DIHYDROXYALUMINUM AMINOACETATE|DIHYDROXYALUMINUM AMINOACETATE
C2728181|T129|1012134|RXNORM|SOUR CHERRY ALLERGENIC EXTRACT|SOUR CHERRY ALLERGENIC EXTRACT
C0772342|T121|237005|RXNORM|LEVOMETHADYL|LEVOMETHADYL
C0361275|T129|108542|RXNORM|MENINGITIS VACCINE|MENINGITIS VACCINE
C0318391|T005|1435396|RXNORM|HUMAN COXSACKIEVIRUS B3|HUMAN COXSACKIEVIRUS B3
C2080441|T121|812415|RXNORM|PHENAZOPYRIDINE / SULFAMETHOXAZOLE / TRIMETHOPRIM|PHENAZOPYRIDINE / SULFAMETHOXAZOLE / TRIMETHOPRIM
C3256271|T109|1305662|RXNORM|ROSA MOSCHATA OIL|ROSA MOSCHATA OIL
C3486699|T121|1310261|RXNORM|BOS TAURUS HYPOTHALAMUS PREPARATION|BOVINE HYPOTHALAMUS PREPARATION
C0011279|T121|3155|RXNORM|NORDAZEPAM|NORDAZEPAM
C0011276|T195|3154|RXNORM|DEMECLOCYCLINE|DEMECLOCYCLINE
C3282427|T121|1251312|RXNORM|ALGINIC ACID / CALCIUM CARBONATE / MAGNESIUM TRISILICATE / SODIUM BICARBONATE|ALGINIC ACID / CALCIUM CARBONATE / MAGNESIUM TRISILICATE / SODIUM BICARBONATE
C3695934|T129|1484986|RXNORM|WHITE WILLOW POLLEN EXTRACT|SALIX ALBA POLLEN EXTRACT
C3695935|T129|1484985|RXNORM|BULBOUS BUTTERCUP POLLEN EXTRACT|RANUNCULUS BULBOSUS POLLEN EXTRACT
C0000946|T121|149|RXNORM|ACEBUTOLOL|ACEBUTOLOL
C2827611|T129|1484983|RXNORM|BROADLEAF PLANTAIN POLLEN EXTRACT|GREATER PLANTAIN POLLEN EXTRACT
C3695936|T129|1484982|RXNORM|ASH POLLEN EXTRACT|FRAXINUS EXCELSIOR POLLEN EXTRACT
C3695937|T129|1484981|RXNORM|EUROPEAN BEECH POLLEN EXTRACT|FAGUS SYLVATICA POLLEN EXTRACT
C3256268|T109|1305665|RXNORM|RIBES NIGRUM SEED OIL|RIBES NIGRUM SEED OIL
C0054672|T121|20220|RXNORM|CARBINOXAMINE|CARBINOXAMINE
C0066351|T121|29844|RXNORM|METHYLENE DIPHOSPHONATE|METHYLENE DIPHOSPHONATE
C1541483|T129|591781|RXNORM|ECULIZUMAB|ECULIZUMAB
C1721194|T121|1544124|RXNORM|ECAMSULE|ECAMSULE
C0025912|T121|6929|RXNORM|MIANSERIN|MIANSERIN
C0772411|T121|1427056|RXNORM|POTATO STARCH|POTATO STARCH
C3848598|T121|1545042|RXNORM|VERBASCUM THAPSUS LEAF EXTRACT|VERBASCUM THAPSUS LEAF EXTRACT
C2722030|T129|894987|RXNORM|DOG SKIN EXTRACT|CANIS LUPUS FAMILIARIS DANDER EXTRACT
C0061559|T121|1311689|RXNORM|GLYCEROL FORMAL|GLYCEROL FORMAL
C3475127|T121|1311688|RXNORM|ZANTHOXYLUM ARMATUM VAR. ARMATUM FRUIT EXTRACT|ZANTHOXYLUM ARMATUM VAR. ARMATUM FRUIT EXTRACT
C3472974|T109|1311687|RXNORM|XANTHIUM STRUMARIUM FRUIT EXTRACT|XANTHIUM STRUMARIUM FRUIT EXTRACT
C3488979|T121|1311686|RXNORM|VITEX TRIFOLIA FRUIT EXTRACT|VITEX TRIFOLIA FRUIT EXTRACT
C3256741|T121|1311685|RXNORM|VACCINIUM MYRTILLUS FRUITING TOP EXTRACT|VACCINIUM MYRTILLUS FRUITING TOP EXTRACT
C3256562|T121|1311684|RXNORM|TETRADIUM RUTICARPUM FRUIT EXTRACT|TETRADIUM RUTICARPUM FRUIT EXTRACT
C3256561|T121|1311683|RXNORM|TERMINALIA CHEBULA FRUIT EXTRACT|TERMINALIA CHEBULA FRUIT EXTRACT
C3485017|T121|1311682|RXNORM|STAR ANISE FRUIT EXTRACT|STAR ANISE FRUIT EXTRACT
C3488420|T121|1311681|RXNORM|SCUTELLARIA LATERIFLORA TOP EXTRACT|SCUTELLARIA LATERIFLORA TOP EXTRACT
C3864835|T109|1596767|RXNORM|CYMBOPOGON CITRATUS WHOLE EXTRACT|CYMBOPOGON CITRATUS WHOLE EXTRACT
C3857964|T109|1551421|RXNORM|ETHYL PYRROLIDONE|ETHYL PYRROLIDONE
C0058056|T121|23088|RXNORM|DIHYDROCODEINE|DIHYDROCODEINE
C3666507|T121|1437222|RXNORM|QUERCUS MARILANDICA POLLEN EXTRACT|QUERCUS MARILANDICA POLLEN EXTRACT
C3864834|T129|1596768|RXNORM|ISOMERIZED SAFFLOWER ACID|ISOMERIZED SAFFLOWER ACID
C2928554|T121|1007638|RXNORM|CAMPHOR / CAPSICUM EXTRACT / METHYL SALICYLATE|CAMPHOR / CAPSICUM EXTRACT / METHYL SALICYLATE
C2928555|T121|1007639|RXNORM|ECHINACEA ROOT EXTRACT / GOLDEN SEAL ROOT|ECHINACEA ROOT EXTRACT / GOLDEN SEAL ROOT
C3857963|T121|1551422|RXNORM|NUPHAR JAPONICA ROOT EXTRACT|NUPHAR JAPONICA ROOT EXTRACT
C2928547|T121|1007630|RXNORM|CALCIUM PHOSPHATE / MAGNESIUM CARBONATE / POTASSIUM CHLORIDE|CALCIUM PHOSPHATE / MAGNESIUM CARBONATE / POTASSIUM CHLORIDE
C2928548|T121|1007631|RXNORM|ALUMINUM HYDROXIDE / MAGNESIUM TRISILICATE / SODIUM BICARBONATE|ALUMINUM HYDROXIDE / MAGNESIUM TRISILICATE / SODIUM BICARBONATE
C2928550|T121|1007633|RXNORM|DIHYDROERGOCRISTINE / LOMIFYLLINE|DIHYDROERGOCRISTINE / LOMIFYLLINE
C2016176|T121|1007634|RXNORM|BROMHEXINE / OXYTETRACYCLINE|BROMHEXINE / OXYTETRACYCLINE
C2928551|T121|1007635|RXNORM|BENZOCAINE / CHLORAMPHENICOL|BENZOCAINE / CHLORAMPHENICOL
C2928552|T121|1007636|RXNORM|BENZALKONIUM / BORIC ACID|BENZALKONIUM / BORIC ACID
C2946033|T121|1038763|RXNORM|BENZALKONIUM / BENZETHONIUM|BENZALKONIUM / BENZETHONIUM
C1690432|T129|993449|RXNORM|DENOSUMAB|DENOSUMAB
C0065517|T197|29155|RXNORM|MAGNESIUM CARBONATE|MAGNESIUM CARBONATE
C0065512|T197|29151|RXNORM|MAGALDRATE|MAGALDRATE
C1875111|T121|691231|RXNORM|EPHEDRINE / PHENOBARBITAL|EPHEDRINE / PHENOBARBITAL
C1875112|T121|691232|RXNORM|EPHEDRINE / PHENOBARBITAL / POTASSIUM IODIDE / THEOPHYLLINE|EPHEDRINE / PHENOBARBITAL / POTASSIUM IODIDE / THEOPHYLLINE
C1875113|T121|691235|RXNORM|EPHEDRINE / SECOBARBITAL|EPHEDRINE / SECOBARBITAL
C1960128|T121|729581|RXNORM|LAMIVUDINE / STAVUDINE|LAMIVUDINE / STAVUDINE
C3499442|T121|1312084|RXNORM|YUCCA GLAUCA ROOT EXTRACT|YUCCA GLAUCA ROOT EXTRACT
C3499443|T121|1312085|RXNORM|CONVALLARIA MAJALIS BULB EXTRACT|CONVALLARIA MAJALIS BULB EXTRACT
C2343926|T121||RXNORM|NIACIN / SIMVASTATIN
C0032623|T122|8570|RXNORM|POLYVINYL ALCOHOL|POLYVINYL ALCOHOL
C0982156|T121|314623|RXNORM|FIBRINOGEN,I-125|FIBRINOGEN (125I)
C0072076|T121|34568|RXNORM|PROGABIDE|PROGABIDE
C2722020|T129|971849|RXNORM|LAMB ALLERGENIC EXTRACT|LAMB ALLERGENIC EXTRACT
C0045093|T121|12574|RXNORM|GEMCITABINE|GEMCITABINE
C3832722|T109|1539418|RXNORM|MAGNOLIA GRANDIFLORA LEAF EXTRACT|MAGNOLIA GRANDIFLORA LEAF EXTRACT
C3535656|T121|1369690|RXNORM|ZANTHOXYLUM BUNGEANUM WHOLE EXTRACT|ZANTHOXYLUM BUNGEANUM WHOLE EXTRACT
C0727050|T121|577312|RXNORM|MINERAL OIL, LIGHT|MINERAL OIL, LIGHT
C0961485|T121|298869|RXNORM|EPLERENONE|EPLERENONE
C0028027|T127|7405|RXNORM|NIACINAMIDE|NIACINAMIDE
C0028027|T127|7405|RXNORM|NIACINAMIDE|NIACINAMIDE
C2931926|T121|1193326|RXNORM|RUXOLITINIB|RUXOLITINIB
C0028017|T121|7402|RXNORM|NICLOSAMIDE|NICLOSAMIDE
C3832792|T121|1539636|RXNORM|TRIISOSTEARYL CITRATE|TRIISOSTEARYL CITRATE
C1301990|T121|687258|RXNORM|CLIOQUINOL / FLUMETHASONE|CLIOQUINOL / FLUMETHASONE
C1827451|T121|687259|RXNORM|CLIOQUINOL / FLUOCINOLONE|CLIOQUINOL / FLUOCINOLONE
C0383429|T129|117055|RXNORM|ALEMTUZUMAB|ALEMTUZUMAB
C0049579|T121|16054|RXNORM|KINETIN|KINETIN
C0054094|T121|19737|RXNORM|BROMFENAC|BROMFENAC
C0054094|T121|19737|RXNORM|BROMFENAC|BROMFENAC
C3848523|T196|1546434|RXNORM|RUBIDIUM CATION RB-82|RUBIDIUM CATION RB-82
C3832723|T109|1539419|RXNORM|PRUNUS X YEDOENSIS LEAF EXTRACT|PRUNUS X YEDOENSIS LEAF EXTRACT
C0118538|T130|1421151|RXNORM|GADOTERATE MEGLUMINE|GADOTERATE MEGLUMINE
C1533316|T121|1421150|RXNORM|CALCIUM MALATE|CALCIUM MALATE
C3832791|T168|1539635|RXNORM|PASSIFLORA EDULIS FRUIT JUICE|PASSIFLORA EDULIS FRUIT JUICE
C0024730|T121|6628|RXNORM|MANNITOL|MANNITOL
C0024730|T121|6628|RXNORM|MANNITOL|MANNITOL
C0024730|T121|6628|RXNORM|MANNITOL|MANNITOL
C3665153|T121|1435391|RXNORM|GELIDIUM CARTILAGINEUM EXTRACT|GELIDIUM CARTILAGINEUM EXTRACT
C2057752|T121|817117|RXNORM|KETOTIFEN / THEOPHYLLINE|KETOTIFEN / THEOPHYLLINE
C0024706|T196|6623|RXNORM|MANGANESE|MANGANESE
C3700884|T122|1486796|RXNORM|BUTYLOCTYL BENZOATE|BUTYLOCTYL BENZOATE
C2194025|T121|812323|RXNORM|MAGNESIUM CARBONATE / MAGNESIUM OXIDE|MAGNESIUM CARBONATE / MAGNESIUM OXIDE
C0215278|T121|69440|RXNORM|POLICOSANOL|POLICOSANOL
C3848526|T196|1546430|RXNORM|THALLIUM CATION TL-201 (1+)|THALLIUM CATION TL-201 (1+)
C1873969|T121|689584|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE
C2006131|T121|1007721|RXNORM|CALCIUM CHLORIDE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE|CALCIUM CHLORIDE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE
C1873967|T121|689582|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|ACETAMINOPHEN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C1873968|T121|689583|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE
C1873965|T121|689580|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE|ACETAMINOPHEN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE
C3498011|T121|1313689|RXNORM|SOLIDAGO CANADENSIS WHOLE EXTRACT|SOLIDAGO CANADENSIS WHOLE EXTRACT
C3497910|T121|1313688|RXNORM|MOSCHUS MOSCHIFERUS WHOLE EXTRACT|MOSCHUS MOSCHIFERUS WHOLE EXTRACT
C2709768|T129|854964|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 5 VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 5 VACCINE
C0146010|T121|57257|RXNORM|TIXOCORTOL|TIXOCORTOL
C3267306|T121|1313685|RXNORM|STEVIA REBAUDIANA WHOLE EXTRACT|STEVIA REBAUDIANA WHOLE EXTRACT
C0754647|T121|228783|RXNORM|FROVATRIPTAN|FROVATRIPTAN
C3282140|T121|1313686|RXNORM|SAPONARIA OFFICINALIS WHOLE EXTRACT|SAPONARIA OFFICINALIS WHOLE EXTRACT
C3857955|T121|1551627|RXNORM|STEARETH-12|STEARETH-12
C0874052|T121|260025|RXNORM|ECHINACEA PURPUREA EXTRACT|ECHINACEA PURPUREA EXTRACT
C0053881|T121|19551|RXNORM|PEMIROLAST|PEMIROLAST
C0054257|T121|19882|RXNORM|BUTHIAZIDE|BUTHIAZIDE
C0053882|T195|19552|RXNORM|CEFPROZIL|CEFPROZIL
C0054259|T121|19884|RXNORM|BUTOCONAZOLE|BUTOCONAZOLE
C0540623|T121|141366|RXNORM|NARATRIPTAN|NARATRIPTAN
C2980883|T129|1094116|RXNORM|CREEPING BENTGRASS POLLEN EXTRACT|AGROSTIS STOLONIFERA POLLEN EXTRACT
C3848605|T109|1544575|RXNORM|DILAURYLDIMONIUM CHLORIDE|DILAURYLDIMONIUM CHLORIDE
C3832794|T109|1539638|RXNORM|2-AMINO-2-ETHYL-1,3-PROPANEDIOL|2-AMINO-2-ETHYL-1,3-PROPANEDIOL
C0051482|T121|1544577|RXNORM|ALFAXOLONE|ALFAXALONE
C2741590|T129|901511|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP Y OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|NEISSERIA MENINGITIDIS SEROGROUP Y OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C0006972|T121|2011|RXNORM|CARBAZOCHROME|CARBAZOCHROME
C0017237|T122|4716|RXNORM|GELATIN|GELATIN
C0068922|T121|31930|RXNORM|NOMEGESTROL|NOMEGESTROL
C0216194|T121|69627|RXNORM|TEA TREE OIL|TEA TREE OIL
C3154622|T121|1306096|RXNORM|ALUMINUM ZIRCONIUM OCTACHLOROHYDREX GLY|ALUMINUM ZIRCONIUM OCTACHLOROHYDREX GLY
C0017245|T121|4719|RXNORM|GEMFIBROZIL|GEMFIBROZIL
C2954886|T109|1306094|RXNORM|CURCUMA XANTHORRHIZA OIL|CURCUMA ZANTHORRHIZA OIL
C3256645|T109|1306095|RXNORM|POMEGRANATE SEED OIL|POMEGRANATE SEED OIL
C1873978|T121|689775|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / GUAIFENESIN|ACETAMINOPHEN / DEXTROMETHORPHAN / GUAIFENESIN
C2037255|T121|817112|RXNORM|ALPRAZOLAM / SULPIRIDE|ALPRAZOLAM / SULPIRIDE
C2928996|T121|1008088|RXNORM|BORIC ACID / OLEATE|BORIC ACID / OLEATE
C2928994|T121|1008086|RXNORM|GLYCOPYRROLATE / NEOSTIGMINE|GLYCOPYRROLATE / NEOSTIGMINE
C2928995|T121|1008087|RXNORM|LINOLEATE / SUNFLOWER SEED OIL|LINOLEATE / SUNFLOWER OIL
C2928992|T121|1008084|RXNORM|CHROMIUM PICOLINATE / LEVOCARNITINE|CHROMIUM PICOLINATE / LEVOCARNITINE
C2928993|T121|1008085|RXNORM|HEPARINOIDS / SALICYLIC ACID|HEPARINOIDS / SALICYLIC ACID
C2928990|T121|1008082|RXNORM|TERBUTALINE / THEOPHYLLINE|TERBUTALINE / THEOPHYLLINE
C2928991|T121|1008083|RXNORM|ACETAMINOPHEN / LORATADINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / LORATADINE / PSEUDOEPHEDRINE
C2928989|T121|1008080|RXNORM|ASPIRIN / METHYLPREDNISOLONE|ASPIRIN / METHYLPREDNISOLONE
C2193826|T121|1008081|RXNORM|AMBROXOL / AMOXICILLIN|AMBROXOL / AMOXICILLIN
C0013360|T121|3714|RXNORM|DYPHYLLINE|DYPHYLLINE
C1445730|T121|466496|RXNORM|COAL TAR / SALICYLIC ACID / SULFUR|COAL TAR / SALICYLIC ACID / SULFUR
C1445442|T129|968413|RXNORM|TRICHOPHYTON RUBRUM ALLERGENIC EXTRACT|TRICHOPHYTON RUBRUM ALLERGENIC EXTRACT
C3651743|T122|1429395|RXNORM|POLYQUATERNIUM-10 (125 MPA.S AT 2%)|POLYQUATERNIUM-10 (125 MPA.S AT 2%)
C2949346|T121|1046422|RXNORM|CALCIUM GLYCEROPHOSPHATE / MONOFLUOROPHOSPHATE / PYRIDOXINE|CALCIUM GLYCEROPHOSPHATE / MONOFLUOROPHOSPHATE / PYRIDOXINE
C2701568|T129|852404|RXNORM|STEMPHYLIUM EXTRACT|STEMPHYLIUM EXTRACT
C1445344|T121|1355405|RXNORM|ORIGANUM MAJORANA EXTRACT|ORIGANUM MAJORANA EXTRACT
C3663501|T121|1433190|RXNORM|VERNONIA APPENDICULATA LEAF EXTRACT|VERNONIA APPENDICULATA LEAF EXTRACT
C3663502|T121|1433191|RXNORM|CYPERUS ESCULENTUS LEAF EXTRACT|CYPERUS ESCULENTUS LEAF EXTRACT
C2929783|T121|1008886|RXNORM|MEPROBAMATE / TRIHEXYPHENIDYL|MEPROBAMATE / TRIHEXYPHENIDYL
C2929784|T121|1008887|RXNORM|ATROPINE / NITROGLYCERIN / THEOBROMINE|ATROPINE / NITROGLYCERIN / THEOBROMINE
C2930759|T121|1008884|RXNORM|DIETHYLAMINE SALICYLATE / FLUFENAMIC ACID / MYRTECAINE|DIETHYLAMINE SALICYLATE / FLUFENAMIC ACID / MYRTECAINE
C2929782|T121|1008885|RXNORM|FLUFENAMIC ACID / GLYCOL SALICYLATE / HEPARINOIDS|FLUFENAMIC ACID / GLYCOL SALICYLATE / HEPARINOIDS
C2929780|T121|1008882|RXNORM|AMERICAN COCKROACH ALLERGENIC EXTRACT / GERMAN COCKROACH ALLERGENIC EXTRACT|AMERICAN COCKROACH ALLERGENIC EXTRACT / GERMAN COCKROACH ALLERGENIC EXTRACT
C2929781|T121|1008883|RXNORM|HEPARINOIDS / LAURETH-9|HEPARINOIDS / POLIDOCANOL
C2929778|T121|1008880|RXNORM|GUAIACOLSULFONIC ACID / HYDROCODONE|GUAIACOLSULFONIC ACID / HYDROCODONE
C2929779|T121|1008881|RXNORM|IRON,PEPTONIZED / LIVER EXTRACT / VITAMIN B 12|IRON,PEPTONIZED / LIVER EXTRACT / VITAMIN B 12
C0017845|T121|4903|RXNORM|GLUTETHIMIDE|GLUTETHIMIDE
C2702431|T121|854130|RXNORM|PENICILLIUM CHRYSOGENUM VAR. CHRYSOGENUM EXTRACT|PENICILLIUM CHRYSOGENUM VAR. CHRYSOGENUM EXTRACT
C2929786|T121|1008889|RXNORM|CODEINE / PHENIRAMINE / PHENYLEPHRINE / SODIUM CITRATE|CODEINE / PHENIRAMINE / PHENYLEPHRINE / SODIUM CITRATE
C0947613|T121|1367117|RXNORM|STARCH, RICE|STARCH, RICE
C0788658|T121|1367110|RXNORM|POLYETHYLENE GLYCOL 1450|POLYETHYLENE GLYCOL 1450
C0912295|T116|1367111|RXNORM|NEOTAME|NEOTAME
C0018880|T196|5140|RXNORM|HELIUM|HELIUM
C0049104|T121|1367119|RXNORM|5-CHLORO-2-METHYL-4-ISOTHIAZOLIN-3-ONE|METHYLCHLOROISOTHIAZOLINONE
C3535689|T121|1368328|RXNORM|AMBROSIA PSILOSTACHYA TOP EXTRACT|AMBROSIA PSILOSTACHYA TOP EXTRACT
C2740815|T129|899770|RXNORM|MILLET SEED ALLERGENIC EXTRACT|PANICUM MILIACEUM ALLERGENIC EXTRACT
C3695983|T122|1482914|RXNORM|HYDROXYPROPYLCOCOATE PEG-8 DIMETHICONE|HYDROXYPROPYLCOCOATE PEG-8 DIMETHICONE
C0055332|T121|20762|RXNORM|CHLORAMINE-T|TOSYLCHLORAMIDE SODIUM
C3535692|T121|1368325|RXNORM|TEUCRIUM MARUM TOP EXTRACT|TEUCRIUM MARUM TOP EXTRACT
C3535691|T121|1368326|RXNORM|VERBASCUM DENSIFLORUM FLOWERING TOP EXTRACT|VERBASCUM DENSIFLORUM FLOWERING TOP EXTRACT
C3535690|T121|1368327|RXNORM|GALPHIMIA GLAUCA WHOLE EXTRACT|GALPHIMIA GLAUCA WHOLE EXTRACT
C0008196|T121|2358|RXNORM|AMINO ACIDS 5.4%|CHLORHEXIDINE
C0008196|T121|2358|RXNORM|AMINO ACIDS 4%|CHLORHEXIDINE
C0008196|T121|2358|RXNORM|AMINO ACIDS 15%|CHLORHEXIDINE
C0008196|T121|2358|RXNORM|AMINO ACIDS 11.4%|CHLORHEXIDINE
C3695953|T109|1484502|RXNORM|VANILLA PLANIFOLIA OIL|VANILLA PLANIFOLIA OIL
C1611331|T121|1309703|RXNORM|MALVIN|MALVIN
C3486861|T121|1309702|RXNORM|AVENA SATIVA FLOWERING TOP EXTRACT|AVENA SATIVA FLOWERING TOP EXTRACT
C3488212|T121|1309701|RXNORM|JATROPHA CURCAS SEED EXTRACT|JATROPHA CURCAS SEED EXTRACT
C3488211|T121|1309706|RXNORM|IPOMOEA PURGA ROOT EXTRACT|IPOMOEA PURGA ROOT EXTRACT
C0008196|T121|2358|RXNORM|AMINO ACIDS 5%|CHLORHEXIDINE
C3488213|T121|1309704|RXNORM|JUSTICIA ADHATODA LEAF EXTRACT|JUSTICIA ADHATODA LEAF EXTRACT
C2726765|T121|885183|RXNORM|AGKISTRODON PISCIVORUS ANTIVENIN|AGKISTRODON PISCIVORUS ANTIVENIN
C2726767|T121|885185|RXNORM|CROTALUS ADAMANTEUS ANTIVENIN|CROTALUS ADAMANTEUS ANTIVENIN
C0369723|T195|618425|RXNORM|NALIDIXATE|NALIDIXATE
C2726769|T121|885187|RXNORM|CROTALUS ATROX ANTIVENIN|CROTALUS ATROX ANTIVENIN
C2726771|T121|885189|RXNORM|CROTALUS SCUTULATUS ANTIVENIN|CROTALUS SCUTULATUS ANTIVENIN
C2980749|T121|1426392|RXNORM|DIETHYLAMINO HYDROXYBENZOYL HEXYL BENZOATE|DIETHYLAMINO HYDROXYBENZOYL HEXYL BENZOATE
C3644409|T121|1424863|RXNORM|ADANSONIA DIGITATA FRUIT EXTRACT|ADANSONIA DIGITATA FRUIT EXTRACT
C3644410|T122|1424864|RXNORM|DIMETHYLSILANOL HYALURONATE|DIMETHYLSILANOL HYALURONATE
C3257517|T109|1424865|RXNORM|APPLE EXTRACT|APPLE EXTRACT
C0724441|T121|220982|RXNORM|YOHIMBINE|YOHIMBINE
C3644412|T122|1424868|RXNORM|CHOLESTERYL-BEHENYL-OCTYLDODECYL LAUROYL GLUTAMATE|CHOLESTERYL-BEHENYL-OCTYLDODECYL LAUROYL GLUTAMATE
C1138626|T121|1373895|RXNORM|COCOA EXTRACT|COCOA EXTRACT
C3859159|T121|1592262|RXNORM|PALM KERNEL GLYCERIDES|PALM KERNEL GLYCERIDES
C2701774|T129|852746|RXNORM|EASTERN SYCAMORE POLLEN EXTRACT|PLATANUS OCCIDENTALIS POLLEN EXTRACT
C0072393|T123|34822|RXNORM|VITAMIN K-DEPENDENT PROTEIN S|PROTEIN S
C0654360|T121|186010|RXNORM|AMBROXOL-THEOPHYLLINE-7-ACETATE|AMBROXOL-THEOPHYLLINE-7-ACETATE
C0027373|T121|7247|RXNORM|NAPHAZOLINE|NAPHAZOLINE
C0027373|T121|7247|RXNORM|NAPHAZOLINE|NAPHAZOLINE
C3190736|T121|1145062|RXNORM|ALUMINUM SULFATE / LIDOCAINE|ALUMINUM SULFATE / LIDOCAINE
C0288171|T121|83818|RXNORM|IRBESARTAN|IRBESARTAN
C0027360|T121|7243|RXNORM|NALTREXONE|NALTREXONE
C0027360|T121|7243|RXNORM|NALTREXONE|NALTREXONE
C0027358|T109|7242|RXNORM|NALOXONE|NALOXONE
C2702430|T129|967111|RXNORM|PENICILLIUM EXPANSUM EXTRACT|PENICILLIUM EXPANSUM EXTRACT
C0874078|T121|260051|RXNORM|WASP VENOM PROTEIN|WASP VENOM PROTEIN
C0874080|T121|260053|RXNORM|ELDERBERRY FRUIT|ELDERBERRY FRUIT
C0074732|T121|36685|RXNORM|SODIUM CARBONATE|SODIUM CARBONATE
C0288165|T121|83816|RXNORM|DELAVIRDINE|DELAVIRDINE
C2929922|T121|1009027|RXNORM|ACETAMINOPHEN / ANTIPYRINE / CAFFEINE|ACETAMINOPHEN / ANTIPYRINE / CAFFEINE
C2929921|T121|1009026|RXNORM|ALTERNARIA ALTERNATA ALLERGENIC EXTRACT / CLADOSPORIUM CLADOSPORIOIDES ALLERGENIC EXTRACT|ALTERNARIA ALTERNATA ALLERGENIC EXTRACT / CLADOSPORIUM CLADOSPORIOIDES ALLERGENIC EXTRACT
C2929920|T121|1009025|RXNORM|LIDOCAINE / TRIAMCINOLONE|LIDOCAINE / TRIAMCINOLONE
C2929919|T121|1009024|RXNORM|CHLORHEXIDINE / DEXPANTHENOL|CHLORHEXIDINE / DEXPANTHENOL
C2929918|T121|1009023|RXNORM|FOLIC ACID / NIACINAMIDE / ZINC OXIDE|FOLIC ACID / NIACINAMIDE / ZINC OXIDE
C2929917|T121|1009022|RXNORM|BEE POLLEN / GINSENG PREPARATION|BEE POLLEN / GINSENG PREPARATION
C2929916|T121|1009021|RXNORM|MILK THISTLE FRUIT / MILK THISTLE FRUIT EXTRACT|MILK THISTLE FRUIT / MILK THISTLE FRUIT EXTRACT
C2929915|T121|1009020|RXNORM|CALCIUM CARBONATE / CALCIUM GLUCONATE / VITAMIN D|CALCIUM CARBONATE / CALCIUM GLUCONATE / VITAMIN D
C3489015|T121|1311207|RXNORM|SUS SCROFA ARTERY PREPARATION|PORCINE ARTERY PREPARATION
C2929924|T121|1009029|RXNORM|CORIANDER EXTRACT / SENNOSIDES, USP|CORIANDER EXTRACT / SENNOSIDES, USP
C2929923|T121|1009028|RXNORM|ASCORBIC ACID / HYDROQUINONE|ASCORBIC ACID / HYDROQUINONE
C2929940|T121|1009045|RXNORM|FLORFENICOL / SULFACETAMIDE|FLORFENICOL / SULFACETAMIDE
C0025625|T121|6822|RXNORM|METHAPYRILENE|METHAPYRILENE
C0025627|T121|6823|RXNORM|METHAQUALONE|METHAQUALONE
C2927952|T121|1007029|RXNORM|DIBASIC POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC|DIBASIC POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE, MONOBASIC
C2927951|T121|1007028|RXNORM|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / TAURINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / TAURINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C0025631|T121|6826|RXNORM|METHAZOLAMIDE|METHAZOLAMIDE
C2929939|T121|1009044|RXNORM|CHOLESTYRAMINE RESIN / DICLOFENAC|CHOLESTYRAMINE RESIN / DICLOFENAC
C2927948|T121|1007025|RXNORM|ALUMINUM ACETOTARTRATE / NONOXYNOL-9|ALUMINUM ACETOTARTRATE / NONOXYNOL-9
C2927950|T121|1007027|RXNORM|RHUBARB PREPARATION / SODIUM BICARBONATE|RHUBARB PREPARATION / SODIUM BICARBONATE
C2927944|T121|1007021|RXNORM|DIHYDRALAZINE / OXPRENOLOL|DIHYDRALAZINE / OXPRENOLOL
C2929942|T121|1009047|RXNORM|EVENING PRIMROSE EXTRACT / GAMMA-LINOLENATE / LINOLEATE|EVENING PRIMROSE EXTRACT / GAMMA-LINOLENATE / LINOLEATE
C2927946|T121|1007023|RXNORM|COAL TAR / LACTATE / SALICYLIC ACID|COAL TAR / LACTATE / SALICYLIC ACID
C2929941|T121|1009046|RXNORM|NEOMYCIN / PROPIONIC ACID|NEOMYCIN / PROPIONIC ACID
C2948090|T121|1426391|RXNORM|DIACETYL BENZOYL LATHYROL|DIACETYL BENZOYL LATHYROL
C1875567|T121|689343|RXNORM|NYSTATIN / OXYTETRACYCLINE|NYSTATIN / OXYTETRACYCLINE
C0304147|T109|1309372|RXNORM|OIL OF PATCHOULI|OIL OF PATCHOULI
C2929936|T121|1009041|RXNORM|BENZOCAINE / CALAMINE|BENZOCAINE / CALAMINE
C3256432|T121|1309370|RXNORM|PLANTAGO LANCEOLATA LEAF EXTRACT|PLANTAGO LANCEOLATA LEAF EXTRACT
C0304113|T109|1309371|RXNORM|ROSE OIL|ROSE OIL
C0172379|T109|1309376|RXNORM|CITRONELLA OIL|CITRONELLA OIL
C1533371|T168|1309377|RXNORM|LIME OIL|LIME OIL
C1656676|T109|1309374|RXNORM|PALMAROSA OIL|PALMAROSA OIL
C2929935|T121|1009040|RXNORM|BILBERRY EXTRACT / GRAPE SEED|BILBERRY EXTRACT / GRAPE SEED
C0950483|T121|288331|RXNORM|DICOBALT EDETATE|DICOBALT EDETATE
C0003438|T121|1009|RXNORM|DIPHTHERIA TOXOID VACCINE, INACTIVATED / H INFLUENZAE TYPE B / PERTUSSIS, WHOLE CELL / TETANUS TOXOID VACCINE, INACTIVATED|ANTITHROMBIN III
C0982015|T197|314494|RXNORM|AMMONIUM SILICOFLUORIDE|AMMONIUM SILICOFLUORIDE
C2929937|T121|1009042|RXNORM|BETA CAROTENE / BILBERRY EXTRACT|BETA CAROTENE / BILBERRY EXTRACT
C3854118|T121|1593854|RXNORM|SHEEP WOOL PREPARATION|SHEEP WOOL PREPARATION
C0136568|T121|54620|RXNORM|PHENOBARBITAL QUINIDINE|PHENOBARBITAL QUINIDINE
C3495447|T197|1311308|RXNORM|STRONTIUM CARBONATE PREPARATION|STRONTIUM CARBONATE PREPARATION
C0033567|T123|8814|RXNORM|EPOPROSTENOL|EPOPROSTENOL
C2729481|T129|895552|RXNORM|ALLSPICE ALLERGENIC EXTRACT|PIMENTA OFFICINALIS ALLERGENIC EXTRACT
C3486812|T121|1311302|RXNORM|ONONIS CAMPESTRIS EXTRACT|ONONIS SPINOSA WHOLE EXTRACT
C0070592|T121|33309|RXNORM|PHENSUXIMIDE|PHENSUXIMIDE
C3486776|T121|1311301|RXNORM|PORCINE HEART PREPARATION|PORCINE HEART PREPARATION
C1622989|T007|1311307|RXNORM|PEPTOSTREPTOCOCCUS ANAEROBIUS|PEPTOSTREPTOCOCCUS ANAEROBIUS
C3484495|T197|1311304|RXNORM|CALCIUM HEXAFLUOROSILICATE|CALCIUM HEXAFLUOROSILICATE
C3486299|T121|1311305|RXNORM|TARAXACUM OFFICINALE WHOLE EXTRACT|TARAXACUM OFFICINALE WHOLE EXTRACT
C2928211|T121|1007289|RXNORM|CALAMINE / DIMETHICONE / ZINC OXIDE|CALAMINE / DIMETHICONE / ZINC OXIDE
C2346990|T121|1326077|RXNORM|BELLIS PERENNIS EXTRACT|BELLIS PERENNIS EXTRACT
C2928203|T121|1007281|RXNORM|DOCUSATE / SORBITOL|DOCUSATE / SORBITOL
C2928205|T121|1007283|RXNORM|ECHINACEA ANGUSTIFOLIA ROOT EXTRACT / ECHINACEA PALLIDA ROOT EXTRACT|ECHINACEA ANGUSTIFOLIA ROOT EXTRACT / ECHINACEA PALLIDA ROOT EXTRACT
C2928204|T121|1007282|RXNORM|CYCLAMATE / SACCHARIN|CYCLAMATE / SACCHARIN
C2928207|T121|1007285|RXNORM|ERGOCALCIFEROL / VITAMIN A|ERGOCALCIFEROL / VITAMIN A
C2928206|T121|1007284|RXNORM|KELP PREPARATION / VITAMIN A|KELP PREPARATION / VITAMIN A
C2928209|T121|1007287|RXNORM|INSULIN, PROMPT ZINC, HUMAN / ULTRALENTE INSULIN, HUMAN|INSULIN, PROMPT ZINC, HUMAN / ULTRALENTE INSULIN, HUMAN
C2928208|T121|1007286|RXNORM|EPHEDRINE / ETHYLMORPHINE|EPHEDRINE / ETHYLMORPHINE
C0982404|T121|1426397|RXNORM|SORBITAN TRISTEARATE|SORBITAN TRISTEARATE
C3555503|T121|1376147|RXNORM|CAPRYLIC-CAPRIC-LINOLEIC TRIGLYCERIDE|CAPRYLIC-CAPRIC-LINOLEIC TRIGLYCERIDE
C3531439|T121|1366798|RXNORM|MICONAZOLE / TRICLOSAN|MICONAZOLE / TRICLOSAN
C3555502|T121|1376149|RXNORM|ALPHA-TOCOPHERYLQUINONE|ALPHA-TOCOPHERYLQUINONE
C0388013|T129|119246|RXNORM|RESPIRATORY SYNCYTIAL VIRUS IMMUNE GLOBULIN INTRAVENOUS|RESPIRATORY SYNCYTIAL VIRUS IMMUNE GLOBULIN INTRAVENOUS
C3486393|T121|1345677|RXNORM|RUMEX CRISPUS ROOT EXTRACT|RUMEX CRISPUS ROOT EXTRACT
C0378366|T121|114934|RXNORM|DESIRUDIN|DESIRUDIN
C2726147|T129|975763|RXNORM|DILL ALLERGENIC EXTRACT|ANETHUM GRAVEOLENS ALLERGENIC EXTRACT
C1444934|T121|465711|RXNORM|CIPROFLOXACIN / HYDROCORTISONE|CIPROFLOXACIN / HYDROCORTISONE
C3486693|T121|1345678|RXNORM|GALIUM APARINE EXTRACT|GALIUM APARINE EXTRACT
C1874897|T121|690085|RXNORM|CODEINE / GUAIFENESIN / PSEUDOEPHEDRINE / TRIPROLIDINE|CODEINE / GUAIFENESIN / PSEUDOEPHEDRINE / TRIPROLIDINE
C1533412|T122|1314379|RXNORM|POLOXAMER 124|POLOXAMER 124
C3834056|T109|1543081|RXNORM|CERTEARETH-100|CERTEARETH-100
C3715207|T109|1543082|RXNORM|BERGAMOT ORANGE EXTRACT|BERGAMOT ORANGE EXTRACT
C1874896|T121|690082|RXNORM|CODEINE / GUAIFENESIN / PHENYLEPHRINE|CODEINE / GUAIFENESIN / PHENYLEPHRINE
C0068443|T121|1314370|RXNORM|NARASIN|NARASIN
C1572727|T129|1314371|RXNORM|FANOLESOMAB|FANOLESOMAB
C1725176|T130|1314372|RXNORM|INDIUM IN-111 OXYQUINOLINE|INDIUM IN-111 OXYQUINOLINE
C1509666|T121|1314373|RXNORM|PALMITOYL OLIGOPEPTIDE|PALMITOYL OLIGOPEPTIDE
C1874901|T121|690089|RXNORM|CODEINE / PAPAVERINE|CODEINE / PAPAVERINE
C1874900|T121|690088|RXNORM|CODEINE / MENTHOL / PHENIRAMINE / PHENYLEPHRINE|CODEINE / MENTHOL / PHENIRAMINE / PHENYLEPHRINE
C1509637|T121|1314376|RXNORM|POLACRILIN|POLACRILIN
C3486664|T121|1309958|RXNORM|CAMELLIA SINENSIS FLOWER EXTRACT|CAMELLIA SINENSIS FLOWER EXTRACT
C3486665|T121|1309959|RXNORM|ALPINIA GALANGA LEAF EXTRACT|ALPINIA GALANGA LEAF EXTRACT
C3489380|T121|1309956|RXNORM|VETIVERIA ZIZANIOIDES ROOT EXTRACT|VETIVERIA ZIZANIOIDES ROOT EXTRACT
C0938478|T121|284153|RXNORM|MILK THISTLE FRUIT EXTRACT|MILK THISTLE FRUIT EXTRACT
C3486638|T121|1309954|RXNORM|ARISAEMA TRIPHYLLUM ROOT EXTRACT|ARISAEMA TRIPHYLLUM ROOT EXTRACT
C3486661|T121|1309955|RXNORM|VIBURNUM PRUNIFOLIUM BARK EXTRACT|VIBURNUM PRUNIFOLIUM BARK EXTRACT
C3486659|T121|1309952|RXNORM|VERONICA OFFICINALIS FLOWERING TOP EXTRACT|VERONICA OFFICINALIS FLOWERING TOP EXTRACT
C3282410|T121|1309953|RXNORM|PRUNUS SPECIOSA LEAF EXTRACT|PRUNUS SPECIOSA LEAF EXTRACT
C3486652|T121|1309950|RXNORM|ALETRIS FARINOSA ROOT EXTRACT|ALETRIS FARINOSA ROOT EXTRACT
C3486657|T121|1309951|RXNORM|ABRUS PRECATORIUS SEED EXTRACT|ABRUS PRECATORIUS SEED EXTRACT
C2740746|T130|899637|RXNORM|CARAWAY SEED ALLERGENIC EXTRACT|CARUS CARVI SEED ALLERGENIC EXTRACT
C0949647|T127|578285|RXNORM|TOCOTRIENOLS|TOCOTRIENOLS
C1875235|T121|692796|RXNORM|HELIUM / OXYGEN|HELIUM / OXYGEN
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C0037494|T197|9863|RXNORM|SODIUM CHLORIDE|SODIUM CHLORIDE
C1875224|T121|692794|RXNORM|GRAMICIDIN / NEOMYCIN / POLYMYXIN B|GRAMICIDIN / NEOMYCIN / POLYMYXIN B
C1875168|T121|692792|RXNORM|FOLLICLE STIMULATING HORMONE / LUTEINIZING HORMONE|FOLLICLE STIMULATING HORMONE / LUTEINIZING HORMONE
C2929481|T121|1008578|RXNORM|GLUCOSE / LACTATE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM CHLORIDE|GLUCOSE / LACTATE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM CHLORIDE
C2929482|T121|1008579|RXNORM|CARBINOXAMINE / PSEUDOEPHEDRINE / SCOPOLAMINE|CARBINOXAMINE / PSEUDOEPHEDRINE / SCOPOLAMINE
C2929479|T121|1008576|RXNORM|ACETYLCARNITINE / THIOCTATE|ACETYLCARNITINE / THIOCTATE
C2929480|T121|1008577|RXNORM|CLORAZEPATE / DOMPERIDONE|CLORAZEPATE / DOMPERIDONE
C2929477|T121|1008574|RXNORM|SODIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC|SODIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC
C2929477|T121|1008574|RXNORM|SODIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC|SODIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC
C2929477|T121|1008574|RXNORM|SODIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC|SODIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC
C2929478|T121|1008575|RXNORM|NOSCAPINE / POLYSORBATES / PROMETHAZINE|NOSCAPINE / POLYSORBATES / PROMETHAZINE
C2929475|T121|1008572|RXNORM|PSEUDOEPHEDRINE / SCOPOLAMINE|PSEUDOEPHEDRINE / SCOPOLAMINE
C2929476|T121|1008573|RXNORM|ALGINIC ACID / CALCIUM CARBONATE / MAGNESIUM CARBONATE|ALGINIC ACID / CALCIUM CARBONATE / MAGNESIUM CARBONATE
C2929473|T121|1008570|RXNORM|GLYCOLATE / PYRUVATE|GLYCOLATE / PYRUVATE
C1705480|T125|11149|RXNORM|VASOPRESSIN (USP)|VASOPRESSIN (USP)
C0076456|T121|38085|RXNORM|THIOCOLCHICOSIDE|THIOCOLCHICOSIDE
C1874668|T121|691032|RXNORM|CALCIUM IODIDE / CODEINE|CALCIUM IODIDE / CODEINE
C1875736|T121|690339|RXNORM|SALICYLIC ACID / ZINC PYRITHIONE|SALICYLIC ACID / ZINC PYRITHIONE
C1875735|T121|690337|RXNORM|SALICYLIC ACID / SODIUM THIOSULFATE|SALICYLIC ACID / SODIUM THIOSULFATE
C0005308|T125|1514|RXNORM|BETAMETHASONE|BETAMETHASONE
C0005308|T125|1514|RXNORM|BETAMETHASONE|BETAMETHASONE
C0005301|T121|1511|RXNORM|BETAHISTINE|BETAHISTINE
C0005304|T121|1512|RXNORM|BETAINE|BETAINE
C0771742|T121|236466|RXNORM|PYGEUM AFRICANUM PREPARATION|PYGEUM AFRICANUM PREPARATION
C0795680|T121|253210|RXNORM|ZINC, CHELATED|ZINC, CHELATED
C2929029|T121|1008122|RXNORM|HOPS EXTRACT / SKULLCAP PREPARATION / VALERIAN ROOT EXTRACT|HOPS EXTRACT / SKULLCAP PREPARATION / VALERIAN ROOT EXTRACT
C2348241|T121|1000082|RXNORM|ALCAFTADINE|ALCAFTADINE
C0813622|T123|258347|RXNORM|HYALURONAN|HYALURONAN
C3833362|T121|1541248|RXNORM|PEG-PPG-25-25 DIMETHICONE|PEG-PPG-25-25 DIMETHICONE
C2350656|T126|1011650|RXNORM|PEGLOTICASE|PEG-URICASE
C3255685|T109|1310092|RXNORM|HIPPOPHAE RHAMNOIDES FRUIT OIL|HIPPOPHAE RHAMNOIDES FRUIT OIL
C3275166|T109|1541240|RXNORM|GEUM URBANUM ROOT EXTRACT|GEUM URBANUM ROOT EXTRACT
C3486768|T121|1310095|RXNORM|PINUS SYLVESTRIS LEAFY TWIG|PINUS SYLVESTRIS LEAFY TWIG
C3812378|T121|1541242|RXNORM|QUERCUS ROBUR WHOLE EXTRACT|QUERCUS ROBUR WHOLE EXTRACT
C3833358|T121|1541243|RXNORM|RHEUM TANGUTICUM WHOLE EXTRACT|RHEUM TANGUTICUM WHOLE EXTRACT
C3833359|T121|1541244|RXNORM|SPHAGNUM SQUARROSUM EXTRACT|SPHAGNUM SQUARROSUM EXTRACT
C0061418|T123|1541246|RXNORM|GLUCOSE-6-PHOSPHATE|GLUCOSE-6-PHOSPHATE
C3833361|T121|1541247|RXNORM|ETHYL PERFLUOROISOBUTYL ETHER|ETHYL PERFLUOROISOBUTYL ETHER
C0772295|T121|236962|RXNORM|BENZOXONIUM|BENZOXONIUM
C1328724|T121|403712|RXNORM|MORINDA CITRIFOLIA EXTRACT|MORINDA CITRIFOLIA EXTRACT
C0064286|T121|28165|RXNORM|KERACYANIN|KERACYANIN
C0304554|T121|91263|RXNORM|ALOE EXTRACT|ALOE EXTRACT
C0041190|T121|10869|RXNORM|TROPICAMIDE|TROPICAMIDE
C0304561|T121|91266|RXNORM|RHUBARB PREPARATION|RHUBARB PREPARATION
C0304556|T121|91264|RXNORM|MALT SOUP EXTRACT|MALT SOUP EXTRACT
C0138666|T121|55175|RXNORM|PROPIVERINE|PROPIVERINE
C3475129|T121|1313746|RXNORM|DIPENTAERYTHRITYL HEXAHYDROXYSTEARATE|DIPENTAERYTHRITYL HEXAHYDROXYSTEARATE
C3255671|T121|1313747|RXNORM|ERICERUS PELA POLYCOSANOL|ERICERUS PELA POLYCOSANOL
C3256035|T121|1313740|RXNORM|DIETHYLHEXYL SUCCINATE|DIETHYLHEXYL SUCCINATE
C2699174|T168|1313217|RXNORM|CHICKEN LIVER PREPARATION|CHICKEN LIVER PREPARATION
C3474465|T121|1313742|RXNORM|DIMETHICONE PEG-7 ISOSTEARATE|DIMETHICONE PEG-7 ISOSTEARATE
C3257768|T121|1313743|RXNORM|DIMETHYL LAURAMINE|DIMETHYL LAURAMINE
C3498008|T121|1313218|RXNORM|BOS TAURUS CEREBELUM PREPARATION|BOS TAURUS CEREBELUM PREPARATION
C0163036|T109|1313219|RXNORM|1-HEXADECENE|1-HEXADECENE
C2717553|T109|1313748|RXNORM|ETHYL LEVULINATE|ETHYL LEVULINATE
C3473226|T121|1313749|RXNORM|ETHYLHEXYL ACETATE|ETHYLHEXYL ACETATE
C3530612|T121|1364948|RXNORM|HEPTYLUNDECYL HYDROXYSTEARATE|HEPTYLUNDECYL HYDROXYSTEARATE
C3530613|T121|1364949|RXNORM|LINOLEAMIDOPROPYL DIMETHYLAMINE|LINOLEAMIDOPROPYL DIMETHYLAMINE
C2929076|T121|1008169|RXNORM|HORSE CHESTNUT PREPARATION / MENTHOL|HORSE CHESTNUT PREPARATION / MENTHOL
C2929075|T121|1008168|RXNORM|UREA / VITAMIN E|UREA / VITAMIN E
C2929072|T121|1008165|RXNORM|ALLANTOIN / BENZALKONIUM / LIDOCAINE|ALLANTOIN / BENZALKONIUM / LIDOCAINE
C2929071|T121|1008164|RXNORM|BENZOXONIUM / LIDOCAINE|BENZOXONIUM / LIDOCAINE
C2929074|T121|1008167|RXNORM|CLONIXIN / SCOPOLAMINE|CLONIXIN / SCOPOLAMINE
C2929073|T121|1008166|RXNORM|RUSCOGENIN / TRIMEBUTINE|RUSCOGENIN / TRIMEBUTINE
C2929068|T121|1008161|RXNORM|PHENIRAMINE / PHENYLTOLOXAMINE / PSEUDOEPHEDRINE / PYRILAMINE|PHENIRAMINE / PHENYLTOLOXAMINE / PSEUDOEPHEDRINE / PYRILAMINE
C2929067|T121|1008160|RXNORM|GUINEA PIG HAIR EXTRACT / GUINEA PIG SKIN EXTRACT|GUINEA PIG HAIR EXTRACT / GUINEA PIG SKIN EXTRACT
C2929070|T121|1008163|RXNORM|ALVERINE / KARAYA GUM|ALVERINE / KARAYA GUM
C2929069|T121|1008162|RXNORM|DOMESTIC COW HAIR EXTRACT / DOMESTIC COW SKIN EXTRACT|DOMESTIC COW HAIR EXTRACT / DOMESTIC COW SKIN EXTRACT
C0123043|T121|51253|RXNORM|IBOPAMINE|IBOPAMINE
C0069810|T121|32680|RXNORM|OXYCHLOROSENE|OXYCHLOROSENE
C0022032|T130|5970|RXNORM|IOTHALAMATE|IOTHALAMATE
C0796545|T129|253453|RXNORM|PEGINTERFERON ALFA-2B|PEGINTERFERON ALFA-2B
C2756528|T129|968467|RXNORM|VERTICILLIUM ALBO-ATRUM EXTRACT|VERTICILLIUM ALBO-ATRUM EXTRACT
C0085319|T204|1322778|RXNORM|CRYPTOSPORIDIUM PARVUM|CRYPTOSPORIDIUM PARVUM
C0073578|T130|1535513|RXNORM|BASIC FUCHSIN|BASIC FUCHSIN
C0041165|T195|10864|RXNORM|TROLEANDOMYCIN|TROLEANDOMYCIN
C1869686|T195|1591901|RXNORM|CEFOVECIN|CEFOVECIN
C0795633|T125|253181|RXNORM|NPH INSULIN, HUMAN|INSULIN HUMAN, ISOPHANE
C1873946|T121|689556|RXNORM|ACETAMINOPHEN / ASPIRIN / PHENYLPROPANOLAMINE|ACETAMINOPHEN / ASPIRIN / PHENYLPROPANOLAMINE
C0795643|T197|253187|RXNORM|MANGANESE ASPARTATE|MANGANESE ASPARTATE
C3667759|T121|1440006|RXNORM|COD LIVER OIL / PETROLATUM|COD LIVER OIL / PETROLATUM
C2370007|T121|827167|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / METHSCOPOLAMINE|CHLORPHENIRAMINE / DEXTROMETHORPHAN / METHSCOPOLAMINE
C0005099|T121|1425|RXNORM|FD&C YELLOW #5|BENZYDAMINE
C0873046|T121|259385|RXNORM|GINSENG ROOT|GINSENG ROOT
C2194288|T121|821588|RXNORM|BROMHEXINE / METAPROTERENOL|BROMHEXINE / METAPROTERENOL
C0873041|T121|259380|RXNORM|VERBENA EXTRACT|VERBENA EXTRACT
C0873051|T121|259389|RXNORM|MILK THISTLE FRUIT|MILK THISTLE FRUIT
C0376892|T121|1373041|RXNORM|POLYHEXANIDE|POLIHEXANIDE
C3848603|T121|1544967|RXNORM|2-BUTYLOCTYL METHACRYLATE|2-BUTYLOCTYL METHACRYLATE
C1700874|T121|1242999|RXNORM|AXITINIB|AXITINIB
C1337299|T129|892484|RXNORM|STRAWBERRY ALLERGENIC EXTRACT|FRAGARIA ANANASSA ALLERGENIC EXTRACT
C3692845|T121|1442702|RXNORM|DICTAMNUS DASYCARPUS WHOLE EXTRACT|DICTAMNUS DASYCARPUS WHOLE EXTRACT
C3692844|T121|1442701|RXNORM|COMMIPHORA MYRRHA WHOLE EXTRACT|COMMIPHORA MYRRHA WHOLE EXTRACT
C0131956|T126|53553|RXNORM|NATTOKINASE|NATTOKINASE
C3486737|T121|1343597|RXNORM|CYPRIPEDIUM PARVIFOLUM ROOT EXTRACT|CYPRIPEDIUM PARVIFOLUM ROOT EXTRACT
C0069021|T121|32022|RXNORM|CATHINE|CATHINE
C0051033|T121|17205|RXNORM|AJMALICINE|AJMALICINE
C3245197|T121|1190559|RXNORM|ETHANOL / LIDOCAINE|ETHANOL / LIDOCAINE
C1563133|T121|597142|RXNORM|BRIMONIDINE / TIMOLOL|BRIMONIDINE / TIMOLOL
C0027599|T196|1311480|RXNORM|NEODYMIUM|NEODYMIUM
C0022154|T121|6011|RXNORM|ISOCARBOXAZID|ISOCARBOXAZID
C0297635|T121|88014|RXNORM|RIZATRIPTAN|RIZATRIPTAN
C0696679|T121|1309814|RXNORM|ASTRAGALUS PROPINQUUS ROOT EXTRACT|ASTRAGALUS PROPINQUUS ROOT EXTRACT
C3500452|T121|1314582|RXNORM|DRYOPTERIS CRASSIRHIZOMA WHOLE EXTRACT|DRYOPTERIS CRASSIRHIZOMA WHOLE EXTRACT
C3660765|T109|1489294|RXNORM|2-BENZYLHEPTANOL|2-BENZYLHEPTANOL
C3495133|T121|1368139|RXNORM|BRUGIA MALAYI PREPARATION|BRUGIA MALAYI PREPARATION
C3500451|T121|1314581|RXNORM|BOS TAURUS PEYER'S PATCH PREPARATION|BOS TAURUS PEYER'S PATCH PREPARATION
C1614561|T121|578377|RXNORM|POLYPODIUM LEUCOTOMOS|POLYPODIUM LEUCOTOMOS
C0075785|T109|1368135|RXNORM|BEEF TALLOW PREPARATION|BEEF TALLOW PREPARATION
C0052934|T121|1368134|RXNORM|BAKUCHIOL|BAKUCHIOL
C3257444|T121|1368137|RXNORM|BIOTINOYL TRIPEPTIDE-1|BIOTINOYL TRIPEPTIDE-1
C3488358|T121|1309810|RXNORM|THUJA OCCIDENTALIS LEAF EXTRACT|THUJA OCCIDENTALIS LEAF EXTRACT
C1612883|T109|1368131|RXNORM|ARACHIDYL ALCOHOL|ARACHIDYL ALCOHOL
C0912024|T121|1368130|RXNORM|APIGENIN|APIGENIN
C3643653|T121|1423803|RXNORM|GLYCERYL PHOSPHATE|GLYCERYL PHOSPHATE
C1612331|T109|1368132|RXNORM|ARACHIDYL GLUCOSIDE|ARACHIDYL GLUCOSIDE
C0725584|T121|221916|RXNORM|CHAMOMILE FLOWERS|CHAMOMILE FLOWERS
C0035179|T121|9260|RXNORM|RESERPINE|RESERPINE
C0771678|T121|236407|RXNORM|TRICARBAURINIUM|TRICARBAURINIUM
C0074926|T123|36853|RXNORM|SOY PROTEINS|SOY PROTEINS
C0040805|T121|10737|RXNORM|TRAZODONE|TRAZODONE
C0040778|T121|10734|RXNORM|TRANYLCYPROMINE|TRANYLCYPROMINE
C0040779|T121|10735|RXNORM|TRAPIDIL|TRAPIDIL
C0038179|T123|10046|RXNORM|STARCH|STARCH
C3535834|T197|1370660|RXNORM|TETRACHLOROAURATE|TETRACHLOROAURATE
C3535833|T109|1370661|RXNORM|URSOLATE|URSOLATE
C3535832|T121|1370662|RXNORM|N-(CARBONYL-METHOXYPOLYETHYLENE GLYCOL 2000)-1,2-DISTEAROYL-SN-GLYCERO-3-PHOSPHOETHANOLAMINE|N-(CARBONYL-METHOXYPOLYETHYLENE GLYCOL 2000)-1,2-DISTEAROYL-SN-GLYCERO-3-PHOSPHOETHANOLAMINE
C3535831|T121|1370663|RXNORM|2,5-DIMETHYLBENZENE-1-SULFONATE|2,5-DIMETHYLBENZENE-1-SULFONATE
C3535830|T109|1370664|RXNORM|ACRYLOYLDIMETHYLTAURATE|ACRYLOYLDIMETHYLTAURATE
C3535829|T121|1370665|RXNORM|ACRYLOYLDIMETHYLTAURATE-ACRYLAMIDE COPOLYMER|ACRYLOYLDIMETHYLTAURATE-ACRYLAMIDE COPOLYMER
C3535828|T121|1370666|RXNORM|ANISATE|ANISATE
C3535827|T121|1370667|RXNORM|OCTOXYNOL-2 ETHANE SULFONATE|OCTOXYNOL-2 ETHANE SULFONATE
C3535826|T109|1370669|RXNORM|POLARCRILLIN|POLARCRILLIN
C0061323|T121|25789|RXNORM|GLIMEPIRIDE|GLIMEPIRIDE
C2609578|T121|834769|RXNORM|CODEINE / DIPHENHYDRAMINE / PHENYLEPHRINE|CODEINE / DIPHENHYDRAMINE / PHENYLEPHRINE
C1719858|T121|645335|RXNORM|MAGNESIUM CARBONATE / SODIUM BICARBONATE|MAGNESIUM CARBONATE / SODIUM BICARBONATE
C1710622|T121|1317116|RXNORM|VELAFERMIN|VELAFERMIN
C3488590|T121|1426377|RXNORM|TAENIA SAGINATA PREPARATION|TAENIA SAGINATA PREPARATION
C1445764|T121|466530|RXNORM|ACETIC ACID / HYDROCORTISONE|ACETIC ACID / HYDROCORTISONE
C0073994|T125|36118|RXNORM|SALMON CALCITONIN|CALCITONIN (SALMON SYNTHETIC)
C0722704|T121|219314|RXNORM|POLYMYXIN B / TRIMETHOPRIM|POLYMYXIN B / TRIMETHOPRIM
C0722705|T121|219315|RXNORM|IRON POLYSACCHARIDE|IRON POLYSACCHARIDE
C2183064|T121|821542|RXNORM|CYPROHEPTADINE / DEXAMETHASONE|CYPROHEPTADINE / DEXAMETHASONE
C3818778|T109|1492036|RXNORM|DIMER DILINOLEYL DIMER DILINOLEATE|DIMER DILINOLEYL DIMER DILINOLEATE
C0717888|T121|214677|RXNORM|LIDOCAINE / OXYTETRACYCLINE|LIDOCAINE / OXYTETRACYCLINE
C2606637|T121|1306286|RXNORM|ELVITEGRAVIR|ELVITEGRAVIR
C3177235|T121|1306284|RXNORM|COBICISTAT|COBICISTAT
C2073899|T121|821019|RXNORM|CHLORPHENIRAMINE / SALICYLAMIDE|CHLORPHENIRAMINE / SALICYLAMIDE
C1699236|T125|618365|RXNORM|SYNTHETIC CONJUGATED ESTROGENS, B|SYNTHETIC CONJUGATED ESTROGENS, B
C2978390|T121|1088795|RXNORM|BLACK PEPPER PREPARATION / GUGGUL LIPIDS|BLACK PEPPER PREPARATION / GUGGUL LIPIDS
C0145055|T197|1431726|RXNORM|TECHNETIUM TC 99M EXAMETAZIME|TECHNETIUM (99MTC) EXAMETAZIME
C2978393|T121|1088798|RXNORM|CALCIUM CARBONATE / ERGOCALCIFEROL / SOY PROTEIN ISOLATE|CALCIUM CARBONATE / ERGOCALCIFEROL / SOY PROTEIN ISOLATE
C2726134|T129|1006258|RXNORM|APIOSPORA MONTAGNEI ALLERGENIC EXTRACT|APIOSPORA MONTAGNEI ALLERGENIC EXTRACT
C3179535|T121|1547099|RXNORM|SUVOREXANT|SUVOREXANT
C3256973|T130|1314215|RXNORM|TROLAMINE STEARATE|TROLAMINE STEARATE
C2927514|T129|1006250|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-CALIFORNIA-07-2009 X-181 (H1N1) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-CALIFORNIA-07-2009 X-181 (H1N1) STRAIN
C3658706|T129|1547545|RXNORM|PEMBROLIZUMAB|PEMBROLIZUMAB
C3488981|T109|1342493|RXNORM|GLYCYRRHIZA URALENSIS EXTRACT|GLYCYRRHIZA URALENSIS EXTRACT
C3486616|T121|1342490|RXNORM|CHENOPODIUM AMBROSIOIDES EXTRACT|CHENOPODIUM AMBROSIOIDES EXTRACT
C3486654|T121|1342491|RXNORM|BALLOTA FOETIDA EXTRACT|BALLOTA FOETIDA EXTRACT
C0614278|T121|164423|RXNORM|LOMIFYLLINE|LOMIFYLLINE
C0209368|T121|68149|RXNORM|MYCOPHENOLATE MOFETIL|MYCOPHENOLATE MOFETIL
C0012525|T121|3500|RXNORM|DIPHENOXYLATE|DIPHENOXYLATE
C0209366|T121|68147|RXNORM|CETRORELIX|CETRORELIX
C0057799|T121|22865|RXNORM|DIBROMPROPAMIDINE|DIBROMPROPAMIDINE
C2719424|T129|860168|RXNORM|ABOBOTULINUMTOXINA|ABOBOTULINUMTOXINA
C0009214|T121|2670|RXNORM|CODEINE|CODEINE
C0009214|T121|2670|RXNORM|CODEINE|CODEINE
C2344066|T129|797629|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP A CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE|NEISSERIA MENINGITIDIS SEROGROUP A CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE
C0215717|T121|69528|RXNORM|PARNAPARIN|PARNAPARIN
C2194151|T121|816530|RXNORM|CITICOLINE / NIMODIPINE|CITICOLINE / NIMODIPINE
C2929662|T121|1008763|RXNORM|CHLOPHEDIANOL / DEXCHLORPHENIRAMINE / PSEUDOEPHEDRINE|CHLOPHEDIANOL / DEXCHLORPHENIRAMINE / PSEUDOEPHEDRINE
C2929660|T121|1008761|RXNORM|CHOLECALCIFEROL / GLUCOSAMINE|CHOLECALCIFEROL / GLUCOSAMINE
C2929659|T121|1008760|RXNORM|BENZALKONIUM / MENTHOL|BENZALKONIUM / MENTHOL
C2929666|T121|1008767|RXNORM|FLUMETHIAZIDE / POTASSIUM CHLORIDE / RAUWOLFIA PREPARATION|FLUMETHIAZIDE / POTASSIUM CHLORIDE / RAUWOLFIA PREPARATION
C2929665|T121|1008766|RXNORM|CALCIUM CARBONATE / DOCOSAHEXAENOATE|CALCIUM CARBONATE / DOCOSAHEXAENOATE
C2929664|T121|1008765|RXNORM|ACEXAMIC ACID / CHLORHEXIDINE|ACEXAMIC ACID / CHLORHEXIDINE
C2929663|T121|1008764|RXNORM|AMYLMETACRESOL / DICHLOROBENZYL ALCOHOL / LIDOCAINE|AMYLMETACRESOL / DICHLOROBENZYL ALCOHOL / LIDOCAINE
C0010347|T121|2921|RXNORM|CROMOGLYCATE|CROMOGLYCATE
C2929668|T121|1008769|RXNORM|BENZOYL PEROXIDE / SALICYLIC ACID|BENZOYL PEROXIDE / SALICYLIC ACID
C2929667|T121|1008768|RXNORM|CHOLECALCIFEROL / VITAMIN K 2|CHOLECALCIFEROL / VITAMIN K 2
C1964492|T121|728498|RXNORM|DEXCHLORPHENIRAMINE / PHENYLEPHRINE|DEXCHLORPHENIRAMINE / PHENYLEPHRINE
C0019588|T123|5333|RXNORM|HISTAMINE|HISTAMINE
C0772283|T121|236953|RXNORM|GUARANA PREPARATION|GUARANA PREPARATION
C3535873|T121|1370610|RXNORM|METHYL COCOYL TAURATE|METHYL COCOYL TAURATE
C1337133|T121|1368869|RXNORM|DIPROPYLENE GLYCOL|DIPROPYLENE GLYCOL
C3486398|T109|1368868|RXNORM|SANGUISORBA OFFICINALIS TOP EXTRACT|SANGUISORBA OFFICINALIS TOP EXTRACT
C0358590|T121|106637|RXNORM|MISOPROSTOL / NAPROXEN|MISOPROSTOL / NAPROXEN
C0030773|T122|1368863|RXNORM|POLYETHYLENE GLYCOL 1000|POLYETHYLENE GLYCOL 1000
C0007289|T123|1368862|RXNORM|CARRAGEENAN|CARRAGEENAN
C0982351|T122|1368867|RXNORM|POLYSORBATE 60|POLYSORBATE 60
C3256556|T121|1368866|RXNORM|POLYETHYLENE GLYCOL 3000|POLYETHYLENE GLYCOL 3000
C3531583|T121|1367305|RXNORM|SORBUS AUCUPARIA FRUIT EXTRACT|SORBUS AUCUPARIA FRUIT EXTRACT
C0982313|T122|1368864|RXNORM|POLYETHYLENE GLYCOL 200|POLYETHYLENE GLYCOL 200
C1576805|T121|1364379|RXNORM|GLYCERYL STEARATE SE|GLYCERYL STEARATE SE
C1509280|T121|1364378|RXNORM|CETYL ACETATE|CETYL ACETATE
C3484452|T131|1310460|RXNORM|MICRURUS CORALLINUS VENOM|MICRURUS CORALLINUS VENOM
C3484453|T131|1310461|RXNORM|NAJA NAJA VENOM|NAJA NAJA VENOM
C3484456|T131|1310462|RXNORM|VIPERA BERUS VENOM|VIPERA BERUS VENOM
C0772357|T121|237020|RXNORM|WILD YAM EXTRACT|WILD YAM EXTRACT
C0772360|T121|237023|RXNORM|SPIKE LAVENDER OIL|SPIKE LAVENDER OIL
C1509211|T121|1364377|RXNORM|HYDROGENATED COCO-GLYCERIDES|HYDROGENATED COCO-GLYCERIDES
C1433693|T121|1364376|RXNORM|N-(3-(DIMETHYLAMINO)PROPYL)OCTADECANAMIDE|STEARAMIDOPROPYL DIMETHYLAMINE
C0772364|T121|237027|RXNORM|LOTEPREDNOL|LOTEPREDNOL
C0260195|T121|78678|RXNORM|RAUWOLFIA PREPARATION|RAUWOLFIA PREPARATION
C3818795|T122|1490690|RXNORM|POLYGLYCERYL-3 LAURATE|POLYGLYCERYL-3 LAURATE
C3818794|T122|1490691|RXNORM|METHYL HYDROGENATED ROSINATE|METHYL HYDROGENATED ROSINATE
C0076126|T121|37815|RXNORM|TERODILINE|TERODILINE
C0053787|T197|1311517|RXNORM|BISMUTH OXYCHLORIDE|BISMUTH OXYCHLORIDE
C0053291|T121|1311516|RXNORM|BENZYL CHLORIDE|BENZYL CHLORIDE
C3488943|T121|1311512|RXNORM|PFAFFIA PANICULATA ROOT EXTRACT|PFAFFIA PANICULATA ROOT EXTRACT
C3488942|T121|1311511|RXNORM|PEUCEDANUM OSTRUTHIUM LEAF EXTRACT|PEUCEDANUM OSTRUTHIUM LEAF EXTRACT
C3488941|T121|1311510|RXNORM|PETROSELINUM CRISPUM ROOT EXTRACT|PETROSELINUM CRISPUM ROOT EXTRACT
C0051750|T121|17813|RXNORM|AMPHETAMINIL|AMPHETAMINIL
C0304721|T121|91413|RXNORM|ADRENAL CORTEX EXTRACT|ADRENAL CORTEX EXTRACT
C3858057|T121|1551279|RXNORM|CAMPHOR / MENTHOL / TURPENTINE|CAMPHOR / MENTHOL / TURPENTINE
C2702329|T129|892565|RXNORM|ORANGE ALLERGENIC EXTRACT|CITRUS AURANTIUM DULCIS ALLERGENIC EXTRACT
C3652805|T121|1430892|RXNORM|FENOFIBRATE / SIMVASTATIN|FENOFIBRATE / SIMVASTATIN
C2928081|T121|1007159|RXNORM|PUMPKIN SEED EXTRACT / PYGEUM AFRICANUM PREPARATION / SAW PALMETTO EXTRACT|PUMPKIN SEED EXTRACT / PYGEUM AFRICANUM PREPARATION / SAW PALMETTO EXTRACT
C0072868|T121|1344799|RXNORM|QUINHYDRONE|QUINHYDRONE
C3495094|T121|1344798|RXNORM|LILIUM LANCIFOLIUM FLOWERING TOP EXTRACT|LILIUM LANCIFOLIUM FLOWERING TOP EXTRACT
C0007545|T195|2179|RXNORM|CEFATRIZINE|CEFATRIZINE
C2364569|T129|805573|RXNORM|ROTAVIRUS VACCINE, LIVE ATTENUATED, G1P[8] HUMAN 89-12 STRAIN|ROTAVIRUS VACCINE, LIVE ATTENUATED, G1P[8] HUMAN 89-12 STRAIN
C3256125|T109|1309207|RXNORM|BORAGO OFFICINALIS FLOWER EXTRACT|BORAGO OFFICINALIS FLOWER EXTRACT
C0771537|T121|236279|RXNORM|DEVIL'S CLAW PREPARATION|HARPAGOPHYTUM PROCUMBENS ROOT PREPARATION
C0061863|T121|26237|RXNORM|GRANISETRON|GRANISETRON
C0002658|T123|725|RXNORM|AMPHETAMINE|AMPHETAMINE
C0002644|T121|722|RXNORM|AMOXAPINE|AMOXAPINE
C0002645|T195|723|RXNORM|AMOXICILLIN|AMOXICILLIN
C0002645|T195|723|RXNORM|AMOXICILLIN|AMOXICILLIN
C0002641|T121|720|RXNORM|AMODIAQUINE|AMODIAQUINE
C3832875|T121|1539817|RXNORM|N-ALKYL DIMETHYL BENZYL AMMONIUM (C12-C18)|N-ALKYL DIMETHYL BENZYL AMMONIUM (C12-C18)
C3692729|T121|1442517|RXNORM|POLYQUATERNIUM-22 (4500 MPA.S)|POLYQUATERNIUM-22 (4500 MPA.S)
C3669287|T121|1442514|RXNORM|HUMAN HAIR PREPARATION|CRINIS CARBONISATUS
C0066335|T121|29829|RXNORM|METHYLBENZETHONIUM|METHYLBENZETHONIUM
C0066335|T121|29829|RXNORM|METHYLBENZETHONIUM|METHYLBENZETHONIUM
C3665568|T121|1442512|RXNORM|PELARGONIUM GRAVEOLENS WHOLE EXTRACT|PELARGONIUM GRAVEOLENS WHOLE EXTRACT
C3832872|T121|1539814|RXNORM|TRIMETHYL PENTAPHENYL TRISILOXANE|TRIMETHYL PENTAPHENYL TRISILOXANE
C3692725|T109|1442510|RXNORM|WHITE PEPPER OIL|WHITE PEPPER OIL
C3668955|T121|1442511|RXNORM|SALVIA OFFICINALIS WHOLE EXTRACT|SALVIA OFFICINALIS WHOLE EXTRACT
C0004011|T123|1167|RXNORM|ASPARTATE MAGNESIUM HYDROCHLORIDE|ASPARTATE MAGNESIUM HYDROCHLORIDE
C0054769|T121|20298|RXNORM|CARBOXYPOLYMETHYLENE|CARBOXYPOLYMETHYLENE
C0004015|T123|1169|RXNORM|ASPARTIC ACID|ASPARTIC ACID
C1450334|T121|1539813|RXNORM|SULFOBETAINE|SULFOBETAINE
C2928266|T121|1007344|RXNORM|TAURINE / VITAMIN B6|TAURINE / VITAMIN B6
C2928531|T121|1007613|RXNORM|ASPIRIN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE|ASPIRIN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE
C2928528|T121|1007610|RXNORM|NICKEL SULFATE / POTASSIUM BROMIDE / ZINC BROMIDE|NICKEL SULFATE / POTASSIUM BROMIDE / ZINC BROMIDE
C2928269|T121|1007347|RXNORM|CHLOROXYLENOL / PRAMOXINE / ZINC ACETATE|CHLOROXYLENOL / PRAMOXINE / ZINC ACETATE
C2928534|T121|1007616|RXNORM|FOLIC ACID / TEFERROL / VITAMIN B 12|FOLIC ACID / TEFERROL / VITAMIN B 12
C2928535|T121|1007617|RXNORM|CLIOQUINOL / FLUOCINONIDE|CLIOQUINOL / FLUOCINONIDE
C2928532|T121|1007614|RXNORM|IVERMECTIN / PRAZIQUANTEL|IVERMECTIN / PRAZIQUANTEL
C2928533|T121|1007615|RXNORM|CALCIUM CITRATE / MAGNESIUM OXIDE / VITAMIN E|CALCIUM CITRATE / MAGNESIUM OXIDE / VITAMIN E
C2928536|T121|1007618|RXNORM|CAMPHOR / CAPSAICIN / MENTHOL|CAMPHOR / CAPSAICIN / MENTHOL
C2928537|T121|1007619|RXNORM|AMPICILLIN / BROMHEXINE|AMPICILLIN / BROMHEXINE
C2928270|T121|1007348|RXNORM|ESTROGENS, ESTERIFIED (USP) / METHYLTESTOSTERONE|ESTROGENS, ESTERIFIED (USP) / METHYLTESTOSTERONE
C2928271|T121|1007349|RXNORM|GINSENG PREPARATION / ROYAL JELLY / VITAMIN B 12|GINSENG PREPARATION / ROYAL JELLY / VITAMIN B 12
C2033084|T121|818964|RXNORM|OXAZEPAM / PANCREATIN / SIMETHICONE|OXAZEPAM / PANCREATIN / SIMETHICONE
C0061387|T121|25842|RXNORM|GLUCONOLACTONE|GLUCONOLACTONE
C3464058|T109|1427231|RXNORM|CETETH-23|CETETH-23
C1874713|T121|691217|RXNORM|CARBINOXAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|CARBINOXAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C3833230|T109|1540871|RXNORM|ETHYL PERFLUOROBUTYL ETHER|ETHYL PERFLUOROBUTYL ETHER
C3848540|T121|1546397|RXNORM|SEA SNAIL PREPARATION|SEA SNAIL PREPARATION
C3282679|T025|1427138|RXNORM|FORESKIN KERATINOCYTE, NEONATAL|FORESKIN KERATINOCYTE, NEONATAL
C3264599|T121|1243019|RXNORM|LINAGLIPTIN / METFORMIN|LINAGLIPTIN / METFORMIN
C0070040|T121|1427237|RXNORM|PANTOLACTONE|PANTOLACTONE
C3700888|T109|1486759|RXNORM|KIWI SEED OIL|KIWI SEED OIL
C0458160|T168|1309208|RXNORM|GRAPE SEED OIL|GRAPE SEED OIL
C3555509|T109|1376088|RXNORM|OLEA EUROPAEA BARK EXTRACT|OLEA EUROPAEA BARK EXTRACT
C1516119|T121|495881|RXNORM|SORAFENIB|SORAFENIB
C0301248|T168|1309209|RXNORM|NUTMEG OIL|NUTMEG OIL
C0065533|T197|29170|RXNORM|MAGNESIUM TRISILICATE|MAGNESIUM TRISILICATE
C2722040|T129|862478|RXNORM|GREEN BELL PEPPER ALLERGENIC EXTRACT|GREEN BELL PEPPER ALLERGENIC EXTRACT
C3490258|T123|1545792|RXNORM|CHRYSOSPLENETIN|CHRYSOSPLENETIN
C3848589|T121|1545790|RXNORM|DAPHNE MEZEREUM WHOLE EXTRACT|DAPHNE MEZEREUM WHOLE EXTRACT
C3833235|T109|1540877|RXNORM|CHONDRUS CRISPUS CARRAGEENAN|CHONDRUS CRISPUS CARRAGEENAN
C3268295|T121|1248594|RXNORM|DOG HAIR EXTRACT / EUROPEAN HOUSE DUST MITE EXTRACT|DOG HAIR EXTRACT / EUROPEAN HOUSE DUST MITE EXTRACT
C0030883|T121|8004|RXNORM|PENTOBARBITAL|PENTOBARBITAL
C0032600|T121|8559|RXNORM|POLYSORBATE 20|POLYSORBATE 20
C0030873|T121|8001|RXNORM|PENTAZOCINE|PENTAZOCINE
C0256103|T126|76895|RXNORM|RETEPLASE|RETEPLASE
C3831895|T121|1538098|RXNORM|FLURALANER|FLURALANER
C1874400|T121|689615|RXNORM|ATROPINE / PREDNISOLONE|ATROPINE / PREDNISOLONE
C1874397|T121|689610|RXNORM|ATROPINE / MORPHINE|ATROPINE / MORPHINE
C1874398|T121|689611|RXNORM|ATROPINE / NEOSTIGMINE|ATROPINE / NEOSTIGMINE
C3538175|T121|1372309|RXNORM|C12-15 PARETH-7|C12-15 PARETH-7
C0051591|T121|17684|RXNORM|AMIDOLINE|AMIDOLINE
C3555496|T197|1376155|RXNORM|POTASSIUM TRIIODIDE|POTASSIUM TRIIODIDE
C0121772|T007|50937|RXNORM|HAEMOPHILUS INFLUENZAE TYPE B|HAEMOPHILUS INFLUENZAE TYPE B
C3249527|T121|1232660|RXNORM|BERMUDA GRASS SMUT EXTRACT / JOHNSON GRASS SMUT EXTRACT|BERMUDA GRASS SMUT EXTRACT / JOHNSON GRASS SMUT EXTRACT
C0054066|T121|19711|RXNORM|AMOXICILLIN / CLAVULANATE|AMOXICILLIN / CLAVULANATE
C3505485|T121|1358479|RXNORM|PLATOSTOMA CHINENSIS WHOLE EXTRACT|PLATOSTOMA CHINENSIS WHOLE EXTRACT
C0002006|T125|1312358|RXNORM|ALDOSTERONE|ALDOSTERONE
C0002865|T125|1312359|RXNORM|ANDROSTERONE|ANDROSTERONE
C0718010|T121|214788|RXNORM|POLYTHIAZIDE / RESERPINE|POLYTHIAZIDE / RESERPINE
C3505484|T121|1358478|RXNORM|IMPATIENS BALSAMINA LEAF EXTRACT|IMPATIENS BALSAMINA LEAF EXTRACT
C0718009|T121|214787|RXNORM|POLYTHIAZIDE / PRAZOSIN|POLYTHIAZIDE / PRAZOSIN
C3499503|T121|1312357|RXNORM|(C10-C30)ALKYL METHACRYLATE ESTER|(C10-C30)ALKYL METHACRYLATE ESTER
C0059752|T121|24506|RXNORM|VINPOCETINE|VINPOCETINE
C0724672|T121|221147|RXNORM|POLYETHYLENE GLYCOL 3350|POLYETHYLENE GLYCOL 3350
C0724672|T121|221147|RXNORM|POLYETHYLENE GLYCOL 3350|POLYETHYLENE GLYCOL 3350
C3832958|T109|1539998|RXNORM|BIXA ORELLANA SEED OIL|BIXA ORELLANA SEED OIL
C0041236|T126|10890|RXNORM|TRYPSIN|TRYPSIN
C3254757|T121|1370784|RXNORM|CHLORELLA VULGARIS EXTRACT|CHLORELLA VULGARIS EXTRACT
C0717446|T121|214254|RXNORM|ASPIRIN / MEPROBAMATE|ASPIRIN / MEPROBAMATE
C0717447|T121|214255|RXNORM|ASPIRIN / METHOCARBAMOL|ASPIRIN / METHOCARBAMOL
C0717448|T121|214256|RXNORM|ASPIRIN / OXYCODONE|ASPIRIN / OXYCODONE
C0717726|T195|214525|RXNORM|DOXORUBICIN LIPOSOME|DOXORUBICIN LIPOSOME
C0717442|T121|214250|RXNORM|ASPIRIN / CAFFEINE|ASPIRIN / CAFFEINE
C0717443|T121|214251|RXNORM|ASPIRIN / CARISOPRODOL|ASPIRIN / CARISOPRODOL
C0717721|T121|214520|RXNORM|DOCUSATE / PHENOLPHTHALEIN|DOCUSATE / PHENOLPHTHALEIN
C0717445|T121|214253|RXNORM|ASPIRIN / HYDROCODONE|ASPIRIN / HYDROCODONE
C3505483|T121|1358477|RXNORM|CISTUS INCANUS WHOLE EXTRACT|CISTUS INCANUS WHOLE EXTRACT
C0717450|T121|214258|RXNORM|ASPIRIN / PHENYLTOLOXAMINE|ASPIRIN / PHENYLTOLOXAMINE
C0717451|T121|214259|RXNORM|ASPIRIN / PSEUDOEPHEDRINE|ASPIRIN / PSEUDOEPHEDRINE
C0717729|T121|214528|RXNORM|DYPHYLLINE / GUAIFENESIN|DYPHYLLINE / GUAIFENESIN
C2194071|T121|816015|RXNORM|ACTIVATED CHARCOAL / SIMETHICONE|ACTIVATED CHARCOAL / SIMETHICONE
C0377265|T121|114477|RXNORM|LEVETIRACETAM|LEVETIRACETAM
C0068897|T121|31914|RXNORM|TIAGABINE|TIAGABINE
C3486814|T121|1347561|RXNORM|ONOSMODIUM VIRGINIANUM ROOT EXTRACT|ONOSMODIUM VIRGINIANUM ROOT EXTRACT
C2928256|T121|1007335|RXNORM|ALUMINUM ACETATE / BENZETHONIUM|ALUMINUM ACETATE / BENZETHONIUM
C0376337|T125|1537799|RXNORM|MELENGESTROL|MELENGESTROL
C0051556|T121|17652|RXNORM|AMCINONIDE|AMCINONIDE
C2928255|T121|1007334|RXNORM|HYDROCORTISONE / LACTATE|HYDROCORTISONE / LACTATE
C3488227|T121|1311365|RXNORM|SUS SCROFA INTERVERTEBRAL DISC PREPARATION|PORCINE INTERVERTEBRAL DISC PREPARATION
C2928759|T121|1007845|RXNORM|VIBRIO CHOLERAE SEROTYPE INABA / VIBRIO CHOLERAE SEROTYPE OGAWA|VIBRIO CHOLERAE SEROTYPE INABA / VIBRIO CHOLERAE SEROTYPE OGAWA
C3488005|T121|1347564|RXNORM|EUPHORBIA HIRTA EXTRACT|EUPHORBIA HIRTA EXTRACT
C2928758|T121|1007844|RXNORM|ECHINACEA PREPARATION / VITAMIN E / ZINC GLUCONATE|ECHINACEA PREPARATION / VITAMIN E / ZINC GLUCONATE
C1659023|T109|1492190|RXNORM|POLOXAMER 237|POLOXAMER 237
C2928253|T121|1007331|RXNORM|METRONIDAZOLE / SCOPOLAMINE|METRONIDAZOLE / SCOPOLAMINE
C0051241|T121|17381|RXNORM|APROBARBITAL|APROBARBITAL
C0051247|T121|17387|RXNORM|ALMINOPROFEN|ALMINOPROFEN
C1956280|T121|1482680|RXNORM|LULICONAZOLE|LULICONAZOLE
C2928252|T121|1007330|RXNORM|PENTAERYTHRITOL / PHENOBARBITAL|PENTAERYTHRITOL / PHENOBARBITAL
C3488085|T121|1309499|RXNORM|AGATHOSMA BETULINA LEAF EXTRACT|AGATHOSMA BETULINA LEAF EXTRACT
C3257672|T121|1309498|RXNORM|AESCULUS HIPPOCASTANUM LEAF EXTRACT|AESCULUS HIPPOCASTANUM LEAF EXTRACT
C2057683|T121|1007333|RXNORM|TETRACYCLINE / TROLEANDOMYCIN|TETRACYCLINE / TROLEANDOMYCIN
C3255711|T121|1309493|RXNORM|PERILLA FRUTESCENS LEAF EXTRACT|PERILLA FRUTESCENS LEAF EXTRACT
C3255845|T109|1309492|RXNORM|LEMON BALM OIL|MELISSA OFFICINALIS SEED OIL
C3255709|T109|1309491|RXNORM|PASSIFLORA INCARNATA SEED OIL|PASSIFLORA INCARNATA SEED OIL
C3255859|T109|1309490|RXNORM|PANAX GINSENG ROOT WATER EXTRACT|PANAX GINSENG ROOT WATER EXTRACT
C3486864|T121|1309497|RXNORM|AESCULUS HIPPOCASTANUM FLOWER EXTRACT|AESCULUS HIPPOCASTANUM FLOWER EXTRACT
C3486863|T121|1309496|RXNORM|ACTAEA SPICATA ROOT EXTRACT|ACTAEA SPICATA ROOT EXTRACT
C3488940|T121|1309495|RXNORM|PETIVERIA ALLIACEA ROOT EXTRACT|PETIVERIA ALLIACEA ROOT EXTRACT
C3256245|T109|1309494|RXNORM|PERSEA AMERICANA SEED BUTTER EXTRACT|AVOCADO SEED BUTTER
C2723772|T129|867361|RXNORM|WHEAT POLLEN EXTRACT|TRITICUM AESTIVUM POLLEN EXTRACT
C0030304|T126|7880|RXNORM|PANCREATIN|PANCREATIN
C0030310|T121|7883|RXNORM|PANCURONIUM|PANCURONIUM
C1509960|T121|477053|RXNORM|CINNAMON BARK|CINNAMON BARK
C0030314|T127|7886|RXNORM|PANGAMIC ACID|PANGAMIC ACID
C0047317|T121|1367170|RXNORM|METACRESOL|METACRESOL
C3256180|T109|1367171|RXNORM|QUARTERNIUM-15|QUARTERNIUM-15
C3531536|T109|1367173|RXNORM|CAPRYL-CAPRAMIDOPROPYL BETAINE|CAPRYL-CAPRAMIDOPROPYL BETAINE
C3531537|T121|1367174|RXNORM|TREPONEMIC SKIN CANKER PREPARATION, HUMAN|TREPONEMIC SKIN CANKER PREPARATION, HUMAN
C0003729|T121|1367175|RXNORM|ARBUTIN|ARBUTIN
C0004717|T195|1367176|RXNORM|BAMBERMYCINS|BAMBERMYCINS
C0007404|T121|1367177|RXNORM|CATECHIN|CATECHIN
C0007828|T196|1367178|RXNORM|CERIUM|CERIUM
C0009028|T121|1367179|RXNORM|CLOPIDOL|CLOPIDOL
C2826080|T122|1309724|RXNORM|METHACRYLIC ACID - METHYL METHACRYLATE COPOLYMER (1:2)|METHACRYLIC ACID - METHYL METHACRYLATE COPOLYMER (1:2)
C3488418|T121|1309727|RXNORM|ROSMARINUS OFFICINALIS FLOWERING TOP EXTRACT|ROSMARINUS OFFICINALIS FLOWERING TOP EXTRACT
C0071599|T122|1309726|RXNORM|POLYLACTIC ACID-POLYGLYCOLIC ACID COPOLYMER|POLYLACTIC ACID-POLYGLYCOLIC ACID COPOLYMER
C3256320|T122|1309721|RXNORM|METHACRYLIC ACID COPOLYMER|METHACRYLIC ACID COPOLYMER
C2698206|T122|1309720|RXNORM|METHACRYLIC ACID - METHYL METHACRYLATE COPOLYMER (1:1)|METHACRYLIC ACID - METHYL METHACRYLATE COPOLYMER (1:1)
C2938851|T121|1309723|RXNORM|INULA HELENIUM ROOT EXTRACT|INULA HELENIUM ROOT EXTRACT
C3488417|T121|1309722|RXNORM|ALCHEMILLA XANTHOCHLORA FLOWERING TOP EXTRACT|ALCHEMILLA XANTHOCHLORA FLOWERING TOP EXTRACT
C0000618|T121|103|RXNORM|MERCAPTOPURINE|MERCAPTOPURINE
C0593880|T121|153154|RXNORM|AMILORIDE / ATENOLOL / HYDROCHLOROTHIAZIDE|AMILORIDE / ATENOLOL / HYDROCHLOROTHIAZIDE
C3488423|T121|1309729|RXNORM|ARGENTINA ANSERINA FLOWERING TOP EXTRACT|POTENTILLA ANSERINA FLOWERING TOP EXTRACT
C0663655|T121|190521|RXNORM|ABACAVIR|ABACAVIR
C3695982|T109|1483080|RXNORM|SORBITYL LAURATE|SORBITYL LAURATE
C3487964|T121|1311360|RXNORM|SUS SCROFA UTERUS PREPARATION|PORCINE UTERUS PREPARATION
C0937628|T121|283568|RXNORM|GUGGUL LIPIDS|GUGGUL LIPIDS
C0770684|T197|235569|RXNORM|SULFURATED LIME|SULFURATED LIME
C2049071|T121|817635|RXNORM|INDOMETHACIN / THIAMINE|INDOMETHACIN / THIAMINE
C0055942|T121|21290|RXNORM|CLOROPHENE|CLOROPHENE
C1384247|T121|452651|RXNORM|OXYQUINOLINE / POTASSIUM SULFATE|OXYQUINOLINE / POTASSIUM SULFATE
C0023142|T109|1362875|RXNORM|DODECANOL|DODECANOL
C2929282|T121|1008377|RXNORM|CALCIUM CHLORIDE / LACTATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CHLORIDE / LACTATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C2929282|T121|1008377|RXNORM|CALCIUM CHLORIDE / LACTATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CHLORIDE / LACTATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C3644423|T121|1424888|RXNORM|FLUTICASONE / VILANTEROL|FLUTICASONE / VILANTEROL
C2935023|T121|1424884|RXNORM|VILANTEROL|VILANTEROL
C0244560|T109|1424880|RXNORM|ISOSTEARATE|ISOSTEARATE
C3256195|T121|1424881|RXNORM|JUGLANS REGIA SHELL EXTRACT|ENGLISH WALNUT SHELL EXTRACT
C3255936|T121|1310582|RXNORM|HYDROGENATED PALM GLYCERIDES|HYDROGENATED PALM GLYCERIDES
C3256169|T109|1310581|RXNORM|MENTHYL LACTATE|MENTHYL LACTATE
C0066258|T121|1310580|RXNORM|METHYL LACTATE|METHYL LACTATE
C0349375|T168|1310587|RXNORM|SKIM MILK|SKIM MILK
C1741925|T109|1310586|RXNORM|OCTYLTRIETHOXYSILANE|OCTYLTRIETHOXYSILANE
C2949375|T121|1310585|RXNORM|PHENYL TRIMETHICONE|PHENYL TRIMETHICONE
C3255780|T121|1310584|RXNORM|LAMINARIA DIGITATA PREPARATION|LAMINARIA DIGITATA PREPARATION
C0004589|T007|1595882|RXNORM|ANTHRAX BACTERIUM|BACILLUS ANTHRACIS
C2927368|T129|1005911|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-PERTH-16-2009 (H3N2) STRAIN|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-PERTH-16-2009 (H3N2) STRAIN
C0887117|T123|314709|RXNORM|ORNITHINE, (L)-ISOMER|ORNITHINE, (L)-ISOMER
C0027444|T195|7268|RXNORM|NATAMYCIN|NATAMYCIN
C0982252|T121|314705|RXNORM|LANOLIN / PETROLATUM|LANOLIN / PETROLATUM
C2168802|T121|812814|RXNORM|DIPIVEFRIN / LEVOBUNOLOL|DIPIVEFRIN / LEVOBUNOLOL
C3538279|T121|1372479|RXNORM|OLEOYL TYROSINE|OLEOYL TYROSINE
C0022938|T007|6204|RXNORM|LACTOBACILLUS|LACTOBACILLUS
C0022939|T007|6205|RXNORM|LACTOBACILLUS ACIDOPHILUS|LACTOBACILLUS ACIDOPHILUS
C2929898|T121|1009003|RXNORM|BENZYL BENZOATE / MONOSULFIRAM|BENZYL BENZOATE / MONOSULFIRAM
C2929897|T121|1009002|RXNORM|CHLORAMPHENICOL / OXYPHENBUTAZONE|CHLORAMPHENICOL / OXYPHENBUTAZONE
C2929900|T121|1009005|RXNORM|ACETYLCARNITINE / TYROSINE|ACETYLCARNITINE / TYROSINE
C2927862|T121|1006939|RXNORM|HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE / NEISSERIA MENINGITIDIS|HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE / NEISSERIA MENINGITIDIS
C2929902|T121|1009007|RXNORM|GLUTAMATE / VITAMIN B6|GLUTAMATE / VITAMIN B6
C2929901|T121|1009006|RXNORM|MAGNESIUM HYDROXIDE / SIMETHICONE|MAGNESIUM HYDROXIDE / SIMETHICONE
C2927857|T121|1006934|RXNORM|HAWTHORN BERRY / HAWTHORN BERRY EXTRACT|HAWTHORN BERRY / HAWTHORN BERRY EXTRACT
C2929903|T121|1009008|RXNORM|COBALT GLUCONATE / MANGANESE GLUCONATE|COBALT GLUCONATE / MANGANESE GLUCONATE
C2927860|T121|1006937|RXNORM|GRIFFONIA PREPARATION / KAVA ROOT / MELATONIN|GRIFFONIA PREPARATION / KAVA ROOT / MELATONIN
C2927853|T121|1006930|RXNORM|COENZYME Q10 / LEVOCARNITINE|COENZYME Q10 / LEVOCARNITINE
C2927854|T121|1006931|RXNORM|BORON / CALCIUM CARBONATE|BORON / CALCIUM CARBONATE
C2927855|T121|1006932|RXNORM|MENTHOL / SALICYLIC ACID|MENTHOL / SALICYLIC ACID
C2927856|T121|1006933|RXNORM|BENZYDAMINE / CETYLPYRIDINIUM|BENZYDAMINE / CETYLPYRIDINIUM
C0770985|T121|1311363|RXNORM|POTASSIUM SODIUM TARTRATE|POTASSIUM SODIUM TARTRATE
C3848578|T121|1546208|RXNORM|BARIUM CITRATE|BARIUM CITRATE
C1659521|T121|605999|RXNORM|CHLORPHENIRAMINE / METHSCOPOLAMINE|CHLORPHENIRAMINE / METHSCOPOLAMINE
C1659521|T121|605999|RXNORM|CHLORPHENIRAMINE / METHSCOPOLAMINE|CHLORPHENIRAMINE / METHSCOPOLAMINE
C1659520|T121|605998|RXNORM|CHLORPHENIRAMINE / CODEINE|CHLORPHENIRAMINE / CODEINE
C0025598|T121|6809|RXNORM|METFORMIN|METFORMIN
C2364496|T129|805467|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED, A-H1N1 (A-BRISBANE-59-2007) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED, A-H1N1 (A-BRISBANE-59-2007) STRAIN
C0025575|T121|6805|RXNORM|METARAMINOL|METARAMINOL
C0019573|T123|1546205|RXNORM|HIRUDIN|HIRUDIN
C3848579|T121|1546206|RXNORM|CROTON TIGLIUM WHOLE EXTRACT|CROTON TIGLIUM WHOLE EXTRACT
C0040112|T123|10562|RXNORM|THYMUS EXTRACTS|THYMUS EXTRACTS
C0040108|T121|10561|RXNORM|MOXISYLYTE|MOXISYLYTE
C3256182|T121|1307944|RXNORM|SEDUM ROSEUM ROOT EXTRACT|RHODIOLA ROSEA ROOT EXTRACT
C0065767|T121|29365|RXNORM|CALCIPOTRIENE|CALCIPOTRIOL
C0040123|T125|10565|RXNORM|THYROGLOBULIN|THYROGLOBULIN
C3255613|T109|1366228|RXNORM|TRIACONTANYL PVP (WP-660)|TRIACONTANYL PVP (WP-660)
C0282351|T122|1366227|RXNORM|DIMETHICONE 20|DIMETHICONE 20
C3531179|T109|1366226|RXNORM|OXACYCLOHEPTADEC-8-EN-2-ONE, (8Z)-|OXACYCLOHEPTADEC-8-EN-2-ONE, (8Z)-
C3531177|T121|1366223|RXNORM|CARBOMER INTERPOLYMER TYPE B (ALLYL PENTAERYTHRITOL CROSSLINKED)|CARBOMER INTERPOLYMER TYPE B (ALLYL PENTAERYTHRITOL CROSSLINKED)
C3255708|T121|1307942|RXNORM|NYMPHAEA CAERULEA FLOWER EXTRACT|NYMPHAEA CAERULEA FLOWER EXTRACT
C2608637|T121|833079|RXNORM|SMALLPOX VACCINE LIVE VACCINIA VIRUS|SMALLPOX VACCINE LIVE VACCINIA VIRUS
C3538277|T121|1372477|RXNORM|VOACANGA AFRICANA SEED EXTRACT|VOACANGA AFRICANA SEED EXTRACT
C0526354|T121|1362933|RXNORM|2,2,4,4,6,8,8-HEPTAMETHYLNONANE|ISOHEXADECANE
C0259568|T109|1362932|RXNORM|LAURIC ACID METHYL ESTER|METHYL LAURATE
C0073589|T130|1362931|RXNORM|ROSIN|ROSIN
C3256079|T121|1307098|RXNORM|PEG-7 GLYCERYL COCOATE|PEG-7 GLYCERYL COCOATE
C0075503|T121|37319|RXNORM|SULCONAZOLE|SULCONAZOLE
C2036577|T121|823128|RXNORM|ACETAMINOPHEN / STYRAMATE|ACETAMINOPHEN / STYRAMATE
C0028369|T125|7519|RXNORM|NORGESTRIENONE|NORGESTRIENONE
C0053152|T121|18923|RXNORM|BENZARONE|BENZARONE
C0033621|T123|8834|RXNORM|PROTEIN C|PROTEIN C
C0075501|T127|37317|RXNORM|SULBUTIAMINE|SULBUTIAMINE
C1509684|T121|1367129|RXNORM|POLYVINYL ACETATE PHTHALATE|POLYVINYL ACETATE PHTHALATE
C0022516|T121|6111|RXNORM|KARAYA GUM|STERCULIA
C0066923|T121|30320|RXNORM|MUCOPOLYSACCHARIDE POLYSULFATE|MUCOPOLYSACCHARIDE POLYSULFATE
C0065023|T195|1111103|RXNORM|FIDAXOMICIN|FIDAXOMICIN
C3857945|T121|1552451|RXNORM|DIDECYL ETHER|DIDECYL ETHER
C0010621|T121|3014|RXNORM|CYPROTERONE|CYPROTERONE
C0029112|T121|7676|RXNORM|OPIUM|OPIUM
C0029112|T121|7676|RXNORM|OPIUM|OPIUM
C0029105|T121|7674|RXNORM|OPIPRAMOL|OPIPRAMOL
C1171274|T121|353497|RXNORM|LEVOBETAXOLOL|LEVOBETAXOLOL
C0059693|T131|1314352|RXNORM|ETHANETHIOL|ETHANETHIOL
C0062640|T130|1311540|RXNORM|HEXAMETHYLDISILOXANE|HEXAMETHYLDISILOXANE
C0014713|T123|1314350|RXNORM|ERGOTHIONEINE|ERGOTHIONEINE
C0014839|T130|1314351|RXNORM|ESCULIN|ESCULIN
C0059755|T109|1314356|RXNORM|ETHYL BUTYRATE|ETHYL BUTYRATE
C1259844|T109|1314357|RXNORM|ETHYL ISOVALERATE|ETHYL ISOVALERATE
C2827224|T121|1311186|RXNORM|LAURAMIDOPROPYL BETAINE|LAURAMIDOPROPYL BETAINE
C3500342|T121|1314245|RXNORM|LAPSANA COMMUNIS WHOLE EXTRACT|LAPSANA COMMUNIS WHOLE EXTRACT
C2917636|T121|1311188|RXNORM|PULSATILLA VULGARIS EXTRACT|ANEMONE PULSATILLA EXTRACT
C3255756|T121|1314358|RXNORM|ETHYL MACADAMIATE|ETHYL MACADAMIATE
C0059773|T121|1314359|RXNORM|ETHYL MALTOL|ETHYL MALTOL
C0053407|T122|1362685|RXNORM|BETADEX|BETADEX
C0057717|T196|1362686|RXNORM|DIAMOND|DIAMOND
C3256065|T109|1305728|RXNORM|PEG-150 DISETEARATE|PEG-150 DISETEARATE
C3500344|T121|1314247|RXNORM|PHYTOLACCA AMERICANA FRUIT EXTRACT|PHYTOLACCA AMERICANA FRUIT EXTRACT
C0055370|T197|20799|RXNORM|CHLORINE DIOXIDE|CHLORINE DIOXIDE
C3255748|T109|1305720|RXNORM|CHINESE CINNAMON EXTRACT|CHINESE CINNAMON EXTRACT
C3257526|T109|1305725|RXNORM|LIME (CITRUS) EXTRACT|LIME (CITRUS) EXTRACT
C0006217|T126|1752|RXNORM|BROMELAINS|BROMELAINS
C2827175|T121|1305727|RXNORM|HYDROXYETHYL CELLULOSE (140 CPS AT 5%)|HYDROXYETHYL CELLULOSE (140 MPA.S AT 5 % )
C3500340|T121|1314241|RXNORM|GLYCERETH-17 STEARATE|GLYCERETH-17 STEARATE
C0669247|T122|1000577|RXNORM|MICROCRYSTALLINE CELLULOSE|MICROCRYSTALLINE CELLULOSE
C3486747|T121|1311246|RXNORM|RAPHANUS SATIVA EXTRACT|RAPHANUS SATIVA EXTRACT
C0379149|T121|115243|RXNORM|TEMOPORFIN|TEMOPORFIN
C2345471|T121|1314243|RXNORM|PPG 12 BUTETH 16|PPG 12 BUTETH 16
C3488058|T121|1309934|RXNORM|FRANGULA CALIFORNICA BARK EXTRACT|FRANGULA CALIFORNICA BARK EXTRACT
C3486631|T121|1309936|RXNORM|CASTANEA SATIVA FLOWER EXTRACT|CASTANEA SATIVA FLOWER EXTRACT
C3488087|T121|1309937|RXNORM|LATHYRUS SATIVAS SEED EXTRACT|LATHYRUS SATIVAS SEED EXTRACT
C0059772|T121|24524|RXNORM|ETHYL LOFLAZEPATE|ETHYL LOFLAZEPATE
C2740754|T129|899650|RXNORM|PIGNUT HICKORY POLLEN EXTRACT|CARYA GLABRA POLLEN EXTRACT
C0059770|T121|24522|RXNORM|ETHYL LINOLEATE|ETHYL LINOLEATE
C0117899|T121|50097|RXNORM|FLUINDIONE|FLUINDIONE
C3528919|T121|1363729|RXNORM|EUCALYPTUS GLOBULUS WHOLE EXTRACT|EUCALYPTUS GLOBULUS WHOLE EXTRACT
C2929423|T121|1008519|RXNORM|GUAIACOLSULFONATE / HYDROCODONE|GUAIACOLSULFONATE / HYDROCODONE
C0771653|T121|1310350|RXNORM|DATURA STRAMONIUM EXTRACT|DATURA STRAMONIUM EXTRACT
C2929414|T121|1008510|RXNORM|MAGNESIUM LACTATE / VITAMIN B6|MAGNESIUM LACTATE / VITAMIN B6
C2929415|T121|1008511|RXNORM|CAMPHOR / MENTHOL / NIACIN|CAMPHOR / MENTHOL / NIACIN
C2929416|T121|1008512|RXNORM|DIMETHICONE / PETROLATUM|DIMETHICONE / PETROLATUM
C2929416|T121|1008512|RXNORM|DIMETHICONE / PETROLATUM|DIMETHICONE / PETROLATUM
C2929417|T121|1008513|RXNORM|DIISOPROMINE / SORBITOL|DIISOPROMINE / SORBITOL
C2929419|T121|1008515|RXNORM|CALCIUM CARBONATE / FOLIC ACID / PYRIDOXINE / VITAMIN B 12|CALCIUM CARBONATE / FOLIC ACID / PYRIDOXINE / VITAMIN B 12
C2929420|T121|1008516|RXNORM|IODINE POVACRYLEX / ISOPROPYL ALCOHOL|IODINE POVACRYLEX / ISOPROPYL ALCOHOL
C2929421|T121|1008517|RXNORM|PHENOL / ZINC OXIDE|PHENOL / ZINC OXIDE
C3247695|T121|1192792|RXNORM|EUROPEAN HOUSE DUST MITE EXTRACT / WHITE OAK POLLEN EXTRACT|EUROPEAN HOUSE DUST MITE EXTRACT / WHITE OAK POLLEN EXTRACT
C3464653|T121|1312987|RXNORM|DIMETHYL PALMITAMINE|DIMETHYL PALMITAMINE
C0033459|T121|8766|RXNORM|PERICIAZINE|PERICIAZINE
C0033447|T121|8761|RXNORM|PROPANTHELINE|PROPANTHELINE
C1875751|T121|690353|RXNORM|SILICONES / STARCH|SILICONES / STARCH
C1720236|T121|645555|RXNORM|BACITRACIN / POLYMYXIN B|BACITRACIN / POLYMYXIN B
C1720236|T121|645555|RXNORM|BACITRACIN / POLYMYXIN B|BACITRACIN / POLYMYXIN B
C0002563|T123|683|RXNORM|AMINOLEVULINIC ACID|AMINOLEVULINIC ACID
C2049070|T121|814504|RXNORM|DEXAMETHASONE / INDOMETHACIN|DEXAMETHASONE / INDOMETHACIN
C0771350|T121|1363721|RXNORM|NIACINAMIDE ASCORBATE|NIACINAMIDE ASCORBATE
C0526737|T109|1363720|RXNORM|MYRISTYL LACTATE|MYRISTYL LACTATE
C2728192|T129|1011633|RXNORM|WHITE PEPPER ALLERGENIC EXTRACT|WHITE PEPPER ALLERGENIC EXTRACT
C0293273|T123|85982|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 6|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 6
C2938758|T121|1012890|RXNORM|ASARUM EUROPAEUM EXTRACT|ASARUM EUROPAEUM EXTRACT
C2726205|T129|883459|RXNORM|PUMPKIN ALLERGENIC EXTRACT|CUCURBITA PEPO ALLERGENIC EXTRACT
C0064304|T121|28181|RXNORM|KETAZOLAM|KETAZOLAM
C0220838|T123|1426907|RXNORM|GLUCURONATE|GLUCURONATE
C0009968|T196|2837|RXNORM|HCG ALPHA,RECOMBINANT|COPPER
C3864848|T121|1595582|RXNORM|CORDYCEPS GUNNII FRUITING BODY EXTRACT|CORDYCEPS GUNNII FRUITING BODY EXTRACT
C0910661|T121|1426903|RXNORM|DROMETRIZOLE|DROMETRIZOLE
C3542458|T121|1428218|RXNORM|ERECHTITES HIERACIIFOLIUS EXTRACT|ERECHTITES HIERACIIFOLIUS EXTRACT
C3282506|T121|1426901|RXNORM|DECYLENE GLYCOL|DECYLENE GLYCOL
C3281578|T122|1426900|RXNORM|SILK, BASE HYDROLYZED (1000 MW)|SILK, BASE HYDROLYZED (1000 MW)
C3651788|T121|1428215|RXNORM|POLYQUATERNIUM-10 (30000 MPA.S AT 2%)|POLYQUATERNIUM-10 (30000 MPA.S AT 2%)
C3651789|T121|1428214|RXNORM|ALISMA PLANTAGO-AQUATICA TOP EXTRACT|ALISMA PLANTAGO-AQUATICA TOP EXTRACT
C0056595|T121|1428217|RXNORM|CUPRIC GLYCINATE|CUPRIC GLYCINATE
C3542446|T121|1428216|RXNORM|CHENOPODIUM VULVARIA EXTRACT|CHENOPODIUM VULVARIA EXTRACT
C3256743|T109|1426909|RXNORM|DIISOPROPYL DILINOLEATE|DIISOPROPYL DILINOLEATE
C3256826|T109|1426908|RXNORM|CAPSOSIPHON FULVESCENS EXTRACT|CAPSOSIPHON FULVESCENS EXTRACT
C0936126|T121|282436|RXNORM|FENUGREEK SEED MEAL|FENUGREEK SEED MEAL
C0051928|T121|1313764|RXNORM|ANNATTO EXTRACT|ANNATTO EXTRACT
C0072857|T121|35208|RXNORM|QUINAPRIL|QUINAPRIL
C3500063|T197|1313762|RXNORM|YTTRIUM FLUORIDE|YTTRIUM FLUORIDE
C3500064|T197|1313763|RXNORM|YTTRIUM IODIDE|YTTRIUM IODIDE
C3500062|T197|1313761|RXNORM|YTTRIUM BROMIDE|YTTRIUM BROMIDE
C0065295|T195|28981|RXNORM|LORACARBEF|LORACARBEF
C2928329|T121|1007407|RXNORM|ASCORBIC ACID / ASPIRIN / CYSTEINE|ASCORBIC ACID / ASPIRIN / CYSTEINE
C2928328|T121|1007406|RXNORM|ISOMYRTOL / PHOLCODINE|ISOMYRTOL / PHOLCODINE
C2928327|T121|1007405|RXNORM|INSULIN, PROMPT ZINC, HUMAN / INSULIN, ZINC, HUMAN|INSULIN, PROMPT ZINC, HUMAN / INSULIN, ZINC, HUMAN
C2928326|T121|1007404|RXNORM|CALCIUM CARBONATE / SOY PROTEIN ISOLATE / VITAMIN D|CALCIUM CARBONATE / SOY PROTEIN ISOLATE / VITAMIN D
C2928325|T121|1007403|RXNORM|CALCIUM CHLORIDE / GLUCOSE / POTASSIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CHLORIDE / GLUCOSE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C3256662|T121|1307645|RXNORM|ASPALATHUS LINEARIS LEAF EXTRACT|ASPALATHUS LINEARIS LEAF EXTRACT
C3474200|T121|1307646|RXNORM|POGOSTEMON CABLIN TOP EXTRACT|POGOSTEMON CABLIN TOP EXTRACT
C2928322|T121|1007400|RXNORM|DIHYDROERGOCORNINE / DIHYDROERGOCRISTINE / DIHYDROERGOCRYPTINE|DIHYDROERGOCORNINE / DIHYDROERGOCRISTINE / DIHYDROERGOCRYPTINE
C3256410|T121|1307648|RXNORM|ANNICKIA CHLORANTHA BARK EXTRACT|ANNICKIA CHLORANTHA BARK EXTRACT
C3256505|T121|1307649|RXNORM|ARTEMISIA ARGYI LEAF EXTRACT|ARTEMISIA ARGYI LEAF EXTRACT
C0123091|T121|51272|RXNORM|QUETIAPINE|QUETIAPINE
C2928331|T121|1007409|RXNORM|LACTATE / PYRROLIDONECARBOXYLIC ACID / UREA|LACTATE / PYRROLIDONECARBOXYLIC ACID / UREA
C2928330|T121|1007408|RXNORM|FERROUS FUMARATE / VITAMIN B 12|FERROUS FUMARATE / VITAMIN B 12
C1874648|T121|691006|RXNORM|CALCIUM CARBONATE / FERROUS FUMARATE / VITAMIN D|CALCIUM CARBONATE / FERROUS FUMARATE / VITAMIN D
C1874647|T121|691005|RXNORM|CALCIUM CARBONATE / FAMOTIDINE / MAGNESIUM HYDROXIDE|CALCIUM CARBONATE / FAMOTIDINE / MAGNESIUM HYDROXIDE
C1655137|T121|606640|RXNORM|CHLORDIAZEPOXIDE / METHSCOPOLAMINE|CHLORDIAZEPOXIDE / METHSCOPOLAMINE
C1656695|T121|606642|RXNORM|FENTANYL / ROPIVACAINE|FENTANYL / ROPIVACAINE
C2014106|T121|819758|RXNORM|NIMESULIDE / ORPHENADRINE|NIMESULIDE / ORPHENADRINE
C0041111|T109|1368872|RXNORM|TRISTEARIN|GLYCERYL TRISTEARATE
C1874650|T121|691008|RXNORM|CALCIUM CARBONATE / GLYCINE|CALCIUM CARBONATE / GLYCINE
C3651726|T109|1430130|RXNORM|PEG-20 METHYL GLUCOSE SESQUISTEARATE|PEG-20 METHYL GLUCOSE SESQUISTEARATE
C1720624|T121|644513|RXNORM|SODIUM BICARBONATE / SODIUM CHLORIDE|SODIUM BICARBONATE / SODIUM CHLORIDE
C3667810|T121|1440064|RXNORM|CAMPHOR / CAPSAICIN / METHYL SALICYLATE|CAMPHOR / CAPSAICIN / METHYL SALICYLATE
C1874069|T121|687195|RXNORM|ALLANTOIN / COAL TAR|ALLANTOIN / COAL TAR
C1874170|T121|687198|RXNORM|ALUMINUM HYDROXIDE / MAGNESIUM TRISILICATE|ALUMINUM HYDROXIDE / MAGNESIUM TRISILICATE
C3832793|T121|1539637|RXNORM|TRIMETHYLOLPROPANE TRIISOSTEARATE|TRIMETHYLOLPROPANE TRIISOSTEARATE
C0025503|T121|6781|RXNORM|MESTEROLONE|MESTEROLONE
C0025506|T121|6782|RXNORM|MESTRANOL|MESTRANOL
C2729799|T129|891776|RXNORM|ARTICHOKE ALLERGENIC EXTRACT|ARTICHOKE ALLERGENIC EXTRACT
C0006034|T007|1426882|RXNORM|BORRELIA BURGDORFERI|BORRELIA BURGDORFERI
C1875202|T121|689425|RXNORM|GLYCERIN / KAOLIN / SODIUM FLUORIDE|GLYCERIN / KAOLIN / SODIUM FLUORIDE
C1875205|T121|689428|RXNORM|GLYCERIN / LYSINE|GLYCERIN / LYSINE
C3651795|T121|1427412|RXNORM|DIPENTAERYTHRITYL HEXA C5-10 ACID ESTERS|DIPENTAERYTHRITYL HEXA C5-10 ACID ESTERS
C3541351|T121|1427413|RXNORM|LINGONBERRY EXTRACT|LINGONBERRY EXTRACT
C2168926|T121|817286|RXNORM|AMINOPHYLLINE / QUININE|AMINOPHYLLINE / QUININE
C0385178|T121|117896|RXNORM|BENZQUERCIN|BENZQUERCIN
C0069008|T121|32009|RXNORM|NORMETHADONE|NORMETHADONE
C0596019|T196|153974|RXNORM|CHLORIDE ION|CL -
C0001187|T130|249|RXNORM|ACRIFLAVINE|EUFLAVINE
C0044295|T109|1427076|RXNORM|GLYCERYL ARACHIDONATE|GLYCERYL ARACHIDONATE
C3191304|T121|1306119|RXNORM|BLACKFOOT ABALONE EXTRACT|BLACKFOOT ABALONE EXTRACT
C3154338|T121|1306118|RXNORM|NEW ZEALAND GREEN MUSSEL EXTRACT|NEW ZEALAND GREEN MUSSEL EXTRACT
C2955065|T125|1306117|RXNORM|GONADOTROPIN RELEASING HORMONE, D-ARG(6) ETHYL AMIDE ACETATE|GONADOTROPIN RELEASING HORMONE, D-ARG(6) ETHYL AMIDE ACETATE
C2698346|T121|1306115|RXNORM|BEMOTRIZINOL|BEMOTRIZINOL
C3282449|T121|1306112|RXNORM|2,2'-DITHIOBISBENZOTHIAZOLE|2,2'-DITHIOBISBENZOTHIAZOLE
C0038711|T195|1306111|RXNORM|SULFAQUINOXALINE|SULFAQUINOXALINE
C0220853|T196|1314279|RXNORM|HYDROXIDE ION|HYDROXIDE ION
C0035100|T126|9248|RXNORM|CHYMOSIN|CHYMOSIN
C3643354|T109|1422485|RXNORM|MELALEUCA ERICIFOLIA LEAF OIL|MELALEUCA ERICIFOLIA LEAF OIL
C1445748|T121|466514|RXNORM|CHLORPHENIRAMINE / HYDROCODONE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / HYDROCODONE / PSEUDOEPHEDRINE
C3535845|T121|1370648|RXNORM|LAUROAMPHODIACETATE|LAUROAMPHODIACETATE
C1445751|T121|466517|RXNORM|ACETAMINOPHEN / DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE
C0060229|T197|24898|RXNORM|FERRIC CHLORIDE|FERRIC CHLORIDE
C1445746|T121|466512|RXNORM|CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE / POTASSIUM IODIDE|CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE / POTASSIUM IODIDE
C1445747|T121|466513|RXNORM|CARBETAPENTANE / CHLORPHENIRAMINE / EPHEDRINE / PHENYLEPHRINE|CARBETAPENTANE / CHLORPHENIRAMINE / EPHEDRINE / PHENYLEPHRINE
C2700159|T130|1370642|RXNORM|VERSETAMIDE|VERSETAMIDE
C3535848|T121|1370643|RXNORM|2,2'-DIHYDROXY-4,4'-DIMETHOXY-5,5'-DISULFOBENZOPHENONE|2,2'-DIHYDROXY-4,4'-DIMETHOXY-5,5'-DISULFOBENZOPHENONE
C3535850|T197|1370640|RXNORM|STANNATE|STANNATE
C0060228|T121|24897|RXNORM|FERRIC AMMONIUM CITRATE|FERRIC AMMONIUM CITRATE
C3535846|T121|1370646|RXNORM|LAURETH SULFOSUCCINATE|LAURETH SULFOSUCCINATE
C3535847|T121|1370644|RXNORM|C12-14 SEC-PARETH-12 SULFOSUCCINATE|C12-14 SEC-PARETH-12 SULFOSUCCINATE
C0540776|T195|141440|RXNORM|ALATROFLOXACIN|ALATROFLOXACIN
C3710015|T121|1488819|RXNORM|LACHESIS MUTA WHOLE EXTRACT|LACHESIS MUTA WHOLE EXTRACT
C0055729|T121|21107|RXNORM|CILOSTAZOL|CILOSTAZOL
C2080532|T121|818576|RXNORM|METHAPYRILENE / PHENYLEPHRINE|METHAPYRILENE / PHENYLEPHRINE
C2741492|T129|901307|RXNORM|SWEET POTATO ALLERGENIC EXTRACT|SWEET POTATO ALLERGENIC EXTRACT
C3282117|T121|1426949|RXNORM|PEG-PPG-105-5 COPOLYMER|PEG-PPG-105-5 COPOLYMER
C2741489|T129|901303|RXNORM|SWEET CHERRY ALLERGENIC EXTRACT|PRUNUS AVIUM ALLERGENIC EXTRACT
C3474802|T121|1301858|RXNORM|TURPENTINE / WHITE SPIRIT TYPE 1|TURPENTINE / WHITE SPIRIT TYPE 1
C3267752|T122|1301854|RXNORM|WHITE SPIRIT TYPE 1|WHITE SPIRIT TYPE 1
C3651702|T121|1431709|RXNORM|RUBUS IDAEUS SEED EXTRACT|RUBUS IDAEUS SEED EXTRACT
C0052971|T197|1305530|RXNORM|BARIUM CARBONATE|BARIUM CARBONATE
C2146619|T121|820749|RXNORM|ACETAMINOPHEN / DIPYRONE|ACETAMINOPHEN / DIPYRONE
C3256004|T121|1363588|RXNORM|HYPROMELLOSE 2208|HYPROMELLOSE 2208
C3651703|T121|1431705|RXNORM|MAURITIA FLEXUOSA WHOLE EXTRACT|MAURITIA FLEXUOSA WHOLE EXTRACT
C0592532|T121|152610|RXNORM|CERTOPARIN|CERTOPARIN
C0012586|T121|3523|RXNORM|DIPYRONE|DIPYRONE
C0012582|T121|3521|RXNORM|DIPYRIDAMOLE|DIPYRIDAMOLE
C0012582|T121|3521|RXNORM|DIPYRIDAMOLE|DIPYRIDAMOLE
C0025446|T131|6774|RXNORM|MERSALYL|MERSALYL
C1875028|T121|690691|RXNORM|DIPHENHYDRAMINE / HYDROCORTISONE|DIPHENHYDRAMINE / HYDROCORTISONE
C3255777|T121|1311635|RXNORM|LYCIUM CHINENSE FRUIT EXTRACT|LYCIUM CHINENSE FRUIT EXTRACT
C3475290|T109|1305536|RXNORM|APRICOT KERNAL OIL PEG-6 ESTERS|APRICOT KERNAL OIL PEG-6 ESTERS
C0071832|T121|1423683|RXNORM|GLYCERYL PALMITOSTEARATE|GLYCERYL PALMITOSTEARATE
C3194726|T129|1117083|RXNORM|WEAKLEAF BUR RAGWEED POLLEN EXTRACT|AMBROSIA CONFERTIFLORA POLLEN EXTRACT
C0771787|T121|1423684|RXNORM|HYPOPHOSPHORUS ACID|HYPOPHOSPHORUS ACID
C2731673|T109|895808|RXNORM|PHENYL SALICYATE|PHENYL SALICYATE
C2344271|T129|798226|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 23F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 23F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C3256100|T121|1363583|RXNORM|HYPROMELLOSE 2910-5CP|HYPROMELLOSE 2910-5CP
C0137984|T121|54987|RXNORM|POTASSIUM ACETATE|POTASSIUM ACETATE
C2929648|T121|1008749|RXNORM|CALCIUM CARBONATE / MAGNESIUM OXIDE / ZINC SULFATE|CALCIUM CARBONATE / MAGNESIUM OXIDE / ZINC SULFATE
C0717520|T121|214326|RXNORM|BROMPHENIRAMINE / PSEUDOEPHEDRINE|BROMPHENIRAMINE / PSEUDOEPHEDRINE
C2929644|T121|1008745|RXNORM|DEXTROMETHORPHAN / EPHEDRINE|DEXTROMETHORPHAN / EPHEDRINE
C2929643|T121|1008744|RXNORM|MINERAL OIL / PROPYLENE GLYCOL / TRIETHANOLAMINE|MINERAL OIL / PROPYLENE GLYCOL / TRIETHANOLAMINE
C2929646|T121|1008747|RXNORM|FORMALDEHYDE / ISOPROPYL ALCOHOL|FORMALDEHYDE / ISOPROPYL ALCOHOL
C2929645|T121|1008746|RXNORM|SALICYLIC ACID / UNDECYLENATE|SALICYLIC ACID / UNDECYLENATE
C2929640|T121|1008741|RXNORM|DIMETHICONE / MINERAL OIL / ZINC OXIDE|DIMETHICONE / MINERAL OIL / ZINC OXIDE
C2929639|T121|1008740|RXNORM|CHROMIC CHLORIDE / NIACIN|CHROMIC CHLORIDE / NIACIN
C0074726|T197|36679|RXNORM|SODIUM BISULFITE|SODIUM BISULFITE
C3834054|T109|1543185|RXNORM|SUCROSE OCTASTEARATE|SUCROSE OCTASTEARATE
C1875714|T121|690185|RXNORM|QUINETHAZONE / RESERPINE|QUINETHAZONE / RESERPINE
C1615657|T126|578033|RXNORM|GALSULFASE|GALSULFASE
C3528820|T121|1363434|RXNORM|ISOPROPYL LAURATE|ISOPROPYL LAURATE
C2928900|T121|1007988|RXNORM|ASCORBIC ACID / VITAMIN B6 / ZINC CITRATE|ASCORBIC ACID / VITAMIN B6 / ZINC CITRATE
C2928901|T121|1007989|RXNORM|FOLIC ACID / IRON POLYSACCHARIDE / VITAMIN B 12|FOLIC ACID / IRON POLYSACCHARIDE / VITAMIN B 12
C3486820|T109|1358860|RXNORM|SESAME EXTRACT|SESAME EXTRACT
C3528819|T121|1363430|RXNORM|ATROPA BELLADONNA WHOLE EXTRACT|ATROPA BELLADONNA WHOLE EXTRACT
C2928894|T121|1007982|RXNORM|CALCIUM HYDROXIDE / ZINC OXIDE|CALCIUM HYDROXIDE / ZINC OXIDE
C2928895|T121|1007983|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-10-2007 (H3N2)-LIKE VIRUS (A-URUGUAY-716-2007 NYMC X-175C) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007, IVR-148 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED, B-FLORIDA-4-2006-LIKE VIRUS (B-FLORIDA-4-2006) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-10-2007 (H3N2)-LIKE VIRUS (A-URUGUAY-716-2007 NYMC X-175C) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-59-2007, IVR-148 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, INACTIVATED, B-FLORIDA-4-2006-LIKE VIRUS (B-FLORIDA-4-2006) STRAIN
C2928892|T121|1007980|RXNORM|ALANINE / ARGININE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2928893|T121|1007981|RXNORM|CLOTRIMAZOLE / UREA|CLOTRIMAZOLE / UREA
C2928898|T121|1007986|RXNORM|BETA SITOSTEROL / CAMPESTEROL / STIGMASTEROL|BETA SITOSTEROL / CAMPESTEROL / STIGMASTEROL
C2928899|T121|1007987|RXNORM|BLACK CURRANT OIL / VITAMIN E|BLACK CURRANT OIL / VITAMIN E
C2928896|T121|1007984|RXNORM|ASCORBIC ACID / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / SODIUM FLUORIDE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D / VITAMIN E|ASCORBIC ACID / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / SODIUM FLUORIDE / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN D / VITAMIN E
C2073921|T121|816659|RXNORM|ACEMETACIN / CHLORZOXAZONE|ACEMETACIN / CHLORZOXAZONE
C3497576|T121|1310119|RXNORM|MYOSOTIS SYLVATICA FLOWERING TOP EXTRACT|MYOSOTIS SYLVATICA FLOWERING TOP EXTRACT
C0006213|T121|1749|RXNORM|BROMAZEPAM|BROMAZEPAM
C3497573|T109|1310114|RXNORM|BALANITES ROXBURGHII SEED OIL|BALANITES ROXBURGHII SEED OIL
C3497574|T121|1310115|RXNORM|ORNITHOGALUM UMBELLATUM FLOWERING TOP EXTRACT|ORNITHOGALUM UMBELLATUM FLOWERING TOP EXTRACT
C3497575|T121|1310117|RXNORM|CITRUS AURANTIIFOLIA FLOWER EXTRACT|CITRUS AURANTIIFOLIA FLOWER EXTRACT
C3486809|T121|1310110|RXNORM|SCLERANTHUS ANNUUS FLOWERING TOP EXTRACT|SCLERANTHUS ANNUUS FLOWERING TOP EXTRACT
C3489390|T121|1310111|RXNORM|AMANITA MUSCARIA VAR. MUSCARIA FRUITING BODY EXTRACT|AMANITA MUSCARIA VAR. MUSCARIA FRUITING BODY EXTRACT
C3474095|T121|1300188|RXNORM|BORDETELLA PERTUSSIS FILAMENTOUS HEMAGGLUTININ VACCINE, INACTIVATED / BORDETELLA PERTUSSIS FIMBRIAE 2/3 VACCINE, INACTIVATED / BORDETELLA PERTUSSIS PERTACTIN VACCINE, INACTIVATED / BORDETELLA PERTUSSIS TOXOID VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCI|BORDETELLA PERTUSSIS FILAMENTOUS HEMAGGLUTININ VACCINE, INACTIVATED / BORDETELLA PERTUSSIS FIMBRIAE 2/3 VACCINE, INACTIVATED / BORDETELLA PERTUSSIS PERTACTIN VACCINE, INACTIVATED / BORDETELLA PERTUSSIS TOXOID VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED
C3497572|T121|1310113|RXNORM|PAULOWNIA TOMENTOSA LEAF EXTRACT|PAULOWNIA TOMENTOSA LEAF EXTRACT
C0939809|T121|285160|RXNORM|POKEWEED PREPARATION|POKEWEED PREPARATION
C3484625|T121|1311538|RXNORM|ANGELICA KEISKEI TOP EXTRACT|ANGELICA KEISKEI TOP EXTRACT
C0939812|T121|285162|RXNORM|RUTA GRAVEOLENS PREPARATION|RUTA GRAVEOLENS PREPARATION
C0939814|T121|285164|RXNORM|SPIGELIA MARILANDICA PREPARATION|SPIGELIA MARILANDICA PREPARATION
C3818804|T121|1490679|RXNORM|ANGELICA DAHURICA WHOLE EXTRACT|ANGELICA DAHURICA WHOLE EXTRACT
C0939817|T121|285166|RXNORM|TOXICODENDRON PREPARATION|TOXICODENDRON PREPARATION
C0939818|T121|285167|RXNORM|URTICA URENS HOMEOPATHIC PREPARATION|URTICA URENS HOMEOPATHIC PREPARATION
C3256824|T121|1311531|RXNORM|EUROPEAN ELDERBERRY EXTRACT|EUROPEAN ELDERBERRY EXTRACT
C0065088|T197|1311533|RXNORM|LITHIUM CHLORIDE|LITHIUM CHLORIDE
C3527982|T121|1361491|RXNORM|BIDENS TRIPARTITA FLOWERING TOP EXTRACT|BIDENS TRIPARTITA FLOWERING TOP EXTRACT
C0025748|T131|1311537|RXNORM|METHYLENE CHLORIDE|METHYLENE CHLORIDE
C2928104|T121|1007182|RXNORM|VITAMIN A / VITAMIN E|VITAMIN A / VITAMIN E
C2928105|T121|1007183|RXNORM|GINKGO BILOBA EXTRACT / GINSENG PREPARATION / GOTU KOLA EXTRACT / LECITHIN|GINKGO BILOBA EXTRACT / GINSENG PREPARATION / GOTU KOLA EXTRACT / LECITHIN
C2928102|T121|1007180|RXNORM|LYSINE / POTASSIUM BICARBONATE / POTASSIUM CHLORIDE|LYSINE / POTASSIUM BICARBONATE / POTASSIUM CHLORIDE
C2928103|T121|1007181|RXNORM|HYOSCYAMUS EXTRACT / PHENAZOPYRIDINE / SULFAMETHIZOLE|HYOSCYAMUS EXTRACT / PHENAZOPYRIDINE / SULFAMETHIZOLE
C2928108|T121|1007186|RXNORM|ACETAMINOPHEN / BROMELAINS|ACETAMINOPHEN / BROMELAINS
C2928109|T121|1007187|RXNORM|MAGNESIUM OXIDE / VITAMIN E|MAGNESIUM OXIDE / VITAMIN E
C2928106|T121|1007184|RXNORM|INSULIN, ASPART PROTAMINE, HUMAN / INSULIN, ASPART, HUMAN|INSULIN, ASPART PROTAMINE, HUMAN / INSULIN, ASPART, HUMAN
C2928107|T121|1007185|RXNORM|CARBON DIOXIDE / NITROUS OXIDE|CARBON DIOXIDE / NITROUS OXIDE
C2830183|T121|996051|RXNORM|CABAZITAXEL|CABAZITAXEL
C2928110|T121|1007188|RXNORM|ACTIVATED CHARCOAL / METHENAMINE|ACTIVATED CHARCOAL / METHENAMINE
C2928111|T121|1007189|RXNORM|BENZOCAINE / CETYLPYRIDINIUM / ZINC CHLORIDE|BENZOCAINE / CETYLPYRIDINIUM / ZINC CHLORIDE
C0056060|T168|1309239|RXNORM|COCONUT OIL|COCONUT OIL
C0061240|T121|1309238|RXNORM|GERMANIUM DIOXIDE|GERMANIUM DIOXIDE
C0873034|T109|1309237|RXNORM|HYSSOPUS OFFICINALIS EXTRACT|HYSSOPUS OFFICINALIS FLOWERING TOP EXTRACT
C0304146|T168|1309236|RXNORM|PARSELY SEED OIL|PARSELY SEED OIL
C0767026|T109|1309235|RXNORM|1,10-DECANEDIOL|1,10-DECANEDIOL
C1647196|T109|1309233|RXNORM|CLOVE LEAF OIL|CLOVE LEAF OIL
C1366079|T109|1309232|RXNORM|CLARY SAGE OIL|CLARY SAGE OIL
C0141927|T197|1309231|RXNORM|SELENIUM DIOXIDE|SELENIUM DIOXIDE
C0254751|T168|1309230|RXNORM|ORANGE OIL|ORANGE OIL
C0058765|T121|23687|RXNORM|CALCIUM GLUCONATE M-HYDRATE|DROXICAM
C0982034|T007|314513|RXNORM|BCG, LIVE, MONTREAL STRAIN|BCG, LIVE, MONTREAL STRAIN
C0982038|T121|314517|RXNORM|BELLADONNA LEAF|BELLADONNA LEAF
C0771909|T121|236614|RXNORM|BUTCHER'S BROOM PREPARATION|BUTCHER'S BROOM PREPARATION
C2979094|T121|1090062|RXNORM|ASCORBIC ACID / BIOTIN / FOLIC ACID / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE|ASCORBIC ACID / BIOTIN / FOLIC ACID / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE
C0795594|T197|253160|RXNORM|CHROMIUM, CHELATED|CHROMIUM, CHELATED
C0058004|T121|23043|RXNORM|DIFLUPREDNATE|DIFLUPREDNATE
C2928290|T121|1007368|RXNORM|ANISOTROPINE / PHENOBARBITAL|ANISOTROPINE / PHENOBARBITAL
C2928291|T121|1007369|RXNORM|CARBOXYMETHYLCELLULOSE / POVIDONE|CARBOXYMETHYLCELLULOSE / POVIDONE
C2928288|T121|1007366|RXNORM|BARBITAL / VALERIAN ROOT EXTRACT|BARBITAL / VALERIAN ROOT EXTRACT
C2928289|T121|1007367|RXNORM|ALUMINUM HYDROXIDE / CARBENOXOLONE|ALUMINUM HYDROXIDE / CARBENOXOLONE
C2928286|T121|1007364|RXNORM|BROMPHENIRAMINE / GUAIFENESIN / PHENYLEPHRINE|BROMPHENIRAMINE / GUAIFENESIN / PHENYLEPHRINE
C2928287|T121|1007365|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-SOUTH DAKOTA-6-2007 (H1N1) (A-BRISBANE-59-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-URUGUAY -716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-BRISBANE-60-2008 STRAIN|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-SOUTH DAKOTA-6-2007 (H1N1) (A-BRISBANE-59-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-URUGUAY -716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-BRISBANE-60-2008 STRAIN
C2928284|T121|1007362|RXNORM|FLUMETHASONE / NEOMYCIN|FLUMETHASONE / NEOMYCIN
C2928285|T121|1007363|RXNORM|BENZOYL PEROXIDE / OXYQUINOLINE|BENZOYL PEROXIDE / OXYQUINOLINE
C2928282|T121|1007360|RXNORM|HYDROCHLOROTHIAZIDE / PINDOLOL|HYDROCHLOROTHIAZIDE / PINDOLOL
C0078299|T121|39580|RXNORM|VIQUIDIL|VIQUIDIL
C2929102|T121|1008195|RXNORM|ALGINIC ACID / MAGNESIUM CARBONATE|ALGINIC ACID / MAGNESIUM CARBONATE
C3555515|T121|1374852|RXNORM|ACETYL DIPEPTIDE-1 CETYL ESTER|ACETYL TYROSYLARGININE CETYL ESTER
C3556197|T121|1374850|RXNORM|BENZALKONIUM / CAMPHOR|BENZALKONIUM / CAMPHOR
C0058646|T121|1362744|RXNORM|DODICIN|DODICIN
C3486464|T121|1314314|RXNORM|PPG-3 BENZYL ETHER MYRISTATE|PPG-3 BENZYL ETHER MYRISTATE
C0061231|T121|1362746|RXNORM|GERANYLGERANYLACETONE|TEPRENONE
C2728193|T129|1011404|RXNORM|MANGO ALLERGENIC EXTRACT|MANGO ALLERGENIC EXTRACT
C0055086|T121|1362741|RXNORM|CERAMIDE 3|CERAMIDE NP
C3464686|T121|1292893|RXNORM|ALLANTOIN / BENZALKONIUM / BENZYL ALCOHOL|ALLANTOIN / BENZALKONIUM / BENZYL ALCOHOL
C0058435|T121|1362743|RXNORM|DIPYRITHIONE|DIPYRITHIONE
C2241670|T121|818852|RXNORM|CODEINE / PHENYLEPHRINE|CODEINE / PHENYLEPHRINE
C0220832|T130|1362748|RXNORM|FORMATE|FORMATE
C0077379|T121|38868|RXNORM|TROMANTADINE|TROMANTADINE
C3848587|T121|1545912|RXNORM|SEDUM ROSEUM WHOLE EXTRACT|SEDUM ROSEUM WHOLE EXTRACT
C2080594|T121|815616|RXNORM|PHENIRAMINE / PHENYLPROPANOLAMINE|PHENIRAMINE / PHENYLPROPANOLAMINE
C2364522|T129|805520|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-10-2007 (H3N2)-LIKE VIRUS (A-URUGUAY-716-2007 NYMC X-175C) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-BRISBANE-10-2007 (H3N2)-LIKE VIRUS (A-URUGUAY-716-2007 NYMC X-175C) STRAIN
C0030940|T126|8028|RXNORM|PEPTIDE HYDROLASES|PEPTIDE HYDROLASES
C3818695|T127|1536458|RXNORM|1.ALPHA.,24S-DIHYDROXYVITAMIN D2|1.ALPHA.,24S-DIHYDROXYVITAMIN D2
C0171462|T121|1012534|RXNORM|MELARSOMINE|MELARSOMINE
C0032535|T195|8536|RXNORM|POLYMYXIN B|POLYMYXIN B
C0771913|T121|236617|RXNORM|FERROUS ASPARTATE|FERROUS ASPARTATE
C1874833|T121|689638|RXNORM|CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLTOLOXAMINE|CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLTOLOXAMINE
C3255113|T121|1236141|RXNORM|CHONDROITIN SULFATES / GLUCOSAMINE / METHYLSULFONYLMETHANE / TOCOPHEROL|CHONDROITIN SULFATES / GLUCOSAMINE / METHYLSULFONYLMETHANE / TOCOPHEROL
C3256661|T121|1306933|RXNORM|ASCORBYL GLUCOSIDE|ASCORBYL GLUCOSIDE
C0028128|T197|7442|RXNORM|NITRIC OXIDE|NITRIC OXIDE
C3256205|T109|1306935|RXNORM|BRAZILLIAN PEPPER EXTRACT|BRAZILLIAN PEPPER EXTRACT
C0129533|T123|1313976|RXNORM|MYRISTATE|MYRISTATE
C0054302|T130|1306937|RXNORM|BUTYLPARABEN|BUTYLPARABEN
C2194251|T121|816693|RXNORM|HOMATROPINE / SIMETHICONE|HOMATROPINE / SIMETHICONE
C0059780|T121|1306938|RXNORM|ETHYL PALMITATE|ETHYL PALMITATE
C1874828|T121|689632|RXNORM|CHLORPHENIRAMINE / METHSCOPOLAMINE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / METHSCOPOLAMINE / PSEUDOEPHEDRINE
C1874829|T121|689633|RXNORM|CHLORPHENIRAMINE / PHENINDAMINE / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / PHENINDAMINE / PHENYLPROPANOLAMINE
C1874830|T121|689635|RXNORM|CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C1874832|T121|689637|RXNORM|CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PYRILAMINE|CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PYRILAMINE
C2928365|T121|1007443|RXNORM|FERROUS SUCCINATE / SUCCINIC ACID|FERROUS SUCCINATE / SUCCINIC ACID
C0001521|T121|333|RXNORM|ADIPHENINE|ADIPHENINE
C3499509|T121|1312372|RXNORM|THUJOPSIS DOLABRATA LEAFY TWIG EXTRACT|THUJOPSIS DOLABRATA LEAFY TWIG EXTRACT
C3499510|T121|1312373|RXNORM|TETRASODIUM GLUTAMATE DIACETATE|TETRASODIUM GLUTAMATE DIACETATE
C3499507|T121|1312370|RXNORM|HUMAN SPUTUM, BORDETELLA PERTUSSIS INFECTED|HUMAN SPUTUM, BORDETELLA PERTUSSIS INFECTED
C3499508|T121|1312371|RXNORM|THUJOPSIS DOLABRATA WHOLE EXTRACT|THUJOPSIS DOLABRATA WHOLE EXTRACT
C0029348|T005|1312376|RXNORM|INFLUENZA B VIRUS|INFLUENZA B VIRUS
C3499514|T121|1312377|RXNORM|MAGNOLIA KOBUS BARK EXTRACT|MAGNOLIA KOBUS BARK EXTRACT
C3643365|T109|1421445|RXNORM|CASEIN, STREPTOCOCCUS THERMOPHILUS CULTURED, PROPIONIBACTERIUM FREUDENREICHII SUBSP. SHERMANII CULTURED, AGED PREPARATION|CASEIN, STREPTOCOCCUS THERMOPHILUS CULTURED, PROPIONIBACTERIUM FREUDENREICHII SUBSP. SHERMANII CULTURED, AGED PREPARATION
C0029347|T005|1312375|RXNORM|INFLUENZA A VIRUS|INFLUENZA A VIRUS
C3499515|T121|1312378|RXNORM|RUBUS CHAMAEMORUS SEED EXTRACT|RUBUS CHAMAEMORUS SEED EXTRACT
C3499516|T121|1312379|RXNORM|HEXAPLEX TRUNCULUS HYPOBRANCHIAL GLAND JUICE|HEXAPLEX TRUNCULUS HYPOBRANCHIAL GLAND JUICE
C0872913|T126|259280|RXNORM|TENECTEPLASE|TENECTEPLASE
C0872916|T196|259282|RXNORM|XENON-133|XENON-133
C3505518|T121|1358698|RXNORM|BOS TAURUS BRAIN PREPARATION|BOVINE BRAIN PREPARATION
C0052276|T121|1425353|RXNORM|GALACTOARABINAN|GALACTOARABINAN
C0991770|T130|317177|RXNORM|ALBUMIN,IODINATED I-125 SERUM|ALBUMIN,IODINATED I-125 SERUM
C2073916|T121|822470|RXNORM|ACETAMINOPHEN / CHLORPHENOXAMINE / PHENYLEPHRINE|ACETAMINOPHEN / CHLORPHENOXAMINE / PHENYLEPHRINE
C0031507|T121|8183|RXNORM|PHENYTOIN|PHENYTOIN
C3644623|T109|1425354|RXNORM|HYDROGENATED TALLOW ACID|HYDROGENATED TALLOW ACID
C3818711|T121|1535492|RXNORM|HUMULUS LUPULUS WHOLE EXTRACT|HUMULUS LUPULUS WHOLE EXTRACT
C3818697|T121|1536454|RXNORM|TABEBUIA IMPETIGINOSA LEAF EXTRACT|TABEBUIA IMPETIGINOSA LEAF EXTRACT
C1654733|T121|606253|RXNORM|GLIMEPIRIDE / ROSIGLITAZONE|GLIMEPIRIDE / ROSIGLITAZONE
C2929624|T121|1008725|RXNORM|CALCIUM IODIZED / PEPTONE,DRIED / THYROID (USP)|CALCIUM IODIZED / PEPTONE,DRIED / THYROID (USP)
C3256648|T121|1358898|RXNORM|PORTULACA OLERACEA WHOLE EXTRACT|PORTULACA OLERACEA WHOLE EXTRACT
C0599532|T121|154876|RXNORM|THIOPHENE|THIOPHENE
C0886584|T121|266604|RXNORM|METYROSINE|METYROSINE
C0060243|T197|24910|RXNORM|FERRIC PHOSPHATE|FERRIC PHOSPHATE
C3643346|T121|1424267|RXNORM|SEMECARPUS ANACARDIUM FRUIT EXTRACT|SEMECARPUS ANACARDIUM FRUIT EXTRACT
C1367202|T129|1094833|RXNORM|IPILIMUMAB|IPILIMUMAB
C1165353|T121|349730|RXNORM|ANHYDROUS DEXTROSE|ANHYDROUS DEXTROSE
C0717703|T121|214502|RXNORM|DICLOFENAC / MISOPROSTOL|DICLOFENAC / MISOPROSTOL
C3485010|T121|1358896|RXNORM|FORSYTHIA SUSPENSA WHOLE EXTRACT|FORSYTHIA SUSPENSA WHOLE EXTRACT
C0029904|T121|7762|RXNORM|OUABAIN|OUABAIN
C0078814|T197|39972|RXNORM|ZIRCONIUM OXIDE|ZIRCONIUM OXIDE
C0717708|T121|214507|RXNORM|DILTIAZEM / ENALAPRIL|DILTIAZEM / ENALAPRIL
C3255612|T121|1358890|RXNORM|TREMELLA FUCIFORMIS FRUITING BODY EXTRACT|TREMELLA FUCIFORMIS FRUITING BODY EXTRACT
C3488424|T121|1309735|RXNORM|ARISTOLOCHIA CLEMATITIS ROOT EXTRACT|ARISTOLOCHIA CLEMATITIS ROOT EXTRACT
C0605984|T121|159085|RXNORM|HEXADECANAMIDE|HEXADECANAMIDE
C0035839|T121|1535498|RXNORM|RONIDAZOLE|RONIDAZOLE
C0246689|T121|73044|RXNORM|REPAGLINIDE|REPAGLINIDE
C2701396|T129|852197|RXNORM|GRAMA GRASS POLLEN EXTRACT|BOUTELOUA GRACILIS POLLEN EXTRACT
C2701701|T129|852627|RXNORM|SWEET GUM POLLEN EXTRACT|LIQUIDAMBAR STYRACIFLUA POLLEN EXTRACT
C2701392|T129|852193|RXNORM|WHITE HICKORY POLLEN EXTRACT|CARYA ALBA POLLEN EXTRACT
C2701697|T129|852622|RXNORM|PRIVET POLLEN EXTRACT|LIGUSTRUM VULGARE POLLEN EXTRACT
C3692850|T130|1442708|RXNORM|NATURAL RED 26|NATURAL RED 26
C3700992|T121|1486325|RXNORM|CAMPHOR / LEVOMENTHOL / METHYL SALICYLATE|CAMPHOR / LEVOMENTHOL / METHYL SALICYLATE
C0065185|T121|28894|RXNORM|LORMETAZEPAM|LORMETAZEPAM
C3486582|T121|1348449|RXNORM|MYOSOTIS ARVENSIS EXTRACT|FORGET-ME-NOT EXTRACT
C0054138|T121|19777|RXNORM|BROMPERIDOL|BROMPERIDOL
C2709742|T129|854938|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 14 VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 14 VACCINE
C2709740|T129|854936|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 12F VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 12F VACCINE
C0021734|T129|5879|RXNORM|INTERFERON ALFA-2A|INTERFERON ALFA-2A
C2709736|T129|854932|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 10A VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 10A VACCINE
C0043047|T197|11295|RXNORM|WATER|WATER
C0043047|T197|11295|RXNORM|WATER|WATER
C0043047|T197|11295|RXNORM|WATER|WATER
C0043047|T197|11295|RXNORM|WATER|WATER
C2701729|T129|852673|RXNORM|BAHIA GRASS POLLEN EXTRACT|PASPALUM NOTATUM POLLEN EXTRACT
C3256598|T109|1425982|RXNORM|C20-40 ACID|C20-40 ACID
C0013615|T121|3752|RXNORM|EDROPHONIUM|EDROPHONIUM
C0013618|T121|3755|RXNORM|EDETIC ACID|EDETIC ACID
C0072651|T130|1426464|RXNORM|D&C GREEN NO. 8|D&C GREEN NO. 8
C0007559|T195|2191|RXNORM|CEFTAZIDIME|CEFTAZIDIME
C0007560|T195|2192|RXNORM|CEFTIZOXIME|CEFTIZOXIME
C0007561|T195|2193|RXNORM|CEFTRIAXONE|CEFTRIAXONE
C0007562|T195|2194|RXNORM|CEFUROXIME|CEFUROXIME
C0067748|T121|1426463|RXNORM|N-ACETYL-METHIONINE|N-ACETYLMETHIONINE
C0165703|T121|60245|RXNORM|IMIDAPRIL|IMIDAPRIL
C0597277|T196|1318915|RXNORM|POTASSIUM ION|POTASSIUM ION
C0016971|T121|4638|RXNORM|GALLAMINE|GALLAMINE
C0069592|T130|1426468|RXNORM|D&C ORANGE NO. 4|D&C ORANGE NO. 4
C3486644|T121|1426469|RXNORM|ANTI-INTERLEUKIN-1.ALPHA. IMMUNOGLOBULIN G RABBIT|ANTI-INTERLEUKIN-1.ALPHA. IMMUNOGLOBULIN G RABBIT
C0993639|T109|317702|RXNORM|ROSMARINUS OFFICINALIS PREPARATION|ROSMARINUS OFFICINALIS PREPARATION
C0068314|T195|31435|RXNORM|ALLERGENIC EXTRACT, CURVULARIA LUNATA MOLD|VALRUBICIN
C0122922|T196|1483317|RXNORM|HYPOCHLORITE|HYPOCHLORITE
C0068314|T195|31435|RXNORM|ALLERGENIC EXTRACT, COTTONWOOD, WESTERN|VALRUBICIN
C0068314|T195|31435|RXNORM|ALLERGENIC EXTRACT, DUST, AUTOGENOUS|VALRUBICIN
C2702346|T129|854025|RXNORM|CANIS LUPUS FAMILIARIS HAIR EXTRACT|CANIS LUPUS FAMILIARIS HAIR EXTRACT
C1703206|T121|618974|RXNORM|4-AMINOBENZOATE|4-AMINOBENZOATE
C0053931|T197|19596|RXNORM|BONE MEAL|BONE MEAL
C1703665|T121|618970|RXNORM|CANRENOATE|CANRENOATE
C0055477|T121|20890|RXNORM|LORNOXICAM|LORNOXICAM
C0055478|T121|20891|RXNORM|CHLORTHENOXAZIN|CHLORTHENOXAZIN
C0070619|T130|1367159|RXNORM|PHENYLACETALDEHYDE|PHENYLACETALDEHYDE
C2930029|T121|1009134|RXNORM|AMBROXOL / THEOPHYLLINE|AMBROXOL / THEOPHYLLINE
C3255966|T109|1367152|RXNORM|PEG-12 DIMETHICONE (300 CST)|PEG-12 DIMETHICONE (300 CST)
C0075476|T109|1367150|RXNORM|SUCROSE PALMITATE|SUCROSE PALMITATE
C0066237|T109|1367156|RXNORM|METHYL CINNAMATE|METHYL CINNAMATE
C0066223|T109|1367155|RXNORM|METHYL ACRYLATE|METHYL ACRYLATE
C0074246|T121|36314|RXNORM|SECNIDAZOLE|SECNIDAZOLE
C2193984|T121|817612|RXNORM|BROMPHENIRAMINE / GUAIFENESIN / HYDROCODONE|BROMPHENIRAMINE / GUAIFENESIN / HYDROCODONE
C0000983|T130|168|RXNORM|ACETIC ACID|ACETIC ACID
C0000983|T130|168|RXNORM|ACETIC ACID|ACETIC ACID
C0000983|T130|168|RXNORM|ACETIC ACID|ACETIC ACID
C0021544|T121|5832|RXNORM|INOSINIC ACID|INOSINIC ACID
C0000975|T121|164|RXNORM|ACETATE|ACETATE
C0000981|T121|167|RXNORM|ACETAZOLAMIDE|ACETAZOLAMIDE
C0000970|T121|161|RXNORM|ACETAMINOPHEN|ACETAMINOPHEN
C0000973|T121|162|RXNORM|ACETANILIDE|ACETANILIDE
C0086140|T121|42635|RXNORM|DEXTRAN|DEXTRAN
C1828194|T121|687386|RXNORM|IBUPROFEN / LEVOMENTHOL|IBUPROFEN / LEVOMENTHOL
C0947604|T121|287513|RXNORM|BLUE COHOSH EXTRACT|BLUE COHOSH EXTRACT
C2930027|T121|1009132|RXNORM|ALLANTOIN / CHLOROCRESOL / NEOMYCIN|ALLANTOIN / CHLOROCRESOL / NEOMYCIN
C0981888|T129|894795|RXNORM|GRAIN MILL DUST ALLERGENIC EXTRACT|GRAIN MILL DUST ALLERGENIC EXTRACT
C2740731|T129|899611|RXNORM|BLUE BEECH POLLEN EXTRACT|CARPINUS CAROLINIANA POLLEN EXTRACT
C0085170|T121|42328|RXNORM|ASTEMIZOLE|ASTEMIZOLE
C0085161|T195|42322|RXNORM|FLEROXACIN|FLEROXACIN
C0068942|T121|31945|RXNORM|NONIVAMIDE|NONIVAMIDE
C3505633|T121|1358981|RXNORM|CAMPHOR / DIMETHICONE / MENTHOL / PHENOL|CAMPHOR / DIMETHICONE / MENTHOL / PHENOL
C2146603|T121|821601|RXNORM|ACETAMINOPHEN / ASPIRIN / CAFFEINE / CODEINE|ACETAMINOPHEN / ASPIRIN / CAFFEINE / CODEINE
C1260298|T195|384455|RXNORM|TIGECYCLINE|TIGECYCLINE
C3500830|T121|1356130|RXNORM|SIMABA CEDRON SEED EXTRACT|SIMABA CEDRON SEED EXTRACT
C0982277|T121|314726|RXNORM|MENTHOL / PHENOL|MENTHOL / PHENOL
C3500832|T121|1356132|RXNORM|2-(3-OXAZOLIDINYL)ETHYL METHACRYLATE|2-(3-OXAZOLIDINYL)ETHYL METHACRYLATE
C3500833|T121|1356133|RXNORM|C12-15 ALKYL LACTATE|C12-15 ALKYL LACTATE
C3500834|T121|1356134|RXNORM|CAPRYLIC-CAPRIC-SUCCINIC TRIGLYERCIDE|CAPRYLIC-CAPRIC-SUCCINIC TRIGLYERCIDE
C0039542|T121|10368|RXNORM|TERBUTALINE|TERBUTALINE
C0039542|T121|10368|RXNORM|TERBUTALINE|TERBUTALINE
C0039542|T121|10368|RXNORM|TERBUTALINE|TERBUTALINE
C3500836|T121|1356136|RXNORM|HYDROXYPROPYL CELLULOSE (TYPE E)|HYDROXYPROPYL CELLULOSE (80000 MW)
C3500837|T121|1356137|RXNORM|HYDROXYPROPYL CELLULOSE (TYPE L)|HYDROXYPROPYL CELLULOSE (120000 MW)
C2927385|T129|1005931|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-VICTORIA-210-2009 X-187 (H3N2) (A-PERTH-16-2009) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-VICTORIA-210-2009 X-187 (H3N2) (A-PERTH-16-2009) STRAIN
C3500838|T109|1356139|RXNORM|PEG-25 HYDROGENATED CASTOR OIL|PEG-25 HYDROGENATED CASTOR OIL
C0039512|T121|10362|RXNORM|TENIPOSIDE|TENIPOSIDE
C2927840|T121|1006916|RXNORM|BENZOCAINE / ISOPROPYL ALCOHOL|BENZOCAINE / ISOPROPYL ALCOHOL
C2927841|T121|1006917|RXNORM|ESTROGENS, CONJUGATED (USP) / MEDROXYPROGESTERONE|ESTROGENS, CONJUGATED (USP) / MEDROXYPROGESTERONE
C2927838|T121|1006914|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL / FERROUS FUMARATE|CALCIUM CARBONATE / CHOLECALCIFEROL / FERROUS FUMARATE
C2927839|T121|1006915|RXNORM|POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY) / POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1) / POLIOVIRUS VACCINE INACTIVATED, TYPE 3 (SAUKETT)|POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY) / POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1) / POLIOVIRUS VACCINE INACTIVATED, TYPE 3 (SAUKETT)
C2927836|T121|1006912|RXNORM|BENZOCAINE / PHENYLPROPANOLAMINE|BENZOCAINE / PHENYLPROPANOLAMINE
C2927837|T121|1006913|RXNORM|BIOTIN / DICALCIUM PHOSPHATE|BIOTIN / DICALCIUM PHOSPHATE
C2927834|T121|1006910|RXNORM|CALCIUM PHOSPHATE / VITAMIN D|CALCIUM PHOSPHATE / VITAMIN D
C2927835|T121|1006911|RXNORM|BENZOATE / SALICYLIC ACID|BENZOATE / SALICYLIC ACID
C3535892|T109|1370589|RXNORM|POLACRILLIN|POLACRILLIN
C2927842|T121|1006918|RXNORM|INTRINSIC FACTOR / VITAMIN B 12|INTRINSIC FACTOR / VITAMIN B 12
C2927843|T121|1006919|RXNORM|CAPSICUM OLEORESIN / TURPENTINE|CAPSICUM OLEORESIN / TURPENTINE
C2929964|T121|1009069|RXNORM|ESTROGENS, CONJUGATED (USP) / NORGESTREL|ESTROGENS, CONJUGATED (USP) / NORGESTREL
C2929963|T121|1009068|RXNORM|DEXPANTHENOL / PROCAINE|DEXPANTHENOL / PROCAINE
C0023024|T121|6227|RXNORM|LANOLIN|LANOLIN
C0771492|T121|236238|RXNORM|BURDOCK ROOT EXTRACT|BURDOCK ROOT EXTRACT
C0771880|T121|236587|RXNORM|THENOATE LITHIUM|THENOATE LITHIUM
C2929958|T121|1009063|RXNORM|BISMUTH / PECTIN|BISMUTH / PECTIN
C2929957|T121|1009062|RXNORM|DICHLORODIFLUOROMETHANE / TRICHLOROTRIFLUOROETHANE|DICHLORODIFLUOROMETHANE / TRICHLOROTRIFLUOROETHANE
C2929956|T121|1009061|RXNORM|CHOLINE / GINKGO BILOBA EXTRACT / VITAMIN B 12 / VITAMIN B6|CHOLINE / GINKGO BILOBA EXTRACT / VITAMIN B 12 / VITAMIN B6
C2929955|T121|1009060|RXNORM|BECLOMETHASONE / CLIOQUINOL|BECLOMETHASONE / CLIOQUINOL
C2929962|T121|1009067|RXNORM|BENZOCAINE / DIOSMIN|BENZOCAINE / DIOSMIN
C2929961|T121|1009066|RXNORM|BORIC ACID / CHLOROCRESOL / ZINC OXIDE|BORIC ACID / CHLOROCRESOL / ZINC OXIDE
C2929960|T121|1009065|RXNORM|PHLOROGLUCINOL / TRIMETHYLPHLOROGLUCINOL|PHLOROGLUCINOL / TRIMETHYLPHLOROGLUCINOL
C2929959|T121|1009064|RXNORM|DIOSMIN / HESPERIDIN|DIOSMIN / HESPERIDIN
C0052793|T121|402580|RXNORM|AZINTAMIDE|AZINTAMIDE
C1322002|T121|402583|RXNORM|CLOCINIZINE|CLOCINIZINE
C0002555|T121|677|RXNORM|AMINOGLUTETHIMIDE|AMINOGLUTETHIMIDE
C0021528|T121|1483575|RXNORM|INOSINE|INOSINE
C1322006|T121|402587|RXNORM|DIFETARSONE|DIFETARSONE
C0049289|T121|15842|RXNORM|5-METHOXYPSORALEN|BERGAPTEN
C0076799|T121|38377|RXNORM|TOLFENAMIC ACID|TOLFENAMIC ACID
C0164386|T121|59636|RXNORM|BUCLIZINE|BUCLIZINE
C0205679|T197|1425919|RXNORM|MONTMORRILLONITE|MONTMORRILLONITE
C2929889|T121|1008994|RXNORM|ALLOIN / APIOLE / ERGOT PREPARATION|ALLOIN / APIOLE / ERGOT PREPARATION
C0147942|T130|1546223|RXNORM|DIATRIZOIC ACID|DIATRIZOIC ACID
C0040377|T121|10636|RXNORM|TOLMETIN|TOLMETIN
C1874806|T121|689380|RXNORM|CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE|CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE
C3531167|T121|1366200|RXNORM|DIMETHYL SULFOXIDE / FLUOCINOLONE|DIMETHYL SULFOXIDE / FLUOCINOLONE
C3256303|T130|1425913|RXNORM|FD&C RED #40 HT ALUMINUM LAKE|FD&C RED #40 HT ALUMINUM LAKE
C1874808|T121|689383|RXNORM|CHLORPHENIRAMINE / CODEINE / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / CODEINE / PHENYLPROPANOLAMINE
C3256165|T130|1425915|RXNORM|FD&C YELLOW #5 ALUMINUM LAKE|FD&C YELLOW #5 ALUMINUM LAKE
C2929891|T121|1008996|RXNORM|BILE SALTS / PANCREATIN / PEPSIN A|BILE SALTS / PANCREATIN / PEPSIN A
C1874810|T121|689387|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE|CHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE
C0040373|T121|10634|RXNORM|TOLAZOLINE|TOLAZOLINE
C3464512|T121|1312621|RXNORM|LAURYL ALDEHYDE|LAURYL ALDEHYDE
C0057919|T121|1362911|RXNORM|DIETHANOLAMINE|DIETHANOLAMINE
C2929885|T121|1008990|RXNORM|DEXTROMETHORPHAN / GUAIACOLSULFONIC ACID / PHENYLEPHRINE|DEXTROMETHORPHAN / GUAIACOLSULFONIC ACID / PHENYLEPHRINE
C3256117|T109|1362913|RXNORM|ISODODECANE|ISODODECANE
C3249694|T121|1233303|RXNORM|DEXTRAN 70 / POLYETHYLENE GLYCOLS|DEXTRAN 70 / POLYETHYLENE GLYCOLS
C0033684|T123|8859|RXNORM|PROTEINS|PROTEINS
C0023582|T121|6377|RXNORM|LEVOPROPOXYPHENE|LEVOPROPOXYPHENE
C2731519|T129|895515|RXNORM|HORSE HAIR EXTRACT|HORSE HAIR EXTRACT
C2928923|T121|1008012|RXNORM|VITAMIN B 12 / VITAMIN B6|VITAMIN B 12 / VITAMIN B6
C0165032|T121|59943|RXNORM|IMIQUIMOD|IMIQUIMOD
C3495434|T121|1363352|RXNORM|HYDROXYETHYL STARCH 130-0.4|HYDROXYETHYL STARCH 130-0.4
C0318392|T005|1427210|RXNORM|HUMAN COXSACKIEVIRUS B4|HUMAN COXSACKIEVIRUS B4
C0019169|T005|1427211|RXNORM|HEPATITIS B VIRUS|HEPATITIS B VIRUS
C0206435|T005|1427212|RXNORM|HUMAN POLIOVIRUS|HUMAN POLIOVIRUS
C3474579|T121|1427215|RXNORM|AMODIMETHICONE (800 CST)|AMODIMETHICONE (800 CST)
C3486807|T121|1427216|RXNORM|SCABIES LESION LYSATE (HUMAN)|PSORINUM LESION LYSATE (HUMAN)
C0076184|T121|37855|RXNORM|TESTOSTERONE 17-PHENYLPROPIONATE|TESTOSTERONE 17-PHENYLPROPIONATE
C3464494|T121|1427218|RXNORM|METHYLSILANOL ACETYLMETHIONATE|METHYLSILANOL ACETYLMETHIONATE
C3474401|T109|1427219|RXNORM|METHYLBENZYL ACETATE|METHYLBENZYL ACETATE
C0062619|T121|26826|RXNORM|HEXAFLUORENIUM|HEXAFLURONIUM
C2929588|T121|1008688|RXNORM|NITROFURANTOIN / SULFAMETHIZOLE|NITROFURANTOIN / SULFAMETHIZOLE
C2929589|T121|1008689|RXNORM|NAPROXEN / THIAMINE|NAPROXEN / THIAMINE
C3464708|T121|1305745|RXNORM|CHAMAECYPARIS OBTUSA LEAF EXTRACT|CHAMAECYPARIS OBTUSA LEAF EXTRACT
C3256216|T121|1305744|RXNORM|CYCLOMETHICONE 5|CYCLOMETHICONE 5
C2929580|T121|1008680|RXNORM|CHOLINE / THIAMINE|CHOLINE / THIAMINE
C2929581|T121|1008681|RXNORM|BENDROFLUMETHIAZIDE / MEPROBAMATE|BENDROFLUMETHIAZIDE / MEPROBAMATE
C2929582|T121|1008682|RXNORM|CALAMINE / RESORCINOL|CALAMINE / RESORCINOL
C2929583|T121|1008683|RXNORM|CHLORQUINALDOL / PROMESTRIENE|CHLORQUINALDOL / PROMESTRIENE
C2929584|T121|1008684|RXNORM|ASPIRIN / LITHIUM / QUININE|ASPIRIN / LITHIUM / QUININE
C2929585|T121|1008685|RXNORM|BENACTYZINE / BENORILATE|BENACTYZINE / BENORILATE
C2929586|T121|1008686|RXNORM|CYCLOBENZAPRINE / NIMESULIDE|CYCLOBENZAPRINE / NIMESULIDE
C1576794|T121|1426610|RXNORM|PEG-PPG-18-18-DIMETHICONE|PEG-PPG-18-18-DIMETHICONE
C2828292|T196|1546266|RXNORM|IODIDE I-125|IODIDE I-125
C3267307|T121|1355807|RXNORM|UNDARIA PINNATIFIDA EXTRACT|UNDARIA PINNATIFIDA EXTRACT
C2346521|T196|1546264|RXNORM|ZINC CATION|ZINC CATION
C3538087|T121|1371988|RXNORM|IODINE / LACTATE|IODINE / LACTATE
C3848576|T196|1546268|RXNORM|THIAMINE ION|THIAMINE ION
C2342732|T121|794252|RXNORM|DIHYDROCODEINE / GUAIFENESIN|DIHYDROCODEINE / GUAIFENESIN
C0072896|T121|35242|RXNORM|QUINUPRAMINE|QUINUPRAMINE
C0080225|T123|40230|RXNORM|THYMOPENTIN|THYMOPENTIN
C2723760|T129|867349|RXNORM|STEMPHYLIUM SOLANI EXTRACT|STEMPHYLIUM SOLANI EXTRACT
C0486268|T131|1371449|RXNORM|2,4-DICHLOROPHENOXYACETATE|2,4-DICHLOROPHENOXYACETATE
C3256551|T121|1313725|RXNORM|POLYBUTENE (1400 MW)|POLYBUTENE (1400 MW)
C0887175|T195|267073|RXNORM|METHICILLIN SODIUM|METHICILLIN SODIUM
C2723754|T130|867341|RXNORM|RED IMPORTED FIRE ANT ALLERGENIC EXTRACT|SOLENOPSIS INVICTA ALLERGENIC EXTRACT
C2052688|T121|1008532|RXNORM|PENICILLIN G PROCAINE / PENICILLIN G SODIUM|PENICILLIN G PROCAINE / PENICILLIN G SODIUM
C2929436|T121|1008533|RXNORM|COENZYME Q10 / RED YEAST RICE|COENZYME Q10 / RED YEAST RICE
C2929434|T121|1008530|RXNORM|GLYCERIN / POLYSORBATE 80|GLYCERIN / POLYSORBATE 80
C2929435|T121|1008531|RXNORM|MEASLES VACCINE / MUMPS VACCINE|MEASLES VACCINE / MUMPS VACCINE
C2929439|T121|1008536|RXNORM|BENZOCAINE / CHLOROXYLENOL / HYDROCORTISONE|BENZOCAINE / CHLOROXYLENOL / HYDROCORTISONE
C2929437|T121|1008534|RXNORM|BILBERRY EXTRACT / LUTEIN|BILBERRY EXTRACT / LUTEIN
C2929438|T121|1008535|RXNORM|GLYCERIN / PETROLATUM / PHENYLEPHRINE / PRAMOXINE|GLYCERIN / PETROLATUM / PHENYLEPHRINE / PRAMOXINE
C2740768|T129|899673|RXNORM|CINNAMON ALLERGENIC EXTRACT|CINNAMON ALLERGENIC EXTRACT
C0611561|T121|162901|RXNORM|SILVER MONO(2-AMINOETHYL)PHOSPHATE|SILVER MONO(2-AMINOETHYL)PHOSPHATE
C2929441|T121|1008538|RXNORM|ACETYLCARNITINE / CARNOSINE / COENZYME Q10|ACETYLCARNITINE / CARNOSINE / COENZYME Q10
C2929442|T121|1008539|RXNORM|CHLOPHEDIANOL / DEXBROMPHENIRAMINE / PHENYLEPHRINE|CHLOPHEDIANOL / DEXBROMPHENIRAMINE / PHENYLEPHRINE
C0076355|T121|37999|RXNORM|TETROXOPRIM|TETROXOPRIM
C3500697|T121|1315123|RXNORM|SNOW CRAB, UNSPECIFIED PREPARATION|SNOW CRAB, UNSPECIFIED PREPARATION
C0174883|T121|62130|RXNORM|CRESOL|CRESOL
C0064636|T121|28439|RXNORM|LAMOTRIGINE|LAMOTRIGINE
C0010682|T123|3036|RXNORM|CYSTINE|CYSTINE
C1113007|T121|324050|RXNORM|MENINGOCOCCAL VACCINE B|MENINGOCOCCAL VACCINE B
C0033228|T121|8703|RXNORM|FENOFIBRATE|FENOFIBRATE
C0304465|T121|91198|RXNORM|CITRIC ACID / SODIUM CITRATE|CITRIC ACID / SODIUM CITRATE
C0033218|T121|8701|RXNORM|PROCAINE|PROCAINE
C0033218|T121|8701|RXNORM|PROCAINE|PROCAINE
C0033216|T121|8700|RXNORM|PROCAINAMIDE|PROCAINAMIDE
C0071772|T197|34316|RXNORM|POTASSIUM NITRATE|POTASSIUM NITRATE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE|PROCHLORPERAZINE
C3256542|T121|1312615|RXNORM|ISODECETH-6|ISODECETH-6
C3464195|T109|1312614|RXNORM|IPOMOEA MAURITIANA TUBER EXTRACT|IPOMOEA MAURITIANA TUBER EXTRACT
C0071774|T197|34318|RXNORM|POTASSIUM PERCHLORATE|POTASSIUM PERCHLORATE
C3256544|T121|1312616|RXNORM|ISONIACINAMIDE|ISONIACINAMIDE
C2825385|T130|1312611|RXNORM|HYDROXYETHYLPIPERAZINE ETHANE SULFONIC ACID|HYDROXYETHYLPIPERAZINE ETHANE SULFONIC ACID
C3499813|T121|1312961|RXNORM|EUCALYPTUS OIL / TEA TREE OIL|EUCALYPTUS OIL / TEA TREE OIL
C2948572|T121|1044415|RXNORM|LANOLIN / ZINC OXIDE|LANOLIN / ZINC OXIDE
C0376266|T121|114203|RXNORM|FEVERFEW EXTRACT|TANACETUM PARTHENIUM EXTRACT
C0376259|T121|114200|RXNORM|CITRATE|CITRATE
C0068485|T121|31565|RXNORM|NEFAZODONE|NEFAZODONE
C0068483|T121|31563|RXNORM|NEDOCROMIL|NEDOCROMIL
C0068483|T121|31563|RXNORM|NEDOCROMIL|NEDOCROMIL
C0001052|T109|200|RXNORM|ACETYLENE|ACETYLENE
C3864821|T109|1597391|RXNORM|THIOCTIC ACID AMIDE|THIOCTIC ACID AMIDE
C3864822|T109|1597390|RXNORM|CARBOXYMETHYLCELLULOSE SODIUM (0.7 CARBOXYMETHYL SUBSTITUTION PER SACCHARIDE; 50-100 MPA.S AT 1% )|CARBOXYMETHYLCELLULOSE SODIUM (0.7 CARBOXYMETHYL SUBSTITUTION PER SACCHARIDE; 50-100 MPA.S AT 1% )
C2702319|T129|995707|RXNORM|EPIDERMOPHYTON FLOCCOSUM ALLERGENIC EXTRACT|EPIDERMOPHYTON FLOCCOSUM ALLERGENIC EXTRACT
C1577314|T109|486120|RXNORM|IRON FUMARATE|IRON FUMARATE
C1577317|T121|486126|RXNORM|ZICONOTIDE ACETATE|ZICONOTIDE ACETATE
C0299792|T121|89013|RXNORM|ARIPIPRAZOLE|ARIPIPRAZOLE
C2928712|T121|1007797|RXNORM|PANTOTHENIC ACID / SENNOSIDES, USP|PANTOTHENIC ACID / SENNOSIDES, USP
C2928711|T121|1007796|RXNORM|POTASSIUM CHLORIDE / RAUWOLFIA PREPARATION|POTASSIUM CHLORIDE / RAUWOLFIA PREPARATION
C2928710|T121|1007795|RXNORM|ASCORBIC ACID / FERROUS SULFATE / NIACIN / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B6 / VITAMIN D / VITAMIN E|ASCORBIC ACID / FERROUS SULFATE / NIACIN / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B6 / VITAMIN D / VITAMIN E
C2928709|T121|1007794|RXNORM|ECONAZOLE / ZINC OXIDE|ECONAZOLE / ZINC OXIDE
C2928708|T121|1007793|RXNORM|MINERAL OIL, LIGHT / PETROLATUM|MINERAL OIL, LIGHT / PETROLATUM
C2928707|T121|1007792|RXNORM|DEHYDROCHOLATE / DOCUSATE / PHENOLPHTHALEIN|DEHYDROCHOLATE / DOCUSATE / PHENOLPHTHALEIN
C2928706|T121|1007791|RXNORM|HYDROCODONE / PHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PYRILAMINE|HYDROCODONE / PHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PYRILAMINE
C3489039|T121|1322554|RXNORM|MERCURIALIS PERENNIS EXTRACT|MERCURIALIS PERENNIS EXTRACT
C2928713|T121|1007798|RXNORM|MINERAL OIL / PETROLATUM / PHENYLEPHRINE|MINERAL OIL / PETROLATUM / PHENYLEPHRINE
C3282507|T121|1426921|RXNORM|LENTIL SEED EXTRACT|LENTIL SEED EXTRACT
C3256726|T109|1426920|RXNORM|SARGASSUM FILIPENDULA EXTRACT|SARGASSUM FILIPENDULA EXTRACT
C3282110|T109|1426923|RXNORM|MENTHA PULEGIUM EXTRACT|MENTHA PULEGIUM EXTRACT
C1875141|T121|691395|RXNORM|EUCALYPTUS OIL / MENTHOL|EUCALYPTUS OIL / MENTHOL
C3465015|T109|1426925|RXNORM|GLYCERYL 1-ADIPATE|GLYCERYL 1-ADIPATE
C2343848|T120|1426924|RXNORM|D&C VIOLET NO. 2|D&C VIOLET NO. 2
C3268188|T122|1426927|RXNORM|GLYCERYL ABIETATE|GLYCERYL ABIETATE
C0379199|T121|115264|RXNORM|IBANDRONATE|IBANDRONATE
C3257703|T109|1314305|RXNORM|TRIDECETH-10|TRIDECETH-10
C3267229|T121|1314304|RXNORM|DIMETHYL CAPRAMIDE|DIMETHYL CAPRAMIDE
C0043406|T007|1426679|RXNORM|YERSINIA ENTEROCOLITICA|YERSINIA ENTEROCOLITICA
C3497607|T121|1313709|RXNORM|HYDROGENATED PALM KERNEL GLYCERIDES|HYDROGENATED PALM KERNEL GLYCERIDES
C3530629|T121|1364988|RXNORM|FICUS CARICA WHOLE EXTRACT|FICUS CARICA WHOLE EXTRACT
C3530630|T121|1364989|RXNORM|ROSA CENTIFOLIA FLOWER EXTRACT|ROSA CENTIFOLIA FLOWER EXTRACT
C3256241|T122|1313700|RXNORM|METHYLCELLULOSE (1500 CPS)|METHYLCELLULOSE (1500 CPS)
C3256242|T121|1313701|RXNORM|METHYLCELLULOSE (25 CPS)|METHYLCELLULOSE (25 CPS)
C3255823|T121|1313702|RXNORM|METHYLCELLULOSE (400 CPS)|METHYLCELLULOSE (400 CPS)
C3255652|T109|1313703|RXNORM|CETYL HYDROXYETHYLCELLULOSE (350000 MW)|CETYL HYDROXYETHYLCELLULOSE (350000 MW)
C3255760|T121|1313704|RXNORM|ETHYLCELLULOSE (10 MPA.S)|ETHYLCELLULOSE (10 MPA.S)
C3256611|T121|1313705|RXNORM|DODECYL BENZOATE|DODECYL BENZOATE
C3489289|T121|1309949|RXNORM|STRYCHNOS WALLICHIANA BARK EXTRACT|STRYCHNOS WALLICHIANA BARK EXTRACT
C2605128|T109|1313707|RXNORM|3,7-DIMETHYLOCTANE-1,7-DIOL|3,7-DIMETHYLOCTANE-1,7-DIOL
C3833239|T109|1540881|RXNORM|HYDROGENATED JOJOBA OIL, RANDOMIZED|HYDROGENATED JOJOBA OIL, RANDOMIZED
C3474077|T121|1314309|RXNORM|OCIMUM BASILICUM WHOLE EXTRACT|OCIMUM BASILICUM WHOLE EXTRACT
C3833240|T109|1540882|RXNORM|GLYCOLIDE|GLYCOLIDE
C1959896|T121|729601|RXNORM|MUCINS / XYLITOL|MUCINS / XYLITOL
C2138496|T121|812238|RXNORM|CROMOLYN / XYLOMETAZOLINE|CROMOLYN / XYLOMETAZOLINE
C3465032|T121|1314308|RXNORM|METHYLSILANOL ASCORBATE|METHYLSILANOL ASCORBATE
C3555463|T121|1420981|RXNORM|SENNA ALATA WHOLE EXTRACT|SENNA ALATA WHOLE EXTRACT
C2073893|T121|812237|RXNORM|CHLORPHENIRAMINE / PYRILAMINE|CHLORPHENIRAMINE / PYRILAMINE
C0388844|T121|1420983|RXNORM|ETHYL FERULATE|ETHYL FERULATE
C0041964|T121|1420982|RXNORM|URETHANE|URETHANE
C2116318|T121|812232|RXNORM|PILOCARPINE / TIMOLOL|PILOCARPINE / TIMOLOL
C3485572|T121|1310076|RXNORM|PHYSOSTIGMA VENENOSUM SEED EXTRACT|PHYSOSTIGMA VENENOSUM SEED EXTRACT
C2928343|T121|1007421|RXNORM|VITAMIN B6 / ZINC GLUCONATE|VITAMIN B6 / ZINC GLUCONATE
C2928342|T121|1007420|RXNORM|LACTATE / ZINC GLUCONATE|LACTATE / ZINC GLUCONATE
C2928345|T121|1007423|RXNORM|DEXAMETHASONE / OXYTETRACYCLINE|DEXAMETHASONE / OXYTETRACYCLINE
C2928344|T121|1007422|RXNORM|CHLORAMPHENICOL / ICTASOL|CHLORAMPHENICOL / ICTASOL
C2928347|T121|1007425|RXNORM|FLUFENAMIC ACID / HEPARINOIDS / SALICYLIC ACID|FLUFENAMIC ACID / HEPARINOIDS / SALICYLIC ACID
C2928346|T121|1007424|RXNORM|ASCORBIC ACID / ASPIRIN / DIPHENYLPYRALINE|ASCORBIC ACID / ASPIRIN / DIPHENYLPYRALINE
C2928349|T121|1007427|RXNORM|PANGAMIC ACID / PROCAINE|PANGAMIC ACID / PROCAINE
C2928348|T121|1007426|RXNORM|HEXYLRESORCINOL / LAURETH-9|HEXYLRESORCINOL / POLIDOCANOL
C2928351|T121|1007429|RXNORM|CAFFEINE / PROCAINE|CAFFEINE / PROCAINE
C2928350|T121|1007428|RXNORM|ACETAMINOPHEN / PHENYLEPHRINE / TERFENADINE|ACETAMINOPHEN / PHENYLEPHRINE / TERFENADINE
C3255776|T121|1307660|RXNORM|LYCIUM CHINENSE ROOT BARK EXTRACT|LYCIUM CHINENSE ROOT BARK EXTRACT
C0795571|T121||RXNORM|AMPHETAMINE / DEXTROAMPHETAMINE
C3255609|T121|1307667|RXNORM|PULSATILLA KOREANA ROOT EXTRACT|PULSATILLA KOREANA ROOT EXTRACT
C3256342|T121|1307664|RXNORM|ANGELICA GIGAS ROOT EXTRACT|ANGELICA GIGAS ROOT EXTRACT
C3268108|T121|1307665|RXNORM|PRUNUS DULCIS BARK EXTRACT|PRUNUS DULCIS BARK EXTRACT
C3818723|T109|1535221|RXNORM|KALANCHOE DAIGREMONTIANA LEAF EXTRACT|KALANCHOE DAIGREMONTIANA LEAF EXTRACT
C2080527|T121|819002|RXNORM|ACETAMINOPHEN / DIPHENHYDRAMINE / GUAIFENESIN / PHENYLEPHRINE|ACETAMINOPHEN / DIPHENHYDRAMINE / GUAIFENESIN / PHENYLEPHRINE
C0061446|T121|1535222|RXNORM|GLUCURONOLACTONE|GLUCURONOLACTONE
C1874662|T121|691025|RXNORM|CALCIUM CITRATE / VITAMIN A / VITAMIN D|CALCIUM CITRATE / VITAMIN A / VITAMIN D
C1874664|T121|691027|RXNORM|CALCIUM CREOSOTATE / IODINE|CALCIUM CREOSOTATE / IODINE
C3858051|T121|1591942|RXNORM|LEDIPASVIR / SOFOSBUVIR|LEDIPASVIR / SOFOSBUVIR
C3256789|T109|1309448|RXNORM|NELUMBO NUCIFERA SEED EXTRACT|NELUMBO NUCIFERA SEED EXTRACT
C0075477|T121|1363060|RXNORM|SUCROSE MONOSTEARATE|SUCROSE MONOSTEARATE
C3505293|T121|1358207|RXNORM|MEDRONATE|MEDRONATE
C0076141|T109|1363061|RXNORM|TERT-BUTYL ALCOHOL|TERT-BUTYL ALCOHOL
C0082286|T121|3142|RXNORM|ACETIC|DEHYDROEMETINE
C1620287|T121|613391|RXNORM|PRASUGREL|PRASUGREL
C0981814|T130|314299|RXNORM|ALBUMIN,CHROMATED CR-51 SERUM|ALBUMIN,CHROMATED CR-51 SERUM
C0981813|T121|314298|RXNORM|ADRENOCORTICOTROPIN (ACTH 1-18),I-125 (TYR)|ADRENOCORTICOTROPIN (ACTH 1-18),I-125 (TYR)
C3256368|T109|1309444|RXNORM|MORUS ALBA BARK EXTRACT|MORUS ALBA BARK EXTRACT
C3854888|T109|1546870|RXNORM|CETEARETH-10 PHOSPHATE|CETEARETH-10 PHOSPHATE
C2351138|T121|1426432|RXNORM|POLYOXYL 40 STEARATE|POLYOXYL 40 STEARATE
C3640212|T129|1440046|RXNORM|LIPEGFILGRASTIM|LIPEGFILGRASTIM
C3257238|T121|1426431|RXNORM|MACROCYSTIS PYRIFERA EXTRACT|MACROCYSTIS PYRIFERA EXTRACT
C3256640|T109|1426430|RXNORM|POLYMETHYLSILSESQUIOXANE (4.5 MICRONS)|POLYMETHYLSILSESQUIOXANE (4.5 MICRONS)
C0025424|T196|6769|RXNORM|MERCURY|MERCURY
C0062585|T121|1314255|RXNORM|HESPERETIN|HESPERETIN
C3499864|T121|1313054|RXNORM|MYRISTOYL PENTAPEPTIDE-4|MYRISTOYL PENTAPEPTIDE-4
C0025405|T121|6765|RXNORM|TIOPRONIN|TIOPRONIN
C0756081|T195|229367|RXNORM|QUINUPRISTIN|QUINUPRISTIN
C0025397|T121|6762|RXNORM|MERBROMIN|MERBROMIN
C0025387|T121|6761|RXNORM|MEPTAZINOL|MEPTAZINOL
C0025386|T121|6760|RXNORM|MEPROBAMATE|MEPROBAMATE
C1636662|T121|608054|RXNORM|FUROSEMIDE / POTASSIUM CHLORIDE|FUROSEMIDE / POTASSIUM CHLORIDE
C0054425|T121|20024|RXNORM|CERULETIDE DIETHYLAMINE|CERULETIDE DIETHYLAMINE
C2701482|T129|852298|RXNORM|GUINEA PIG SKIN EXTRACT|CAVIA PORCELLUS DANDER PREPARATION
C0063088|T197|1366859|RXNORM|HYDROGEN SULFITE|HYDROGEN SULFITE
C2701478|T129|852294|RXNORM|WHITE OAK POLLEN EXTRACT|QUERCUS ALBA POLLEN EXTRACT
C0142785|T121|56443|RXNORM|SODIUM ACETATE|SODIUM ACETATE
C1874821|T121|689401|RXNORM|CHLORPHENIRAMINE / GUAIFENESIN / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / GUAIFENESIN / PHENYLPROPANOLAMINE
C2702424|T129|892599|RXNORM|BEEF ALLERGENIC EXTRACT|BEEF ALLERGENIC EXTRACT
C0050458|T121|16735|RXNORM|ACETOPHENAZINE|ACETOPHENAZINE
C2726148|T129|972601|RXNORM|EGGPLANT ALLERGENIC EXTRACT|EGGPLANT ALLERGENIC EXTRACT
C3244974|T121|1190048|RXNORM|CHLORCYCLIZINE / PHENYLEPHRINE|CHLORCYCLIZINE / PHENYLEPHRINE
C0143961|T121|56790|RXNORM|SUCCINYLATED GELATIN|SUCCINYLATED GELATIN
C2939723|T129|1013913|RXNORM|SCRUB PINE POLLEN EXTRACT|PINUS VIRGINIANA POLLEN EXTRACT
C0054275|T121|19900|RXNORM|BUTYL CHLORIDE|BUTYL CHLORIDE
C3669133|T121|1442997|RXNORM|DICTYOPTERIS POLYPODIOIDES EXTRACT|DICTYOPTERIS POLYPODIOIDES EXTRACT
C0303835|T130|1435572|RXNORM|N-BUTYL LACTATE|N-BUTYL LACTATE
C3818808|T121|1489920|RXNORM|ROSA MULTIFLORA FLOWER WAX|ROSA MULTIFLORA FLOWER WAX
C3818807|T121|1489921|RXNORM|EICOSYL POVIDONE (2 EICOSYL BRANCHES-REPEAT)|EICOSYL POVIDONE (2 EICOSYL BRANCHES-REPEAT)
C2194312|T121|813187|RXNORM|CAFFEINE / DIMENHYDRINATE / ERGOTAMINE|CAFFEINE / DIMENHYDRINATE / ERGOTAMINE
C3255922|T109|1306154|RXNORM|CITRUS MAXIMA FRUIT RIND OIL|CITRUS MAXIMA FRUIT RIND OIL
C1317494|T121|714785|RXNORM|ISOLEUCINE / LEUCINE / VALINE|ISOLEUCINE / LEUCINE / VALINE
C3819170|T121|1489929|RXNORM|PALMITAMIDOPROPYLTRIMONIUM|PALMITAMIDOPROPYLTRIMONIUM
C1638413|T121|608349|RXNORM|CALCIUM PHOSPHATE / CHOLECALCIFEROL|CALCIUM PHOSPHATE / CHOLECALCIFEROL
C3256152|T109|1306138|RXNORM|CRAMBE HISPANICA SUBSP. ABYSSINICA SEED OIL|CRAMBE HISPANICA SUBSP. ABYSSINICA SEED OIL
C0037473|T196|9853|RXNORM|SODIUM|SODIUM
C2726357|T121|1312707|RXNORM|POLYETHYLENE GLYCOL 3500|POLYETHYLENE GLYCOL 3500
C3255926|T109|1306131|RXNORM|CITRUS RETICULATA FRUIT OIL|CITRUS RETICULATA FRUIT OIL
C3256844|T109|1306130|RXNORM|GRAPEFRUIT SEED OIL|GRAPEFRUIT SEED OIL
C3255928|T109|1306133|RXNORM|CITRUS SINENSIS FLOWER OIL|CITRUS SINENSIS FLOWER OIL
C3255927|T109|1306132|RXNORM|CITRUS RETICULATA LEAF OIL|CITRUS RETICULATA LEAF OIL
C3256141|T109|1306135|RXNORM|COLEUS FORSKOHLII ROOT OIL|COLEUS FORSKOHLII ROOT OIL
C3256022|T109|1306134|RXNORM|CLADANTHUS MIXTUS FLOWER VOLATILE OIL|CLADANTHUS MIXTUS FLOWER VOLATILE OIL
C3256151|T109|1306137|RXNORM|CORYMBIA CITRIODORA LEAF OIL|CORYMBIA CITRIODORA LEAF OIL
C3256143|T109|1306136|RXNORM|COPIBA OIL|COPAIBA OIL
C1509513|T121|1427180|RXNORM|GENTISIC ACID ETHANOLAMIDE|GENTISIC ACID ETHANOLAMIDE
C3645276|T121|1427185|RXNORM|OCTADECENEDIOATE|OCTADECENEDIOATE
C2354965|T109|1427186|RXNORM|LAURYL PEG-PPG-18-18 METHICONE|LAURYL PEG-PPG-18-18 METHICONE
C3282683|T121|1427188|RXNORM|HYDROXYPHENYL PROPAMIDOBENZOIC ACID|HYDROXYPHENYL PROPAMIDOBENZOIC ACID
C3282458|T121|1427189|RXNORM|P-TERT-BUTYLPHENOL-FORMALDEHYDE RESIN (LOW MOLECULAR WEIGHT)|P-TERT-BUTYLPHENOL-FORMALDEHYDE RESIN (LOW MOLECULAR WEIGHT)
C1831796|T121|714438|RXNORM|PAZOPANIB|PAZOPANIB
C3858055|T121|1551411|RXNORM|9-FLUOROPREDNISOLONE / NEOMYCIN / TETRACAINE|ISOFLUPREDONE / NEOMYCIN / TETRACAINE
C2741510|T129|901329|RXNORM|RED BELL PEPPER ALLERGENIC EXTRACT|RED BELL PEPPER ALLERGENIC EXTRACT
C1720480|T121|645371|RXNORM|AMILORIDE / BUMETANIDE|AMILORIDE / BUMETANIDE
C2978884|T121|1089733|RXNORM|CHOLECALCIFEROL / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / VITAMIN E|CHOLECALCIFEROL / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / VITAMIN E
C1532485|T121|484259|RXNORM|IBUPROFEN / OXYCODONE|IBUPROFEN / OXYCODONE
C0008593|T121|2508|RXNORM|CHROMONAR|CHROMONAR
C0061632|T121|26051|RXNORM|GLYCOL SALICYLATE|GLYCOL SALICYLATE
C0115137|T197|49334|RXNORM|DURAPATITE|DURAPATITE
C0001143|T195|239|RXNORM|ACLARUBICIN|ACLARUBICIN
C1874579|T121|690610|RXNORM|BISMUTH SUBSALICYLATE / CALCIUM CARBONATE|BISMUTH SUBSALICYLATE / CALCIUM CARBONATE
C3529024|T121|1363985|RXNORM|ACTINIDIA CHINENSIS ROOT EXTRACT|ACTINIDIA CHINENSIS ROOT EXTRACT
C0077039|T131|38578|RXNORM|TRICHLOROFLUOROMETHANE|TRICHLOROMONOFLUOROMETHANE
C0146706|T109|1363986|RXNORM|TRIETHANOLAMINE LAURYL SULFATE|TRIETHANOLAMINE LAURYL SULFATE
C0208225|T121|1539968|RXNORM|ETHYL PYRUVATE|ETHYL PYRUVATE
C3832943|T121|1539969|RXNORM|QUATERNIUM-24|QUATERNIUM-24
C0077034|T121|38574|RXNORM|TRICHLOROACETALDEHYDE|TRICHLOROACETALDEHYDE
C2756406|T129|968114|RXNORM|WHITE-ROT FUNGUS EXTRACT|SPOROTRICHUM PRUINOSUM EXTRACT
C0036048|T168|9515|RXNORM|SAFFLOWER OIL|SAFFLOWER OIL
C0771139|T121|235935|RXNORM|DOBESILIC ACID|DOBESILIC ACID
C0036025|T004|9511|RXNORM|SACCHAROMYCES CEREVISIAE|SACCHAROMYCES CEREVISIAE
C0796396|T196|253341|RXNORM|IODINE-125|IODINE-125
C3832942|T121|1539967|RXNORM|DIOCTYLDIMONIUM CHLORIDE|DIOCTYLDIMONIUM CHLORIDE
C0303542|T196|90611|RXNORM|82 STRONTIUM|82 STRONTIUM
C0303544|T196|90613|RXNORM|85 STRONTIUM|85 STRONTIUM
C3255941|T121|1307311|RXNORM|HYDROLYZED JOJOBA ESTERS (ACID FORM)|HYDROLYZED JOJOBA ESTERS (ACID FORM)
C0036071|T121|9518|RXNORM|SALICYLAMIDE|SALICYLAMIDE
C2740655|T129|899470|RXNORM|PLUM ALLERGENIC EXTRACT|PRUNUS DOMESTICA ALLERGENIC EXTRACT
C0772241|T121|236913|RXNORM|LEVOMETHADONE|LEVOMETHADONE
C0048045|T121|14852|RXNORM|4-AMINOMETHYLBENZOIC ACID|AMINOMETHYLBENZOIC ACID
C0048044|T123|14851|RXNORM|VIGABATRIN|VIGABATRIN
C0172021|T121|61609|RXNORM|ARBUTAMINE|ARBUTAMINE
C0071098|T121|33739|RXNORM|PIPAMPERONE|PIPAMPERONE
C0071097|T121|33738|RXNORM|PIOGLITAZONE|PIOGLITAZONE
C0134235|T129|54214|RXNORM|OSPA PROTEIN|OSPA PROTEIN
C0053105|T121|18880|RXNORM|BENFLUOREX|BENFLUOREX
C3535675|T121|1368530|RXNORM|PANAX GINSENG WHOLE EXTRACT|PANAX GINSENG WHOLE EXTRACT
C0061720|T116|1368533|RXNORM|PREZATIDE|GLY-HIS-LYS-OH
C2346854|T197|1485046|RXNORM|ARSENIC CATION|ARSENIC CATION (3+)
C3535672|T121|1368534|RXNORM|SNAIL PREPARATION|SNAIL PREPARATION
C0077081|T121|38617|RXNORM|TRIDIHEXETHYL|TRIDIHEXETHYL
C0077073|T121|38610|RXNORM|TRICLOFOS|TRICLOFOS
C3535902|T121|1370578|RXNORM|STEARALKONIUM|STEARALKONIUM
C3486822|T121|1310134|RXNORM|ELYMUS REPENS ROOT EXTRACT|ELYMUS REPENS ROOT EXTRACT
C2080567|T121|817405|RXNORM|ASPIRIN / PHENYLPROPANOLAMINE|ASPIRIN / PHENYLPROPANOLAMINE
C1632844|T121|608343|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL|CALCIUM CARBONATE / CHOLECALCIFEROL
C1321598|T121|1044977|RXNORM|PANTHENOL|PANTHENOL
C2194257|T121|817400|RXNORM|ESTROGENS / TESTOSTERONE|ESTROGENS / TESTOSTERONE
C0027270|T123|1044975|RXNORM|NICOTINAMIDE ADENINE DINUCLEOTIDE (NAD)|NICOTINAMIDE ADENINE DINUCLEOTIDE (NAD)
C3264704|T121|1358846|RXNORM|ALARIA ESCULENTA EXTRACT|ALARIA ESCULENTA EXTRACT
C0633963|T121|1358844|RXNORM|1-PROPOXY-2-PROPANOL|1-PROPOXY-2-PROPANOL
C0054631|T121|1358845|RXNORM|2-MERCAPTOBENZOTHIAZOLE|2-MERCAPTOBENZOTHIAZOLE
C0772397|T121|237060|RXNORM|TORMENTIL|TORMENTIL
C0772399|T129|237062|RXNORM|HEPATITIS A IMMUNE GLOBULIN,HU|HEPATITIS A IMMUNE GLOBULIN,HU
C0073983|T121|36108|RXNORM|SALSALATE|SALSALATE
C2747686|T129|966943|RXNORM|PENICILLIUM CAMEMBERTI ALLERGENIC EXTRACT|PENICILLIUM CAMEMBERTI ALLERGENIC EXTRACT
C0073969|T121|36100|RXNORM|SALICIN|SALICIN
C3535901|T121|1370579|RXNORM|BEHENTRIMONIUM|BEHENTRIMONIUM
C1869488|T123|1435864|RXNORM|METHYLINOSITOL|METHYLINOSITOL
C3666150|T121|1435865|RXNORM|PEG-20 GLYCERYL ISOSTEARATE|PEG-20 GLYCERYL ISOSTEARATE
C3666151|T121|1435866|RXNORM|POLYGONATUM MULTIFLORUM WHOLE EXTRACT|POLYGONATUM MULTIFLORUM WHOLE EXTRACT
C3666152|T121|1435867|RXNORM|RHEUM OFFICINALE WHOLE EXTRACT|RHEUM OFFICINALE WHOLE EXTRACT
C0065520|T197|1435860|RXNORM|MAGNESIUM FLUORIDE|MAGNESIUM FLUORIDE
C3666148|T121|1435861|RXNORM|ANGELICA ATROPURPUREA ROOT EXTRACT|ANGELICA ATROPURPUREA ROOT EXTRACT
C3666149|T121|1435862|RXNORM|JUGLANS REGIA WHOLE EXTRACT|JUGLANS REGIA WHOLE EXTRACT
C2702356|T129|892517|RXNORM|CANTALOUPE ALLERGENIC EXTRACT|CUCUMIS MELO ALLERGENIC EXTRACT
C0004475|T121|1251|RXNORM|AZACITIDINE|AZACITIDINE
C3666153|T121|1435868|RXNORM|SAURURUS CHINENSIS WHOLE EXTRACT|SAURURUS CHINENSIS WHOLE EXTRACT
C3666154|T121|1435869|RXNORM|BABESIA MICROTI PREPARATION|BABESIA MICROTI PREPARATION
C0301503|T129|89886|RXNORM|RABIES IMMUNE GLOBULIN, HUMAN|RABIES IMMUNE GLOBULIN, HUMAN
C3153044|T121|1098500|RXNORM|HOG HAIR EXTRACT / HOG SKIN EXTRACT|HOG HAIR EXTRACT / HOG SKIN EXTRACT
C3538156|T121|1372272|RXNORM|GREEN PEPPERCORN EXTRACT|GREEN PEPPERCORN EXTRACT
C2928090|T121|1007168|RXNORM|BORAGE EXTRACT / RED CLOVER PREPARATION / SALICIN EXTRACT|BORAGE EXTRACT / RED CLOVER PREPARATION / SALICIN EXTRACT
C2928091|T121|1007169|RXNORM|CALCIUM CARBONATE / CHASTE TREE PREPARATION / MAGNESIUM OXIDE|CALCIUM CARBONATE / CHASTE TREE PREPARATION / MAGNESIUM OXIDE
C0700607|T129|203223|RXNORM|DIGOXIN ANTIBODIES FAB FRAGMENTS|DIGOXIN ANTIBODIES FAB FRAGMENTS
C0109669|T121|48064|RXNORM|CHROMOCARB DIETHYLAMINE|CHROMOCARB DIETHYLAMINE
C3834088|T122|1541726|RXNORM|CANANGA ODORATA FLOWER WAX|CANANGA ODORATA FLOWER WAX
C2928087|T121|1007165|RXNORM|FRUCTOOLIGOSACCHARIDE / LACTOBACILLUS / PECTIN|FRUCTOOLIGOSACCHARIDE / LACTOBACILLUS / PECTIN
C2928088|T121|1007166|RXNORM|CALCIUM CARBONATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CARBONATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C2928089|T121|1007167|RXNORM|METHAPYRILENE / PYRILAMINE|METHAPYRILENE / PYRILAMINE
C2928083|T121|1007161|RXNORM|BENZYDAMINE / DIPYRONE|BENZYDAMINE / DIPYRONE
C2928084|T121|1007162|RXNORM|ATROPINE / HYOSCYAMINE / PHENYLEPHRINE / PSEUDOEPHEDRINE / SCOPOLAMINE|ATROPINE / HYOSCYAMINE / PHENYLEPHRINE / PSEUDOEPHEDRINE / SCOPOLAMINE
C2928085|T121|1007163|RXNORM|NITRAZEPAM / OXAZEPAM / SCOPOLAMINE|NITRAZEPAM / OXAZEPAM / SCOPOLAMINE
C1874332|T121|689245|RXNORM|APROBARBITAL / BUTABARBITAL / PHENOBARBITAL|APROBARBITAL / BUTABARBITAL / PHENOBARBITAL
C0982060|T109|1309218|RXNORM|HYDROGENATED CASTOR OIL|HYDROGENATED CASTOR OIL
C1874319|T121|689241|RXNORM|ANTIPYRINE / HYDROCORTISONE / NEOMYCIN / POLYMYXIN B|ANTIPYRINE / HYDROCORTISONE / NEOMYCIN / POLYMYXIN B
C0038722|T121|10193|RXNORM|SULFATHIAZOLE|SULFATHIAZOLE
C0965390|T121|301739|RXNORM|ABARELIX|ABARELIX
C0376274|T109|1309211|RXNORM|CAJUPUT OIL|CAJUPUT OIL
C1802750|T168|1309210|RXNORM|OIL OF GARLIC|OIL OF GARLIC
C0070247|T109|1309213|RXNORM|PENNYROYAL OIL|PENNYROYAL OIL
C3254749|T109|1309212|RXNORM|GRAPEFRUIT OIL|GRAPEFRUIT OIL
C3255681|T121|1309215|RXNORM|HIBISCUS SABDARIFFA FLOWER EXTRACT|HIBISCUS SABDARIFFA FLOWER EXTRACT
C0439966|T109|1309214|RXNORM|CANANGA OIL|CANANGA OIL
C0304100|T121|1309217|RXNORM|CEDAR LEAF OIL|CEDAR LEAF OIL
C1509464|T109|1309216|RXNORM|POLYOXYL 40 CASTOR OIL|PEG-40 CASTOR OIL
C3255979|T109|1305655|RXNORM|SWEET MARJORAM OIL|SWEET MARJORAM OIL
C2052852|T121|818530|RXNORM|DIMENHYDRINATE / NIACIN / PENTYLENETETRAZOLE|DIMENHYDRINATE / NIACIN / PENTYLENETETRAZOLE
C0767316|T121|1362584|RXNORM|1,2-HEXANEDIOL|1,2-HEXANEDIOL
C0064745|T109|1305654|RXNORM|WEST INDIAN LEMONGRASS OIL|WEST INDIAN LEMONGRASS OIL
C3497625|T121|1310294|RXNORM|BOS TAURUS SPINAL CORD PREPARATION|BOVINE SPINAL CORD PREPARATION
C3848613|T116|1544275|RXNORM|ETHYL GLUTAMATE|ETHYL GLUTAMATE
C2928230|T121|1007308|RXNORM|BORAGE OIL / GAMMA LINOLEIC ACID|BORAGE OIL / GAMMA LINOLEIC ACID
C2928231|T121|1007309|RXNORM|CHOLINE / GLYCERIN|CHOLINE / GLYCERIN
C0206232|T121|67031|RXNORM|NADROPARIN|NADROPARIN
C2928222|T121|1007300|RXNORM|ALLANTOIN / BENZOCAINE / DIMETHICONE / PETROLATUM|ALLANTOIN / BENZOCAINE / DIMETHICONE / PETROLATUM
C2928223|T121|1007301|RXNORM|GUAIACOLSULFONATE / ZIPEPROL|GUAIACOLSULFONATE / ZIPEPROL
C2928224|T121|1007302|RXNORM|GUAIFENESIN / PHENOBARBITAL / THEOPHYLLINE|GUAIFENESIN / PHENOBARBITAL / THEOPHYLLINE
C2928225|T121|1007303|RXNORM|PHENYLTOLOXAMINE / PHOLCODINE|PHENYLTOLOXAMINE / PHOLCODINE
C2928226|T121|1007304|RXNORM|FENNEL SEED PREPARATION / SENNA LEAVES / SENNOSIDES, USP|FENNEL SEED PREPARATION / SENNA LEAVES / SENNOSIDES, USP
C2928229|T121|1007307|RXNORM|BUTHIAZIDE / DIHYDRALAZINE / METIPRANOLOL|BUTHIAZIDE / DIHYDRALAZINE / METIPRANOLOL
C3487974|T121|1314257|RXNORM|JUNIPERUS VIRGINIANA TWIG EXTRACT|JUNIPERUS VIRGINIANA TWIG EXTRACT
C3486689|T121|1314256|RXNORM|HERRING SPERM DNA|HERRING SPERM DNA
C3473142|T121|1298205|RXNORM|APPLE CIDER VINEGAR / CALCIUM CARBONATE|APPLE CIDER VINEGAR / CALCIUM CARBONATE
C0058261|T121|1311550|RXNORM|DISTEARYLDIMONIUM|DISTEARYLDIMONIUM
C3474040|T121|1311557|RXNORM|BENINCASA HISPIDA FRUIT EXTRACT|BENINCASA HISPIDA FRUIT EXTRACT
C3255603|T121|1311556|RXNORM|NONOXYNOL-10|NONOXYNOL-10
C0068787|T121|1311555|RXNORM|NITARSONE|NITARSONE
C0035780|T121|1311554|RXNORM|ROBENIDINE|ROBENIDINE
C1445797|T121|466563|RXNORM|POLYETHYLENE GLYCOLS / PROPYLENE GLYCOL|POLYETHYLENE GLYCOLS / PROPYLENE GLYCOL
C3255606|T121|1311559|RXNORM|NONOXYNOL-30|NONOXYNOL-30
C3255604|T109|1311558|RXNORM|NONOXYNOL-100|NONOXYNOL-100
C2728184|T130|1011426|RXNORM|PAPAYA ALLERGENIC EXTRACT|CARICA PAPAYA ALLERGENIC EXTRACT
C3486771|T121|1326503|RXNORM|POA PRATENSIS TOP EXTRACT|POA PRATENSIS TOP EXTRACT
C3282675|T121|1314259|RXNORM|1-TETRACOSANOL|1-TETRACOSANOL
C3265711|T121|1314258|RXNORM|(2-CARBETHOXYETHYL)DIETHOXY(METHYL)SILANE|(2-CARBETHOXYETHYL)DIETHOXY(METHYL)SILANE
C0030966|T130|8040|RXNORM|PEPTONES|PEPTONES
C0032478|T121|8514|RXNORM|POLYETHYLENE GLYCOL 400|POLYETHYLENE GLYCOL 400
C0032478|T121|8514|RXNORM|POLYETHYLENE GLYCOL 400|POLYETHYLENE GLYCOL 400
C2348479|T121|1337279|RXNORM|EVERLASTING EXTRACT|EVERLASTING EXTRACT
C0032477|T121|8513|RXNORM|POLYETHYLENE GLYCOL 300|POLYETHYLENE GLYCOL 300
C0031007|T121|8047|RXNORM|PERGOLIDE|PERGOLIDE
C3709647|T122|1487927|RXNORM|BETA-SITOSTERYL SULFATE|BETA-SITOSTERYL SULFATE
C0873181|T121|259511|RXNORM|BLACK COHOSH ROOT EXTRACT|BLACK COHOSH ROOT EXTRACT
C0873183|T121|259513|RXNORM|ECHINACEA PURPUREA ROOT EXTRACT|ECHINACEA PURPUREA ROOT EXTRACT
C0053950|T121|1370421|RXNORM|BOROGLUCONATE|BOROGLUCONATE
C0171473|T121|1091919|RXNORM|ROMIFIDINE|ROMIFIDINE
C0050402|T121|16688|RXNORM|ACECARBROMAL|ACECARBROMAL
C3819177|T121|1494183|RXNORM|ALPHA-D-GALACTOSIDASE ENZYME / LACTASE|ALPHA-D-GALACTOSIDASE ENZYME / LACTASE
C2722024|T129|975119|RXNORM|TURKEY ALLERGENIC EXTRACT|MELEAGRIS GALLOPAVO ALLERGENIC EXTRACT
C3500184|T121|1313956|RXNORM|CHROMIUM PICOLINATE / CINNAMON BARK|CHROMIUM PICOLINATE / CINNAMON BARK
C0359156|T129|107044|RXNORM|RABBIT ANTI-HUMAN T-LYMPHOCYTE GLOBULIN|RABBIT ANTI-HUMAN T-LYMPHOCYTE GLOBULIN
C2144535|T121|814985|RXNORM|IBUPROFEN / TOLPERISONE|IBUPROFEN / TOLPERISONE
C0058031|T121|23066|RXNORM|DIHEMATOPORPHYRIN ETHER|DIHEMATOPORPHYRIN ETHER
C2183733|T121|815052|RXNORM|ASPIRIN / DIPHENHYDRAMINE / PHENYLPROPANOLAMINE|ASPIRIN / DIPHENHYDRAMINE / PHENYLPROPANOLAMINE
C3833354|T109|1541235|RXNORM|BIOSACCHARIDE GUM-2|BIOSACCHARIDE GUM-2
C0966107|T121|302285|RXNORM|CONIVAPTAN|CONIVAPTAN
C0059483|T121|24285|RXNORM|EPSIPRANTEL|EPSIPRANTEL
C3153926|T121|1100466|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / BETA CAROTENE / CALCIUM CARBONATE / CHOLECALCIFEROL / CUPRIC OXIDE / FERROUS BISGLYCINATE / FOLIC ACID / IRON PROTEIN SUCCINYLATE / MAGNESIUM OXIDE / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC OXIDE|ALPHA TOCOPHEROL / ASCORBIC ACID / BETA CAROTENE / CALCIUM CARBONATE / CHOLECALCIFEROL / CUPRIC OXIDE / FERROUS BISGLYCINATE / FOLIC ACID / IRON PROTEIN SUCCINYLATE / MAGNESIUM OXIDE / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC OXIDE
C0555881|T121|144377|RXNORM|ARNICA EXTRACT|ARNICA EXTRACT
C3813320|T121|1541237|RXNORM|EUPOLYPHAGA SINENSIS EXTRACT|EUPOLYPHAGA SINENSIS PREPARATION
C2928667|T121|1007752|RXNORM|COENZYME Q10 / THIOCTATE / VITAMIN E|COENZYME Q10 / THIOCTATE / VITAMIN E
C3499525|T121|1312394|RXNORM|HYDROXYPROPYL DISTARCH PHOSPHATE, HIGH AMYLOSE CORN|HYDROXYPROPYL DISTARCH PHOSPHATE, HIGH AMYLOSE CORN
C3499526|T121|1312395|RXNORM|POLYGLYCERYL-10 STEARATE|POLYGLYCERYL-10 STEARATE
C3499527|T121|1312396|RXNORM|PEG-9 DIMETHICONE|PEG-9 DIMETHICONE
C2980094|T121|1312397|RXNORM|REGORAFENIB|REGORAFENIB
C3254664|T121|1312390|RXNORM|METHYL METHACRYLATE-GLYCOL DIMETHACRYLATE CROSSPOLYMER|METHYL METHACRYLATE-GLYCOL DIMETHACRYLATE CROSSPOLYMER
C2928888|T121|1007975|RXNORM|CHLORPHENIRAMINE / GUAIFENESIN|CHLORPHENIRAMINE / GUAIFENESIN
C3499524|T121|1312392|RXNORM|GLYCERYL CAPRYLATE-CAPRATE|GLYCERYL CAPRYLATE-CAPRATE
C2928887|T121|1007974|RXNORM|HYDROCHLOROTHIAZIDE / VERAPAMIL|HYDROCHLOROTHIAZIDE / VERAPAMIL
C3833356|T196|1541238|RXNORM|FERROUS CATION|FERROUS CATION
C2928886|T121|1007973|RXNORM|ASCORBIC ACID / QUININE|ASCORBIC ACID / QUININE
C0141982|T121|56161|RXNORM|SENNOSIDE B|SENNOSIDE B
C3710068|T109|1489000|RXNORM|DAVANA OIL|DAVANA OIL
C2928885|T121|1007972|RXNORM|ALLANTOIN / BENZALKONIUM|ALLANTOIN / BENZALKONIUM
C2981098|T121|1094500|RXNORM|CHLOPHEDIANOL / PHENYLEPHRINE / TRIPROLIDINE|CHLOPHEDIANOL / PHENYLEPHRINE / TRIPROLIDINE
C0724724|T129|221182|RXNORM|YELLOW-FEVER VIRUS|YELLOW-FEVER VIRUS
C2928883|T121|1007970|RXNORM|CLONIDINE / HYDROCHLOROTHIAZIDE / TRIAMTERENE|CLONIDINE / HYDROCHLOROTHIAZIDE / TRIAMTERENE
C3535905|T109|1370571|RXNORM|LAUROAMPHOACETATE|LAUROAMPHOACETATE
C2194180|T121|813995|RXNORM|ALLOPURINOL / COLCHICINE|ALLOPURINOL / COLCHICINE
C2183095|T121|815631|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN / SODIUM CITRATE|DEXTROMETHORPHAN / GUAIFENESIN / SODIUM CITRATE
C0065180|T121|28889|RXNORM|LORATADINE|LORATADINE
C0050236|T121|1546449|RXNORM|ISOFLUPREDONE|ISOFLUPREDONE
C2724201|T129|892368|RXNORM|CARROT ALLERGENIC EXTRACT|DAUCUS CAROTA SATIVA ALLERGENIC EXTRACT
C0717492|T121|214298|RXNORM|BENZOCAINE / DEXTROMETHORPHAN|BENZOCAINE / DEXTROMETHORPHAN
C0717493|T121|214299|RXNORM|BENZOCAINE / DOCUSATE|BENZOCAINE / DOCUSATE
C2701681|T129|852605|RXNORM|KOELERS GRASS POLLEN EXTRACT|KOELERIA MACRANTHA POLLEN EXTRACT
C2930202|T121|814394|RXNORM|BETAMETHASONE ACETATE / BETAMETHASONE SODIUM PHOSPHATE|BETAMETHASONE ACETATE / BETAMETHASONE SODIUM PHOSPHATE
C2701677|T129|852601|RXNORM|ROCKY MOUNTAIN JUNIPER POLLEN EXTRACT|JUNIPERUS SCOPULORUM POLLEN EXTRACT
C0023591|T121|6379|RXNORM|LEVULINIC ACID|LEVULINIC ACID
C2194313|T121|818740|RXNORM|CAFFEINE / DIPHENHYDRAMINE / ERGOTAMINE|CAFFEINE / DIPHENHYDRAMINE / ERGOTAMINE
C1619838|T121|611854|RXNORM|CHLORDIAZEPOXIDE / CLIDINIUM|CHLORDIAZEPOXIDE / CLIDINIUM
C2701685|T129|852609|RXNORM|RED CEDAR POLLEN EXTRACT|JUNIPERUS VIRGINIANA POLLEN EXTRACT
C0717769|T121|214565|RXNORM|FEXOFENADINE / PSEUDOEPHEDRINE|FEXOFENADINE / PSEUDOEPHEDRINE
C0075783|T121|37546|RXNORM|TALINOLOL|TALINOLOL
C3665150|T121|1435387|RXNORM|CENTAUREA BENEDICTA FLOWERING TOP EXTRACT|CENTAUREA BENEDICTA FLOWERING TOP EXTRACT
C3252566|T197|1364533|RXNORM|PYROPHOSPHATE|PYROPHOSPHATE
C0061930|T121|26288|RXNORM|GUAIACOLSULFONIC ACID|GUAIACOLSULFONIC ACID
C0017440|T130|4778|RXNORM|GENTIAN VIOLET|GENTIAN VIOLET
C0017440|T130|4778|RXNORM|GENTIAN VIOLET|GENTIAN VIOLET
C0068955|T121|31958|RXNORM|THEODRENALINE|THEODRENALINE
C2928939|T121|1008028|RXNORM|GUAIACOLSULFONATE / PROMETHAZINE|GUAIACOLSULFONATE / PROMETHAZINE
C2928940|T121|1008029|RXNORM|ORMETOPRIM / SULFADIMETHOXINE|ORMETOPRIM / SULFADIMETHOXINE
C1870115|T121|720825|RXNORM|SILODOSIN|SILODOSIN
C3464500|T121|1292439|RXNORM|MEASLES VIRUS VACCINE LIVE, ENDERS' ATTENUATED EDMONSTON STRAIN / MUMPS VIRUS VACCINE LIVE, JERYL LYNN STRAIN / RUBELLA VIRUS VACCINE LIVE (WISTAR RA 27-3 STRAIN) / VARICELLA-ZOSTER VIRUS VACCINE LIVE (OKA-MERCK) STRAIN|MEASLES VIRUS VACCINE LIVE, ENDERS' ATTENUATED EDMONSTON STRAIN / MUMPS VIRUS VACCINE LIVE, JERYL LYNN STRAIN / RUBELLA VIRUS VACCINE LIVE (WISTAR RA 27-3 STRAIN) / VARICELLA-ZOSTER VIRUS VACCINE LIVE (OKA-MERCK) STRAIN
C2928935|T121|1008024|RXNORM|ASCORBIC ACID / BIOTIN / CALCIUM CARBONATE / CUPRIC OXIDE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM OXIDE / NIACINAMIDE / PANTOTHENIC ACID / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / BIOTIN / CALCIUM CARBONATE / CUPRIC OXIDE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM OXIDE / NIACINAMIDE / PANTOTHENIC ACID / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN E / ZINC OXIDE
C2928936|T121|1008025|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL / SOY PROTEIN ISOLATE|CALCIUM CARBONATE / CHOLECALCIFEROL / SOY PROTEIN ISOLATE
C2928937|T121|1008026|RXNORM|BENZYL ALCOHOL / ZINC ACETATE|BENZYL ALCOHOL / ZINC ACETATE
C2928938|T121|1008027|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIACOLSULFONATE / GUAIFENESIN / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIACOLSULFONATE / GUAIFENESIN / PSEUDOEPHEDRINE
C2928931|T121|1008020|RXNORM|BENZOCAINE / PECTIN|BENZOCAINE / PECTIN
C2928932|T121|1008021|RXNORM|ASCORBIC ACID / PECTIN / ZINC GLUCONATE|ASCORBIC ACID / PECTIN / ZINC GLUCONATE
C2928933|T121|1008022|RXNORM|BENZOCAINE / MENTHOL / METHYL SALICYLATE|BENZOCAINE / MENTHOL / METHYL SALICYLATE
C2928934|T121|1008023|RXNORM|ASCORBIC ACID / VITAMIN B 12 / ZINC GLUCONATE|ASCORBIC ACID / VITAMIN B 12 / ZINC GLUCONATE
C3541342|T197|1424174|RXNORM|RADIUM CHLORIDE RA-223|RADIUM CHLORIDE RA-223
C2709762|T129|854958|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 3 VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 3 VACCINE
C0123903|T121|51487|RXNORM|IPRIFLAVONE|IPRIFLAVONE
C0123902|T121|51486|RXNORM|IPRAZOCHROME|IPRAZOCHROME
C0054120|T121|19759|RXNORM|BROMODIPHENHYDRAMINE|BROMAZINE
C3643347|T121|1424173|RXNORM|DIMETHICONE PEG-7 PHOSPHATE|DIMETHICONE PEG-7 PHOSPHATE
C2709754|T129|854950|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 2 VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 2 VACCINE
C0143559|T121|56701|RXNORM|STANNOUS TARTRATE|STANNOUS TARTRATE
C0010843|T123|1372540|RXNORM|CYTOSINE|CYTOSINE
C2709758|T129|854954|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 22F VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 22F VACCINE
C2709760|T129|854956|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 23F VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 23F VACCINE
C0051519|T197|17618|RXNORM|ALUMINUM PHOSPHATE|ALUMINIUM PHOSPHATE
C2701591|T129|852466|RXNORM|EPICOCCUM NIGRUM EXTRACT|EPICOCCUM NIGRUM EXTRACT
C0126777|T121|52358|RXNORM|MAGNESIUM GLUCONATE|MAGNESIUM GLUCONATE
C0126774|T121|52356|RXNORM|MAGNESIUM CITRATE|MAGNESIUM CITRATE
C2364539|T129|805539|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-URUGUAY -716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-URUGUAY -716-2007 (H3N2) (A-BRISBANE-10-2007-LIKE) STRAIN
C0051515|T197|17614|RXNORM|ALUMINUM MAGNESIUM SILICATE|ALMASILATE
C3256650|T109|1309459|RXNORM|SALIX ALBA LEAF EXTRACT|SALIX ALBA LEAF EXTRACT
C3256864|T121|1309458|RXNORM|PRUNUS ARMENIACA SEED EXTRACT|PRUNUS ARMENIACA SEED EXTRACT
C3256633|T109|1309457|RXNORM|POLYGONUM CUSPIDATUM ROOT EXTRACT|REYNOUTRIA JAPONICA ROOT EXTRACT
C2929800|T121|1008903|RXNORM|ASCORBIC ACID / VITAMIN A / VITAMIN D|ASCORBIC ACID / VITAMIN A / VITAMIN D
C3256436|T109|1309455|RXNORM|PLUM SEED OIL|PLUM SEED OIL
C3256434|T109|1309454|RXNORM|PLECTRANTHUS BARBATUS ROOT EXTRACT|PLECTRANTHUS BARBATUS ROOT EXTRACT
C3256433|T121|1309453|RXNORM|PLATYCLADUS ORIENTALIS LEAF EXTRACT|PLATYCLADUS ORIENTALIS LEAF EXTRACT
C3488654|T121|1309452|RXNORM|PIPER METHYSTICUM ROOT EXTRACT|MACROPIPER METHYSTICUM ROOT
C3256798|T109|1309451|RXNORM|OPUNTIA FICUS-INDICA STEM EXTRACT|OPUNTIA FICUS-INDICA STEM EXTRACT
C3256711|T109|1309450|RXNORM|OENOTHERA BIENNIS ROOT EXTRACT|OENOTHERA BIENNIS ROOT EXTRACT
C1701455|T121|641465|RXNORM|ARMODAFINIL|ARMODAFINIL
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, GRASS, BROME|PRASTERONE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, GRASS, JOHNSON|PRASTERONE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, GRASS, KENTUCKY BLUE|PRASTERONE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, GRASS, ORCHARD|PRASTERONE
C0028094|T121|7426|RXNORM|NIMODIPINE|NIMODIPINE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, RYE GRASS PERENNIAL|PRASTERONE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, GRASS, SWEET VERNAL|PRASTERONE
C0063103|T121|27220|RXNORM|HYDROQUINIDINE|HYDROQUINIDINE
C0063105|T197|27221|RXNORM|HYDROTALCITE|HYDROTALCITE
C3709597|T121|1487833|RXNORM|PRIMULA VERIS FLOWER EXTRACT|COWSLIP FLOWER EXTRACT
C2701737|T129|852687|RXNORM|MUCOR EXTRACT|MUCOR RACEMOSUS EXTRACT
C0055463|T121|20877|RXNORM|CHLOROXYLENOL|CHLOROXYLENOL
C0055463|T121|20877|RXNORM|CHLOROXYLENOL|CHLOROXYLENOL
C0055461|T121|20875|RXNORM|CHLOROXINE|CHLOROXINE
C0126177|T121|52177|RXNORM|LOTEPREDNOL ETABONATE|LOTEPREDNOL ETABONATE
C0126174|T121|52175|RXNORM|LOSARTAN|LOSARTAN
C3858058|T121|1550956|RXNORM|DIPHENHYDRAMINE / NAPROXEN|DIPHENHYDRAMINE / NAPROXEN
C3190827|T121|1145207|RXNORM|CHLORAMPHENICOL / DEOXYRIBONUCLEASES / PLASMIN|CHLORAMPHENICOL / DEOXYRIBONUCLEASES / PLASMIN
C0003524|T121|1029|RXNORM|CORYNEBACTERIUM PARVUM VACCINE|APAZONE
C2927818|T121|1006894|RXNORM|HYDROCHLOROTHIAZIDE / SOTALOL|HYDROCHLOROTHIAZIDE / SOTALOL
C2194099|T121|819833|RXNORM|METHENAMINE / SODIUM PHOSPHATE|METHENAMINE / SODIUM PHOSPHATE
C0178834|T121|618482|RXNORM|RICINOLEATE|RICINOLEATE
C0050409|T121|16695|RXNORM|ACEMETACIN|ACEMETACIN
C3474165|T121|1307870|RXNORM|PISTACHIO OIL|PISTACHIO OIL
C1302961|T121|392677|RXNORM|CYCLIZINE / DIPIPANONE|CYCLIZINE / DIPIPANONE
C0009325|T121|2714|RXNORM|COLLAGEN|COLLAGEN
C0220833|T121|70598|RXNORM|FUMARATE|FUMARATE
C0220836|T123|70599|RXNORM|GLUCONATE|GLUCONATE
C0078622|T121|39823|RXNORM|XIBORNOL|XIBORNOL
C0039418|T197|10349|RXNORM|SODIUM PERTECHNETATE TC 99M|SODIUM PERTECHNETATE TC 99M
C0027289|T123|7222|RXNORM|NADH|NADH
C0027302|T121|7226|RXNORM|NADOLOL|NADOLOL
C0040613|T121|10691|RXNORM|TRANEXAMIC ACID|TRANEXAMIC ACID
C2962827|T121|1087244|RXNORM|CALCIUM ASCORBATE / CALCIUM THREONATE / FERROUS ASPARTO GLYCINATE / FOLIC ACID / POLYSACCHARIDE IRON COMPLEX / SUCCINIC ACID / VITAMIN B 12|CALCIUM ASCORBATE / CALCIUM THREONATE / FERROUS ASPARTO GLYCINATE / FOLIC ACID / POLYSACCHARIDE IRON COMPLEX / SUCCINIC ACID / VITAMIN B 12
C2927893|T121|1006970|RXNORM|ACETAMINOPHEN / DIMENHYDRINATE|ACETAMINOPHEN / DIMENHYDRINATE
C2927894|T121|1006971|RXNORM|COUMARIN / RUTIN|COUMARIN / RUTIN
C2927895|T121|1006972|RXNORM|BISMUTH SUBGALLATE / BUTOXYCAINE / ZINC OXIDE|BISMUTH SUBGALLATE / BUTOXYCAINE / ZINC OXIDE
C2927896|T121|1006973|RXNORM|ATROPINE / EPINEPHRINE / TYRAMINE|ATROPINE / EPINEPHRINE / TYRAMINE
C2927897|T121|1006974|RXNORM|LIDOCAINE / LINDANE|LIDOCAINE / LINDANE
C2927898|T121|1006975|RXNORM|SULFAMERAZINE / TRIMETHOPRIM|SULFAMERAZINE / TRIMETHOPRIM
C2927899|T121|1006976|RXNORM|CELLULOSE / METHYLCELLULOSE|CELLULOSE / METHYLCELLULOSE
C2927900|T121|1006977|RXNORM|MEPROBAMATE / THEOPHYLLINE|MEPROBAMATE / THEOPHYLLINE
C2927901|T121|1006978|RXNORM|METHOCARBAMOL / METHYLNICOTINATE|METHOCARBAMOL / METHYLNICOTINATE
C2701782|T129|852756|RXNORM|PHOMA EXTRACT|PHOMA EXTRACT
C2929944|T121|1009049|RXNORM|FERROUS SULFATE / PHENOLPHTHALEIN|FERROUS SULFATE / PHENOLPHTHALEIN
C2929943|T121|1009048|RXNORM|CHLOROBUTANOL / PYROGALLOL|CHLOROBUTANOL / PYROGALLOL
C2725890|T129|972037|RXNORM|DUCK ALLERGENIC EXTRACT|DUCK ALLERGENIC EXTRACT
C3668757|T121|1441382|RXNORM|BACILLUS COAGULANS / INULIN|BACILLUS COAGULANS / INULIN
C0771472|T121|236219|RXNORM|ALIBENDOL|ALIBENDOL
C2346970|T121|1441386|RXNORM|BAZEDOXIFENE|BAZEDOXIFENE
C2723573|T129|867142|RXNORM|PRAIRIE SAGEBRUSH POLLEN EXTRACT|ARTEMISIA FRIGIDA POLLEN EXTRACT
C0036751|T123|1311214|RXNORM|SEROTONIN|SEROTONIN
C3848609|T109|1544483|RXNORM|BIS-PEG-10 DIMETHICONE DIMER DILINOLEATE COPOLYMER|BIS-PEG-10 DIMETHICONE DIMER DILINOLEATE COPOLYMER
C3485578|T121|1310091|RXNORM|SYZYGIUM CUMINI SEED EXTRACT|SYZYGIUM CUMINI SEED EXTRACT
C0218633|T121|70161|RXNORM|MOLGRAMOSTIM|RECOMBINANT HUMAN GM-CSF
C3485579|T121|1310093|RXNORM|HABERLEA RHODOPENSIS LEAF EXTRACT|HABERLEA RHODOPENSIS LEAF EXTRACT
C0040005|T123|10524|RXNORM|THREONINE|THREONINE
C0753678|T121|679314|RXNORM|PALIPERIDONE|PALIPERIDONE
C3255698|T121|1310094|RXNORM|LOPHATHERUM GRACILE LEAF EXTRACT|LOPHATHERUM GRACILE LEAF EXTRACT
C3255699|T109|1310097|RXNORM|LOVAGE OIL|LOVAGE OIL
C3486005|T109|1310096|RXNORM|RUBUS CHAMAEMORUS SEED OIL|RUBUS CHAMAEMORUS SEED OIL
C3486772|T121|1310099|RXNORM|PODOPHYLLUM PELTATUM ROOT EXTRACT|PODOPHYLLUM PELTATUM ROOT EXTRACT
C3486012|T121|1310098|RXNORM|KAEMPFERIA GALANGA ROOT EXTRACT|KAEMPFERIA GALANGA ROOT EXTRACT
C0040018|T126|10528|RXNORM|THROMBIN|THROMBIN
C2929951|T121|1009056|RXNORM|FENTANYL / ROPIVACAINE / SODIUM CHLORIDE|FENTANYL / ROPIVACAINE / SODIUM CHLORIDE
C3848606|T109|1544486|RXNORM|MYRETH-4|MYRETH-4
C2929952|T121|1009057|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL / INULIN|CALCIUM CARBONATE / CHOLECALCIFEROL / INULIN
C0033705|T121|8871|RXNORM|PROTHIONAMIDE|PROTHIONAMIDE
C0727538|T121|223779|RXNORM|POTASSIUM BITARTRATE|POTASSIUM HYDROGEN TARTRATE
C0048215|T121|14997|RXNORM|4-CRESYL ACETATE|4-CRESYL ACETATE
C0070585|T121|33303|RXNORM|PHENOTHRIN|PHENOTHRIN
C3464062|T121|1313189|RXNORM|VANILLYL BUTYL ETHER|4-(BUTOXYMETHYL)-2-METHOXYPHENOL
C2725883|T129|895538|RXNORM|WHITE-TAILED DEER HAIR EXTRACT|WHITE-TAILED DEER HAIR ALLERGENIC EXTRACT
C3486288|T109|1313229|RXNORM|CLADOSIPHON OKAMURANUS PREPARATION|CLADOSIPHON OKAMURANUS PREPARATION
C3666880|T121|1437910|RXNORM|HAEMOPHILUS INFLUENZAE TYPE B, CAPSULAR POLYSACCHARIDE INACTIVATED TETANUS TOXOID CONJUGATE VACCINE / MENINGOCOCCAL GROUP C POLYSACCHARIDE / MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP Y|HAEMOPHILUS INFLUENZAE TYPE B, CAPSULAR POLYSACCHARIDE INACTIVATED TETANUS TOXOID CONJUGATE VACCINE / MENINGOCOCCAL GROUP C POLYSACCHARIDE / MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP Y
C0075639|T168|37422|RXNORM|SUNFLOWER SEED OIL|SUNFLOWER OIL
C0541315|T121|141704|RXNORM|EVEROLIMUS|EVEROLIMUS
C3465211|T197|1313228|RXNORM|CALCIUM ALUMINOSILICATE|CALCIUM ALUMINOSILICATE
C0597265|T122|1370575|RXNORM|POLYACRYLATE|POLYACRYLATE
C2929953|T121|1009058|RXNORM|FOLIC ACID / HEME IRON POLYPEPTIDE / POLYSACCHARIDE IRON COMPLEX / VITAMIN B 12|FOLIC ACID / HEME IRON POLYPEPTIDE / POLYSACCHARIDE IRON COMPLEX / VITAMIN B 12
C0050407|T121|1426379|RXNORM|ACEGLUTAMIDE|ACEGLUTAMIDE
C2927869|T121|1006946|RXNORM|ALOE EXTRACT / CASCARA SAGRADA|ALOE EXTRACT / CASCARA SAGRADA
C2080525|T121|814648|RXNORM|CITRIC ACID / DEXTROMETHORPHAN / PHENYLEPHRINE / SODIUM CITRATE|CITRIC ACID / DEXTROMETHORPHAN / PHENYLEPHRINE / SODIUM CITRATE
C0062648|T121|26849|RXNORM|HEXAMIDINE|HEXAMIDINE
C3535906|T195|1370570|RXNORM|LAIDLOMYCIN PROPIONATE|LAIDLOMYCIN PROPIONATE
C3256061|T109|1363610|RXNORM|MELON EXTRACT|MELON EXTRACT
C3253516|T121|1427238|RXNORM|CETYLDIMETHYLETHYLAMMONIUM BROMIDE|MECETRONIUM BROMIDE
C1968272|T122|748794|RXNORM|INERT INGREDIENTS|INERT INGREDIENTS
C3535904|T121|1370572|RXNORM|3-HYDROXY-4-METHOXYBENZENESULFONATE|3-HYDROXY-4-METHOXYBENZENESULFONATE
C2928421|T121|1007499|RXNORM|CHLORPHENIRAMINE / GUAIFENESIN / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / GUAIFENESIN / PHENYLPROPANOLAMINE / PSEUDOEPHEDRINE
C3488589|T121|1426375|RXNORM|ECHINOCOCCUS GRANULOSUS PREPARATION|HYDATID WORM PREPARATION
C0524704|T109|1427233|RXNORM|QUINATE|QUINATE
C3473504|T121|1427230|RXNORM|N,N-BIS(2-HYDROXYETHYL)-P-PHENYLENEDIAMINE SULFATE|N,N-BIS(2-HYDROXYETHYL)-P-PHENYLENEDIAMINE SULFATE
C3535903|T121|1370573|RXNORM|BUTEDRONATE|BUTEDRONATE
C1137427|T126|338817|RXNORM|AGALSIDASE BETA|AGALSIDASE BETA
C3256488|T121|1426376|RXNORM|3-HEXENYL ACETATE, (3Z)-|3-HEXENYL ACETATE, CIS-
C3500350|T121|1314398|RXNORM|DEXPANTHENOL / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|DEXPANTHENOL / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C0520442|T121|132871|RXNORM|ACETYLDIGITOXIN|ACETYLDIGITOXIN
C0006050|T131|1712|RXNORM|BOTULINUM TOXIN TYPE A|BOTULINUM TOXIN TYPE A
C3486554|T121|1330087|RXNORM|HEDERA HELIX FLOWERING TWIG EXTRACT|HEDERA HELIX FLOWERING TWIG EXTRACT
C0019223|T121|5254|RXNORM|HEPTAMINOL|HEPTAMINOL
C0218499|T131|1251576|RXNORM|IMIDACLOPRID|IMIDACLOPRID
C3538174|T121|1372308|RXNORM|HUMAN MAMMARY GLAND PREPARATION|HUMAN MAMMARY GLAND PREPARATION
C3256091|T109|1305761|RXNORM|SAPOSHNIKOVIA DIVARICATA ROOT EXTRACT|SAPOSHNIKOVIA DIVARICATA ROOT EXTRACT
C3256606|T121|1305763|RXNORM|MILK FAT, COW|MILK FAT, COW
C3256142|T109|1305762|RXNORM|COLOCASIA ESCULENTA ROOT EXTRACT|COLOCASIA ESCULENTA ROOT EXTRACT
C3864840|T121|1596138|RXNORM|HYDROXYPROPYL CORN AMYLOPECTIN, PHOSPHATE CROSSLINKED (4000 MPA.S AT 5%)|HYDROXYPROPYL CORN AMYLOPECTIN, PHOSPHATE CROSSLINKED (4000 MPA.S AT 5%)
C3864839|T131|1596139|RXNORM|MONOSODIUM METHYLARSONATE|MONOSODIUM METHYLARSONATE
C3496936|T121|1371968|RXNORM|GLYCERYL BEHENATE-EICOSADIOATE|GLYCERYL BEHENATE-EICOSADIOATE
C3473975|T121|1313225|RXNORM|ARTEMISIA ABROTANUM WHOLE EXTRACT|ARTEMISIA ABROTANUM WHOLE EXTRACT
C3198869|T109|1313224|RXNORM|ALUMINUM CHLOROHYDREX PROPYLENE GLYCOL|ALUMINUM CHLOROHYDREX PROPYLENE GLYCOL
C3864965|T109|1596136|RXNORM|BEHENOYL HYDROXYPROLINE|BEHENOYL HYDROXYPROLINE
C3864841|T109|1596137|RXNORM|DEHYDROXANTHAN GUM|DEHYDROXANTHAN GUM
C3255614|T121|1312647|RXNORM|TRIBEHENIN PEG-20 ESTERS|TRIBEHENIN PEG-20 ESTERS
C3834077|T122|1541738|RXNORM|STEARETH-20 METHACRYLATE|STEARETH-20 METHACRYLATE
C3834076|T122|1541739|RXNORM|STEARETH-7|STEARETH-7
C3834080|T122|1541734|RXNORM|BIOSACCHARIDE GUM-4|BIOSACCHARIDE GUM-4
C3834079|T121|1541735|RXNORM|BLACK CATECHU EXTRACT|BLACK CATECHU EXTRACT
C3834044|T121|1541736|RXNORM|QUATERNIUM-82|QUATERNIUM-82
C3834078|T122|1541737|RXNORM|CAPRAMIDOPROPYL BETAINE|CAPRAMIDOPROPYL BETAINE
C3834084|T122|1541730|RXNORM|CINNAMOMUM CAMPHORA RESIN|CINNAMOMUM CAMPHORA RESIN
C3834083|T121|1541731|RXNORM|EUCALYPTUS GUM EXTRACT|EUCALYPTUS GUM EXTRACT
C3834082|T109|1541732|RXNORM|COIX LACRYMA-JOBI VAR. MA-YUEN SEED OIL|COIX LACRYMA-JOBI VAR. MA-YUEN SEED OIL
C3834081|T122|1541733|RXNORM|4-HYDROXY ACETOPHENONE|4-HYDROXY ACETOPHENONE
C0052429|T121|18343|RXNORM|ARTEMETHER|ARTEMETHER
C0042306|T196|11121|RXNORM|VANADIUM|VANADIUM
C0042313|T195|11124|RXNORM|VANCOMYCIN|VANCOMYCIN
C0052432|T121|18346|RXNORM|ARTESUNATE|ARTESUNATE
C0047506|T130|14448|RXNORM|3-IODOBENZYLGUANIDINE|3-IODOBENZYLGUANIDINE
C3848593|T121|1545680|RXNORM|CERVUS ELAPHUS WHOLE PREPARATION|CERVUS ELAPHUS WHOLE PREPARATION
C0070313|T121|33086|RXNORM|PENTIFYLLINE|PENTIFYLLINE
C3256251|T121|1307947|RXNORM|PHELLODENDRON AMURENSE BARK EXTRACT|PHELLODENDRON AMURENSE BARK EXTRACT
C3256471|T121|1307946|RXNORM|COLA NUT EXTRACT|COLA NUT EXTRACT
C3255632|T121|1307945|RXNORM|GENTIANA LUTEA ROOT EXTRACT|GENTIANA LUTEA ROOT EXTRACT
C0040845|T131|10753|RXNORM|TRETINOIN|TRETINOIN
C0040845|T131|10753|RXNORM|TRETINOIN|TRETINOIN
C3256189|T121|1307943|RXNORM|BETULA PUBESCENS BARK EXTRACT|BETULA PUBESCENS BARK EXTRACT
C3247664|T121|1192753|RXNORM|BERMUDA GRASS POLLEN EXTRACT / TIMOTHY GRASS POLLEN EXTRACT|BERMUDA GRASS POLLEN EXTRACT / TIMOTHY GRASS POLLEN EXTRACT
C3665069|T121|1435256|RXNORM|BENZOCAINE / CAMPHOR / PHENOL|BENZOCAINE / CAMPHOR / PHENOL
C3668868|T109|1484860|RXNORM|LARREA TRIDENTATA WHOLE EXTRACT|LARREA TRIDENTATA WHOLE EXTRACT
C0010620|T121|3013|RXNORM|CYPROHEPTADINE|CYPROHEPTADINE
C0895222|T109|1484865|RXNORM|NERAL|NERAL
C2348160|T121|1307949|RXNORM|SAXIFRAGA STOLONIFERA LEAF EXTRACT|SAXIFRAGA STOLONIFERA LEAF EXTRACT
C2346607|T109|1307948|RXNORM|JUNIPERUS VIRGINIANA OIL|JUNIPERUS VIRGINIANA OIL
C0020350|T125|5530|RXNORM|HYDROXYESTRONES|HYDROXYESTRONES
C1960121|T121|753346|RXNORM|SINECATECHINS|SINECATECHINS
C0649350|T121|183379|RXNORM|RIVASTIGMINE|RIVASTIGMINE
C3488451|T121|1334750|RXNORM|VERBASCUM THAPSUS EXTRACT|VERBASCUM THAPSUS EXTRACT
C0033294|T121|8723|RXNORM|PROFLAVINE|PROFLAVINE
C0033308|T125|8727|RXNORM|PROGESTERONE|PROGESTERONE
C3859424|T121|1592895|RXNORM|DILAURYL CITRATE|DILAURYL CITRATE
C3464466|T121|1292333|RXNORM|FOLIC ACID / INOSITOL|FOLIC ACID / INOSITOL
C0733609|T126|227410|RXNORM|SULTILAINS|SULTILAINS
C0015137|T121|4182|RXNORM|ETRETINATE|ETRETINATE
C0015153|T121|4186|RXNORM|EUGENOL|EUGENOL
C3651725|T121|1430131|RXNORM|PERFLUOROPOLYMETHYLISOPROPYL ETHER|PERFLUOROPOLYMETHYLISOPROPYL ETHER
C0020852|T129|5666|RXNORM|IMMUNOGLOBULIN G|IMMUNOGLOBULIN G
C0015502|T123|4254|RXNORM|FACTOR VII|FACTOR VII
C0301352|T197|89767|RXNORM|COLLOID SULFUR|COLLOID SULFUR
C0937931|T121|581398|RXNORM|CITRUS PECTIN|CITRUS PECTIN
C3486743|T121|1350212|RXNORM|STAR ANISE EXTRACT|ILLICIUM VERUM SEED EXTRACT
C3486733|T121|1350211|RXNORM|PHLEUM PRATENSE TOP EXTRACT|PHLEUM PRATENSE TOP EXTRACT
C3486400|T121|1350210|RXNORM|TRIPE PREPARATION|TRIPE PREPARATION
C3486818|T168|1350214|RXNORM|SEMECARPUS ANACARDIUM JUICE EXTRACT|SEMECARPUS ANACARDIUM JUICE
C3645208|T109|1426943|RXNORM|DIBUTYLDITHIOCARBAMATE|DIBUTYLDITHIOCARBAMATE
C0035609|T195|9385|RXNORM|RIFAMYCINS|RIFAMYCINS
C0065988|T197|1426941|RXNORM|MERCURIC IODIDE|MERCURIC IODIDE
C3153835|T121|1100257|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / CALCIUM CITRATE / CHOLECALCIFEROL / CUPRIC OXIDE / DOCUSATE / FOLIC ACID / IRON CARBONYL / NIACINAMIDE / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / ZINC OXIDE|ALPHA TOCOPHEROL / ASCORBIC ACID / CALCIUM CITRATE / CHOLECALCIFEROL / CUPRIC OXIDE / DOCUSATE / FOLIC ACID / IRON CARBONYL / NIACINAMIDE / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / ZINC OXIDE
C3265816|T122|1426947|RXNORM|PEG-PPG-30-160 COPOLYMER|PEG-PPG-30-160 COPOLYMER
C3282583|T122|1426946|RXNORM|PPG-11 STEARYL ETHER|PPG-11 STEARYL ETHER
C3282690|T121|1426945|RXNORM|PPG-15 STEARYL ETHER BENZOATE|PPG-15 STEARYL ETHER BENZOATE
C3267653|T121|1426944|RXNORM|GLYCERETH-18 ETHYLHEXANOATE|GLYCERETH-18 ETHYLHEXANOATE
C3818787|T122|1491738|RXNORM|TOXICODENDRON SUCCEDANEUM WHOLE EXTRACT|TOXICODENDRON SUCCEDANEUM WHOLE EXTRACT
C3256406|T109|1424658|RXNORM|1,2-DIPALMITOYL-SN-GLYCERO-3-(PHOSPHO-RAC-(1-GLYCEROL))|1,2-DIPALMITOYL-SN-GLYCERO-3-(PHOSPHO-RAC-(1-GLYCEROL))
C0717712|T121|668797|RXNORM|DIPHENHYDRAMINE / MAGNESIUM SALICYLATE|DIPHENHYDRAMINE / MAGNESIUM SALICYLATE
C0795604|T125|253166|RXNORM|SYNTHETIC CONJUGATED ESTROGENS, A|SYNTHETIC CONJUGATED ESTROGENS, A
C0795600|T121|253165|RXNORM|DIDESMETHYLTOCOTRIENOL|DIDESMETHYLTOCOTRIENOL
C2740668|T129|899490|RXNORM|BLACK-EYED PEA ALLERGENIC EXTRACT|BLACK-EYED PEA ALLERGENIC EXTRACT
C0795598|T197|253163|RXNORM|DICALCIUM PHOSPHATE|DICALCIUM PHOSPHATE
C0795595|T121|253161|RXNORM|COLLAGEN HEMOSTAT|COLLAGEN HEMOSTAT
C3645163|T131|1426779|RXNORM|PHENYLMERCURY|PHENYLMERCURY
C0106127|T121|47070|RXNORM|BETA SITOSTEROL|BETA SITOSTEROL
C0877778|T121|262263|RXNORM|SKULLCAP PREPARATION|SKULLCAP PREPARATION
C0795610|T121|253168|RXNORM|GARCINIA CAMBOGIA PREPARATION|GARCINIA CAMBOGIA PREPARATION
C0044955|T121|12473|RXNORM|PREDNYLIDENE|PREDNYLIDENE
C2928371|T121|1007449|RXNORM|CETYLPYRIDINIUM / DIPHENHYDRAMINE|CETYLPYRIDINIUM / DIPHENHYDRAMINE
C2928370|T121|1007448|RXNORM|LIDOCAINE / NITROMERSOL|LIDOCAINE / NITROMERSOL
C0023764|T126|6406|RXNORM|LIPASE|LIPASE
C0023754|T168|6404|RXNORM|LINSEED OIL|LINSEED
C3818749|T109|1494198|RXNORM|1,3,3,3-TETRAFLUOROPROPENE, (1E)-|1,3,3,3-TETRAFLUOROPROPENE, (1E)-
C3152896|T129|1098274|RXNORM|SMOOTH SUMAC POLLEN EXTRACT|RHUS GLABRA POLLEN EXTRACT
C2928364|T121|1007442|RXNORM|CAPSICUM OLEORESIN / METHYLNICOTINATE|CAPSICUM OLEORESIN / METHYLNICOTINATE
C2928363|T121|1007441|RXNORM|CLOTRIMAZOLE / PHENYLETHYL ALCOHOL|CLOTRIMAZOLE / PHENYLETHYL ALCOHOL
C2928362|T121|1007440|RXNORM|DOBESILIC ACID / LIDOCAINE|DOBESILIC ACID / LIDOCAINE
C2928369|T121|1007447|RXNORM|FLUFENAMIC ACID / NIACIN / SULFATED MUCOPOLYSACCHARIDES|FLUFENAMIC ACID / NIACIN / SULFATED MUCOPOLYSACCHARIDES
C2928368|T121|1007446|RXNORM|AZINTAMIDE / SCOPOLAMINE|AZINTAMIDE / SCOPOLAMINE
C2928367|T121|1007445|RXNORM|ACETIC ACID / PYRETHRINS|ACETIC ACID / PYRETHRINS
C2928366|T121|1007444|RXNORM|ASPARTIC ACID / MAGNESIUM CHLORIDE|ASPARTIC ACID / MAGNESIUM CHLORIDE
C2193904|T121|819068|RXNORM|AMILORIDE / HYDROCHLOROTHIAZIDE / METHYLDOPA|AMILORIDE / HYDROCHLOROTHIAZIDE / METHYLDOPA
C0008241|T121|2382|RXNORM|PROGUANIL|PROGUANIL
C3192790|T121|1147841|RXNORM|CODEINE / PHENIRAMINE / PHENYLEPHRINE|CODEINE / PHENIRAMINE / PHENYLEPHRINE
C0754011|T121|1100072|RXNORM|ABIRATERONE|ABIRATERONE
C1169987|T121|352362|RXNORM|ACETAMINOPHEN / TRAMADOL|ACETAMINOPHEN / TRAMADOL
C1169990|T121|352365|RXNORM|CARBETAPENTANE / CHLORPHENIRAMINE|CARBETAPENTANE / CHLORPHENIRAMINE
C1169989|T121|352364|RXNORM|BUPRENORPHINE / NALOXONE|BUPRENORPHINE / NALOXONE
C1169992|T121|352367|RXNORM|CETIRIZINE / PSEUDOEPHEDRINE|CETIRIZINE / PSEUDOEPHEDRINE
C1169991|T121|352366|RXNORM|CARBINOXAMINE / METHSCOPOLAMINE / PSEUDOEPHEDRINE|CARBINOXAMINE / METHSCOPOLAMINE / PSEUDOEPHEDRINE
C0669388|T121|1424652|RXNORM|DECAN-4-OLIDE|DECAN-4-OLIDE
C0056852|T121|22051|RXNORM|CYPRODENATE|CYPRODENATE
C3504803|T121|1356680|RXNORM|CAMELLIA SINENSIS WHOLE EXTRACT|CAMELLIA SINENSIS WHOLE EXTRACT
C3504804|T121|1356686|RXNORM|HIPPOPHAE RHAMNOIDES WHOLE EXTRACT|HIPPOPHAE RHAMNOIDES WHOLE EXTRACT
C0909839|T121|276237|RXNORM|EMTRICITABINE|EMTRICITABINE
C0069717|T121|32592|RXNORM|OXALIPLATIN|OXALIPLATIN
C0142825|T121|56466|RXNORM|SODIUM CITRATE|SODIUM CITRATE
C0142825|T121|56466|RXNORM|SODIUM CITRATE|SODIUM CITRATE
C0142825|T121|56466|RXNORM|SODIUM CITRATE|SODIUM CITRATE
C3666307|T121|1436168|RXNORM|RHEUM PALMATUM ROOT EXTRACT|TURKEY RHUBARB ROOT EXTRACT
C2825688|T121|1313722|RXNORM|REGRELOR|REGRELOR
C3256255|T121|1313723|RXNORM|PHENOXYISOPROPANOL|PHENOXYISOPROPANOL
C3265176|T121|1313720|RXNORM|METHICONE (20 CST)|METHICONE (20 CST)
C3256628|T109|1313721|RXNORM|POLYGLYCERIN-6|POLYGLYCERIN-6
C3818750|T109|1494197|RXNORM|PEG-PPG-15-15 DIMETHICONE|PEG-PPG-15-15 DIMETHICONE
C1741338|T121|1313724|RXNORM|PHENYLETHYL RESORCINOL|PHENYLETHYL RESORCINOL
C1678805|T121|1492727|RXNORM|APREMILAST|APREMILAST
C0717800|T121|689460|RXNORM|GUAIFENESIN / HYDROMORPHONE|GUAIFENESIN / HYDROMORPHONE
C3255975|T109|1426619|RXNORM|PROPYLENE GLYCOL DICAPRYLATE|PROPYLENE GLYCOL DICAPRYLATE
C0005100|T121|1426|RXNORM|PROPYLENE GLYCOL MONOSTEARATE|BENZYL ALCOHOL
C1875600|T121|689467|RXNORM|OXYTETRACYCLINE / POLYMYXIN B|OXYTETRACYCLINE / POLYMYXIN B
C1875600|T121|689467|RXNORM|OXYTETRACYCLINE / POLYMYXIN B|OXYTETRACYCLINE / POLYMYXIN B
C1875600|T121|689467|RXNORM|OXYTETRACYCLINE / POLYMYXIN B|OXYTETRACYCLINE / POLYMYXIN B
C1875599|T121|689466|RXNORM|OXYTETRACYCLINE / PHENAZOPYRIDINE / SULFAMETHIZOLE|OXYTETRACYCLINE / PHENAZOPYRIDINE / SULFAMETHIZOLE
C0053526|T121|19257|RXNORM|BETHANECHOL|BETHANECHOL
C1302041|T121|392499|RXNORM|ASPIRIN / GLYCINE|ASPIRIN / GLYCINE
C0054306|T121|19928|RXNORM|BUTYLVINAL|BUTYLVINAL
C1302031|T121|392492|RXNORM|BENZTHIAZIDE / TRIAMTERENE|BENZTHIAZIDE / TRIAMTERENE
C1302034|T121|392494|RXNORM|ERYTHROMYCIN / ISOTRETINOIN|ERYTHROMYCIN / ISOTRETINOIN
C3255846|T121|1314594|RXNORM|LEMON PEEL EXTRACT|LEMON PEEL EXTRACT
C0717360|T129|214177|RXNORM|LYME DISEASE VACCINE|LYME DISEASE VACCINE
C1327841|T121|1426872|RXNORM|HEXYL 5-AMINOLEVULINATE|HEXYL 5-AMINOLEVULINATE
C0717363|T121|214179|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE|ACETAMINOPHEN / CHLORPHENIRAMINE
C0717361|T121|214178|RXNORM|ACETAMINOPHEN / BUTALBITAL|ACETAMINOPHEN / BUTALBITAL
C0073999|T121|36122|RXNORM|PHENYL SALICYLATE|PHENYL SALICYLATE
C2142855|T121|818689|RXNORM|CARBINOXAMINE / GUAIFENESIN / PSEUDOEPHEDRINE|CARBINOXAMINE / GUAIFENESIN / PSEUDOEPHEDRINE
C3255920|T109|1306152|RXNORM|CITRUS LIMON FRUIT OIL|CITRUS LIMON FRUIT OIL
C3255916|T109|1306151|RXNORM|CITRUS AURANTIUM FRUIT OIL|CITRUS AURANTIUM FRUIT OIL
C3255915|T109|1306150|RXNORM|CITRUS AURANTIUM FLOWER OIL|CITRUS AURANTIUM FLOWER OIL
C3256351|T109|1306157|RXNORM|CEDRUS ATLANTICA BARK OIL|CEDRUS ATLANTICA BARK OIL
C3256204|T109|1306156|RXNORM|BRAZIL NUT OIL|BRAZIL NUT OIL
C3256130|T109|1306155|RXNORM|BRASSICA RAPA VAR. RAPA OIL|BRASSICA RAPA VAR. RAPA OIL
C0143993|T121|56795|RXNORM|SUFENTANIL|SUFENTANIL
C3693106|T121|1482537|RXNORM|MALUS DOMESTICA WHOLE EXTRACT|MALUS DOMESTICA WHOLE EXTRACT
C0072982|T168|1306159|RXNORM|BRASSICA NAPUS OIL|BRASSICA NAPUS OIL
C3256492|T109|1306158|RXNORM|ABIES SIBIRICA LEAF OIL|ABIES SIBIRICA LEAF OIL
C2194085|T121|818685|RXNORM|DIAZEPAM / METOCLOPRAMIDE / SIMETHICONE|DIAZEPAM / METOCLOPRAMIDE / SIMETHICONE
C1527251|T121|498855|RXNORM|DOCUSATE / GLYCERIN|DOCUSATE / GLYCERIN
C1956796|T130|1426874|RXNORM|IOFLUPANE I-123|IODINE IOFLUPANE
C0771711|T121|236439|RXNORM|PANCREAS EXTRACT|PANCREAS EXTRACT
C3249289|T121|1235015|RXNORM|ALLANTOIN / COLLOIDAL OATMEAL|ALLANTOIN / COLLOIDAL OATMEAL
C3693107|T121|1482538|RXNORM|ACAI FRUIT PULP|ACAI FRUIT PULP
C2727018|T129|972480|RXNORM|RED CURRANT ALLERGENIC EXTRACT|RIBES RUBRUM ALLERGENIC EXTRACT
C0717405|T121|214217|RXNORM|AMINOPHYLLINE / AMOBARBITAL / EPHEDRINE|AMINOPHYLLINE / AMOBARBITAL / EPHEDRINE
C1738934|T121|1102129|RXNORM|BOCEPREVIR|BOCEPREVIR
C3848616|T109|1544272|RXNORM|ANEMARRHENA ASPHODELOIDES WHOLE EXTRACT|ANEMARRHENA ASPHODELOIDES WHOLE EXTRACT
C1874205|T121|690804|RXNORM|AMMONIUM CHLORIDE / CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE|AMMONIUM CHLORIDE / CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE
C3840273|T121|1544270|RXNORM|SYZYGIUM AROMATICUM FRUIT EXTRACT|SYZYGIUM AROMATICUM FRUIT EXTRACT
C3840272|T121|1544271|RXNORM|SWEET MARJORAM EXTRACT|SWEET MARJORAM EXTRACT
C3848612|T109|1544276|RXNORM|PROPYLENE GLYCOL 1-ALLYL ETHER|PROPYLENE GLYCOL 1-ALLYL ETHER
C0000956|T121|154|RXNORM|GELLAN GUM (HIGH ACYL)|ACENOCOUMAROL
C3848614|T116|1544274|RXNORM|HYDROLYZED SERICIN (ENZYMATIC; 2500 MW)|HYDROLYZED SERICIN (ENZYMATIC; 2500 MW)
C1874203|T121|690802|RXNORM|AMMONIUM CHLORIDE / ANTIMONY POTASSIUM TARTRATE / IPECAC|AMMONIUM CHLORIDE / ANTIMONY POTASSIUM TARTRATE / IPECAC
C1874614|T121|690808|RXNORM|BROMPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|BROMPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C1874614|T121|690808|RXNORM|BROMPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|BROMPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C0008736|T126|2525|RXNORM|CHYMOPAPAIN|CHYMOPAPAIN
C3542946|T121|1428420|RXNORM|JACOBAEA VULGARIS EXTRACT|JACOBAEA VULGARIS EXTRACT
C3818710|T121|1535493|RXNORM|LEPIDIUM SATIVUM SEED EXTRACT|LEPIDIUM SATIVUM SEED EXTRACT
C3256259|T109|1309502|RXNORM|ROSA GALLICA FLOWER EXTRACT|ROSA GALLICA FLOWER EXTRACT
C3665328|T109|1482539|RXNORM|PARSLEY OIL|PARSLEY OIL
C3254801|T121|1235449|RXNORM|ALUMINUM MAGNESIUM SILICATE / MAGNESIUM HYDROXIDE / SIMETHICONE|ALUMINUM MAGNESIUM SILICATE / MAGNESIUM HYDROXIDE / SIMETHICONE
C2006140|T121|817172|RXNORM|CALCIUM GLUCONATE / CALCIUM LACTOBIONATE|CALCIUM GLUCONATE / CALCIUM LACTOBIONATE
C2701814|T129|852814|RXNORM|ARIZONA CYPRESS POLLEN EXTRACT|CUPRESSUS ARIZONICA POLLEN EXTRACT
C0008183|T121|2354|RXNORM|THYROID STRONG|CHLORCYCLIZINE
C0770558|T125|235481|RXNORM|HUMAN CALCITONIN|HUMAN CALCITONIN
C2347832|T121|1343346|RXNORM|COMFREY ROOT EXTRACT|COMFREY ROOT EXTRACT
C0043597|T121|11469|RXNORM|MOFEZOLAC|MOFEZOLAC
C2927823|T121|1006899|RXNORM|GAMMA-LINOLENATE / VITAMIN E|GAMMA-LINOLENATE / VITAMIN E
C2927822|T121|1006898|RXNORM|CEREBRAL PHOSPHOLIPIDS / DOCOSAHEXAENOATE|CEREBRAL PHOSPHOLIPIDS / DOCOSAHEXAENOATE
C2927817|T121|1006893|RXNORM|ACETAMINOPHEN / CARBINOXAMINE / PHENYLPROPANOLAMINE|ACETAMINOPHEN / CARBINOXAMINE / PHENYLPROPANOLAMINE
C2927816|T121|1006892|RXNORM|BELLADONNA ALKALOIDS / KAOLIN / PHENOBARBITAL|BELLADONNA ALKALOIDS / KAOLIN / PHENOBARBITAL
C2927815|T121|1006891|RXNORM|CHLORPHENIRAMINE / HYDROCORTISONE / PYRILAMINE|CHLORPHENIRAMINE / HYDROCORTISONE / PYRILAMINE
C2927814|T121|1006890|RXNORM|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE / PSEUDOEPHEDRINE
C2927820|T121|1006896|RXNORM|BORAGE OIL / DOCOSAHEXAENOATE / EICOSAPENTAENOATE|BORAGE OIL / DOCOSAHEXAENOATE / EICOSAPENTAENOATE
C2927819|T121|1006895|RXNORM|FLUOCORTOLONE CAPROATE / FLUOCORTOLONE PIVALATE|FLUOCORTOLONE CAPROATE / FLUOCORTOLONE PIVALATE
C2937579|T121|1009451|RXNORM|COFFEE FRUIT PREPARATION|COFFEE FRUIT PREPARATION
C0077304|T121|38802|RXNORM|TRISULFAPYRIMIDINE|TRISULFAPYRIMIDINE
C0077013|T121|38555|RXNORM|TRIAZULENONE|LOPRAZOLAM
C0077015|T121|38557|RXNORM|TRIBENOSIDE|TRIBENOSIDE
C0041350|T129|1534774|RXNORM|TUFTSIN|TUFTSIN
C1996230|T121|834774|RXNORM|BROMPHENIRAMINE / DIPHENHYDRAMINE / PHENYLEPHRINE|BROMPHENIRAMINE / DIPHENHYDRAMINE / PHENYLEPHRINE
C0304116|T109|1309664|RXNORM|SASSAFRAS OIL|SASSAFRAS OIL
C0010372|T131|1309665|RXNORM|CROTON OIL|CROTON OIL
C0771571|T121|1309666|RXNORM|CINCHONA BARK EXTRACT|CINCHONA BARK EXTRACT
C3488586|T121|1309667|RXNORM|CINCHONA PUBESCENS BARK EXTRACT|CINCHONA PUBESCENS BARK EXTRACT
C0982323|T109|1363619|RXNORM|PEG-75 LANOLIN|PEG-75 LANOLIN
C3256078|T109|1363618|RXNORM|PEG-60 ALMOND GLYCERIDES|PEG-60 ALMOND GLYCERIDES
C0218640|T121|70167|RXNORM|LENOGRASTIM|LENOGRASTIM
C0982316|T109|1363615|RXNORM|PEG-40 SORBITAN DIISOSTEARATE|PEG-40 SORBITAN DIISOSTEARATE
C3256071|T109|1363614|RXNORM|PEG-4 LAURATE|PEG-4 LAURATE
C0982320|T109|1363617|RXNORM|PEG-6 LAURAMIDE|PEG-6 LAURAMIDE
C3256075|T109|1363616|RXNORM|PEG-5 OLEATE|PEG-5 OLEATE
C3256064|T121|1363611|RXNORM|PEG-15 GLYCERYL STEARATE|PEG-15 GLYCERYL STEARATE
C3488379|T121|1309669|RXNORM|EPHEDRA DISTACHYA FLOWERING TWIG EXTRACT|EPHEDRA DISTACHYA FLOWERING TWIG EXTRACT
C0982314|T121|1363613|RXNORM|PEG-4 DILAURATE|PEG-4 DILAURATE
C3256067|T121|1363612|RXNORM|PEG-20 STEARATE|PEG-20 STEARATE
C0040864|T121|10759|RXNORM|TRIAMCINOLONE|TRIAMCINOLONE
C0040864|T121|10759|RXNORM|TRIAMCINOLONE|TRIAMCINOLONE
C0040864|T121|10759|RXNORM|TRIAMCINOLONE|TRIAMCINOLONE
C0040864|T121|10759|RXNORM|TRIAMCINOLONE|TRIAMCINOLONE
C0040864|T121|10759|RXNORM|TRIAMCINOLONE|TRIAMCINOLONE
C0040864|T121|10759|RXNORM|TRIAMCINOLONE|TRIAMCINOLONE
C1874894|T121|689888|RXNORM|CODEINE / EPHEDRINE / GUAIFENESIN|CODEINE / EPHEDRINE / GUAIFENESIN
C3464489|T121|1331688|RXNORM|AGARUM CLATHRATUM EXTRACT|AGARUM CLATHRATUM EXTRACT
C0048897|T123|753340|RXNORM|SAPROPTERIN|SAPROPTERIN
C0048897|T123|753340|RXNORM|SAPROPTERIN|SAPROPTERIN
C1874889|T121|689881|RXNORM|COAL TAR / SALICYLIC ACID|COAL TAR / SALICYLIC ACID
C1874888|T121|689880|RXNORM|COAL TAR / POLYSORBATE 80|COAL TAR / POLYSORBATE 80
C0040853|T121|10756|RXNORM|TRIACETIN|TRIACETIN
C0040854|T130|10757|RXNORM|TRIACETONEAMINE-N-OXYL|TRIACETONEAMINE-N-OXYL
C3535889|T109|1370592|RXNORM|LAUROYL LACTYLATE|LAUROYL LACTYLATE
C0071069|T121|33712|RXNORM|PIMETHIXENE|PIMETHIXENE
C0885511|T121|1311289|RXNORM|LACTUCA VIROSA EXTRACT|WILD LETTUCE EXTRACT
C0071074|T121|33717|RXNORM|PINACIDIL|PINACIDIL
C0134337|T121|54236|RXNORM|OXATOMIDE|OXATOMIDE
C2714003|T109|1368889|RXNORM|TETRAFLUOROMETHANE|TETRAFLUOROMETHANE
C1739800|T109|1368888|RXNORM|THIOTAURINE|THIOTAURINE
C3666306|T121|1436167|RXNORM|PROPANEDIOL DICAPRYLATE|PROPANEDIOL DICAPRYLATE
C3281370|T121|1248730|RXNORM|ALFALFA PREPARATION / CHLOROPHYLL|ALFALFA PREPARATION / CHLOROPHYLL
C1875458|T121|705029|RXNORM|MAGNESIUM CHLORIDE / SODIUM CHLORIDE|MAGNESIUM CHLORIDE / SODIUM CHLORIDE
C0077190|T121|1368881|RXNORM|TRIMETHYLOLPROPANE|TRIMETHYLOLPROPANE
C0077140|T109|1368880|RXNORM|TRILAURIN|TRILAURIN
C0377344|T121|1368883|RXNORM|OLEYLAMIDE|OLEYLAMIDE
C0077214|T121|1368882|RXNORM|TRIMYRISTIN|TRIMYRISTIN
C0982210|T121|1368885|RXNORM|IMIDUREA|IMIDUREA
C0068051|T109|1368884|RXNORM|N-HYDROXYSUCCINIMIDE|N-HYDROXYSUCCINIMIDE
C0982352|T122|1368887|RXNORM|POLYSORBATE 85|POLYSORBATE 85
C0772483|T109|1368886|RXNORM|2-ETHYLHEXYL STEARATE|OCTYL STEARATE
C3486839|T121|1310150|RXNORM|PAPAVER RHOEAS FLOWER EXTRACT|PAPAVER RHOEAS FLOWER EXTRACT
C3487965|T121|1310151|RXNORM|SYMPHYTUM TUBEROSUM ROOT EXTRACT|SYMPHYTUM TUBEROSUM ROOT EXTRACT
C2981069|T121|1310152|RXNORM|DACTYLIS GLOMERATA TOP EXTRACT|DACTYLIS GLOMERATA TOP EXTRACT
C0085484|T007|1491010|RXNORM|ENTEROBACTER CLOACAE|ENTEROBACTER CLOACAE
C3486681|T121|1310154|RXNORM|SYZYGIUM JAMBOS SEED EXTRACT|SYZYGIUM JAMBOS SEED EXTRACT
C3487968|T121|1310155|RXNORM|ZANTHOXYLUM AMERICANUM BARK EXTRACT|ZANTHOXYLUM AMERICANUM BARK EXTRACT
C3487970|T121|1310157|RXNORM|JATEORHIZA CALUMBA ROOT EXTRACT|JATEORHIZA CALUMBA ROOT EXTRACT
C1097115|T109|1442718|RXNORM|1-NAPHTHALENESULFONIC ACID|1-NAPHTHALENESULFONIC ACID
C3487971|T121|1310159|RXNORM|JUGLANS REGIA FLOWERING TOP EXTRACT|JUGLANS REGIA FLOWERING TOP EXTRACT
C0023082|T195|1364397|RXNORM|LASALOCID|LASALOCID
C2698111|T121|1440972|RXNORM|ANAZOLENE ACID|ANAZOLENE ACID
C2194166|T121|820701|RXNORM|ACETAMINOPHEN / ASPIRIN / SALICYLAMIDE|ACETAMINOPHEN / ASPIRIN / SALICYLAMIDE
C0967817|T123|1440971|RXNORM|1-PALMITOYL-2-OLEOYL-SN-GLYCERO-3-(PHOSPHO-RAC-(1-GLYCEROL))|1-PALMITOYL-2-OLEOYL-SN-GLYCERO-3-(PHOSPHO-RAC-(1-GLYCEROL))
C3194702|T129|1116977|RXNORM|AMERICAN HOUSE DUST MITE EXTRACT|AMERICAN HOUSE DUST MITE EXTRACT
C0007332|T121|1440974|RXNORM|CASEINS|CASEINS
C3194704|T129|1116979|RXNORM|EUROPEAN HOUSE DUST MITE EXTRACT|EUROPEAN HOUSE DUST MITE EXTRACT
C2928068|T121|1007146|RXNORM|SHARK LIVER OIL / VITAMIN E|SHARK LIVER OIL / VITAMIN E
C2928069|T121|1007147|RXNORM|HOMATROPINE / PHENOBARBITAL|HOMATROPINE / PHENOBARBITAL
C2928067|T121|1007145|RXNORM|ECHINACEA ANGUSTIFOLIA EXTRACT / GOLDENSEAL EXTRACT|ECHINACEA ANGUSTIFOLIA EXTRACT / GOLDENSEAL EXTRACT
C2928064|T121|1007142|RXNORM|BENZALKONIUM / SALICYLIC ACID|BENZALKONIUM / SALICYLIC ACID
C2928065|T121|1007143|RXNORM|PERUVIAN BALSAM / TRYPSIN|PERUVIAN BALSAM / TRYPSIN
C2928062|T121|1007140|RXNORM|ESTROGENS, CONJUGATED (USP) / MEPROBAMATE|ESTROGENS, CONJUGATED (USP) / MEPROBAMATE
C2928063|T121|1007141|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / PSEUDOEPHEDRINE / PYRILAMINE|ACETAMINOPHEN / DEXTROMETHORPHAN / PSEUDOEPHEDRINE / PYRILAMINE
C2702418|T129|892575|RXNORM|PEACH ALLERGENIC EXTRACT|PRUNUS PERSICA ALLERGENIC EXTRACT
C2928070|T121|1007148|RXNORM|SALICYLIC ACID / TRIAMCINOLONE|SALICYLIC ACID / TRIAMCINOLONE
C2928071|T121|1007149|RXNORM|CHLORHEXIDINE / SIMETHICONE|CHLORHEXIDINE / SIMETHICONE
C3848544|T196|1546388|RXNORM|CEROUS CATION|CEROUS CATION
C0109398|T131|48008|RXNORM|CHLOROACETATE|CHLOROACETATE
C0016016|T126|4388|RXNORM|PLASMIN|PLASMIN
C0673093|T123|1546380|RXNORM|4-HYDROXYBUTYRIC ACID|4-HYDROXYBUTYRIC ACID
C3848547|T121|1546381|RXNORM|AMARANTH ACID|AMARANTH ACID
C3488985|T121|1309279|RXNORM|WITHANIA SOMNIFERA ROOT EXTRACT|WITHANIA SOMNIFERA ROOT EXTRACT
C0904505|T123|274403|RXNORM|MECASERMIN|MECASERMIN
C3848545|T121|1546386|RXNORM|BROMOTHEOPHYLLINE|BROMOTHEOPHYLLINE
C3535890|T121|1370591|RXNORM|METHYL AMINOMETHYLCYCLOHEXANE CARBOXAMIDE|METHYL AMINOMETHYLCYCLOHEXANE CARBOXAMIDE
C0002860|T125|784|RXNORM|ANDROSTENEDIONE|ANDROSTANEDIONE
C0061328|T121|25793|RXNORM|GLIQUIDONE|GLIQUIDONE
C0035668|T114|9394|RXNORM|RNA|RNA
C0035661|T121|9392|RXNORM|RITODRINE|RITODRINE
C0982076|T197|314553|RXNORM|CHLORIDE HEXAHYDRATE|CHLORIDE HEXAHYDRATE
C0795674|T121|253206|RXNORM|VALERIAN ROOT EXTRACT|VALERIAN ROOT EXTRACT
C0286738|T121|83395|RXNORM|SAQUINAVIR|SAQUINAVIR
C0043506|T196|1534771|RXNORM|ZIRCONIUM|ZIRCONIUM
C3833363|T121|1541249|RXNORM|POLIGNATE SODIUM|POLIGNATE SODIUM
C0883242|T121|265323|RXNORM|MYCOPHENOLATE|MYCOPHENOLATE
C3535886|T121|1370596|RXNORM|C14-16 OLEFIN SULFONATE|C14-16 OLEFIN SULFONATE
C3473135|T121|1298198|RXNORM|CHOLECALCIFEROL / FOLIC ACID / PYRIDOXINE / RIBOFLAVIN / VITAMIN B 12|CHOLECALCIFEROL / FOLIC ACID / PYRIDOXINE / RIBOFLAVIN / VITAMIN B 12
C2928244|T121|1007322|RXNORM|BENZOCAINE / CETYLPYRIDINIUM / MENTHOL / ZINC CHLORIDE|BENZOCAINE / CETYLPYRIDINIUM / MENTHOL / ZINC CHLORIDE
C0071751|T121|34296|RXNORM|POTASSIUM BICARBONATE|POTASSIUM BICARBONATE
C2928242|T121|1007320|RXNORM|ASCORBIC ACID / BIOTIN / FOLIC ACID / NIACIN / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|ASCORBIC ACID / BIOTIN / FOLIC ACID / NIACIN / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C2928243|T121|1007321|RXNORM|LOMBARD POPLAR POLLEN EXTRACT / WHITE POPLAR POLLEN EXTRACT|LOMBARD POPLAR POLLEN EXTRACT / WHITE POPLAR POLLEN EXTRACT
C2928248|T121|1007326|RXNORM|ASCORBIC ACID / FOLIC ACID / POLYSACCHARIDE IRON COMPLEX / VITAMIN B 12|ASCORBIC ACID / FOLIC ACID / POLYSACCHARIDE IRON COMPLEX / VITAMIN B 12
C2928249|T121|1007327|RXNORM|FOLIC ACID / IRON CARBONYL|FOLIC ACID / IRON CARBONYL
C2928766|T121|1007852|RXNORM|ALUMINUM CHLORHYDRATE / NEOMYCIN|ALUMINUM CHLOROHYDRATE / NEOMYCIN
C2928767|T121|1007853|RXNORM|CAFFEINE / SALICYLAMIDE / SALICYLIC ACID|CAFFEINE / SALICYLAMIDE / SALICYLIC ACID
C2928497|T121|1007577|RXNORM|CARBOXYMETHYLCELLULOSE / CASANTHRANOL|CARBOXYMETHYLCELLULOSE / CASANTHRANOL
C2928250|T121|1007328|RXNORM|BENZETHONIUM / MENTHOL|BENZETHONIUM / MENTHOL
C1172636|T195|1539239|RXNORM|DALBAVANCIN|DALBAVANCIN
C2928772|T121|1007858|RXNORM|CHLORHEXIDINE / SILVER SULFADIAZINE|CHLORHEXIDINE / SILVER SULFADIAZINE
C2928773|T121|1007859|RXNORM|MENTHOL / ZINC PYRITHIONE|MENTHOL / ZINC PYRITHIONE
C0071754|T197|34299|RXNORM|POTASSIUM BROMIDE|POTASSIUM BROMIDE
C0071753|T197|34298|RXNORM|POTASSIUM BROMATE|POTASSIUM BROMATE
C1012087|T004|1343912|RXNORM|CANDIDA TORRESII|CANDIDA TORRESII
C0078257|T121|39541|RXNORM|VINORELBINE|VINORELBINE
C0168706|T121|60906|RXNORM|TOCAMPHYL|TOCAMPHYL
C3535885|T121|1370597|RXNORM|MYRISTOYL SARCOSINATE|MYRISTOYL SARCOSINATE
C3464931|T121|1293412|RXNORM|5-HYDROXYTRYPTOPHAN / MAGNESIUM OXIDE / MELATONIN / TRYPTOPHAN / VITAMIN B6|5-HYDROXYTRYPTOPHAN / MAGNESIUM OXIDE / MELATONIN / TRYPTOPHAN / VITAMIN B6
C3651954|T121|1427391|RXNORM|DEXTROMETHORPHAN / PHENYLEPHRINE / THONZYLAMINE|DEXTROMETHORPHAN / PHENYLEPHRINE / THONZYLAMINE
C3505161|T121|1357998|RXNORM|AESCULUS GLABRA NUT EXTRACT|AESCULUS GLABRA NUT EXTRACT
C0067942|T121|1314271|RXNORM|N-DODECANE|N-DODECANE
C3497848|T109|1314270|RXNORM|LUFFA AEGYPTIACA SEED OIL|LUFFA AEGYPTIACA SEED OIL
C3465036|T121|1314273|RXNORM|N-ACETYL DIPEPTIDE-1|N-ACETYL DIPEPTIDE-1
C3474400|T121|1314272|RXNORM|ISOAMYL BUTYRATE|ISOAMYL BUTYRATE
C3489144|T121|1311579|RXNORM|TRIBULUS TERRESTRIS FRUIT EXTRACT|TRIBULUS TERRESTRIS FRUIT EXTRACT
C3282784|T121|1314274|RXNORM|STANNOUS 2-ETHYLHEXANOATE|STANNOUS 2-ETHYLHEXANOATE
C3255856|T121|1314277|RXNORM|PALMITOYL TETRAPEPTIDE-7|PALMITOYL TETRAPEPTIDE-7
C3256621|T109|1314276|RXNORM|ISOPENTYLDIOL|ISOPENTYLDIOL
C1509253|T109|1311575|RXNORM|C13-14 ISOPARAFFIN|C13-14 ISOPARAFFIN
C2954419|T121|1314278|RXNORM|SACCHARIDE ISOMERATE|SACCHARIDE ISOMERATE
C3474201|T121|1311577|RXNORM|CRATAEGUS MONOGYNA FRUIT EXTRACT|CRATAEGUS MONOGYNA FRUIT EXTRACT
C0173050|T121|1311576|RXNORM|COCAMIDOPROPYL BETAINE|COCAMIDOPROPYL BETAINE
C0624698|T121|1311571|RXNORM|ETHYL VANILLIN|ETHYL VANILLIN
C0939773|T121|285129|RXNORM|GLYBURIDE / METFORMIN|GLYBURIDE / METFORMIN
C3267737|T121|1311573|RXNORM|CITRUS AURANTIUM FRUIT EXTRACT|CITRUS AURANTIUM FRUIT EXTRACT
C1509204|T121|1311572|RXNORM|DECYL GLUCOSIDE|DECYL GLUCOSIDE
C0066531|T195|30005|RXNORM|MIDECAMYCIN|MIDECAMYCIN
C0359052|T121|106991|RXNORM|LIDOCAINE / METHYLPREDNISOLONE|LIDOCAINE / METHYLPREDNISOLONE
C0359051|T121|106990|RXNORM|CHLORQUINALDOL / HYDROCORTISONE|CHLORQUINALDOL / HYDROCORTISONE
C0066535|T121|30009|RXNORM|MIGLITOL|MIGLITOL
C0028215|T197|7486|RXNORM|NITROUS OXIDE|NITROUS OXIDE
C1874858|T121|689678|RXNORM|CITRIC ACID / MAGNESIUM OXIDE / SODIUM CARBONATE|CITRIC ACID / MAGNESIUM OXIDE / SODIUM CARBONATE
C0081580|T121|40660|RXNORM|AMYLOCAINE|AMYLOCAINE
C2726152|T129|971379|RXNORM|GREEN OLIVE ALLERGENIC EXTRACT|GREEN OLIVE ALLERGENIC EXTRACT
C0073096|T121|1000492|RXNORM|RESVERATROL|RESVERATROL
C2929381|T121|1008477|RXNORM|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E
C2929380|T121|1008476|RXNORM|METFORMIN / ROPINIROLE|METFORMIN / ROPINIROLE
C2929379|T121|1008475|RXNORM|FLUMETHASONE / TRIIODOTHYRONINE|FLUMETHASONE / LIOTHYRONINE
C2929378|T121|1008474|RXNORM|CLOTRIMAZOLE / HEXAMIDINE / PREDNISOLONE|CLOTRIMAZOLE / HEXAMIDINE / PREDNISOLONE
C2929377|T121|1008473|RXNORM|PHENYLEPHRINE / PRAMOXINE|PHENYLEPHRINE / PRAMOXINE
C2929376|T121|1008472|RXNORM|GINKGO BILOBA EXTRACT / KOREAN GINSENG ROOT EXTRACT|GINKGO BILOBA EXTRACT / KOREAN GINSENG ROOT EXTRACT
C2929375|T121|1008471|RXNORM|CALCIUM ASCORBATE / CALCIUM CARBONATE / CHOLECALCIFEROL / FOLIC ACID / PYRIDOXINE|CALCIUM ASCORBATE / CALCIUM CARBONATE / CHOLECALCIFEROL / FOLIC ACID / PYRIDOXINE
C2929374|T121|1008470|RXNORM|BENZALKONIUM / IDOXURIDINE / LIDOCAINE|BENZALKONIUM / IDOXURIDINE / LIDOCAINE
C2740793|T129|899734|RXNORM|CRANBERRY ALLERGENIC EXTRACT|VACCINIUM MACROCARPON ALLERGENIC EXTRACT
C0010192|T130|2890|RXNORM|COSYNTROPIN|COSYNTROPIN
C2929383|T121|1008479|RXNORM|AFRICAN PYGEUM EXTRACT / BEARBERRY PREPARATION / PUMPKIN SEED OIL / SAW PALMETTO EXTRACT|AFRICAN PYGEUM EXTRACT / BEARBERRY PREPARATION / PUMPKIN SEED OIL / SAW PALMETTO EXTRACT
C2929382|T121|1008478|RXNORM|DORNASE ALFA / STREPTOKINASE|DORNASE ALFA / STREPTOKINASE
C0064164|T123|28068|RXNORM|OXACEPROL|OXACEPROL
C0031404|T121|8129|RXNORM|PHENFORMIN|PHENFORMIN
C0717989|T121|214769|RXNORM|PHENYLEPHRINE / PROMETHAZINE|PHENYLEPHRINE / PROMETHAZINE
C0015824|T121|4327|RXNORM|FENDILINE|FENDILINE
C3153908|T121|1100448|RXNORM|PENTOBARBITAL / PHENYTOIN|PENTOBARBITAL / PHENYTOIN
C0717982|T121|214762|RXNORM|PHENIRAMINE / PHENYLTOLOXAMINE / PYRILAMINE|PHENIRAMINE / PHENYLTOLOXAMINE / PYRILAMINE
C3281555|T121|1249116|RXNORM|CALAMINE / MENTHOL / PETROLATUM / ZINC OXIDE|CALAMINE / MENTHOL / PETROLATUM / ZINC OXIDE
C0051607|T121|17698|RXNORM|AMINEPTIN|AMINEPTINE
C1874169|T121|692568|RXNORM|ALUMINUM HYDROXIDE / MAGNESIUM HYDROXIDE / MAGNESIUM TRISILICATE|ALUMINUM HYDROXIDE / MAGNESIUM HYDROXIDE / MAGNESIUM TRISILICATE
C3268167|T121|1248141|RXNORM|ASCORBIC ACID / BETA CAROTENE / CALCIUM CARBONATE / CHOLECALCIFEROL / CUPRIC OXIDE / DOCUSATE / FOLIC ACID / IRON CARBONYL / MAGNESIUM OXIDE / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / BETA CAROTENE / CALCIUM CARBONATE / CHOLECALCIFEROL / CUPRIC OXIDE / DOCUSATE / FOLIC ACID / IRON CARBONYL / MAGNESIUM OXIDE / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN E / ZINC OXIDE
C0062220|T126|26514|RXNORM|HEMICELLULASE|HEMICELLULASE
C2740848|T129|899883|RXNORM|PEAR ALLERGENIC EXTRACT|PYRUS COMMUNIS ALLERGENIC EXTRACT
C0994494|T121|317857|RXNORM|PARSLEY EXTRACT|PARSLEY EXTRACT
C3535884|T109|1370598|RXNORM|COCOYL SARCOSINATE|COCOYL SARCOSINATE
C0076625|T123|38233|RXNORM|THYMOSTIMULIN|THYMOSTIMULIN
C1445240|T121|1370790|RXNORM|ASTACUS ASTACUS EXTRACT|ASTACUS ASTACUS EXTRACT
C3709636|T121|1487909|RXNORM|EPERUA FALCATA BARK EXTRACT|EPERUA FALCATA BARK EXTRACT
C0961780|T121|1371313|RXNORM|ISOXAFLUTOLE|ISOXAFLUTOLE
C3537693|T121|1371312|RXNORM|GRIFOLA FRONDOSA WHOLE EXTRACT|GRIFOLA FRONDOSA WHOLE EXTRACT
C3537692|T122|1371311|RXNORM|GLYCERETH-7|GLYCERETH-7
C2711031|T121|859393|RXNORM|ADAPALENE / BENZOYL PEROXIDE|ADAPALENE / BENZOYL PEROXIDE
C0388762|T130|1371317|RXNORM|N,N-DIMETHYLACRYLAMIDE|N,N-DIMETHYLACRYLAMIDE
C3495101|T121|1370792|RXNORM|URTICA URENS EXTRACT|URTICA URENS EXTRACT
C3537694|T168|1371314|RXNORM|VANILLIN 2,3-BUTANEDIOL ACETAL, CIS-|VANILLIN 2,3-BUTANEDIOL ACETAL, CIS-
C2701725|T129|852669|RXNORM|WHITE MULBERRY POLLEN EXTRACT|MORUS ALBA POLLEN EXTRACT
C0717602|T121|214405|RXNORM|CHLORPHENIRAMINE / EPHEDRINE / GUAIFENESIN|CHLORPHENIRAMINE / EPHEDRINE / GUAIFENESIN
C3537696|T122|1371318|RXNORM|PPG-25-LAURETH-25|PPG-25-LAURETH-25
C3556198|T121|1374794|RXNORM|SILICON DIOXIDE / TRICALCIUM PHOSPHATE|SILICON DIOXIDE / TRICALCIUM PHOSPHATE
C2747605|T129|966696|RXNORM|ORANGE PEKOE TEA ALLERGENIC EXTRACT|CAMELLIA SINENSIS ALLERGENIC EXTRACT
C2928917|T121|1008006|RXNORM|ASPIRIN / CAFFEINE / MAGNESIUM SALICYLATE|ASPIRIN / CAFFEINE / MAGNESIUM SALICYLATE
C2928918|T121|1008007|RXNORM|DIMETHICONE / PRAMOXINE|DIMETHICONE / PRAMOXINE
C2928916|T121|1008004|RXNORM|CALCIUM CARBONATE / SOY PROTEIN ISOLATE|CALCIUM CARBONATE / SOY PROTEIN ISOLATE
C2736424|T121|1008005|RXNORM|LEUCINE / PHENYLALANINE|LEUCINE / PHENYLALANINE
C2928914|T121|1008002|RXNORM|BROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE|BROMPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN / PHENYLEPHRINE
C2928915|T121|1008003|RXNORM|BISMUTH ALUMINATE / DOCUSATE|BISMUTH ALUMINATE / DOCUSATE
C2928912|T121|1008000|RXNORM|AMMONIUM CHLORIDE / BENZOATE / CLOBUTINOL|AMMONIUM CHLORIDE / BENZOATE / CLOBUTINOL
C2928913|T121|1008001|RXNORM|GLUCOSE / MAGNESIUM ACETATE / POTASSIUM ACETATE / SODIUM CHLORIDE|GLUCOSE / MAGNESIUM ACETATE / POTASSIUM ACETATE / SODIUM CHLORIDE
C2928530|T121|1007612|RXNORM|CALCIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C2928530|T121|1007612|RXNORM|CALCIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C0017505|T125|4791|RXNORM|GESTONORONE CAPROATE|GESTONORONE CAPROATE
C2928919|T121|1008008|RXNORM|ALLANTOIN / DIMETHICONE|ALLANTOIN / DIMETHICONE
C2928920|T121|1008009|RXNORM|ASCORBIC ACID / IRON CARBONYL|ASCORBIC ACID / IRON CARBONYL
C3538339|T121|1372565|RXNORM|LAMINARIA DIGITATA HYDROLIZED ALGINIC ACID|LAMINARIA DIGITATA HYDROLIZED ALGINIC ACID
C1365533|T121|1372564|RXNORM|COLTSFOOT LEAF EXTRACT|TUSSILAGO FARFARA LEAF EXTRACT
C3538340|T122|1372567|RXNORM|POLYQUATERNIUM-37 (25000 MPA.S)|POLYQUATERNIUM-37 (25000 MPA.S)
C2709774|T129|854970|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 8 VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 8 VACCINE
C3538336|T121|1372561|RXNORM|PINUS SYLVESTRIS CONE EXTRACT|PINUS SYLVESTRIS CONE EXTRACT
C0021547|T127|5833|RXNORM|INOSITOL|INOSITOL
C0042878|T127|11258|RXNORM|VITAMIN K|VITAMIN K
C2709778|T129|854974|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 9V VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 9V VACCINE
C0042874|T127|11256|RXNORM|VITAMIN E|VITAMIN E
C0042874|T127|11256|RXNORM|VITAMIN E|VITAMIN E
C3537529|T109|1370986|RXNORM|DULACIA INOPIFLORA WOOD EXTRACT|DULACIA INOPIFLORA WOOD EXTRACT
C0042866|T127|11253|RXNORM|VITAMIN D|VITAMIN D
C0042849|T127|11251|RXNORM|VITAMIN B COMPLEX|VITAMIN B COMPLEX
C0140591|T121|55679|RXNORM|RILMENIDINE|RILMENIDINE
C0053245|T121|19008|RXNORM|BENZTHIAZIDE|BENZTHIAZIDE
C3651780|T121|1428422|RXNORM|POPULUS BALSAMIFERA LEAF BUD EXTRACT|POPULUS BALSAMIFERA LEAF BUD EXTRACT
C3651779|T121|1428423|RXNORM|SASSAFRA ALBIDUM ROOT BARK EXTRACT|SASSAFRA ALBIDUM ROOT BARK EXTRACT
C0452460|T168|1307149|RXNORM|TOMATO JUICE|TOMATO JUICE
C3255706|T109|1307148|RXNORM|NEOPENTYL GLYCOL DIETHYLHEXANOATE|NEOPENTYL GLYCOL DIETHYLHEXANOATE
C0140575|T195|55672|RXNORM|RIFABUTIN|RIFABUTIN
C3255663|T121|1307144|RXNORM|ELAEIS GUINEENSIS FRUIT BUTTER|ELAEIS GUINEENSIS FRUIT BUTTER
C2365142|T116|1307143|RXNORM|SILK AMINO ACIDS|SILK AMINO ACIDS
C0070108|T121|32926|RXNORM|PAREGORIC|PAREGORIC
C0385231|T121|1307141|RXNORM|DIBENZYLIDENE SORBITOL|DIBENZYLIDENE SORBITOL
C2928768|T121|1007854|RXNORM|CLOTRIMAZOLE / DEXAMETHASONE|CLOTRIMAZOLE / DEXAMETHASONE
C0873084|T121|259421|RXNORM|KAVA ROOT|KAVA ROOT
C0165590|T121|60207|RXNORM|DORZOLAMIDE|DORZOLAMIDE
C2928245|T121|1007323|RXNORM|BUTABARBITAL / METHAMPHETAMINE|BUTABARBITAL / METHAMPHETAMINE
C2928770|T121|1007856|RXNORM|NIFURZIDE / PECTIN|NIFURZIDE / PECTIN
C2348785|T109|1309479|RXNORM|THYMUS OIL|THYMUS OIL
C3255734|T109|1309478|RXNORM|HYDROGENATED COTTONSEED OIL|HYDROGENATED COTTONSEED OIL
C2928771|T121|1007857|RXNORM|FRAMYCETIN / GRAMICIDIN|FRAMYCETIN / GRAMICIDIN
C3488977|T121|1309471|RXNORM|SINAPSIS ARVENSIS FLOWERING-FRUITING TOP EXTRACT|SINAPSIS ARVENSIS FLOWERING-FRUITING TOP EXTRACT
C2928764|T121|1007850|RXNORM|PANCREATIN / PEPSIN A|PANCREATIN / PEPSIN A
C3256809|T109|1309473|RXNORM|SMILAX ARISTOLOCHIAEFOLIA ROOT EXTRACT|SMILAX ARISTOLOCHIAEFOLIA ROOT EXTRACT
C3255844|T121|1309472|RXNORM|HUMULUS LUPULUS STEM EXTRACT|HUMULUS LUPULUS STEM EXTRACT
C3488917|T121|1309475|RXNORM|HYDRANGEA ARBORESCENS ROOT EXTRACT|HYDRANGEA ARBORESCENS ROOT EXTRACT
C3256448|T109|1309474|RXNORM|TAGETES ERECTA FLOWER EXTRACT|TAGETES ERECTA FLOWER EXTRACT
C3254762|T109|1309477|RXNORM|TEA LEAF OIL|TEA LEAF OIL
C2928765|T121|1007851|RXNORM|BACITRACIN / LIDOCAINE|BACITRACIN / LIDOCAINE
C0051043|T121|17214|RXNORM|CAFEDRINE / THEODRENALINE|CAFEDRINE / THEODRENALINE
C2727872|T129|895195|RXNORM|EUROPEAN RABBIT SKIN EXTRACT|ORYCTOLAGUS CUNICULUS SKIN EXTRACT
C2344265|T129|798220|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 14 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 14 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C2726215|T129|968123|RXNORM|STACHYBOTRYS CHARTARUM ALLERGENIC EXTRACT|STACHYBOTRYS CHARTARUM ALLERGENIC EXTRACT
C2741285|T129|900754|RXNORM|RED PINE POLLEN EXTRACT|PINUS RESINOSA POLLEN EXTRACT
C3268305|T121|1248604|RXNORM|GIANT RAGWEED POLLEN EXTRACT / SHORT RAGWEED POLLEN EXTRACT|GIANT RAGWEED POLLEN EXTRACT / SHORT RAGWEED POLLEN EXTRACT
C2741282|T129|900750|RXNORM|AUSTRIAN PINE POLLEN EXTRACT|PINUS NIGRA POLLEN EXTRACT
C2746972|T109|968631|RXNORM|CHIA SEED OIL|CHIA SEED OIL
C0025815|T125|6902|RXNORM|METHYLPREDNISOLONE|METHYLPREDNISOLONE
C0025815|T125|6902|RXNORM|METHYLPREDNISOLONE|METHYLPREDNISOLONE
C0025815|T125|6902|RXNORM|METHYLPREDNISOLONE|METHYLPREDNISOLONE
C0717747|T121|214545|RXNORM|EPINEPHRINE / ETIDOCAINE|EPINEPHRINE / ETIDOCAINE
C0717750|T121|214547|RXNORM|EPINEPHRINE / PRILOCAINE|EPINEPHRINE / PRILOCAINE
C0063090|T197|27208|RXNORM|HYDROIODIC ACID|HYDROIODIC ACID
C0718037|T121|214813|RXNORM|RESERPINE / TRICHLORMETHIAZIDE|RESERPINE / TRICHLORMETHIAZIDE
C0717744|T121|214542|RXNORM|EPHEDRINE / PHENOBARBITAL / THEOPHYLLINE|EPHEDRINE / PHENOBARBITAL / THEOPHYLLINE
C0043408|T007|1432993|RXNORM|YERSINIA PESTIS|YERSINIA PESTIS
C0796392|T129|253337|RXNORM|BEVACIZUMAB|BEVACIZUMAB
C3485068|T121|1309783|RXNORM|EUPATORIUM PERFOLIATUM FLOWERING TOP EXTRACT|EUPATORIUM PERFOLIATUM FLOWERING TOP EXTRACT
C3488557|T121|1309782|RXNORM|COLLINSONIA CANADENSIS ROOT EXTRACT|COLLINSONIA CANADENSIS ROOT EXTRACT
C3488555|T121|1309781|RXNORM|SANICULA EUROPAEA LEAF EXTRACT|SANICULA EUROPAEA LEAF EXTRACT
C2928251|T121|1007329|RXNORM|IBUPROFEN / PHENYLEPHRINE|IBUPROFEN / PHENYLEPHRINE
C3853724|T121|1594581|RXNORM|PHELLODENDRON AMURENSE WHOLE EXTRACT|PHELLODENDRON AMURENSE WHOLE EXTRACT
C3152944|T121|1309786|RXNORM|PLATYCODON GRANDIFLORUM LEAF EXTRACT|PLATYCODON GRANDIFLORUM LEAF EXTRACT
C3487957|T121|1309785|RXNORM|GOSSYPIUM HERBACEUM ROOT BARK EXTRACT|GOSSYPIUM HERBACEUM ROOT BARK EXTRACT
C3860110|T121|1594582|RXNORM|SCOPOLIA CARNIOLICA WHOLE EXTRACT|SCOPOLIA CARNIOLICA WHOLE EXTRACT
C3488667|T121|1309789|RXNORM|ARUM MACULATUM ROOT EXTRACT|ARUM MACULATUM ROOT EXTRACT
C3160309|T121|1309788|RXNORM|EUCOMMIA ULMOIDES BARK EXTRACT|EUCOMMIA ULMOIDES BARK EXTRACT
C2344273|T129|798228|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 4 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 4 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C0057383|T121|22503|RXNORM|DENAVERINE|DENAVERINE
C2828213|T130|1546452|RXNORM|IOTHALAMIC ACID I-125|IOTHALAMIC ACID I-125
C0085251|T121|42368|RXNORM|ENCAINIDE|ENCAINIDE
C0966225|T129|302379|RXNORM|OMALIZUMAB|OMALIZUMAB
C0031422|T121|8136|RXNORM|PHENYLEPHRINE / THENYLDIAMINE|OXYPHENISATIN
C3538639|T121|1373216|RXNORM|2-BUTANOYLOXYBENZOATE|2-BUTANOYLOXYBENZOATE
C3668870|T121|1484856|RXNORM|CICUTA VIROSA WHOLE EXTRACT|CICUTA VIROSA WHOLE EXTRACT
C0041073|T121|1368168|RXNORM|TRIOLEIN|GLYCERYL TRIOLEATE
C3864832|T129|1596930|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 31 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 31 VACCINE
C0041087|T121|1368169|RXNORM|TRIPALMITIN|TRIPALMITIN
C3538641|T121|1373218|RXNORM|3-BROMOCAMPHOR, (+-)-|3-BROMOCAMPHOR, (+-)-
C2929248|T121|1008343|RXNORM|LACTATE / UREA|LACTATE / UREA
C2929248|T121|1008343|RXNORM|LACTATE / UREA|LACTATE / UREA
C2929811|T121|1008914|RXNORM|GLYCOL SALICYLATE / NIACIN|GLYCOL SALICYLATE / NIACIN
C2929812|T121|1008915|RXNORM|CAMPHOR / LIDOCAINE|CAMPHOR / LIDOCAINE
C2929813|T121|1008916|RXNORM|BENZOCAINE / BUTETAMATE|BENZOCAINE / BUTETAMATE
C2929814|T121|1008917|RXNORM|HYDROCORTISONE / TETRACYCLINE|HYDROCORTISONE / TETRACYCLINE
C2929807|T121|1008910|RXNORM|ETHAMIVAN / HEPTAMINOL / NORFENEFRINE|ETHAMIVAN / HEPTAMINOL / NORFENEFRINE
C2929808|T121|1008911|RXNORM|ASCORBIC ACID / CRANBERRY PREPARATION / VITAMIN E|ASCORBIC ACID / CRANBERRY PREPARATION / VITAMIN E
C2929809|T121|1008912|RXNORM|MAGNESIUM OXIDE / VITAMIN B6 / VITAMIN E|MAGNESIUM OXIDE / VITAMIN B6 / VITAMIN E
C2929810|T121|1008913|RXNORM|BENZALKONIUM / CHLOROXYLENOL / HYDROCORTISONE|BENZALKONIUM / CHLOROXYLENOL / HYDROCORTISONE
C0043355|T121|11371|RXNORM|XIPAMIDE|XIPAMIDE
C3695950|T109|1484852|RXNORM|C12-16 PARETH-9|C12-16 PARETH-9
C2929815|T121|1008918|RXNORM|CHLOROXYLENOL / TRICLOSAN|CHLOROXYLENOL / TRICLOSAN
C2929816|T121|1008919|RXNORM|SILICONES / SIMETHICONE|SILICONES / SIMETHICONE
C2183091|T121|821647|RXNORM|AMMONIUM CHLORIDE / DEXTROMETHORPHAN|AMMONIUM CHLORIDE / DEXTROMETHORPHAN
C3818735|T109|1495456|RXNORM|HYRIOPSIS CUMINGII WHOLE EXTRACT|HYRIOPSIS CUMINGII WHOLE EXTRACT
C3818737|T109|1495454|RXNORM|CARYOCAR BRASILIENSE FRUIT OIL|CARYOCAR BRASILIENSE FRUIT OIL
C0030817|T121|7975|RXNORM|PENICILLAMINE|PENICILLAMINE
C0034665|T121|9143|RXNORM|RANITIDINE|RANITIDINE
C0034665|T121|9143|RXNORM|RANITIDINE|RANITIDINE
C0030812|T121|7973|RXNORM|PENBUTOLOL|PENBUTOLOL
C0071773|T197|1365705|RXNORM|POTASSIUM NITRITE|POTASSIUM NITRITE
C2927881|T121|1006958|RXNORM|CAPSICUM EXTRACT / GARLIC PREPARATION|CAPSICUM EXTRACT / GARLIC PREPARATION
C2927882|T121|1006959|RXNORM|DEHYDROSANOL / TRIAMTERENE|DEHYDROSANOL / TRIAMTERENE
C1876818|T121|700807|RXNORM|DEXBROMPHENIRAMINE / PYRILAMINE|DEXBROMPHENIRAMINE / PYRILAMINE
C0023175|T196|6260|RXNORM|LEAD|LEAD
C2927875|T121|1006952|RXNORM|MEPROBAMATE / PENTAERYTHRITOL|MEPROBAMATE / PENTAERYTHRITOL
C2927876|T121|1006953|RXNORM|EUCALYPTUS EXTRACT / PEPPERMINT OIL|EUCALYPTUS EXTRACT / PEPPERMINT OIL
C2927873|T121|1006950|RXNORM|SODIUM NITRITE / VERATRUM VIRIDE PREPARATION|SODIUM NITRITE / VERATRUM VIRIDE PREPARATION
C2927874|T121|1006951|RXNORM|CAMPHOR / EUCALYPTOL / MENTHOL|CAMPHOR / EUCALYPTOL / MENTHOL
C2927879|T121|1006956|RXNORM|HYDROXYZINE / PENTAERYTHRITOL|HYDROXYZINE / PENTAERYTHRITOL
C2927880|T121|1006957|RXNORM|SWEETLEAF PREPARATION / ZINC ACETATE|SWEETLEAF PREPARATION / ZINC ACETATE
C2927877|T121|1006954|RXNORM|CARBON DIOXIDE / HELIUM / NITROGEN / OXYGEN|CARBON DIOXIDE / HELIUM / NITROGEN / OXYGEN
C2927878|T121|1006955|RXNORM|RUTIN / VINCAMINE|RUTIN / VINCAMINE
C0126120|T121|52151|RXNORM|LODOXAMIDE|LODOXAMIDE
C1827180|T121|687428|RXNORM|LAMIVUDINE / NEVIRAPINE / ZIDOVUDINE|LAMIVUDINE / NEVIRAPINE / ZIDOVUDINE
C3818746|T109|1494854|RXNORM|DECYLAMINE OXIDE|DECYLAMINE OXIDE
C0055435|T123|20852|RXNORM|CHLOROPHYLLIN|CHLOROPHYLLIN
C3488226|T121|1311361|RXNORM|SUS SCROFA EYE PREPARATION|PORCINE EYE PREPARATION
C0055443|T121|20859|RXNORM|CHLOROPROCAINE|CHLOROPROCAINE
C0304955|T197|91510|RXNORM|SODIUM CHROMATE CR51|SODIUM CHROMATE CR51
C0036860|T131|9724|RXNORM|CARBARYL|CARBARYL
C3256286|T109|1307956|RXNORM|MACADAMIA OIL|MACADAMIA OIL
C0087296|T197|42987|RXNORM|INDIUM IN-111 CHLORIDE|INDIUM IN-111 CHLORIDE
C0114873|T121|49276|RXNORM|DOXAZOSIN|DOXAZOSIN
C1706668|T129|997261|RXNORM|SIPULEUCEL-T|SIPULEUCEL-T
C3484455|T121|1427134|RXNORM|USTILAGO MAYDIS EXTRACT|USTILAGO MAYDIS EXTRACT
C0033798|T121|8896|RXNORM|PSEUDOEPHEDRINE|PSEUDOEPHEDRINE
C0543448|T123|142131|RXNORM|MAGNESIUM ASPARTATE|MAGNESIUM ASPARTATE
C3282677|T121|1427137|RXNORM|FORESKIN FIBROBLAST, NEONATAL|FORESKIN FIBROBLAST, NEONATAL
C3538265|T126|1372465|RXNORM|ACETYLCHOLINESTERASE HUMAN|ACETYLCHOLINESTERASE HUMAN
C1384520|T121|48274|RXNORM|ACETAMINOPHEN / PROPOXYPHENE|ACETAMINOPHEN / PROPOXYPHENE
C3535918|T109|1368618|RXNORM|GUAR HYDROXYPROPYLTRIMONIUM (1.7 SUBSTITUENTS PER SACCHARIDE)|GUAR HYDROXYPROPYLTRIMONIUM (1.7 SUBSTITUENTS PER SACCHARIDE)
C0055355|T121|20785|RXNORM|CHLORFENETHAZINE|CHLORFENETHAZINE
C0123163|T121|51296|RXNORM|IDEBENONE|IDEBENONE
C2080574|T121|820115|RXNORM|CAFFEINE / PHENYLPROPANOLAMINE|CAFFEINE / PHENYLPROPANOLAMINE
C0973456|T121|307387|RXNORM|PLUM PREPARATION|PLUM PREPARATION
C3858052|T121|1552342|RXNORM|NETUPITANT / PALONOSETRON|NETUPITANT / PALONOSETRON
C0062674|T121|26867|RXNORM|HEXOCYCLIUM|HEXOCYCLIUM
C0732290|T130|226724|RXNORM|[13C] UREA|UREA C-13
C2929548|T121|1008648|RXNORM|CAFFEINE / MECLIZINE|CAFFEINE / MECLIZINE
C2929549|T121|1008649|RXNORM|ANTIPYRINE / LIDOCAINE|ANTIPYRINE / LIDOCAINE
C2929544|T121|1008644|RXNORM|ACETAMINOPHEN / ATROPINE / CHLORPHENIRAMINE / PHENYLEPHRINE|ACETAMINOPHEN / ATROPINE / CHLORPHENIRAMINE / PHENYLEPHRINE
C2929545|T121|1008645|RXNORM|KAOLIN / SALICYLIC ACID|KAOLIN / SALICYLIC ACID
C2929546|T121|1008646|RXNORM|CLEMASTINE / CLOCORTOLONE|CLEMASTINE / CLOCORTOLONE
C2929547|T121|1008647|RXNORM|AJMALINE / DIHYDROERGOCRISTINE|AJMALINE / DIHYDROERGOCRISTINE
C2929540|T121|1008640|RXNORM|DIHYDRO-ALPHA-ERGOCRYPTINE / DIHYDRO-BETA-ERGOCRYPTINE / DIHYDROERGOCORNINE / DIHYDROERGOCRISTINE|DIHYDRO-ALPHA-ERGOCRYPTINE / DIHYDRO-BETA-ERGOCRYPTINE / DIHYDROERGOCORNINE / DIHYDROERGOCRISTINE
C2929541|T121|1008641|RXNORM|LIDOCAINE / NOREPINEPHRINE|LIDOCAINE / NOREPINEPHRINE
C2929542|T121|1008642|RXNORM|BETAMETHASONE / DIPHENYLPYRALINE|BETAMETHASONE / DIPHENYLPYRALINE
C2929543|T121|1008643|RXNORM|BETAINE / PEPSIN A|BETAINE / PEPSIN A
C0526783|T121|1367265|RXNORM|POLYSORBATE 40|POLYSORBATE 40
C2949504|T121|1046697|RXNORM|HEXYLRESORCINOL / MENTHOL|HEXYLRESORCINOL / MENTHOL
C0052944|T121|18751|RXNORM|BAMBUTEROL|BAMBUTEROL
C3535683|T109|1368342|RXNORM|PRICKLY PEAR FRUIT EXTRACT|PRICKLY PEAR FRUIT EXTRACT
C1690852|T195|1367269|RXNORM|PRADOFLOXACIN|PRADOFLOXACIN
C3538055|T121|1371948|RXNORM|DROSERA INTERMEDIA EXTRACT|DROSERA INTERMEDIA EXTRACT
C3256647|T109|1368343|RXNORM|PORPHYRA UMBILICALIS EXTRACT|PORPHYRA UMBILICALIS EXTRACT
C0076513|T121|38133|RXNORM|THIOPROPAZATE|THIOPROPAZATE
C0052946|T121|18753|RXNORM|BAMIPINE|BAMIPINE
C2739894|T129|897332|RXNORM|GROUNDSEL POLLEN EXTRACT|BACCHARIS HALIMIFOLIA POLLEN EXTRACT
C3496084|T121|1314275|RXNORM|THIOREDOXIN|THIOREDOXIN
C0050876|T121|17073|RXNORM|ADRENALONE|ADRENALONE
C3535866|T121|1370619|RXNORM|MYRISTOYL ISETHIONATE|MYRISTOYL ISETHIONATE
C2684343|T130|851906|RXNORM|BERMUDA GRASS POLLEN EXTRACT|CYNODON DACTYLON POLLEN EXTRACT
C0981980|T130|851902|RXNORM|TAG ALDER POLLEN EXTRACT|ALNUS INCANA SUBSP. RUGOSA POLLEN EXTRACT
C0085295|T129|1311299|RXNORM|INTERLEUKIN-10|INTERLEUKIN-10
C2741339|T129|900991|RXNORM|BUR OAK POLLEN EXTRACT|QUERCUS MACROCARPA POLLEN EXTRACT
C0005632|T121|1596|RXNORM|BISACODYL|BISACODYL
C0005632|T121|1596|RXNORM|BISACODYL|BISACODYL
C2741342|T129|900995|RXNORM|CHESNUT OAK POLLEN EXTRACT|QUERCUS MUEHLENBERGII POLLEN EXTRACT
C3486748|T121|1311291|RXNORM|DANIO RERIO EGG PREPARATION|DANIO RERIO EGG PREPARATION
C3486548|T197|1311292|RXNORM|CHROMIUM GLUCONATE|CHROMIUM GLUCONATE
C1950058|T197|1311293|RXNORM|FERROSOFERRIC PHOSPHATE|FERRUM PHOSPHORICUM PREPARATION
C2348724|T109|1307685|RXNORM|GALBANUM OIL|GALBANUM OIL
C0005640|T121|1598|RXNORM|DICUMAROL|DICUMAROL
C2828269|T197|1311296|RXNORM|FERROUS IODIDE|FERROUS IODIDE
C3486635|T197|1311297|RXNORM|GOLD TRICHLORIDE|GOLD TRICHLORIDE
C3256389|T121|1307961|RXNORM|CENTELLA ASIATICA LEAF EXTRACT|CENTELLA ASIATICA LEAF EXTRACT
C3255849|T121|1307960|RXNORM|LONICERA CAPRIFOLIUM FLOWER EXTRACT|LONICERA CAPRIFOLIUM FLOWER EXTRACT
C3528608|T121|1362703|RXNORM|BENZOCAINE / CETYLPYRIDINIUM / MENTHOL|BENZOCAINE / CETYLPYRIDINIUM / MENTHOL
C3495978|T121|1307965|RXNORM|CENTELLA ASIATICA LEAF HOMEOPATHIC PREPARATION|HYDROCOTYLE ASIATICA EXTRACT HOMEOPATHIC PREPARATION
C3256504|T121|1307964|RXNORM|ARNICA CORDIFOLIA FLOWER EXTRACT|ARNICA CORDIFOLIA FLOWER EXTRACT
C3257434|T121|1307967|RXNORM|FILIPENDULA ULMARIA ROOT EXTRACT|FILIPENDULA ULMARIA ROOT EXTRACT
C3256816|T121|1307966|RXNORM|VITIS VINIFERA SEED EXTRACT|VITIS VINIFERA SEED EXTRACT
C3256450|T121|1307969|RXNORM|TAMARIND SEED EXTRACT|TAMARIND SEED EXTRACT
C0304712|T121|91405|RXNORM|ERGOT PREPARATION|ERGOT PREPARATION
C1950689|T121|705259|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / PHENYLEPHRINE|ACETAMINOPHEN / DEXTROMETHORPHAN / PHENYLEPHRINE
C0175158|T121|62174|RXNORM|DESERPIDINE|DESERPIDINE
C0982073|T109|1311570|RXNORM|CETYL ESTERS WAX|CETYL ESTERS WAX
C3488066|T121|1310217|RXNORM|SOLANUM NIGRUM TOP EXTRACT|SOLANUM NIGRUM TOP EXTRACT
C3266928|T121|1310216|RXNORM|BLACK WIDOW SPIDER PREPARATION|BLACK WIDOW SPIDER PREPARATION
C3489324|T121|1310215|RXNORM|RUTA GRAVEOLENS WHOLE EXTRACT|RUTA GRAVEOLENS WHOLE EXTRACT
C2938581|T121|1310213|RXNORM|AMERICAN ELDERBERRY EXTRACT|AMERICAN ELDERBERRY EXTRACT
C3488688|T121|1309768|RXNORM|ASTRAGALUS NUTTALLII LEAF EXTRACT|ASTRAGALUS NUTTALLII LEAF EXTRACT
C2726135|T129|999384|RXNORM|ASPERGILLUS FLAVUS ALLERGENIC EXTRACT|ASPERGILLUS FLAVUS ALLERGENIC EXTRACT
C0013900|T123|1043181|RXNORM|ELLAGIC ACID|ELLAGIC ACID
C2947973|T121|1043184|RXNORM|ELLAGIC ACID / POMEGRANATE EXTRACT|ELLAGIC ACID / POMEGRANATE EXTRACT
C3538338|T109|1372563|RXNORM|ZINGIBER OFFICINALE WHOLE EXTRACT|ZINGIBER OFFICINALE WHOLE EXTRACT
C0781804|T121|242874|RXNORM|CONSTANT ALBICANS EXTRACT|CONSTANT ALBICANS EXTRACT
C0083220|T121|1311744|RXNORM|DESLORELIN|DESLORELIN
C0068451|T121|31538|RXNORM|NARINGIN|NARINGIN
C3535869|T130|1370615|RXNORM|BIS(1-METHYLAMYL) SULFOSUCCINATE|BIS(1-METHYLAMYL) SULFOSUCCINATE
C0076516|T121|38136|RXNORM|TISOPURINE|TISOPURINE
C3484574|T121|1311039|RXNORM|AMANITA MUSCARIA EXTRACT|AMANITA MUSCARIA EXTRACT
C3535870|T121|1370614|RXNORM|LAUROYL GLUTAMATE|LAUROYL GLUTAMATE
C0068978|T121|47589|RXNORM|CAFEDRINE|CAFEDRINE
C0293153|T121|85929|RXNORM|TELMESTEINE|TELMESTEINE
C0020740|T121|5640|RXNORM|IBUPROFEN|IBUPROFEN
C0020740|T121|5640|RXNORM|IBUPROFEN|IBUPROFEN
C1095803|T121|319780|RXNORM|CAPSICUM EXTRACT|CAPSICUM EXTRACT
C1095804|T121|319781|RXNORM|EUCALYPTUS EXTRACT|EUCALYPTUS EXTRACT
C0020752|T121|5645|RXNORM|ICHTHAMMOL|ICHTHAMMOL
C3695971|T122|1483690|RXNORM|DISODIUM (ETHOXYCARBONYL)PHOSPHONATE|DISODIUM (ETHOXYCARBONYL)PHOSPHONATE
C1620263|T121|614348|RXNORM|METFORMIN / ROSIGLITAZONE|METFORMIN / ROSIGLITAZONE
C3651761|T130|1428858|RXNORM|TETRADECAMETHYLHEXASILOXANE|TETRADECAMETHYLHEXASILOXANE
C3651762|T122|1428857|RXNORM|TRIS-BHT MESITYLENE|TRIS-BHT MESITYLENE
C0146556|T109|1428856|RXNORM|TREHALULOSE|TREHALULOSE
C3651763|T121|1428855|RXNORM|DESERT DATE EXTRACT|DESERT DATE EXTRACT
C0971023|T121|306266|RXNORM|ENTECAVIR|ENTECAVIR
C3540735|T109|1428853|RXNORM|CURCUMA LONGA WHOLE EXTRACT|CURCUMA LONGA EXTRACT
C3205127|T121|1150171|RXNORM|ASCORBIC ACID / CALCIUM CARBONATE|ASCORBIC ACID / CALCIUM CARBONATE
C3651766|T121|1428851|RXNORM|MONARDA DIDYMA LEAF EXTRACT|MONARDA DIDYMA LEAF EXTRACT
C2987510|T121|1428850|RXNORM|ARTEMISIA ABSINTHIUM EXTRACT|ARTEMISIA ABSINTHIUM EXTRACT
C3715210|T121|1541716|RXNORM|CORIANDRUM SATIVUM WHOLE EXTRACT|CORIANDRUM SATIVUM WHOLE EXTRACT
C0719849|T121||RXNORM|GLUCOSE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C3834096|T121|1541714|RXNORM|CIMICIFUGA SIMPLEX ROOT EXTRACT|CIMICIFUGA SIMPLEX ROOT EXTRACT
C3834095|T121|1541715|RXNORM|CITRUS AURANTIIFOLIA WHOLE EXTRACT|CITRUS AURANTIIFOLIA WHOLE EXTRACT
C3834097|T109|1541712|RXNORM|ZINGIBER CASSUMUNAR ROOT OIL|ZINGIBER CASSUMUNAR ROOT OIL
C3834099|T109|1541710|RXNORM|RUBUS IDAEUS FRUIT VOLATILE OIL|RUBUS IDAEUS FRUIT VOLATILE OIL
C3834098|T109|1541711|RXNORM|SANTALUM ALBUM SEED OIL|SANTALUM ALBUM SEED OIL
C3485042|T129|1304122|RXNORM|INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS|INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS
C3834093|T122|1541718|RXNORM|EREMOCITRUS GLAUCA FRUIT EXTRACT|EREMOCITRUS GLAUCA FRUIT EXTRACT
C3485046|T121|1304127|RXNORM|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-WISCONSIN-1-2010-LIKE VIRUS|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-WISCONSIN-1-2010-LIKE VIRUS
C3490348|T121|1545653|RXNORM|EMPAGLIFLOZIN|EMPAGLIFLOZIN
C0058831|T121|23744|RXNORM|DYCLONINE|DYCLONINE
C2016123|T121|812278|RXNORM|CHLORTHALIDONE / OXPRENOLOL|CHLORTHALIDONE / OXPRENOLOL
C2928387|T121|1007465|RXNORM|LACTOSE / MAGNESIUM PHOSPHATE|LACTOSE / MAGNESIUM PHOSPHATE
C2928386|T121|1007464|RXNORM|OXYPHENCYCLIMINE / PHENOBARBITAL|OXYPHENCYCLIMINE / PHENOBARBITAL
C3152885|T121|1098254|RXNORM|EASTERN COTTONWOOD POLLEN EXTRACT / PLAINS COTTONWOOD POLLEN EXTRACT|EASTERN COTTONWOOD POLLEN EXTRACT / PLAINS COTTONWOOD POLLEN EXTRACT
C2928388|T121|1007466|RXNORM|LYSINE / PHENYLALANINE|LYSINE / PHENYLALANINE
C2928383|T121|1007461|RXNORM|CLOCORTOLONE / SALICYLIC ACID|CLOCORTOLONE / SALICYLIC ACID
C2928382|T121|1007460|RXNORM|ASCORBIC ACID / DEQUALINIUM|ASCORBIC ACID / DEQUALINIUM
C2928384|T121|1007462|RXNORM|MAGNESIUM CITRATE / MAGNESIUM PHOSPHATE|MAGNESIUM CITRATE / MAGNESIUM PHOSPHATE
C2353951|T121|1488564|RXNORM|DAPAGLIFLOZIN|DAPAGLIFLOZIN
C2928391|T121|1007469|RXNORM|ETHAMIVAN / HEXOBENDINE|ETHAMIVAN / HEXOBENDINE
C2928390|T121|1007468|RXNORM|GUAIAZULENE / PANTOTHENIC ACID|GUAIAZULENE / PANTOTHENIC ACID
C0002026|T121|480|RXNORM|ALFENTANIL|ALFENTANIL
C0023992|T121|6468|RXNORM|LOPERAMIDE|LOPERAMIDE
C0023929|T121|6464|RXNORM|LOBELINE|LOBELINE
C0023961|T121|6465|RXNORM|LOFEPRAMINE|LOFEPRAMINE
C0023972|T121|6466|RXNORM|LOMUSTINE|LOMUSTINE
C3255299|T121|1236648|RXNORM|BIFIDOBACTERIUM BIFIDUM / BIFIDOBACTERIUM LONGUM|BIFIDOBACTERIUM BIFIDUM / BIFIDOBACTERIUM LONGUM
C3848546|T196|1546382|RXNORM|ARSENITE ION|ARSENITE ION
C1165386|T121|349762|RXNORM|EGG YOLK PHOSPHATIDES|EGG YOLK PHOSPHATIDES
C0014277|T121|3920|RXNORM|ENFLURANE|ENFLURANE
C3651723|T121|1430389|RXNORM|METHANOLAMINE|METHANOLAMINE
C0014310|T121|3925|RXNORM|ENOXACIN|ENOXACIN
C0053817|T121|19499|RXNORM|BITOLTEROL|BITOLTEROL
C0031855|T130|8302|RXNORM|PHYTIC ACID|PHYTIC ACID
C0072245|T121|34710|RXNORM|PROPYPHENAZONE|PROPYPHENAZONE
C3495428|T197|1362917|RXNORM|ALUMINUM SILICATE|ALUMINUM SILICATE
C0025270|T127|6728|RXNORM|VITAMIN K 3|VITAMIN K 3
C0031862|T127|8308|RXNORM|VITAMIN K 1|VITAMIN K 1
C1875218|T121|689443|RXNORM|IODINATED GLYCEROL / THEOPHYLLINE|IODINATED GLYCEROL / THEOPHYLLINE
C1875217|T121|689441|RXNORM|GLYCERIN / SODIUM CHLORIDE|GLYCERIN / SODIUM CHLORIDE
C0142931|T121|56524|RXNORM|SODIUM TARTRATE|SODIUM TARTRATE
C1509236|T121|1366817|RXNORM|ACETYLTRYPTOPHANATE|ACETYLTRYPTOPHANATE
C2727860|T129|889591|RXNORM|MACKEREL ALLERGENIC EXTRACT|SCOMBER SCOMBRUS ALLERGENIC EXTRACT
C0037659|T125|9939|RXNORM|SOMATOSTATIN|SOMATOSTATIN
C0118168|T121|50166|RXNORM|FOSINOPRIL|FOSINOPRIL
C0724544|T197|221069|RXNORM|CALCIUM CHLORIDE, DIHYDRATION|CALCIUM CHLORIDE, DIHYDRATION
C3192573|T121|1426635|RXNORM|STYPOCAULON SCOPARIUM PREPARATION|STYPOCAULON SCOPARIUM PREPARATION
C0036766|T007|1426634|RXNORM|SERRATIA MARCESCENS|SERRATIA MARCESCENS
C2981351|T121|1426636|RXNORM|LUTRELIN|LUTRELIN
C3486587|T121|1426631|RXNORM|RINFABATE|RINFABATE
C3256770|T109|1426630|RXNORM|GLYCERETH-26|GLYCERETH-26
C2955479|T121|1050324|RXNORM|HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / SODIUM PHOSPHATE, MONOBASIC|HYOSCYAMINE / METHENAMINE / METHYLENE BLUE / SODIUM PHOSPHATE, MONOBASIC
C3153178|T129|1426632|RXNORM|ULMUS RUBRA POLLEN ALLERGENIC EXTRACT|SLIPPERY ELM POLLEN ALLERGENIC EXTRACT
C3256057|T109|1307775|RXNORM|MAURITIA FLEXUOSA FRUIT OIL|MAURITIA FLEXUOSA FRUIT OIL
C2348030|T121|1307777|RXNORM|CYPERUS ROTUNDUS ROOT EXTRACT|CYPERUS ROTUNDUS ROOT EXTRACT
C3256020|T109|1307770|RXNORM|BETULA PUBESCENS RESIN|BETULA PUBESCENS RESIN
C3256144|T121|1307772|RXNORM|COPAIFERA OFFICINALIS RESIN|COPAIFERA OFFICINALIS RESIN
C3256336|T121|1307773|RXNORM|AMMONIUM LAURETH-3 SULFATE|AMMONIUM LAURETH-3 SULFATE
C3256120|T121|1307778|RXNORM|ALUMINUM DISTEARATE|ALUMINUM DISTEARATE
C3256279|T121|1307779|RXNORM|C14-22 ALCOHOLS|C14-22 ALCOHOLS
C0022487|T195|6099|RXNORM|KANAMYCIN|KANAMYCIN
C3857938|T121|1591895|RXNORM|BACKHOUSIA CITRIODORA WHOLE EXTRACT|BACKHOUSIA CITRIODORA WHOLE EXTRACT
C0018330|T121|1591890|RXNORM|GUANOSINE|GUANOSINE
C1572778|T121|1591891|RXNORM|PENTAFLUOROPROPANE|PENTAFLUOROPROPANE
C0717338|T121||RXNORM|ASPIRIN / BUTALBITAL / CAFFEINE
C3857939|T121|1591893|RXNORM|3-NONYLPHENOL|3-NONYLPHENOL
C0717335|T121|214156|RXNORM|ACETAMINOPHEN / PAMABROM / PYRILAMINE|ACETAMINOPHEN / PAMABROM / PYRILAMINE
C0044410|T127|12062|RXNORM|ALFACALCIDOL|ALFACALCIDOL
C0717332|T121|214153|RXNORM|ACETAMINOPHEN / DICHLORALPHENAZONE / ISOMETHEPTENE|ACETAMINOPHEN / DICHLORALPHENAZONE / ISOMETHEPTENE
C0010206|T121|2898|RXNORM|COUMARIN|COUMARIN
C3255651|T109|1306179|RXNORM|CETYL GLUCOSIDE|CETYL GLUCOSIDE
C3255650|T109|1306178|RXNORM|CETYL ETHYLHEXANOATE|CETYL ETHYLHEXANOATE
C0214439|T195|69256|RXNORM|MARBOFLOXACIN|MARBOFLOXACIN
C3255649|T109|1306175|RXNORM|CETYL BETAINE|CETYL BETAINE
C3255648|T109|1306174|RXNORM|CETETH-25|CETETH-25
C0360537|T121|108091|RXNORM|FLUCLOROLONE|FLUCLOROLONE
C3255645|T109|1306171|RXNORM|BAMBUSA VULGARIS STEM EXTRACT|BAMBUSA VULGARIS STEM EXTRACT
C3255644|T109|1306170|RXNORM|BAMBUSA VULGARIS SAP EXTRACT|BAMBUSA VULGARIS SAP EXTRACT
C3255647|T109|1306173|RXNORM|CETETH-24|CETETH-24
C3255646|T109|1306172|RXNORM|CETETH-16|CETETH-16
C1172734|T129|354770|RXNORM|NATALIZUMAB|NATALIZUMAB
C0982294|T121|314743|RXNORM|NUX VOMICA EXTRACT|NUX VOMICA EXTRACT
C0951745|T121|289497|RXNORM|ALPHA-GLUCOHEPTONIC ACID, MAGNESIUM SALT (2:1)|ALPHA-GLUCOHEPTONIC ACID, MAGNESIUM SALT (2:1)
C1532516|T121|483593|RXNORM|FLUPREDNIDENE / MICONAZOLE|FLUPREDNIDENE / MICONAZOLE
C3853658|T121|1551454|RXNORM|EPHEDRA SINICA STEM EXTRACT|EPHEDRA SINICA STEM EXTRACT
C0074799|T195|1551455|RXNORM|SOLASULFONE|SOLASULFONE
C3857962|T121|1551456|RXNORM|LYCOPODIUM COMPLANATUM SPORE EXTRACT|LYCOPODIUM COMPLANATUM SPORE EXTRACT
C3857961|T109|1551457|RXNORM|POTASSIUM METHOXYSALICYLATE|POTASSIUM METHOXYSALICYLATE
C3857960|T121|1551458|RXNORM|FORMALDEHYDE-SODIUM NAPHTHALENESULFONATE COPOLYMER (3000 MW)|FORMALDEHYDE-SODIUM NAPHTHALENESULFONATE COPOLYMER (3000 MW)
C0600175|T121|1546387|RXNORM|CARBAMOYLCHOLINE|CARBAMOYLCHOLINE
C2684348|T129|852834|RXNORM|KENTUCKY BLUEGRASS POLLEN EXTRACT|POA PRATENSIS POLLEN EXTRACT
C2741534|T129|901369|RXNORM|CULTIVATED MUSHROOM ALLERGENIC EXTRACT|CULTIVATED MUSHROOM ALLERGENIC EXTRACT
C2701522|T129|852343|RXNORM|QUACKGRASS POLLEN EXTRACT|ELYMUS REPENS POLLEN EXTRACT
C1874631|T121|690828|RXNORM|BUTABARBITAL / PHENOBARBITAL / SECOBARBITAL|BUTABARBITAL / PHENOBARBITAL / SECOBARBITAL
C1176315|T121|358262|RXNORM|FOSAMPRENAVIR|FOSAMPRENAVIR
C1176316|T121|358263|RXNORM|TADALAFIL|TADALAFIL
C1176316|T121|358263|RXNORM|TADALAFIL|TADALAFIL
C1874629|T121|690825|RXNORM|BUTABARBITAL / EPINEPHRINE / THEOPHYLLINE|BUTABARBITAL / EPINEPHRINE / THEOPHYLLINE
C1874628|T121|690824|RXNORM|BUTABARBITAL / EPHEDRINE / GUAIFENESIN / THEOPHYLLINE|BUTABARBITAL / EPHEDRINE / GUAIFENESIN / THEOPHYLLINE
C2701821|T129|852839|RXNORM|HOG SKIN EXTRACT|SUS SCROFA EPITHELIAL EXTRACT
C2701526|T129|852348|RXNORM|LOMBARD POPLAR POLLEN EXTRACT|POPULUS NIGRA POLLEN EXTRACT
C0008783|T121|2541|RXNORM|CIMETIDINE|CIMETIDINE
C0008777|T121|2540|RXNORM|CILASTATIN|CILASTATIN
C2741336|T129|900987|RXNORM|GARRYS OAK POLLEN EXTRACT|QUERCUS GARRYANA POLLEN EXTRACT
C1532737|T121|484211|RXNORM|EZETIMIBE / SIMVASTATIN|EZETIMIBE / SIMVASTATIN
C0533363|T123|1314424|RXNORM|FU LING|FU LING
C0770524|T121|235461|RXNORM|ALUMINUM SUBACETATE|ALUMINUM SUBACETATE
C0035823|T195|9462|RXNORM|ROLITETRACYCLINE|ROLITETRACYCLINE
C2928066|T121|1251740|RXNORM|LINSEED OIL / VITAMIN E|LINSEED OIL / VITAMIN E
C0527316|T121|135447|RXNORM|DONEPEZIL|DONEPEZIL
C0877777|T131|854163|RXNORM|EUROPEAN HONEY BEE VENOM PROTEIN|APIS MELLIFERA VENOM
C3256797|T121|1426950|RXNORM|OPUNTIA FICUS-INDICA EXTRACT|OPUNTIA FICUS-INDICA EXTRACT
C1720502|T121|645080|RXNORM|CHLORHEXIDINE / TETRACAINE|CHLORHEXIDINE / TETRACAINE
C2006345|T121|821890|RXNORM|CARBINOXAMINE / PHENYLPROPANOLAMINE / PYRILAMINE|CARBINOXAMINE / PHENYLPROPANOLAMINE / PYRILAMINE
C1572770|T121|1367077|RXNORM|NONOXYNOL-4 SULFATE|NONOXYNOL-4 SULFATE
C0074769|T197|36721|RXNORM|SODIUM SULFATE|SODIUM SULFATE
C0074771|T197|36723|RXNORM|SODIUM SULFITE|SODIUM SULFITE
C0012757|T121|3551|RXNORM|DISTIGMINE|DISTIGMINE
C0074774|T197|36726|RXNORM|SODIUM THIOSULFATE|THIOSULFURIC ACID, DISODIUM SALT
C0026794|T126|7094|RXNORM|MURAMIDASE|MURAMIDASE
C2741034|T129|900148|RXNORM|GIANT WILD RYE POLLEN EXTRACT|LEYMUS CONDENSATUS POLLEN EXTRACT
C2270172|T004|1324086|RXNORM|ASPERGILLUS RUBER|ASPERGILLUS RUBER
C0163655|T197|1423914|RXNORM|SILVER IODIDE|SILVER IODIDE
C0772387|T197|1423913|RXNORM|ANTIMONY TRIIODIDE|ANTIMONY TRIIODIDE
C2740606|T129|899390|RXNORM|BRUSSELS SPROUT ALLERGENIC EXTRACT|BRUSSELS SPROUT ALLERGENIC EXTRACT
C2702387|T129|1297535|RXNORM|WESTERN YELLOWJACKET VENOM PROTEIN|VESPULA PENSYLVANICA VENOM PROTEIN
C0178626|T121|62349|RXNORM|ETHACRYNATE|ETHACRYNATE
C2702385|T129|1297531|RXNORM|GERMAN WASP VENOM PROTEIN|VESPULA GERMANICA VENOM PROTEIN
C2702388|T129|1297533|RXNORM|SOUTHERN YELLOWJACKET VENOM PROTEIN|VESPULA SQUAMOSA VENOM PROTEIN
C1165560|T121|349908|RXNORM|CALCIUM CARBONATE, PRECIPITATED|CALCIUM CARBONATE, PRECIPITATED
C0054568|T121|20136|RXNORM|CAMYLOFINE|CAMYLOFIN
C0078839|T121|39993|RXNORM|ZOLPIDEM|ZOLPIDEM
C0078836|T121|39990|RXNORM|ZOFENOPRIL|ZOFENOPRIL
C0078840|T121|39994|RXNORM|ZOMEPIRAC|ZOMEPIRAC
C3831936|T109|1538143|RXNORM|PALMITOYLLYSYLVALYLDIAMINOBUTYRIC ACID|PALMITOYLLYSYLVALYLDIAMINOBUTYRIC ACID
C3486677|T121|1310173|RXNORM|RHUS GLABRA TOP EXTRACT|RHUS GLABRA TOP EXTRACT
C0078844|T121|39998|RXNORM|ZONISAMIDE|ZONISAMIDE
C3264823|T121|1243467|RXNORM|ACETONE / TEA TREE OIL|ACETONE / TEA TREE OIL
C0304597|T121|694012|RXNORM|UNDECYLENIC ACID / ZINC UNDECYLENATE|UNDECYLENIC ACID / ZINC UNDECYLENATE
C0453269|T121|125929|RXNORM|BILBERRY EXTRACT|BILBERRY EXTRACT
C0991800|T121|317206|RXNORM|CALCIUM CREOSOTATE|CALCIUM CREOSOTATE
C1660713|T121|604984|RXNORM|DEXTRAN / SODIUM CHLORIDE|DEXTRAN / SODIUM CHLORIDE
C0453260|T121|125921|RXNORM|GINGER ROOT|GINGER ROOT
C0913246|T121|278567|RXNORM|VALDECOXIB|VALDECOXIB
C2928042|T121|1007120|RXNORM|MAGNESIUM OXIDE / VITAMIN B6|MAGNESIUM OXIDE / VITAMIN B6
C2928043|T121|1007121|RXNORM|CHOLECALCIFEROL / VITAMIN A|CHOLECALCIFEROL / VITAMIN A
C2928044|T121|1007122|RXNORM|CAPSAICIN / MENTHOL|CAPSAICIN / MENTHOL
C1690962|T121|1007123|RXNORM|FERRIC AMMONIUM CITRATE / FOLIC ACID|FERRIC AMMONIUM CITRATE / FOLIC ACID
C2928047|T121|1007125|RXNORM|AMDINOCILLIN PIVOXIL / PIVAMPICILLIN|AMDINOCILLIN PIVOXIL / PIVAMPICILLIN
C2928048|T121|1007126|RXNORM|CLORAZEPATE / MAZINDOL|CLORAZEPATE / MAZINDOL
C2928049|T121|1007127|RXNORM|TRYPTOPHAN / VITAMIN B6|TRYPTOPHAN / VITAMIN B6
C2928050|T121|1007128|RXNORM|ALANINE / GLUTAMATE / GLYCINE|ALANINE / GLUTAMATE / GLYCINE
C2928051|T121|1007129|RXNORM|CALCIUM CITRATE / GLUTAMATE|CALCIUM CITRATE / GLUTAMATE
C3255615|T121|1314421|RXNORM|TRICAPRYLYL CITRATE|TRICAPRYLYL CITRATE
C0771936|T121|1309259|RXNORM|YARROW FLOWER EXTRACT|YARROW FLOWER EXTRACT
C0064161|T121|1309258|RXNORM|JOJOBA WAX|JOJOBA OIL
C2983857|T121|1309255|RXNORM|QUININE ARSENATE|QUININE ARSENATE
C2983862|T121|1309254|RXNORM|TETRAHEXYLDECYL ASCORBATE|TETRAHEXYLDECYL ASCORBATE
C3256742|T109|1309257|RXNORM|VACCINIUM MYRTILLUS LEAF EXTRACT|VACCINIUM MYRTILLUS LEAF EXTRACT
C1738282|T109|1309256|RXNORM|MEADOWFOAM OIL|MEADOWFOAM OIL
C0069449|T168|1309250|RXNORM|OLIVE OIL|OLIVE OIL
C0304108|T168|1309253|RXNORM|LEMON OIL|LEMON OIL
C0982306|T168|1309252|RXNORM|PALM KERNEL OIL|PALM KERNEL OIL
C3504634|T121|1356329|RXNORM|CAMPHOR / CAPSAICIN / MENTHOL / METHYL SALICYLATE / PEPPERMINT OIL / ZINC OXIDE|CAMPHOR / CAPSAICIN / MENTHOL / METHYL SALICYLATE / PEPPERMINT OIL / ZINC OXIDE
C1446936|T129|467329|RXNORM|USTILAGO MAYDIS ANTIGEN|USTILAGO MAYDIS ANTIGEN
C3256137|T109|1311605|RXNORM|CODIUM TOMENTOSUM EXTRACT|CODIUM TOMENTOSUM EXTRACT
C0071132|T121|33770|RXNORM|PIRETANIDE|PIRETANIDE
C0052657|T197|18516|RXNORM|ATTAPULGITE|ATTAPULGITE
C2928614|T121|1007698|RXNORM|ACETYLCYSTEINE / CEFUROXIME|ACETYLCYSTEINE / CEFUROXIME
C2928615|T121|1007699|RXNORM|CLOPAMIDE / RESERPINE|CLOPAMIDE / RESERPINE
C2928792|T121|1007878|RXNORM|HYDROXYZINE / LABETALOL|HYDROXYZINE / LABETALOL
C2928793|T121|1007879|RXNORM|ASCORBIC ACID / PHENOL|ASCORBIC ACID / PHENOL
C2928608|T121|1007692|RXNORM|PHENAZOPYRIDINE / SULFANILYLUREA|PHENAZOPYRIDINE / SULFANILYLUREA
C2928609|T121|1007693|RXNORM|ACETAMINOPHEN / FURSULTIAMIN|ACETAMINOPHEN / FURSULTIAMIN
C2928606|T121|1007690|RXNORM|BENZETHONIUM / LAURETH-9 / UREA|BENZETHONIUM / POLIDOCANOL / UREA
C2928607|T121|1007691|RXNORM|BROMHEXINE / CHLORPHENIRAMINE / ERYTHROMYCIN|BROMHEXINE / CHLORPHENIRAMINE / ERYTHROMYCIN
C2928786|T121|1007872|RXNORM|CLONIXIN / ERGOTAMINE|CLONIXIN / ERGOTAMINE
C2928613|T121|1007697|RXNORM|ALGINIC ACID / ZINC GLUCONATE|ALGINIC ACID / ZINC GLUCONATE
C2928784|T121|1007870|RXNORM|CINNARIZINE / DIHYDROERGOCRISTINE|CINNARIZINE / DIHYDROERGOCRISTINE
C2928611|T121|1007695|RXNORM|DIFEBARBAMATE / FEBARBAMATE / PHENOBARBITAL|DIFEBARBAMATE / FEBARBAMATE / PHENOBARBITAL
C0082607|T121|41126|RXNORM|FLUTICASONE|FLUTICASONE
C0082607|T121|41126|RXNORM|FLUTICASONE|FLUTICASONE
C0082607|T121|41126|RXNORM|FLUTICASONE|FLUTICASONE
C0443434|T109|1487139|RXNORM|1,1,2,2-TETRAFLUOROETHANE|1,1,2,2-TETRAFLUOROETHANE
C0034625|T196|1546450|RXNORM|RADIUM|RADIUM
C3256325|T109|1311603|RXNORM|ACETYLTRIETHYL CITRATE|ACETYLTRIETHYL CITRATE
C0068689|T197|31738|RXNORM|NICKEL SULFATE|NICKEL SULFATE
C1444901|T121|465678|RXNORM|FLUOROMETHOLONE / TOBRAMYCIN|FLUOROMETHOLONE / TOBRAMYCIN
C2001767|T197|1314219|RXNORM|LAPONITE|LAPONITE
C2954898|T121|1049136|RXNORM|COCOA BUTTER / ZINC OXIDE|COCOA BUTTER / ZINC OXIDE
C3256858|T109|1314212|RXNORM|PROPYLENE GLYCOL DIBENZOATE|PROPYLENE GLYCOL DIBENZOATE
C3256847|T121|1314211|RXNORM|LAURYL BETAINE|LAURYL BETAINE
C3256802|T109|1314210|RXNORM|PPG-9|PPG-9
C3256980|T121|1314216|RXNORM|NONOXYNOL-12|NONOXYNOL-12
C0301554|T121|89916|RXNORM|TERPIN HYDRATE|TERPIN HYDRATE
C0086008|T123|1314214|RXNORM|CHONDROITIN 4-SULFATE|CHONDROITIN 4-SULFATE
C0022034|T130|1546451|RXNORM|IOTHALAMIC ACID|IOTHALAMIC ACID
C3256486|T109|1311602|RXNORM|3,7-DIMETHYLOCTANAL|3,7-DIMETHYLOCTANAL
C0066548|T130|30021|RXNORM|MILD SILVER PROTEIN|MILD SILVER PROTEIN
C0006351|T121|1796|RXNORM|BUFEXAMAC|BUFEXAMAC
C0359075|T121|107005|RXNORM|METHYLPREDNISOLONE / NEOMYCIN|METHYLPREDNISOLONE / NEOMYCIN
C2974289|T121|1148495|RXNORM|CRIZOTINIB|CRIZOTINIB
C2929355|T121|1008451|RXNORM|ASCORBIC ACID / TETRACAINE / TYROTHRICIN|ASCORBIC ACID / TETRACAINE / TYROTHRICIN
C2929354|T121|1008450|RXNORM|BLACK IMPORTED FIRE ANT ALLERGENIC EXTRACT / RED IMPORTED FIRE ANT ALLERGENIC EXTRACT|BLACK IMPORTED FIRE ANT ALLERGENIC EXTRACT / RED IMPORTED FIRE ANT ALLERGENIC EXTRACT
C2929357|T121|1008453|RXNORM|BENZALKONIUM / MINERAL OIL / TRICLOSAN|BENZALKONIUM / MINERAL OIL / TRICLOSAN
C2929356|T121|1008452|RXNORM|CARISOPRODOL / DICLOFENAC|CARISOPRODOL / DICLOFENAC
C2929359|T121|1008455|RXNORM|AMINOQUINURIDE / TETRACAINE|AMINOQUINURIDE / TETRACAINE
C2929358|T121|1008454|RXNORM|DIHYDROCODEINE / PHENYLTOLOXAMINE|DIHYDROCODEINE / PHENYLTOLOXAMINE
C2929361|T121|1008457|RXNORM|GLYCINE / MAGNESIUM CHLORIDE|GLYCINE / MAGNESIUM CHLORIDE
C2929360|T121|1008456|RXNORM|HORSE HAIR EXTRACT / HORSE SKIN EXTRACT|HORSE HAIR EXTRACT / HORSE SKIN EXTRACT
C0529813|T121|1006619|RXNORM|EPRINOMECTIN|EPRINOMECTIN
C2929362|T121|1008458|RXNORM|ACRIFLAVINE / BENZOCAINE|ACRIFLAVINE / BENZOCAINE
C0059438|T121|24246|RXNORM|EPIGALLOCATECHIN GALLATE|EPIGALLOCATECHIN GALLATE
C1874018|T121|690212|RXNORM|ACETONE / ISOPROPYL ALCOHOL / POLYSORBATE 80|ACETONE / ISOPROPYL ALCOHOL / POLYSORBATE 80
C0005214|T121|1476|RXNORM|BETA-ESCIN|BETA-ESCIN
C0211011|T121|68503|RXNORM|ZICONOTIDE|ZICONOTIDE
C0057977|T121|23020|RXNORM|DIFEBARBAMATE|DIFEBARBAMATE
C3819175|T121|1534418|RXNORM|ACETAMINOPHEN / CARBIDOPA|ACETAMINOPHEN / CARBIDOPA
C0057981|T121|23024|RXNORM|DIFENOXIN|DIFENOXIN
C3848518|T121|1546453|RXNORM|ISOSULFAN BLUE INNER SALT|ISOSULFAN BLUE INNER SALT
C1962556|T121|725123|RXNORM|CARBOXYMETHYLCELLULOSE / GLYCERIN|CARBOXYMETHYLCELLULOSE / GLYCERIN
C3488982|T109|1309357|RXNORM|LEPTOSPERMUM PETERSONII LEAF OIL EXTRACT|LEPTOSPERMUM PETERSONII LEAF OIL EXTRACT
C3474072|T121|1358888|RXNORM|EUTERPE OLERACEA WHOLE EXTRACT|EUTERPE OLERACEA WHOLE EXTRACT
C0057233|T131|22374|RXNORM|DECAMETHRIN|DECAMETHRIN
C3163155|T121|1115788|RXNORM|ASCORBIC ACID / COPPER GLUCONATE / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / LUTEIN / VITAMIN E / ZEAXANTHIN / ZINC OXIDE|ASCORBIC ACID / COPPER GLUCONATE / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / LUTEIN / VITAMIN E / ZEAXANTHIN / ZINC OXIDE
C3485008|T121|1358889|RXNORM|EPIMEDIUM GRANDIFLORUM WHOLE EXTRACT|EPIMEDIUM GRANDIFLORUM WHOLE EXTRACT
C3152878|T129|1098247|RXNORM|PACIFIC SALMON ALLERGENIC EXTRACT|PINK SALMON ALLERGENIC EXTRACT
C3535655|T121|1369897|RXNORM|QUASSIA AMARA WHOLE EXTRACT|QUASSIA AMARA WHOLE EXTRACT
C1876824|T121|700821|RXNORM|HYDROCODONE / PSEUDOEPHEDRINE / TRIPROLIDINE|HYDROCODONE / PSEUDOEPHEDRINE / TRIPROLIDINE
C3535654|T121|1369898|RXNORM|LAURYL-MYRISTYL BENZOATE|LAURYL-MYRISTYL BENZOATE
C0068263|T123|1546454|RXNORM|VALERIC ACID|VALERIC ACID
C0064870|T121|28627|RXNORM|LEVOCABASTINE|LEVOCABASTINE
C0012458|T121|1487907|RXNORM|DINITOLMIDE|DINITOLMIDE
C0077857|T121|39230|RXNORM|URAPIDIL|URAPIDIL
C0059506|T121|24305|RXNORM|ERDOSTEINE|ERDOSTEINE
C0076607|T123|38217|RXNORM|THYMOMODULIN|THYMOMODULIN
C2949275|T121|1046312|RXNORM|BENZOCAINE / ETHANOL|BENZOCAINE / ETHANOL
C0063220|T121|1546455|RXNORM|HYPERICIN|HYPERICIN
C0063817|T130|27781|RXNORM|IOPROMIDE|IOPROMIDE
C2701339|T129|852136|RXNORM|JOHNSON GRASS POLLEN EXTRACT|SORGHUM HALEPENSE POLLEN EXTRACT
C0981977|T130|852132|RXNORM|SUGAR BEET POLLEN EXTRACT|BETA VULGARIS POLLEN EXTRACT
C2928971|T121|1008060|RXNORM|BUTALBITAL / CAFFEINE / CODEINE|BUTALBITAL / CAFFEINE / CODEINE
C2928972|T121|1008061|RXNORM|DEHYDROCHOLATE / HOMATROPINE|DEHYDROCHOLATE / HOMATROPINE
C2928973|T121|1008062|RXNORM|DEXTROMETHORPHAN / GUAIACOLSULFONIC ACID / PROMETHAZINE|DEXTROMETHORPHAN / GUAIACOLSULFONIC ACID / PROMETHAZINE
C2928974|T121|1008063|RXNORM|CARELESS WEED POLLEN EXTRACT / REDROOT PIGWEED POLLEN EXTRACT|CARELESS WEED POLLEN EXTRACT / REDROOT PIGWEED POLLEN EXTRACT
C2928975|T121|1008064|RXNORM|FOLIC ACID / VITAMIN B 12 / VITAMIN B6|FOLIC ACID / VITAMIN B 12 / VITAMIN B6
C0717768|T121|1008065|RXNORM|FERROUS SULFATE / FOLIC ACID|FERROUS SULFATE / FOLIC ACID
C2928977|T121|1008066|RXNORM|KETOCONAZOLE / SECNIDAZOLE|KETOCONAZOLE / SECNIDAZOLE
C2928978|T121|1008067|RXNORM|AMINOHYDROXYBUTYRIC ACID / PYRITHIOXIN|AMINOHYDROXYBUTYRIC ACID / PYRITHIOXIN
C2193914|T121|1008068|RXNORM|NAPHAZOLINE / NEOMYCIN|NAPHAZOLINE / NEOMYCIN
C2928979|T121|1008069|RXNORM|INDOMETHACIN / METHOCARBAMOL|INDOMETHACIN / METHOCARBAMOL
C0073393|T121|35636|RXNORM|RISPERIDONE|RISPERIDONE
C2728182|T129|1011021|RXNORM|OKRA ALLERGENIC EXTRACT|OKRA ALLERGENIC EXTRACT
C0070126|T121|32941|RXNORM|PARTHENOLIDE|PARTHENOLIDE
C2741251|T129|900704|RXNORM|BLUE SPRUCE POLLEN EXTRACT|PICEA PUNGENS POLLEN EXTRACT
C0058762|T121|23684|RXNORM|DROTAVERIN|DROTAVERINE
C1135662|T126|337623|RXNORM|DORNASE ALFA|DORNASE ALFA (DESOXYRIBONUCLEASE)
C3833143|T121|1540662|RXNORM|ALLANTOIN / LIDOCAINE / PETROLATUM|ALLANTOIN / LIDOCAINE / PETROLATUM
C0717916|T121|214703|RXNORM|METHYCLOTHIAZIDE / RESERPINE|METHYCLOTHIAZIDE / RESERPINE
C0078752|T121|39918|RXNORM|ZEAXANTHIN|ZEAXANTHIN
C0019468|T121|5301|RXNORM|HEXETIDINE|HEXETIDINE
C0717922|T121|214709|RXNORM|MINERAL OIL / PHENOLPHTHALEIN|MINERAL OIL / PHENOLPHTHALEIN
C3488966|T121|1309413|RXNORM|ASCLEPIAS TUBEROSA ROOT EXTRACT|ASCLEPIAS TUBEROSA ROOT EXTRACT
C3256291|T109|1309412|RXNORM|BUPLEURUM FALCATUM ROOT EXTRACT|BUPLEURUM FALCATUM ROOT EXTRACT
C3256657|T109|1309411|RXNORM|ARTEMISIA PRINCEPS LEAF EXTRACT|ARTEMISIA PRINCEPS LEAF EXTRACT
C0060787|T125|25357|RXNORM|FOLLITROPIN BETA|FOLLITROPIN BETA
C3256829|T109|1309417|RXNORM|CAREX HUMILIS ROOT EXTRACT|CAREX HUMILIS ROOT EXTRACT
C3464785|T109|1426407|RXNORM|PPG-2 MYRISTYL ETHER PROPIONATE|PPG-2 MYRISTYL ETHER PROPIONATE
C3256348|T109|1309415|RXNORM|CARICA PAPAYA LEAF EXTRACT|CARICA PAPAYA LEAF EXTRACT
C3256668|T109|1309414|RXNORM|CAMELLIA JAPONICA SEED EXTRACT|CAMELLIA JAPONICA SEED EXTRACT
C3644973|T121|1426158|RXNORM|GRINDELIA SQUARROSA FLOWERING TOP EXTRACT|GRINDELIA SQUARROSA FLOWERING TOP EXTRACT
C3644974|T122|1426159|RXNORM|DI-PPG-2 MYRETH-10 ADIPATE|DI-PPG-2 MYRETH-10 ADIPATE
C3256833|T109|1309419|RXNORM|DIOSCOREA COLLETTII VAR. HYPOGLAUCA ROOT EXTRACT|DIOSCOREA COLLETTII VAR. HYPOGLAUCA ROOT EXTRACT
C3256353|T109|1309418|RXNORM|CENTAUREA CYANUS FLOWER EXTRACT|CENTAUREA CYANUS FLOWER EXTRACT
C0165631|T121|60223|RXNORM|ADAPALENE|ADAPALENE
C2701721|T129|852663|RXNORM|SYRIAN HAMSTER SKIN EXTRACT|MESOCRICETUS AURATUS SKIN EXTRACT
C0032896|T121|8620|RXNORM|PRACTOLOL|PRACTOLOL
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, CALIFORNIA HAZELNUT POLLEN|PRASTERONE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, CALIFORNIA LIVE OAK|PRASTERONE
C3537691|T109|1371310|RXNORM|C12-15 ALCOHOLS|C12-15 ALCOHOLS
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, BOX ELDER|PRASTERONE
C2741294|T129|900770|RXNORM|LOBLOLLY PINE POLLEN EXTRACT|PINUS TAEDA POLLEN EXTRACT
C0206679|T005|1316105|RXNORM|HUMAN HERPESVIRUS 1|HUMAN HERPESVIRUS 1
C0205725|T005|1316104|RXNORM|HUMAN HERPESVIRUS 5 SPECIES|HUMAN HERPESVIRUS 5 SPECIES
C1880288|T121|734064|RXNORM|DESVENLAFAXINE|DESVENLAFAXINE
C0002937|T121|820|RXNORM|ANETHOLE TRITHIONE|ANETHOLE TRITHIONE
C2073887|T121|817322|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE
C0771402|T121|236156|RXNORM|FUMITORY EXTRACT|FUMITORY EXTRACT
C0032899|T121|8622|RXNORM|PRAJMALINE|PRAJMALINE
C0007903|T121|2284|RXNORM|CETRIMIDES|CETRIMIDES
C0007906|T121|2286|RXNORM|CETYLPYRIDINIUM|CETYLPYRIDINIUM
C0007906|T121|2286|RXNORM|CETYLPYRIDINIUM|CETYLPYRIDINIUM
C0054040|T121|19685|RXNORM|BRETYLIUM|BRETYLIUM
C0771400|T121|236154|RXNORM|BLACK CURRANT PREPARATION|BLACK CURRANT PREPARATION
C2344398|T121|798467|RXNORM|SMALLPOX VACCINE LIVE, NEW YORK CITY BOARD OF HEALTH VACCINIA STRAIN|SMALLPOX VACCINE LIVE, NEW YORK CITY BOARD OF HEALTH VACCINIA STRAIN
C1302059|T121|392512|RXNORM|CLOPAMIDE / PINDOLOL|CLOPAMIDE / PINDOLOL
C3864974|T121|1595248|RXNORM|HYALURONATE / LIDOCAINE|HYALURONATE / LIDOCAINE
C0085210|T121|42348|RXNORM|CANTHAXANTHIN|CANTHAXANTHIN
C3500588|T121|1314850|RXNORM|DIGITALIS PURPUREA WHOLE EXTRACT|DIGITALIS PURPUREA WHOLE EXTRACT
C3500590|T121|1314853|RXNORM|ELETTARIA CARDAMOMUM WHOLE EXTRACT|ELETTARIA CARDAMOMUM WHOLE EXTRACT
C3500592|T121|1314855|RXNORM|MENTHA ARVENSIS LEAF EXTRACT|MENTHA ARVENSIS LEAF EXTRACT
C3500591|T121|1314854|RXNORM|HAMAMELIS VIRGINIANA WHOLE EXTRACT|HAMAMELIS VIRGINIANA WHOLE EXTRACT
C0035549|T109|1314858|RXNORM|RIBOSE|RIBOSE
C2919955|T121|1370424|RXNORM|TETRADECYL HYDROGEN SULFATE (ESTER)|TETRADECYL HYDROGEN SULFATE (ESTER)
C2930154|T121|1370425|RXNORM|ALUMINUM ZIRCONIUM TRICHLOROHYDREX GLY|ALUMINUM ZIRCONIUM TRICHLOROHYDREX GLY
C1802535|T197|1370422|RXNORM|POTASH|POTASH
C2343882|T121|1370423|RXNORM|TRILAURETH-4 PHOSPHATE|TRILAURETH-4 PHOSPHATE
C0085208|T121|42347|RXNORM|BUPROPION|BUPROPION
C0085208|T121|42347|RXNORM|BUPROPION|BUPROPION
C0077497|T121|38967|RXNORM|TULOBUTEROL|TULOBUTEROL
C0051150|T121|17300|RXNORM|ALFUZOSIN|ALFUZOSIN
C0051150|T121|17300|RXNORM|ALFUZOSIN|ALFUZOSIN
C3474131|T121|1369702|RXNORM|COCO-CAPRYLATE-CAPRATE|COCO-CAPRYLATE-CAPRATE
C0051156|T121|17305|RXNORM|ALGINIC ACID|ALGINIC ACID
C0041289|T130|10908|RXNORM|TUBERCULIN|TUBERCULIN
C0982112|T109|314584|RXNORM|D-GLUCURONIC ACID|D-GLUCURONIC ACID
C0016576|T130|4537|RXNORM|FORMIC ACID|HYDROGEN CARBOXYLIC ACID
C0059771|T121|1483807|RXNORM|ETHYL LINOLENATE|ETHYL LINOLENATE
C2929835|T121|1008938|RXNORM|BELLADONNA ALKALOIDS / SIMETHICONE|BELLADONNA ALKALOIDS / SIMETHICONE
C2929836|T121|1008939|RXNORM|ASCORBIC ACID / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID|ASCORBIC ACID / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID
C2929833|T121|1008936|RXNORM|CALCIUM PHOSPHATE / GAMBOGE|CALCIUM PHOSPHATE / GAMBOGE
C2929834|T121|1008937|RXNORM|LACTATE / RESORCINOL / SALICYLIC ACID|LACTATE / RESORCINOL / SALICYLIC ACID
C2929831|T121|1008934|RXNORM|NIFLUMIC ACID / ORPHENADRINE|NIFLUMIC ACID / ORPHENADRINE
C2929832|T121|1008935|RXNORM|ACETAMINOPHEN / KETOPROFEN|ACETAMINOPHEN / KETOPROFEN
C2929829|T121|1008932|RXNORM|AMYLASES / CELLULASE / ENDOPEPTIDASES / LIPASE|AMYLASES / CELLULASE / ENDOPEPTIDASES / LIPASE
C2929830|T121|1008933|RXNORM|ACELLULAR PERTUSSIS VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / HAEMOPHILUS INFLUENZAE TYPE B, CAPSULAR POLYSACCHARIDE INACTIVATED TETANUS TOXOID CONJUGATE VACCINE / POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY) / POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1) / POLIOVIRUS VACCINE INACTIVATED, TYPE 3 (SAUKETT) / TETANUS TOXOID VACCINE, INACTIVATED|ACELLULAR PERTUSSIS VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / HAEMOPHILUS INFLUENZAE TYPE B, CAPSULAR POLYSACCHARIDE INACTIVATED TETANUS TOXOID CONJUGATE VACCINE / POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY) / POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1) / POLIOVIRUS VACCINE INACTIVATED, TYPE 3 (SAUKETT) / TETANUS TOXOID VACCINE, INACTIVATED
C2929827|T121|1008930|RXNORM|DEXAMETHASONE / PHENYLEPHRINE|DEXAMETHASONE / PHENYLEPHRINE
C2929828|T121|1008931|RXNORM|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / SCOPOLAMINE|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / SCOPOLAMINE
C2948906|T121|1045323|RXNORM|ALLANTOIN / GLYCERIN|ALLANTOIN / GLYCERIN
C3818734|T109|1495477|RXNORM|BIS-PEG PPG-16-16 PEG-PPG-16-16 DIMETHICONE|BIS-PEG PPG-16-16 PEG-PPG-16-16 DIMETHICONE
C3818733|T109|1495478|RXNORM|DIETHANOLAMINE OLETH-3 PHOSPHATE|DIETHANOLAMINE OLETH-3 PHOSPHATE
C0030454|T121|7910|RXNORM|PARAMETHASONE|PARAMETHASONE
C2929984|T121|1009089|RXNORM|BENZALKONIUM / BENZOCAINE|BENZALKONIUM / BENZOCAINE
C2929984|T121|1009089|RXNORM|BENZALKONIUM / BENZOCAINE|BENZALKONIUM / BENZOCAINE
C2929983|T121|1009088|RXNORM|GINSENG PREPARATION / ROYAL JELLY|GINSENG PREPARATION / ROYAL JELLY
C3834049|T109|1543455|RXNORM|METHOXY PEG PPG-7-3 AMINOPROPYL DIMETHICONE|METHOXY PEG PPG-7-3 AMINOPROPYL DIMETHICONE
C1874574|T121|690452|RXNORM|BISMUTH SUBCARBONATE / MORPHINE|BISMUTH SUBCARBONATE / MORPHINE
C0771514|T121|236259|RXNORM|POTASSIUM GLUCOHEPTONATE|POTASSIUM GLUCOHEPTONATE
C1874573|T121|690451|RXNORM|BISMUTH SUBCARBONATE / KAOLIN / PECTIN|BISMUTH SUBCARBONATE / KAOLIN / PECTIN
C2929976|T121|1009081|RXNORM|ALUMINUM HYDROXIDE / CALCIUM CARBONATE|ALUMINUM HYDROXIDE / CALCIUM CARBONATE
C2929975|T121|1009080|RXNORM|DICLOFENAC / TROXERUTIN|DICLOFENAC / TROXERUTIN
C2929978|T121|1009083|RXNORM|CALCIUM CITRATE / CALCIUM PHOSPHATE|CALCIUM CITRATE / CALCIUM PHOSPHATE
C2929977|T121|1009082|RXNORM|FERROUS FUMARATE / FERROUS GLUCONATE|FERROUS FUMARATE / FERROUS GLUCONATE
C2929980|T121|1009085|RXNORM|DEHYDROEPIANDROSTERONE / DICALCIUM PHOSPHATE|DICALCIUM PHOSPHATE / PRASTERONE
C2929979|T121|1009084|RXNORM|AMOXICILLIN / CLONIXIN|AMOXICILLIN / CLONIXIN
C0937917|T121|283810|RXNORM|BIMATOPROST|BIMATOPROST
C0937917|T121|283810|RXNORM|BIMATOPROST|BIMATOPROST
C2929981|T121|1009086|RXNORM|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / SODIUM METABISULFITE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / ASPARTATE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / SODIUM METABISULFITE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C0017507|T125|4792|RXNORM|GESTRINONE|GESTRINONE
C0017508|T121|4793|RXNORM|GESTRONOL|GESTRONOL
C3535926|T121|1368384|RXNORM|ALOGLIPTIN / METFORMIN|ALOGLIPTIN / METFORMIN
C3695968|T109|1483735|RXNORM|C11-15 PARETH-7|C11-15 PARETH-7
C3695967|T109|1483736|RXNORM|GLYCERETH-5 LACTATE|GLYCERETH-5 LACTATE
C0015821|T121|4325|RXNORM|FENBENDAZOLE|FENBENDAZOLE
C3273401|T126|1291609|RXNORM|TALIGLUCERASE ALFA|TALIGLUCERASE ALFA
C3535665|T197|1369404|RXNORM|COBALT ACETATE|COBALT ACETATE
C0064992|T121|28730|RXNORM|LIMONENE|LIMONENE
C0392428|T197|121070|RXNORM|CHROMIC PHOSPHATE P32|CHROMIC PHOSPHATE P32
C3256175|T109|1369405|RXNORM|PENTAERYTHRITOL TETRAKIS(3-(3,5-DI-TERT-BUTYL-4-HYDROXYPHENYL)PROPIONATE)|PENTAERYTHRITOL TETRAKIS(3-(3,5-DI-TERT-BUTYL-4-HYDROXYPHENYL)PROPIONATE)
C0076891|T121|38454|RXNORM|TRANDOLAPRIL|TRANDOLAPRIL
C0012390|T121|3449|RXNORM|DIMETHINDENE|DIMETHINDENE
C3160077|T121|1112447|RXNORM|HYDROQUINONE / LANOLIN|HYDROQUINONE / LANOLIN
C0057916|T125|22968|RXNORM|DIENOGEST|DIENOGEST
C0012383|T121|3445|RXNORM|DIMERCAPROL|DIMERCAPROL
C0012381|T121|3444|RXNORM|DIMENHYDRINATE|DIMENHYDRINATE
C0012384|T121|3446|RXNORM|SUCCIMER|MESO-2,3-DIMERCAPTOSUCCINIC ACID
C0003143|T121|865|RXNORM|ANTAZOLINE|ANTAZOLINE
C0012373|T121|3443|RXNORM|DILTIAZEM|DILTIAZEM
C0006983|T121|2020|RXNORM|CARBIMAZOLE|CARBIMAZOLE
C0006992|T121|2023|RXNORM|CARBOCYSTEINE|CARBOCYSTEINE
C0353946|T121|104129|RXNORM|ISPAGHULA HUSK|ISPAGHULA HUSK
C2146470|T121|814303|RXNORM|PHENYLEPHRINE / TROPICAMIDE|PHENYLEPHRINE / TROPICAMIDE
C2929566|T121|1008666|RXNORM|NIACINAMIDE / VITAMIN B6|NIACINAMIDE / VITAMIN B6
C2929567|T121|1008667|RXNORM|MAGNESIUM LACTATE / VITAMIN E|MAGNESIUM LACTATE / VITAMIN E
C2929564|T121|1008664|RXNORM|BENZALKONIUM / IDOXURIDINE|BENZALKONIUM / IDOXURIDINE
C2929565|T121|1008665|RXNORM|TROXERUTIN / VITAMIN E|TROXERUTIN / VITAMIN E
C2929562|T121|1008662|RXNORM|IODOQUINOL / SIMETHICONE|IODOQUINOL / SIMETHICONE
C2929563|T121|1008663|RXNORM|BISMUTH ALUMINATE / MAGNESIUM TRISILICATE|BISMUTH ALUMINATE / MAGNESIUM TRISILICATE
C2929560|T121|1008660|RXNORM|HYDROCORTISONE / LACTATE / UREA|HYDROCORTISONE / LACTATE / UREA
C2929561|T121|1008661|RXNORM|ICTASOL / SALICYLIC ACID|ICTASOL / SALICYLIC ACID
C0094813|T121|44532|RXNORM|TREPIBUTONE|TREPIBUTONE
C2701351|T129|852148|RXNORM|RIVER BIRCH POLLEN EXTRACT|RIVER BIRCH POLLEN EXTRACT
C2929568|T121|1008668|RXNORM|AMBROXOL / CEPHALEXIN|AMBROXOL / CEPHALEXIN
C2929569|T121|1008669|RXNORM|SULFACETAMIDE / VITAMIN B6|SULFACETAMIDE / VITAMIN B6
C2075715|T121|819757|RXNORM|AMBROXOL / CLENBUTEROL|AMBROXOL / CLENBUTEROL
C3272698|T121|1547220|RXNORM|ELIGLUSTAT|ELIGLUSTAT
C1875278|T121|689937|RXNORM|HYDROXYZINE / OXYPHENCYCLIMINE|HYDROXYZINE / OXYPHENCYCLIMINE
C1675411|T007|1372568|RXNORM|BACILLUS POLYFERMENTICUS|BACILLUS POLYFERMENTICUS
C3244899|T121|1370777|RXNORM|BIRD PEPPER EXTRACT|BIRD PEPPER EXTRACT
C1875275|T121|689934|RXNORM|HYDROXYETHYL CELLULOSE / POVIDONE|HYDROXYETHYL CELLULOSE / POVIDONE
C2928156|T121|1007234|RXNORM|DOLOMITE / MAGNESIUM SALT|DOLOMITE / MAGNESIUM SALT
C0302583|T196|90176|RXNORM|IRON|IRON
C0772462|T121|237124|RXNORM|SODIUM PHENOLSULFONATE|SODIUM PHENOLSULFONATE
C3668954|T121|1442699|RXNORM|MELILOTUS INDICUS WHOLE EXTRACT|MELILOTUS INDICUS WHOLE EXTRACT
C0772461|T121|237123|RXNORM|DIPOTASSIUM ADIPATE|DIPOTASSIUM ADIPATE
C2929493|T121|1008590|RXNORM|ALUMINUM HYDROXIDE / CALCIUM CARBONATE / MAGNESIUM HYDROXIDE / SIMETHICONE|ALUMINUM HYDROXIDE / CALCIUM CARBONATE / MAGNESIUM HYDROXIDE / SIMETHICONE
C2929494|T121|1008591|RXNORM|CYSTEINE / INOSITOL / METHIONINE / SODIUM PROPIONATE / UREA|CYSTEINE / INOSITOL / METHIONINE / SODIUM PROPIONATE / UREA
C2929495|T121|1008592|RXNORM|GUAIACOLSULFONATE / PHENYLEPHRINE|GUAIACOLSULFONATE / PHENYLEPHRINE
C2057681|T121|1008593|RXNORM|PAPAIN / TETRACYCLINE|PAPAIN / TETRACYCLINE
C2929496|T121|1008594|RXNORM|PROGLUMIDE / SULPIRIDE|PROGLUMIDE / SULPIRIDE
C2929497|T121|1008595|RXNORM|COAL TAR / TRIAMCINOLONE|COAL TAR / TRIAMCINOLONE
C2929498|T121|1008596|RXNORM|D-TRANSALLETHRIN / PIPERONYL BUTOXIDE|D-TRANSALLETHRIN / PIPERONYL BUTOXIDE
C2929499|T121|1008597|RXNORM|ASCORBIC ACID / PANTOTHENIC ACID|ASCORBIC ACID / PANTOTHENIC ACID
C2929500|T121|1008598|RXNORM|DICALCIUM PHOSPHATE / VITAMIN D|DICALCIUM PHOSPHATE / VITAMIN D
C2929501|T121|1008599|RXNORM|ASCORBIC ACID / PANTOTHENIC ACID / QUERCETIN|ASCORBIC ACID / PANTOTHENIC ACID / QUERCETIN
C3651781|T121|1428421|RXNORM|PLATANUS X ACERIFOLIA WHOLE EXTRACT|PLATANUS X ACERIFOLIA WHOLE EXTRACT
C0075470|T121|37289|RXNORM|SUCCINYLSULFATHIAZOLE|SUCCINYLSULFATHIAZOLE
C0076383|T121|38025|RXNORM|THENYLDIAMINE|THENYLDIAMINE
C3256121|T121|1372008|RXNORM|BITTER FENNEL EXTRACT|BITTER FENNEL EXTRACT
C0175035|T121|62153|RXNORM|EXAMETAZIME|EXAMETAZIME
C0076379|T121|38021|RXNORM|THEAFLAVIN|THEAFLAVIN
C0076380|T123|38022|RXNORM|THEANINE|THEANINE
C1337200|T168|1372002|RXNORM|BLACKBERRY FLAVOR|BLACKBERRY FLAVOR
C1337281|T109|1372003|RXNORM|BAMBOO EXTRACT|BAMBOO EXTRACT
C0772334|T121|1372000|RXNORM|CANADA BALSAM EXTRACT|CANADA BALSAM EXTRACT
C1095880|T109|1372001|RXNORM|HYDRANGEA EXTRACT|HYDRANGEA EXTRACT
C2980688|T121|1372006|RXNORM|ELM EXTRACT|ELM EXTRACT
C3256295|T109|1307145|RXNORM|CAPRYLHYDROXAMIC ACID|CAPRYLHYDROXAMIC ACID
C1576800|T121|1372004|RXNORM|MINT EXTRACT|MINT EXTRACT
C1644606|T109|1372005|RXNORM|DRAGON'S BLOOD EXTRACT|DRAGON'S BLOOD EXTRACT
C2756297|T129|967921|RXNORM|HOUSE FLY EXTRACT|HOUSE FLY EXTRACT
C1950715|T121|705279|RXNORM|OREGANO OIL|OREGANO OIL
C3854860|T121|1546706|RXNORM|PANDANUS TECTORIUS ROOT EXTRACT|PANDANUS TECTORIUS ROOT EXTRACT
C0304433|T121|91171|RXNORM|DIHYDRO-BETA-ERGOCRYPTINE|DIHYDRO-BETA-ERGOCRYPTINE
C0304432|T121|91170|RXNORM|DIHYDRO-ALPHA-ERGOCRYPTINE|DIHYDRO-ALPHA-ERGOCRYPTINE
C3485575|T121|1307142|RXNORM|RICINOLEAMIDOPROPYL ETHYLDIMONIUM ETHOSULFATE|RICINOLEAMIDOPROPYL ETHYLDIMONIUM ETHOSULFATE
C2608750|T121|1310235|RXNORM|SPIGELIA ANTHELMIA PREPARATION|SPIGELIA ANTHELMIA PREPARATION
C3495979|T121|1310238|RXNORM|BOS TAURUS ACHILLES TENDON PREPARATION|BOVINE ACHILLES TENDON PREPARATION
C3505486|T121|1358480|RXNORM|UNCARIA TOMENTOSA LEAF EXTRACT|UNCARIA TOMENTOSA LEAF EXTRACT
C0286185|T121|83213|RXNORM|MIBEFRADIL|MIBEFRADIL
C0007648|T123|2221|RXNORM|CELLULOSE|CELLULOSE
C2701347|T129|852144|RXNORM|CHERRY BIRCH POLLEN EXTRACT|BETULA LENTA POLLEN EXTRACT
C0042118|T121|1546707|RXNORM|USNIC ACID|USNIC ACID
C0252725|T197|1427055|RXNORM|COPPER CARBONATE|CUPRIC CARBONATE
C3832704|T197|1539374|RXNORM|UREA SULFATE|UREA SULFATE
C3205112|T121|1150152|RXNORM|QUERCETIN / RESVERATROL|QUERCETIN / RESVERATROL
C3864836|T109|1596688|RXNORM|SCLEROCARYA BIRREA SEED OIL|SCLEROCARYA BIRREA SEED OIL
C1633995|T121|608649|RXNORM|AMILORIDE / CYCLOPENTHIAZIDE|AMILORIDE / CYCLOPENTHIAZIDE
C3651749|T109|1428878|RXNORM|D-GLUTAMIC ACID|D-GLUTAMIC ACID
C0055561|T109|1368200|RXNORM|CHOLESTERYL OLEATE|CHOLESTERYL OLEATE
C2725875|T129|1098353|RXNORM|ORRIS ROOT ALLERGENIC EXTRACT|IRIS GERMANICA VAR. FLORENTINA ROOT ALLERGENIC EXTRACT
C3651753|T109|1428870|RXNORM|GLYCOL CETEARATE|GLYCOL CETEARATE
C0059737|T121|1358000|RXNORM|ETHYBENZTROPINE|ETHYBENZTROPINE
C3505163|T121|1358001|RXNORM|GAULTHERIA PROCUMBENS LEAF EXTRACT|GAULTHERIA PROCUMBENS LEAF EXTRACT
C3651751|T122|1428875|RXNORM|PEG-32 OLEATE|PEG-32 OLEATE
C3651752|T109|1428874|RXNORM|LAURYL GLYCOL HYDROXYPROPYL ETHER|LAURYL GLYCOL HYDROXYPROPYL ETHER
C3651750|T109|1428877|RXNORM|PPG-10 METHYL GLUCOSE ETHER|PPG-10 METHYL GLUCOSE ETHER
C1608551|T121|611247|RXNORM|FLUOXETINE / OLANZAPINE|FLUOXETINE / OLANZAPINE
C3864970|T121|1596454|RXNORM|BETAMETHASONE / CLOTRIMAZOLE / GENTAMICIN|BETAMETHASONE / CLOTRIMAZOLE / GENTAMICIN
C0080356|T121|40254|RXNORM|VALPROATE|VALPROATE
C2093603|T129|813859|RXNORM|RABBIT ALLERGENIC EXTRACT|RABBIT ALLERGENIC EXTRACT
C2723738|T129|867325|RXNORM|BLACK LOCUST POLLEN EXTRACT|ROBINIA PSEUDOACACIA POLLEN EXTRACT
C0065942|T129|29501|RXNORM|MENINGOCOCCAL GROUP A POLYSACCHARIDE|MENINGOCOCCAL GROUP A POLYSACCHARIDE
C2723734|T129|867321|RXNORM|RHODOTORULA RUBRA ALLERGENIC EXTRACT|RHODOTORULA RUBRA ALLERGENIC EXTRACT
C0065944|T129|29503|RXNORM|MENINGOCOCCAL GROUP C POLYSACCHARIDE|MENINGOCOCCAL GROUP C POLYSACCHARIDE
C0065199|T121|28908|RXNORM|LOXOPROFEN|LOXOPROFEN
C1176320|T130|1540828|RXNORM|PERFLEXANE|PERFLEXANE
C3833194|T109|1540827|RXNORM|CARDIOSPERMUM HALICACBUM WHOLE EXTRACT|CARDIOSPERMUM HALICACBUM WHOLE EXTRACT
C3833193|T109|1540826|RXNORM|BEHENYL ERUCATE|BEHENYL ERUCATE
C2744850|T121|1540825|RXNORM|TEDIZOLID|TEDIZOLID
C2194297|T121|812525|RXNORM|ASPIRIN / PHENOBARBITAL|ASPIRIN / PHENOBARBITAL
C3833192|T197|1540823|RXNORM|ESCARGOT SHELL, COOKED|ESCARGOT SHELL, COOKED
C0006304|T007|1540822|RXNORM|BRUCELLA ABORTUS|BRUCELLA ABORTUS
C0023863|T121|6446|RXNORM|LISURIDE|LISURIDE
C0025853|T121|6915|RXNORM|METOCLOPRAMIDE|METOCLOPRAMIDE
C0025854|T121|6916|RXNORM|METOLAZONE|METOLAZONE
C0025840|T121|6910|RXNORM|METHYPRYLON|METHYPRYLON
C0025842|T121|6911|RXNORM|METHYSERGIDE|METHYSERGIDE
C2928411|T121|1007489|RXNORM|FELODIPINE / METOPROLOL|FELODIPINE / METOPROLOL
C2928410|T121|1007488|RXNORM|DIPHENHYDRAMINE / PENTAERYTHRITOL|DIPHENHYDRAMINE / PENTAERYTHRITOL
C2928409|T121|1007487|RXNORM|FLUOCORTOLONE / SALICYLIC ACID|FLUOCORTOLONE / SALICYLIC ACID
C2928408|T121|1007486|RXNORM|CALCIUM ASCORBATE / CALCIUM THREONATE / FERROUS ASPARTO GLYCINATE / FERROUS FUMARATE / FOLIC ACID / SUCCINIC ACID / VITAMIN B 12|CALCIUM ASCORBATE / CALCIUM THREONATE / FERROUS ASPARTO GLYCINATE / FERROUS FUMARATE / FOLIC ACID / SUCCINIC ACID / VITAMIN B 12
C2928407|T121|1007485|RXNORM|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2928407|T121|1007485|RXNORM|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2928407|T121|1007485|RXNORM|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2928406|T121|1007484|RXNORM|DIHYDRALAZINE / PROPRANOLOL|DIHYDRALAZINE / PROPRANOLOL
C0025859|T121|6918|RXNORM|METOPROLOL|METOPROLOL
C2928404|T121|1007482|RXNORM|IBUPROFEN / LIDOCAINE|IBUPROFEN / LIDOCAINE
C2928403|T121|1007481|RXNORM|COLLAGEN / TRETINOIN|COLLAGEN / TRETINOIN
C2928402|T121|1007480|RXNORM|LIPASE / SIMETHICONE|LIPASE / SIMETHICONE
C3556199|T121|1373759|RXNORM|MONOFLUOROPHOSPHATE / SILICON DIOXIDE|MONOFLUOROPHOSPHATE / SILICON DIOXIDE
C3255863|T121|1426428|RXNORM|POLYGLYCERIN-3|POLYGLYCERIN-3
C3693000|T121|1442994|RXNORM|POTENTILLA ANSERINA WHOLE EXTRACT|POTENTILLA ANSERINA WHOLE EXTRACT
C3256639|T109|1426429|RXNORM|POLYMETHYLSILSESQUIOXANE (11 MICRONS)|POLYMETHYLSILSESQUIOXANE (11 MICRONS)
C3473982|T121|1314312|RXNORM|GLYCOL OLEATE|GLYCOL OLEATE
C3669288|T121|1442995|RXNORM|PRUNUS SPINOSA WHOLE EXTRACT|PRUNUS SPINOSA WHOLE EXTRACT
C2726164|T129|968502|RXNORM|TETRACOCCOSPORIUM PAXIANUM ALLERGENIC EXTRACT|TETRACOCCOSPORIUM PAXIANUM ALLERGENIC EXTRACT
C3474299|T121|1314313|RXNORM|SISYMBRIUM OFFICIANALE WHOLE EXTRACT|SISYMBRIUM OFFICIANALE WHOLE EXTRACT
C3529025|T121|1363991|RXNORM|LIMONENE, ()-|LIMONENE, ()-
C0060814|T121|1314310|RXNORM|FULVIC ACID|FULVIC ACID
C0981984|T129|867357|RXNORM|TRICHOPHYTON MENTAGROPHYTES EXTRACT|TRICHOPHYTON MENTAGROPHYTES EXTRACT
C0022237|T121|797541|RXNORM|ISOPROPYL ALCOHOL|ISOPROPYL ALCOHOL
C0022237|T121|797541|RXNORM|ISOPROPYL ALCOHOL|ISOPROPYL ALCOHOL
C0022237|T121|797541|RXNORM|ISOPROPYL ALCOHOL|ISOPROPYL ALCOHOL
C0053792|T121|19478|RXNORM|BISMUTH SUBSALICYLATE|BISMUTH SUBSALICYLATE
C0053792|T121|19478|RXNORM|BISMUTH SUBSALICYLATE|BISMUTH SUBSALICYLATE
C0872973|T121|259320|RXNORM|PLANT STANOL ESTER|PLANT STANOL ESTER
C0053790|T121|19476|RXNORM|BISMUTH SUBGALLATE|BISMUTH SUBGALLATE
C0053791|T197|19477|RXNORM|BISMUTH SUBNITRATE|BISMUTH SUBNITRATE
C0053789|T121|19475|RXNORM|BISMUTH SUBCARBONATE|BISMUTH SUBCARBONATE
C0053786|T197|19472|RXNORM|BISMUTH OXIDE|BISMUTH OXIDE
C3529028|T121|1363996|RXNORM|ISOSTEARYL ISOSTEARATE|ISOSTEARYL ISOSTEARATE
C1653588|T125|606396|RXNORM|HUMAN SECRETIN|HUMAN SECRETIN
C3489051|T121|1426420|RXNORM|LOXOSCELES RECLUSA PREPARATION|LOXOSCELES RECLUSA PREPARATION
C0031923|T121|8328|RXNORM|PILOCARPINE|PILOCARPINE
C0031923|T121|8328|RXNORM|PILOCARPINE|PILOCARPINE
C3256807|T121|1309470|RXNORM|SIMMONDSIA CHINESIS SEED EXTRACT|SIMMONDSIA CHINESIS SEED EXTRACT
C0025175|T125|6703|RXNORM|MEGESTROL|MEGESTROL
C1136867|T130|1426422|RXNORM|ACID VIOLET 43|EXT. D&C VIOLET NO. 2
C0071553|T125|34119|RXNORM|POLYESTRADIOL|POLYESTRADIOL
C3195253|T121|1119568|RXNORM|ASCORBIC ACID / CHOLECALCIFEROL / CUPROUS OXIDE / FOLIC ACID / MAGNESIUM OXIDE / NIACIN / POLYSACCHARIDE IRON COMPLEX / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / CHOLECALCIFEROL / CUPROUS OXIDE / FOLIC ACID / MAGNESIUM OXIDE / NIACIN / POLYSACCHARIDE IRON COMPLEX / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC OXIDE
C0037556|T121|9913|RXNORM|SODIUM TETRADECYL SULFATE|SODIUM TETRADECYL SULFATE
C3255815|T109|1426423|RXNORM|ZIZIPHUS EXTRACT|ZIZYPHUS
C0077656|T121|39085|RXNORM|UBIQUINOL|UBIQUINOL
C3255942|T109|1426424|RXNORM|HYDROLYZED WHEAT PROTEIN (ENZYMATIC, 3000 MW)|HYDROLYZED WHEAT PROTEIN (ENZYMATIC, 3000 MW)
C3486679|T121|1309973|RXNORM|RUBIA TINCTORUM ROOT EXTRACT|RUBIA TINCTORUM ROOT EXTRACT
C3529029|T121|1363997|RXNORM|TRIETHANOLAMINE BENZOATE|TRIETHANOLAMINE BENZOATE
C3255980|T109|1426425|RXNORM|SYNTHETIC WAX (1200 MW)|SYNTHETIC WAX (1200 MW)
C0059714|T121|24474|RXNORM|ETHINAMATE|ETHINAMATE
C3255865|T109|1426426|RXNORM|POLYISOBUTYLENE (1300 MW)|POLYISOBUTYLENE (1300 MW)
C2731902|T129|896246|RXNORM|DARK LEAVED MUGWORT POLLEN EXTRACT|ARTEMISIA LUDOVICIANA POLLEN EXTRACT
C3256462|T109|1309476|RXNORM|TANACETUM PARTHENIUM FLOWER EXTRACT|TANACETUM PARTHENIUM FLOWER EXTRACT
C3256403|T121|1307758|RXNORM|1,2-BUTANEDIOL|1,2-BUTANEDIOL
C3257506|T109|1307759|RXNORM|JUNIPERUS DEPPEANA WOOD OIL|JUNIPERUS DEPPEANA WOOD OIL
C3255597|T121|1307756|RXNORM|HAMAMELIS VIRGINIANA TOP EXTRACT|HAMAMELIS VIRGINIANA TOP EXTRACT
C3255889|T121|1307757|RXNORM|AMBROSIA PERUVIANA LEAF EXTRACT|AMBROSIA PERUVIANA LEAF EXTRACT
C3257503|T121|1307754|RXNORM|CINNAMOMUM CAMPHORA LEAF EXTRACT|CINNAMOMUM CAMPHORA LEAF EXTRACT
C3486290|T121|1307755|RXNORM|ILEX AQUIFOLIUM LEAF EXTRACT|ILEX AQUIFOLIUM LEAF EXTRACT
C3256166|T121|1307752|RXNORM|HAMAMELIS VIRGINIANA BARK EXTRACT|HAMAMELIS VIRGINIANA BARK EXTRACT
C3255697|T121|1307753|RXNORM|LONICERA JAPONICA FLOWER EXTRACT|LONICERA JAPONICA FLOWER EXTRACT
C3256092|T121|1307750|RXNORM|SCUTELLARIA BAICALENSIS ROOT EXTRACT|SCUTELLARIA BAICALENSIS ROOT EXTRACT
C2947522|T121|1041795|RXNORM|CHOLECALCIFEROL / OMEGA-3 ACID ETHYL ESTERS (USP)|CHOLECALCIFEROL / OMEGA-3 ACID ETHYL ESTERS (USP)
C2701661|T129|852585|RXNORM|CALIFORNIA JUNIPER POLLEN EXTRACT|JUNIPERUS CALIFORNICA POLLEN EXTRACT
C2939841|T129|1014191|RXNORM|CEDAR ELM POLLEN EXTRACT|ULMUS CRASSIFOLIA POLLEN EXTRACT
C2701657|T129|852581|RXNORM|MOUNTAIN CEDAR POLLEN EXTRACT|JUNIPERUS ASHEI POLLEN EXTRACT
C0717309|T121|214130|RXNORM|ACETAMINOPHEN / BUTALBITAL / CAFFEINE|ACETAMINOPHEN / BUTALBITAL / CAFFEINE
C2168930|T121|813694|RXNORM|QUININE / VITAMIN E|QUININE / VITAMIN E
C2701665|T129|852589|RXNORM|WESTERN JUNIPER POLLEN EXTRACT|JUNIPERUS OCCIDENTALIS POLLEN EXTRACT
C0717316|T121|214137|RXNORM|ACETAMINOPHEN / CAFFEINE / PYRILAMINE|ACETAMINOPHEN / CAFFEINE / PYRILAMINE
C2741287|T129|900758|RXNORM|PITCH PINE POLLEN EXTRACT|PINUS RIGIDA POLLEN EXTRACT
C0014806|T195|4053|RXNORM|ERYTHROMYCIN|ERYTHROMYCIN
C0014806|T195|4053|RXNORM|ERYTHROMYCIN|ERYTHROMYCIN
C0014806|T195|4053|RXNORM|ERYTHROMYCIN|ERYTHROMYCIN
C3692232|T122|1441535|RXNORM|SODIUM LAURETH-2 PHOSPHATE|SODIUM LAURETH-2 PHOSPHATE
C2723764|T129|867353|RXNORM|QUEEN PALM POLLEN EXTRACT|SYAGRUS ROMANZOFFIANA POLLEN EXTRACT
C0058636|T121|1094060|RXNORM|DODECYLBENZENESULFONIC ACID|DODECYLBENZENESULFONIC ACID
C2980850|T121|1094063|RXNORM|DODECYLBENZENESULFONIC ACID / LACTATE|DODECYLBENZENESULFONIC ACID / LACTATE
C0718207|T121|214970|RXNORM|ACETIC ACID / ALUMINUM ACETATE|ACETIC ACID / ALUMINUM ACETATE
C0284941|T121|82819|RXNORM|ACAMPROSATE|ACAMPROSATE
C0012963|T121|3616|RXNORM|DOBUTAMINE|DOBUTAMINE
C1445828|T121|466594|RXNORM|BENZOCAINE / TRICLOSAN|BENZOCAINE / TRICLOSAN
C1445827|T121|466593|RXNORM|BENZOCAINE / PHENOL|BENZOCAINE / PHENOL
C1875031|T121|690848|RXNORM|DIPHENHYDRAMINE / ZINC OXIDE|DIPHENHYDRAMINE / ZINC OXIDE
C2080621|T121|813109|RXNORM|PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE|PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE
C0073194|T130|1362930|RXNORM|RHODAMINE B|RHODAMINE B
C1815281|T121|669396|RXNORM|CARBETAPENTANE / DIPHENHYDRAMINE|CARBETAPENTANE / DIPHENHYDRAMINE
C1874642|T121|690841|RXNORM|CALAMINE / PHENOL / ZINC OXIDE|CALAMINE / PHENOL / ZINC OXIDE
C1875030|T121|690847|RXNORM|DIPHENHYDRAMINE / TRIPELENNAMINE|DIPHENHYDRAMINE / TRIPELENNAMINE
C0717898|T121|486895|RXNORM|MAGNESIUM AMINO ACID CHELATE|MAGNESIUM AMINO ACID CHELATE
C0000477|T121|897018|RXNORM|DALFAMPRIDINE|FAMPRIDINE
C3528960|T121|1363827|RXNORM|DISTEAROYLETHYL HYDROXYETHYLMONIUM METHOSULFATE|DISTEAROYLETHYL HYDROXYETHYLMONIUM METHOSULFATE
C0008864|T123|2567|RXNORM|CITRULLINE|CITRULLINE
C1816264|T121|672626|RXNORM|DEXBROMPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE|DEXBROMPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE
C3256233|T130|1425504|RXNORM|FD&C BLUE #10 ALUMINUM LAKE|FD&C BLUE #10 ALUMINUM LAKE
C0717742|T121|214540|RXNORM|EPHEDRINE / GUAIFENESIN / THEOPHYLLINE|EPHEDRINE / GUAIFENESIN / THEOPHYLLINE
C0043491|T197|11423|RXNORM|ZINC OXIDE|ZINC OXIDE
C0043491|T197|11423|RXNORM|ZINC OXIDE|ZINC OXIDE
C0043491|T197|11423|RXNORM|ZINC OXIDE|ZINC OXIDE
C0043490|T121|11422|RXNORM|ZINC OROTATE|ZINC OROTATE
C1872963|T121|718967|RXNORM|PAFURAMIDINE|PAFURAMIDINE
C0717743|T121|214541|RXNORM|EPHEDRINE / HYDROXYZINE / THEOPHYLLINE|EPHEDRINE / HYDROXYZINE / THEOPHYLLINE
C1453102|T121|473298|RXNORM|FIROCOXIB|FIROCOXIB
C3488426|T121|1424920|RXNORM|ATLANTIC HALIBUT PREPARATION|ATLANTIC HALIBUT PREPARATION
C2929608|T121|1191375|RXNORM|ALOE POLYSACCHARIDE / HYDROCORTISONE / IODOQUINOL|ALOE POLYSACCHARIDE / HYDROCORTISONE / IODOQUINOL
C0018242|T121|5021|RXNORM|GRISEOFULVIN|GRISEOFULVIN
C0771461|T121|236209|RXNORM|DIHEXYVERINE|DIHEXYVERINE
C0982276|T129|314725|RXNORM|MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP Y|MENINGOCOCCAL POLYSACCHARIDE VACCINE GROUP Y
C0016225|T121|4440|RXNORM|FLAVOXATE|FLAVOXATE
C0016229|T121|4441|RXNORM|FLECAINIDE|FLECAINIDE
C3811625|T109|1492326|RXNORM|EHRLICHIA CHAFFEENSIS EXTRACT|EHRLICHIA CHAFFEENSIS EXTRACT
C0038409|T007|1363920|RXNORM|STREPTOCOCCUS MUTANS|STREPTOCOCCUS MUTANS
C0016245|T121|4444|RXNORM|FLOCTAFENINE|FLOCTAFENINE
C0016267|T195|4448|RXNORM|FLOXACILLIN|FLOXACILLIN
C0771210|T126|235996|RXNORM|ERWINIA ASPARAGINASE|ERWINIA ASPARAGINASE
C0074757|T197|36709|RXNORM|SODIUM PHOSPHATE|SODIUM PHOSPHATE
C3244430|T121|1188531|RXNORM|CHLOPHEDIANOL / CHLORPHENIRAMINE / PSEUDOEPHEDRINE|CHLOPHEDIANOL / CHLORPHENIRAMINE / PSEUDOEPHEDRINE
C0633267|T109|1356759|RXNORM|RETINYL PROPIONATE|RETINYL PROPIONATE
C0717752|T125|214549|RXNORM|ESTROGENS, ESTERIFIED (USP)|ESTROGENS, ESTERIFIED (USP)
C2928541|T121|1007623|RXNORM|CLEMIZOLPENICILLIN / PENICILLIN G|CLEMIZOLPENICILLIN / PENICILLIN G
C0060135|T121|24812|RXNORM|FELBAMATE|FELBAMATE
C0600157|T123|155002|RXNORM|AMINOLEVULINATE|AMINOLEVULINATE
C1875775|T121|705062|RXNORM|SODIUM FLUORIDE / SODIUM PHOSPHATE|SODIUM FLUORIDE / SODIUM PHOSPHATE
C2194160|T121|819817|RXNORM|ASPIRIN / CYCLIZINE|ASPIRIN / CYCLIZINE
C2927924|T121|1007001|RXNORM|MEFRUSIDE / NIFEDIPINE|MEFRUSIDE / NIFEDIPINE
C3530536|T121|1364573|RXNORM|BENZYL ALCOHOL / MENTHOL|BENZYL ALCOHOL / MENTHOL
C0082966|T121|41289|RXNORM|IBUTILIDE|IBUTILIDE
C1875797|T121|705068|RXNORM|SULFUR / ZINC OXIDE / ZINC SULFATE|SULFUR / ZINC OXIDE / ZINC SULFATE
C2083540|T121|817466|RXNORM|ACETAMINOPHEN / THIOCOLCHICOSIDE|ACETAMINOPHEN / THIOCOLCHICOSIDE
C3486592|T121|1309780|RXNORM|CLERODENDRANTHUS SPICATUS LEAF EXTRACT|CLERODENDRANTHUS SPICATUS LEAF EXTRACT
C0163055|T121|59078|RXNORM|METAXALONE|METAXALONE
C1737290|T121|647235|RXNORM|GLIMEPIRIDE / PIOGLITAZONE|GLIMEPIRIDE / PIOGLITAZONE
C3860109|T121|1594580|RXNORM|MOMORDICA CHARANTIA WHOLE EXTRACT|MOMORDICA CHARANTIA WHOLE EXTRACT
C3555485|T122|1376451|RXNORM|C9-11 PARETH-6|C9-11 PARETH-6
C3555484|T109|1376452|RXNORM|HYDROXYETHYL CELLULOSE (1800 MPA.S AT 2%)|HYDROXYETHYL CELLULOSE (1800 MPA.S AT 2%)
C0078789|T197|1594583|RXNORM|ZINC PHOSPHIDE|ZINC PHOSPHIDE
C0076723|T121|38315|RXNORM|TIROPRAMIDE|TIROPRAMIDE
C3495351|T121|42662|RXNORM|EDETATE|EDETATE
C0991824|T121|317229|RXNORM|FERRIC CACODYLATE|FERRIC CACODYLATE
C2930035|T121|1009140|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLTOLOXAMINE|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLTOLOXAMINE
C2930036|T121|1009141|RXNORM|GLUCOSE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE / SODIUM PHOSPHATE, DIBASIC|GLUCOSE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM ACETATE / SODIUM CHLORIDE / SODIUM GLUCONATE / SODIUM PHOSPHATE, DIBASIC
C2930037|T121|1009142|RXNORM|LOTEPREDNOL ETABONATE / TOBRAMYCIN|LOTEPREDNOL ETABONATE / TOBRAMYCIN
C2930038|T121|1009143|RXNORM|UBIQUINONE / VITAMIN E|UBIQUINONE / VITAMIN E
C0002503|T130|645|RXNORM|AMINACRINE|AMINACRINE
C0069679|T121|1547630|RXNORM|OSTHOL|OSTHOL
C2930041|T121|1009148|RXNORM|AMPICILLIN / SULBACTAM|AMPICILLIN / SULBACTAM
C2930042|T121|1009149|RXNORM|ALUMINUM HYDROXIDE / MAGNESIUM HYDROXIDE|ALUMINUM HYDROXIDE / MAGNESIUM HYDROXIDE
C0301499|T121|1440290|RXNORM|FERROUS CARBONATE|FERROUS CARBONATE
C2928030|T121|1007108|RXNORM|DICLOFENAC / PRIDINOL|DICLOFENAC / PRIDINOL
C2928031|T121|1007109|RXNORM|CHLORAMPHENICOL / RESORCINOL / SALICYLIC ACID|CHLORAMPHENICOL / RESORCINOL / SALICYLIC ACID
C0903898|T121|274332|RXNORM|NATEGLINIDE|NATEGLINIDE
C2928024|T121|1007102|RXNORM|ISOPROPAMIDE / TRIFLUOPERAZINE|ISOPROPAMIDE / TRIFLUOPERAZINE
C2928025|T121|1007103|RXNORM|MENINGOCOCCAL GROUP C POLYSACCHARIDE / MENINGOCOCCAL VACCINE B|MENINGOCOCCAL GROUP C POLYSACCHARIDE / MENINGOCOCCAL VACCINE B
C2928023|T121|1007100|RXNORM|CHOLINE / POLYETHYLENE GLYCOLS|CHOLINE / POLYETHYLENE GLYCOLS
C2057675|T121|1007101|RXNORM|DIPYRONE / TETRACYCLINE|DIPYRONE / TETRACYCLINE
C2928029|T121|1007107|RXNORM|MENINGOCOCCAL GROUP A POLYSACCHARIDE / MENINGOCOCCAL GROUP C POLYSACCHARIDE|MENINGOCOCCAL GROUP A POLYSACCHARIDE / MENINGOCOCCAL GROUP C POLYSACCHARIDE
C2928026|T121|1007104|RXNORM|CAMYLOFINE / DIPYRONE|CAMYLOFINE / DIPYRONE
C2928027|T121|1007105|RXNORM|ASTEMIZOLE / DEXAMETHASONE|ASTEMIZOLE / DEXAMETHASONE
C0287573|T121|83682|RXNORM|CEFDITOREN|CEFDITOREN
C1875672|T121|689954|RXNORM|POLYETHYLENE GLYCOLS / POLYVINYL ALCOHOL|POLYETHYLENE GLYCOLS / POLYVINYL ALCOHOL
C0039855|T121|10464|RXNORM|THIAMYLAL|THIAMYLAL
C0023025|T123|1442199|RXNORM|LANOSTEROL|LANOSTEROL
C0065642|T197|29261|RXNORM|MANGANESE CHLORIDE|MANGANESE CHLORIDE
C1875671|T121|689953|RXNORM|POLYETHYLENE GLYCOL 400 / PROPYLENE GLYCOL|POLYETHYLENE GLYCOL 400 / PROPYLENE GLYCOL
C0065644|T197|29263|RXNORM|MANGANESE DIOXIDE|MANGANESE DIOXIDE
C3555492|T121|1376213|RXNORM|CARTHAMUS TINCTORIUS FLOWER BUD EXTRACT|CARTHAMUS TINCTORIUS FLOWER BUD EXTRACT
C0065649|T197|29268|RXNORM|MANGANESE SULFATE|MANGANESE SULFATE
C1875673|T121|689958|RXNORM|POLYVINYL ALCOHOL / POVIDONE|POLYVINYL ALCOHOL / POVIDONE
C3555493|T121|1376212|RXNORM|GARCINIA INDICA FRUIT EXTRACT|GARCINIA INDICA FRUIT EXTRACT
C2722896|T126|1427034|RXNORM|PANCRELIPASE PROTEASE|PANCRELIPASE PROTEASE
C0982128|T121|314599|RXNORM|DISOFENIN|DISOFENIN
C2740590|T129|899363|RXNORM|BLACK PEPPER ALLERGENIC EXTRACT|PIPER NIGRUM ALLERGENIC EXTRACT
C2722894|T126|1427033|RXNORM|PANCRELIPASE AMYLASE|PANCRELIPASE AMYLASE
C2722043|T129|975509|RXNORM|SQUASH ALLERGENIC EXTRACT|CUCURBITA MAXIMA ALLERGENIC EXTRACT
C0982121|T121|314592|RXNORM|DILTIAZEM MALEATE|DILTIAZEM MALEATE
C0597206|T121|1495318|RXNORM|PHENOLATE|PHENOLATE
C3818738|T109|1495319|RXNORM|P-DODECYLBENZENESULFONIC ACID|P-DODECYLBENZENESULFONIC ACID
C3695964|T121|1484143|RXNORM|ACACIA SENEGAL FLOWER EXTRACT|ACACIA SENEGAL FLOWER EXTRACT
C3535895|T121|1370585|RXNORM|PALMITOYL GLUTAMATE|PALMITOYL GLUTAMATE
C0772067|T121|236757|RXNORM|PHOSPHOLIPID,BEEF|PHOSPHOLIPID,BEEF
C0137757|T121|54908|RXNORM|POLICRESULEN|POLICRESULEN
C3692542|T121|1442193|RXNORM|BOS TAURUS EYE PREPARATION|BOS TAURUS EYE PREPARATION
C0162745|T126|58939|RXNORM|COLLAGENASE|COLLAGENASE
C0075210|T121|37075|RXNORM|ETHINYL ESTRADIOL / NORGESTREL|ETHINYL ESTRADIOL / NORGESTREL
C0071115|T121|33753|RXNORM|PIPERONAL|PIPERONAL
C3256429|T121|1372264|RXNORM|EASTERN WHITE PINE EXTRACT|PINUS STROBUS EXTRACT
C0939905|T121|285251|RXNORM|OATS PREPARATION|OATS PREPARATION
C2928733|T121|1007818|RXNORM|CALCIUM GLUCEPTATE / CALCIUM GLUCONATE|CALCIUM GLUCEPTATE / CALCIUM GLUCONATE
C2928734|T121|1007819|RXNORM|CALCIUM CARBONATE / CALCIUM GLUBIONATE|CALCIUM CARBONATE / CALCIUM GLUBIONATE
C2344297|T129|798268|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 6 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 6 VACCINE
C3665364|T121|1442191|RXNORM|ARGEMONE MEXICANA WHOLE EXTRACT|ARGEMONE MEXICANA WHOLE EXTRACT
C0163069|T121|59087|RXNORM|EUCALYPTUS OIL|EUCALYPTUS OIL
C0163069|T121|59087|RXNORM|EUCALYPTUS OIL|EUCALYPTUS OIL
C2728177|T129|1012026|RXNORM|VEAL ALLERGENIC EXTRACT|VEAL ALLERGENIC EXTRACT
C2928728|T121|1007813|RXNORM|AMOXICILLIN / BROMHEXINE|AMOXICILLIN / BROMHEXINE
C2928729|T121|1007814|RXNORM|CYPROTERONE / ETHINYL ESTRADIOL|CYPROTERONE / ETHINYL ESTRADIOL
C2928730|T121|1007815|RXNORM|ACETAMINOPHEN / CAFFEINE / SALICYLIC ACID|ACETAMINOPHEN / CAFFEINE / SALICYLIC ACID
C2928731|T121|1007816|RXNORM|PHENOBARBITAL / PROPANTHELINE|PHENOBARBITAL / PROPANTHELINE
C2928732|T121|1007817|RXNORM|SULFALENE / TRIMETHOPRIM|SULFALENE / TRIMETHOPRIM
C2730252|T129|892661|RXNORM|RICE (WHOLE GRAIN) ALLERGENIC EXTRACT|RICE (WHOLE GRAIN) ALLERGENIC EXTRACT
C3255812|T121|1372260|RXNORM|SPANISH CHESTNUT EXTRACT|SPANISH CHESTNUT EXTRACT
C1699439|T121|617772|RXNORM|ACETAMINOPHEN / PHENIRAMINE / PHENYLEPHRINE|ACETAMINOPHEN / PHENIRAMINE / PHENYLEPHRINE
C0006837|T004|1963|RXNORM|CANDIDA ALBICANS|CANDIDA ALBICANS
C0915082|T121|1314235|RXNORM|ISOPULEGOL|ISOPULEGOL
C3282687|T121|1314234|RXNORM|POLYQUATERNIUM 37 (200 MPA.S)|POLYQUATERNIUM 37 (200 MPA.S)
C3496037|T121|1314237|RXNORM|BOS TAURUS BONE MARROW PREPARATION|BOVINE BONE MARROW PREPARATION
C0766326|T121|233698|RXNORM|DRONEDARONE|DRONEDARONE
C3282852|T122|1314231|RXNORM|PYRIDOXINE DIPALMITATE|PYRIDOXINE DIPALMITATE
C3473398|T121|1314230|RXNORM|PEG-4 DIHEPTANOATE|PEG-4 DIHEPTANOATE
C3496663|T121|1314233|RXNORM|PREZATIDE COPPER|PREZATIDE COPPER
C3474240|T109|1314232|RXNORM|UNDECYLENIC ACID MONOETHANOLAMIDE|UNDECYLENIC ACID MONOETHANOLAMIDE
C2080605|T121|815641|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN / PHENYLPROPANOLAMINE / PYRILAMINE|DEXTROMETHORPHAN / GUAIFENESIN / PHENYLPROPANOLAMINE / PYRILAMINE
C0072221|T130|1314239|RXNORM|PROPYLENE|PROPYLENE
C3500338|T121|1314238|RXNORM|VACCINIUM VITIS-IDAEA LEAF EXTRACT|VACCINIUM VITIS-IDAEA LEAF EXTRACT
C0001159|T121|1441664|RXNORM|ACONITINE|ACONITINE
C3669135|T121|1441660|RXNORM|OXALATE|OXALATE
C3486147|T121|1305199|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / BIOTIN / DEXPANTHENOL / ERGOCALCIFEROL / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN K 1|ALPHA TOCOPHEROL / ASCORBIC ACID / BIOTIN / DEXPANTHENOL / ERGOCALCIFEROL / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN K 1
C0075870|T195|37617|RXNORM|TAZOBACTAM|TAZOBACTAM
C2978568|T121|1089112|RXNORM|BACITRACIN / DIMETHICONE / ZINC OXIDE|BACITRACIN / DIMETHICONE / ZINC OXIDE
C1657828|T121|605570|RXNORM|CARBINOXAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE|CARBINOXAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE
C0066522|T126|29998|RXNORM|OCRIPLASMIN|OCRIPLASMIN
C3851350|T121|1591922|RXNORM|LEDIPASVIR|LEDIPASVIR
C0071114|T121|33752|RXNORM|PIPEROCAINE|PIPEROCAINE
C0066520|T121|29996|RXNORM|MICRONOMICIN|MICRONOMICIN
C0005324|T121|1523|RXNORM|BETHANIDINE|BETHANIDINE
C3473401|T121|1352512|RXNORM|ABELMOSCHUS MOSCHATUS SEED EXTRACT|ABELMOSCHUS MOSCHATUS SEED EXTRACT
C2929343|T121|1008439|RXNORM|ASCORBIC ACID / NIACINAMIDE|ASCORBIC ACID / NIACINAMIDE
C2929342|T121|1008438|RXNORM|HESPERIDIN / RUTIN|HESPERIDIN / RUTIN
C2929337|T121|1008433|RXNORM|BENZOCAINE / BISMUTH SUBGALLATE / ZINC OXIDE|BENZOCAINE / BISMUTH SUBGALLATE / ZINC OXIDE
C2929336|T121|1008432|RXNORM|FORMALDEHYDE / SODIUM FLUORIDE|FORMALDEHYDE / SODIUM FLUORIDE
C2929335|T121|1008431|RXNORM|ADRENALONE / TETRACAINE|ADRENALONE / TETRACAINE
C2929334|T121|1008430|RXNORM|COAL TAR / PYRITHIONE|COAL TAR / PYRITHIONE
C2929341|T121|1008437|RXNORM|DIHYDROERGOTAMINE / TROXERUTIN|DIHYDROERGOTAMINE / TROXERUTIN
C2929340|T121|1008436|RXNORM|GLYCOPYRROLATE / PHENOBARBITAL|GLYCOPYRROLATE / PHENOBARBITAL
C2929339|T121|1008435|RXNORM|LICORICE / UNDECYLENATE|LICORICE / UNDECYLENATE
C2929338|T121|1008434|RXNORM|METHYLNICOTINATE / PHENYLBUTAZONE / PIPERAZINE|METHYLNICOTINATE / PHENYLBUTAZONE / PIPERAZINE
C0005088|T121|1418|RXNORM|BENZOYL PEROXIDE|BENZOYL PEROXIDE
C3848581|T196|1546167|RXNORM|ANTIMONY CATION (3+)|ANTIMONY CATION (3+)
C1874521|T121|690271|RXNORM|BENZOCAINE / METHYL SALICYLATE|BENZOCAINE / METHYL SALICYLATE
C1874524|T121|690276|RXNORM|BENZOCAINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE|BENZOCAINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C2928877|T121|1007964|RXNORM|LYSINE / ZINC OXIDE|LYSINE / ZINC OXIDE
C2701804|T129|852802|RXNORM|CALIFORNIA SCRUB OAK POLLEN EXTRACT|QUERCUS DUMOSA POLLEN EXTRACT
C0063204|T121|27306|RXNORM|HYLAN|HYLAN
C2928878|T121|1007965|RXNORM|ACETAMINOPHEN / CAFFEINE / HOMATROPINE|ACETAMINOPHEN / CAFFEINE / HOMATROPINE
C2928879|T121|1007966|RXNORM|ALUMINUM OXIDE / SIMETHICONE|ALUMINUM OXIDE / SIMETHICONE
C3503778|T121|1364849|RXNORM|BOS TAURUS INTESTINAL MUCOSA PREPARATION|BOVINE INTESTINAL MUCOSA PREPARATION
C3864824|T121|1597373|RXNORM|PARITAPREVIR|PARITAPREVIR
C2928880|T121|1007967|RXNORM|METHIONINE / SILYMARIN|METHIONINE / SILYMARIN
C3282848|T109|1314265|RXNORM|ARABIDOPSIS THALIANA EXTRACT|ARABIDOPSIS THALIANA EXTRACT
C2928873|T121|1007960|RXNORM|BENDROFLUMETHIAZIDE / RESERPINE|BENDROFLUMETHIAZIDE / RESERPINE
C0014757|T123|1369563|RXNORM|ERYTHRITOL|ERYTHRITOL
C3535663|T109|1369565|RXNORM|THYMUS MASTICHINA FLOWERING TOP OIL|THYMUS MASTICHINA FLOWERING TOP OIL
C3535664|T121|1369564|RXNORM|PHYSALIS ALKEKENGI CALYX EXTRACT|PHYSALIS ALKEKENGI CALYX EXTRACT
C0137904|T122|1546437|RXNORM|POLYSTYRENE SULFONATE|POLYSTYRENE SULFONATE
C2928874|T121|1007961|RXNORM|NORFENEFRINE / PENTYLENETETRAZOLE|NORFENEFRINE / PENTYLENETETRAZOLE
C2928875|T121|1007962|RXNORM|ARGININE / GINSENG PREPARATION|ARGININE / GINSENG PREPARATION
C2928876|T121|1007963|RXNORM|FOLIC ACID / POTASSIUM GLUCONATE|FOLIC ACID / POTASSIUM GLUCONATE
C0145942|T121|57230|RXNORM|TILUDRONATE|TILUDRONATE
C0301387|T121|89795|RXNORM|XANTHINOL|XANTHINOL
C3848700|T121|1546458|RXNORM|PICOSULFURATE|PICOSULFURATE
C2193955|T121|823181|RXNORM|BROMPHENIRAMINE / CODEINE|BROMPHENIRAMINE / CODEINE
C0359010|T121|106955|RXNORM|HYDROCORTISONE / PRAMOXINE|HYDROCORTISONE / PRAMOXINE
C0359010|T121|106955|RXNORM|HYDROCORTISONE / PRAMOXINE|HYDROCORTISONE / PRAMOXINE
C0359012|T121|106957|RXNORM|CROTAMITON / HYDROCORTISONE|CROTAMITON / HYDROCORTISONE
C0305070|T121|91613|RXNORM|SQUILL EXTRACT|SQUILL EXTRACT
C0770578|T197|235496|RXNORM|SODIUM PHOSPHATE, MONOBASIC|SODIUM PHOSPHATE, MONOBASIC
C0017963|T125|1427201|RXNORM|GLYCOPROTEIN HORMONES, ALPHA SUBUNIT|GLYCOPROTEIN HORMONES, ALPHA SUBUNIT
C1615665|T126|578350|RXNORM|HYALURONIDASE, BOVINE|HYALURONIDASE, BOVINE
C3486622|T121|1313319|RXNORM|AVENS EXTRACT|AVENS EXTRACT
C0073372|T195|35617|RXNORM|RIFAPENTINE|RIFAPENTINE
C0073374|T121|35619|RXNORM|RIFAXIMIN|RIFAXIMIN
C3488140|T197|1313315|RXNORM|ARSENIC TRIBROMIDE|ARSENIC TRIBROMIDE
C2939742|T129|1013944|RXNORM|WATER OAK POLLEN EXTRACT|QUERCUS NIGRA POLLEN EXTRACT
C3486627|T121|1313312|RXNORM|ANGUILLA ROSTRATA BLOOD SERUM|ANGUILLA ROSTRATA BLOOD SERUM
C0997758|T204|1313311|RXNORM|AMOEBA PROTEUS|AMOEBA PROTEUS
C3488947|T196|1313310|RXNORM|AMMONIUM ION|AMMONIUM CATION
C2728176|T129|1011049|RXNORM|CHICKPEA ALLERGENIC EXTRACT|CHICKPEA ALLERGENIC EXTRACT
C2928959|T121|1008048|RXNORM|ERGOLOID MESYLATES, USP / VITAMIN B6|ERGOLOID MESYLATES, USP / VITAMIN B6
C2928960|T121|1008049|RXNORM|PENICILLIN G BENZATHINE / PENICILLIN G SODIUM|PENICILLIN G BENZATHINE / PENICILLIN G SODIUM
C2928953|T121|1008042|RXNORM|CHOLECALCIFEROL / CHROMIUM PICOLINATE|CHOLECALCIFEROL / CHROMIUM PICOLINATE
C2928954|T121|1008043|RXNORM|CONIVAPTAN / GLUCOSE|CONIVAPTAN / GLUCOSE
C2928951|T121|1008040|RXNORM|BENZOCAINE / DEXTROMETHORPHAN / GLYCERIN|BENZOCAINE / DEXTROMETHORPHAN / GLYCERIN
C2928957|T121|1008046|RXNORM|CINNARIZINE / ERGOLOID MESYLATES, USP|CINNARIZINE / ERGOLOID MESYLATES, USP
C2928958|T121|1008047|RXNORM|METHYLSULFONYLMETHANE / MOLYBDENUM|METHYLSULFONYLMETHANE / MOLYBDENUM
C2928955|T121|1008044|RXNORM|BENZOCAINE / COMPOUND BENZOIN TINCTURE (USP)|BENZOCAINE / COMPOUND BENZOIN TINCTURE (USP)
C2948480|T121|1044247|RXNORM|MENTHOL / SODIUM CHLORIDE|MENTHOL / SODIUM CHLORIDE
C0012091|T121|3355|RXNORM|DICLOFENAC|DICLOFENAC
C0012091|T121|3355|RXNORM|DICLOFENAC|DICLOFENAC
C0012091|T121|3355|RXNORM|DICLOFENAC|DICLOFENAC
C1684371|T121|1307101|RXNORM|NEOPENTYL GLY DCAPRYL-DCAPRATE|NEOPENTYL GLY DCAPRYL-DCAPRATE
C3268107|T109|1307100|RXNORM|NEOPENTYL GLYCOL DICAPRYLATE-DICAPRATE|NEOPENTYL GLYCOL DICAPRYLATE-DICAPRATE
C0123677|T125|51428|RXNORM|INSULIN, ASPART, HUMAN|INSULIN, ASPART, HUMAN
C3667869|T122|1440228|RXNORM|HYDROGENATED METHYL ABIETATE|HYDROGENATED METHYL ABIETATE
C0070166|T121|32968|RXNORM|CLOPIDOGREL|CLOPIDOGREL
C3667868|T121|1440226|RXNORM|FICUS CARICA LEAF EXTRACT|FICUS CARICA LEAF EXTRACT
C0043456|T123|1440227|RXNORM|ZEATIN|ZEATIN
C3667866|T121|1440224|RXNORM|BOSWELLIA SACRA WHOLE EXTRACT|BOSWELLIA SACRA WHOLE EXTRACT
C3667867|T121|1440225|RXNORM|CORN COB EXTRACT|CORN COB EXTRACT
C0053284|T121|19041|RXNORM|BENZQUINAMIDE|BENZQUINAMIDE
C3855129|T121|1547458|RXNORM|CALCIUM CHLORIDE / MAGNESIUM CHLORIDE / POTASSIUM ACETATE / SODIUM ACETATE / SODIUM CHLORIDE|CALCIUM CHLORIDE / MAGNESIUM CHLORIDE / POTASSIUM ACETATE / SODIUM ACETATE / SODIUM CHLORIDE
C2700227|T130|1546432|RXNORM|GADOPENTETATE|GADOPENTETATE
C0063829|T130|27793|RXNORM|IOXILAN|IOXILAN
C0600692|T121|155164|RXNORM|ETHOSUXIMIDE / QUINACRINE|ETHOSUXIMIDE / QUINACRINE
C0717936|T121|214721|RXNORM|NALOXONE / PENTAZOCINE|NALOXONE / PENTAZOCINE
C3256855|T109|1309439|RXNORM|LEONTOPODIUM ALPINUM FLOWERING TOP EXTRACT|LEONTOPODIUM ALPINUM FLOWERING TOP EXTRACT
C3256854|T109|1309438|RXNORM|LEONTOPODIUM ALPINUM FLOWER EXTRACT|LEONTOPODIUM ALPINUM FLOWER EXTRACT
C0018165|T195|5011|RXNORM|GRAMICIDIN|GRAMICIDIN
C3256779|T109|1309435|RXNORM|LAPSANA COMMUNIS FLOWERING TOP EXTRACT|LAPSANA COMMUNIS FLOWERING TOP EXTRACT
C3256778|T109|1309434|RXNORM|LAMIUM ALBUM FLOWER EXTRACT|LAMIUM ALBUM FLOWER EXTRACT
C3256851|T109|1309437|RXNORM|LAVANDULA STOECHAS FLOWERING TOP EXTRACT|LAVANDULA STOECHAS FLOWERING TOP EXTRACT
C3256783|T109|1309436|RXNORM|LATHYRUS ODORATUS FLOWER EXTRACT|LATHYRUS ODORATUS FLOWER EXTRACT
C0718704|T121|215451|RXNORM|ASPIRIN / OXYCODONE HYDROCHLORIDE / OXYCODONE TEREPHTHALATE|ASPIRIN / OXYCODONE HYDROCHLORIDE / OXYCODONE TEREPHTHALATE
C0039267|T197|10323|RXNORM|TALC|TALC
C0039267|T197|10323|RXNORM|TALC|TALC
C3256417|T109|1309433|RXNORM|IMPERATA CYLINDRICA ROOT EXTRACT|IMPERATA CYLINDRICA ROOT EXTRACT
C3256416|T109|1309432|RXNORM|ILEX PUBESCENS ROOT EXTRACT|ILEX PUBESCENS ROOT EXTRACT
C0531104|T121|847728|RXNORM|LUMEFANTRINE|LUMEFANTRINE
C0039266|T195|10322|RXNORM|TALAMPICILLIN|TALAMPICILLIN
C2194270|T121|812750|RXNORM|ETHINYL ESTRADIOL / ETHISTERONE|ETHINYL ESTRADIOL / ETHISTERONE
C3848524|T121|1546433|RXNORM|MONOMETHYL FUMARATE|MONOMETHYL FUMARATE
C0036006|T123|9506|RXNORM|S-ADENOSYLMETHIONINE SULFATE TOSYLATE|S-ADENOSYLMETHIONINE SULFATE TOSYLATE
C2146455|T121|812759|RXNORM|SULFAMOXOLE / TRIMETHOPRIM|SULFAMOXOLE / TRIMETHOPRIM
C0039286|T121|10324|RXNORM|TAMOXIFEN|TAMOXIFEN
C0537894|T121|140108|RXNORM|CASPOFUNGIN|CASPOFUNGIN
C0063131|T122|27244|RXNORM|HYDROXYETHYL CELLULOSE|HYDROXYETHYL CELLULOSE
C1110619|T109|324030|RXNORM|PAPAYA PREPARATION|PAPAYA PREPARATION
C3535908|T122|1370196|RXNORM|C18 OLEFIN SULFONATE|C18 OLEFIN SULFONATE
C3535639|T121|1370197|RXNORM|SORGHUM BICOLOR WHOLE EXTRACT|SORGHUM BICOLOR WHOLE EXTRACT
C3535641|T121|1370194|RXNORM|SALVIA OFFICINALIS FLOWERING TOP EXTRACT|SALVIA OFFICINALIS FLOWERING TOP EXTRACT
C1962523|T121|729455|RXNORM|AMLODIPINE / VALSARTAN|AMLODIPINE / VALSARTAN
C3535642|T121|1370193|RXNORM|PROPYLENE GLYCOL 1,2-DISTEARATE|PROPYLENE GLYCOL 1,2-DISTEARATE
C3535644|T121|1370191|RXNORM|ACACIA ANGUSTISSIMA BARK EXTRACT|ACACIA ANGUSTISSIMA BARK EXTRACT
C1873975|T121|689767|RXNORM|ACETAMINOPHEN / CINNAMEDRINE / PAMABROM|ACETAMINOPHEN / CINNAMEDRINE / PAMABROM
C1873973|T121|689764|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / SALICYLAMIDE|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE / SALICYLAMIDE
C1873974|T121|689765|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / CHLORPHENIRAMINE / PSEUDOEPHEDRINE
C1873971|T121|689762|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE
C3531463|T109|1366990|RXNORM|GELATIN HYDROLYSATE (PORCINE SKIN, MW 3000)|GELATIN HYDROLYSATE (PORCINE SKIN, MW 3000)
C3531465|T109|1366993|RXNORM|PEG:PPG-4-12:DIMETHICONE|PEG:PPG-4-12:DIMETHICONE
C0039294|T121|10328|RXNORM|TANNIC ACID|TANNIC ACID
C0717787|T121|214582|RXNORM|GLATIRAMER|GLATIRAMER
C3531469|T129|1366998|RXNORM|INFLUENZA B VIRUS ANTIGEN, HONG KONG 330-2001|INFLUENZA B VIRUS ANTIGEN, HONG KONG 330-2001
C1873976|T121|689769|RXNORM|ACETAMINOPHEN / CODEINE / GUAIFENESIN / PHENYLPROPANOLAMINE|ACETAMINOPHEN / CODEINE / GUAIFENESIN / PHENYLPROPANOLAMINE
C0017817|T123|4890|RXNORM|GLUTATHIONE|GLUTATHIONE
C1110620|T121|324031|RXNORM|CARICA PAPAYA PREPARATION|CARICA PAPAYA PREPARATION
C1122962|T121|328134|RXNORM|GEFITINIB|GEFITINIB
C0004969|T121|1367|RXNORM|BETAMETHASONE / CLOTRIMAZOLE / GENTAMICIN SULFATE (USP)|BENCYCLANE
C2928279|T121|1007357|RXNORM|PRAMOXINE / ZINC ACETATE|PRAMOXINE / ZINC ACETATE
C1874979|T121|687306|RXNORM|DEXTRAN 70 / HYPROMELLOSE|DEXTRAN 70 / HYPROMELLOSE
C1302082|T121|392531|RXNORM|ERYTHROMYCIN / ZINC ACETATE|ERYTHROMYCIN / ZINC ACETATE
C1827640|T121|687304|RXNORM|DEXAMETHASONE / TRAMAZOLINE|DEXAMETHASONE / TRAMAZOLINE
C2927811|T121|1006887|RXNORM|ACETAMINOPHEN / DOXYLAMINE / PHENYLEPHRINE|ACETAMINOPHEN / DOXYLAMINE / PHENYLEPHRINE
C1302086|T121|392534|RXNORM|BUMETANIDE / POTASSIUM|BUMETANIDE / POTASSIUM
C1695970|T125|631657|RXNORM|INSULIN HUMAN, RDNA ORIGIN|INSULIN HUMAN, RDNA ORIGIN
C3643659|T121|1422070|RXNORM|BENZALKONIUM / CHLORHEXIDINE / N-ALKYL ETHYLBENZYL DIMETHYL AMMONIUM (C12-C14)|BENZALKONIUM / CHLORHEXIDINE / N-ALKYL ETHYLBENZYL DIMETHYL AMMONIUM (C12-C14)
C0028070|T121|7419|RXNORM|NIFURATEL|NIFURATEL
C3473248|T121|1298466|RXNORM|BENZYL ALCOHOL / CALAMINE / DIPHENHYDRAMINE|BENZYL ALCOHOL / CALAMINE / DIPHENHYDRAMINE
C2928278|T121|1007356|RXNORM|ASCORBIC ACID / BROMELAINS|ASCORBIC ACID / BROMELAINS
C2918009|T121|994202|RXNORM|ESOMEPRAZOLE / NAPROXEN|ESOMEPRAZOLE / NAPROXEN
C2936902|T121|994203|RXNORM|DIENOGEST / ESTRADIOL|DIENOGEST / ESTRADIOL
C0301513|T129|597392|RXNORM|HUMAN VACCINIA IMMUNE GLOBULIN|HUMAN VACCINIA IMMUNE GLOBULIN
C3834053|T121|1543293|RXNORM|ASPLENIUM SCOLOPENDRIUM WHOLE EXTRACT|ASPLENIUM SCOLOPENDRIUM WHOLE EXTRACT
C2929854|T121|1008958|RXNORM|HYDROCORTISONE / POTASSIUM OXYQUINOLONE|HYDROCORTISONE / POTASSIUM OXYQUINOLONE
C0030557|T121|7930|RXNORM|PARGYLINE|PARGYLINE
C0030576|T195|7934|RXNORM|PAROMOMYCIN|PAROMOMYCIN
C0027556|T121|7285|RXNORM|NEFOPAM|NEFOPAM
C2929847|T121|1008950|RXNORM|CITRIC ACID / STEVIOSIDE / TARTARIC ACID|CITRIC ACID / STEVIOSIDE / TARTARIC ACID
C2929848|T121|1008951|RXNORM|BENZOCAINE / CETYLPYRIDINIUM / SULFACHRYSOIDINE|BENZOCAINE / CETYLPYRIDINIUM / SULFACHRYSOIDINE
C2929849|T121|1008952|RXNORM|BISMUTH HYDROXIDE / PECTIN|BISMUTH HYDROXIDE / PECTIN
C0027575|T007|7288|RXNORM|NEISSERIA MENINGITIDIS|NEISSERIA MENINGITIDIS
C2929851|T121|1008954|RXNORM|CODEINE / ERYSIMUM PREPARATION|CODEINE / ERYSIMUM PREPARATION
C2929852|T121|1008955|RXNORM|GUAIACOLSULFONATE / HYDROCODONE / PSEUDOEPHEDRINE|GUAIACOLSULFONATE / HYDROCODONE / PSEUDOEPHEDRINE
C2929853|T121|1008956|RXNORM|ASCORBIC ACID / UBIQUINOL|ASCORBIC ACID / UBIQUINOL
C3834052|T121|1543294|RXNORM|ROSA DAMASCENA WHOLE EXTRACT|ROSA DAMASCENA WHOLE EXTRACT
C1699911|T121|617777|RXNORM|OMEPRAZOLE / SODIUM BICARBONATE|OMEPRAZOLE / SODIUM BICARBONATE
C0055775|T121|21149|RXNORM|CIPROFIBRATE|CIPROFIBRATE
C3538032|T121|1371903|RXNORM|BOS TAURUS PLACENTA PREPARATION|BOS TAURUS PLACENTA PREPARATION
C0030815|T121|7974|RXNORM|PENFLURIDOL|PENFLURIDOL
C0937950|T121|283838|RXNORM|DARBEPOETIN ALFA|DARBEPOETIN ALFA
C3668731|T121|1441322|RXNORM|IRESINE CALEA EXTRACT|IRESINE CALEA EXTRACT
C0075429|T121|37255|RXNORM|SUCCINIC ACID|SUCCINIC ACID
C1874980|T121|690474|RXNORM|DEXTRAN 70 / SODIUM CHLORIDE|DEXTRAN 70 / SODIUM CHLORIDE
C1874985|T121|690479|RXNORM|DEXTROMETHORPHAN / DYPHYLLINE / PSEUDOEPHEDRINE|DEXTROMETHORPHAN / DYPHYLLINE / PSEUDOEPHEDRINE
C0771782|T197|236502|RXNORM|TRIBASIC POTASSIUM PHOSPHATE|TRIBASIC POTASSIUM PHOSPHATE
C3651706|T121|1431310|RXNORM|OPUNTIA TUNA FLOWERING TOP EXTRACT|OPUNTIA TUNA FLOWERING TOP EXTRACT
C3530899|T121|1365707|RXNORM|PANAX NOTOGINSENG ROOT EXTRACT|PANAX NOTOGINSENG ROOT EXTRACT
C3530898|T121|1365706|RXNORM|LIGUSTICUM WALLICHII ROOT EXTRACT|LIGUSTICUM WALLICHII ROOT EXTRACT
C0138037|T197|55018|RXNORM|DIBASIC POTASSIUM PHOSPHATE|DIBASIC POTASSIUM PHOSPHATE
C3813123|T121|1544392|RXNORM|EPIGAEA REPENS EXTRACT|EPIGAEA REPENS EXTRACT
C3256540|T121|1313238|RXNORM|ISOAMYL LAURATE|ISOAMYL LAURATE
C0012319|T127|3429|RXNORM|DIHYDROTACHYSTEROL|DIHYDROTACHYSTEROL
C2222740|T121|814380|RXNORM|BIOALLETHRIN / PIPERONYL BUTOXIDE|BIOALLETHRIN / PIPERONYL BUTOXIDE
C0144576|T121|56946|RXNORM|PACLITAXEL|PACLITAXEL
C2949423|T121|1046533|RXNORM|DEXPANTHENOL / LEVOMENTHOL / SALICYLIC ACID|DEXPANTHENOL / LEVOMENTHOL / SALICYLIC ACID
C0012306|T121|3423|RXNORM|HYDROMORPHONE|HYDROMORPHONE
C2741435|T129|901191|RXNORM|CONCORD GRAPE ALLERGENIC EXTRACT|VITIS LABRUSCA ALLERGENIC EXTRACT
C2741438|T129|901195|RXNORM|SAFFLOWER SEED ALLERGENIC EXTRACT|SAFFLOWER SEED ALLERGENIC EXTRACT
C3256235|T130|1425505|RXNORM|FD&C BLUE #2 HT ALUMINUM LAKE|FD&C BLUE #2 HT ALUMINUM LAKE
C0006949|T121|2002|RXNORM|CARBAMAZEPINE|CARBAMAZEPINE
C0055819|T123|21183|RXNORM|CITRIC ACID|CITRIC ACID
C0017725|T123|4850|RXNORM|GLUCOSE|GLUCOSE
C0017725|T123|4850|RXNORM|GLUCOSE|GLUCOSE
C0017725|T123|4850|RXNORM|GLUCOSE|GLUCOSE
C0017725|T123|4850|RXNORM|GLUCOSE|GLUCOSE
C2929502|T121|1008600|RXNORM|BLACK COHOSH EXTRACT / MAGNESIUM OXIDE / ST. JOHN'S WORT EXTRACT|BLACK COHOSH EXTRACT / MAGNESIUM OXIDE / ST. JOHN'S WORT EXTRACT
C2929503|T121|1008601|RXNORM|PYGEUM AFRICANUM PREPARATION / URTICA PREPARATION|PYGEUM AFRICANUM PREPARATION / URTICA PREPARATION
C2929504|T121|1008602|RXNORM|ASCORBIC ACID / ECHINACEA PURPUREA EXTRACT / ZINC GLUCONATE|ASCORBIC ACID / ECHINACEA PURPUREA EXTRACT / ZINC GLUCONATE
C2193837|T121|1008603|RXNORM|AMOXICILLIN / NYSTATIN|AMOXICILLIN / NYSTATIN
C2929505|T121|1008604|RXNORM|DANTHRON / PANTOTHENATE|DANTHRON / PANTOTHENATE
C2929506|T121|1008605|RXNORM|MAGNESIUM SULFATE / PHENOLPHTHALEIN|MAGNESIUM SULFATE / PHENOLPHTHALEIN
C2193854|T121|1008606|RXNORM|AMOXICILLIN / PIROXICAM|AMOXICILLIN / PIROXICAM
C3247775|T129|1192968|RXNORM|HYPOMYCES PERNICIOSUS EXTRACT|HYPOMYCES PERNICIOSUS EXTRACT
C2929508|T121|1008608|RXNORM|ARGININE / GINKGO BILOBA EXTRACT / YOHIMBINE|ARGININE / GINKGO BILOBA EXTRACT / YOHIMBINE
C2929509|T121|1008609|RXNORM|NAPHAZOLINE / POLYETHYLENE GLYCOLS|NAPHAZOLINE / POLYETHYLENE GLYCOLS
C0003380|T196|1311407|RXNORM|ANTIMONY|ANTIMONY
C3530900|T121|1365708|RXNORM|ZANTHOXYLUM NITIDUM ROOT EXTRACT|ZANTHOXYLUM NITIDUM ROOT EXTRACT
C3645142|T121|1426693|RXNORM|CHONDROITIN SULFATES / GLUCOSAMINE / HYALURONATE / METHYLSULFONYLMETHANE|CHONDROITIN SULFATES / GLUCOSAMINE / HYALURONATE / METHYLSULFONYLMETHANE
C3152989|T129|1311406|RXNORM|SORGHUM BICOLOR POLLEN EXTRACT|SORGHUM BICOLOR SUBSP. BICOLOR POLLEN EXTRACT
C1519991|T121|1304991|RXNORM|VINCRISTINE LIPOSOME|VINCRISTINE LIPOSOME
C0057380|T109|1313232|RXNORM|DENATONIUM BENZOATE|DENATONIUM BENZOATE
C0026088|T121|6964|RXNORM|MIFEPRISTONE|MIFEPRISTONE
C0026088|T121|6964|RXNORM|MIFEPRISTONE|MIFEPRISTONE
C3538036|T109|1371908|RXNORM|ANGELICA ACUTILOBA ROOT OIL|ANGELICA ACUTILOBA ROOT OIL
C3267476|T168|1313233|RXNORM|PEAR JUICE|PEAR JUICE
C3814772|T121|1546438|RXNORM|GLYCOPYRRONIUM|GLYCOPYRRONIUM
C0026534|T121|1368900|RXNORM|MORANTEL|MORANTEL
C1314952|T121|400674|RXNORM|DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE|DEXBROMPHENIRAMINE / PSEUDOEPHEDRINE
C1572729|T121|1368902|RXNORM|ELEUTHERO PREPARATION|ELEUTHERO PREPARATION
C3487961|T197|1368903|RXNORM|MERCURIC CATION|MERCURIC CATION
C3535669|T121|1368905|RXNORM|C12-13 PARETH-23|C12-13 PARETH-23
C3538033|T121|1371904|RXNORM|BOS TAURUS VEIN PREPARATION|BOS TAURUS VEIN PREPARATION
C3535668|T121|1368907|RXNORM|C12-13 PARETH-3|C12-13 PARETH-3
C0040162|T125|10580|RXNORM|THYROTROPIN-RELEASING HORMONE|THYROTROPIN-RELEASING HORMONE
C0040165|T125|10582|RXNORM|THYROXINE|LEVOTHYROXINE
C3486569|T121|1310039|RXNORM|TRIFOLIUM PRATENSE FLOWER EXTRACT|TRIFOLIUM PRATENSE FLOWER EXTRACT
C3474081|T121|1310037|RXNORM|PRUNUS SERRULATA FLOWER EXTRACT|PRUNUS SERRULATA FLOWER EXTRACT
C0040180|T121|10588|RXNORM|TIAPRIDE|TIAPRIDE
C3486557|T121|1310035|RXNORM|SOLANUM DULCAMARA STEM EXTRACT|SOLANUM DULCAMARA STEM EXTRACT
C3474076|T121|1310034|RXNORM|MAGNOLIA LILIIFLORA FLOWER EXTRACT|MAGNOLIA LILIIFLORA FLOWER EXTRACT
C3484423|T121|1310033|RXNORM|PIMPINELLA SAXIFRAGA ROOT EXTRACT|PIMPINELLA SAXIFRAGA ROOT EXTRACT
C3486550|T121|1310032|RXNORM|TURNERA DIFFUSA LEAFY TWIG EXTRACT|TURNERA DIFFUSA LEAFY TWIG EXTRACT
C3484408|T121|1310031|RXNORM|NERIUM OLEANDER LEAF EXTRACT|NERIUM OLEANDER LEAF EXTRACT
C3473993|T109|1310030|RXNORM|SPANISH THYME OIL|SPANISH THYME OIL
C2684757|T129|851949|RXNORM|CAT SKIN EXTRACT|FELIS CATUS SKIN EXTRACT
C3267654|T121|1306885|RXNORM|MOMORDICA CHARANTIA FRUIT EXTRACT|MOMORDICA CHARANTIA FRUIT EXTRACT
C3486833|T121|1311258|RXNORM|SUS SCROFA SYMPATHETIC NERVE PREPARATION|PORCINE SYMPATHETIC NERVE PREPARATION
C0070525|T121|33253|RXNORM|PHENACEMIDE|PHENACEMIDE
C0071324|T121|33926|RXNORM|POLDINE|POLDINE
C3496030|T121|1311254|RXNORM|SUS SCROFA MESENCHYME PREPARATION|PORCINE MESENCHYME PREPARATION
C3496031|T121|1311255|RXNORM|SUS SCROFA RED BLOOD CELL PREPARATION|PORCINE ERYTHROCYTE PREPARATION
C3496032|T121|1311256|RXNORM|SUS SCROFA SOLAR PLEXUS PREPARATION|PORCINE SOLAR PLEXUS PREPARATION
C0360665|T121|108190|RXNORM|GLUCOSE / SODIUM CHLORIDE|GLUCOSE / SODIUM CHLORIDE
C3496027|T121|1311250|RXNORM|SUS SCROFA HIP JOINT PREPARATION|PORCINE HIP JOINT PREPARATION
C3496028|T121|1311251|RXNORM|SUS SCROFA HIPPOCAMPUS PREPARATION|PORCINE HIPPOCAMPUS PREPARATION
C3496029|T121|1311252|RXNORM|SUS SCROFA JOINT CAPSULE PREPARATION|PORCINE JOINT CAPSULE PREPARATION
C3486802|T121|1311253|RXNORM|SUS SCROFA LYMPH PREPARATION|PORCINE LYMPH PREPARATION
C3282460|T121|1306886|RXNORM|N-CYCLOHEXYL-2-BENZOTHIAZOSULFENAMIDE|N-CYCLOHEXYL-2-BENZOTHIAZOSULFENAMIDE
C0075932|T130|37665|RXNORM|TECHNETIUM TC 99M DISOFENIN|TECHNETIUM (99MTC) DISOFENIN
C0083381|T121|41493|RXNORM|MELOXICAM|MELOXICAM
C2980840|T129|1306881|RXNORM|ABSIDIA CAPILLATA ALLERGENIC EXTRACT|ABSIDIA CAPILLATA ALLERGENIC EXTRACT
C0101700|T121|45938|RXNORM|ADRAFINIL|ADRAFINIL
C3486617|T121|1318231|RXNORM|CHIMAPHILA UMBELLATA EXTRACT|CHIMAPHILA UMBELLATA EXTRACT
C0063340|T121|27403|RXNORM|IFENPRODIL|IFENPRODIL
C3486662|T121|1318233|RXNORM|VINCA MINOR EXTRACT|VINCA MINOR EXTRACT
C0041090|T121|10847|RXNORM|TRIPELENNAMINE|TRIPELENNAMINE
C0041090|T121|10847|RXNORM|TRIPELENNAMINE|TRIPELENNAMINE
C3488032|T121|1318235|RXNORM|COMFREY LEAF EXTRACT|COMFREY LEAF EXTRACT
C3486838|T121|1318234|RXNORM|XEROPHYLLUM ASPHODELOIDES EXTRACT|XEROPHYLLUM ASPHODELOIDES EXTRACT
C3488986|T121|1318237|RXNORM|XANTHIUM EXTRACT|XANTHIUM EXTRACT
C3488946|T121|1318236|RXNORM|ACHYROCLINE SATUREIOIDES EXTRACT|ACHYROCLINE SATUREIOIDES EXTRACT
C0982208|T121|314674|RXNORM|HYOSCYAMUS EXTRACT|HYOSCYAMUS EXTRACT
C3486723|T121|1310259|RXNORM|CRATAEGUS LAEVIGATA FRUIT|CRATAEGUS LAEVIGATA FRUIT
C3495983|T121|1310258|RXNORM|BOS TAURUS HIP JOINT PREPARATION|BOVINE HIP JOINT PREPARATION
C2727910|T129|889646|RXNORM|RED SNAPPER ALLERGENIC EXTRACT|RED SNAPPER ALLERGENIC EXTRACT
C3256127|T121|1310253|RXNORM|BOS TAURUS COLOSTRUM PREPARATION|BOVINE COLOSTRUM PREPARATION
C0005139|T196|1310252|RXNORM|BERYLLIUM|BERYLLIUM
C2962946|T121|1087405|RXNORM|ASCORBIC ACID / BIOTIN / COPPER SULFATE / DOCUSATE / FOLIC ACID / IRON CARBONYL / VITAMIN B 12 / VITAMIN E|ASCORBIC ACID / BIOTIN / COPPER SULFATE / DOCUSATE / FOLIC ACID / IRON CARBONYL / VITAMIN B 12 / VITAMIN E
C3486287|T121|1310256|RXNORM|BOS TAURUS GALLBLADDER PREPARATION|BOVINE GALLBLADDER PREPARATION
C3495982|T121|1310255|RXNORM|BOS TAURUS FRONTAL LOBE PREPARATION|BOVINE FRONTAL LOBE PREPARATION
C3486836|T121|1311078|RXNORM|SUS SCROFA PINEAL GLAND PREPARATION|PORCINE PINEAL GLAND PREPARATION
C3484597|T121|1311079|RXNORM|SANGUINARIA CANADENSIS EXTRACT|SANGUINARIA CANADENSIS EXTRACT
C3555479|T168|1420960|RXNORM|COCONUT JUICE|COCONUT JUICE
C0023031|T196|1311070|RXNORM|LANTHANUM|LANTHANUM
C3486585|T121|1311071|RXNORM|PORK LIVER PREPARATION|PORK LIVER PREPARATION
C0873186|T197|1311072|RXNORM|BARIUM IODIDE|BARIUM IODIDE
C3485062|T121|1311073|RXNORM|CAIRINA MOSHCATA HEART-LIVER PREPARATION|CAIRINA MOSHCATA HEART-LIVER PREPARATION
C3488333|T197|1311076|RXNORM|RADIUM BROMIDE|RADIUM BROMIDE
C3484593|T121|1311077|RXNORM|CLAVICEPS PURPUREA SCLEROTIUM|CLAVICEPS PURPUREA SCLEROTIUM
C2928635|T121|1007719|RXNORM|FLUOXYMESTERONE / GINSENOSIDE / VITAMIN E|FLUOXYMESTERONE / GINSENOSIDE / VITAMIN E
C2928634|T121|1007718|RXNORM|CHLORAMPHENICOL / NEOMYCIN|CHLORAMPHENICOL / NEOMYCIN
C2928633|T121|1007717|RXNORM|DIPERODON / HYDROCORTISONE|DIPERODON / HYDROCORTISONE
C2928632|T121|1007716|RXNORM|ACETAMINOPHEN / THIAMINE|ACETAMINOPHEN / THIAMINE
C2928631|T121|1007715|RXNORM|ESTRADIOL / ESTRIOL|ESTRADIOL / ESTRIOL
C2928630|T121|1007714|RXNORM|IODINE / POTASSIUM GLUCONATE|IODINE / POTASSIUM GLUCONATE
C2928629|T121|1007713|RXNORM|DIPHENHYDRAMINE / OXELADIN / SALICYLAMIDE|DIPHENHYDRAMINE / OXELADIN / SALICYLAMIDE
C2928628|T121|1007712|RXNORM|MEBENDAZOLE / NICLOSAMIDE / TINIDAZOLE|MEBENDAZOLE / NICLOSAMIDE / TINIDAZOLE
C2928627|T121|1007711|RXNORM|ISOSORBIDE DINITRATE / VERAPAMIL|ISOSORBIDE DINITRATE / VERAPAMIL
C2928626|T121|1007710|RXNORM|CALCIUM CARBONATE / MAGNESIUM CARBONATE / SIMETHICONE|CALCIUM CARBONATE / MAGNESIUM CARBONATE / SIMETHICONE
C1579345|T121|591533|RXNORM|SULFADIAZINE / TRIMETHOPRIM|SULFADIAZINE / TRIMETHOPRIM
C3256916|T109|1309999|RXNORM|GANODERMA LUCIDUM STEM EXTRACT|GANODERMA LUCIDUM STEM EXTRACT
C3256105|T109|1368890|RXNORM|HYPROMELLOSE PHTHALATE (24% PHTHALATE, 55 CST)|HYPROMELLOSE PHTHALATE (24% PHTHALATE, 55 CST)
C1874221|T121|691318|RXNORM|AMOBARBITAL / EPHEDRINE|AMOBARBITAL / EPHEDRINE
C0876769|T197|262150|RXNORM|IRON CARBONYL|IRON CARBONYL
C3465267|T121|1309993|RXNORM|ULMUS DAVIDIANA ROOT EXTRACT|ULMUS DAVIDIANA ROOT EXTRACT
C3486688|T121|1309990|RXNORM|HELLEBORUS NIGER ROOT EXTRACT|HELLEBORUS NIGER ROOT EXTRACT
C3488655|T121|1309991|RXNORM|THUJA OCCIDENTALIS ROOT EXTRACT|THUJA OCCIDENTALIS ROOT EXTRACT
C3465271|T121|1309996|RXNORM|FRAXINUS EXCELSIOR BARK EXTRACT|FRAXINUS EXCELSIOR BARK EXTRACT
C3256899|T109|1309997|RXNORM|CEDRELOPSIS GREVEI BARK EXTRACT|CEDRELOPSIS GREVEI BARK EXTRACT
C3488987|T121|1309994|RXNORM|CARPINUS BETULUS FLOWER EXTRACT|CARPINUS BETULUS FLOWER EXTRACT
C0055559|T109|1362887|RXNORM|CHOLESTERYL NONANOATE|CHOLESTERYL NONANOATE
C0055465|T195|1362886|RXNORM|CHLOROZOTOCIN|CHLOROZOTOCIN
C0053183|T109|1362885|RXNORM|BENZIMIDAZOLE|BENZIMIDAZOLE
C0051719|T197|1362884|RXNORM|AMMONIUM HYDROXIDE|AMMONIUM HYDROXIDE
C0051704|T130|1362883|RXNORM|AMMONIUM ACETATE|AMMONIUM ACETATE
C0051348|T121|1362882|RXNORM|ALPHA-CYCLODEXTRIN|ALPHA-CYCLODEXTRIN
C0045801|T121|1362881|RXNORM|2-ACETYLTRIBUTYLCITRATE|2-ACETYLTRIBUTYLCITRATE
C0044041|T121|1362880|RXNORM|1,5-PENTANEDIOL|PENTYLENE GLYCOL
C0065967|T125|29523|RXNORM|MEPREDNISONE|MEPREDNISONE
C0612777|T121|1541750|RXNORM|GLYCERAN POLYRICINOLEIC ACID ESTER|GLYCERAN POLYRICINOLEIC ACID ESTER
C0055762|T109|1362889|RXNORM|CINNAMYL ALCOHOL|CINNAMYL ALCOHOL
C0055661|T121|1362888|RXNORM|CHRYSIN|CHRYSIN
C3709490|T121|1487532|RXNORM|SUNFLOWER LECITHIN|SUNFLOWER LECITHIN
C0062636|T197|1487531|RXNORM|HEXAMETAPHOSPHATE|HEXAMETAPHOSPHATE
C0001962|T121|448|RXNORM|ETHANOL|ETHANOL
C0001962|T121|448|RXNORM|ETHANOL|ETHANOL
C0001962|T121|448|RXNORM|ETHANOL|ETHANOL
C0146894|T197|1487534|RXNORM|TRIPHOSPHATE|TRIPHOSPHATE
C2003424|T121|1040028|RXNORM|LURASIDONE|LURASIDONE
C3666444|T121|1436961|RXNORM|PPG-3 BENZYL ETHER ETHYLHEXANOATE|PPG-3 BENZYL ETHER ETHYLHEXANOATE
C0004754|T197|1331|RXNORM|BARIUM SULFATE|BARIUM SULFATE
C2142877|T121|818931|RXNORM|DEXTROMETHORPHAN / PSEUDOEPHEDRINE / TRIPROLIDINE|DEXTROMETHORPHAN / PSEUDOEPHEDRINE / TRIPROLIDINE
C1170013|T121||RXNORM|LOVASTATIN / NIACIN
C2079438|T121|814321|RXNORM|ETHAMBUTOL / ISONIAZID / RIFAMPIN|ETHAMBUTOL / ISONIAZID / RIFAMPIN
C0937645|T121|283583|RXNORM|RHUS TOXICODENDRON|RHUS TOXICODENDRON EXTRACT
C0033215|T121|8699|RXNORM|PROBUCOL|PROBUCOL
C0033209|T121|8698|RXNORM|PROBENECID|PROBENECID
C1170007|T121|352381|RXNORM|GLIPIZIDE / METFORMIN|GLIPIZIDE / METFORMIN
C3256565|T121|1307605|RXNORM|THEOBROMA GRANDIFLORUM SEED BUTTER EXTRACT|THEOBROMA GRANDIFLORUM SEED BUTTER EXTRACT
C0075246|T121|37106|RXNORM|STEVIOSIDE|STEVIOSIDE
C2726179|T129|1192992|RXNORM|MICROASCUS BREVICAULIS ALLERGENIC EXTRACT|MICROASCUS BREVICAULIS ALLERGENIC EXTRACT
C0031392|T121|8123|RXNORM|PHENELZINE|PHENELZINE
C3152855|T121|1098214|RXNORM|ETHANOL / POVIDONE-IODINE|ETHANOL / POVIDONE-IODINE
C2726184|T129|1192997|RXNORM|GLIOCLADIUM ALLERGENIC EXTRACT|MYROTHECIUM VERRUCARIA ALLERGENIC EXTRACT
C0029277|T123|7704|RXNORM|ORNITHINE|ORNITHINE
C1722449|T109|1424270|RXNORM|N-LACTOYLETHANOLAMINE|N-LACTOYLETHANOLAMINE
C0029276|T121|7703|RXNORM|ORNIPRESSIN|ORNIPRESSIN
C0029274|T121|7701|RXNORM|ORNIDAZOLE|ORNIDAZOLE
C2743583|T109|1428039|RXNORM|CALENDULOSIDE E|CALENDULOSIDE E
C1304571|T121|392938|RXNORM|BUTETHAMATE|BUTETHAMATE
C0142822|T197|992920|RXNORM|SODIUM CHLORITE|SODIUM CHLORITE
C0120726|T121|50749|RXNORM|HALOFANTRINE|HALOFANTRINE
C3666987|T121|1438114|RXNORM|BEHENAMIDOPROPYLTRIMONIUM METHOSULFATE|BEHENAMIDOPROPYLTRIMONIUM METHOSULFATE
C3256084|T121|1307851|RXNORM|PRUNUS SEROTINA BARK EXTRACT|PRUNUS SEROTINA BARK EXTRACT
C1658225|T121|581386|RXNORM|WHORTLEBERRY SUBSTANCE|WHORTLEBERRY SUBSTANCE
C0059725|T121|24484|RXNORM|ETHOHEPTAZINE|ETHOHEPTAZINE
C3535637|T197|1370299|RXNORM|FERROUS ARSENATE|FERROUS ARSENATE
C3535638|T121|1370298|RXNORM|ANTIARIS TOXICARA RESIN EXTRACT|ANTIARIS TOXICARA RESIN
C0171023|T121|61381|RXNORM|OLANZAPINE|OLANZAPINE
C3832870|T121|1539811|RXNORM|DIMETHYLMETHOXY CHROMANOL|DIMETHYLMETHOXY CHROMANOL
C3531289|T121|1366507|RXNORM|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / GUAIFENESIN / N-METHYLEPHEDRINE|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / GUAIFENESIN / N-METHYLEPHEDRINE
C1276338|T121|389103|RXNORM|EPINEPHRINE / MEPIVACAINE|EPINEPHRINE / MEPIVACAINE
C0031968|T121|8348|RXNORM|PIPOTHIAZINE|PIPOTHIAZINE
C2348901|T109|1307850|RXNORM|BULNESIA SARMIENTOI WOOD OIL|BULNESIA SARMIENTOI WOOD OIL
C0031957|T121|8340|RXNORM|PIPERAZINE|PIPERAZINE
C0031965|T121|8347|RXNORM|PIPOBROMAN|PIPOBROMAN
C1874347|T121|689489|RXNORM|ASCORBIC ACID / DOCUSATE / FERROUS FUMARATE|ASCORBIC ACID / DOCUSATE / FERROUS FUMARATE
C0057257|T121|1311089|RXNORM|DEFIBROTIDE|DEFIBROTIDE
C0752378|T121|228080|RXNORM|PIRENOXINE|PIRENOXINE
C0063075|T197|1426869|RXNORM|HYDROBROMIC ACID|HYDROBROMIC ACID
C0318253|T007|100534|RXNORM|VIBRIO CHOLERAE SEROTYPE OGAWA|VIBRIO CHOLERAE SEROTYPE OGAWA
C0318252|T007|100533|RXNORM|VIBRIO CHOLERAE SEROTYPE INABA|VIBRIO CHOLERAE SEROTYPE INABA
C0079134|T007|1534764|RXNORM|CLOSTRIDIUM DIFFICILE (BACTERIA)|CLOSTRIDIUM DIFFICILE (BACTERIA)
C1876654|T122|1364388|RXNORM|LAURAMINE OXIDE|LAURAMINE OXIDE
C3542455|T121|1435392|RXNORM|SARGASSUM FUSIFORME EXTRACT|SARGASSUM FUSIFORME EXTRACT
C0059696|T130|24457|RXNORM|ETHANOLAMINE|ETHANOLAMINE
C3858056|T121|1551285|RXNORM|CHLOPHEDIANOL / DEXBROMPHENIRAMINE|CHLOPHEDIANOL / DEXBROMPHENIRAMINE
C0059692|T121|24453|RXNORM|ETHAMIVAN|ETAMIVAN
C0717645|T121|214445|RXNORM|CODEINE / PSEUDOEPHEDRINE|CODEINE / PSEUDOEPHEDRINE
C0717644|T121|214444|RXNORM|CODEINE / PROMETHAZINE|CODEINE / PROMETHAZINE
C0717647|T121|214447|RXNORM|CODEINE / GUAIFENESIN / PHENYLPROPANOLAMINE|CODEINE / GUAIFENESIN / PHENYLPROPANOLAMINE
C0303296|T197|1544125|RXNORM|SILVER FLUORIDE|SILVER FLUORIDE
C0717643|T121|214443|RXNORM|CODEINE / IODINATED GLYCEROL|CODEINE / IODINATED GLYCEROL
C0717642|T121|214442|RXNORM|CODEINE / GUAIFENESIN|CODEINE / GUAIFENESIN
C3256056|T121|1307730|RXNORM|MATRICARIA RECUTITA FLOWERING TOP EXTRACT|MATRICARIA RECUTITA FLOWERING TOP EXTRACT
C3255854|T121|1307731|RXNORM|PAEONIA LACTIFLORA ROOT EXTRACT|PAEONIA LACTIFLORA ROOT EXTRACT
C3282453|T025|1307732|RXNORM|HUMAN CORD BLOOD HEMATOPOIETIC PROGENITOR CELL|HUMAN CORD BLOOD HEMATOPOIETIC PROGENITOR CELL
C3256211|T121|1307733|RXNORM|CUCUMBER SEED EXTRACT|CUCUMBER SEED EXTRACT
C0717649|T121|214449|RXNORM|CODEINE / PHENYLEPHRINE / PROMETHAZINE|CODEINE / PHENYLEPHRINE / PROMETHAZINE
C3256672|T121|1307735|RXNORM|CYATHULA OFFICINALIS ROOT EXTRACT|CYATHULA OFFICINALIS ROOT EXTRACT
C3256509|T121|1307736|RXNORM|BUPLEURUM CHINENSE ROOT EXTRACT|BUPLEURUM CHINENSE ROOT EXTRACT
C3256715|T121|1307737|RXNORM|POTENTILLA ERECTA ROOT EXTRACT|POTENTILLA ERECTA ROOT EXTRACT
C3665583|T121|1486391|RXNORM|BOSWELLIA SERRATA WHOLE EXTRACT|BOSWELLIA SERRATA WHOLE EXTRACT
C3486628|T121|1309830|RXNORM|APOCYNUM ANDROSAEMIFOLIUM ROOT EXTRACT|APOCYNUM ANDROSAEMIFOLIUM ROOT EXTRACT
C3268187|T121|1426862|RXNORM|ETHYLHEXYL OLEATE|ETHYLHEXYL OLEATE
C2701645|T129|852561|RXNORM|CALIFORNIA BLACK WALNUT POLLEN EXTRACT|JUGLANS CALIFORNICA POLLEN EXTRACT
C2929289|T121|1008385|RXNORM|APPLE PECTIN / GUAR GUM|APPLE PECTIN / GUAR GUM
C2929288|T121|1008384|RXNORM|ATTAPULGITE / SALICYLIC ACID / SULFUR,COLLOIDAL|ATTAPULGITE / SALICYLIC ACID / SULFUR,COLLOIDAL
C2929291|T121|1008387|RXNORM|GINSENG PREPARATION / SAW PALMETTO EXTRACT|GINSENG PREPARATION / SAW PALMETTO EXTRACT
C1874349|T121|1008386|RXNORM|ASCORBIC ACID / FERROUS SULFATE / FOLIC ACID|ASCORBIC ACID / FERROUS SULFATE / FOLIC ACID
C2929286|T121|1008381|RXNORM|CHROMIUM PICOLINATE / GAMBOGE|CHROMIUM PICOLINATE / GAMBOGE
C2929285|T121|1008380|RXNORM|GLUCOSAMINE / POTASSIUM|GLUCOSAMINE / POTASSIUM
C2929287|T121|1008383|RXNORM|BENZETHONIUM / DIPHENHYDRAMINE / ZINC ACETATE|BENZETHONIUM / DIPHENHYDRAMINE / ZINC ACETATE
C3505678|T121|1359085|RXNORM|OLETH-3|OLETH-3
C3159546|T121|1111420|RXNORM|ASPIRIN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE|ASPIRIN / CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE
C0014892|T121|4077|RXNORM|ESTAZOLAM|ESTAZOLAM
C3505679|T121|1359086|RXNORM|PALMITOYL GLYCINE|PALMITOYL GLYCINE
C2929293|T121|1008389|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / FERROUS FUMARATE / FOLIC ACID / PYRIDOXINE / TRICALCIUM PHOSPHATE|ALPHA TOCOPHEROL / ASCORBIC ACID / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / FERROUS FUMARATE / FOLIC ACID / PYRIDOXINE / TRICALCIUM PHOSPHATE
C0014479|T121|3966|RXNORM|EPHEDRINE|EPHEDRINE
C0014479|T121|3966|RXNORM|EPHEDRINE|EPHEDRINE
C0014479|T121|3966|RXNORM|EPHEDRINE|EPHEDRINE
C3535897|T121|1370583|RXNORM|DODECAHYDROXYCYCLOHEXANE|DODECAHYDROXYCYCLOHEXANE
C0034392|T127|9060|RXNORM|QUERCETIN|QUERCETIN
C2948088|T121|1310164|RXNORM|CENTELLA ASIATICA EXTRACT|HYDROCOTYLE ASIATICA EXTRACT
C1875702|T121|690169|RXNORM|PROPYLENE GLYCOL / SODIUM CHLORIDE|PROPYLENE GLYCOL / SODIUM CHLORIDE
C3487977|T121|1310166|RXNORM|PELARGONIUM SIDOIDES ROOT EXTRACT|PELARGONIUM SIDOIDES ROOT EXTRACT
C0013085|T121|3638|RXNORM|DOXEPIN|DOXEPIN
C0013085|T121|3638|RXNORM|DOXEPIN|DOXEPIN
C0013089|T195|3639|RXNORM|DOXORUBICIN|DOXORUBICIN
C3857958|T122|1551570|RXNORM|VINYLPYRROLIDONE-HEXADECENE COPOLYMER|VINYLPYRROLIDONE-HEXADECENE COPOLYMER
C0013084|T121|3637|RXNORM|DOXAPRAM|DOXAPRAM
C0013065|T121|3634|RXNORM|DOTHIEPIN|DOTHIEPIN
C0717396|T121|214208|RXNORM|ALUMINUM HYDROXIDE / MINERAL OIL|ALUMINUM HYDROXIDE / MINERAL OIL
C2702393|T129|854082|RXNORM|ASPERGILLUS NIGER VAR. NIGER EXTRACT|ASPERGILLUS NIGER VAR. NIGER EXTRACT
C0281563|T121|81782|RXNORM|SHARK CARTILAGE EXTRACT|SHARK CARTILAGE EXTRACT
C3487975|T121|1310163|RXNORM|KALMIA ANGUSTIFOLIA LEAF EXTRACT|KALMIA ANGUSTIFOLIA LEAF EXTRACT
C2006342|T121|817061|RXNORM|CARBINOXAMINE / OXELADIN|CARBINOXAMINE / OXELADIN
C2701486|T129|852302|RXNORM|COAST LIVE OAK POLLEN EXTRACT|QUERCUS AGRIFOLIA POLLEN EXTRACT
C2146612|T121|817430|RXNORM|ACETAMINOPHEN / CAFFEINE / CODEINE / MEPROBAMATE|ACETAMINOPHEN / CAFFEINE / CODEINE / MEPROBAMATE
C2701490|T129|852306|RXNORM|SILVER RAGWEED POLLEN EXTRACT|DICORIA CANESCENS POLLEN EXTRACT
C0771692|T197|236420|RXNORM|MAGNESIUM THIOSULFATE|MAGNESIUM THIOSULFATE
C3245225|T121|1190599|RXNORM|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C0303294|T121|1306066|RXNORM|SILVER CITRATE|SILVER CITRATE
C0303212|T196|1306065|RXNORM|CHROMIUM CR-51|CHROMIUM CR-51
C0078781|T121|1306063|RXNORM|ZINC GLYCINATE|ZINC GLYCINATE
C0077375|T121|38865|RXNORM|TROFOSFAMIDE|TROFOSFAMIDE
C0077376|T121|38866|RXNORM|TROLAMINE SALICYLATE|TROLAMINE SALICYLATE
C3475152|T121|1306060|RXNORM|THERMUS THERMOPHILUS LYSATE|THERMUS THERMOPHILUS LYSATE
C2961540|T121|1053132|RXNORM|HYPROMELLOSE / NAPHAZOLINE / POLYSORBATE 80 / ZINC SULFATE|HYPROMELLOSE / NAPHAZOLINE / POLYSORBATE 80 / ZINC SULFATE
C3255959|T109|1424904|RXNORM|MASTOCARPUS STELLATUS EXTRACT|MASTOCARPUS STELLATUS ALGAE EXTRACT
C2828373|T130|1424906|RXNORM|METHACRYLATE|METHACRYLATE
C1572775|T121|1306068|RXNORM|OXIDRONATE|OXIDRONATE
C1576847|T121|994438|RXNORM|CALCIUM AMINO ACID CHELATE|CALCIUM AMINO ACID CHELATE
C0008163|T121|2346|RXNORM|CHLORAMBUCIL|CHLORAMBUCIL
C0016299|T121|4462|RXNORM|FLUOCINONIDE|FLUOCINONIDE
C0016301|T121|4463|RXNORM|FLUOCORTOLONE|FLUOCORTOLONE
C2700141|T129|1492300|RXNORM|VACCINIA VIRUS STRAIN NEW YORK CITY BOARD OF HEALTH LIVE ANTIGEN|VACCINIA VIRUS STRAIN NEW YORK CITY BOARD OF HEALTH LIVE ANTIGEN
C0078847|T121|40001|RXNORM|ZOPICLONE|ZOPICLONE
C3486032|T109|1426673|RXNORM|PEG-PPG-14-4 DIMETHICONE|PEG-PPG-14-4 DIMETHICONE
C2741006|T129|900108|RXNORM|ONESEED JUNIPER POLLEN EXTRACT|JUNIPERUS MONOSPERMA POLLEN EXTRACT
C0036147|T196|9549|RXNORM|SAMARIUM|SAMARIUM
C2987648|T121|1430438|RXNORM|AFATINIB|AFATINIB
C3651719|T122|1430439|RXNORM|HYDROXYETHYL CELLULOSE (5500 MPA.S AT 2%)|HYDROXYETHYL CELLULOSE (5500 MPA.S AT 2%)
C0060203|T121|24876|RXNORM|FENTICONAZOLE|FENTICONAZOLE
C2937545|T121|1009387|RXNORM|DEXAMETHASONE / NEOMYCIN / THIABENDAZOLE|DEXAMETHASONE / NEOMYCIN / THIABENDAZOLE
C2740956|T129|900031|RXNORM|ATLANTIC SALMON ALLERGENIC EXTRACT|ATLANTIC SALMON ALLERGENIC EXTRACT
C2739878|T129|897304|RXNORM|ALLSCALE POLLEN EXTRACT|ATRIPLEX POLYCARPA POLLEN EXTRACT
C3832727|T109|1539423|RXNORM|ARTEMISIA UMBELLIFORMIS WHOLE EXTRACT|ARTEMISIA UMBELLIFORMIS WHOLE EXTRACT
C3474239|T109|1426672|RXNORM|PEG-PPG-20-20 DIMETHICONE|PEG-PPG-20-20 DIMETHICONE
C3832726|T109|1539422|RXNORM|AMARANTHUS HYPOCHONDRIACUS WHOLE EXTRACT|AMARANTHUS HYPOCHONDRIACUS WHOLE EXTRACT
C1165607|T121|349948|RXNORM|SARRACENIA PURPUREA PREPARATION|SARRACENIA PURPUREA PREPARATION
C3853839|T129|1597258|RXNORM|BLINATUMOMAB|BLINATUMOMAB
C1875387|T121|705040|RXNORM|IODINE / SODIUM IODIDE|IODINE / SODIUM IODIDE
C3832725|T109|1539421|RXNORM|ADANSONIA DIGIATA WHOLE EXTRACT|ADANSONIA DIGIATA WHOLE EXTRACT
C3487972|T121|1324597|RXNORM|JUGLANS REGIA LEAF EXTRACT|JUGLANS REGIA LEAF EXTRACT
C3486722|T121|1324596|RXNORM|BUFO BUFO CUTANEOUS GLAND PREPARATION|COMMON TOAD CUTANEOUS GLAND PREPARATION
C3486656|T121|1324595|RXNORM|CALIFORNIA SHEEPHEAD PREPARATION|CALIFORNIA SHEEPHEAD PREPARATION
C3486655|T121|1324594|RXNORM|ULEX EUROPAEUS FLOWER EXTRACT|ULEX EUROPAEUS FLOWER EXTRACT
C2080591|T121|817486|RXNORM|IODINATED GLYCEROL / PHENYLPROPANOLAMINE|IODINATED GLYCEROL / PHENYLPROPANOLAMINE
C3832731|T109|1539427|RXNORM|SCUTELLARIA ALPINA FLOWERING TOP EXTRACT|SCUTELLARIA ALPINA FLOWERING TOP EXTRACT
C2106236|T121|817482|RXNORM|COAL TAR / JUNIPER TAR / PINE TAR|COAL TAR / JUNIPER TAR / PINE TAR
C2106231|T121|812483|RXNORM|BORIC ACID / COAL TAR|BORIC ACID / COAL TAR
C3832730|T109|1539426|RXNORM|MAGNOLIA X ALBA FLOWER OIL|MAGNOLIA X ALBA FLOWER OIL
C3832729|T109|1539425|RXNORM|KALANCHOE PINNATA LEAF EXTRACT|KALANCHOE PINNATA LEAF EXTRACT
C1875678|T121|689963|RXNORM|POTASSIUM ACETATE / POTASSIUM BICARBONATE / POTASSIUM CITRATE|POTASSIUM ACETATE / POTASSIUM BICARBONATE / POTASSIUM CITRATE
C3832728|T109|1539424|RXNORM|EPILOBIUM ANGUSTIFOLIUM WHOLE EXTRACT|EPILOBIUM ANGUSTIFOLIUM WHOLE EXTRACT
C0063815|T121|27779|RXNORM|IOPENTOL|IOPENTOL
C2364933|T121|806626|RXNORM|GLYCINE ZINC CHELATE|GLYCINE ZINC CHELATE
C0771447|T121|236196|RXNORM|FERROUS OXALATE|FERROUS OXALATE
C0281385|T196|81638|RXNORM|STRONTIUM-89|STRONTIUM-89
C0086024|T127|42604|RXNORM|COBALAMINS|COBALAMINS
C3266927|T121|1342455|RXNORM|ERIODICTYON CALIFORNICUM LEAF EXTRACT|ERIODICTYON CALIFORNICUM LEAF EXTRACT
C2193944|T121|816812|RXNORM|ACETANILIDE / ASPIRIN / CAFFEINE / EPHEDRINE|ACETANILIDE / ASPIRIN / CAFFEINE / EPHEDRINE
C0770956|T121|235784|RXNORM|CALCIUM LACTOBIONATE|CALCIUM LACTOBIONATE
C0032493|T121|8521|RXNORM|POLYGELINE|POLYGELINE
C0164858|T121|59860|RXNORM|CHLORPROETHAZINE|CHLORPROETHAZINE
C3818757|T130|1492940|RXNORM|FLORBETABEN F-18|FLORBETABEN F-18
C3818756|T121|1492941|RXNORM|SUS SCROFA EAR PREPARATION|SUS SCROFA EAR PREPARATION
C0132326|T121|53654|RXNORM|NEVIRAPINE|NEVIRAPINE
C2946720|T121|1039701|RXNORM|ETHANOL / TRICLOSAN|ETHANOL / TRICLOSAN
C0038432|T195|10114|RXNORM|STREPTOZOCIN|STREPTOZOCIN
C0065583|T123|29209|RXNORM|MALIC ACID|MALIC ACID
C3474186|T121|1300389|RXNORM|BORDETELLA PERTUSSIS FILAMENTOUS HEMAGGLUTININ VACCINE, INACTIVATED / BORDETELLA PERTUSSIS TOXOID VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED|BORDETELLA PERTUSSIS FILAMENTOUS HEMAGGLUTININ VACCINE, INACTIVATED / BORDETELLA PERTUSSIS TOXOID VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED
C3474186|T121|1300389|RXNORM|BORDETELLA PERTUSSIS FILAMENTOUS HEMAGGLUTININ VACCINE, INACTIVATED / BORDETELLA PERTUSSIS TOXOID VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED|BORDETELLA PERTUSSIS FILAMENTOUS HEMAGGLUTININ VACCINE, INACTIVATED / BORDETELLA PERTUSSIS TOXOID VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED
C1455147|T121|475342|RXNORM|DASATINIB|DASATINIB
C3537415|T121|1426677|RXNORM|TRIMETHYLSILOXYSILICATE (M-Q 0.6-0.8)|TRIMETHYLSILOXYSILICATE (M-Q 0.6-0.8)
C3666865|T121|1437851|RXNORM|MELICOPE PTELEIFOLIA LEAF EXTRACT|MELICOPE PTELEIFOLIA LEAF EXTRACT
C3498010|T109|1427016|RXNORM|PEG-3 DISTEAROYLAMIDOETHYLMONIUM METHOSULFATE|PEG-3 DISTEAROYLAMIDOETHYLMONIUM METHOSULFATE
C3486306|T121|1427017|RXNORM|HEXYLDECYL MYRISTOYL METHYLAMINOPROPIONATE|HEXYLDECYL MYRISTOYL METHYLAMINOPROPIONATE
C0521959|T125|1427014|RXNORM|SOMETRIBOVE|SOMETRIBOVE
C3257691|T121|1427015|RXNORM|RICE GERM PREPARATION|RICE GERM PREPARATION
C3256861|T109|1427010|RXNORM|PROPYLENE GLYCOL MONOPALMITOSTEARATE|PROPYLENE GLYCOL MONOPALMITOSTEARATE
C3204993|T109|1427011|RXNORM|PROPYLHEPTYL CAPRYLATE|PROPYLHEPTYL CAPRYLATE
C0939937|T121|285279|RXNORM|HONEY PREPARATION|HONEY PREPARATION
C3643357|T122|1421889|RXNORM|POLYGLYCERYL-10 DECAOLEATE|POLYGLYCERYL-10 DECAOLEATE
C0772089|T121|236778|RXNORM|TROSPIUM|TROSPIUM
C3643358|T121|1421886|RXNORM|FESTUCA PRATENSIS TOP EXTRACT|FESTUCA PRATENSIS TOP EXTRACT
C3643359|T121|1421885|RXNORM|CHENOPODIUM ALBUM WHOLE EXTRACT|CHENOPODIUM ALBUM WHOLE EXTRACT
C0772080|T121|236770|RXNORM|TALNIFLUMATE|TALNIFLUMATE
C0380393|T121|115698|RXNORM|ZIPRASIDONE|ZIPRASIDONE
C3256306|T121|1307957|RXNORM|MIMOSA TENUIFLORA BARK EXTRACT|MIMOSA TENUIFLORA BARK EXTRACT
C3858053|T121|1552240|RXNORM|IODINE / ISOPROPYL ALCOHOL / POTASSIUM IODIDE|IODINE / ISOPROPYL ALCOHOL / POTASSIUM IODIDE
C2722054|T129|891641|RXNORM|LIMA BEAN ALLERGENIC EXTRACT|LIMA BEAN ALLERGENIC EXTRACT
C2726182|T129|891647|RXNORM|MUNG BEAN ALLERGENIC EXTRACT|MUNG BEAN ALLERGENIC EXTRACT
C2006341|T121|819109|RXNORM|AMMONIUM CHLORIDE / CARBINOXAMINE|AMMONIUM CHLORIDE / CARBINOXAMINE
C2702382|T129|892592|RXNORM|SHRIMP ALLERGENIC EXTRACT|SHRIMP ALLERGENIC EXTRACT
C1612894|T121|1305600|RXNORM|CAPRYLOYL GLYCINE|CAPRYLOYL GLYCINE
C3256300|T122|1305601|RXNORM|CARBOMER INTERPOLYMER TYPE A (ALLYL SUCROSE CROSSLINKED)|CARBOMER INTERPOLYMER TYPE A (ALLYL SUCROSE CROSSLINKED)
C3500566|T121|1314785|RXNORM|COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENATE / POLYSACCHARIDE IRON COMPLEX / PYRIDOXINE / RIBOFLAVIN / SODIUM ASCORBATE / THIAMINE / VITAMIN B 12 / ZINC SULFATE|COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENATE / POLYSACCHARIDE IRON COMPLEX / PYRIDOXINE / RIBOFLAVIN / SODIUM ASCORBATE / THIAMINE / VITAMIN B 12 / ZINC SULFATE
C0304105|T109|1305608|RXNORM|FENNEL OIL|FENNEL OIL
C3848555|T196|1546366|RXNORM|SELENATE ION|SELENATE ION
C3848557|T196|1546364|RXNORM|TRIIODIDE ION|TRIIODIDE ION
C1874195|T121|690789|RXNORM|AMINOPHYLLINE / EPHEDRINE / PHENOBARBITAL|AMINOPHYLLINE / EPHEDRINE / PHENOBARBITAL
C3848701|T121|1546362|RXNORM|ZINC PICRATE|ZINC PICRATE
C0209227|T121|68099|RXNORM|FAMCICLOVIR|FAMCICLOVIR
C3848560|T121|1546360|RXNORM|ZINC VALERATE|ZINC VALERATE
C0033706|T123|1441688|RXNORM|PROTHROMBIN|PROTHROMBIN
C3855324|T109|1547713|RXNORM|C12-15 ALKYL ETHYLHEXANOATE|C12-15 ALKYL ETHYLHEXANOATE
C1874193|T121|690787|RXNORM|AMINOPHYLLINE / EPHEDRINE|AMINOPHYLLINE / EPHEDRINE
C0209211|T121|68092|RXNORM|LANREOTIDE|LANREOTIDE
C2717561|T121|1439816|RXNORM|RIOCIGUAT|RIOCIGUAT
C3853719|T121|1593200|RXNORM|TRIGONELLA FOENUM-GRAECUM WHOLE EXTRACT|TRIGONELLA FOENUM-GRAECUM WHOLE EXTRACT
C0285590|T121|83008|RXNORM|BICALUTAMIDE|BICALUTAMIDE
C3256545|T122|1371947|RXNORM|POLOXAMER 181|POLOXAMER 181
C1095907|T121|319828|RXNORM|BUCKTHORN PREPARATION|BUCKTHORN PREPARATION
C2929319|T121|1008415|RXNORM|LIDOCAINE / ZINC SULFATE|LIDOCAINE / ZINC SULFATE
C0002686|T121|1006654|RXNORM|AMPROLIUM|AMPROLIUM
C2929321|T121|1008417|RXNORM|CHLORMADINONE / ETHINYL ESTRADIOL|CHLORMADINONE / ETHINYL ESTRADIOL
C2929320|T121|1008416|RXNORM|ASCORBIC ACID / RIBOFLAVIN|ASCORBIC ACID / RIBOFLAVIN
C2929315|T121|1008411|RXNORM|MEPIVACAINE / NOREPINEPHRINE|MEPIVACAINE / NOREPINEPHRINE
C2929314|T121|1008410|RXNORM|CROTAMITON / FLUOCINOLONE|CROTAMITON / FLUOCINOLONE
C2929317|T121|1008413|RXNORM|FORMALDEHYDE / GLUTARAL|FORMALDEHYDE / GLUTARAL
C2929316|T121|1008412|RXNORM|ALGINIC ACID / ALUMINUM HYDROXIDE|ALGINIC ACID / ALUMINUM HYDROXIDE
C0009968|T196|2837|RXNORM|COPPER|COPPER
C2929323|T121|1008419|RXNORM|RESORCINOL / SULFUR / TRICLOSAN|RESORCINOL / SULFUR / TRICLOSAN
C2929322|T121|1008418|RXNORM|BROMHEXINE / FOMINOBEN|BROMHEXINE / FOMINOBEN
C1874507|T121|690254|RXNORM|BENZOCAINE / CETALKONIUM CHLORIDE|BENZOCAINE / CETALKONIUM CHLORIDE
C0012203|T131|3390|RXNORM|DIETHYLSTILBESTROL|DIETHYLSTILBESTROL
C0012228|T121|3393|RXNORM|DIFLUNISAL|DIFLUNISAL
C0012227|T121|3392|RXNORM|DIFLUCORTOLONE|DIFLUCORTOLONE
C1874503|T121|690250|RXNORM|BENZOCAINE / CALCIUM CARBONATE / MAGNESIUM CARBONATE / PHENOBARBITAL|BENZOCAINE / CALCIUM CARBONATE / MAGNESIUM CARBONATE / PHENOBARBITAL
C0064777|T121|28554|RXNORM|LETOSTEINE|LETOSTEINE
C2928302|T121|1007380|RXNORM|DIAZEPAM / ISOPROPAMIDE|DIAZEPAM / ISOPROPAMIDE
C2928303|T121|1007381|RXNORM|NITROFURANTOIN / TETRACAINE|NITROFURANTOIN / TETRACAINE
C2928745|T121|1007830|RXNORM|DEHYDROCHOLATE / PEPSIN A|DEHYDROCHOLATE / PEPSIN A
C2928305|T121|1007383|RXNORM|ATTAPULGITE / MORPHINE|ATTAPULGITE / MORPHINE
C2928751|T121|1007836|RXNORM|BENZALKONIUM / POLYETHYLENES|BENZALKONIUM / POLYETHYLENES
C2928752|T121|1007837|RXNORM|ARACHIS OIL / CALAMINE|CALAMINE / PEANUT OIL
C2928749|T121|1007834|RXNORM|POTASSIUM BICARBONATE / POTASSIUM TARTRATE|POTASSIUM BICARBONATE / POTASSIUM TARTRATE
C2928750|T121|1007835|RXNORM|CALCIUM CITRATE / CHOLECALCIFEROL|CALCIUM CITRATE / CHOLECALCIFEROL
C2928310|T121|1007388|RXNORM|LACTASE / RENNET|LACTASE / RENNET
C2928311|T121|1007389|RXNORM|ECHINACEA PREPARATION / GOLDEN SEAL ROOT|ECHINACEA PREPARATION / GOLDEN SEAL ROOT
C0077275|T125|38782|RXNORM|TRIPTORELIN|TRIPTORELIN
C2106244|T121|814631|RXNORM|COAL TAR / RESORCINOL / SALICYLIC ACID|COAL TAR / RESORCINOL / SALICYLIC ACID
C0015518|T126|4262|RXNORM|FACTOR X|FACTOR X
C0066165|T121|29704|RXNORM|METHOXYPHENAMINE|METHOXYPHENAMINE
C2698371|T121|863035|RXNORM|BEPOTASTINE|BEPOTASTINE
C3819171|T121|1537197|RXNORM|HYDROCORTISONE / LIDOCAINE / PRAMOXINE|HYDROCORTISONE / LIDOCAINE / PRAMOXINE
C3819172|T121|1537193|RXNORM|BENZETHONIUM / DIPHENHYDRAMINE / HYDROCORTISONE|BENZETHONIUM / DIPHENHYDRAMINE / HYDROCORTISONE
C2169318|T121|818284|RXNORM|HYDROCHLOROTHIAZIDE / RAMIPRIL|HYDROCHLOROTHIAZIDE / RAMIPRIL
C2725876|T129|891502|RXNORM|ARABICA COFFEE BEAN ALLERGENIC EXTRACT|ARABICA COFFEE BEAN ALLERGENIC EXTRACT
C3538056|T121|1371949|RXNORM|ERIODICTYON CALIFORNICUM FLOWERING TOP EXTRACT|ERIODICTYON CALIFORNICUM FLOWERING TOP EXTRACT
C2701586|T129|852440|RXNORM|COTTON SEED ALLERGENIC EXTRACT|COTTON SEED ALLERGENIC EXTRACT
C0076652|T121|38252|RXNORM|TIANEPTINE|TIANEPTINE
C0359028|T121|106970|RXNORM|ECONAZOLE / HYDROCORTISONE|ECONAZOLE / HYDROCORTISONE
C0045010|T125|5542|RXNORM|HYDROXYPROGESTERONE|HYDROXYPROGESTERONE
C2183728|T121|818281|RXNORM|DIPHENHYDRAMINE / MENTHOL|DIPHENHYDRAMINE / MENTHOL
C3538363|T121|1372633|RXNORM|ATRACTYLODES MACROCEPHALA ROOT EXTRACT|ATRACTYLODES MACROCEPHALA ROOT EXTRACT
C3538362|T121|1372632|RXNORM|ALISMA PLANTAGO-AQUATICA SUBSP. ORIENTALE ROOT EXTRACT|ALISMA PLANTAGO-AQUATICA SUBSP. ORIENTALE ROOT EXTRACT
C3538365|T121|1372635|RXNORM|IMMATURE CITRUS AURANTIUM FRUIT EXTRACT|IMMATURE CITRUS AURANTIUM FRUIT EXTRACT
C3538364|T121|1372634|RXNORM|BIDENS PILOSA WHOLE EXTRACT|BIDENS PILOSA WHOLE EXTRACT
C3538367|T121|1372637|RXNORM|POLYGONATUM SIBIRICUM ROOT EXTRACT|POLYGONATUM SIBIRICUM ROOT EXTRACT
C3538366|T121|1372636|RXNORM|ILEX PEDUNCULOSA WHOLE EXTRACT|ILEX PEDUNCULOSA WHOLE EXTRACT
C0110806|T109|1309387|RXNORM|COSTUS ROOT OIL|COSTUS ROOT OIL
C2725886|T129|976711|RXNORM|PERCH ALLERGENIC EXTRACT|PERCH ALLERGENIC EXTRACT
C2341724|T109|1309385|RXNORM|LAVANDIN OIL|LAVANDIN OIL
C0939226|T121|284630|RXNORM|CARBINOXAMINE / HYDROCODONE / PSEUDOEPHEDRINE|CARBINOXAMINE / HYDROCODONE / PSEUDOEPHEDRINE
C0939234|T122|284637|RXNORM|HYLAN G-F 20|HYLAN G-F 20
C0939233|T121|284636|RXNORM|HYDROCHLOROTHIAZIDE / TELMISARTAN|HYDROCHLOROTHIAZIDE / TELMISARTAN
C0939232|T121|284635|RXNORM|FLUTICASONE / SALMETEROL|FLUTICASONE / SALMETEROL
C0032831|T197|8597|RXNORM|POTASSIUM IODIDE|POTASSIUM IODIDE
C0032829|T197|8595|RXNORM|POTASSIUM DICHROMATE|POTASSIUM DICHROMATE
C3645179|T121|1426828|RXNORM|DIMETHICONE PEG-15 ACETATE|DIMETHICONE PEG-15 ACETATE
C2194233|T121|812739|RXNORM|ATTAPULGITE / SALICYLIC ACID|ATTAPULGITE / SALICYLIC ACID
C1337244|T109|1309389|RXNORM|EMU OIL|EMU OIL
C0032825|T197|8591|RXNORM|POTASSIUM CHLORIDE|POTASSIUM CHLORIDE
C0032825|T197|8591|RXNORM|POTASSIUM CHLORIDE|POTASSIUM CHLORIDE
C0032825|T197|8591|RXNORM|POTASSIUM CHLORIDE|POTASSIUM CHLORIDE
C2726177|T129|1011060|RXNORM|LIME ALLERGENIC EXTRACT|LIME ALLERGENIC EXTRACT
C2728187|T129|1011066|RXNORM|MACADAMIA NUT ALLERGENIC EXTRACT|MACADAMIA NUT ALLERGENIC EXTRACT
C0947713|T121|287585|RXNORM|GUANETHIDINE / HYDROCHLOROTHIAZIDE|GUANETHIDINE / HYDROCHLOROTHIAZIDE
C0961275|T121|1044269|RXNORM|SELAMECTIN|SELAMECTIN
C0073057|T126|35360|RXNORM|RENNET|RENNET
C0056245|T123|1313334|RXNORM|CONIINE|CONIINE
C1110459|T121|324014|RXNORM|BORON CITRATE|BORON CITRATE
C3486750|T196|1313336|RXNORM|DICHROMATE ION|DICHROMATE ION
C0021758|T129|5891|RXNORM|INTERLEUKIN-4|INTERLEUKIN-4
C0042754|T195|11232|RXNORM|VIRGINIAMYCIN|VIRGINIAMYCIN
C1714000|T130|637320|RXNORM|GADOXETATE DISODIUM|GADOXETATE DISODIUM
C2928446|T121|1007524|RXNORM|ASCORBIC ACID / BIOTIN / FERROUS FUMARATE / FOLIC ACID / MECOBALAMIN / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE|ASCORBIC ACID / BIOTIN / FERROUS FUMARATE / FOLIC ACID / MECOBALAMIN / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE
C2928447|T121|1007525|RXNORM|DEXTROMETHORPHAN / GUAIACOLSULFONATE / GUAIFENESIN|DEXTROMETHORPHAN / GUAIACOLSULFONATE / GUAIFENESIN
C2928448|T121|1007526|RXNORM|GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC|GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC
C2928449|T121|1007527|RXNORM|DEXTROMETHORPHAN / GUAIACOLSULFONATE / GUAIFENESIN / PSEUDOEPHEDRINE|DEXTROMETHORPHAN / GUAIACOLSULFONATE / GUAIFENESIN / PSEUDOEPHEDRINE
C2928442|T121|1007520|RXNORM|DEXCHLORPHENIRAMINE / PSEUDOEPHEDRINE / PYRILAMINE|DEXCHLORPHENIRAMINE / PSEUDOEPHEDRINE / PYRILAMINE
C2928443|T121|1007521|RXNORM|ACETAMINOPHEN / CAFFEINE / PHENYLTOLOXAMINE / SALICYLIC ACID|ACETAMINOPHEN / CAFFEINE / PHENYLTOLOXAMINE / SALICYLIC ACID
C2928444|T121|1007522|RXNORM|ACETAMINOPHEN / CAFFEINE / MAGNESIUM SALICYLATE / PHENYLTOLOXAMINE|ACETAMINOPHEN / CAFFEINE / MAGNESIUM SALICYLATE / PHENYLTOLOXAMINE
C2928445|T121|1007523|RXNORM|ALANINE / ARGININE / CALCIUM CHLORIDE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / SODIUM ACETATE TRIHYDRATE / SODIUM CHLORIDE / THREON|ALANINE / ARGININE / CALCIUM CHLORIDE / DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / SODIUM ACETATE TRIHYDRATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C3163419|T121|1116241|RXNORM|EPHEDRINE / TOLU BALSAM|EPHEDRINE / TOLU BALSAM
C2928450|T121|1007528|RXNORM|ALANINE / ARGININE / CYSTEINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE|ALANINE / ARGININE / CYSTEINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE
C2928451|T121|1007529|RXNORM|ALANINE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE|ALANINE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE
C3667881|T109|1440247|RXNORM|HYDROGENATED RAPESEED OIL|HYDROGENATED RAPESEED OIL
C1875479|T121|691125|RXNORM|MENTHOL / SULFUR|MENTHOL / SULFUR
C3473400|T121|1310029|RXNORM|SENNA ALEXANDRINA SEED EXTRACT|SENNA ALEXANDRINA SEED EXTRACT
C3700985|T109|1486524|RXNORM|CARBOXYETHYL SILICONATE|CARBOXYETHYL SILICONATE
C1875476|T121|691122|RXNORM|MENTHOL / PRAMOXINE|MENTHOL / PRAMOXINE
C1875482|T121|691129|RXNORM|MEPROBAMATE / TRIDIHEXETHYL|MEPROBAMATE / TRIDIHEXETHYL
C1613391|T121|614534|RXNORM|ABACAVIR / LAMIVUDINE|ABACAVIR / LAMIVUDINE
C2025215|T121|817105|RXNORM|CARISOPRODOL / PIROXICAM|CARISOPRODOL / PIROXICAM
C3695943|T129|1484937|RXNORM|COLONIAL BENT GRASS POLLEN EXTRACT|COMMON BENT POLLEN EXTRACT
C3853878|T121|1549329|RXNORM|BLUEBERRY EXTRACT|BLUEBERRY EXTRACT
C2756449|T129|968184|RXNORM|TRICHODERMA HARZIANAM EXTRACT|TRICHODERMA HARZIANAM EXTRACT
C0304961|T130|91516|RXNORM|CYANOCOBALAMIN CO57|COBALT (57CO) CYANOCOBALAMINE
C2928779|T121|1007865|RXNORM|ASCORBIC ACID / VITAMIN A / VITAMIN E|ASCORBIC ACID / VITAMIN A / VITAMIN E
C2741270|T129|900731|RXNORM|SLASH PINE POLLEN EXTRACT|PINUS ELLIOTTII POLLEN EXTRACT
C0058426|T121|23420|RXNORM|DIPROPYLACETAMIDE|DIPROPYLACETAMIDE
C2928778|T121|1007864|RXNORM|CALCIUM PHOSPHATE / VITAMIN B 12|CALCIUM PHOSPHATE / VITAMIN B 12
C2825257|T121|1250203|RXNORM|ROBENACOXIB|ROBENACOXIB
C0075765|T121|82665|RXNORM|DETAJMIUM|DETAJMIUM
C2344277|T129|798232|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 9V CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 9V CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C3666958|T121|1438056|RXNORM|BOLETUS SATANAS FRUITING BODY EXTRACT|BOLETUS SATANAS FRUITING BODY EXTRACT
C3666959|T121|1438057|RXNORM|BLACK CARROT ANTHOCYANINS EXTRACT|BLACK CARROT ANTHOCYANINS EXTRACT
C0037532|T197|9894|RXNORM|SODIUM NITRITE|SODIUM NITRITE
C2928783|T121|1007869|RXNORM|CALCIUM CARBONATE / VITAMIN A / VITAMIN D|CALCIUM CARBONATE / VITAMIN A / VITAMIN D
C1875647|T121|689742|RXNORM|PHENIRAMINE / PHENYLPROPANOLAMINE / PYRILAMINE|PHENIRAMINE / PHENYLPROPANOLAMINE / PYRILAMINE
C1875648|T121|689744|RXNORM|PHENOBARBITAL / PHENYTOIN|PHENOBARBITAL / PHENYTOIN
C1875649|T121|689745|RXNORM|PHENOBARBITAL / POTASSIUM IODIDE / SODIUM BICARBONATE / THEOBROMINE|PHENOBARBITAL / POTASSIUM IODIDE / SODIUM BICARBONATE / THEOBROMINE
C0037530|T121|9892|RXNORM|SODIUM MORRHUATE|SODIUM MORRHUATE
C2928782|T121|1007868|RXNORM|SULFUR / ZINC PYRITHIONE|SULFUR / ZINC PYRITHIONE
C1875652|T121|689748|RXNORM|PHENOL / RESORCINOL|PHENOL / RESORCINOL
C2701380|T129|852178|RXNORM|GRAY BIRCH POLLEN EXTRACT|GRAY BIRCH POLLEN EXTRACT
C0009002|T121|2594|RXNORM|ASTRAGALUS ROOT|CLOFIBRATE
C0037537|T121|9899|RXNORM|SODIUM OXYBATE|SODIUM OXYBATE
C1302109|T121|392553|RXNORM|TRANYLCYPROMINE / TRIFLUOPERAZINE|TRANYLCYPROMINE / TRIFLUOPERAZINE
C1302114|T121|392556|RXNORM|BENZOYL PEROXIDE / ERYTHROMYCIN|BENZOYL PEROXIDE / ERYTHROMYCIN
C0065972|T121|29528|RXNORM|MEQUITAZINE|MEQUITAZINE
C0938435|T121|802755|RXNORM|LIVER STOMACH CONCENTRATE|LIVER STOMACH CONCENTRATE
C2080625|T121|817816|RXNORM|MEPHOBARBITAL / PHENYTOIN|MEPHOBARBITAL / PHENYTOIN
C3535907|T121|1370462|RXNORM|HYDROXYSTEARATE|HYDROXYSTEARATE
C0178487|T127|1370460|RXNORM|ASCORBATE|ASCORBATE
C3535631|T121|1370466|RXNORM|JUGLANS NIGRA WHOLE EXTRACT|JUGLANS NIGRA WHOLE EXTRACT
C0015833|T121|1370467|RXNORM|FENNEL EXTRACT|FENNEL EXTRACT
C3535633|T121|1370464|RXNORM|BEEF LUNG PREPARATION|BEEF LUNG PREPARATION
C2929787|T121|1008890|RXNORM|DIBUCAINE / PREDNISOLONE|DIBUCAINE / PREDNISOLONE
C3535630|T121|1370468|RXNORM|FLUKE, UNSPECIFIED PREPARATION|FLUKE, UNSPECIFIED PREPARATION
C0949117|T121|1370469|RXNORM|ONION EXTRACT|ONION EXTRACT
C0022614|T121|6130|RXNORM|KETAMINE|KETAMINE
C0771473|T121|236220|RXNORM|AMMONIUM SALICYLATE|AMMONIUM SALICYLATE
C0022625|T121|6135|RXNORM|KETOCONAZOLE|KETOCONAZOLE
C0022625|T121|6135|RXNORM|KETOCONAZOLE|KETOCONAZOLE
C2725341|T121|880350|RXNORM|KRILL OIL|KRILL OIL
C3256394|T109|1425221|RXNORM|CETYL STEARATE|CETYL STEARATE
C3256392|T121|1425220|RXNORM|CETETH-2|CETETH-2
C3855323|T121|1547712|RXNORM|ACMELLA OLERACEA FLOWERING TOP EXTRACT|ACMELLA OLERACEA FLOWERING TOP EXTRACT
C0064474|T121|28303|RXNORM|CLORSULON|CLORSULON
C1828724|T123|1291425|RXNORM|DOCOSAENOIC ACID|DOCOSAENOIC ACID
C0035857|T130|9471|RXNORM|ROSE BENGAL|ROSE BENGAL
C0220893|T121|70619|RXNORM|PHENYLACETATE|PHENYLACETATE
C2731478|T109|895385|RXNORM|SUGAR MAPLE POLLEN EXTRACT|SUGAR MAPLE POLLEN EXTRACT
C0975057|T121|308814|RXNORM|BROWN MIXTURE|BROWN MIXTURE
C0771853|T121|236564|RXNORM|MAGNESIUM GLUCONOGLUCEPTATE|MAGNESIUM GLUCONOGLUCEPTATE
C0717495|T121|214301|RXNORM|BENZOCAINE / TRIMETHOBENZAMIDE|BENZOCAINE / TRIMETHOBENZAMIDE
C2741345|T129|900999|RXNORM|PIN OAK POLLEN EXTRACT|QUERCUS PALUSTRIS POLLEN EXTRACT
C1572407|T129|852797|RXNORM|WHEAT SMUT ALLERGENIC EXTRACT|TILLETIA CARIES ALLERGENIC EXTRACT
C1874547|T121|690419|RXNORM|BETAMETHASONE / CALCIPOTRIENE|BETAMETHASONE / CALCIPOTRIENE
C0018988|T123|5175|RXNORM|HEMIN|HEMIN
C3668715|T121|1441303|RXNORM|CAMPHOR / METHYL SALICYLATE|CAMPHOR / METHYL SALICYLATE
C3663777|T121|1433756|RXNORM|1-PROPANAMINIUM, 2-(ACETYLOXY)-3-CARBOXY-N,N,N-TRIMETHYL-, INNER SALT, (2S)-|(S)-ACETYLCARNITINE
C1874536|T121|690411|RXNORM|BENZYL ALCOHOL / SODIUM CHLORIDE|BENZYL ALCOHOL / SODIUM CHLORIDE
C3834050|T121|1543415|RXNORM|PEG-11 AVOCADO GLYCERIDES|PEG-11 AVOCADO GLYCERIDES
C0005036|T131|1311295|RXNORM|BENZENE|BENZENE
C0012551|T129|798304|RXNORM|DIPHTHERIA TOXOID VACCINE, INACTIVATED|DIPHTHERIA TOXOID VACCINE, INACTIVATED
C0771148|T121|235942|RXNORM|BUTETAMATE|BUTETAMATE
C0281398|T121|81647|RXNORM|PHENYLBUTYRATE|PHENYLBUTYRATE
C0281398|T121|81647|RXNORM|PHENYLBUTYRATE|PHENYLBUTYRATE
C0281666|T127|81864|RXNORM|ALITRETINOIN|ALITRETINOIN
C0007745|T123|2243|RXNORM|CERAMIDES|CERAMIDES
C0686816|T007|1544932|RXNORM|BARTONELLA ELIZABETHAE|BARTONELLA ELIZABETHAE
C0059374|T195|24192|RXNORM|ENROFLOXACIN|ENROFLOXACIN
C0102840|T197|46241|RXNORM|ALUMINUM CHLORIDE|ALUMINIUM CHLORIDE
C0102840|T197|46241|RXNORM|ALUMINUM CHLORIDE|ALUMINIUM CHLORIDE
C0102840|T197|46241|RXNORM|ALUMINUM CHLORIDE|ALUMINIUM CHLORIDE
C0102840|T197|46241|RXNORM|ALUMINUM CHLORIDE|ALUMINIUM CHLORIDE
C0102850|T122|46243|RXNORM|ALUMINUM STEARATE|ALUMINUM STEARATE
C0175163|T121|62178|RXNORM|TYBAMATE|TYBAMATE
C0012258|T121|3403|RXNORM|DIGITOXIN|DIGITOXIN
C0253563|T121|75635|RXNORM|EPTIFIBATIDE|EPTIFIBATIDE
C0012265|T121|3407|RXNORM|DIGOXIN|DIGOXIN
C3160109|T121|1112481|RXNORM|CHONDROITIN SULFATES / COLLAGEN / HYALURONATE|CHONDROITIN SULFATES / COLLAGEN / HYALURONATE
C0012271|T121|3409|RXNORM|DIHYDRALAZINE|DIHYDRALAZINE
C3535915|T121|1368629|RXNORM|12-HYDROXYSTEARATE|12-HYDROXYSTEARATE
C3267305|T121|1427123|RXNORM|SPIRULINA MAXIMA PREPARATION|ARTHROSPIRA MAXIMA PREPARATION
C0076840|T121|38413|RXNORM|TORSEMIDE|TORASEMIDE
C1166257|T121|350532|RXNORM|LUESINUM|LUESINUM
C1166258|T121|350533|RXNORM|MEDORRHINUM|MEDORRHINUM
C1166255|T121|350530|RXNORM|TUSSILAGO PETASITES|TUSSILAGO PETASITES
C2929868|T121|1008972|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / OMEGA-3 ACID ETHYL ESTERS (USP) / PYRIDOXINE / VITAMIN B 12|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / OMEGA-3 ACID ETHYL ESTERS (USP) / PYRIDOXINE / VITAMIN B 12
C2929869|T121|1008973|RXNORM|GUAIFENESIN / TERPIN HYDRATE / TETRACYCLINE|GUAIFENESIN / TERPIN HYDRATE / TETRACYCLINE
C2929867|T121|1008971|RXNORM|MONOFLUOROPHOSPHATE / POTASSIUM NITRATE|MONOFLUOROPHOSPHATE / POTASSIUM NITRATE
C2929872|T121|1008976|RXNORM|LEVONORGESTREL / PROMESTRIENE|LEVONORGESTREL / PROMESTRIENE
C2929873|T121|1008977|RXNORM|METOCLOPRAMIDE / PANCREATIN|METOCLOPRAMIDE / PANCREATIN
C2929870|T121|1008974|RXNORM|ALUMINUM HYDROXIDE / NIFLUMIC ACID / ORPHENADRINE|ALUMINUM HYDROXIDE / NIFLUMIC ACID / ORPHENADRINE
C2929871|T121|1008975|RXNORM|CAMPHOR / EUCALYPTUS EXTRACT / MENTHOL|CAMPHOR / EUCALYPTUS EXTRACT / MENTHOL
C2929874|T121|1008978|RXNORM|CETYLPYRIDINIUM / PHOLCODINE|CETYLPYRIDINIUM / PHOLCODINE
C2929875|T121|1008979|RXNORM|SULFAETHIDOLE / SULFAMETHIZOLE|SULFAETHIDOLE / SULFAMETHIZOLE
C0007077|T121|2067|RXNORM|CARBROMAL|CARBROMAL
C0069803|T121|32673|RXNORM|OXYBENZONE|OXYBENZONE
C2929528|T121|1008628|RXNORM|4-AMINOBENZOIC ACID / SALICYLIC ACID|4-AMINOBENZOIC ACID / SALICYLIC ACID
C2348308|T121|1006469|RXNORM|DOCONEXENT|DOCONEXENT
C3645268|T122|1427124|RXNORM|TRIISONONANOIN|TRIISONONANOIN
C0771648|T121|236381|RXNORM|PORACTANT ALFA|PORACTANT ALFA
C2929522|T121|1008622|RXNORM|LACTATE / PHENOL / SALICYLIC ACID|LACTATE / PHENOL / SALICYLIC ACID
C2929523|T121|1008623|RXNORM|CALCIUM CARBONATE / FOLIC ACID / VITAMIN B COMPLEX|CALCIUM CARBONATE / FOLIC ACID / VITAMIN B COMPLEX
C2929521|T121|1008621|RXNORM|POTASSIUM NITRATE / SODIUM FLUORIDE|POTASSIUM NITRATE / SODIUM FLUORIDE
C2929526|T121|1008626|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / OMEGA-3 ACID ETHYL ESTERS (USP)|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / OMEGA-3 ACID ETHYL ESTERS (USP)
C2929527|T121|1008627|RXNORM|HELIUM / NITROGEN / OXYGEN|HELIUM / NITROGEN / OXYGEN
C2929524|T121|1008624|RXNORM|NICKEL SULFATE / POTASSIUM BROMIDE / SULFUR|NICKEL SULFATE / POTASSIUM BROMIDE / SULFUR
C2929525|T121|1008625|RXNORM|CHITOSAN / CHROMIUM PICOLINATE|CHITOSAN / CHROMIUM PICOLINATE
C0021761|T129|1367202|RXNORM|INTERLEUKIN-7|INTERLEUKIN-7
C3486574|T121|1367200|RXNORM|TREPONEMA PALLIDUM IMMUNOSERUM RABBIT|TREPONEMA PALLIDUM IMMUNOSERUM RABBIT
C3486581|T129|1367201|RXNORM|STAPHYLOCOCCUS EPIDERMIDIS IMMUNOSERUM RABBIT|STAPHYLOCOCCUS EPIDERMIDIS IMMUNOSERUM RABBIT
C0392144|T197|1367207|RXNORM|SODIUM BISULFATE|SODIUM BISULFATE
C3535917|T121|1368620|RXNORM|CAPRYLOAMPHOPROPIONATE|CAPRYLOAMPHOPROPIONATE
C3535916|T121|1368623|RXNORM|10-HYDROXYDECANOATE|10-HYDROXYDECANOATE
C3495387|T121|1363040|RXNORM|ISOBUTANE|ISOBUTANE
C3651949|T121|1432137|RXNORM|BENZYL ALCOHOL / ISOPROPYL ALCOHOL / PICRATE / TANNIC ACID|BENZYL ALCOHOL / ISOPROPYL ALCOHOL / PICRATE / TANNIC ACID
C0014994|T121|1363043|RXNORM|ETHYL ETHER|ETHYL ETHER
C0012528|T121|1363044|RXNORM|DIPHENYLAMINE|DIPHENYLAMINE
C3256063|T109|1307691|RXNORM|MENTHA ARVENSIS LEAF OIL|MENTHA ARVENSIS LEAF OIL
C0060238|T197|1363046|RXNORM|FERRIC NITRATE|FERRIC NITRATE
C0060279|T197|1363047|RXNORM|FERROUS OXIDE|FERROUS OXIDE
C0063922|T121|1363048|RXNORM|ISOBUTYL ALCOHOL|ISOBUTYL ALCOHOL
C0065600|T121|1363049|RXNORM|MALTITOL|MALTITOL
C3256313|T109|1311568|RXNORM|CARNUBA WAX|CARNUBA WAX
C3473230|T121|1310019|RXNORM|PRUNUS PERSICA LEAF EXTRACT|PRUNUS PERSICA LEAF EXTRACT
C3486720|T121|1310018|RXNORM|ANAMIRTA COCCULUS SEED EXTRACT|ANAMIRTA COCCULUS SEED EXTRACT
C1366036|T130|1311569|RXNORM|TETROFOSMIN|TETROFOSMIN
C0947651|T122|9785|RXNORM|SILVER PREPARATION|SILVER PREPARATION
C3257596|T109|1310011|RXNORM|ROSA MOSCHATA SEED OIL|ROSA MOSCHATA SEED OIL
C0037129|T197|9789|RXNORM|SILVER NITRATE|SILVER NITRATE
C0037129|T197|9789|RXNORM|SILVER NITRATE|SILVER NITRATE
C0074493|T121|36514|RXNORM|SIBUTRAMINE|SIBUTRAMINE
C3486716|T121|1310015|RXNORM|MARSDENIA CONDURANGO BARK EXTRACT|MARSDENIA CONDURANGO BARK EXTRACT
C3486714|T121|1310014|RXNORM|MANDRAGORA OFFICINARUM ROOT EXTRACT|MANDRAGORA OFFICINARUM ROOT EXTRACT
C3486718|T121|1310017|RXNORM|PRUNUS LAUROCERASUS LEAF EXTRACT|PRUNUS LAUROCERASUS LEAF EXTRACT
C3484466|T121|1310016|RXNORM|ROSA DAMASCENA FLOWERING TOP EXTRACT|ROSA DAMASCENA FLOWERING TOP EXTRACT
C3664996|T121|1435103|RXNORM|SACCHARUM OFFICINARUM WHOLE EXTRACT|SACCHARUM OFFICINARUM WHOLE EXTRACT
C3664995|T121|1435102|RXNORM|CORYDALIS DECUMBENS ROOT EXTRACT|CORYDALIS DECUMBENS ROOT EXTRACT
C3664994|T121|1435101|RXNORM|ALTHAEA OFFICINALIS FLOWER EXTRACT|ALTHAEA OFFICINALIS FLOWER EXTRACT
C3664993|T121|1435100|RXNORM|ARGANIA SPINOSA SEED EXTRACT|ARGANIA SPINOSA SEED EXTRACT
C3665000|T122|1435107|RXNORM|CHOLESTERYL-OCTYLDODECYL LAUROYL GLUTAMATE|CHOLESTERYL-OCTYLDODECYL LAUROYL GLUTAMATE
C3664999|T130|1435106|RXNORM|ACID BLACK 52|ACID BLACK 52
C2733073|T121|900937|RXNORM|ALISKIREN / VALSARTAN|ALISKIREN / VALSARTAN
C3664997|T121|1435104|RXNORM|SOPHORA TETRAPTERA FLOWER EXTRACT|SOPHORA TETRAPTERA FLOWER EXTRACT
C3665002|T122|1435109|RXNORM|DIPENTAERYTHRITYL HEXA C5-9 ACID ESTERS|DIPENTAERYTHRITYL HEXA C5-9 ACID ESTERS
C3665001|T122|1435108|RXNORM|DIETHYLENE GLYCOL DIETHYL ETHER|DIETHYLENE GLYCOL DIETHYL ETHER
C0070549|T121|33272|RXNORM|PHENDIMETRAZINE|PHENDIMETRAZINE
C2929927|T121|1009032|RXNORM|BETAINE / ENDOPEPTIDASES|BETAINE / ENDOPEPTIDASES
C0054826|T121|20342|RXNORM|CARPIPRAMINE|CARPIPRAMINE
C0054827|T121|20343|RXNORM|CARPROFEN|CARPROFEN
C3474039|T121|1314267|RXNORM|ASCLEPIAS QUADRIFOLIA WHOLE EXTRACT|ASCLEPIAS QUADRIFOLIA WHOLE EXTRACT
C3488935|T121|1310275|RXNORM|BOS TAURUS PANCREAS PREPARATION|BOVINE PANCREAS PREPARATION
C3488091|T121|1310276|RXNORM|VIROLA SEBIFERA RESIN EXTRACT|VIROLA SEBIFERA RESIN
C3695951|T121|1484765|RXNORM|SALICYLOYL PHYTOSPHINGOSINE|SALICYLOYL PHYTOSPHINGOSINE
C3497622|T121|1310273|RXNORM|BOS TAURUS OVARY PREPARATION|BOVINE OVARY PREPARATION
C2723310|T121|866459|RXNORM|HYDROXYPROPYL CHITOSAN|HYDROXYPROPYL CHITOSAN
C0073987|T195|1311566|RXNORM|SALINOMYCIN|SALINOMYCIN
C3282348|T121|1250990|RXNORM|PROPIONIC ACID / UNDECYLENATE|PROPIONIC ACID / UNDECYLENATE
C3488415|T121|1310279|RXNORM|POLYGONUM AVICULARE TOP EXTRACT|POLYGONUM AVICULARE TOP EXTRACT
C1874649|T121|1009033|RXNORM|CALCIUM CARBONATE / FOLIC ACID / MAGNESIUM CARBONATE|CALCIUM CARBONATE / FOLIC ACID / MAGNESIUM CARBONATE
C3529104|T109|1364131|RXNORM|CAMELLIA SINENSIS SEED OIL|CAMELLIA SINENSIS SEED OIL
C3464059|T121|1314260|RXNORM|3-((L-MENTHYL)OXY)PROPANE-1,2-DIOL|3-((L-MENTHYL)OXY)PROPANE-1,2-DIOL
C2183709|T121|820172|RXNORM|AMMONIUM CHLORIDE / DIPHENHYDRAMINE / SODIUM CITRATE|AMMONIUM CHLORIDE / DIPHENHYDRAMINE / SODIUM CITRATE
C3485561|T121|1310339|RXNORM|CYCLAMEN PURPURASCENS TUBER EXTRACT|CYCLAMEN PURPURASCENS TUBER EXTRACT
C2605120|T121|1314261|RXNORM|4-METHYL-1-(1-METHYLETHYL)-3-CYCLOHEXEN-1-OL|4-METHYL-1-(1-METHYLETHYL)-3-CYCLOHEXEN-1-OL
C1435738|T109|1364132|RXNORM|TALL OIL|TALL OIL
C2928654|T121|1007739|RXNORM|CAMPHOR / MENTHOL / PETROLATUM / PHENOL|CAMPHOR / MENTHOL / PETROLATUM / PHENOL
C2928653|T121|1007738|RXNORM|LUTEIN / VITAMIN E / ZEAXANTHIN|LUTEIN / VITAMIN E / ZEAXANTHIN
C3651774|T121|1428839|RXNORM|MELIA AZEDERACH LEAF EXTRACT|MELIA AZEDERACH LEAF EXTRACT
C3495981|T121|1310251|RXNORM|BOS TAURUS CARTILAGE PREPARATION|BOVINE CARTILAGE PREPARATION
C3273430|T126|1546420|RXNORM|CONDOLIASE|CONDOLIASE
C2928648|T121|1007733|RXNORM|MINERAL OIL / MINERAL OIL, LIGHT|MINERAL OIL / MINERAL OIL, LIGHT
C2928647|T121|1007732|RXNORM|ALBUTEROL / CROMOLYN|ALBUTEROL / CROMOLYN
C2928650|T121|1007735|RXNORM|CAMPHOR / MENTHOL / METHYL SALICYLATE / TURPENTINE|CAMPHOR / MENTHOL / METHYL SALICYLATE / TURPENTINE
C2928649|T121|1007734|RXNORM|ASCORBIC ACID / CRANBERRY PREPARATION|ASCORBIC ACID / CRANBERRY PREPARATION
C2928652|T121|1007737|RXNORM|LECITHIN / VITAMIN A / VITAMIN E|LECITHIN / VITAMIN A / VITAMIN E
C2928651|T121|1007736|RXNORM|AMYLASES / ENDOPEPTIDASES / PAPAIN / PAPAYA PREPARATION|AMYLASES / ENDOPEPTIDASES / PAPAIN / PAPAYA PREPARATION
C0058218|T121|1373478|RXNORM|DIMETHYL FUMARATE|DIMETHYL FUMARATE
C1874235|T121|691339|RXNORM|AMYLASES / PAPAIN|AMYLASES / PAPAIN
C0108245|T121|30193|RXNORM|CAMPHORIC ACID 1-METHYL ESTER|CAMPHORIC ACID 1-METHYL ESTER
C0065986|T197|29542|RXNORM|MERCURY, AMMONIATED|MERCURY CHLORIDE, AMMONIATED
C0065989|T197|29545|RXNORM|MERCURIC OXIDE|MERCURIC OXIDE
C3531142|T121|1366154|RXNORM|ARGININE / FOLIC ACID / PIPERINE / VITAMIN B 12 / VITAMIN B6|ARGININE / FOLIC ACID / PIPERINE / VITAMIN B 12 / VITAMIN B6
C3486781|T121|1311276|RXNORM|SUS SCROFA BONE MARROW PREPARATION|PORCINE BONE MARROW PREPARATION
C2728190|T129|1010926|RXNORM|KIWI FRUIT ALLERGENIC EXTRACT|KIWI FRUIT ALLERGENIC EXTRACT
C0038172|T007|1311275|RXNORM|STAPHYLOCOCCUS AUREUS|STAPHYLOCOCCUS AUREUS
C3486779|T121|1311272|RXNORM|SUS SCROFA BLOOD PREPARATION|PORCINE BLOOD PREPARATION
C0036274|T196|1311273|RXNORM|SCANDIUM|SCANDIUM
C0981919|T129|851965|RXNORM|JUNE GRASS POLLEN EXTRACT|JUNE GRASS POLLEN EXTRACT
C3488210|T121|1311271|RXNORM|GUAIACUM SANCTUM RESIN|GUAIACUM SANCTUM RESIN
C2701198|T129|851969|RXNORM|RABBIT BUSH POLLEN EXTRACT|AMBROSIA DELTOIDEA POLLEN EXTRACT
C0055749|T197|1311278|RXNORM|MERCURIC SULFIDE|MERCURIO SULFIDE
C0030230|T196|1311279|RXNORM|PALLADIUM|PALLADIUM
C0004954|T123|1359|RXNORM|BELLADONNA ALKALOIDS|BELLADONNA ALKALOIDS
C0004954|T123|1359|RXNORM|BELLADONNA ALKALOIDS|BELLADONNA ALKALOIDS
C0004954|T123|1359|RXNORM|BELLADONNA ALKALOIDS|BELLADONNA ALKALOIDS
C3709478|T121|1487518|RXNORM|UMECLIDINIUM / VILANTEROL|UMECLIDINIUM / VILANTEROL
C3256379|T109|1425936|RXNORM|PHORMIDIUM PERSICINUM EXTRACT|PHORMIDIUM PERSICINUM EXTRACT
C3661274|T121|1487514|RXNORM|UMECLIDINIUM|UMECLIDINIUM
C3709473|T121|1487511|RXNORM|BEHENYL BENZOATE|BEHENYL BENZOATE
C0245514|T121|72610|RXNORM|TROGLITAZONE|TROGLITAZONE
C2001521|T195|1040005|RXNORM|CEFTAROLINE|CEFTAROLINE
C0026924|T007|1310907|RXNORM|MYCOBACTERIUM PHLEI|MYCOBACTERIUM PHLEI
C0320003|T004|1310905|RXNORM|TRICHOPHYTON VERRUCOSUM|TRICHOPHYTON VERRUCOSUM
C0033701|T007|1310903|RXNORM|PROTEUS MIRABILIS|PROTEUS MIRABILIS
C0031618|T123|8215|RXNORM|PHOSPHATIDYLETHANOLAMINES|PHOSPHATIDYLETHANOLAMINES
C0317955|T007|1310909|RXNORM|PROPIONIBACTERIUM AVIDUM|PROPIONIBACTERIUM AVIDUM
C0995674|T007|1310908|RXNORM|BREVIBACTERIUM STATIONIS|BREVIBACTERIUM STATIONIS
C1289957|T121|588003|RXNORM|MECLOFENAMATE|MECLOFENAMATE
C2726185|T129|1193003|RXNORM|NEUROSPORA CRASSA ALLERGENIC EXTRACT|NEUROSPORA CRASSA ALLERGENIC EXTRACT
C3486067|T121|1311052|RXNORM|QUERCUS ROBUR NUT EXTRACT|QUERCUS ROBUR NUT EXTRACT
C3489003|T121|1311050|RXNORM|OENANTHE AQUATICA FRUIT EXTRACT|OENANTHE AQUATICA FRUIT EXTRACT
C3485573|T121|1311051|RXNORM|PICEA MARIANA RESIN EXTRACT|PICEA MARIANA RESIN
C1451381|T197|1311056|RXNORM|CAUSTICUM PREPARATION|CAUSTICUM PREPARATION
C3484409|T121|1311057|RXNORM|LYCOPODIUM CLAVATUM SPORE EXTRACT|LYCOPODIUM CLAVATUM SPORE EXTRACT
C3488383|T121|1311054|RXNORM|TANACETUM VULGARE TOP EXTRACT|TANACETUM VULGARE TOP EXTRACT
C1509329|T130|1311059|RXNORM|BRUCINE SULFATE|BRUCINE SULFATE
C0717893|T121|214682|RXNORM|LORATADINE / PSEUDOEPHEDRINE|LORATADINE / PSEUDOEPHEDRINE
C0717892|T121|214681|RXNORM|LOPERAMIDE / SIMETHICONE|LOPERAMIDE / SIMETHICONE
C0717899|T121|214687|RXNORM|MAGNESIUM HYDROXIDE / MINERAL OIL|MAGNESIUM HYDROXIDE / MINERAL OIL
C0717897|T121|214685|RXNORM|MAGALDRATE / SIMETHICONE|MAGALDRATE / SIMETHICONE
C0032017|T125|8366|RXNORM|POSTERIOR PITUITARY HORMONES|POSTERIOR PITUITARY HORMONES
C0717901|T121|214689|RXNORM|MAGNESIUM SALICYLATE / PHENYLTOLOXAMINE|MAGNESIUM SALICYLATE / PHENYLTOLOXAMINE
C0717900|T121|214688|RXNORM|MAGNESIUM LACTATE|MAGNESIUM LACTATE
C0873028|T121|259367|RXNORM|VERONICASTRUM VIRGINICUM ROOT EXTRACT|VERONICASTRUM VIRGINICUM ROOT EXTRACT
C0873027|T121|259366|RXNORM|EYEBRIGHT PREPARATION|EYEBRIGHT PREPARATION
C3540768|T121|1425412|RXNORM|HELIANTHUS ANNUUS WHOLE EXTRACT|HELIANTHUS ANNUUS WHOLE EXTRACT
C3644644|T121|1425413|RXNORM|ELAEIS GUINEENSIS WHOLE EXTRACT|ELAEIS GUINEENSIS WHOLE EXTRACT
C2717174|T129|1366567|RXNORM|RAXIBACUMAB|RAXIBACUMAB
C2698585|T196|1425419|RXNORM|CHOLINE C-11|CHOLINE C-11
C1619962|T129|1112973|RXNORM|BELATACEPT|BELATACEPT
C3204645|T121|1148649|RXNORM|TOCOTRIENOLS / VITAMIN E|TOCOTRIENOLS / VITAMIN E
C3848558|T121|1546363|RXNORM|VERBASCUM DENSIFLORUM WHOLE EXTRACT|VERBASCUM DENSIFLORUM WHOLE EXTRACT
C0059867|T121|24607|RXNORM|ETOFAMIDE|ETOFAMIDE
C2349012|T121|1338620|RXNORM|ULVA LACTUCA EXTRACT|ULVA LACTUCA EXTRACT
C1095894|T121|319815|RXNORM|BRYONIA PREPARATION|BRYONIA PREPARATION
C1095891|T121|319812|RXNORM|SIBERIAN GINSENG PREPARATION|SIBERIAN GINSENG PREPARATION
C1095889|T121|319810|RXNORM|CABBAGE PREPARATION|CABBAGE PREPARATION
C3692880|T121|1442791|RXNORM|BOS TAURUS INTERVERTEBRAL DISC PREPARATION|BOS TAURUS INTERVERTEBRAL DISC PREPARATION
C0066770|T121|30198|RXNORM|MONOOCTANOIN|MONOOCTANOIN
C3833228|T109|1540869|RXNORM|JASMINUM SAMBAC FLOWER EXTRACT|JASMINUM SAMBAC FLOWER EXTRACT
C1095897|T121|319818|RXNORM|ASTRAGALUS PREPARATION|ASTRAGALUS PREPARATION
C0072733|T197|1544140|RXNORM|FERROUS DISULFIDE|FERROUS DISULFIDE
C0876229|T121|261713|RXNORM|MONASCUS PURPUREUS WEST|MONASCUS PURPUREUS WEST
C2000088|T121|784649|RXNORM|ASENAPINE|ASENAPINE
C0043603|T121|11473|RXNORM|LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS SP|PAMIDRONATE
C0043603|T121|11473|RXNORM|LACTOBACILLUS SP|PAMIDRONATE
C0717668|T195|214468|RXNORM|DAUNORUBICIN LIPOSOMAL|DAUNORUBICIN LIPOSOMAL
C0010132|T125|214461|RXNORM|CORTICOTROPIN-RELEASING HORMONE|CORTICORELIN
C2189663|T121|819609|RXNORM|CINNARIZINE / VINCAMINE|CINNARIZINE / VINCAMINE
C3257206|T121|1241763|RXNORM|BIFIDOBACTERIUM BIFIDUM / BIFIDOBACTERIUM LACTIS / LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS CASEI RHAMNOSUS|BIFIDOBACTERIUM BIFIDUM / BIFIDOBACTERIUM LACTIS / LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS CASEI RHAMNOSUS
C0073591|T195|35797|RXNORM|ROSOXACIN|ROSOXACIN
C0061999|T121|26346|RXNORM|GUGULU EXTRACT|GUGULU EXTRACT
C0061996|T121|26344|RXNORM|GUAR GUM|GUAR GUM
C2701294|T109|852091|RXNORM|HOG EPITHELIA EXTRACT|HOG EPITHELIA EXTRACT
C2701299|T129|852096|RXNORM|LENS SCALE POLLEN EXTRACT|ATRIPLEX LENTIFORMIS POLLEN EXTRACT
C0061081|T109|25608|RXNORM|GAMMA-ORYZANOL|GAMMA-ORYZANOL
C0014695|T127|4018|RXNORM|ERGOCALCIFEROL|ERGOCALCIFEROL
C0014695|T127|4018|RXNORM|ERGOCALCIFEROL|ERGOCALCIFEROL
C3651760|T109|1428859|RXNORM|2-ETHYL-1,6-HEXANEDIOL|2-ETHYL-1,6-HEXANEDIOL
C2929274|T121|1008369|RXNORM|ETHYNODIOL / QUINESTROL|ETHYNODIOL / QUINESTROL
C2929273|T121|1008368|RXNORM|KOREAN GINSENG PREPARATION / SIBERIAN GINSENG PREPARATION / VITAMIN B 12|KOREAN GINSENG PREPARATION / SIBERIAN GINSENG PREPARATION / VITAMIN B 12
C2929272|T121|1008367|RXNORM|ATROPINE / HYOSCYAMINE / SCOPOLAMINE|ATROPINE / HYOSCYAMINE / SCOPOLAMINE
C2929270|T121|1008365|RXNORM|ALGINIC ACID / POTASSIUM BICARBONATE|ALGINIC ACID / POTASSIUM BICARBONATE
C2929269|T121|1008364|RXNORM|BENZALKONIUM / ETHANOL|BENZALKONIUM / ETHANOL
C2929268|T121|1008363|RXNORM|CLOSTEBOL / NEOMYCIN|CLOSTEBOL / NEOMYCIN
C2929267|T121|1008362|RXNORM|DIPYRONE / SCOPOLAMINE|DIPYRONE / SCOPOLAMINE
C2929265|T121|1008360|RXNORM|ADIPHENINE / PHENOBARBITAL|ADIPHENINE / PHENOBARBITAL
C1827168|T121|687403|RXNORM|IODINE / ISOPROPYL ALCOHOL|IODINE / ISOPROPYL ALCOHOL
C1827353|T121|687408|RXNORM|ACETAMINOPHEN / ISOMETHEPTENE|ACETAMINOPHEN / ISOMETHEPTENE
C1720527|T121|758455|RXNORM|COD LIVER OIL / ZINC OXIDE|COD LIVER OIL / ZINC OXIDE
C2701506|T129|852324|RXNORM|HACKBERRY POLLEN EXTRACT|CELTIS OCCIDENTALIS POLLEN EXTRACT
C3651764|T109|1428854|RXNORM|APRICOT FRUIT OIL|APRICOT FRUIT OIL
C2701502|T129|852320|RXNORM|MESQUITE POLLEN EXTRACT|PROSOPIS JULIFLORA POLLEN EXTRACT
C2701863|T121|852897|RXNORM|AMLODIPINE / HYDROCHLOROTHIAZIDE / VALSARTAN|AMLODIPINE / HYDROCHLOROTHIAZIDE / VALSARTAN
C3666443|T121|1436960|RXNORM|SIRAITIA GROSVENORII FRUIT EXTRACT|SIRAITIA GROSVENORII FRUIT EXTRACT
C1329989|T121|852898|RXNORM|CARBETAPENTANE / DIPHENHYDRAMINE / PHENYLEPHRINE|CARBETAPENTANE / DIPHENHYDRAMINE / PHENYLEPHRINE
C2747097|T129|904859|RXNORM|BARLEY (WHOLE GRAIN) ALLERGENIC EXTRACT|BARLEY (WHOLE GRAIN) ALLERGENIC EXTRACT
C2701510|T129|852329|RXNORM|SALT GRASS POLLEN EXTRACT|DISTICHLIS SPICATA POLLEN EXTRACT
C3651765|T109|1428852|RXNORM|NELUMBO NUCIFERA GERM EXTRACT|NELUMBO NUCIFERA GERM EXTRACT
C3265532|T121|1426781|RXNORM|DIETHYLHEXYL SEBACATE|DIETHYLHEXYL SEBACATE
C3257699|T121|1426780|RXNORM|PEG-PPG-20-6 DIMETHICONE|PEG-PPG-20-6 DIMETHICONE
C3536780|T121|1426783|RXNORM|PANTOLACTONE, (+-)-|PANTOLACTONE, (+-)-
C3495131|T121|1333420|RXNORM|ENTEROBIUS VERMICULARIS PREPARATION|ENTEROBIUS VERMICULARIS PREPARATION
C0164321|T197|1333425|RXNORM|CALCIUM ARSENATE|CALCIUM ARSENATE
C0012052|T121|1362873|RXNORM|DIBUTYL PHTHALATE|DIBUTYL PHTHALATE
C1588587|T197|543375|RXNORM|ALUMINUM SESQUICHLOROHYDRATE|ALUMINUM SESQUICHLOROHYDRATE
C2183726|T121|815866|RXNORM|DIPHENHYDRAMINE / GUAIFENESIN|DIPHENHYDRAMINE / GUAIFENESIN
C0770393|T121|235408|RXNORM|CLORAZEPIC ACID|CLORAZEPIC ACID
C3834094|T121|1541717|RXNORM|CUCURBITA PEPO WHOLE EXTRACT|CUCURBITA PEPO WHOLE EXTRACT
C0758542|T130|230435|RXNORM|TECHNETIUM TC 99M ARCITUMOMAB|TECHNETIUM (99MTC) ARCITUMONMAB
C3256369|T121|1307712|RXNORM|MORUS ALBA ROOT EXTRACT|MORUS ALBA ROOT EXTRACT
C3474133|T121|1307713|RXNORM|KALOPANAX SEPTEMLOBUS BARK EXTRACT|KALOPANAX SEPTEMLOBUS BARK EXTRACT
C3496937|T109|1307710|RXNORM|CRYPTHECODINIUM COHNII DHA OIL|CRYPTHECODINIUM COHNII DHA OIL
C3474281|T121|1307711|RXNORM|JUGLANS NIGRA BARK EXTRACT|JUGLANS NIGRA BARK EXTRACT
C3256463|T121|1307716|RXNORM|TILIA CORDATA FLOWER EXTRACT|TILIA CORDATA FLOWER EXTRACT
C0982074|T168|1307717|RXNORM|CHERRY JUICE|CHERRY JUICE
C3255689|T121|1307714|RXNORM|LILIUM CANDIDUM FLOWER EXTRACT|LILIUM CANDIDUM FLOWER EXTRACT
C3256498|T121|1307715|RXNORM|AQUILARIA MALACCENSIS STEM EXTRACT|AQUILARIA MALACCENSIS STEM EXTRACT
C0001367|T121|281|RXNORM|ACYCLOVIR|ACYCLOVIR
C0001367|T121|281|RXNORM|ACYCLOVIR|ACYCLOVIR
C3257535|T121|1307718|RXNORM|WINE GRAPE EXTRACT|WINE GRAPE EXTRACT
C3256597|T121|1307719|RXNORM|ATRACTYLODES LANCEA ROOT EXTRACT|ATRACTYLODES JAPONICA ROOT EXTRACT
C0063041|T121|27169|RXNORM|LEFLUNOMIDE|LEFLUNOMIDE
C2739934|T129|897403|RXNORM|ORANGE POLLEN EXTRACT|CITRUS SINENSIS POLLEN EXTRACT
C1699163|T121|617568|RXNORM|DEXTROMETHORPHAN / PHENIRAMINE / PHENYLEPHRINE|DEXTROMETHORPHAN / PHENIRAMINE / PHENYLEPHRINE
C0055628|T197|1363045|RXNORM|CHROMIUM OXIDE|CHROMIUM OXIDE
C2980404|T121|1092391|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / OMEGA-3 ACID ETHYL ESTERS (USP) / VITAMIN E|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / OMEGA-3 ACID ETHYL ESTERS (USP) / VITAMIN E
C1958126|T121|1368001|RXNORM|ALOGLIPTIN|ALOGLIPTIN
C2828294|T196|1546415|RXNORM|IODIDE ION I-131|IODIDE ION I-131
C0125654|T121|52014|RXNORM|DIPROPIZINE, (S)-ISOMER|LEVODROPROPIZINE
C2701709|T129|903913|RXNORM|BROAD LEAVED PAPERBARK POLLEN EXTRACT|MELALEUCA QUINQUENERVIA POLLEN EXTRACT
C0125656|T121|52016|RXNORM|MEDETOMIDINE|MEDETOMIDINE
C3663405|T121|1432990|RXNORM|PTYCHOPETALUM OLACOIDES ROOT EXTRACT|PTYCHOPETALUM OLACOIDES ROOT EXTRACT
C2080526|T121|817716|RXNORM|DIMETHINDENE / PHENYLEPHRINE|DIMETHINDENE / PHENYLEPHRINE
C3486623|T121|1352521|RXNORM|HELIANTHEMUM NUMMULARIUM FLOWER EXTRACT|HELIANTHEMUM NUMMULARIUM FLOWER EXTRACT
C0982185|T121|1426255|RXNORM|GLYCOL STEARATE|GLYCOL STEARATE
C3848516|T121|1546416|RXNORM|CHLORTHEOPHYLLINE|CHLORTHEOPHYLLINE
C3504821|T121|1356711|RXNORM|PALMATE|PALMATE
C0004924|T122|1356|RXNORM|METHYL PYRROLIDINE CARBOXYLATE, (-),DL-|BEESWAX
C1720020|T121|645079|RXNORM|CETYLPYRIDINIUM / MENTHOL|CETYLPYRIDINIUM / MENTHOL
C3502818|T109|1356714|RXNORM|THERMUS THERMOPHILUS EXTRACT|THERMUS THERMOPHILUS EXTRACT
C3855805|T121|1549105|RXNORM|LEONURUS CARDIACA FLOWERING TOP EXTRACT|LEONURUS CARDIACA FLOWERING TOP EXTRACT
C3486571|T121|1310042|RXNORM|TOXICODENDRON DIVERSILOBUM LEAF EXTRACT|TOXICODENDRON DIVERSILOBUM LEAF EXTRACT
C0982026|T129|485234|RXNORM|ANTIRABIES SERUM,EQUINE|ANTIRABIES SERUM,EQUINE
C0060180|T121|24853|RXNORM|FENOLDOPAM|FENOLDOPAM
C0060182|T121|24855|RXNORM|FENOVERINE|FENOVERINE
C0060183|T121|24856|RXNORM|FENOXAZOLINE|FENOXAZOLINE
C0008466|T123|2473|RXNORM|CHONDROITIN SULFATES|CHONDROITIN SULFATES
C3818714|T121|1535489|RXNORM|FRITILLARIA CIRRHOSA BULB EXTRACT|FRITILLARIA CIRRHOSA BULB EXTRACT
C3818715|T121|1535488|RXNORM|EUGENIA UNIFLORA WHOLE EXTRACT|EUGENIA UNIFLORA WHOLE EXTRACT
C3833051|T109|1540273|RXNORM|PEG-10 GLYCERYL TRIISOSTEARATE|PEG-10 GLYCERYL TRIISOSTEARATE
C2724903|T121|880341|RXNORM|COCKLEBUR EXTRACT|COCKLEBUR EXTRACT
C0078772|T130|39935|RXNORM|ZINC CARBONATE|ZINC CARBONATE
C0078774|T197|39937|RXNORM|ZINC CHLORIDE|ZINC CHLORIDE
C0086123|T125|42627|RXNORM|DEOXYCHOLATE|DEOXYCHOLATE
C0086108|T130|42625|RXNORM|DEHYDROCHOLATE|DEHYDROCHOLATE
C0076651|T121|1546410|RXNORM|TIAMULIN|TIAMULIN
C0873099|T121|259436|RXNORM|DANDELION ROOT EXTRACT|TARAXACUM OFFICINALE ROOT EXTRACT
C2930003|T121|1009108|RXNORM|HEXETIDINE / NIFLUMIC ACID|HEXETIDINE / NIFLUMIC ACID
C2930004|T121|1009109|RXNORM|GREEN TEA EXTRACT / THEAFLAVIN|GREEN TEA EXTRACT / THEAFLAVIN
C0717539|T121|214344|RXNORM|CALCIUM ACETATE / MAGNESIUM CARBONATE|CALCIUM ACETATE / MAGNESIUM CARBONATE
C2929995|T121|1009100|RXNORM|ASCORBIC ACID / CUPROUS OXIDE / LUTEIN / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / CUPROUS OXIDE / LUTEIN / VITAMIN E / ZINC OXIDE
C2929996|T121|1009101|RXNORM|ALUMINUM OXIDE / MAGNESIUM HYDROXIDE|ALUMINUM OXIDE / MAGNESIUM HYDROXIDE
C2929997|T121|1009102|RXNORM|ERGOTAMINE / LEVOROTATORY ALKALOIDS OF BELLADONNA / PHENOBARBITAL|ERGOTAMINE / LEVOROTATORY ALKALOIDS OF BELLADONNA / PHENOBARBITAL
C2929998|T121|1009103|RXNORM|AMYLASES / ENDOPEPTIDASES|AMYLASES / ENDOPEPTIDASES
C2929999|T121|1009104|RXNORM|CERAMIDES / TRIAMCINOLONE|CERAMIDES / TRIAMCINOLONE
C2930000|T121|1009105|RXNORM|4-AMINOBENZOIC ACID / METHOXSALEN|4-AMINOBENZOIC ACID / METHOXSALEN
C2930001|T121|1009106|RXNORM|CALCIUM BROMIDE / CALCIUM LACTATE|CALCIUM BROMIDE / CALCIUM LACTATE
C2930002|T121|1009107|RXNORM|ASCORBIC ACID / TYROTHRICIN|ASCORBIC ACID / TYROTHRICIN
C0872896|T121|259266|RXNORM|HOPS EXTRACT|HOPS EXTRACT
C3848534|T196|1546411|RXNORM|THIOSULFATE ION|THIOSULFATE ION
C1695579|T126|629565|RXNORM|ALGLUCOSIDASE ALFA|ALGLUCOSIDASE ALFA
C1330001|T121|668889|RXNORM|DIPHENHYDRAMINE / HYDROCODONE / PHENYLEPHRINE|DIPHENHYDRAMINE / HYDROCODONE / PHENYLEPHRINE
C1875261|T121|689910|RXNORM|HYDROCODONE / PHENYLTOLOXAMINE|HYDROCODONE / PHENYLTOLOXAMINE
C0036581|T196|9641|RXNORM|SELENIUM|SELENIUM
C1875262|T121|689914|RXNORM|HYDROCORTISONE / ISOPROPYL ALCOHOL / RESORCINOL / SULFUR|HYDROCORTISONE / ISOPROPYL ALCOHOL / RESORCINOL / SULFUR
C0078442|T121|39684|RXNORM|EPINASTINE|EPINASTINE
C0061629|T109|1427078|RXNORM|GLYCOFUROL|GLYCOFUROL
C1880991|T121|1427079|RXNORM|GLYCOL DIMETHACRYLATE|GLYCOL DIMETHACRYLATE
C3485671|T121|1426654|RXNORM|POLYQUATERNIUM-11 (1000000 MW)|POLYQUATERNIUM-11 (1000000 MW)
C0053091|T121|18867|RXNORM|BENAZEPRIL|BENAZEPRIL
C3152887|T129|1098257|RXNORM|DOUGLAS FIR POLLEN EXTRACT|PSEUDOTSUGA MENZIESII POLLEN EXTRACT
C2949056|T121|1045531|RXNORM|BENZOCAINE / DEXTROMETHORPHAN / MENTHOL|BENZOCAINE / DEXTROMETHORPHAN / MENTHOL
C0259497|T121|1363699|RXNORM|STEARAMIDOETHYL DIETHYLAMINE|STEARAMIDOETHYL DIETHYLAMINE
C0059769|T121|1427072|RXNORM|ETHYL LACTATE|ETHYL LACTATE
C2955001|T121|1049378|RXNORM|BENZALKONIUM / TYLOXAPOL|BENZALKONIUM / TYLOXAPOL
C2928389|T121|1007467|RXNORM|DI-ISOPROPYLAMMONIUM / PROCAINE|DI-ISOPROPYLAMMONIUM / PROCAINE
C0722613|T121|219228|RXNORM|ACETAMINOPHEN / PHENYLTOLOXAMINE|ACETAMINOPHEN / PHENYLTOLOXAMINE
C2697509|T121|1427077|RXNORM|GLYCERYL RICINOLEATE|GLYCERYL RICINOLEATE
C0772024|T197|236719|RXNORM|SODIUM PHOSPHATE, DIBASIC|SODIUM PHOSPHATE, DIBASIC
C0772023|T121|236718|RXNORM|SULFONATED PHENOL|SULFONATED PHENOL
C2741453|T129|901258|RXNORM|WATERMELON ALLERGENIC EXTRACT|WATERMELON ALLERGENIC EXTRACT
C0772018|T121|236713|RXNORM|THEOFIBRATE|THEOFIBRATE
C2927934|T121|1007011|RXNORM|DEQUALINIUM / DIBUNATE|DEQUALINIUM / DIBUNATE
C2702409|T129|891668|RXNORM|SOYBEAN ALLERGENIC EXTRACT|SOYBEAN ALLERGENIC EXTRACT
C0025688|T121|6857|RXNORM|METHOXYFLURANE|METHOXYFLURANE
C2356367|T129|804179|RXNORM|MEASLES VIRUS VACCINE LIVE, ENDERS' ATTENUATED EDMONSTON STRAIN|MEASLES VIRUS VACCINE LIVE, ENDERS' ATTENUATED EDMONSTON STRAIN
C0025677|T121|6851|RXNORM|METHOTREXATE|METHOTREXATE
C3256723|T109|1305660|RXNORM|SANTALUM SPICATUM OIL|SANTALUM SPICATUM OIL
C1177183|T168|1305661|RXNORM|SAGE OIL|SAGE OIL
C0006886|T131|1984|RXNORM|CANTHARIDIN|CANTHARIDIN
C3256258|T109|1305663|RXNORM|ROSA DAMASCENA FLOWER OIL|ROSA DAMASCENA FLOWER OIL
C3256256|T109|1305664|RXNORM|ROSA CENTIFOLIA FLOWER OIL|ROSA CENTIFOLIA FLOWER OIL
C2927939|T121|1007016|RXNORM|ACEPROMAZINE / ACEPROMETAZINE / CLORAZEPIC ACID|ACEPROMAZINE / ACEPROMETAZINE / CLORAZEPIC ACID
C2827309|T109|1305669|RXNORM|POLYOXYL 40 HYDROGENATED CASTOR OIL|POLYOXYL 40 HYDROGENATED CASTOR OIL
C2927940|T121|1007017|RXNORM|NIACINAMIDE / RIBOFLAVIN|NIACINAMIDE / RIBOFLAVIN
C3257521|T121|1372248|RXNORM|COCONUT EXTRACT|COCONUT EXTRACT
C3256023|T121|1372249|RXNORM|CLUSTER FIG EXTRACT|CLUSTER FIG EXTRACT
C1142985|T121|341248|RXNORM|EZETIMIBE|EZETIMIBE
C2979411|T121|1090823|RXNORM|ASCORBIC ACID / BETA CAROTENE / COPPER SULFATE / SELENITE / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / BETA CAROTENE / COPPER SULFATE / SELENITE / VITAMIN E / ZINC OXIDE
C2224242|T121|822929|RXNORM|AMPHETAMINE ASPARTATE / AMPHETAMINE SULFATE / DEXTROAMPHETAMINE SACCHARATE / DEXTROAMPHETAMINE SULFATE|AMPHETAMINE ASPARTATE / AMPHETAMINE SULFATE / DEXTROAMPHETAMINE SACCHARATE / DEXTROAMPHETAMINE SULFATE
C0002260|T121|569|RXNORM|EFLORNITHINE|EFLORNITHINE
C0002260|T121|569|RXNORM|EFLORNITHINE|EFLORNITHINE
C2194328|T121|814386|RXNORM|ACETAMINOPHEN / METHOCARBAMOL|ACETAMINOPHEN / METHOCARBAMOL
C0032487|T122|8519|RXNORM|POLYETHYLENES|POLYETHYLENES
C3853624|T126|560|RXNORM|ALPHA-AMYLASES|ALPHA-AMYLASE
C3819169|T109|1491980|RXNORM|CAPROYL LACTATE|CAPROYL LACTATE
C0066469|T121|29954|RXNORM|METOPIMAZINE|METOPIMAZINE
C2723679|T129|867260|RXNORM|SOUTHERN BAYBERRY POLLEN EXTRACT|MORELLA CERIFERA POLLEN EXTRACT
C0066465|T121|29950|RXNORM|METOCURINE|METOCURINE
C0135166|T121|54365|RXNORM|PAMABROM|PAMABROM
C0071038|T121|33684|RXNORM|PICOLINIC ACID|PICOLINIC ACID
C0071042|T121|33688|RXNORM|PICOSULFATE SODIUM|PICOSULFATE SODIUM
C0212750|T168|68905|RXNORM|BORAGE OIL|STARFLOWER OIL
C0162680|T197|1482913|RXNORM|TECHNETIUM TC 99M SESTAMIBI|TECHNETIUM (99MTC) SESTAMIBI
C2106240|T121|815521|RXNORM|BENZOCAINE / COAL TAR / SALICYLIC ACID|BENZOCAINE / COAL TAR / SALICYLIC ACID
C2586803|T129|830464|RXNORM|RABIES VIRUS VACCINE WISTAR STRAIN PM-1503-3M (HUMAN), INACTIVATED|RABIES VIRUS VACCINE WISTAR STRAIN PM-1503-3M (HUMAN), INACTIVATED
C0004037|T004|1182|RXNORM|ASPERGILLUS FUMIGATUS|ASPERGILLUS FUMIGATUS
C0064803|T123|28574|RXNORM|LEUCOCYANIDIN|LEUCOCYANIDIN
C0025132|T121|6686|RXNORM|MEDIGOXIN|MEDIGOXIN
C2746103|T129|901620|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 1 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 1 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C2006116|T121|821119|RXNORM|CALCIUM CARBONATE / MAGNESIUM OXIDE|CALCIUM CARBONATE / MAGNESIUM OXIDE
C3257595|T109|1356713|RXNORM|MENTHYL PYRROLIDONE CARBOXYLATE, (-),DL-|MENTHYL DL-PYRROLIDONECARBOXYLATE
C0015491|T123|4249|RXNORM|FACTOR IX|FACTOR IX
C2194230|T121|814652|RXNORM|BENZOYL PEROXIDE / MICONAZOLE|BENZOYL PEROXIDE / MICONAZOLE
C0072804|T121|35163|RXNORM|PYRVINIUM|PYRVINIUM
C2194019|T121|819049|RXNORM|BETAMETHASONE / LORATADINE|BETAMETHASONE / LORATADINE
C0020336|T121|5521|RXNORM|HYDROXYCHLOROQUINE|HYDROXYCHLOROQUINE
C2726157|T129|892317|RXNORM|WINE GRAPE ALLERGENIC EXTRACT|WINE GRAPE ALLERGENIC EXTRACT
C0081592|T109|1424668|RXNORM|ANISYL ALCOHOL|ANISYL ALCOHOL
C3256292|T109|1424669|RXNORM|BUTETH-3|BUTETH-3
C0246330|T121|72937|RXNORM|TOLCAPONE|TOLCAPONE
C3256332|T109|1424665|RXNORM|AMMONIO METHACRYLATE COPOLYMER TYPE A|AMMONIO METHACRYLATE COPOLYMER TYPE A
C0000294|T121|44|RXNORM|MESNA|MESNA
C0000294|T121|44|RXNORM|MESNA|MESNA
C0103076|T121|1424667|RXNORM|AMMONIUM LAURYL SULFATE|AMMONIUM LAURYL SULFATE
C3256407|T109|1424661|RXNORM|1,3-DIMETHYLBUTYL SALICYLATE|1,3-DIMETHYLBUTYL SALICYLATE
C3256408|T109|1424662|RXNORM|GLYCERYL 1,3-DIOLEATE|GLYCERYL 1,3-DIOLEATE
C2827302|T109|1486516|RXNORM|POLOXAMER 331|POLOXAMER 331
C3486614|T121|1309819|RXNORM|BETULA PUBESCENS LEAF EXTRACT|BETULA PUBESCENS LEAF EXTRACT
C3488360|T121|1309818|RXNORM|CARPINUS BETULUS FLOWERING TOP EXTRACT|CARPINUS BETULUS FLOWERING TOP EXTRACT
C1950313|T121|1309816|RXNORM|PRUNUS SPINOSA FLOWER BUD EXTRACT|PRUNUS SPINOSA FLOWER BUD EXTRACT
C3486613|T121|1309815|RXNORM|BETULA PENDULA BARK EXTRACT|BETULA PENDULA BARK EXTRACT
C3488928|T109|1309362|RXNORM|HYPERICUM PERFORATUM FLOWER EXTRACT|HYPERICUM PERFORATUM FLOWER EXTRACT
C3488359|T121|1309813|RXNORM|TSUGA CANADENSIS FLOWER BUD EXTRACT|TSUGA CANADENSIS FLOWER BUD EXTRACT
C3486611|T121|1309812|RXNORM|ASPIDOSPERMA QUEBRACHO-BLANCO BARK EXTRACT|ASPIDOSPERMA QUEBRACHO-BLANCO BARK EXTRACT
C3256917|T121|1309811|RXNORM|GARCINIA INDICA SEED BUTTER EXTRACT|GARCINIA INDICA SEED BUTTER EXTRACT
C3153858|T121|1100370|RXNORM|ALPHA TOCOPHEROL / CALCIUM CITRATE / CHOLECALCIFEROL / DOCOSAHEXAENOATE / DOCUSATE / FOLIC ACID / IRON CARBONYL / PYRIDOXINE|ALPHA TOCOPHEROL / CALCIUM CITRATE / CHOLECALCIFEROL / DOCOSAHEXAENOATE / DOCUSATE / FOLIC ACID / IRON CARBONYL / PYRIDOXINE
C1719855|T121|645081|RXNORM|CHLORHEXIDINE / TOLNAFTATE|CHLORHEXIDINE / TOLNAFTATE
C3693004|T197|1443002|RXNORM|DITHIONATE|DITHIONATE
C0137033|T130|1443000|RXNORM|PICRATE|PICRATE
C0072980|T195|35302|RXNORM|SIROLIMUS|SIROLIMUS
C3700895|T109|1486517|RXNORM|MANGIFERA INDICA SEED EXTRACT|MANGIFERA INDICA SEED EXTRACT
C2948509|T121|1044283|RXNORM|ALLANTOIN / BENZOCAINE|ALLANTOIN / BENZOCAINE
C0052929|T121|1440261|RXNORM|BAICALIN|BAICALIN
C0301544|T121|1440266|RXNORM|AMINOMETRADINE|AMINOMETRADINE
C0002583|T131|1440264|RXNORM|AMINOPTERIN|AMINOPTERIN
C2826082|T121|1440268|RXNORM|AMINOPROPAZINE FUMARATE|AMINOPROPAZINE FUMARATE
C0058676|T197|23622|RXNORM|DOLOMITE|DOLOMITE
C0058677|T121|23623|RXNORM|DOMIPHEN|DOMIPHEN
C0172907|T121|61773|RXNORM|FLUTRIMAZOLE|FLUTRIMAZOLE
C2918519|T129|995738|RXNORM|BLACK IMPORTED FIRE ANT ALLERGENIC EXTRACT|SOLENOPSIS RICHTERI ALLERGENIC EXTRACT
C0048306|T125|15070|RXNORM|FORMESTANE|FORMESTANE
C2928431|T121|1007509|RXNORM|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM OXIDE / NIACIN / POTASSIUM IODIDE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM OXIDE / NIACIN / POTASSIUM IODIDE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN E / ZINC OXIDE
C2928428|T121|1007506|RXNORM|EPHEDRINE / GUAIACOLSULFONIC ACID|EPHEDRINE / GUAIACOLSULFONIC ACID
C2928429|T121|1007507|RXNORM|IVERMECTIN / PRAZIQUANTEL / PYRANTEL|IVERMECTIN / PRAZIQUANTEL / PYRANTEL
C2928426|T121|1007504|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / DOCUSATE / FERROUS FUMARATE / FOLIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|ALPHA TOCOPHEROL / ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / DOCUSATE / FERROUS FUMARATE / FOLIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C2928427|T121|1007505|RXNORM|ASCORBIC ACID / BIOTIN / DOCUSATE / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|ASCORBIC ACID / BIOTIN / DOCUSATE / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C3832871|T121|1539812|RXNORM|SODIUM DECYLGLUCOSIDE HYDROXYPROPYLSULFONATE|SODIUM DECYLGLUCOSIDE HYDROXYPROPYLSULFONATE
C2928425|T121|1007503|RXNORM|ACETATE / CYSTEINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / SODIUM BISULFITE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / VALINE|ACETATE / CYSTEINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / SODIUM BISULFITE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / VALINE
C2928422|T121|1007500|RXNORM|ALUMINUM CHLORHYDRATE / ETHANOL|ALUMINUM CHLOROHYDRATE / ETHANOL
C2928423|T121|1007501|RXNORM|ALLANTOIN / PRAMOXINE|ALLANTOIN / PRAMOXINE
C1874798|T121|689371|RXNORM|CHLOROXYLENOL / HYDROCORTISONE / PRAMOXINE|CHLOROXYLENOL / HYDROCORTISONE / PRAMOXINE
C3651700|T121|1431718|RXNORM|HARRISIA POMANENSIS STEM EXTRACT|HARRISIA POMANENSIS STEM EXTRACT
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, HORSE DANDER|PRASTERONE
C3855903|T121|1549307|RXNORM|TRICLOSAN / ZINC OXIDE|TRICLOSAN / ZINC OXIDE
C0011185|T125|3143|RXNORM|ALLERGENIC EXTRACT, HOUSE DUST EXTRACT CONCENTRATE|PRASTERONE
C0084453|T121|41967|RXNORM|SALMON OIL|SALMON OIL
C3537685|T121|1371301|RXNORM|EUPHORBIA THYMIFOLIA WHOLE EXTRACT|EUPHORBIA THYMIFOLIA WHOLE EXTRACT
C1172628|T109|1426415|RXNORM|ALUMINUM STARCH OCTENYLSUCCINATE|ALUMINUM STARCH OCTENYLSUCCINATE
C1874802|T121|689375|RXNORM|CHLOROXYLENOL / RESORCINOL / SULFUR|CHLOROXYLENOL / RESORCINOL / SULFUR
C0068334|T121|31448|RXNORM|ALLERGENIC EXTRACT,FULIGO SEPTICA|NABUMETONE
C2701286|T121|852083|RXNORM|SALT CEDAR POLLEN|SALT CEDAR POLLEN
C2366367|T129|809864|RXNORM|C1 INHIBITOR (HUMAN)|C1 ESTERASE INHIBITOR (HUMAN)
C0876716|T121|262100|RXNORM|RAPACURONIUM|RAPACURONIUM
C1959889|T121|729490|RXNORM|CALCIUM CARBONATE / MAGNESIUM CHLORIDE|CALCIUM CARBONATE / MAGNESIUM CHLORIDE
C3199350|T121|1125499|RXNORM|CALCIUM CARBONATE / CHOLECALCIFEROL / MAGNESIUM OXIDE / ZINC OXIDE|CALCIUM CARBONATE / CHOLECALCIFEROL / MAGNESIUM OXIDE / ZINC OXIDE
C2701331|T129|852128|RXNORM|JOHNSON GRASS SMUT EXTRACT|JOHNSON GRASS SMUT ALLERGENIC EXTRACT
C0206824|T130|1426414|RXNORM|LACTOBIONATE|LACTOBIONATE
C0028365|T195|7517|RXNORM|NORFLOXACIN|NORFLOXACIN
C0028365|T195|7517|RXNORM|NORFLOXACIN|NORFLOXACIN
C0028360|T125|7515|RXNORM|NORETHYNODREL|NORETHYNODREL
C0028356|T125|7514|RXNORM|NORETHINDRONE|NORETHINDRONE
C0028356|T125|7514|RXNORM|NORETHINDRONE|NORETHINDRONE
C0028355|T125|7513|RXNORM|NORETHANDROLONE|NORETHANDROLONE
C0028351|T125|7512|RXNORM|NOREPINEPHRINE|NOREPINEPHRINE
C2701355|T129|852152|RXNORM|GREASEWOOD POLLEN EXTRACT|SARCOBATUS VERMICULATUS POLLEN EXTRACT
C1572720|T121|1366957|RXNORM|ENTSUFON|ENTSUFON
C0028368|T125|7518|RXNORM|NORGESTREL|NORGESTREL
C1827410|T121|687342|RXNORM|FENOTEROL / IPRATROPIUM|FENOTEROL / IPRATROPIUM
C2928468|T121|1007547|RXNORM|ASCORBIC ACID / FERROUS FUMARATE / NIACINAMIDE / POLYSACCHARIDE IRON COMPLEX|ASCORBIC ACID / FERROUS FUMARATE / NIACINAMIDE / POLYSACCHARIDE IRON COMPLEX
C0069359|T122|32301|RXNORM|OCTOXYNOL|OCTOXYNOL
C1302135|T121|392575|RXNORM|NYSTATIN / TETRACYCLINE|NYSTATIN / TETRACYCLINE
C1302137|T121|392576|RXNORM|BENDROFLUMETHIAZIDE / POTASSIUM|BENDROFLUMETHIAZIDE / POTASSIUM
C1302130|T121|392570|RXNORM|FUROSEMIDE / TRIAMTERENE|FUROSEMIDE / TRIAMTERENE
C0069787|T121|32658|RXNORM|OXOLAMINE|OXOLAMINE
C0772344|T121|237007|RXNORM|SCOPARIUM|SCOPARIUM
C3700989|T121|1487092|RXNORM|LUFENURON / MILBEMYCIN OXIME / PRAZIQUANTEL|LUFENURON / MILBEMYCIN OXIME / PRAZIQUANTEL
C3644548|T121|1425205|RXNORM|CHOLECALCIFEROL / COD LIVER OIL / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / VITAMIN A|CHOLECALCIFEROL / COD LIVER OIL / DOCOSAHEXAENOATE / EICOSAPENTAENOATE / VITAMIN A
C0041485|T123|10962|RXNORM|TYROSINE|TYROSINE
C0041483|T130|10960|RXNORM|TYROPANOATE|TYROPANOATE
C2937996|T129|1011033|RXNORM|RHUBARB ALLERGENIC EXTRACT|RHUBARB ALLERGENIC EXTRACT
C0041499|T195|10968|RXNORM|TYROTHRICIN|TYROTHRICIN
C3651731|T121|1429953|RXNORM|PULSATILLA KOREANA WHOLE EXTRACT|PULSATILLA KOREANA WHOLE EXTRACT
C3651730|T121|1429955|RXNORM|THEOBROMA CACAO WHOLE EXTRACT|THEOBROMA CACAO WHOLE EXTRACT
C1443664|T121|465370|RXNORM|ATROPINE / PRALIDOXIME|ATROPINE / PRALIDOXIME
C2724931|T121|880374|RXNORM|CHLOPHEDIANOL / PSEUDOEPHEDRINE|CHLOPHEDIANOL / PSEUDOEPHEDRINE
C3813540|T121|1492174|RXNORM|PINEAPPLE EXTRACT|PINEAPPLE EXTRACT
C3818776|T109|1492171|RXNORM|STROPHANTHUS KOMBE WHOLE EXTRACT|STROPHANTHUS KOMBE WHOLE EXTRACT
C0596004|T121|153970|RXNORM|HYOSCYAMINE|HYOSCYAMINE
C2724930|T121|880373|RXNORM|CARBETAPENTANE / GUAIFENESIN / PSEUDOEPHEDRINE|CARBETAPENTANE / GUAIFENESIN / PSEUDOEPHEDRINE
C0055723|T121|21102|RXNORM|CILAZAPRIL|CILAZAPRIL
C2928984|T121|1008075|RXNORM|BENZETHONIUM / BENZOCAINE|BENZETHONIUM / BENZOCAINE
C1876229|T121|1102261|RXNORM|TELAPREVIR|TELAPREVIR
C3819176|T121|1495187|RXNORM|PRAMOXINE / SALICYLOYL PHYTOSPHINGOSINE|PRAMOXINE / SALICYLOYL PHYTOSPHINGOSINE
C3651775|T121|1428838|RXNORM|MELIA AZEDARACH FRUIT EXTRACT|MELIA AZEDARACH FRUIT EXTRACT
C3256085|T121|1363624|RXNORM|PUMMELO EXTRACT|POMELO EXTRACT
C0717517|T121|214323|RXNORM|BROMODIPHENHYDRAMINE / CODEINE|BROMODIPHENHYDRAMINE / CODEINE
C0717518|T121|214324|RXNORM|BROMPHENIRAMINE / PHENYLEPHRINE|BROMPHENIRAMINE / PHENYLEPHRINE
C0717519|T121|214325|RXNORM|BROMPHENIRAMINE / PHENYLPROPANOLAMINE|BROMPHENIRAMINE / PHENYLPROPANOLAMINE
C0057626|T121|22713|RXNORM|DEZOCINE|DEZOCINE
C0717521|T121|214327|RXNORM|BROMPHENIRAMINE / CODEINE / PHENYLPROPANOLAMINE|BROMPHENIRAMINE / CODEINE / PHENYLPROPANOLAMINE
C0001134|T197|236|RXNORM|LAURETH-9|ACIDULATED PHOSPHATE FLUORIDE
C1509940|T121|476786|RXNORM|ALOE POLYSACCHARIDE|ALOE POLYSACCHARIDE
C0073379|T121|35623|RXNORM|RILUZOLE|RILUZOLE
C0017479|T196|4784|RXNORM|GERMANIUM|GERMANIUM
C0991769|T130|317176|RXNORM|ALBUMIN,AGGREGATED|ALBUMIN,AGGREGATED
C0937640|T121|283579|RXNORM|MILK THISTLE EXTRACT|MILK THISTLE EXTRACT
C0982413|T197|314853|RXNORM|STANNOUS CHLORIDE,ANHYDROUS|STANNOUS CHLORIDE,ANHYDROUS
C3256088|T121|1363625|RXNORM|QUATERNIUM-18|QUATERNIUM-18
C2929101|T121|1008194|RXNORM|BENZOCAINE / ZINC SULFATE|BENZOCAINE / ZINC SULFATE
C0033429|T121|8754|RXNORM|PROPAFENONE|PROPAFENONE
C2929103|T121|1008196|RXNORM|CAFFEINE / HORDENINE|CAFFEINE / HORDENINE
C2929104|T121|1008197|RXNORM|CHLORZOXAZONE / KETOPROFEN|CHLORZOXAZONE / KETOPROFEN
C2929097|T121|1008190|RXNORM|DIHYDROXYBUTYL ETHER / SIMETHICONE|DIHYDROXYBUTYL ETHER / SIMETHICONE
C2929098|T121|1008191|RXNORM|FERRIC AMMONIUM CITRATE / FOLIC ACID / VITAMIN B 12|FERRIC AMMONIUM CITRATE / FOLIC ACID / VITAMIN B 12
C2929099|T121|1008192|RXNORM|ATROPINE / HYDROCORTISONE|ATROPINE / HYDROCORTISONE
C2929100|T121|1008193|RXNORM|GLYCOL SALICYLATE / NIACIN / NONIVAMIDE|GLYCOL SALICYLATE / NIACIN / NONIVAMIDE
C0606070|T127|159151|RXNORM|TOCOPHERSOLAN|TOCOFERSOLAN
C0051917|T121|17939|RXNORM|ANIRACETAM|ANIRACETAM
C2929105|T121|1008198|RXNORM|ATENOLOL / CHLORTHALIDONE / HYDRALAZINE|ATENOLOL / CHLORTHALIDONE / HYDRALAZINE
C2929106|T121|1008199|RXNORM|CLOFEXAMIDE / CLOFEZONE|CLOFEXAMIDE / CLOFEZONE
C0248719|T121|73494|RXNORM|TELMISARTAN|TELMISARTAN
C3700399|T121|1551777|RXNORM|NALOXEGOL|NALOXEGOL
C0064009|T123|1423782|RXNORM|ISOMETHYLEUGENOL|ISOMETHYLEUGENOL
C3643351|T121|1423780|RXNORM|C30-50 ALCOHOLS|C30-50 ALCOHOLS
C0675372|T109|1423781|RXNORM|4-ALLYL-2,6-DIMETHOXYPHENOL|4-ALLYL-2,6-DIMETHOXYPHENOL
C3668637|T121|1441186|RXNORM|ISODECYL LAURATE|ISODECYL LAURATE
C0770735|T129|235614|RXNORM|HYMENOPTERA ALLERGENIC EXTRACT|HYMENOPTERA ALLERGENIC EXTRACT
C0057846|T121|22906|RXNORM|DICHLOROBENZYL ALCOHOL|DICHLOROBENZYL ALCOHOL
C0017631|T121|4816|RXNORM|GLICLAZIDE|GLICLAZIDE
C0017628|T121|4815|RXNORM|GLYBURIDE|GLYBURIDE
C3256097|T109|1363627|RXNORM|ASPARAGOPSIS ARMATA EXTRACT|ASPARAGOPSIS ARMATA EXTRACT
C3486394|T121|1340181|RXNORM|SMILAX REGELII ROOT EXTRACT|SMILAX REGELII ROOT EXTRACT
C2929893|T121|1008998|RXNORM|CYSTINE / INOSITOL / RACEMETHIONINE / SODIUM PROPIONATE / UREA|CYSTINE / INOSITOL / RACEMETHIONINE / SODIUM PROPIONATE / UREA
C2929894|T121|1008999|RXNORM|BENZALKONIUM / LIDOCAINE / UREA|BENZALKONIUM / LIDOCAINE / UREA
C0040382|T121|10639|RXNORM|TOLPERISONE|TOLPERISONE
C0040380|T130|10638|RXNORM|TOLONIUM CHLORIDE|TOLONIUM CHLORIDE
C0040379|T121|10637|RXNORM|TOLNAFTATE|TOLNAFTATE
C2929890|T121|1008995|RXNORM|CAMPHOR / EUCALYPTUS OIL / METHYL SALICYLATE|CAMPHOR / EUCALYPTUS OIL / METHYL SALICYLATE
C0040374|T121|10635|RXNORM|TOLBUTAMIDE|TOLBUTAMIDE
C0040374|T121|10635|RXNORM|TOLBUTAMIDE|TOLBUTAMIDE
C2929892|T121|1008997|RXNORM|ANGELICA SINENSIS PREPARATION / BLACK COHOSH EXTRACT|ANGELICA SINENSIS PREPARATION / BLACK COHOSH EXTRACT
C0040372|T121|10633|RXNORM|TOLAZAMIDE|TOLAZAMIDE
C2929886|T121|1008991|RXNORM|AMINOBUTYRATE / PHENOBARBITAL / PHENYTOIN|AMINOBUTYRATE / PHENOBARBITAL / PHENYTOIN
C2929887|T121|1008992|RXNORM|ANTIPYRINE / BENZOCAINE / UREA|ANTIPYRINE / BENZOCAINE / UREA
C2929888|T121|1008993|RXNORM|SHARK LIVER OIL / TISSUE RESPIRATORY FACTOR|SHARK LIVER OIL / TISSUE RESPIRATORY FACTOR
C3645112|T109|1426613|RXNORM|DIETHYLAMINOETHYL-DEXTRAN|DIETHYLAMINOETHYL-DEXTRAN
C3864972|T121|1595783|RXNORM|BENZOCAINE / CAPSAICIN / LIDOCAINE / METHYL SALICYLATE|BENZOCAINE / CAPSAICIN / LIDOCAINE / METHYL SALICYLATE
C2730261|T129|892679|RXNORM|BREWER'S YEAST ALLERGENIC EXTRACT|BREWER'S YEAST ALLERGENIC EXTRACT
C0772133|T121|236816|RXNORM|NEO-HOMOSALATE|NEO-HOMOSALATE
C0052565|T121|18451|RXNORM|ASTAXANTHIN|ASTAXANTHIN
C0136123|T121|54552|RXNORM|PERINDOPRIL|PERINDOPRIL
C3535927|T121|1368279|RXNORM|NEOMYCIN / NYSTATIN / THIOSTREPTON / TRIAMCINOLONE|NEOMYCIN / NYSTATIN / THIOSTREPTON / TRIAMCINOLONE
C2702421|T129|1294632|RXNORM|NORTHERN PAPER WASP VENOM PROTEIN|POLISTES FUSCATUS VENOM
C3486740|T121|1310073|RXNORM|SALIX ALBA FLOWERING TOP EXTRACT|SALIX ALBA FLOWERING TOP EXTRACT
C3485006|T121|1310072|RXNORM|CUSCUTA CHINENSIS SEED EXTRACT|CUSCUTA CHINENSIS SEED EXTRACT
C3485003|T121|1310071|RXNORM|ACONITUM CARMICHAELII ROOT EXTRACT|ACONITUM CARMICHAELII ROOT EXTRACT
C3484830|T109|1310070|RXNORM|BETULA PENDULA TAR OIL|BETULA PENDULA TAR OIL
C3501358|T121|1442981|RXNORM|IBRUTINIB|IBRUTINIB
C0035527|T127|9346|RXNORM|RIBOFLAVIN|RIBOFLAVIN (VIT B2)
C3485007|T121|1310075|RXNORM|DIPSACUS ASPER ROOT EXTRACT|DIPSACUS ASPER ROOT EXTRACT
C0076470|T121|1363062|RXNORM|THIOGLYCEROL|THIOGLYCEROL
C3486752|T121|1310079|RXNORM|LESPEDEZA CAPITATA FLOWERING TOP EXTRACT|LESPEDEZA CAPITATA FLOWERING TOP EXTRACT
C3485011|T121|1310078|RXNORM|JUSTICIA GENDARUSSA LEAF EXTRACT|JUSTICIA GENDARUSSA LEAF EXTRACT
C0772484|T121|237144|RXNORM|THURFYL SALICYLATE|THURFYL SALICYLATE
C0055568|T123|1440856|RXNORM|CHOLIC ACID|CHOLIC ACID
C3695938|T129|1484980|RXNORM|CRESTED DOGSTAIL POLLEN EXTRACT|CYNOSURUS CRISTATUS POLLEN EXTRACT
C3256148|T109|1426611|RXNORM|MODIFIED CORN STARCH (3-E-DOCECENYL SUCCINIC ANHYDRIDE)|MODIFIED CORN STARCH (3-E-DOCECENYL SUCCINIC ANHYDRIDE)
C0070477|T109|33219|RXNORM|PERUVIAN BALSAM|PERUVIAN BALSAM
C1609165|T129|612865|RXNORM|TOCILIZUMAB|TOCILIZUMAB
C2344317|T129|798294|RXNORM|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN P1A[8] VACCINE|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN P1A[8] VACCINE
C3465362|T121|1294638|RXNORM|COMMON PAPER WASP VENOM PROTEIN / METRICUS PAPER WASP VENOM PROTEIN / NORTHERN PAPER WASP VENOM PROTEIN / RED PAPER WASP VENOM PROTEIN|COMMON PAPER WASP VENOM PROTEIN / METRICUS PAPER WASP VENOM PROTEIN / NORTHERN PAPER WASP VENOM PROTEIN / RED PAPER WASP VENOM PROTEIN
C0314977|T007|1150096|RXNORM|BIFIDOBACTERIUM LONGUM|BIFIDOBACTERIUM LONGUM
C1264802|T007|1150094|RXNORM|BIFIDOBACTERIUM LACTIS|BIFIDOBACTERIUM LACTIS
C3205064|T121|1150092|RXNORM|CHROMIUM PICOLINATE / INULIN|CHROMIUM PICOLINATE / INULIN
C0065870|T121|29444|RXNORM|MEFENOREX|MEFENOREX
C2739927|T129|897391|RXNORM|MEXICAN TEA POLLEN EXTRACT|CHENOPODIUM AMBROSIOIDES POLLEN EXTRACT
C3497628|T121|1310299|RXNORM|BOS TAURUS TONSIL PREPARATION|BOVINE TONSIL PREPARATION
C3489092|T121|1310298|RXNORM|BOS TAURUS TESTICLE PREPARATION|BOVINE TESTICLE PREPARATION
C3497627|T121|1310297|RXNORM|BOS TAURUS TENDON PREPARATION|BOVINE TENDON PREPARATION
C3497626|T121|1310296|RXNORM|BOS TAURUS SYMPATHETIC NERVE PREPARATION|BOVINE SYMPATHETIC NERVE PREPARATION
C3486700|T121|1310295|RXNORM|BOS TAURUS SPLEEN PREPARATION|BOVINE SPLEEN PREPARATION
C0038404|T007|10098|RXNORM|ENTEROCOCCUS FAECALIS|ENTEROCOCCUS FAECALIS
C3497624|T121|1310293|RXNORM|BOS TAURUS SOLAR PLEXUS PREPARATION|BOVINE SOLAR PLEXUS PREPARATION
C3497623|T121|1310292|RXNORM|BOS TAURUS RED BLOOD CELL PREPARATION|BOVINE ERYTHROCYTE PREPARATION
C3488236|T121|1310291|RXNORM|BOS TAURUS PITUITARY GLAND PREPARATION|BOVINE PITUITARY GLAND PREPARATION
C3488235|T121|1310290|RXNORM|BOS TAURUS PINEAL GLAND PREPARATION|BOVINE PINEAL GLAND PREPARATION
C0982172|T197|314639|RXNORM|GALLIUM CHLORIDE,GA-67|GALLIUM CHLORIDE,GA-67
C0965618|T121|1091836|RXNORM|ROFLUMILAST|ROFLUMILAST
C0031404|T121|8129|RXNORM|HYDROCORTISONE / NAPHAZOLINE|PHENFORMIN
C0949307|T131|314636|RXNORM|FORMALIN|FORMALIN
C2928889|T121|1007976|RXNORM|DEOXYRIBONUCLEASES / PLASMIN|DEOXYRIBONUCLEASES / PLASMIN
C2928666|T121|1007751|RXNORM|OMEGA-3 ACID ETHYL ESTERS (USP) / PYRIDOXINE / VITAMIN B 12|OMEGA-3 ACID ETHYL ESTERS (USP) / PYRIDOXINE / VITAMIN B 12
C2928665|T121|1007750|RXNORM|GLYCERIN / HYPROMELLOSE / POLYETHYLENE GLYCOL 400 / TETRAHYDROZOLINE / ZINC SULFATE|GLYCERIN / HYPROMELLOSE / POLYETHYLENE GLYCOL 400 / TETRAHYDROZOLINE / ZINC SULFATE
C2928672|T121|1007757|RXNORM|NARATRIPTAN / SUMATRIPTAN|NARATRIPTAN / SUMATRIPTAN
C2928671|T121|1007756|RXNORM|GLYCERIN / HYPROMELLOSE / POLYETHYLENE GLYCOL 400 / TETRAHYDROZOLINE|GLYCERIN / HYPROMELLOSE / POLYETHYLENE GLYCOL 400 / TETRAHYDROZOLINE
C2928669|T121|1007754|RXNORM|DOCUSATE / PIPERAZINE|DOCUSATE / PIPERAZINE
C2928674|T121|1007759|RXNORM|DEXTROMETHORPHAN / GUAIACOLSULFONATE / PHENYLEPHRINE / PYRILAMINE|DEXTROMETHORPHAN / GUAIACOLSULFONATE / PHENYLEPHRINE / PYRILAMINE
C2928673|T121|1007758|RXNORM|LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS SPOROGENES|BACILLUS COAGULANS / LACTOBACILLUS ACIDOPHILUS
C3256155|T109|1426417|RXNORM|DIMETHICONE 1000|DIMETHICONE 1000
C2928891|T121|1007979|RXNORM|CHLORPHENIRAMINE / NOSCAPINE / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / NOSCAPINE / PHENYLPROPANOLAMINE
C2193838|T121|1007978|RXNORM|AMOXICILLIN / SULFINPYRAZONE|AMOXICILLIN / SULFINPYRAZONE
C3256174|T109|1426416|RXNORM|PELVETIA CANALICULATA EXTRACT|CHANNEL WRACK EXTRACT
C2343589|T129|763450|RXNORM|RILONACEPT|RILONACEPT
C3255594|T109|1426411|RXNORM|GLYCERYL STEARATE CITRATE|GLYCERYL STEARATE CITRATE
C2974540|T121|1373458|RXNORM|CANAGLIFLOZIN|CANAGLIFLOZIN
C0982302|T121|1426410|RXNORM|OLETH-2|OLETH-2
C2731559|T129|895574|RXNORM|APRICOT ALLERGENIC EXTRACT|PRUNUS ARMENIACA ALLERGENIC EXTRACT
C0026682|T123|7076|RXNORM|MUCINS|MUCINS
C3256635|T109|1426412|RXNORM|POLYISOBUTYLENE (1100000 MW)|POLYISOBUTYLENE (1200000 MW)
C0066005|T195|29561|RXNORM|MEROPENEM|MEROPENEM
C0051675|T121|17747|RXNORM|AMINOQUINURIDE|AMINOQUINURIDE
C3489017|T121|1311210|RXNORM|SUS SCROFA VEIN PREPARATION|PORCINE VEIN PREPARATION
C3488292|T121|1311212|RXNORM|SUS SCROFA BRAINSTEM PREPARATION|PORCINE BRAINSTEM PREPARATION
C0076080|T121|37776|RXNORM|TEMOZOLOMIDE|TEMOZOLOMIDE
C0076075|T195|37771|RXNORM|TEMAFLOXACIN|TEMAFLOXACIN
C3488293|T121|1311215|RXNORM|SUS SCROFA CEREBRUM PREPARATION|PORCINE BRAIN PREPARATION
C0052796|T195|18631|RXNORM|AZITHROMYCIN|AZITHROMYCIN
C0052796|T195|18631|RXNORM|AZITHROMYCIN|AZITHROMYCIN
C2701206|T130|851985|RXNORM|WESTERN RAGWEED POLLEN EXTRACT|AMBROSIA PSILOSTACHYA POLLEN EXTRACT
C0950387|T121|288262|RXNORM|CINOXATE|CINOXATE
C2701202|T129|851981|RXNORM|DESERT RAGWEED POLLEN EXTRACT|AMBROSIA DUMOSA POLLEN EXTRACT
C0000473|T127|74|RXNORM|NILOTINIB HYDROCHLORIDE|AMINOBENZOIC ACID
C0031469|T121|8163|RXNORM|PHENYLEPHRINE|PHENYLEPHRINE
C0031469|T121|8163|RXNORM|PHENYLEPHRINE|PHENYLEPHRINE
C0031469|T121|8163|RXNORM|PHENYLEPHRINE|PHENYLEPHRINE
C0031469|T121|8163|RXNORM|PHENYLEPHRINE|PHENYLEPHRINE
C0031469|T121|8163|RXNORM|PHENYLEPHRINE|PHENYLEPHRINE
C0031463|T121|8160|RXNORM|PHENYLBUTAZONE|PHENYLBUTAZONE
C0026156|T121|6972|RXNORM|MINERAL OIL|MINERAL OIL
C0026156|T121|6972|RXNORM|MINERAL OIL|MINERAL OIL
C2344313|T129|798290|RXNORM|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G3 VACCINE|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G3 VACCINE
C3474080|T122|1312743|RXNORM|PERFLUOROOCTYL TRIETHOXYSILANE|PERFLUOROOCTYL TRIETHOXYSILANE
C3282850|T122|1312742|RXNORM|POLYACRYLAMIDE (1500 MW)|POLYACRYLAMIDE (1500 MW)
C0068517|T121|1312741|RXNORM|NEOHESPERIDIN DIHYDROCHALCONE|NEOHESPERIDIN DIHYDROCHALCONE
C3465041|T121|1312740|RXNORM|SILANETRIOL|SILANETRIOL
C0939882|T121|285228|RXNORM|KAVA PREPARATION|KAVA
C3669202|T121|1485066|RXNORM|LYCOPODIUM CLAVATUM WHOLE EXTRACT|LYCOPODIUM CLAVATUM WHOLE EXTRACT
C3695932|T121|1485065|RXNORM|COLCHICUM AUTUMNALE SEED EXTRACT|COLCHICUM AUTUMNALE SEED EXTRACT
C3669153|T121|1485064|RXNORM|BAMBUSA BAMBOS WHOLE EXTRACT|BAMBUSA BAMBOS WHOLE EXTRACT
C3490290|T116|1591894|RXNORM|ADVANTAME|ADVANTAME
C1143528|T109|1314360|RXNORM|ETHYL NITRATE|ETHYL NITRATE
C3159402|T121|1111077|RXNORM|METHYL SALICYLATE / TURPENTINE|METHYL SALICYLATE / TURPENTINE
C0006388|T121|1813|RXNORM|LEVOBUNOLOL|LEVOBUNOLOL
C1445421|T129|466192|RXNORM|ASPERGILLUS FUMIGATUS EXTRACT|ASPERGILLUS FUMIGATUS EXTRACT
C1313052|T121|1490468|RXNORM|TASIMELTEON|TASIMELTEON
C1445426|T129|466197|RXNORM|CHAETOMIUM GLOBOSUM EXTRACT|CHAETOMIUM GLOBOSUM EXTRACT
C1445427|T129|466198|RXNORM|CLADOSPORIUM HERBARUM EXTRACT|CLADOSPORIUM HERBARUM EXTRACT
C3485054|T121|1314595|RXNORM|AGRIMONIA EUPATORIA EXTRACT|AGRIMONIA EUPATORIA EXTRACT
C3256803|T121|1314596|RXNORM|PREZATIDE COPPER ACETATE|PREZATIDE COPPER ACETATE
C0939869|T121|1314597|RXNORM|ROSEMARY EXTRACT|ROSEMARY EXTRACT
C3502538|T109|1420141|RXNORM|LYRAL|LYRAL
C2726173|T129|1314591|RXNORM|JUNIPERUS VIRGINIANA ALLERGENIC EXTRACT|JUNIPERUS VIRGINIANA ALLERGENIC EXTRACT
C2726217|T129|1314592|RXNORM|STREPTOMYCES GRISEUS ALLERGENIC EXTRACT|STREPTOMYCES GRISEUS ALLERGENIC EXTRACT
C0029923|T123|1314593|RXNORM|OVALBUMIN|OVALBUMIN
C3255752|T121|1312568|RXNORM|ETHYL 2-METHYLBUTYRATE|ETHYL 2-METHYLBUTYRATE
C0068946|T109|1591892|RXNORM|N-NONYLPHENOL|NONYLPHENOL
C0717874|T121|214665|RXNORM|KAOLIN / PECTIN|KAOLIN / PECTIN
C0717873|T121|214664|RXNORM|ISOPROTERENOL / PHENYLEPHRINE|ISOPROTERENOL / PHENYLEPHRINE
C3267311|T121|1312560|RXNORM|DISTEARYL PHTHALAMIC ACID|DISTEARYL PHTHALAMIC ACID
C3643363|T109|1421547|RXNORM|PEG-9 DIGLYCIDYL ETHER AND SODIUM HYALURONATE CROSS POLYMER|PEG-9 DIGLYCIDYL ETHER AND SODIUM HYALURONATE CROSS POLYMER
C0717871|T121|214662|RXNORM|ISONIAZID / PYRAZINAMIDE / RIFAMPIN|ISONIAZID / PYRAZINAMIDE / RIFAMPIN
C2080475|T121|817824|RXNORM|ACETAMINOPHEN / ASCORBIC ACID / PHENYLEPHRINE|ACETAMINOPHEN / ASCORBIC ACID / PHENYLEPHRINE
C0303232|T197|1545043|RXNORM|LEAD CARBONATE|LEAD CARBONATE
C2929111|T121|1008204|RXNORM|PRIDINOL / ROFECOXIB|PRIDINOL / ROFECOXIB
C2929112|T121|1008205|RXNORM|HYDROCHLOROTHIAZIDE / MAGNESIUM CHLORIDE / METHOTRIMEPRAZINE|HYDROCHLOROTHIAZIDE / MAGNESIUM CHLORIDE / METHOTRIMEPRAZINE
C2929113|T121|1008206|RXNORM|ACTIVATED CHARCOAL / PAPAVERINE|ACTIVATED CHARCOAL / PAPAVERINE
C2929114|T121|1008207|RXNORM|CAFFEINE / ETHENZAMIDE|CAFFEINE / ETHENZAMIDE
C2929107|T121|1008200|RXNORM|MENTHOL / SIMETHICONE|MENTHOL / SIMETHICONE
C2929108|T121|1008201|RXNORM|BETA-ALANINE / OXAZEPAM|BETA-ALANINE / OXAZEPAM
C2929109|T121|1008202|RXNORM|CALCIUM LACTATE / MAGNESIUM OXIDE|CALCIUM LACTATE / MAGNESIUM OXIDE
C2929110|T121|1008203|RXNORM|CARNITINE / RACEMETHIONINE / THIAMINE|CARNITINE / RACEMETHIONINE / THIAMINE
C0022478|T126|6095|RXNORM|KININOGENASE|KININOGENASE
C0015980|T129|4381|RXNORM|INTERFERON-BETA|INTERFERON BETA NATURAL
C3848599|T121|1545041|RXNORM|OVIS ARIES TESTICLE PREPARATION|OVIS ARIES TESTICLE PREPARATION
C2929115|T121|1008208|RXNORM|METOLAZONE / TRIAMTERENE|METOLAZONE / TRIAMTERENE
C2929116|T121|1008209|RXNORM|AMILORIDE / TRICHLORMETHIAZIDE|AMILORIDE / TRICHLORMETHIAZIDE
C0016006|T123|4385|RXNORM|FIBRINOGEN|FIBRINOGEN
C3505162|T121|1357999|RXNORM|AMARANTHUS VIRIDIS LEAF EXTRACT|AMARANTHUS VIRIDIS LEAF EXTRACT
C0379135|T123|115238|RXNORM|BECAPLERMIN|BECAPLERMIN
C0005013|T121|1373|RXNORM|BENPERIDOL|BENPERIDOL
C0005011|T121|1372|RXNORM|BENORILATE|BENORILATE
C0005018|T197|1375|RXNORM|BENTONITE|BENTONITE
C0005014|T121|1374|RXNORM|BENSERAZIDE|BENSERAZIDE
C0018488|T196|1534767|RXNORM|HAFNIUM|HAFNIUM
C1095916|T121|319837|RXNORM|GOTU KOLA EXTRACT|GOTU KOLA EXTRACT
C2183092|T121|812544|RXNORM|BROMHEXINE / DEXTROMETHORPHAN|BROMHEXINE / DEXTROMETHORPHAN
C0005025|T121|1378|RXNORM|BENZALKONIUM|BENZALKONIUM
C0005025|T121|1378|RXNORM|BENZALKONIUM|BENZALKONIUM
C2183764|T121|817157|RXNORM|DIPYRONE / PAPAVERINE|DIPYRONE / PAPAVERINE
C3505160|T109|1357997|RXNORM|CURED FAT, PORK SIDE BACON|CURED FAT, PORK SIDE BACON
C0717606|T121|214409|RXNORM|CHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE|CHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE
C1827991|T121|818629|RXNORM|BISMUTH BISKALCITRATE / METRONIDAZOLE / TETRACYCLINE|BISMUTH BISKALCITRATE / METRONIDAZOLE / TETRACYCLINE
C2701625|T129|852526|RXNORM|BURROBRUSH POLLEN EXTRACT|HYMENOCLEA SALSOLA POLLEN EXTRACT
C0055153|T109|1368150|RXNORM|CETYL LACTATE|CETYL LACTATE
C0717604|T121|214407|RXNORM|CHLORPHENIRAMINE / GUAIFENESIN / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / GUAIFENESIN / PSEUDOEPHEDRINE
C0717603|T121|214406|RXNORM|CHLORPHENIRAMINE / GUAIFENESIN / PHENYLEPHRINE|CHLORPHENIRAMINE / GUAIFENESIN / PHENYLEPHRINE
C1720375|T121|646781|RXNORM|BENZOYL PEROXIDE / CLINDAMYCIN|BENZOYL PEROXIDE / CLINDAMYCIN
C2929254|T121|1008349|RXNORM|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE|DEXBROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE
C2929253|T121|1008348|RXNORM|ASTEMIZOLE / CLORAZEPATE|ASTEMIZOLE / CLORAZEPATE
C0043375|T123|11378|RXNORM|XYLOSE|XYLOSE
C2929246|T121|1008341|RXNORM|FUSIDATE / HYDROCORTISONE|FUSIDATE / HYDROCORTISONE
C2929245|T121|1008340|RXNORM|DOCUSATE / SENNOSIDES, USP|DOCUSATE / SENNOSIDES, USP
C2929245|T121|1008340|RXNORM|DOCUSATE / SENNOSIDES, USP|DOCUSATE / SENNOSIDES, USP
C0043369|T121|11377|RXNORM|XYLITOL|XYLITOL
C2929247|T121|1008342|RXNORM|LAURETH-9 / OLEATE|OLEATE / POLIDOCANOL
C2929250|T121|1008345|RXNORM|GAMMA-LINOLENATE / LINOLEATE|GAMMA-LINOLENATE / LINOLEATE
C2929249|T121|1008344|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 14 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 18C CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 19F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 23F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 4 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 6B CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 9V CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 14 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 18C CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 19F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 23F CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 4 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 6B CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE / STREPTOCOCCUS PNEUMONIAE SEROTYPE 9V CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C2929252|T121|1008347|RXNORM|FUROSEMIDE / PENBUTOLOL|FUROSEMIDE / PENBUTOLOL
C2929251|T121|1008346|RXNORM|THIAMINE / THIOCTATE|THIAMINE / THIOCTATE
C3255876|T109|1307083|RXNORM|STEARYL ETHYLHEXANOATE|STEARYL ETHYLHEXANOATE
C0772202|T121|1307080|RXNORM|CYCLOMETHICONE|CYCLOMETHICONE
C3256217|T109|1307081|RXNORM|CYCLOMETHICONE 6|CYCLOMETHICONE 6
C3256083|T109|1307086|RXNORM|PEG-9 STEARATE|PEG-9 STEARATE
C3256600|T109|1307087|RXNORM|CAESALPINIA SPINOSA RESIN|CAESALPINIA SPINOSA RESIN
C3268186|T121|1307085|RXNORM|2-(4-(DIETHYLAMINO)-2-HYDROXYBENZOYL)BENZOIC ACID|2-(4-(DIETHYLAMINO)-2-HYDROXYBENZOYL)BENZOIC ACID
C0138045|T121|55024|RXNORM|POTASSIUM TARTRATE|POTASSIUM TARTRATE
C3256624|T109|1307088|RXNORM|ISOTRIDECYL ISONONANOATE|ISOTRIDECYL ISONONANOATE
C0069647|T121|32533|RXNORM|ORMETOPRIM|ORMETOPRIM
C0053396|T127|19143|RXNORM|BETA CAROTENE|BETA CAROTENE
C0053396|T127|19143|RXNORM|BETA CAROTENE|BETA CAROTENE
C3538266|T121|1372466|RXNORM|HIBISCUS SYRIACUS SEED EXTRACT|HIBISCUS SYRIACUS SEED EXTRACT
C0939871|T121|285219|RXNORM|APIS MELLIFERA PREPARATION|APIS MELLIFERA PREPARATION
C2242156|T129|763096|RXNORM|POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY)|POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY)
C2194291|T121|812663|RXNORM|PIPENZOLATE / SIMETHICONE|PIPENZOLATE / SIMETHICONE
C0991776|T129|999438|RXNORM|CURVULARIA INEQUALIS ALLERGENIC EXTRACT|CURVULARIA INEQUALIS ALLERGENIC EXTRACT
C2142868|T121|814512|RXNORM|DEXBROMPHENIRAMINE / GUAIFENESIN / PSEUDOEPHEDRINE|DEXBROMPHENIRAMINE / GUAIFENESIN / PSEUDOEPHEDRINE
C1959893|T121|729536|RXNORM|DYDROGESTERONE / ESTRADIOL|DYDROGESTERONE / ESTRADIOL
C2073821|T121|815844|RXNORM|CHLORCYCLIZINE / PSEUDOEPHEDRINE|CHLORCYCLIZINE / PSEUDOEPHEDRINE
C3504693|T121|1356480|RXNORM|LUFFA OPERCULATA WHOLE EXTRACT|LUFFA OPERCULATA WHOLE EXTRACT
C3504694|T121|1356481|RXNORM|2-PROPOXY-1-PROPANOL|2-PROPOXY-1-PROPANOL
C3504695|T121|1356482|RXNORM|ACTINIDIA CHINENSIS WHOLE EXTRACT|ACTINIDIA CHINENSIS WHOLE EXTRACT
C3504696|T121|1356483|RXNORM|ISOPROPYL BEHENATE|ISOPROPYL BEHENATE
C0620926|T121|1356484|RXNORM|PANTHENYL ETHYL ETHER|PANTHENYL ETHYL ETHER
C0717754|T121|214551|RXNORM|ESTRADIOL / NORETHINDRONE|ESTRADIOL / NORETHINDRONE
C0009148|T196|1310300|RXNORM|COBALT|COBALT
C2709756|T129|854952|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 20 VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 20 VACCINE
C3255593|T121|1307262|RXNORM|GLYCERYL LINOLENATE|GLYCERYL LINOLENATE
C3256524|T121|1307263|RXNORM|DISTEARYL ETHER|DISTEARYL ETHER
C3256001|T109|1367169|RXNORM|HYDROXYOCTACOSANYL HYDROXYSTEARATE|HYDROXYOCTACOSANYL HYDROXYSTEARATE
C0917147|T121|1492341|RXNORM|EQUOL, (+-)-|EQUOL, (+-)-
C3815502|T121|1492439|RXNORM|SYMPHYTUM OFFICINALE WHOLE EXTRACT|SYMPHYTUM OFFICINALE WHOLE EXTRACT
C0770228|T125|235282|RXNORM|ULTRALENTE INSULIN, BEEF|ULTRALENTE INSULIN, BEEF
C0770230|T125|235283|RXNORM|INSULIN, PROMPT ZINC, BEEF-PORK|INSULIN, PROMPT ZINC, BEEF-PORK
C0770221|T125|235280|RXNORM|LENTE INSULIN, BEEF|LENTE INSULIN, BEEF
C0770226|T125|235281|RXNORM|ULTRALENTE INSULIN, BEEF-PORK|ULTRALENTE INSULIN, BEEF-PORK
C0770234|T125|235286|RXNORM|INSULIN, PROMPT ZINC, PORK|INSULIN, PROMPT ZINC, PORK
C0770232|T125|235284|RXNORM|INSULIN, PROMPT ZINC, BEEF|INSULIN, PROMPT ZINC, BEEF
C0770233|T125|235285|RXNORM|INSULIN, PROMPT ZINC, HUMAN|INSULIN, PROMPT ZINC, HUMAN
C0060502|T121|25121|RXNORM|FLUNIXIN|FLUNIXIN
C0060501|T121|25120|RXNORM|FLUNISOLIDE|FLUNISOLIDE
C0060501|T121|25120|RXNORM|FLUNISOLIDE|FLUNISOLIDE
C0060508|T121|25127|RXNORM|FLUOCORTIN BUTYL ESTER|FLUOCORTIN BUTYL ESTER
C0060507|T121|25126|RXNORM|FLUOCINOLONE|FLUOCINOLONE
C0060507|T121|25126|RXNORM|FLUOCINOLONE|FLUOCINOLONE
C0060507|T121|25126|RXNORM|FLUOCINOLONE|FLUOCINOLONE
C0060879|T195|25437|RXNORM|FUSAFUNGIN|FUSAFUNGIN
C0069763|T121|1009342|RXNORM|OXIBENDAZOLE|OXIBENDAZOLE
C1721498|T121|1102188|RXNORM|FERROUS BISGLYCINATE|FERROUS BISGLYCINATE
C1636671|T121|608838|RXNORM|DROSPIRENONE / ESTRADIOL|DROSPIRENONE / ESTRADIOL
C1641847|T121|608835|RXNORM|AMMONIUM CHLORIDE / DIPHENHYDRAMINE|AMMONIUM CHLORIDE / DIPHENHYDRAMINE
C2929735|T121|1008837|RXNORM|HEPATITIS A VACCINE (INACTIVATED) STRAIN HM175 / HEPATITIS B SURFACE ANTIGEN VACCINE|HEPATITIS A VACCINE (INACTIVATED) STRAIN HM175 / HEPATITIS B SURFACE ANTIGEN VACCINE
C2929734|T121|1008836|RXNORM|GUAIFENESIN / PHENYLEPHRINE / PSEUDOEPHEDRINE|GUAIFENESIN / PHENYLEPHRINE / PSEUDOEPHEDRINE
C2929733|T121|1008835|RXNORM|VITAMIN E / ZINC CITRATE|VITAMIN E / ZINC CITRATE
C2929732|T121|1008834|RXNORM|BENZOCAINE / NITROFURAZONE / TYROTHRICIN|BENZOCAINE / NITROFURAZONE / TYROTHRICIN
C2929731|T121|1008833|RXNORM|BUZEPIDE METIODIDE / CLOCINIZINE / PHENYLPROPANOLAMINE|BUZEPIDE METIODIDE / CLOCINIZINE / PHENYLPROPANOLAMINE
C2929730|T121|1008832|RXNORM|ASPIRIN / SULFUR|ASPIRIN / SULFUR
C2929729|T121|1008831|RXNORM|CALCIUM LACTATE / MAGNESIUM CITRATE|CALCIUM LACTATE / MAGNESIUM CITRATE
C2929728|T121|1008830|RXNORM|ITRACONAZOLE / SECNIDAZOLE|ITRACONAZOLE / SECNIDAZOLE
C3474136|T121|1358886|RXNORM|ZANTHOXYLUM SCHINIFOLIUM WHOLE EXTRACT|ZANTHOXYLUM SCHINIFOLIUM WHOLE EXTRACT
C3475119|T109|1358887|RXNORM|EUONYMUS ALATUS WHOLE EXTRACT|EUONYMUS ALATUS WHOLE EXTRACT
C2929737|T121|1008839|RXNORM|DIMETHICONE / LANOLIN|DIMETHICONE / LANOLIN
C2929736|T121|1008838|RXNORM|GREEN TEA EXTRACT / GREEN TEA LEAF EXTRACT|GREEN TEA EXTRACT / GREEN TEA LEAF EXTRACT
C2962887|T121|1087329|RXNORM|ALPHA TOCOPHEROL / FOLIC ACID / HYDROXOCOBALAMIN / MAGNESIUM OXIDE / PYRIDOXINE|ALPHA TOCOPHEROL / FOLIC ACID / HYDROXOCOBALAMIN / MAGNESIUM OXIDE / PYRIDOXINE
C0671970|T121|194000|RXNORM|CAPECITABINE|CAPECITABINE
C0001050|T121|199|RXNORM|ACETYLDIGOXINS|ACETYLDIGOXINS
C2928553|T121|1007637|RXNORM|PHENYLEPHRINE / WITCH HAZEL|PHENYLEPHRINE / WITCH HAZEL
C3818772|T121|1492299|RXNORM|LOLIUM TEMULENTUM TOP EXTRACT|LOLIUM TEMULENTUM TOP EXTRACT
C2930017|T121|1009122|RXNORM|BETAMETHASONE / MAGNESIUM TRISILICATE|BETAMETHASONE / MAGNESIUM TRISILICATE
C2930018|T121|1009123|RXNORM|ACETAMINOPHEN / DOMPERIDONE|ACETAMINOPHEN / DOMPERIDONE
C2930015|T121|1009120|RXNORM|HOMATROPINE / IODOQUINOL / PHTHALYLSULFACETAMIDE|HOMATROPINE / IODOQUINOL / PHTHALYLSULFACETAMIDE
C2930016|T121|1009121|RXNORM|CALCIUM CARBONATE / PHENYTOIN|CALCIUM CARBONATE / PHENYTOIN
C2930021|T121|1009126|RXNORM|ANTHRAQUINONE GLYCOSIDE / SALICYLIC ACID|ANTHRAQUINONE GLYCOSIDE / SALICYLIC ACID
C2930022|T121|1009127|RXNORM|ANTHRALIN / COAL TAR / SALICYLIC ACID|ANTHRALIN / COAL TAR / SALICYLIC ACID
C2930019|T121|1009124|RXNORM|ASCORBIC ACID / COLLAGEN, HYDROLYZED|ASCORBIC ACID / COLLAGEN, HYDROLYZED
C2930020|T121|1009125|RXNORM|BENZALKONIUM / DIMETHICONE|BENZALKONIUM / DIMETHICONE
C2930023|T121|1009128|RXNORM|CAFFEINE / ERGOTAMINE / IBUPROFEN|CAFFEINE / ERGOTAMINE / IBUPROFEN
C2930024|T121|1009129|RXNORM|MECOBALAMIN / VITAMIN B 12|MECOBALAMIN / VITAMIN B 12
C0001044|T126|195|RXNORM|ACETYLCHOLINESTERASE|ACETYLCHOLINESTERASE
C3538468|T121|1372889|RXNORM|HYDROCORTISONE / PHENOL|HYDROCORTISONE / PHENOL
C3819167|T121|1494975|RXNORM|BISHYDROXYETHYL DIHYDROXYPROPYL STEARAMMONIUM|BISHYDROXYETHYL DIHYDROXYPROPYL STEARAMMONIUM
C3488906|T121|1309799|RXNORM|LIGUSTICUM PORTERI ROOT EXTRACT|LIGUSTICUM PORTERI ROOT EXTRACT
C1966236|T121|745510|RXNORM|CARBETAPENTANE / PYRILAMINE|CARBETAPENTANE / PYRILAMINE
C3255715|T121|1372259|RXNORM|PICEA ABIES WOOD EXTRACT|PICEA ABIES WOOD EXTRACT
C0039663|T121|10402|RXNORM|TETRAHYDROCANNABINOL|TETRAHYDROCANNABINOL
C1875271|T121|689930|RXNORM|HYDROGEN PEROXIDE / SODIUM BICARBONATE|HYDROGEN PEROXIDE / SODIUM BICARBONATE
C0038633|T121|10156|RXNORM|SUCRALFATE|SUCRALFATE
C0038627|T121|10154|RXNORM|SUCCINYLCHOLINE|SUCCINYLCHOLINE
C3818706|T109|1535514|RXNORM|DIPHENYL DIMETHICONE (100 CST)|DIPHENYL DIMETHICONE (100 CST)
C1874783|T121|689289|RXNORM|CHLORCYCLIZINE / HYDROCORTISONE|CHLORCYCLIZINE / HYDROCORTISONE
C1874782|T121|689288|RXNORM|CHLORAMPHENICOL / HYDROCORTISONE / POLYMYXIN B|CHLORAMPHENICOL / HYDROCORTISONE / POLYMYXIN B
C0038636|T123|10159|RXNORM|SUCROSE|SUCROSE
C0225326|T121|70727|RXNORM|FIBER|FIBER
C0982140|T121|314611|RXNORM|ETHYL DIHYDROXYPROPYL PABA|ETHYL DIHYDROXYPROPYL PABA
C0771017|T121|235829|RXNORM|METHOSERPIDINE|METHOSERPIDINE
C2702422|T129|1294628|RXNORM|COMMON PAPER WASP VENOM PROTEIN|POLISTES EXCLAMANS VENOM
C3535623|T121|1370734|RXNORM|TOXICODENDRON PUBESCENS SHOOT EXTRACT|EASTERN POISON OAK SHOOT EXTRACT
C3535625|T121|1370732|RXNORM|SODIUM LAUROYL 1-METHYL ISETHIONATE|SODIUM LAUROYL 1-METHYL ISETHIONATE
C3535624|T121|1370733|RXNORM|TRIMETHYLSILOXYSILICATE (M-Q 1.0-1.2)|TRIMETHYLSILOXYSILICATE (M-Q 1.0-1.2)
C3535626|T109|1370731|RXNORM|POLYGLYCERYL-3 OLEATE|POLYGLYCERYL-3 OLEATE
C0069715|T130|1427058|RXNORM|OXALIC ACID|OXALIC ACID
C1165733|T129|1427059|RXNORM|LOLIUM PERENNE ALLERGENIC EXTRACT|PERENNIAL RYEGRASS ALLERGENIC EXTRACT
C0036534|T125|9627|RXNORM|SECRETIN|SECRETIN
C0036516|T121|9624|RXNORM|SECOBARBITAL|SECOBARBITAL
C2701542|T129|852367|RXNORM|RUSSIAN OLIVE POLLEN EXTRACT|OLEASTER POLLEN EXTRACT
C0001134|T197|236|RXNORM|ROSE HIPS|ACIDULATED PHOSPHATE FLUORIDE
C0772035|T121|236730|RXNORM|SIMALDRATE|SIMALDRATE
C0772041|T129|236736|RXNORM|TICK-BORN ENCEPHALITIS VACC|TICK-BORN ENCEPHALITIS VACC
C0020274|T197|5496|RXNORM|HYDROFLUORIC ACID|HYDROFLUORIC ACID
C0056480|T121|21732|RXNORM|CRESATIN|CRESATIN
C0056480|T121|21732|RXNORM|CRESATIN|CRESATIN
C0056480|T121|21732|RXNORM|CRESATIN|CRESATIN
C0053067|T121|18846|RXNORM|BECLAMIDE|BECLAMIDE
C0006865|T121|1976|RXNORM|CANNABINOL|CANNABINOL
C2222738|T121|1117535|RXNORM|POTASSIUM NITRATE / SILVER NITRATE|POTASSIUM NITRATE / SILVER NITRATE
C3692231|T121|1441534|RXNORM|POLYETHYLENE GLYCOL 900000|POLYETHYLENE GLYCOL 900000
C3692233|T121|1441536|RXNORM|ALLIUM SATIVUM WHOLE EXTRACT|ALLIUM SATIVUM WHOLE EXTRACT
C3651717|T121|1431147|RXNORM|DECYL JOJOBATE|DECYL JOJOBATE
C2722050|T129|891687|RXNORM|ENGLISH WALNUT ALLERGENIC EXTRACT|JUGLANS REGIA ALLERGENIC EXTRACT
C3651715|T121|1431149|RXNORM|METHYL PERFLUOROISOBUTYL ETHER|METHYL PERFLUOROISOBUTYL ETHER
C3651716|T121|1431148|RXNORM|METHYL PERFLUOROBUTYL ETHER|METHYL PERFLUOROBUTYL ETHER
C1827393|T121|687104|RXNORM|BENZOCAINE / DEQUALINIUM|BENZOCAINE / DEQUALINIUM
C3819180|T121|1491617|RXNORM|CALCIUM CARBONATE / MAGNESIUM OXIDE / ZINC OXIDE|CALCIUM CARBONATE / MAGNESIUM OXIDE / ZINC OXIDE
C3256388|T121|1314293|RXNORM|TRIMETHOXYCAPRYLYLSILANE|TRIMETHOXYCAPRYLYLSILANE
C3256386|T109|1314292|RXNORM|TRIHYDROXYPALMITAMIDOHYDROXYPROPYL MYRISTYL ETHER|TRIHYDROXYPALMITAMIDOHYDROXYPROPYL MYRISTYL ETHER
C3256288|T121|1314291|RXNORM|MAGNESIUM ALUMINOMETASILICATE TYPE I-B|MAGNESIUM ALUMINOMETASILICATE TYPE I-B
C3256222|T121|1314290|RXNORM|DIMETHICONOL (250000 MW)|DIMETHICONOL (250000 MW)
C3256643|T121|1314297|RXNORM|POLYQUATERNIUM-7 (70-30 ACRYLAMIDE-DADMAC; 900 KD)|POLYQUATERNIUM-7 (70-30 ACRYLAMIDE-DADMAC; 900 KD)
C3256563|T121|1314296|RXNORM|TETRAPEPTIDE-21|TETRAPEPTIDE-21
C3256453|T109|1314295|RXNORM|TRIMETHYLOLPROPANE TRIETHYLHEXANOATE|TRIMETHYLOLPROPANE TRIETHYLHEXANOATE
C3256452|T109|1314294|RXNORM|TRIMETHYLOLPROPANE TRICAPRATE|TRIMETHYLOLPROPANE TRICAPRATE
C3256682|T109|1314299|RXNORM|GARDEN LADY'S MANTLE EXTRACT|GARDEN LADY'S MANTLE EXTRACT
C1656494|T109|1547632|RXNORM|SODIUM DIACETATE|SODIUM DIACETATE
C2927565|T129|1006340|RXNORM|CAYENNE PEPPER ALLERGENIC EXTRACT|CAYENNE PEPPER ALLERGENIC EXTRACT
C3486323|T109|1305648|RXNORM|AZADIRACHTA INDICA SEED OIL|AZADIRACHTA INDICA SEED OIL
C2346950|T168|1305649|RXNORM|BABASSU OIL|BABASSU OIL
C2194026|T121|812357|RXNORM|MAGNESIUM SULFATE / PEPTONES|MAGNESIUM SULFATE / PEPTONES
C3834236|T121|1543748|RXNORM|CAPSAICIN / HISTAMINE|CAPSAICIN / HISTAMINE
C2975054|T168|1305642|RXNORM|ARGAN OIL|ARGAN OIL
C2980709|T109|1305643|RXNORM|ATRACTYLODES JAPONICA ROOT OIL|ATRACTYLODES LANCEA ROOT OIL
C3256343|T109|1305640|RXNORM|ANGELICA ROOT OIL|ANGELICA ROOT OIL
C3473403|T109|1305641|RXNORM|ANGELICA SEED OIL|ANGELICA SEED OIL
C3256185|T121|1372262|RXNORM|SNOW PEA EXTRACT|SNOW PEA EXTRACT
C3256274|T121|1372263|RXNORM|SALICORNIA EUROPAEA EXTRACT|GLASSWORT EXTRACT
C1875791|T121|690740|RXNORM|SULFACETAMIDE / SULFUR|SULFACETAMIDE / SULFUR
C1875791|T121|690740|RXNORM|SULFACETAMIDE / SULFUR|SULFACETAMIDE / SULFUR
C1875792|T121|690741|RXNORM|SULFADIAZINE / SULFAMERAZINE / SULFAMETHAZINE|SULFADIAZINE / SULFAMERAZINE / SULFAMETHAZINE
C3644496|T122|1425089|RXNORM|POLAWAX POLYSORBATE|POLAWAX POLYSORBATE
C3854051|T121|1592735|RXNORM|PHAEODACTYLUM TRICORNUTUM|PHAEODACTYLUM TRICORNUTUM EXTRACT
C2930789|T121|1592737|RXNORM|NINTEDANIB|NINTEDANIB
C3859335|T121|1592733|RXNORM|CLOVE OIL / EUCALYPTUS OIL / MENTHOL|CLOVE OIL / EUCALYPTUS OIL / MENTHOL
C0612470|T121|163406|RXNORM|DIFEMERINE|DIFEMERINE
C0010137|T125|2878|RXNORM|CORTISONE|CORTISONE
C2194089|T121|814417|RXNORM|METOCLOPRAMIDE / PANCREATIN / SIMETHICONE|METOCLOPRAMIDE / PANCREATIN / SIMETHICONE
C0360470|T121|108038|RXNORM|ACETAMINOPHEN / CAFFEINE|ACETAMINOPHEN / CAFFEINE
C0012093|T195|3356|RXNORM|DICLOXACILLIN|DICLOXACILLIN
C0012082|T121|3351|RXNORM|DICHLOROPHEN|DICHLOROPHEN
C0012081|T121|3350|RXNORM|CLODRONIC ACID|CLODRONIC ACID
C0012086|T121|3353|RXNORM|DICHLORPHENAMIDE|DICLOFENAMIDE
C3528056|T109|1361658|RXNORM|PHENOXYETHYL CAPRYLATE|PHENOXYETHYL CAPRYLATE
C3495673|T196|1361657|RXNORM|IODIDE ION I-123|IODIDE ION I-123
C0163981|T122|1361656|RXNORM|PROPYLENE GLYCOL ALGINATE ESTER|PROPYLENE GLYCOL ALGINATE ESTER
C3528055|T109|1361655|RXNORM|HYDROXYPROPYL GUAR (2500-4500 MPA.S AT 1%)|HYDROXYPROPYL GUAR (2500-4500 MPA.S AT 1%)
C3528054|T121|1361654|RXNORM|ETHYLENEDIAMINE TETRAETHANOL|ETHYLENEDIAMINE TETRAETHANOL
C3256016|T121|1307864|RXNORM|ALTHAEA OFFICINALIS LEAF EXTRACT|ALTHAEA OFFICINALIS LEAF EXTRACT
C1879704|T121|1307866|RXNORM|ANGELICA SINENSIS ROOT EXTRACT|ANGELICA SINENSIS ROOT EXTRACT
C3709688|T121|1488055|RXNORM|DIHEPTYL SUCCINATE|DIHEPTYL SUCCINATE
C3709687|T121|1488054|RXNORM|CETYL HYDROXYETHYLCELLULOSE (550000 MW)|CETYL HYDROXYETHYLCELLULOSE (550000 MW)
C0054480|T121|20063|RXNORM|CALCIUM POLYCARBOPHIL|CALCIUM POLYCARBOPHIL
C0054480|T121|20063|RXNORM|CALCIUM POLYCARBOPHIL|CALCIUM POLYCARBOPHIL
C3255904|T109|1307863|RXNORM|KUKUI NUT EXTRACT|ALEURITES MOLUCCANA SEED EXTRACT
C2146602|T121|813990|RXNORM|ACETAMINOPHEN / CINNAMEDRINE / PAMABROM / PYRILAMINE|ACETAMINOPHEN / CINNAMEDRINE / PAMABROM / PYRILAMINE
C0768119|T121|234416|RXNORM|LANTHANUM CARBONATE|LANTHANUM CARBONATE
C3864833|T121|1596929|RXNORM|ETHYLHEXYL GALLATE|ETHYLHEXYL GALLATE
C3499444|T121|1312086|RXNORM|TRIETHANOLAMINE LACTATE|TEA-LACTATE
C1874934|T121|690296|RXNORM|CRESOL / FORMALDEHYDE|CRESOL / FORMALDEHYDE
C2344311|T129|798288|RXNORM|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G2 VACCINE|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G2 VACCINE
C0008803|T121|2549|RXNORM|CINNARIZINE|CINNARIZINE
C2344309|T129|798286|RXNORM|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G1 VACCINE|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G1 VACCINE
C3486738|T121|1311404|RXNORM|LARIX DECIDUA RESIN EXTRACT|LARIX DECIDUA RESIN
C0982182|T121|1311155|RXNORM|GLYCERYL STEARATE|GLYCERYL STEARATE
C3486862|T121|1311154|RXNORM|PULSATILLA PATENS EXTRACT|PULSATILLA PATENS EXTRACT
C2928521|T121|1007603|RXNORM|CAFFEINE / ERGOTAMINE / LEVOROTATORY ALKALOIDS OF BELLADONNA / PENTOBARBITAL|CAFFEINE / ERGOTAMINE / LEVOROTATORY ALKALOIDS OF BELLADONNA / PENTOBARBITAL
C1095899|T121|1311152|RXNORM|HYOSCYAMUS NIGER EXTRACT|HYOSCYAMUS NIGER EXTRACT
C2940254|T121|1311151|RXNORM|PULEX IRRITANS PREPARATION|PULEX IRRITANS PREPARATION
C0035493|T196|1311402|RXNORM|RHODIUM|RHODIUM
C3464610|T121|1292748|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / PHYTOSTEROLS|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / PHYTOSTEROLS
C0301366|T121|89778|RXNORM|ECHOTHIOPHATE|ECHOTHIOPHATE
C3488253|T197|1311159|RXNORM|LEAD IODIDE PREPARATION|LEAD IODIDE PREPARATION
C3256396|T109|1424646|RXNORM|(PHTHALOCYANINATO(2-)) COPPER|(PHTHALOCYANINATO(2-)) COPPER
C3256399|T121|1424647|RXNORM|ALPHA-GLUCAN OLIGOSACCHARIDE|ALPHA-GLUCAN OLIGOSACCHARIDE
C3644331|T121|1424644|RXNORM|COCETH-7 CARBOXYLIC ACID|COCETH-7 CARBOXYLIC ACID
C3495485|T121|1424645|RXNORM|PURSLANE EXTRACT|PURSLANE EXTRACT
C0020306|T121|5509|RXNORM|HYDROQUINONE|HYDROQUINONE
C0020306|T121|5509|RXNORM|HYDROQUINONE|HYDROQUINONE
C2928868|T121|1007955|RXNORM|NAFTAZONE / RUTIN|NAFTAZONE / RUTIN
C3538397|T121|1372677|RXNORM|AMYLASES / ENDOPEPTIDASES / PAPAIN|AMYLASES / ENDOPEPTIDASES / PAPAIN
C2730104|T129|892332|RXNORM|PECAN ALLERGENIC EXTRACT|PECAN ALLERGENIC EXTRACT
C0217873|T121|1424648|RXNORM|TOCOTRIENOL, ALPHA|TOCOTRIENOL, ALPHA
C2928867|T121|1007954|RXNORM|ENSULIZOLE / ZINC OXIDE|ENSULIZOLE / ZINC OXIDE
C2343853|T121|797195|RXNORM|FESOTERODINE|FESOTERODINE
C2722774|T129|1098455|RXNORM|SUDAN GRASS POLLEN EXTRACT|SORGHUM BICOR SSP. DRUMMONDII POLLEN EXTRACT
C0076705|T121|38298|RXNORM|TIOCONAZOLE|TIOCONAZOLE
C0078595|T121|39801|RXNORM|XAMOTEROL|XAMOTEROL
C2054225|T121|813441|RXNORM|PHENOL / TANNIC ACID|PHENOL / TANNIC ACID
C0071166|T109|1426868|RXNORM|PIVALIC ACID|PIVALIC ACID
C2928872|T121|1007959|RXNORM|ETHAMIVAN / ETOFYLLINE / HEXOBENDINE|ETHAMIVAN / ETOFYLLINE / HEXOBENDINE
C2928689|T121|1007774|RXNORM|CALCIUM STEARATE / CHOLECALCIFEROL|CALCIUM STEARATE / CHOLECALCIFEROL
C3489261|T121|1309831|RXNORM|OCIMUM AMERICANUM LEAF EXTRACT|OCIMUM AMERICANUM LEAF EXTRACT
C3485650|T121|1304510|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / CUPRIC OXIDE / DOCUSATE / FOLIC ACID / IRON CARBONYL / MAGNESIUM OXIDE / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC OXIDE|ALPHA TOCOPHEROL / ASCORBIC ACID / CALCIUM CARBONATE / CHOLECALCIFEROL / CUPRIC OXIDE / DOCUSATE / FOLIC ACID / IRON CARBONYL / MAGNESIUM OXIDE / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC OXIDE
C3486629|T121|1309833|RXNORM|ARALIA RACEMOSA ROOT EXTRACT|ARALIA RACEMOSA ROOT EXTRACT
C3267744|T121|1309832|RXNORM|IRIS PALLIDA ROOT EXTRACT|IRIS PALLIDA ROOT EXTRACT
C0053170|T121|993243|RXNORM|BENZENESULFONIC ACID|BENZENESULFONIC ACID
C3541379|T126|1426865|RXNORM|LYSOZYME|LYSOZYME
C0079633|T129|1426866|RXNORM|INTERLEUKIN-8|INTERLEUKIN-8
C0028101|T196|1426867|RXNORM|NIOBIUM|NIOBIUM
C0301042|T121|89552|RXNORM|PHENOXYETHANOL|PHENOXYETHANOL
C3848595|T121|1545170|RXNORM|APIS CERANA WHOLE PREPARATION|APIS CERANA WHOLE PREPARATION
C0301404|T121|89808|RXNORM|CHLORAL BETAINE|CHLORAL BETAINE
C1646045|T121|607278|RXNORM|CALCIUM CARBONATE / RISEDRONATE|CALCIUM CARBONATE / RISEDRONATE
C0754923|T123|1440288|RXNORM|SINAPULTIDE|SINAPULTIDE
C3667902|T121|1440289|RXNORM|TRIPTERYGIUM WILFORDII WHOLE EXTRACT|TRIPTERYGIUM WILFORDII WHOLE EXTRACT
C1948466|T121|705701|RXNORM|PETIVERIA ALLIACEA PREPARATION|PETIVERIA ALLIACEA PREPARATION
C3190457|T121|1144760|RXNORM|BETAINE / FOLIC ACID / MECOBALAMIN / PYRIDOXINE|BETAINE / FOLIC ACID / MECOBALAMIN / PYRIDOXINE
C3667900|T131|1440286|RXNORM|OXYURANUS SCUTELLATUS CANNI VENOM EXTRACT|OXYURANUS SCUTELLATUS CANNI VENOM EXTRACT
C3667901|T131|1440287|RXNORM|CROTALUS DURISSUS TERRIFICUS VENOM EXTRACT|CROTALUS DURISSUS TERRIFICUS VENOM EXTRACT
C0528926|T121|136034|RXNORM|FERROUS LACTATE|FERROUS LACTATE
C2928488|T121|1007568|RXNORM|CODEINE / GUAIACOLSULFONIC ACID / PHENYLEPHRINE / PROMETHAZINE|CODEINE / GUAIACOLSULFONIC ACID / PHENYLEPHRINE / PROMETHAZINE
C2928489|T121|1007569|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / CODEINE|ACETAMINOPHEN / CHLORPHENIRAMINE / CODEINE
C1655131|T121|1007560|RXNORM|ALENDRONATE / CHOLECALCIFEROL|ALENDRONATE / CHOLECALCIFEROL
C2928481|T121|1007561|RXNORM|ATROPINE / HYDROMORPHONE|ATROPINE / HYDROMORPHONE
C2928482|T121|1007562|RXNORM|ECHINACEA PURPUREA EXTRACT / PECTIN|ECHINACEA PURPUREA EXTRACT / PECTIN
C2928483|T121|1007563|RXNORM|CALCIUM LACTATE / GLUCOSE / MAGNESIUM CITRATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE|CALCIUM LACTATE / GLUCOSE / MAGNESIUM CITRATE / POTASSIUM CHLORIDE / SODIUM CHLORIDE
C3664991|T121|1435097|RXNORM|PHYSALIS ALKEKENGI FRUIT EXTRACT|PHYSALIS ALKEKENGI FRUIT EXTRACT
C2928486|T121|1007566|RXNORM|BENZENESULFONIC ACID / HYDROGEN PEROXIDE / LACTATE|BENZENESULFONIC ACID / HYDROGEN PEROXIDE / LACTATE
C2928487|T121|1007567|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-CALIFORNIA-7-2009 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-PERTH-16-2009 (H3N2) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-BRISBANE-60-2008 STRAIN|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-CALIFORNIA-7-2009 (H1N1) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-PERTH-16-2009 (H3N2) STRAIN / INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-BRISBANE-60-2008 STRAIN
C1874246|T121|691169|RXNORM|ANTAZOLINE / NAPHAZOLINE|ANTAZOLINE / NAPHAZOLINE
C3664990|T121|1435096|RXNORM|MELALEUCA ALTERNIFOLIA FLOWERING TOP EXTRACT|MELALEUCA ALTERNIFOLIA FLOWERING TOP EXTRACT
C1875867|T121|691161|RXNORM|YOHIMBINE / ZINC SULFATE|YOHIMBINE / ZINC SULFATE
C0061516|T121|25953|RXNORM|GLUTATHIONE DISULFIDE|GLUTATHIONE DISULFIDE
C2183385|T121|821410|RXNORM|DIAZEPAM / DIETHYLPROPION / FENPROPOREX|DIAZEPAM / DIETHYLPROPION / FENPROPOREX
C0249582|T127|73710|RXNORM|PARICALCITOL|PARICALCITOL
C0014025|T121|3827|RXNORM|ENALAPRIL|ENALAPRIL
C0078643|T121|39841|RXNORM|XYLOMETAZOLINE|XYLOMETAZOLINE
C2194286|T121|812737|RXNORM|ALBUTEROL / GUAIFENESIN|ALBUTEROL / GUAIFENESIN
C0013974|T121|3820|RXNORM|EMETINE|EMETINE
C3848594|T109|1545358|RXNORM|PEG-20 GLYCERYL TRIISOSTEARATE|PEG-20 GLYCERYL TRIISOSTEARATE
C0770963|T129|1099933|RXNORM|ADENOVIRUS TYPE 4 VACCINE LIVE|ADENOVIRUS TYPE 4 VACCINE LIVE
C0014027|T121|3829|RXNORM|ENALAPRILAT|ENALAPRILAT
C0770964|T129|1099937|RXNORM|ADENOVIRUS TYPE 7 VACCINE LIVE|ADENOVIRUS TYPE 7 VACCINE LIVE
C0012024|T195|3328|RXNORM|DIBEKACIN|DIBEKACIN
C2241636|T121|761177|RXNORM|BROMPHENIRAMINE / DIHYDROCODEINE / PHENYLEPHRINE|BROMPHENIRAMINE / DIHYDROCODEINE / PHENYLEPHRINE
C0072159|T121|34633|RXNORM|PROPAMIDINE|PROPAMIDINE
C0873113|T121|259449|RXNORM|GRAPEFRUIT SEED EXTRACT|CITRUS PARADISI SEED EXTRACT
C2929821|T121|1008924|RXNORM|ASCORBIC ACID / CALCIUM SULFATE / CHOLECALCIFEROL / CUPRIC OXIDE / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / CALCIUM SULFATE / CHOLECALCIFEROL / CUPRIC OXIDE / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC OXIDE
C1875250|T121|689704|RXNORM|HEXACHLOROPHENE / HYDROCORTISONE / MENTHOL|HEXACHLOROPHENE / HYDROCORTISONE / MENTHOL
C0937873|T121|283767|RXNORM|MANGANESE CITRATE|MANGANESE CITRATE
C2722023|T129|971932|RXNORM|OAT ALLERGENIC EXTRACT|OAT ALLERGENIC EXTRACT
C3664992|T121|1435099|RXNORM|CITRUS MEDICA FRUIT EXTRACT|CITRUS MEDICA FRUIT EXTRACT
C0960501|T130|1366938|RXNORM|IMINODISUCCINATE|IMINODISUCCINATE
C1875253|T121|689708|RXNORM|HOMATROPINE / OPIUM / PECTIN|HOMATROPINE / OPIUM / PECTIN
C3542462|T121|1435098|RXNORM|SOURSOP EXTRACT|ANNONA MURICATA FRUIT EXTRACT
C0028458|T195|7538|RXNORM|NOVOBIOCIN|NOVOBIOCIN
C0028420|T121|7531|RXNORM|NORTRIPTYLINE|NORTRIPTYLINE
C1337242|T121|407990|RXNORM|CINACALCET|CINACALCET
C0028426|T121|7533|RXNORM|NOSCAPINE|NOSCAPINE
C3256267|T121|1307697|RXNORM|RUBES NIGRUM SEED EXTRACT|RUBES NIGRUM SEED EXTRACT
C3256630|T121|1307696|RXNORM|POLYGONATUM MULTIFLORUM ROOT EXTRACT|POLYGONATUM MULTIFLORUM ROOT EXTRACT
C0060124|T130|1307695|RXNORM|FD&C BLUE #2 LAKE|FD&C BLUE #2 LAKE
C3257191|T130|1307694|RXNORM|FD&C BLUE #1 ALUMINUM LAKE|FD&C BLUE #1 ALUMINUM LAKE
C2347980|T109|1307693|RXNORM|ROSEWOOD OIL|ROSEWOOD OIL
C3256792|T121|1307692|RXNORM|ONONIS CAMPESTRIS ROOT EXTRACT|ONONIS SPINOSA ROOT EXTRACT
C0069805|T121|32675|RXNORM|OXYBUTYNIN|OXYBUTYNIN
C3256290|T121|1307690|RXNORM|AMARANTHUS CAUDATUS SEED EXTRACT|AMARANTHUS CAUDATUS SEED EXTRACT
C0053941|T121|19605|RXNORM|BOPINDOLOL|BOPINDOLOL
C3255948|T121|1307853|RXNORM|MAGNOLIA OFFICINALIS BARK EXTRACT|MAGNOLIA OFFICINALIS BARK EXTRACT
C3256853|T121|1307699|RXNORM|LAWSONIA INERMIS LEAF EXTRACT|LAWSONIA INERMIS LEAF EXTRACT
C3484418|T121|1307698|RXNORM|SAMBUCUS NIGRA FLOWERING TOP|SAMBUCUS NIGRA FLOWERING TOP
C3264697|T121|1307852|RXNORM|MENTHA AQUATICA LEAF EXTRACT|MENTHA AQUATICA LEAF EXTRACT
C0663384|T121|190433|RXNORM|PRAMIVERINE|PRAMIVERINE
C3485014|T121|1307855|RXNORM|PIPER KADSURA STEM EXTRACT|PIPER KADSURA STEM EXTRACT
C1874157|T121|690989|RXNORM|ALUMINUM ACETATE / CAMPHOR / MENTHOL / PHENOL|ALUMINUM ACETATE / CAMPHOR / MENTHOL / PHENOL
C2344315|T129|798292|RXNORM|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G4 VACCINE|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G4 VACCINE
C3257445|T121|1307857|RXNORM|RHUS GLABRA BARK EXTRACT|RHUS GLABRA BARK EXTRACT
C2726437|T121|884629|RXNORM|CALCIUM PYRUVATE|CALCIUM PYRUVATE
C3255686|T121|1307856|RXNORM|HOLARRHENA PUBESCENS BARK EXTRACT|HOLARRHENA PUBESCENS BARK EXTRACT
C0059865|T121|24605|RXNORM|ETODOLAC|ETODOLAC
C0359949|T121|107602|RXNORM|EPINEPHRINE / LIDOCAINE|EPINEPHRINE / LIDOCAINE
C3651734|T121|1429939|RXNORM|MELIA AZEDARACH WHOLE EXTRACT|MELIA AZEDARACH WHOLE EXTRACT
C3651737|T121|1429933|RXNORM|ISOPROPYL ISOBUTYRATE|ISOPROPYL ISOBUTYRATE
C0109497|T123|1426483|RXNORM|CHOLATE|CHOLATE
C0303763|T130|1426480|RXNORM|LIQUEFIED PETROLEUM GAS|LIQUEFIED PETROLEUM GAS
C2962064|T129|1426481|RXNORM|CLONOSTACHYS ROSEA F. ROSEA ALLERGENIC EXTRACT|CLONOSTACHYS ROSEA F. ROSEA ALLERGENIC EXTRACT
C3651735|T109|1429937|RXNORM|MACADAMIA SEED OIL GLYCERETH-8 ESTERS|MACADAMIA SEED OIL GLYCERETH-8 ESTERS
C0059868|T121|24608|RXNORM|ETOFENAMATE|ETOFENAMATE
C3651736|T121|1429934|RXNORM|LIMNANTHES ALBA WHOLE EXTRACT|LIMNANTHES ALBA WHOLE EXTRACT
C0065501|T121|1551573|RXNORM|MADECASSIC ACID|MADECASSIC ACID
C3857956|T109|1551572|RXNORM|METHYL LACTATE, (+)-|METHYL LACTATE, (+)-
C3857957|T121|1551571|RXNORM|ACV TRIPEPTIDE|ACV TRIPEPTIDE
C3531639|T109|1367425|RXNORM|RUTA GRAVEOLENS FLOWERING TOP OIL|RUTA GRAVEOLENS FLOWERING TOP OIL
C0081660|T121|1551574|RXNORM|ASIATIC ACID|ASIATIC ACID
C2827183|T121|1376345|RXNORM|HYPROMELLOSE ACETATE SUCCINATE 06081224 (3 MM2-S)|HYPROMELLOSE ACETATE SUCCINATE 06081224 (3 MM2-S)
C0055747|T121|21125|RXNORM|CINITAPRIDE|CINITAPRIDE
C2193911|T121|813460|RXNORM|BUFLOMEDIL / DIOSMIN|BUFLOMEDIL / DIOSMIN
C0717545|T121|214349|RXNORM|CALCIUM CARBONATE / SODIUM FLUORIDE|CALCIUM CARBONATE / SODIUM FLUORIDE
C0717537|T130|214342|RXNORM|CALCIUM ACETATE|CALCIUM ACETATE
C1174840|T121|356834|RXNORM|DERACOXIB|DERACOXIB
C0717542|T121|214346|RXNORM|CALCIUM CARBONATE / MAGNESIUM CARBONATE|CALCIUM CARBONATE / MAGNESIUM CARBONATE
C0717543|T121|214347|RXNORM|CALCIUM CARBONATE / MAGNESIUM HYDROXIDE|CALCIUM CARBONATE / MAGNESIUM HYDROXIDE
C3249317|T121|1235143|RXNORM|AZILSARTAN / CHLORTHALIDONE|AZILSARTAN / CHLORTHALIDONE
C0068771|T121|31805|RXNORM|NILUTAMIDE|NILUTAMIDE
C0949222|T121|287637|RXNORM|CALCIUM ASPARTATE|CALCIUM ASPARTATE
C3818732|T121|1534766|RXNORM|ANDROGRAPHIS PANICULATA WHOLE EXTRACT|ANDROGRAPHIS PANICULATA WHOLE EXTRACT
C0053332|T121|19084|RXNORM|BENZYLTHIOURACIL|BENZYLTHIOURACIL
C0597484|T196|1364429|RXNORM|SODIUM CATION|SODIUM CATION
C0035923|T129|9486|RXNORM|RUBELLA VIRUS VACCINE|RUBELLA, LIVE ATTENUATED
C0064711|T197|1423667|RXNORM|LEAD ACETATE|LEAD ACETATE
C0011522|T126|3210|RXNORM|DEOXYRIBONUCLEASES|DEOXYRIBONUCLEASES
C1263450|T121|386055|RXNORM|LAUROMACROGOLS|LAUROMACROGOLS
C0056057|T121|21389|RXNORM|COCOA BUTTER|COCOA BUTTER
C0772002|T197|1305582|RXNORM|FERRIC OXIDE YELLOW|FERRIC OXIDE YELLOW
C3695984|T109|1482794|RXNORM|CURCUMA AROMATICA ROOT OIL|CURCUMA AROMATICA ROOT OIL
C2605855|T121|1482790|RXNORM|SIMEPREVIR|SIMEPREVIR
C3695986|T121|1482791|RXNORM|DACTYLOPIUS COCCUS WHOLE EXTRACT|DACTYLOPIUS COCCUS WHOLE EXTRACT
C1612168|T109|1482792|RXNORM|PENOXSULAM|PENOXSULAM
C3695985|T121|1482793|RXNORM|TYLOPHORA INDICA LEAF EXTRACT|TYLOPHORA INDICA LEAF EXTRACT
C0043465|T121|1368476|RXNORM|ZERANOL|ZERANOL
C3535676|T109|1368471|RXNORM|DIMETHICONE-VINYL DIMETHICONE CROSSPOLYMER (HARD PARTICLE)|DIMETHICONE-VINYL DIMETHICONE CROSSPOLYMER (HARD PARTICLE)
C2929058|T121|1008151|RXNORM|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / INTRINSIC FACTOR / VITAMIN B 12|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / INTRINSIC FACTOR / VITAMIN B 12
C0017687|T125|4832|RXNORM|GLUCAGON|GLUCAGON
C0030859|T125|7993|RXNORM|PENTAGASTRIN|PENTAGASTRIN
C0770739|T121|235618|RXNORM|MOLD EXTRACT|MOLD EXTRACT
C0178649|T123|618771|RXNORM|GAMMA-AMINOBUTYRATE|GAMMA-AMINOBUTYRATE
C0030863|T121|7994|RXNORM|PENTAMIDINE|PENTAMIDINE
C0030863|T121|7994|RXNORM|PENTAMIDINE|PENTAMIDINE
C3556195|T121|1375959|RXNORM|CHOLECALCIFEROL / GLUCOSE|CHOLECALCIFEROL / GLUCOSE
C0043822|T121|11636|RXNORM|DROSPIRENONE|DROSPIRENONE
C0008188|T121|2356|RXNORM|POLLEN EXTRACTS|CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|STOCK RAGWEED POLLEN MIXTURE|CHLORDIAZEPOXIDE
C0178793|T127|62400|RXNORM|PANTOTHENATE|PANTOTHENATE
C3709747|T109|1488263|RXNORM|VERNICIA FORDII SEED OIL|VERNICIA FORDII SEED OIL
C0019453|T131|5296|RXNORM|ALTRETAMINE|ALTRETAMINE
C0772151|T121|236832|RXNORM|SULFACHRYSOIDINE|SULFACHRYSOIDINE
C2722032|T130|892653|RXNORM|CHICKEN ALLERGENIC EXTRACT|GALLUS GALLUS ALLERGENIC EXTRACT
C0019435|T121|5293|RXNORM|HEXACHLOROPHENE|HEXACHLOROPHENE
C2073895|T121|813110|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PYRILAMINE|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PYRILAMINE
C3709749|T121|1488269|RXNORM|MOXIDECTIN / PRAZIQUANTEL|MOXIDECTIN / PRAZIQUANTEL
C0440459|T131|124427|RXNORM|HONEY BEE VENOM|HONEY BEE VENOM
C3488381|T121|1311411|RXNORM|ANEMONE AMERICANA EXTRACT|ANEMONE AMERICANA EXTRACT
C0282085|T121|81971|RXNORM|CANRENOIC ACID|CANRENOIC ACID
C0069451|T197|1368210|RXNORM|OLIVINE|OLIVINE
C0077030|T121|1314420|RXNORM|TRICAPRYLIN|GLYCEROL TRICAPRYLATE
C0067790|T121|1368212|RXNORM|N-ACETYLTRYPTOPHAN|N-ACETYLTRYPTOPHAN
C0761662|T109|1368213|RXNORM|1-BUTYL OLEATE|1-BUTYL OLEATE
C0982416|T121|1368215|RXNORM|STEARAMIDE AMP|STEARAMIDE AMP
C0028403|T123|1311141|RXNORM|OCTOPAMINE|OCTOPAMINE
C2356074|T121|802683|RXNORM|CHLOPHEDIANOL / GUAIFENESIN / PSEUDOEPHEDRINE|CHLOPHEDIANOL / GUAIFENESIN / PSEUDOEPHEDRINE
C3152925|T121|1310055|RXNORM|MORUS ALBA ROOT BARK EXTRACT|MORUS ALBA ROOT BARK EXTRACT
C3486735|T121|1310057|RXNORM|TEUCRIUM SCORODONIA FLOWERING TOP EXTRACT|TEUCRIUM SCORODONIA FLOWERING TOP EXTRACT
C3484564|T121|1310056|RXNORM|JACARANDA CAROBA FLOWER EXTRACT|JACARANDA CAROBA FLOWER EXTRACT
C3486731|T121|1310051|RXNORM|SOLANUM DULCAMARA FLOWER EXTRACT|SOLANUM DULCAMARA FLOWER EXTRACT
C2981080|T121|1310050|RXNORM|STILLINGIA SYLVATICA ROOT EXTRACT|STILLINGIA SYLVATICA ROOT EXTRACT
C3486734|T121|1310052|RXNORM|NYMPHAEA ODORATA ROOT EXTRACT|NYMPHAEA ODORATA ROOT EXTRACT
C0032949|T121|8637|RXNORM|PREDNIMUSTINE|PREDNIMUSTINE
C0537270|T125|139825|RXNORM|INSULIN DETEMIR|INSULIN DETEMIR
C0071883|T121|34407|RXNORM|PRENYLAMINE LACTATE|PRENYLAMINE LACTATE
C2146629|T121|820354|RXNORM|ACETAMINOPHEN / PYRILAMINE|ACETAMINOPHEN / PYRILAMINE
C1506770|T121|480167|RXNORM|LAPATINIB|LAPATINIB
C0031432|T121|8143|RXNORM|PHENOPERIDINE|PHENOPERIDINE
C2701074|T129|851740|RXNORM|BOX ELDER MAPLE POLLEN EXTRACT|ACER NEGUNDO POLLEN EXTRACT
C3651777|T109|1428833|RXNORM|BENZOPHENONE-5|BENZOPHENONE-5
C1095890|T121|1309324|RXNORM|WORMWOOD EXTRACT|WORMWOOD EXTRACT
C0027780|T195|7337|RXNORM|NETILMICIN|NETILMICIN
C0288672|T129|83929|RXNORM|ABCIXIMAB|ABCIXIMAB
C0672596|T129|194279|RXNORM|PALIVIZUMAB|PALIVIZUMAB
C0069834|T121|32699|RXNORM|OXYPOLYGELATINE|OXYPOLYGELATINE
C3864852|T121|1595034|RXNORM|DODECENE|1-DODECENE
C3555471|T121|1420971|RXNORM|LINDERA AGGREGATA ROOT EXTRACT|LINDERA AGGREGATA ROOT EXTRACT
C0885180|T121|265758|RXNORM|CANTHARIS VESICATORIA PREPARATION|CANTHARIS VESICATORIA PREPARATION
C0036193|T121|9556|RXNORM|SARALASIN|SARALASIN
C2928864|T121|1007951|RXNORM|BENZOCAINE / DEQUALINIUM / TYROTHRICIN|BENZOCAINE / DEQUALINIUM / TYROTHRICIN
C2928863|T121|1007950|RXNORM|TETRACAINE / TYROTHRICIN|TETRACAINE / TYROTHRICIN
C2928866|T121|1007953|RXNORM|CALCIUM GLUCONATE / CALCIUM LACTATE|CALCIUM GLUCONATE / CALCIUM LACTATE
C2928865|T121|1007952|RXNORM|CHLORTHALIDONE / HYDRALAZINE / OXPRENOLOL|CHLORTHALIDONE / HYDRALAZINE / OXPRENOLOL
C2928694|T121|1007779|RXNORM|EPHEDRINE / SODIUM IODIDE|EPHEDRINE / SODIUM IODIDE
C2928693|T121|1007778|RXNORM|BIOTIN / CALCIUM CARBONATE|BIOTIN / CALCIUM CARBONATE
C2928870|T121|1007957|RXNORM|OXELADIN / REPROTEROL|OXELADIN / REPROTEROL
C2928869|T121|1007956|RXNORM|DEQUALINIUM / TYROTHRICIN|DEQUALINIUM / TYROTHRICIN
C2928690|T121|1007775|RXNORM|CALCIUM CARBONATE / MAGNESIUM OXIDE / ZINC GLUCONATE|CALCIUM CARBONATE / MAGNESIUM OXIDE / ZINC GLUCONATE
C2928871|T121|1007958|RXNORM|ASCORBIC ACID / POTASSIUM CITRATE|ASCORBIC ACID / POTASSIUM CITRATE
C2928692|T121|1007777|RXNORM|CARBETAPENTANE / GUAIACOLSULFONATE / PHENYLEPHRINE / PHENYLPROPANOLAMINE|CARBETAPENTANE / GUAIACOLSULFONATE / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C2928691|T121|1007776|RXNORM|DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM CHLORIDE / SODIUM PHOSPHATE, MONOBASIC|DIBASIC POTASSIUM PHOSPHATE / GLUCOSE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM CHLORIDE / SODIUM PHOSPHATE, MONOBASIC
C2928686|T121|1007771|RXNORM|ASCORBIC ACID / CHONDROITIN SULFATES / GLUCOSAMINE|ASCORBIC ACID / CHONDROITIN SULFATES / GLUCOSAMINE
C2928685|T121|1007770|RXNORM|NIACIN / PENTAERYTHRITOL|NIACIN / PENTAERYTHRITOL
C2928687|T121|1007772|RXNORM|ASCORBIC ACID / BIOTIN / FOLIC ACID / MECOBALAMIN / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE|ASCORBIC ACID / BIOTIN / FOLIC ACID / MECOBALAMIN / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE
C3257504|T121|1426863|RXNORM|COCONUT ALCOHOL|COCONUT ALCOHOL
C3538018|T121|1371880|RXNORM|MONOFLUOROPHOSPHATE / POTASSIUM NITRATE / ZINC CITRATE|MONOFLUOROPHOSPHATE / POTASSIUM NITRATE / ZINC CITRATE
C0666743|T129|191831|RXNORM|INFLIXIMAB|INFLIXIMAB
C3531112|T121|1366113|RXNORM|HURA CREPITANS SAP EXTRACT|HURA CREPITANS SAP EXTRACT
C0038753|T130|10212|RXNORM|SULFOBROMOPHTHALEIN|SULFOBROMOPHTHALEIN
C3834063|T109|1542375|RXNORM|PENTAERYTHRITYL TETRABEHENATE|PENTAERYTHRITYL TETRABEHENATE
C2938407|T129|1012183|RXNORM|RED KIDNEY BEAN ALLERGENIC EXTRACT|RED KIDNEY BEAN ALLERGENIC EXTRACT
C3541308|T121|1376349|RXNORM|THYMUS VULGARIS WHOLE EXTRACT|THYMUS VULGARIS WHOLE EXTRACT
C3555487|T109|1376348|RXNORM|ROSMARINUS OFFICINALIS FLOWERING TOP OIL|ROSMARINUS OFFICINALIS FLOWERING TOP OIL
C0359955|T121|107608|RXNORM|FELYPRESSIN / PRILOCAINE|FELYPRESSIN / PRILOCAINE
C0359957|T121|107609|RXNORM|COCAINE / EPINEPHRINE|COCAINE / EPINEPHRINE
C3643652|T121|1424269|RXNORM|STEAROAMPHOACETATE|STEAROAMPHOACETATE
C0026549|T121|7052|RXNORM|MORPHINE|MORPHINE
C0359950|T121|107603|RXNORM|CHLORHEXIDINE / LIDOCAINE|CHLORHEXIDINE / LIDOCAINE
C0603000|T122|1376343|RXNORM|CYCLAMEN ALDEHYDE|CYCLAMEN ALDEHYDE
C0052168|T121|1376342|RXNORM|APOCAROTENAL|APOCAROTENAL
C0359953|T121|107606|RXNORM|BUPIVACAINE / EPINEPHRINE|BUPIVACAINE / EPINEPHRINE
C3555488|T121|1376344|RXNORM|HYDROXYETHYL CELLULOSE (6500 MPA.S AT 2%)|HYDROXYETHYL CELLULOSE (6500 MPA.S AT 2%)
C3539016|T121|1376347|RXNORM|OLEA EUROPAEA WHOLE EXTRACT|OLEA EUROPAEA WHOLE EXTRACT
C3542425|T121|1376346|RXNORM|LAVANDULA ANGUSTIFOLIA WHOLE EXTRACT|LAVANDULA ANGUSTIFOLIA WHOLE EXTRACT
C3256446|T130|1305585|RXNORM|SYNTHETIC YELLOW IRON OXIDE|SYNTHETIC YELLOW IRON OXIDE
C0112458|T120|1305581|RXNORM|D&C YELLOW NO. 11|D&C YELLOW NO. 11
C0078034|T121|39371|RXNORM|VANILLYL-N-NONYLAMIDE|VANILLYL-N-NONYLAMIDE
C3473202|T121|1298309|RXNORM|ASCORBIC ACID / BIOTIN / FOLIC ACID / NIACIN / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN E|ASCORBIC ACID / BIOTIN / FOLIC ACID / NIACIN / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / VITAMIN E
C3489115|T121|1311232|RXNORM|SUS SCROFA ORAL MUCOSA PREPARATION|PORCINE ORAL MUCOSA PREPARATION
C2728183|T129|1010965|RXNORM|OREGANO ALLERGENIC EXTRACT|OREGANO ALLERGENIC EXTRACT
C3486799|T121|1311234|RXNORM|SUS SCROFA GALLBLADDER PREPARATION|PORCINE GALLBLADDER PREPARATION
C3487983|T121|1311235|RXNORM|SUS SCROFA ADRENAL GLAND PREPARATION|PORCINE ADRENAL GLAND PREPARATION
C0031441|T121|8149|RXNORM|PHENOXYBENZAMINE|PHENOXYBENZAMINE
C2740640|T130|899448|RXNORM|LETTUCE ALLERGENIC EXTRACT|LATUCA SATIVA ALLERGENIC EXTRACT
C0939820|T121|1297537|RXNORM|YELLOW HORNET VENOM PROTEIN|DOLICHOVESPULA ARENARIA VENOM PROTEIN
C0032950|T121|8638|RXNORM|PREDNISOLONE|PREDNISOLONE
C0032950|T121|8638|RXNORM|PREDNISOLONE|PREDNISOLONE
C0031430|T130|8141|RXNORM|PHENOLSULFONPHTHALEIN|PHENOLSULFONPHTHALEIN
C0026234|T195|6995|RXNORM|PLICAMYCIN|PLICAMYCIN
C0026236|T121|6996|RXNORM|MITOBRONITOL|MITOBRONITOL
C0006706|T109|1485048|RXNORM|CALCIUM OXALATE|CALCIUM OXALATE
C3489227|T121|1309825|RXNORM|TYLOPHORA INDICA ROOT EXTRACT|TYLOPHORA INDICA ROOT EXTRACT
C3818782|T109|1491868|RXNORM|PIGMENT YELLOW 3|PIGMENT YELLOW 3
C3818781|T109|1491869|RXNORM|3,4,9,10-PERYLENETETRACARBOXYLIC DIIMIDE|3,4,9,10-PERYLENETETRACARBOXYLIC DIIMIDE
C0318143|T007|1491866|RXNORM|STREPTOCOCCUS DYSGALACTIAE|STREPTOCOCCUS DYSGALACTIAE
C3282145|T121|1426948|RXNORM|TRIMETHYLSILOXYSILICATE (M-Q 0.66)|TRIMETHYLSILOXYSILICATE (M-Q 0.66)
C0318150|T007|1491864|RXNORM|STREPTOCOCCUS UBERIS|STREPTOCOCCUS UBERIS
C3163630|T007|1491865|RXNORM|STREPTOCOCCUS EQUINUS|STREPTOCOCCUS EQUINUS
C0376325|T005|1491862|RXNORM|HEPATITIS A VIRUS|HEPATITIS A VIRUS
C0220847|T005|1491863|RXNORM|HEPATITIS C VIRUS|HEPATITIS C VIRUS
C3818784|T109|1491860|RXNORM|RIBES NIGRUM LEAF EXTRACT|RIBES NIGRUM LEAF EXTRACT
C3488691|T121|1309823|RXNORM|TILIA X EUROPAEA FLOWER EXTRACT|TILIA X EUROPAEA FLOWER EXTRACT
C3486070|T121|1311096|RXNORM|VISCUM ALBUM FRUITING TOP EXTRACT|VISCUM ALBUM FRUITING TOP EXTRACT
C1602364|T121|541439|RXNORM|SODIUM GLYCINATE|SODIUM GLYCINATE
C0021344|T005|1311095|RXNORM|HUMAN PAPILLOMAVIRUS|HUMAN PAPILLOMAVIRUS
C3486641|T121|1311092|RXNORM|MOMORDICA BALSAMINA IMMATURE FRUIT EXTRACT|MOMORDICA BALSAMINA IMMATURE FRUIT EXTRACT
C2346927|T196|1426853|RXNORM|MAGNESIUM CATION|MN 2+
C3486658|T197|1311090|RXNORM|BARIUM OXALOSUCCINATE|BARIUM OXALOSUCCINATE
C3489125|T121|1311091|RXNORM|THERIDION CURASSAVICUM PREPARATION|THERIDION CURASSAVICUM PREPARATION
C0724699|T121|221166|RXNORM|STANDARDIZED SENNA CONCENTRATE|STANDARDIZED SENNA CONCENTRATE
C2740659|T129|899476|RXNORM|HONEYDEW MELON ALLERGENIC EXTRACT|HONEYDEW MELON ALLERGENIC EXTRACT
C0075630|T121|37416|RXNORM|SULTOPRIDE|SULTOPRIDE
C0025423|T197|1311098|RXNORM|CALOMEL|CALOMEL
C2983917|T130|1486026|RXNORM|FLUTEMETAMOL|FLUTEMETAMOL
C0209738|T121|68244|RXNORM|LAMIVUDINE|LAMIVUDINE
C3818729|T121|1534776|RXNORM|THREE-LOBE SAGE EXTRACT|THREE-LOBE SAGE EXTRACT
C3818728|T121|1534777|RXNORM|DICENTRA CANADENSIS ROOT EXTRACT|DICENTRA CANADENSIS ROOT EXTRACT
C0043432|T196|1534770|RXNORM|YTTRIUM|YTTRIUM
C3474134|T121|1313687|RXNORM|ELEUTHEROCOCCUS SESSILFLORUS WHOLE EXTRACT|ELEUTHEROCOCCUS SESSILFLORUS WHOLE EXTRACT
C0024170|T197|1534772|RXNORM|LUTETIUM|LUTETIUM
C3642427|T121|1543173|RXNORM|TAVABOROLE|TAVABOROLE
C3163077|T121|1115703|RXNORM|DYCLONINE / GLYCERIN|DYCLONINE / GLYCERIN
C3818727|T122|1534778|RXNORM|LIMONEN-10-OL, (+)-|LIMONEN-10-OL, (+)-
C0025810|T121|6901|RXNORM|PSYLLIUM / SUCROSE|METHYLPHENIDATE
C0220802|T109|596718|RXNORM|BUTYRATE|BUTYRATE
C0014968|T121|4112|RXNORM|ETHAMSYLATE|ETHAMSYLATE
C3645199|T121|1426858|RXNORM|GLYOXAL TRIMER|GLYOXAL TRIMER
C0724561|T197|221083|RXNORM|SULFUR,COLLOIDAL|SULFUR,COLLOIDAL
C0724560|T121|221082|RXNORM|COLLOIDAL OATMEAL|COLLOIDAL OATMEAL
C0724560|T121|221082|RXNORM|COLLOIDAL OATMEAL|COLLOIDAL OATMEAL
C3486626|T121|1309828|RXNORM|ANGELICA ARCHANGELICA ROOT EXTRACT|ANGELICA ARCHANGELICA ROOT EXTRACT
C3265310|T121|1354504|RXNORM|SAGE EXTRACT|SAGE EXTRACT
C0037962|T195|9991|RXNORM|SPIRAMYCIN|SPIRAMYCIN
C3833310|T121|1541116|RXNORM|CAPRYLYL CAPRYLATE-CAPRATE|CAPRYLYL CAPRYLATE-CAPRATE
C3489255|T121|1309829|RXNORM|VERBENA OFFICINALIS FLOWERING TOP EXTRACT|VERBENA OFFICINALIS FLOWERING TOP EXTRACT
C1166065|T121|350374|RXNORM|BETAINE, ANHYDROUS|BETAINE, ANHYDROUS
C0037982|T121|9997|RXNORM|SPIRONOLACTONE|SPIRONOLACTONE
C3700882|T129|1486798|RXNORM|ANDROCTONUS AUSTRALIS VENOM|ANDROCTONUS AUSTRALIS VENOM
C3700881|T197|1486799|RXNORM|GOLD MONOIODIDE|GOLD MONOIODIDE
C3527959|T121|1361461|RXNORM|ATROPA BELLADONA WHOLE EXTRACT|ATROPA BELLADONA WHOLE EXTRACT
C2929135|T121|1008228|RXNORM|MAGNESIUM SULFATE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM CHLORIDE / SODIUM PHOSPHATE DIHYDRATE|MAGNESIUM SULFATE / POTASSIUM CHLORIDE / POTASSIUM PHOSPHATE / SODIUM CHLORIDE / SODIUM PHOSPHATE
C2929136|T121|1008229|RXNORM|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929136|T121|1008229|RXNORM|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2929134|T121|1008227|RXNORM|COENZYME Q10 / LEVOCARNITINE / VITAMIN E|COENZYME Q10 / LEVOCARNITINE / VITAMIN E
C2929131|T121|1008224|RXNORM|DIBASIC POTASSIUM PHOSPHATE / POTASSIUM PHOSPHATE|DIBASIC POTASSIUM PHOSPHATE / POTASSIUM PHOSPHATE
C2929132|T121|1008225|RXNORM|ALOE VERA PREPARATION / UREA|ALOE VERA PREPARATION / UREA
C2929129|T121|1008222|RXNORM|TROXERUTIN / VINCAMINE|TROXERUTIN / VINCAMINE
C2929130|T121|1008223|RXNORM|ALGINIC ACID / SODIUM BICARBONATE|ALGINIC ACID / SODIUM BICARBONATE
C2929127|T121|1008220|RXNORM|DIETHYLAMINE SALICYLATE / GLYCOL SALICYLATE / METHYLNICOTINATE|DIETHYLAMINE SALICYLATE / GLYCOL SALICYLATE / METHYLNICOTINATE
C2929128|T121|1008221|RXNORM|AMMONIUM FERROUS SULFATE / FOLIC ACID|AMMONIUM FERROUS SULFATE / FOLIC ACID
C2756545|T129|968498|RXNORM|TEA LEAF EXTRACT|TEA LEAF EXTRACT
C0064990|T197|28728|RXNORM|CALCIUM OXIDE|CALCIUM OXIDE
C0005059|T121|1399|RXNORM|BENZOCAINE|BENZOCAINE
C0005059|T121|1399|RXNORM|BENZOCAINE|BENZOCAINE
C0005059|T121|1399|RXNORM|BENZOCAINE|BENZOCAINE
C0005059|T121|1399|RXNORM|BENZOCAINE|BENZOCAINE
C0021988|T121|596712|RXNORM|IODOPHORS|IODOPHORS
C0001888|T121|423|RXNORM|AJMALINE|AJMALINE
C2193887|T121|818996|RXNORM|ESTRADIOL / ESTRONE|ESTRADIOL / ESTRONE
C0005041|T121|1390|RXNORM|BENZETHONIUM|BENZETHONIUM
C0005041|T121|1390|RXNORM|BENZETHONIUM|BENZETHONIUM
C3486395|T121|1331702|RXNORM|SOLANUM DULCAMARA TOP EXTRACT|SOLANUM DULCAMARA TOP EXTRACT
C0054255|T121|19880|RXNORM|BUTIBUFEN|BUTIBUFEN
C3486552|T121|1331704|RXNORM|CONYZA CANADENSIS EXTRACT|ERIGERON CANADENSIS EXTRACT
C3486766|T121|1331706|RXNORM|OLEA EUROPAEA FLOWER EXTRACT|OLEA EUROPAEA FLOWER EXTRACT
C0887700|T121|267453|RXNORM|SODIUM ACETATE, ANHYDROUS|SODIUM ACETATE, ANHYDROUS
C2701264|T129|852054|RXNORM|AMERICAN ELM POLLEN EXTRACT|ULMUS AMERICANA POLLEN EXTRACT
C2701609|T129|852503|RXNORM|FUSARIUM EXTRACT|HAEMATONECTRIA HAEMATOCOCCA EXTRACT
C2707536|T121|1008323|RXNORM|AMOXICILLIN / SULBACTAM|AMOXICILLIN / SULBACTAM
C2929229|T121|1008322|RXNORM|DECAMETHRIN / PIPERONYL BUTOXIDE|DECAMETHRIN / PIPERONYL BUTOXIDE
C2929228|T121|1008321|RXNORM|CAFFEINE / PHENYLEPHRINE|CAFFEINE / PHENYLEPHRINE
C2929227|T121|1008320|RXNORM|BIFONAZOLE / UREA|BIFONAZOLE / UREA
C2929233|T121|1008327|RXNORM|DEOXYCHOLATE / PEPSIN A|DEOXYCHOLATE / PEPSIN A
C2929232|T121|1008326|RXNORM|ASCORBIC ACID / RUTIN|ASCORBIC ACID / RUTIN
C2929231|T121|1008325|RXNORM|AMBROXOL / ASTEMIZOLE / BUTETHAMATE / PHENYLEPHRINE|AMBROXOL / ASTEMIZOLE / BUTETHAMATE / PHENYLEPHRINE
C2929230|T121|1008324|RXNORM|BILE SALTS / CYNARA PREPARATION|BILE SALTS / CYNARA PREPARATION
C2929234|T121|1008329|RXNORM|BENZOCAINE / PHENYLEPHRINE|BENZOCAINE / PHENYLEPHRINE
C2057677|T121|1008328|RXNORM|GUAIFENESIN / TETRACYCLINE|GUAIFENESIN / TETRACYCLINE
C0043328|T123|11359|RXNORM|LUTEIN|LUTEIN
C0069962|T168|32809|RXNORM|PALM OIL|PALM OIL
C3692843|T121|1442700|RXNORM|PRUNUS VIRGINIANA BARK EXTRACT|PRUNUS VIRGINIANA BARK EXTRACT
C3818726|T122|1534779|RXNORM|DI-N-OCTYL SODIUM SULFOSUCCINATE|DI-N-OCTYL SODIUM SULFOSUCCINATE
C3282035|T109|1312545|RXNORM|CETEARYL BEHENATE|CETEARYL BEHENATE
C0717852|T121|214646|RXNORM|HYDROFLUMETHIAZIDE / RESERPINE|HYDROFLUMETHIAZIDE / RESERPINE
C2348059|T130|1312547|RXNORM|D&C ORANGE NO. 5|D&C ORANGE NO. 5
C0055625|T197|1312546|RXNORM|CHROMIUM DIOXIDE|CHROMIUM DIOXIDE
C3496934|T121|1312541|RXNORM|ANIBA ROSAEODORA WOOD EXTRACT|ANIBA ROSAEODORA WOOD EXTRACT
C2698095|T121|1312540|RXNORM|AMMONIUM BENZOATE|AMMONIUM BENZOATE
C3473931|T121|1312543|RXNORM|BEHENYL BEHENATE|BEHENYL BEHENATE
C3497689|T121|1312542|RXNORM|ARCTIUM LAPPA WHOLE EXTRACT|ARCTIUM LAPPA WHOLE EXTRACT
C3475230|T121|1312549|RXNORM|DIETHYLENETRIAMINE PENTAMETHYLENE PHOSPHONIC ACID|DIETHYLENETRIAMINE PENTAMETHYLENE PHOSPHONIC ACID
C3465255|T121|1312548|RXNORM|DIACETYL BOLDINE|DIACETYL BOLDINE
C3693114|T109|1482549|RXNORM|BOS TAURUS BRAINSTEM PREPARATION|BOVINE BRAINSTEM PREPARATION
C3668958|T121|1482548|RXNORM|PRUNUS SPINOSA FRUIT EXTRACT|PRUNUS SPINOSA FRUIT EXTRACT
C0073188|T129|35465|RXNORM|RHO(D) IMMUNE GLOBULIN|ANTI-D (RH) IMMUNOGLOBULIN
C0718857|T121|215597|RXNORM|BELLADONNA ALKALOIDS / OPIUM|BELLADONNA ALKALOIDS / OPIUM
C3693109|T121|1482541|RXNORM|ARGANIA SPINOSA WHOLE EXTRACT|ARGANIA SPINOSA WHOLE EXTRACT
C3693108|T109|1482540|RXNORM|PPG-30|PPG-30
C3693111|T121|1482543|RXNORM|LEVISTICUM OFFICINALE ROOT EXTRACT|LEVISTICUM OFFICINALE ROOT EXTRACT
C3693110|T121|1482542|RXNORM|CELOSIA ARGENTEA SEED EXTRACT|CELOSIA ARGENTEA SEED EXTRACT
C0718858|T121|215598|RXNORM|BELLADONNA ALKALOIDS / ERGOTAMINE / PHENOBARBITAL|BELLADONNA ALKALOIDS / ERGOTAMINE / PHENOBARBITAL
C3669136|T121|1482544|RXNORM|PERSICARIA PUNCTATA EXTRACT|POLYGONUM PUNCTATUM EXTRACT
C3693113|T121|1482547|RXNORM|ASPLENIUM SCOLOPENDRIUM TOP EXTRACT|ASPLENIUM SCOLOPENDRIUM TOP EXTRACT
C0035588|T007|1482546|RXNORM|RICKETTSIA RICKETTSII|RICKETTSIA RICKETTSII
C0304925|T121|828529|RXNORM|ALBUMIN HUMAN, USP|ALBUMIN HUMAN, USP
C3859160|T121|1592263|RXNORM|BETA-D-RIBOSE|BETA-D-RIBOSE
C1698162|T109|1368211|RXNORM|3,7,11,15-TETRAMETHYL-1,2,3-HEXADECANETRIOL|3,7,11,15-TETRAMETHYL-1,2,3-HEXADECANETRIOL
C1959890|T121|729512|RXNORM|CINNARIZINE / DIMENHYDRINATE|CINNARIZINE / DIMENHYDRINATE
C1959978|T121|729513|RXNORM|CITRIC ACID / GLUCONOLACTONE / MAGNESIUM CARBONATE|CITRIC ACID / GLUCONOLACTONE / MAGNESIUM CARBONATE
C3256021|T109|1424360|RXNORM|BIOSACCHARIDE GUM-1|BIOSACCHARIDE GUM-1
C0005099|T121|1425|RXNORM|BENZYDAMINE|BENZYDAMINE
C0717618|T121|214421|RXNORM|CHOLINE / DEXPANTHENOL|CHOLINE / DEXPANTHENOL
C0717626|T121|214427|RXNORM|CITRIC ACID / POTASSIUM CITRATE|CITRIC ACID / POTASSIUM CITRATE
C3152834|T129|1098189|RXNORM|OSAGE ORANGE POLLEN EXTRACT|MACLURA POMIFERA POLLEN EXTRACT
C0062970|T123|27120|RXNORM|HORDENINE|HORDENINE
C3692932|T122|1442883|RXNORM|OLEALKONIUM CHLORIDE|OLEALKONIUM CHLORIDE
C2980835|T129|1098183|RXNORM|LARGEMOUTH BASS ALLERGENIC EXTRACT|LARGEMOUTH BASS ALLERGENIC EXTRACT
C0041441|T195|995505|RXNORM|TYLOSIN|TYLOSIN
C2073863|T121|819910|RXNORM|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / PHENYLEPHRINE|ACETAMINOPHEN / CAFFEINE / CHLORPHENIRAMINE / PHENYLEPHRINE
C2351042|T195|819911|RXNORM|BESIFLOXACIN|BESIFLOXACIN
C0991801|T197|317207|RXNORM|CALCIUM IODIZED|CALCIUM IODIZED
C2014107|T121|819919|RXNORM|ORPHENADRINE / PIROXICAM|ORPHENADRINE / PIROXICAM
C3486481|T197|1306098|RXNORM|ALUMINUM SULFATE TETRADECAHYDRATE|ALUMINUM SULFATE TETRADECAHYDRATE
C3256055|T109|1426290|RXNORM|HYPROMELLOSE ACETATE SUCCINATE 12070923 (3 MM2-S)|HYPROMELLOSE ACETATE SUCCINATE 12070923 (3 MM2-S)
C1337243|T121|1549114|RXNORM|ZINC ASCORBATE|ZINC ASCORBATE
C3855810|T121|1549115|RXNORM|1,2-DOCOSAHEXANOYL-SN-GLYCERO-3-PHOSPHOSERINE|1,2-DOCOSAHEXANOYL-SN-GLYCERO-3-PHOSPHOSERINE
C3855811|T121|1549116|RXNORM|1,2-DOCOSAHEXANOYL-SN-GLYCERO-3-PHOSPHOSERINE CALCIUM|1,2-DOCOSAHEXANOYL-SN-GLYCERO-3-PHOSPHOSERINE CALCIUM
C3855812|T121|1549117|RXNORM|1,2-ICOSAPENTOYL-SN-GLYCERO-3-PHOSPHOSERINE|1,2-ICOSAPENTOYL-SN-GLYCERO-3-PHOSPHOSERINE
C0074542|T197|1549110|RXNORM|SILVER SULFIDE|SILVER SULFIDE
C3853723|T121|1549111|RXNORM|TEUCRIUM SCORODONIA WHOLE EXTRACT|TEUCRIUM SCORODONIA WHOLE EXTRACT
C3859158|T121|1592261|RXNORM|SCIADOPITYS VERTICILLATA ROOT EXTRACT|SCIADOPITYS VERTICILLATA ROOT EXTRACT
C1329979|T129|404774|RXNORM|ANTHRAX VACCINE ADSORBED|ANTHRAX VACCINE ADSORBED
C3855813|T121|1549118|RXNORM|1,2-ICOSAPENTOYL-SN-GLYCERO-3-PHOSPHOSERINE CALCIUM|1,2-ICOSAPENTOYL-SN-GLYCERO-3-PHOSPHOSERINE CALCIUM
C2928149|T121|1007227|RXNORM|ACETAMINOPHEN / BUCLIZINE|ACETAMINOPHEN / BUCLIZINE
C0872910|T121|259277|RXNORM|POTASSIUM,CHELATED|POTASSIUM,CHELATED
C0872909|T121|259276|RXNORM|PINE BARK EXTRACT|PINE BARK EXTRACT
C3700876|T122|1487115|RXNORM|TRIDECYL LACTATE|TRIDECYL LACTATE
C0300892|T123|1487114|RXNORM|FARNESYL ACETATE|FARNESYL ACETATE
C3700875|T122|1487116|RXNORM|BENZYL PCA|BENZYL PCA
C0008996|T130|2592|RXNORM|SOY LECITHIN|CLOFAZIMINE
C2928478|T121|1007557|RXNORM|MELITRACEN / PERICIAZINE|MELITRACEN / PERICIAZINE
C2928146|T121|1007224|RXNORM|ASCORBIC ACID / FERROUS CHLORIDE|ASCORBIC ACID / FERROUS CHLORIDE
C1321596|T121|402316|RXNORM|MIGLUSTAT|MIGLUSTAT
C0025147|T125|6691|RXNORM|MEDROXYPROGESTERONE|MEDROXYPROGESTERONE
C0025147|T125|6691|RXNORM|MEDROXYPROGESTERONE|MEDROXYPROGESTERONE
C0025145|T125|6690|RXNORM|MEDROGESTONE|MEDROGESTONE
C0025156|T121|6696|RXNORM|MEFRUSIDE|MEFRUSIDE
C0025153|T121|6694|RXNORM|MEFLOQUINE|MEFLOQUINE
C2929710|T121|1008811|RXNORM|BENZOATE / PHENYLACETATE|BENZOATE / PHENYLACETATE
C2929709|T121|1008810|RXNORM|FORMALDEHYDE / MALACHITE GREEN|FORMALDEHYDE / MALACHITE GREEN
C2929712|T121|1008813|RXNORM|DEXTRAN 70 / POLYETHYLENE GLYCOL 400 / POVIDONE / TETRAHYDROZOLINE|DEXTRAN 70 / POLYETHYLENE GLYCOL 400 / POVIDONE / TETRAHYDROZOLINE
C2929711|T121|1008812|RXNORM|CODEINE / GUAIACOLSULFONIC ACID / PROMETHAZINE|CODEINE / GUAIACOLSULFONIC ACID / PROMETHAZINE
C2929714|T121|1008815|RXNORM|SULFAMETHAZINE / TRIMETHOPRIM|SULFAMETHAZINE / TRIMETHOPRIM
C0113293|T121|48937|RXNORM|DEXMEDETOMIDINE|DEXMEDETOMIDINE
C2929716|T121|1008817|RXNORM|ASCORBIC ACID / ECHINACEA PREPARATION|ASCORBIC ACID / ECHINACEA PREPARATION
C2929715|T121|1008816|RXNORM|CHLORMADINONE / MESTRANOL|CHLORMADINONE / MESTRANOL
C2929718|T121|1008819|RXNORM|CAPSAICIN / TROLAMINE SALICYLATE|CAPSAICIN / TROLAMINE SALICYLATE
C2929717|T121|1008818|RXNORM|LIDOCAINE / MENTHOL|LIDOCAINE / MENTHOL
C2928473|T121|1007552|RXNORM|ALOE POLYSACCHARIDE / IODOQUINOL|ALOE POLYSACCHARIDE / IODOQUINOL
C1871526|T121|719872|RXNORM|RALTEGRAVIR|RALTEGRAVIR
C2979691|T197|1306097|RXNORM|ALUMINUM ZIRCONIUM PENTACHLOROHYDRATE|ALUMINUM ZIRCONIUM PENTACHLOROHYDRATE
C3464349|T121|1291859|RXNORM|AZELASTINE / FLUTICASONE|AZELASTINE / FLUTICASONE
C0030140|T121|7839|RXNORM|P-HYDROXYAMPHETAMINE|P-HYDROXYAMPHETAMINE
C3833033|T121|1540238|RXNORM|BRASSICA RAPA SUBSP. RAPA SEED EXTRACT|BRASSICA RAPA SUBSP. RAPA SEED EXTRACT
C3833034|T121|1540239|RXNORM|LAVANDULA STOECHAS WHOLE EXTRACT|LAVANDULA STOECHAS WHOLE EXTRACT
C0054202|T121|19832|RXNORM|BUDIPINE|BUDIPINE
C0054201|T121|19831|RXNORM|BUDESONIDE|BUDESONIDE
C0054201|T121|19831|RXNORM|BUDESONIDE|BUDESONIDE
C0054201|T121|19831|RXNORM|BUDESONIDE|BUDESONIDE
C0030123|T130|7832|RXNORM|4-AMINOHIPPURIC ACID|4-AMINOHIPPURIC ACID
C0030125|T121|7833|RXNORM|AMINOSALICYLIC ACID|AMINOSALICYLIC ACID
C0771378|T121|236133|RXNORM|SPONGIA TOSTA|SPONGIA TOSTA
C0075518|T121|37333|RXNORM|SULFANILYLUREA|SULFANILYLUREA
C1166067|T121|350376|RXNORM|SEPIA EXTRACT|SEPIA EXTRACT
C0127615|T121|52582|RXNORM|MESALAMINE|MESALAMINE
C0127615|T121|52582|RXNORM|MESALAMINE|MESALAMINE
C0038686|T195|10178|RXNORM|SULFAMETHAZINE|SULFAMETHAZINE
C0038687|T121|10179|RXNORM|SULFAMETHIZOLE|SULFAMETHIZOLE
C3531212|T121|1366328|RXNORM|ORCHIS MASCULA WHOLE EXTRACT|ORCHIS MASCULA WHOLE EXTRACT
C3531213|T121|1366329|RXNORM|ORYZA SATIVA WHOLE EXTRACT|ORYZA SATIVA WHOLE EXTRACT
C3531207|T109|1366322|RXNORM|CERATONIA SILIQUA WHOLE EXTRACT|CERATONIA SILIQUA WHOLE EXTRACT
C0038675|T195|10171|RXNORM|SULFADIAZINE|SULFADIAZINE
C0038676|T195|10172|RXNORM|SULFADIMETHOXINE|SULFADIMETHOXINE
C0038679|T121|10173|RXNORM|SULFADOXINE|SULFADOXINE
C0038681|T195|10174|RXNORM|SULFAGUANIDINE|SULFAGUANIDINE
C0038683|T121|10175|RXNORM|SULFALENE|SULFALENE
C0038684|T121|10176|RXNORM|SULFAMERAZINE|SULFAMERAZINE
C3531209|T109|1366325|RXNORM|COIX LACRYMA-JOBI SEED OIL|COIX LACRYMA-JOBI SEED OIL
C0060926|T121|25480|RXNORM|GABAPENTIN|GABAPENTIN
C0060926|T121|25480|RXNORM|GABAPENTIN|GABAPENTIN
C0055894|T121|21244|RXNORM|CLOBENZOREX|CLOBENZOREX
C0056464|T123|21716|RXNORM|CRATAEGUS EXTRACT|CRATAEGUS EXTRACT
C0055891|T121|21241|RXNORM|CLOBAZAM|CLOBAZAM
C3473104|T121|1298158|RXNORM|CALCIUM CARBONATE / FOLIC ACID|CALCIUM CARBONATE / FOLIC ACID
C0055899|T125|21249|RXNORM|CLOCORTOLONE|CLOCORTOLONE
C2146445|T121|818205|RXNORM|RIFAMPIN / TRIMETHOPRIM|RIFAMPIN / TRIMETHOPRIM
C2733369|T121|901212|RXNORM|AMLODIPINE / TELMISARTAN|AMLODIPINE / TELMISARTAN
C0060930|T130|25483|RXNORM|GADOTERIDOL|GADOTERIDOL
C0047625|T109|1484499|RXNORM|3-BUTYLPHTHALIDE|3-N-BUTYLPHTHALIDE
C3527960|T121|1361462|RXNORM|SUS SCROFA LARGE INTESTINE PREPARATION|SUS SCROFA LARGE INTESTINE PREPARATION
C3818688|T121|1537752|RXNORM|PAPAYA SEED EXTRACT|PAPAYA SEED EXTRACT
C0057236|T109|1484495|RXNORM|DECANAL|DECANAL
C3695958|T109|1484494|RXNORM|BILBERRY SEED OIL|BILBERRY SEED OIL
C0662731|T109|1484497|RXNORM|FARNESAL|FARNESAL
C3527961|T121|1361463|RXNORM|TYLOPHORA INDICA WHOLE EXTRACT|TYLOPHORA INDICA WHOLE EXTRACT
C1873970|T121|689585|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE / SALICYLAMIDE|ACETAMINOPHEN / CHLORPHENIRAMINE / PHENYLEPHRINE / SALICYLAMIDE
C0006376|T121|1808|RXNORM|BUMETANIDE|BUMETANIDE
C0082787|T121|41208|RXNORM|HALOBETASOL|HALOBETASOL
C3486392|T121|1350999|RXNORM|DAPHNE MEZEREUM BARK EXTRACT|DAPHNE MEZEREUM BARK EXTRACT
C1113058|T121|324051|RXNORM|METHYLENEDIOXYCINNAMIC ACID|METHYLENEDIOXYCINNAMIC ACID
C0060934|T130|25486|RXNORM|GADOPENTETATE DIMEGLUMINE|GADOPENTETATE DIMEGLUMINE
C2701066|T129|851732|RXNORM|ACACIA POLLEN EXTRACT|ACACIA POLLEN EXTRACT
C3700887|T168|1486793|RXNORM|LOWBUSH BLUEBERRY JUICE|LOWBUSH BLUEBERRY JUICE
C2701070|T129|851736|RXNORM|COAST MAPLE POLLEN EXTRACT|ACER MACROPHYLLUM POLLEN EXTRACT
C2701132|T129|851882|RXNORM|SISAL FIBER EXTRACT|AGAVE SISALANA FIBER EXTRACT
C2348465|T121|1332872|RXNORM|EQUISETUM HYEMALE EXTRACT|EQUISETUM HYEMALE EXTRACT
C3700886|T168|1486794|RXNORM|STRAWBERRY JUICE|FRAGARIA ANANASSA JUICE
C3700885|T122|1486795|RXNORM|POLYGLYCERIN-4|POLYGLYCERIN-4
C0115510|T121|49428|RXNORM|EDOXUDINE|EDOXUDINE
C3190643|T121|1144963|RXNORM|ASCORBATE MANGANESE / CHONDROITIN SULFATES / GLUCOSAMINE|ASCORBATE MANGANESE / CHONDROITIN SULFATES / GLUCOSAMINE
C0772022|T121|1144960|RXNORM|ASCORBATE MANGANESE|ASCORBATE MANGANESE
C1144403|T121|1547611|RXNORM|ORITAVANCIN|ORITAVANCIN
C1572754|T121|1547610|RXNORM|MORRHUATE|MORRHUATE
C3163249|T121|1115951|RXNORM|WHITE SWEET CLOVER POLLEN EXTRACT / YELLOW SWEET CLOVER POLLEN EXTRACT|WHITE SWEET CLOVER POLLEN EXTRACT / YELLOW SWEET CLOVER POLLEN EXTRACT
C1719936|T121|645168|RXNORM|MAGNESIUM HYDROXIDE / OMEPRAZOLE / SODIUM BICARBONATE|MAGNESIUM HYDROXIDE / OMEPRAZOLE / SODIUM BICARBONATE
C0010566|T109|1367180|RXNORM|CYCLOHEXANE|CYCLOHEXANE
C0020270|T197|1367183|RXNORM|HYDROGEN CYANIDE|HYDROGEN CYANIDE
C0019225|T109|1367182|RXNORM|HEPTANES|HEPTANES
C0021760|T129|1367185|RXNORM|INTERLEUKIN-6|INTERLEUKIN-6
C0021759|T129|1367184|RXNORM|INTERLEUKIN-5|INTERLEUKIN-5
C0087161|T127|1367187|RXNORM|ALL-TRANS-RETINOL|ALL-TRANS-RETINOL
C0039541|T196|1367186|RXNORM|TERBIUM|TERBIUM
C3255605|T109|1367189|RXNORM|NONOXYNOL-20|NONOXYNOL-20
C0011701|T125|3251|RXNORM|DESMOPRESSIN|DESMOPRESSIN
C0011705|T121|3254|RXNORM|DESONIDE|DESONIDE
C0011707|T125|3255|RXNORM|DESOXIMETASONE|DESOXIMETASONE
C0011710|T125|3256|RXNORM|DEOXYCORTICOSTERONE|DESOXYCORTICOSTERONE
C1875825|T121|690767|RXNORM|TETRAHYDROZOLINE / ZINC SULFATE|TETRAHYDROZOLINE / ZINC SULFATE
C3700901|T109|1486029|RXNORM|BEHENAMIDOPROPYL DIMETHYLAMINE BEHENATE|BEHENAMIDOPROPYL DIMETHYLAMINE BEHENATE
C0072864|T125|35215|RXNORM|QUINESTRADOL|QUINESTRADOL
C0062527|T129|797752|RXNORM|HEPATITIS B SURFACE ANTIGEN VACCINE|HEPATITIS B SURFACE ANTIGEN VACCINE
C0054433|T121|1311397|RXNORM|CAFFEIC ACID|CAFFEIC ACID
C0024469|T121|1311396|RXNORM|MAGNESIUM ASCORBATE|MAGNESIUM ASCORBATE
C0068808|T197|1311391|RXNORM|NITRIC ACID|NITRIC ACID
C0036179|T121|1311390|RXNORM|SANTONIN|SANTONIN
C0242864|T109|1311393|RXNORM|AMBER|AMBER
C3486777|T121|1311392|RXNORM|PORK INTESTINE PREPARATION|SUS SCROFA INTESTINE PREPARATION
C3255772|T109|1426436|RXNORM|HOREHOUND EXTRACT|HOREHOUND EXTRACT
C1271556|T121|388053|RXNORM|LATANOPROST / TIMOLOL|LATANOPROST / TIMOLOL
C3472925|T121|1311399|RXNORM|DRIMIA MARITIMA BULB EXTRACT|DRIMIA MARITIMA BULB EXTRACT
C1095900|T121|1311398|RXNORM|LOBELIA SPICATA LEAF EXTRACT|LOBELIA SPICATA LEAF EXTRACT
C2073848|T121|823294|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN|CHLORPHENIRAMINE / DEXTROMETHORPHAN / GUAIFENESIN
C0012030|T121|3332|RXNORM|DIBENZEPIN|DIBENZEPIN
C0019142|T121|5228|RXNORM|HEPARINOIDS|HEPARINOIDS
C0020197|T126|5464|RXNORM|HYALURONIDASE|HYALURONIDASE
C0072865|T121|35216|RXNORM|QUINFAMIDE|QUINFAMIDE
C0012050|T121|3339|RXNORM|DIBUCAINE|DIBUCAINE
C2701766|T129|852738|RXNORM|EASTERN WHITE PINE POLLEN EXTRACT|PINUS STROBUS POLLEN EXTRACT
C2928804|T121|1007890|RXNORM|POTASSIUM IODIDE / THYROXINE|LEVOTHYROXINE / POTASSIUM IODIDE
C2928806|T121|1007892|RXNORM|METHENAMINE / SODIUM PHOSPHATE, MONOBASIC|METHENAMINE / SODIUM PHOSPHATE, MONOBASIC
C2928807|T121|1007893|RXNORM|BELLADONNA ALKALOIDS / CAFFEINE / ERGOTAMINE / PENTOBARBITAL|BELLADONNA ALKALOIDS / CAFFEINE / ERGOTAMINE / PENTOBARBITAL
C2928808|T121|1007894|RXNORM|ASCORBIC ACID / VITAMIN A / VITAMIN E / ZINC SULFATE|ASCORBIC ACID / VITAMIN A / VITAMIN E / ZINC SULFATE
C2928809|T121|1007895|RXNORM|BRYONIA PREPARATION / HYDRASTIS PREPARATION / YELLOW PHENOLPHTHALEIN|BRYONIA PREPARATION / HYDRASTIS PREPARATION / YELLOW PHENOLPHTHALEIN
C2928810|T121|1007896|RXNORM|ASCORBIC ACID / MAGNESIUM SULFATE / VITAMIN E / ZINC SULFATE|ASCORBIC ACID / MAGNESIUM SULFATE / VITAMIN E / ZINC SULFATE
C2928811|T121|1007897|RXNORM|ASCORBIC ACID / FERROUS BISGLYCINATE / FOLIC ACID / VITAMIN B 12|ASCORBIC ACID / FERROUS BISGLYCINATE / FOLIC ACID / VITAMIN B 12
C2928812|T121|1007898|RXNORM|CETYL ALCOHOL / COLFOSCERIL|CETYL ALCOHOL / COLFOSCERIL
C2928813|T121|1007899|RXNORM|ARGININE / CALCIUM CARBONATE / MACA PREPARATION|ARGININE / CALCIUM CARBONATE / MACA PREPARATION
C3256246|T121|1307844|RXNORM|PERSEA AMERICANA LEAF EXTRACT|PERSEA AMERICANA LEAF EXTRACT
C3644290|T121|1424560|RXNORM|PEPPERMINT OIL / SAGE OIL|PEPPERMINT OIL / SAGE OIL
C3256586|T121|1307842|RXNORM|ACTINIDIA CHINENSIS SEED EXTRACT|ACTINIDIA CHINENSIS SEED EXTRACT
C3256365|T109|1307843|RXNORM|MORINDA CITRIFOLIA SEED OIL|MORINDA CITRIFOLIA SEED OIL
C0055149|T122|1307840|RXNORM|CETOSTEARYL ALCOHOL|CETOSTEARYL ALCOHOL
C3255850|T121|1307841|RXNORM|MAACKIA FLORIBUNDA STEM EXTRACT|MAACKIA FLORIBUNDA STEM EXTRACT
C0609416|T121|1310554|RXNORM|ETHYL CITRATE|ETHYL CITRATE
C1273023|T121|1363569|RXNORM|DIMETHICONE 350|DIMETHICONE 350
C1444947|T122|1363568|RXNORM|CARBOMER-974P|CARBOMER-974P
C0006474|T121|1310550|RXNORM|BUTANE|BUTANE
C3528889|T121|1363563|RXNORM|TRIFOLIUM REPENS POLLEN EXTRACT|TRIFOLIUM REPENS POLLEN EXTRACT
C3528888|T121|1363562|RXNORM|RUMEX ACETOSA WHOLE EXTRACT|RUMEX ACETOSA WHOLE EXTRACT
C2827593|T129|1363561|RXNORM|AMARANTHUS HYBRIDUS POLLEN EXTRACT|AMARANTHUS HYBRIDUS POLLEN EXTRACT
C0001898|T123|426|RXNORM|ALANINE|ALANINE
C3256161|T130|1310558|RXNORM|FD & C RED NO. 40 ALUMINUM LAKE|FD & C RED NO. 40 ALUMINUM LAKE
C3257193|T130|1310559|RXNORM|D&C RED NO. 27 ALUMINUM LAKE|D&C RED NO. 27 ALUMINUM LAKE
C3528890|T109|1363565|RXNORM|DECYL PALMITATE|DECYL PALMITATE
C0982100|T120|1311171|RXNORM|D & C GREEN 5|D&C GREEN NO. 5
C3497905|T121|1311170|RXNORM|BEEF KIDNEY PREPARATION|BEEF KIDNEY PREPARATION
C0035890|T121|1314413|RXNORM|ROXARSONE|ROXARSONE
C0205892|T120|1311172|RXNORM|D & C RED NO. 27|D & C RED NO. 27
C1533427|T122|1314415|RXNORM|ISOPROPYL ISOSTEARATE|ISOPROPYL ISOSTEARATE
C0301298|T121|89717|RXNORM|THYMOL IODIDE|THYMOL IODIDE
C3489150|T121|1311177|RXNORM|GONORRHEAL URETHRAL SECRETION HUMAN|GONORRHEAL URETHRAL SECRETION HUMAN
C0982104|T120|1311176|RXNORM|D&C RED NO. 30|D&C RED NO. 30
C0064058|T121|1311179|RXNORM|ISOPROPYL PALMITATE|ISOPROPYL PALMITATE
C1509303|T120|1311178|RXNORM|D&C RED NO. 6|D&C RED NO. 6
C3464615|T121|1292760|RXNORM|DOCOSAHEXAENOATE / LUTEIN / VITAMIN E|DOCOSAHEXAENOATE / LUTEIN / VITAMIN E
C0766026|T121|233562|RXNORM|HELICIDINE|HELICIDINE
C0005098|T121|1424|RXNORM|GENTAMICIN SULFATE (USP)|BENZTROPINE
C0005098|T121|1424|RXNORM|GENTAMICIN SULFATE (USP)|BENZTROPINE
C0005098|T121|1424|RXNORM|GENTAMICIN SULFATE (USP)|BENZTROPINE
C1453100|T121|1433192|RXNORM|GLUCOSYL HESPERIDIN|GLUCOSYL HESPERIDIN
C3163603|T129|1116738|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED A-CHRISTCHURCH-16-2010 NIB-74 (H1N1) (A-CALIFORNIA-7-2009) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED A-CHRISTCHURCH-16-2010 NIB-74 (H1N1) (A-CALIFORNIA-7-2009) STRAIN
C3486698|T121|1331705|RXNORM|BOTRYOGLOSSUM PLATYCARPUM EXTRACT|BOTRYOGLOSSUM PLATYCARPUM EXTRACT
C2928021|T121|1007098|RXNORM|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / LIVER STOMACH CONCENTRATE / VITAMIN B 12|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / LIVER STOMACH CONCENTRATE / VITAMIN B 12
C2928022|T121|1007099|RXNORM|DEHYDROCHOLATE / DIMETHICONE / PANCREATIN|DEHYDROCHOLATE / DIMETHICONE / PANCREATIN
C3645194|T109|1426846|RXNORM|HYPROMELLOSE 2906 (4 MPA.S)|HYPROMELLOSE 2906 (4 MPA.S)
C0005100|T121|1426|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-VICTORIA-361-2011 (H3N2) STRAIN|BENZYL ALCOHOL
C2928013|T121|1007090|RXNORM|POLYETHYLENE GLYCOL 400 / POLYVINYL ALCOHOL|POLYETHYLENE GLYCOL 400 / POLYVINYL ALCOHOL
C2928014|T121|1007091|RXNORM|PECAN POLLEN EXTRACT / WHITE HICKORY POLLEN EXTRACT|PECAN POLLEN EXTRACT / WHITE HICKORY POLLEN EXTRACT
C2928015|T121|1007092|RXNORM|PSYLLIUM / SENNOSIDES, USP|PSYLLIUM / SENNOSIDES, USP
C2928017|T121|1007094|RXNORM|ACETIC ACID / OXYQUINOLINE / RICINOLEATE|ACETIC ACID / OXYQUINOLINE / RICINOLEATE
C2928018|T121|1007095|RXNORM|ACETIC ACID / GLYCERIN / OXYQUINOLINE / RICINOLEATE|ACETIC ACID / GLYCERIN / OXYQUINOLINE / RICINOLEATE
C2928019|T121|1007096|RXNORM|CETYLPYRIDINIUM / SODIUM FLUORIDE|CETYLPYRIDINIUM / SODIUM FLUORIDE
C2928020|T121|1007097|RXNORM|DEHYDROCHOLATE / PANCREATIN / PEPSIN A|DEHYDROCHOLATE / PANCREATIN / PEPSIN A
C3811620|T109|1535698|RXNORM|DANDELION HONEY|DANDELION HONEY
C3811677|T129|1541617|RXNORM|INFLUENZA A VIRUS VACCINE, A-TEXAS-50-2012 (H3N2)-LIKE VIRUS|INFLUENZA A VIRUS VACCINE, A-TEXAS-50-2012 (H3N2)-LIKE VIRUS
C0287721|T195|83719|RXNORM|GREPAFLOXACIN|GREPAFLOXACIN
C0981884|T129|867228|RXNORM|FUSARIUM OXYSPORUM VASINFECTUM EXTRACT|FUSARIUM OXYSPORUM VASINFECTUM EXTRACT
C0002164|T121|528|RXNORM|ALMITRINE|ALMITRINE
C0877880|T129|262323|RXNORM|IBRITUMOMAB TIUXETAN|IBRITUMOMAB TIUXETAN
C0064585|T121|28395|RXNORM|LACTITOL|LACTITOL
C0202474|T131|66422|RXNORM|STRYCHNINE|STRYCHNINE
C0301421|T121|89821|RXNORM|WITCH HAZEL|WITCH HAZEL
C1141247|T121|340398|RXNORM|IOPANOATE SODIUM|IOPANOATE SODIUM
C0063739|T109|27712|RXNORM|INVERT SUGAR|MAIZE INVERT SUGAR
C0063739|T109|27712|RXNORM|INVERT SUGAR|MAIZE INVERT SUGAR
C2928157|T121|1007235|RXNORM|BROMELAINS / PAPAIN / TRYPSIN|BROMELAINS / PAPAIN / TRYPSIN
C2928158|T121|1007236|RXNORM|CYCLOTHIAZIDE / TRIAMTERENE|CYCLOTHIAZIDE / TRIAMTERENE
C2928467|T121|1007546|RXNORM|ALANINE / ARGININE / ASPARTATE / GLUCOSE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / SODIUM PHOSPHATE / THREONINE / TRYPTOP|ALANINE / ARGININE / ASPARTATE / GLUCOSE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / POTASSIUM CHLORIDE / PROLINE / SERINE / SODIUM CHLORIDE / SODIUM PHOSPHATE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2928153|T121|1007231|RXNORM|ASCORBIC ACID / THIAMINE|ASCORBIC ACID / THIAMINE
C2928465|T121|1007544|RXNORM|ASCORBIC ACID / POLYETHYLENE GLYCOL 3350 / POTASSIUM CHLORIDE / SODIUM ASCORBATE / SODIUM CHLORIDE / SODIUM SULFATE|ASCORBIC ACID / POLYETHYLENE GLYCOL 3350 / POTASSIUM CHLORIDE / SODIUM ASCORBATE / SODIUM CHLORIDE / SODIUM SULFATE
C2928466|T121|1007545|RXNORM|ACELLULAR PERTUSSIS VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / HEPATITIS B SURFACE ANTIGEN VACCINE / POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY) / POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1) / POLIOVIRUS VACCINE INACTIVATED, T|ACELLULAR PERTUSSIS VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / HEPATITIS B SURFACE ANTIGEN VACCINE / POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY) / POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1) / POLIOVIRUS VACCINE INACTIVATED, TYPE 3 (SAUKETT) / TETANUS TOXOID VACCINE, INACTIVATED
C2928469|T121|1007548|RXNORM|FE HEME POLYPEPTIDE / POLYSACCHARIDE IRON COMPLEX|FE HEME POLYPEPTIDE / POLYSACCHARIDE IRON COMPLEX
C2928470|T121|1007549|RXNORM|BENZOCAINE / PYRILAMINE / ZINC OXIDE|BENZOCAINE / PYRILAMINE / ZINC OXIDE
C2928160|T121|1007238|RXNORM|ACONITE / CODEINE / ERYSIMUM PREPARATION|ACONITE / CODEINE / ERYSIMUM PREPARATION
C2928161|T121|1007239|RXNORM|FORMALDEHYDE / LIDOCAINE|FORMALDEHYDE / LIDOCAINE
C1875489|T121|691142|RXNORM|METHYCLOTHIAZIDE / PARGYLINE|METHYCLOTHIAZIDE / PARGYLINE
C1875490|T121|691144|RXNORM|METHYL ANTHRANILATE / TITANIUM DIOXIDE|METHYL ANTHRANILATE / TITANIUM DIOXIDE
C0017066|T121|4678|RXNORM|GANCICLOVIR|GANCICLOVIR
C0017066|T121|4678|RXNORM|GANCICLOVIR|GANCICLOVIR
C0066082|T195|29629|RXNORM|METHAMPICILLIN|METAMIPICILLIN
C3864969|T121|1597093|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 11 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 16 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 31 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 33 VACCINE /|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 11 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 16 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 18 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 31 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 33 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 45 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 52 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 58 VACCINE / L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 6 VACCINE
C3248810|T121|1233902|RXNORM|CAFFEINE / DIHYDROERGOCRYPTINE|CAFFEINE / DIHYDROERGOCRYPTINE
C2701170|T129|851930|RXNORM|REDROOT PIGWEED POLLEN EXTRACT|AMARANTHUS RETROFLEXUS POLLEN EXTRACT
C1654195|T121|607464|RXNORM|DEXCHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE|DEXCHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE
C3535646|T109|1370110|RXNORM|ZINC ACETYLMETHIONATE|ZINC ACETYLMETHIONATE
C1178580|T121|360375|RXNORM|FENUGREEK SEED PREPARATION|FENUGREEK SEED PREPARATION
C0032333|T121|8462|RXNORM|PODOPHYLLIN|PODOPHYLLIN
C0032334|T131|8463|RXNORM|PODOFILOX|PODOFILOX
C0937858|T130|283753|RXNORM|PERFLUTREN|PERFLUTREN
C0677667|T121|196239|RXNORM|RALTITREXED|RALTITREXED
C2929490|T121|1008587|RXNORM|CHLOROPHYLLIN / THYMOL|CHLOROPHYLLIN / THYMOL
C0873128|T121|259462|RXNORM|LUTEIN ESTERS|LUTEIN ESTERS
C0245179|T121|72467|RXNORM|TIRILAZAD|TIRILAZAD
C1720087|T121|645184|RXNORM|CYCLIZINE / MORPHINE|CYCLIZINE / MORPHINE
C3195298|T121|1119628|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / PHYTOSTEROL ESTERS|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / PHYTOSTEROL ESTERS
C3531376|T109|1366669|RXNORM|PEG-6 ISOSTEARATE|PEG-6 ISOSTEARATE
C3531375|T109|1366668|RXNORM|PEG-15 COCAMINE|PEG-15 COCAMINE
C0072185|T121|1366667|RXNORM|PROPIONAMIDE|PROPIONAMIDE
C0035871|T131|1366666|RXNORM|ROTENONE|ROTENONE
C3531374|T121|1366665|RXNORM|HESPERETIN LAURATE|HESPERETIN LAURATE
C1881893|T121|1366664|RXNORM|GLYCERYL CAPRATE|GLYCERYL CAPRATE
C2928790|T121|1007876|RXNORM|ESCIN / NYLIDRIN|ESCIN / NYLIDRIN
C0059849|T121|24591|RXNORM|ETHYNODIOL|ETYNODIOL
C3535648|T109|1370107|RXNORM|DIBUTYL ETHYLHEXANOYL GLUTAMIDE|DIBUTYL ETHYLHEXANOYL GLUTAMIDE
C2928791|T121|1007877|RXNORM|CREOSOTE / GUAIACOL / METHYL SALICYLATE|CREOSOTE / GUAIACOL / METHYL SALICYLATE
C2081459|T121|818190|RXNORM|ACETAMINOPHEN / PIROXICAM|ACETAMINOPHEN / PIROXICAM
C0753645|T195|228476|RXNORM|GATIFLOXACIN|GATIFLOXACIN
C0753645|T195|228476|RXNORM|GATIFLOXACIN|GATIFLOXACIN
C0053618|T131|19338|RXNORM|BIOALLETHRIN|BIOALLETHRIN
C2928789|T121|1007875|RXNORM|CALAMINE / RESORCINOL / SULFUR,COLLOIDAL|CALAMINE / RESORCINOL / SULFUR,COLLOIDAL
C2928612|T121|1007696|RXNORM|PAMABROM / PYRILAMINE|PAMABROM / PYRILAMINE
C0069739|T121|32613|RXNORM|OXAPROZIN|OXAPROZIN
C2194207|T121|1007873|RXNORM|FOLIC ACID / LIVER EXTRACT|FOLIC ACID / LIVER EXTRACT
C2928610|T121|1007694|RXNORM|NORFENEFRINE / OCTODRINE|NORFENEFRINE / OCTODRINE
C2348248|T121|816346|RXNORM|DEXLANSOPRAZOLE|DEXLANSOPRAZOLE
C2073885|T121|813265|RXNORM|CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE|CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE
C0129044|T121|52918|RXNORM|MOXAVERINE|MOXAVERINE
C3651741|T121|1429914|RXNORM|ACRYLIC ACID-SODIUM ACRYLATE COPOLYMER (1:1; 600 MPA.S AT 0.2%)|ACRYLIC ACID-SODIUM ACRYLATE COPOLYMER (1:1; 600 MPA.S AT 0.2%)
C0015131|T121|4177|RXNORM|ETOMIDATE|ETOMIDATE
C0015120|T121|4171|RXNORM|ETIDOCAINE|ETIDOCAINE
C0015133|T121|4179|RXNORM|ETOPOSIDE|ETOPOSIDE
C1165801|T129|350141|RXNORM|SACCHAROMYCES CEREVISIAE ALLERGENIC EXTRACT|SACCHAROMYCES CEREVISIAE ALLERGENIC EXTRACT
C3556193|T121|1376005|RXNORM|FOLIC ACID / SUCCINIC ACID|FOLIC ACID / SUCCINIC ACID
C0717561|T121|214364|RXNORM|CARBINOXAMINE / PSEUDOEPHEDRINE|CARBINOXAMINE / PSEUDOEPHEDRINE
C0526513|T121|135098|RXNORM|DALFOPRISTIN / QUINUPRISTIN|DALFOPRISTIN / QUINUPRISTIN
C0717564|T121|214367|RXNORM|CASANTHRANOL / DOCUSATE|CASANTHRANOL / DOCUSATE
C0027999|T121|7394|RXNORM|NIALAMIDE|NIALAMIDE
C3256593|T121|1307543|RXNORM|AGAVE TEQUILANA LEAF EXTRACT|AGAVE TEQUILANA LEAF EXTRACT
C3256098|T121|1307542|RXNORM|ASTROCARYUM MURUMURU SEED BUTTER EXTRACT|ASTROCARYUM MURUMURU SEED BUTTER EXTRACT
C3255949|T121|1307541|RXNORM|MAGNOLIA VIRGINIANA FLOWER EXTRACT|MAGNOLIA VIRGINIANA FLOWER EXTRACT
C3282868|T121|1307540|RXNORM|VIOLA ODORATA FLOWERING TOP EXTRACT|VIOLA ODORATA FLOWERING TOP EXTRACT
C3256666|T121|1307547|RXNORM|CAMELLIA JAPONICA FLOWER EXTRACT|CAMELLIA JAPONICA FLOWER EXTRACT
C3473229|T121|1307545|RXNORM|MORUS ALBA STEM EXTRACT|MORUS ALBA STEM EXTRACT
C0526510|T121|135095|RXNORM|ASPIRIN / CODEINE|ASPIRIN / CODEINE
C0057678|T121|22759|RXNORM|DIACETYLRHEIN|DIACEREIN
C2701459|T129|852264|RXNORM|CURVULARIA EXTRACT|COCHLIOBOLUS LUNATUS EXTRACT
C0875927|T121|261418|RXNORM|HYOSCYAMINE / PHENOBARBITAL|HYOSCYAMINE / PHENOBARBITAL
C2701455|T129|852260|RXNORM|BLACK OAK POLLEN EXTRACT|QUERCUS VELUTINA POLLEN EXTRACT
C2348058|T109|1544393|RXNORM|D&C ORANGE NO. 11|D&C ORANGE NO. 11
C2698692|T121|1544460|RXNORM|IDELALISIB|IDELALISIB
C0875926|T121|261417|RXNORM|HYDROCHLOROTHIAZIDE / QUINAPRIL|HYDROCHLOROTHIAZIDE / QUINAPRIL
C0875921|T121|261414|RXNORM|ESTRADIOL / NORGESTIMATE|ESTRADIOL / NORGESTIMATE
C0875922|T121|261415|RXNORM|FOSINOPRIL / HYDROCHLOROTHIAZIDE|FOSINOPRIL / HYDROCHLOROTHIAZIDE
C3530450|T109|1364403|RXNORM|IRVINGIA GABONENSIS SEED BUTTER EXTRACT|IRVINGIA GABONENSIS SEED BUTTER EXTRACT
C3530451|T121|1364404|RXNORM|LONG PEPPER EXTRACT|LONG PEPPER EXTRACT
C3530453|T121|1364407|RXNORM|VIOLA ODORATA LEAF EXTRACT|VIOLA ODORATA LEAF EXTRACT
C3484626|T109|1312544|RXNORM|BIDENS BIPINNATA WHOLE EXTRACT|BIDENS BIPINNATA WHOLE EXTRACT
C3651698|T122|1431997|RXNORM|QUATERNIUM-18 HECTORITE|QUATERNIUM-18 HECTORITE
C3695952|T129|1484984|RXNORM|ENGLISH OAK POLLEN EXTRACT|QUERCUS ROBUR POLLEN EXTRACT
C0304125|T109|1431992|RXNORM|CALAMUS OIL|CALAMUS OIL
C0257685|T121|77655|RXNORM|ZOLEDRONIC ACID|ZOLEDRONIC ACID
C0021936|T130|5924|RXNORM|INULIN|INULIN
C0021936|T130|5924|RXNORM|INULIN|INULIN
C0600370|T121|155080|RXNORM|METHACHOLINE|METHACHOLINE
C0021918|T123|5920|RXNORM|INTRINSIC FACTOR|INTRINSIC FACTOR
C0304984|T197|91537|RXNORM|IOTHALAMATE SODIUM I125|SODIUM IOTHALAMATE (125I)
C0021961|T130|5928|RXNORM|IODAMIDE|IODAMIDE
C3643364|T109|1421446|RXNORM|PIPER BETLE LEAF EXTRACT|PIPER BETLE LEAF EXTRACT
C3486068|T121|1328307|RXNORM|RANUNCULUS BULBOSUS EXTRACT|RANUNCULUS BULBOSUS EXTRACT
C0304982|T197|91535|RXNORM|SODIUM IODIDE I131|SODIUM IODIDE I131
C3486692|T121|1328308|RXNORM|ALPINE STRAWBERRY EXTRACT|FRAGARIA VESCA FRUIT EXTRACT
C3486764|T121|1328309|RXNORM|LUFFA OPERCULATA FRUIT EXTRACT|LUFFA OPERCULATA FRUIT EXTRACT
C3256363|T121|1368188|RXNORM|MONOSTEARYL CITRATE|MONOSTEARYL CITRATE
C3256385|T109|1368189|RXNORM|TRIETHYLHEXANOIN|TRIETHYLHEXANOIN
C0016383|T121|4507|RXNORM|FLUSPIRILENE|FLUSPIRILENE
C0016375|T121|4501|RXNORM|FLURAZEPAM|FLURAZEPAM
C0016374|T125|4500|RXNORM|FLURANDRENOLIDE|FLURANDRENOLIDE
C0016377|T121|4502|RXNORM|FLURBIPROFEN|FLURBIPROFEN
C0016377|T121|4502|RXNORM|FLURBIPROFEN|FLURBIPROFEN
C0348029|T121|1368180|RXNORM|TERPINEOL|TERPINEOL
C0611044|T109|1368181|RXNORM|ETHYL STEARATE|ETHYL STEARATE
C0982345|T121|1368182|RXNORM|POLOXAMER 184|POLOXAMER 184
C1509674|T121|1368183|RXNORM|PPG-20 METHYL GLUCOSE ETHER|PPG-20 METHYL GLUCOSE ETHER
C0016384|T121|4508|RXNORM|FLUTAMIDE|FLUTAMIDE
C1530834|T109|1368186|RXNORM|ALPHA-ISOMETHYLIONONE|ALPHA-ISOMETHYLIONONE
C1671133|T109|1368187|RXNORM|TRIDECYL STEARATE|TRIDECYL STEARATE
C0060470|T121|25089|RXNORM|FLOSEQUINAN|FLOSEQUINAN
C0060466|T195|25086|RXNORM|FLORFENICOL|FLORFENICOL
C3504802|T121|1356679|RXNORM|GARCINIA MANGOSTANA FRUIT RIND EXTRACT|GARCINIA MANGOSTANA FRUIT RIND EXTRACT
C3504801|T121|1356678|RXNORM|XYLITAN|XYLITAN
C3535825|T121|1370670|RXNORM|DIHYDROXYCETYL PHOSPHATE|DIHYDROXYCETYL PHOSPHATE
C0724595|T121|221105|RXNORM|HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE|HAEMOPHILUS CAPSULAR OLIGOSACCHARIDE
C3464199|T121|1291441|RXNORM|CHLOROXYLENOL / PETROLATUM|CHLOROXYLENOL / PETROLATUM
C3643352|T109|1422929|RXNORM|PRUNUS DOMESTICA SUBSP. INSITITIA SEED OIL|PRUNUS DOMESTICA SUBSP. INSITITIA SEED OIL
C3643353|T121|1422928|RXNORM|ALOE ARBORESCENS LEAF EXTRACT|ALOE ARBORESCENS LEAF EXTRACT
C0051692|T131|17763|RXNORM|AMITRAZ|AMITRAZ
C0051696|T121|17767|RXNORM|AMLODIPINE|AMLODIPINE
C0178882|T123|62427|RXNORM|URSODEOXYCHOLATE|URSODEOXYCHOLATE
C2725899|T129|971166|RXNORM|WHITE CATFISH ALLERGENIC EXTRACT|AMIURUS CATTUS ALLERGENIC EXTRACT
C1952447|T121|1310709|RXNORM|CETETH-20|CETETH-20
C3256111|T197|1310708|RXNORM|IRON OXIDE BLACK|FERROSOFERRIC OXIDE
C1302002|T121|392464|RXNORM|FUROSEMIDE / POTASSIUM|FUROSEMIDE / POTASSIUM
C1302000|T121|392462|RXNORM|FUROSEMIDE / SPIRONOLACTONE|FUROSEMIDE / SPIRONOLACTONE
C0060087|T120|1310705|RXNORM|FAST GREEN FCF STAIN|FAST GREEN FCF STAIN
C1383453|T130|1310707|RXNORM|D&C RED NO. 28|D&C RED NO. 28
C0728803|T121|1310706|RXNORM|CROSPOVIDONE|CROSPOVIDONE
C3864973|T121|1595630|RXNORM|ACETAMINOPHEN / BROMPHENIRAMINE|ACETAMINOPHEN / BROMPHENIRAMINE
C0600614|T121|155155|RXNORM|POLOXAMER 407|POLOXAMER 407
C0086555|T121|42769|RXNORM|LICORICE|LICORICE
C0082689|T121|41157|RXNORM|GEPEFRINE|GEPEFRINE
C3693112|T121|1482545|RXNORM|PTERIDIUM AQUILINUM WHOLE EXTRACT|PTERIDIUM AQUILINUM WHOLE EXTRACT
C0052945|T121|18752|RXNORM|BAMIFYLLINE|BAMIFYLLINE
C0288792|T121|83947|RXNORM|TAZAROTENE|TAZAROTENE
C0301547|T121|89911|RXNORM|FLUMETHIAZIDE|FLUMETHIAZIDE
C0001040|T127|193|RXNORM|PTPNS1 PROTEIN, HUMAN|ACETYLCARNITINE
C2727904|T129|895279|RXNORM|RAT SKIN EXTRACT|RATTUS NORVEGICUS SKIN EXTRACT
C1874886|T121|689878|RXNORM|COAL TAR / MENTHOL|COAL TAR / MENTHOL
C1874887|T121|689879|RXNORM|COAL TAR / MENTHOL / SALICYLIC ACID|COAL TAR / MENTHOL / SALICYLIC ACID
C0034263|T127|9002|RXNORM|PYRIDOXAL|PYRIDOXAL
C3486606|T196|1427153|RXNORM|GERMANIUM CITRATE LACTATE|GERMANIUM CITRATE LACTATE
C3256838|T109|1427150|RXNORM|GLYCEROL 1,2-DIDOCOSANOATE|GLYCERYL 1,2-DIBEHENATE
C0027679|T121|7315|RXNORM|NEOSTIGMINE|NEOSTIGMINE
C2193976|T121|816701|RXNORM|GUAIFENESIN / NOSCAPINE|GUAIFENESIN / NOSCAPINE
C1509685|T121|1246101|RXNORM|POMEGRANATE FRUIT EXTRACT|POMEGRANATE FRUIT EXTRACT
C0242275|T125|1427158|RXNORM|EPIDERMAL GROWTH FACTOR|EPIDERMAL GROWTH FACTOR
C0070743|T121|33432|RXNORM|PHOLEDRINE|PHOLEDRINE
C0046525|T121|236677|RXNORM|2-PHENYLPHENOL|2-PHENYLPHENOL
C0771976|T121|236674|RXNORM|DIENOGEST / ETHINYL ESTRADIOL|DIENOGEST / ETHINYL ESTRADIOL
C0070742|T121|33431|RXNORM|PHOLCODINE|PHOLCODINE
C0732279|T121|226716|RXNORM|ASPIRIN / DIPYRIDAMOLE|ASPIRIN / DIPYRIDAMOLE
C0772177|T007|236855|RXNORM|LACTOBACILLUS BIFIDUS|LACTOBACILLUS BIFIDUS
C1874165|T121|690997|RXNORM|ALUMINUM HYDROXIDE / ASPIRIN / MAGNESIUM HYDROXIDE|ALUMINUM HYDROXIDE / ASPIRIN / MAGNESIUM HYDROXIDE
C2702374|T129|892638|RXNORM|RYE ALLERGENIC EXTRACT|SECALE CEREALE ALLERGENIC EXTRACT
C0031853|T126|1043631|RXNORM|PHYTASE|PHYTASE
C2928853|T121|1007939|RXNORM|CHOLINE / METHIONINE|CHOLINE / METHIONINE
C2928852|T121|1007938|RXNORM|AMILORIDE / METOLAZONE|AMILORIDE / METOLAZONE
C0036584|T121|9644|RXNORM|SELENOMETHIONINE|SELENOMETHIONINE
C2928847|T121|1007933|RXNORM|HYDROCORTISONE / SODIUM CHLORIDE / UREA|HYDROCORTISONE / SODIUM CHLORIDE / UREA
C2928846|T121|1007932|RXNORM|DIPHENHYDRAMINE / FOMOCAIN / TYROTHRICIN|DIPHENHYDRAMINE / FOMOCAIN / TYROTHRICIN
C2928845|T121|1007931|RXNORM|CITRIC ACID / PEPSIN A|CITRIC ACID / PEPSIN A
C2928844|T121|1007930|RXNORM|BAMETHAN / ESCIN|BAMETHAN / ESCIN
C2928851|T121|1007937|RXNORM|PIROCTONE OLAMINE / SALICYLIC ACID|PIROCTONE OLAMINE / SALICYLIC ACID
C2928850|T121|1007936|RXNORM|HYDROCORTISONE / SULFACETAMIDE|HYDROCORTISONE / SULFACETAMIDE
C2355841|T129|798361|RXNORM|HEPATITIS A VACCINE (INACTIVATED) STRAIN HM175|HEPATITIS A VACCINE (INACTIVATED) STRAIN HM175
C2928848|T121|1007934|RXNORM|ESTRADIOL / HEXACHLOROPHENE|ESTRADIOL / HEXACHLOROPHENE
C0038784|T197|10231|RXNORM|SULFURIC ACID|SULFURIC ACID
C0034283|T121|9010|RXNORM|PYRIMETHAMINE|PYRIMETHAMINE
C0038803|T121|10239|RXNORM|SULPIRIDE|SULPIRIDE
C3818816|T121|1489551|RXNORM|ZANTHOXYLUM PIPERITUM WHOLE EXTRACT|ZANTHOXYLUM PIPERITUM WHOLE EXTRACT
C3818817|T121|1489550|RXNORM|SCHIZONEPETA TENUIFOLIA WHOLE EXTRACT|SCHIZONEPETA TENUIFOLIA WHOLE EXTRACT
C1445185|T129|894934|RXNORM|CHICKEN FEATHER EXTRACT|GALLUS GALLUS FEATHER EXTRACT
C0982109|T130|1305567|RXNORM|D&C YELLOW NO. 10, ALUMINUM LAKE|D&C YELLOW NO. 10, ALUMINUM LAKE
C0054391|T120|1305564|RXNORM|QUINOLINE YELLOW|D&C YELLOW NO. 10
C2729981|T129|892181|RXNORM|BLUEFISH ALLERGENIC EXTRACT|BLUEFISH ALLERGENIC EXTRACT
C3256304|T130|1305560|RXNORM|FD&C RED 40 LAKE|FD&C RED 40 LAKE
C0286651|T121|83367|RXNORM|ATORVASTATIN|ATORVASTATIN
C2033089|T121|822009|RXNORM|PANCREATIN / SIMETHICONE|PANCREATIN / SIMETHICONE
C2740646|T129|899456|RXNORM|MUSTARD SEED ALLERGENIC EXTRACT|MUSTARD SEED ALLERGENIC EXTRACT
C2978230|T121|1088442|RXNORM|6-O-PALMITOYLASCORBIC ACID / ALPHA TOCOPHEROL / COENZYME Q10 / LEVOCARNITINE|6-O-PALMITOYLASCORBIC ACID / ALPHA TOCOPHEROL / COENZYME Q10 / LEVOCARNITINE
C2740643|T129|899452|RXNORM|MUSTARD GREENS ALLERGENIC EXTRACT|MUSTARD GREENS ALLERGENIC EXTRACT
C3848703|T121|1545169|RXNORM|CETEARETH-2|CETEARETH-2
C0301037|T121|89548|RXNORM|DICHLOROBENZENE|DICHLOROBENZENE
C0029997|T121|7781|RXNORM|OXAZEPAM|OXAZEPAM
C0950191|T121|288088|RXNORM|CETRIMIDE|CETRIMIDE
C3859663|T121|1593612|RXNORM|PINUS TAEDA BARK EXTRACT|PINUS TAEDA BARK EXTRACT
C2929698|T121|1008799|RXNORM|ASCORBIC ACID / BIOTIN / FOLIC ACID / MECOBALAMIN / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / ZINC CITRATE|ASCORBIC ACID / BIOTIN / FOLIC ACID / MECOBALAMIN / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / ZINC CITRATE
C2929695|T121|1008796|RXNORM|GIANT RAGWEED POLLEN EXTRACT / WESTERN RAGWEED POLLEN EXTRACT|GIANT RAGWEED POLLEN EXTRACT / WESTERN RAGWEED POLLEN EXTRACT
C2929696|T121|1008797|RXNORM|FEBANTEL / PRAZIQUANTEL / PYRANTEL|FEBANTEL / PRAZIQUANTEL / PYRANTEL
C2929694|T121|1008795|RXNORM|CALCIUM PYRUVATE / DIHYDROXYACETONE|CALCIUM PYRUVATE / DIHYDROXYACETONE
C2929691|T121|1008792|RXNORM|CHOLECALCIFEROL / SOY PROTEIN ISOLATE|CHOLECALCIFEROL / SOY PROTEIN ISOLATE
C2929692|T121|1008793|RXNORM|CHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE / PYRILAMINE|CHLORPHENIRAMINE / HYDROCODONE / PHENYLEPHRINE / PYRILAMINE
C2929690|T121|1008791|RXNORM|ASPIRIN / CAFFEINE / MAGNESIUM CARBONATE / MAGNESIUM SALICYLATE|ASPIRIN / CAFFEINE / MAGNESIUM CARBONATE / MAGNESIUM SALICYLATE
C0003438|T121|1009|RXNORM|ANTITHROMBIN III|ANTITHROMBIN III
C0003420|T121|1001|RXNORM|ANTIPYRINE|ANTIPYRINE
C1165993|T121|350312|RXNORM|ASPERGILLUS NIGER PREPARATION|ASPERGILLUS NIGER PREPARATION
C1165991|T121|350310|RXNORM|MUCOR RACEMOSUS PREPARATION|MUCOR RACEMOSUS PREPARATION
C3818692|T109|1537210|RXNORM|AMORPHOPHALLUS KONJAC ROOT EXTRACT|AMORPHOPHALLUS KONJAC ROOT EXTRACT
C3818691|T121|1537211|RXNORM|CERAMIDE EOP|CERAMIDE EOP
C2370010|T121|827172|RXNORM|DEXCHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE|DEXCHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE
C3859481|T121|1593109|RXNORM|ACETAMINOPHEN / ASPIRIN / DIPHENHYDRAMINE|ACETAMINOPHEN / ASPIRIN / DIPHENHYDRAMINE
C0552314|T121|143980|RXNORM|AMINOBENZOATE|AMINOBENZOATE
C3486726|T121|1354524|RXNORM|CUTTLEFISH PREPARATION|ACANTHOSEPION CUTTLEFISH PREPARATION
C3489050|T121|1354527|RXNORM|PHYSALIA PHYSALIS PREPARATION|PHYSALIA PHYSALIS PREPARATION
C3488474|T121|1354526|RXNORM|PUNICA GRANATUM ROOT BARK EXTRACT|PUNICA GRANATUM ROOT BARK EXTRACT
C2929155|T121|1008248|RXNORM|DEHYDROEPIANDROSTERONE / GINKGO BILOBA EXTRACT|GINKGO BILOBA EXTRACT / PRASTERONE
C2929156|T121|1008249|RXNORM|ALUMINUM SUBACETATE / BORIC ACID|ALUMINUM SUBACETATE / BORIC ACID
C3484402|T121|1338933|RXNORM|SORGHUM EXTRACT|SORGHUM EXTRACT
C3484435|T109|1338934|RXNORM|DROSERA ANGLICA EXTRACT|DROSERA ANGLICA EXTRACT
C2976303|T121|1484911|RXNORM|SOFOSBUVIR|SOFOSBUVIR
C3488954|T121|1338937|RXNORM|PHYSALIS ANGULATA EXTRACT|PHYSALIS ANGULATA EXTRACT
C2929147|T121|1008240|RXNORM|ASCORBIC ACID / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE CHLORIDE / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC SULFATE|ASCORBIC ACID / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE CHLORIDE / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC SULFATE
C2929148|T121|1008241|RXNORM|PREDNISOLONE / ZINC OXIDE|PREDNISOLONE / ZINC OXIDE
C2929149|T121|1008242|RXNORM|BENZALKONIUM / CHLOROXYLENOL / PRAMOXINE|BENZALKONIUM / CHLOROXYLENOL / PRAMOXINE
C2929150|T121|1008243|RXNORM|NYSTATIN / TINIDAZOLE|NYSTATIN / TINIDAZOLE
C2929151|T121|1008244|RXNORM|PREDNISOLONE / PROPYLENE GLYCOL SALICYLATE|PREDNISOLONE / PROPYLENE GLYCOL SALICYLATE
C2929152|T121|1008245|RXNORM|MENTHOL / PREDNISOLONE / THYMOL|MENTHOL / PREDNISOLONE / THYMOL
C2929153|T121|1008246|RXNORM|ASCORBIC ACID / CALCIUM SULFATE / CUPRIC OXIDE / NIACINAMIDE / PYRIDOXINE / VITAMIN B 12|ASCORBIC ACID / CALCIUM SULFATE / CUPRIC OXIDE / NIACINAMIDE / PYRIDOXINE / VITAMIN B 12
C2929154|T121|1008247|RXNORM|NIACINAMIDE / PREDNISOLONE|NIACINAMIDE / PREDNISOLONE
C0032857|T121|8611|RXNORM|POVIDONE-IODINE|POVIDONE-IODINE
C0032857|T121|8611|RXNORM|POVIDONE-IODINE|POVIDONE-IODINE
C0032857|T121|8611|RXNORM|POVIDONE-IODINE|POVIDONE-IODINE
C0032857|T121|8611|RXNORM|POVIDONE-IODINE|POVIDONE-IODINE
C0032857|T121|8611|RXNORM|POVIDONE-IODINE|POVIDONE-IODINE
C0032857|T121|8611|RXNORM|POVIDONE-IODINE|POVIDONE-IODINE
C0032856|T122|8610|RXNORM|POVIDONE|POVIDONE
C0358905|T121|106876|RXNORM|ISONIAZID / RIFAMPIN|ISONIAZID / RIFAMPIN
C3255799|T122|1312709|RXNORM|POLISTIREX|POLISTIREX
C3255662|T126|1312708|RXNORM|DEXTRANASE PENICILLIUM|DEXTRANASE PENICILLIUM
C0076531|T121|38150|RXNORM|THIPHENAMIL|THIPHENAMIL
C2701282|T129|852079|RXNORM|DANDELION POLLEN EXTRACT|TARAXACUM OFFICINALE POLLEN EXTRACT
C0982384|T197|314826|RXNORM|SILICON DIOXIDE, COLLOIDAL|SILICON DIOXIDE, COLLOIDAL
C2701275|T129|852070|RXNORM|LINDEN POLLEN EXTRACT|TILIA CORDATA POLLEN EXTRACT
C0246904|T121|73107|RXNORM|LEVOSIMENDAN|LEVOSIMENDAN
C3494482|T121|1334930|RXNORM|MENTHA PIPERITA EXTRACT|MENTHA PIPERITA EXTRACT
C3255819|T121|1311614|RXNORM|METHYL TRIMETHICONE|METHYL TRIMETHICONE
C2980866|T121|1094082|RXNORM|ARGININE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / THREONINE / TRYPTOPHAN / VALINE|ARGININE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / THREONINE / TRYPTOPHAN / VALINE
C3486011|T121|1311616|RXNORM|ETHYLHEXYL METHOXYCRYLENE|ETHYLHEXYL METHOXYCRYLENE
C3267219|T121|1311617|RXNORM|OCTYLDODECYL MYRISTATE|OCTYLDODECYL MYRISTATE
C2929216|T121|1008309|RXNORM|MINERAL OIL / PETROLATUM / PHENYLEPHRINE / SHARK LIVER OIL|MINERAL OIL / PETROLATUM / PHENYLEPHRINE / SHARK LIVER OIL
C2929215|T121|1008308|RXNORM|ENROFLOXACIN / SILVER SULFADIAZINE|ENROFLOXACIN / SILVER SULFADIAZINE
C3256538|T121|1311612|RXNORM|IPOMOEA PURPUREA TOP EXTRACT|IPOMOEA PURPUREA TOP EXTRACT
C3267652|T121|1311613|RXNORM|GLYCERETH-18|GLYCERETH-18
C2929212|T121|1008305|RXNORM|ASCORBIC ACID / CALCIUM PHOSPHATE DIBASIC / ECHINACEA PURPUREA EXTRACT|ASCORBIC ACID / CALCIUM PHOSPHATE DIBASIC / ECHINACEA PURPUREA EXTRACT
C2929211|T121|1008304|RXNORM|ASCORBIC ACID / BETA CAROTENE / CUPROUS OXIDE / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / BETA CAROTENE / CUPROUS OXIDE / VITAMIN E / ZINC OXIDE
C2929214|T121|1008307|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / CHOLECALCIFEROL / COPPER SULFATE / DOCUSATE / FOLIC ACID / IRON CARBONYL / MAGNESIUM OXIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / ZINC SULFATE|ALPHA TOCOPHEROL / ASCORBIC ACID / CHOLECALCIFEROL / COPPER SULFATE / DOCUSATE / FOLIC ACID / IRON CARBONYL / MAGNESIUM OXIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / ZINC SULFATE
C2929213|T121|1008306|RXNORM|PRAZIQUANTEL / PYRANTEL|PRAZIQUANTEL / PYRANTEL
C2929208|T121|1008301|RXNORM|HARD MAPLE POLLEN EXTRACT / RED MAPLE POLLEN EXTRACT / SILVER MAPLE POLLEN EXTRACT|HARD MAPLE POLLEN EXTRACT / RED MAPLE POLLEN EXTRACT / SILVER MAPLE POLLEN EXTRACT
C2929207|T121|1008300|RXNORM|HYDROFLUMETHIAZIDE / POTASSIUM / RAUWOLFIA PREPARATION|HYDROFLUMETHIAZIDE / POTASSIUM / RAUWOLFIA PREPARATION
C2929210|T121|1008303|RXNORM|CYCLOBENZAPRINE / MAGNESIUM OXIDE|CYCLOBENZAPRINE / MAGNESIUM OXIDE
C2929209|T121|1008302|RXNORM|NAPHAZOLINE / POLYSORBATE 20|NAPHAZOLINE / POLYSORBATE 20
C3255867|T109|1307046|RXNORM|POLYOXYL 20 CETOSTEARYL ETHER|POLYOXYL 20 CETOSTEARYL ETHER
C0443412|T121|1435520|RXNORM|METHYL PROPIONATE|METHYL PROPIONATE
C3255824|T109|1307044|RXNORM|METHYLDIBROMO GLUTARONITRILE|METHYLDIBROMO GLUTARONITRILE
C2348057|T130|1307045|RXNORM|D&C ORANGE NO. 10|D&C ORANGE NO. 10
C3255864|T109|1307042|RXNORM|POLYHYDROXYSTEARIC ACID (2300 MW)|POLYHYDROXYSTEARIC ACID (2300 MW)
C3256497|T168|1307043|RXNORM|APRICOT JUICE EXTRACT|APRICOT JUICE
C3257347|T121|1307040|RXNORM|ASPERGILLUS FLAVUS VAR. ORYZAE PROTEASE|BRINOLASE
C3267318|T121|1307041|RXNORM|PEG-6 COCAMIDE|PEG-6 COCAMIDE
C1695876|T121|631647|RXNORM|CARBETAPENTANE / CARBINOXAMINE / PHENYLEPHRINE|CARBETAPENTANE / CARBINOXAMINE / PHENYLEPHRINE
C3256033|T109|1307048|RXNORM|DIETHYLHEXYL CARBONATE|DIETHYLHEXYL CARBONATE
C3255695|T109|1307049|RXNORM|LITCHI FRUIT EXTRACT|LITCHI FRUIT EXTRACT
C0717827|T121|214621|RXNORM|HYDROCHLOROTHIAZIDE / METOPROLOL|HYDROCHLOROTHIAZIDE / METOPROLOL
C0717826|T121|214620|RXNORM|HYDROCHLOROTHIAZIDE / METHYLDOPA|HYDROCHLOROTHIAZIDE / METHYLDOPA
C0717829|T121|214623|RXNORM|HYDROCHLOROTHIAZIDE / PROPRANOLOL|HYDROCHLOROTHIAZIDE / PROPRANOLOL
C0717828|T121|214622|RXNORM|HYDROCHLOROTHIAZIDE / MOEXIPRIL|HYDROCHLOROTHIAZIDE / MOEXIPRIL
C0717831|T121|214625|RXNORM|HYDROCHLOROTHIAZIDE / TIMOLOL|HYDROCHLOROTHIAZIDE / TIMOLOL
C0717830|T121|214624|RXNORM|HYDROCHLOROTHIAZIDE / RESERPINE|HYDROCHLOROTHIAZIDE / RESERPINE
C3651951|T121|1428987|RXNORM|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS|INFLUENZA A VIRUS VACCINE, A-CALIFORNIA-7-2009 (H1N1)-LIKE VIRUS / INFLUENZA A VIRUS VACCINE, A-VICTORIA-361-2011 (H3N2)-LIKE VIRUS / INFLUENZA B VIRUS VACCINE, B-MASSACHUSETTS-2-2012-LIKE VIRUS
C0717832|T121|214626|RXNORM|HYDROCHLOROTHIAZIDE / VALSARTAN|HYDROCHLOROTHIAZIDE / VALSARTAN
C0717835|T121|214629|RXNORM|HYDROCODONE / PHENYLPROPANOLAMINE|HYDROCODONE / PHENYLPROPANOLAMINE
C0717834|T121|214628|RXNORM|HYDROCODONE / PHENYLEPHRINE|HYDROCODONE / PHENYLEPHRINE
C0600334|T121|155067|RXNORM|SILYBIN|SILIBININ
C2987473|T123|1322428|RXNORM|BOS TAURUS THYMUS PREPARATION|BOVINE THYMUS PREPARATION
C0051771|T130|1370452|RXNORM|AMYL ACETATE|AMYL ACETATE
C3488260|T121|1192621|RXNORM|ASTERIAS RUBENS PREPARATION|ASTERIAS RUBENS PREPARATION
C0059869|T121|24609|RXNORM|ETOFIBRATE|ETOFIBRATE
C1170010|T121|352384|RXNORM|IFOSFAMIDE / MESNA|IFOSFAMIDE / MESNA
C2727176|T129|886637|RXNORM|DOG FLEA ALLERGENIC EXTRACT|CTENOCEPHALIDES CANIS ALLERGENIC EXTRACT
C0165921|T121|60307|RXNORM|ENTACAPONE|ENTACAPONE
C0065166|T121|28876|RXNORM|LONAZOLAC|LONAZOLAC
C0060524|T130|25142|RXNORM|FLUORESCEIN DILAURATE|FLUORESCEIN DILAURATE
C0065162|T121|28872|RXNORM|LOMEFLOXACIN|LOMEFLOXACIN
C0102137|T122|1370451|RXNORM|ALGINATE|ALGINATE
C3818806|T121|1489927|RXNORM|ISOBUTYL STEARATE|ISOBUTYL STEARATE
C0064401|T121|1426451|RXNORM|KOJIC ACID|KOJIC ACID
C3666985|T168|1438112|RXNORM|EUROPEAN ELDERBERRY JUICE PREPARATION|EUROPEAN ELDERBERRY JUICE
C3666984|T121|1438111|RXNORM|CETEARETH 8|CETEARETH 8
C3666983|T109|1438110|RXNORM|QUILLAJA SAPONARIA WOOD EXTRACT|QUILLAJA SAPONARIA WOOD EXTRACT
C3666989|T121|1438116|RXNORM|CUPRESSUS SEMPERVIRENS FRUITING LEAFY TWIG EXTRACT|CUPRESSUS SEMPERVIRENS FRUITING LEAFY TWIG EXTRACT
C3666988|T121|1438115|RXNORM|POLYETHYLENE GLYCOL 2000000|POLYETHYLENE GLYCOL 2000000
C0062941|T121|27100|RXNORM|OMACETAXINE MEPESUCCINATE|OMACETAXINE MEPESUCCINATE
C0054616|T121|20178|RXNORM|OCTANOIC ACID|OCTANOIC ACID
C3855222|T109|1547570|RXNORM|PEACH KERNEL OIL GLYCERETH-8 ESTERS|PEACH KERNEL OIL GLYCERETH-8 ESTERS
C3555464|T109|1420980|RXNORM|SCROPHULARIA NINGPOENSIS ROOT EXTRACT|SCROPHULARIA NINGPOENSIS ROOT EXTRACT
C0208322|T120|1426926|RXNORM|D.C. RED NO. 36|D.C. RED NO. 36
C3864847|T121|1595583|RXNORM|CYNANCHUM STAUNTONII ROOT EXTRACT|CYNANCHUM STAUNTONII ROOT EXTRACT
C0060281|T121|24946|RXNORM|FERROUS SUCCINATE|FERROUS SUCCINATE
C0717386|T121|214199|RXNORM|ALBUTEROL / IPRATROPIUM|ALBUTEROL / IPRATROPIUM
C0301524|T121|89900|RXNORM|SODIUM BITARTRATE|SODIUM BITARTRATE
C1001894|T007|1551569|RXNORM|ALTEROMONAS MACLEODII|ALTEROMONAS MACLEODII
C3864849|T109|1595581|RXNORM|BIS-PHENYLPROPYL DIMETHICONE (15 CST)|BIS-PHENYLPROPYL DIMETHICONE (15 CST)
C0717382|T121|214196|RXNORM|ACRIVASTINE / PSEUDOEPHEDRINE|ACRIVASTINE / PSEUDOEPHEDRINE
C3256625|T109|1426450|RXNORM|MESOPHYLLUM LICHENOIDES EXTRACT|MESOPHYLLUM LICHENOIDES EXTRACT
C2983984|T121|1349278|RXNORM|METENKEFALIN|METENKEFALIN
C2057525|T121|817953|RXNORM|GUAIFENESIN / TERBUTALINE|GUAIFENESIN / TERBUTALINE
C2194168|T121|817778|RXNORM|ASPIRIN / CAFFEINE / QUININE|ASPIRIN / CAFFEINE / QUININE
C3485057|T121|1309682|RXNORM|VERATRUM ALBUM ROOT EXTRACT|VERATRUM ALBUM ROOT EXTRACT
C3486604|T121|1309683|RXNORM|GRINDELIA HIRSUTULA FLOWERING TOP EXTRACT|GRINDELIA CAMPORUM TOP EXTRACT
C0123759|T129|1309680|RXNORM|INTERLEUKIN-12|INTERLEUKIN-12
C3489268|T121|1309681|RXNORM|BAMBUSA VULGARIS LEAF EXTRACT|BAMBUSA VULGARIS LEAF EXTRACT
C3254758|T121|1309686|RXNORM|HELIANTHUS ANNUUS FLOWERING TOP EXTRACT|HELIANTHUS ANNUUS FLOWERING TOP EXTRACT
C3488335|T121|1309684|RXNORM|STROPHANTHUS HISPIDUS SEED EXTRACT|STROPHANTHUS HISPIDUS SEED EXTRACT
C3484422|T121|1309685|RXNORM|RUTA GRAVEOLENS FLOWERING TOP EXTRACT|RUTA GRAVEOLENS FLOWERING TOP EXTRACT
C0140610|T121|55685|RXNORM|RISEDRONIC ACID|RISEDRONIC ACID
C0027368|T125|7244|RXNORM|NANDROLONE|NANDROLONE
C0140594|T121|55681|RXNORM|RIMEXOLONE|RIMEXOLONE
C3267460|T121|1246296|RXNORM|ALUMINUM MAGNESIUM SILICATE / MAGNESIUM HYDROXIDE|ALUMINUM MAGNESIUM SILICATE / MAGNESIUM HYDROXIDE
C2963009|T121|1087558|RXNORM|LUTEIN / OMEGA-3 ACID ETHYL ESTERS (USP) / ZEAXANTHIN|LUTEIN / OMEGA-3 ACID ETHYL ESTERS (USP) / ZEAXANTHIN
C0621433|T109|1370303|RXNORM|SUCROSE DISTEARATE|SUCROSE DISTEARATE
C0301250|T168|1370302|RXNORM|BITTER ALMOND OIL|BITTER ALMOND OIL
C3535636|T121|1370301|RXNORM|RUBIA TINCTORUM WHOLE EXTRACT|RUBIA TINCTORUM WHOLE EXTRACT
C1874365|T121|689515|RXNORM|ASPIRIN / CAFFEINE / HYDROCODONE|ASPIRIN / CAFFEINE / HYDROCODONE
C0041038|T121|10827|RXNORM|TRIMETHADIONE|TRIMETHADIONE
C2939981|T129|1014391|RXNORM|HUMICOLA GRISEA EXTRACT|HUMICOLA GRISEA EXTRACT
C0041031|T121|10825|RXNORM|TRIMEPRAZINE|TRIMEPRAZINE
C1874361|T121|689511|RXNORM|ASPIRIN / CAFFEINE / CODEINE|ASPIRIN / CAFFEINE / CODEINE
C2726180|T129|1014395|RXNORM|MICROSPORUM AUDOUINII ALLERGENIC EXTRACT|MICROSPORUM AUDOUINII ALLERGENIC EXTRACT
C1874362|T121|689512|RXNORM|ASPIRIN / CAFFEINE / DIHYDROCODEINE|ASPIRIN / CAFFEINE / DIHYDROCODEINE
C2726181|T129|1014399|RXNORM|MICROSPORUM CANIS ALLERGENIC EXTRACT|MICROSPORUM CANIS ALLERGENIC EXTRACT
C1874368|T121|689519|RXNORM|ASPIRIN / CAFFEINE / SALICYLAMIDE|ASPIRIN / CAFFEINE / SALICYLAMIDE
C1874367|T121|689518|RXNORM|ASPIRIN / CAFFEINE / PROPOXYPHENE|ASPIRIN / CAFFEINE / PROPOXYPHENE
C0041040|T121|10828|RXNORM|TRIMETHAPHAN|TRIMETHAPHAN
C0041041|T195|10829|RXNORM|TRIMETHOPRIM|TRIMETHOPRIM
C0030078|T121|7816|RXNORM|OXYPHENBUTAZONE|OXYPHENBUTAZONE
C2929777|T121|1008879|RXNORM|CAPSICUM EXTRACT / CASCARA SAGRADA / GINGER EXTRACT / NUX VOMICA EXTRACT|CAPSICUM EXTRACT / CASCARA SAGRADA / GINGER EXTRACT / NUX VOMICA EXTRACT
C2929776|T121|1008878|RXNORM|ANETHOLE TRITHIONE / CHOLINE|ANETHOLE TRITHIONE / CHOLINE
C0030071|T121|7812|RXNORM|OXYMETAZOLINE|OXYMETAZOLINE
C0030071|T121|7812|RXNORM|OXYMETAZOLINE|OXYMETAZOLINE
C0030072|T125|7813|RXNORM|OXYMETHOLONE|OXYMETHOLONE
C2939580|T121|1013625|RXNORM|DROSPIRENONE / ETHINYL ESTRADIOL / LEVOMEFOLIC ACID|DROSPIRENONE / ETHINYL ESTRADIOL / LEVOMEFOLATE
C2929771|T121|1008873|RXNORM|GLYBURIDE / PHENFORMIN|GLYBURIDE / PHENFORMIN
C2929770|T121|1008872|RXNORM|BIFONAZOLE / DIPHENHYDRAMINE|BIFONAZOLE / DIPHENHYDRAMINE
C2929769|T121|1008871|RXNORM|ACETAMINOPHEN / CODEINE / GUAIFENESIN / PHENYLEPHRINE|ACETAMINOPHEN / CODEINE / GUAIFENESIN / PHENYLEPHRINE
C0078794|T197|39954|RXNORM|ZINC SULFATE|ZINC SULFATE
C2929775|T121|1008877|RXNORM|ASPIRIN / CHLORPHENIRAMINE / PSEUDOEPHEDRINE|ASPIRIN / CHLORPHENIRAMINE / PSEUDOEPHEDRINE
C2929774|T121|1008876|RXNORM|KELP PREPARATION / VITAMIN B6|KELP PREPARATION / VITAMIN B6
C2929773|T121|1008875|RXNORM|CALCIUM PHOSPHATE / CHROMIUM PICOLINATE|CALCIUM PHOSPHATE / CHROMIUM PICOLINATE
C2929772|T121|1008874|RXNORM|SOY PROTEIN ISOLATE / SOYBEAN PREPARATION|SOY PROTEIN ISOLATE / SOYBEAN PREPARATION
C0086268|T121|42682|RXNORM|ETIDRONATE|ETIDRONATE
C0055738|T121|21116|RXNORM|EUCALYPTOL|CINEOLE
C3475023|T121|1302471|RXNORM|LACTOBACILLUS REUTERI / LACTOBACILLUS RHAMNOSUS GG|LACTOBACILLUS REUTERI / LACTOBACILLUS RHAMNOSUS GG
C1099414|T121|321952|RXNORM|PIMECROLIMUS|PIMECROLIMUS
C0016369|T125|4497|RXNORM|FLUPREDNISOLONE|FLUPREDNISOLONE
C0771722|T121|236449|RXNORM|PROPYLENE GLYCOL SALICYLATE|PROPYLENE GLYCOL SALICYLATE
C3281747|T121|1249671|RXNORM|BIFIDOBACTERIUM LACTIS / LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS CASEI RHAMNOSUS|BIFIDOBACTERIUM LACTIS / LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS CASEI RHAMNOSUS
C2001867|T121|1433693|RXNORM|FERRIC CARBOXYMALTOSE|FERRIC CARBOXYMALTOSE
C3540668|T121|1424266|RXNORM|LOBELIA CARDINALIS EXTRACT|CARDINAL FLOWER EXTRACT
C3245436|T121|1191399|RXNORM|FLUOCINOLONE / ZINC PYRITHIONE|FLUOCINOLONE / ZINC PYRITHIONE
C0001134|T197|236|RXNORM|BIOFLAVONOID, LEMON|ACIDULATED PHOSPHATE FLUORIDE
C2701166|T129|851926|RXNORM|CARELESS WEED POLLEN EXTRACT|AMARANTHUS PALMERI POLLEN EXTRACT
C3818764|T109|1492385|RXNORM|COLCHICUM AUTUMNALE FLOWER EXTRACT|COLCHICUM AUTUMNALE FLOWER EXTRACT
C3818765|T109|1492383|RXNORM|SALIX PURPUREA BARK EXTRACT|SALIX PURPUREA BARK EXTRACT
C0016365|T121|4493|RXNORM|FLUOXETINE|FLUOXETINE
C0141729|T121|56084|RXNORM|SCHIZANDRA PREPARATION|SCHIZANDRA PREPARATION
C0016351|T121|4491|RXNORM|FLUOROMETHOLONE|FLUOROMETHOLONE
C0872906|T121|259274|RXNORM|MILK THISTLE SEED EXTRACT|MILK THISTLE SEED EXTRACT
C1445656|T121|466424|RXNORM|ASPIRIN / CAFFEINE / CINNAMEDRINE|ASPIRIN / CAFFEINE / CINNAMEDRINE
C1445658|T121|466426|RXNORM|BENZOCAINE / MENTHOL|BENZOCAINE / MENTHOL
C1445658|T121|466426|RXNORM|BENZOCAINE / MENTHOL|BENZOCAINE / MENTHOL
C1445659|T121|466427|RXNORM|BENZOCAINE / RESORCINOL|BENZOCAINE / RESORCINOL
C1445655|T121|466423|RXNORM|ANTIPYRINE / BENZOCAINE|ANTIPYRINE / BENZOCAINE
C0055915|T195|21264|RXNORM|CLOFOCTOL|CLOFOCTOL
C2722017|T129|1370773|RXNORM|BEAN EXTRACT|BEAN EXTRACT
C0291216|T130|84990|RXNORM|GADOBUTROL|GADOBUTROL
C1445660|T121|466428|RXNORM|ANTIPYRINE / BENZOCAINE / PHENYLEPHRINE|ANTIPYRINE / BENZOCAINE / PHENYLEPHRINE
C1445661|T121|466429|RXNORM|CAMPHOR / MENTHOL / PHENOL|CAMPHOR / MENTHOL / PHENOL
C2948830|T121|1370774|RXNORM|ASIAN GINSENG EXTRACT|ASIAN GINSENG EXTRACT
C2723553|T129|905070|RXNORM|ACREMONIUM STRICTUM ALLERGENIC EXTRACT|SAROCLADIUM STRICTUM ALLERGENIC EXTRACT
C2315887|T121|754763|RXNORM|FOSAPREPITANT DIMEGLUMINE|FOSAPREPITANT DIMEGLUMINE
C0006466|T121|1829|RXNORM|BUTACAINE|BUTACAINE
C0006463|T131|1828|RXNORM|BUSULFAN|BUSULFAN
C0006456|T121|1825|RXNORM|BUSERELIN|BUSERELIN
C0006462|T121|1827|RXNORM|BUSPIRONE|BUSPIRONE
C2344068|T129|797631|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP C CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE|NEISSERIA MENINGITIDIS SEROGROUP C CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE
C0008296|T121|2410|RXNORM|CHLORZOXAZONE|CHLORZOXAZONE
C2722036|T129|891727|RXNORM|COFFEE BEAN ALLERGENIC EXTRACT|COFFEE BEAN ALLERGENIC EXTRACT
C0008318|T127|2418|RXNORM|CHOLECALCIFEROL|CHOLECALCIFEROL
C0907402|T125|274783|RXNORM|INSULIN GLARGINE|INSULIN GLARGINE
C0117480|T121|49991|RXNORM|DROPERIDOL / FENTANYL|DROPERIDOL / FENTANYL
C0025624|T121|6821|RXNORM|METHANTHELINE|METHANTHELINE
C2701120|T129|851866|RXNORM|SILVER MAPLE POLLEN EXTRACT|ACER SACCHARINUM POLLEN EXTRACT
C3538508|T121|1372934|RXNORM|SODIUM LAURETH-13 CARBOXYLATE|SODIUM LAURETH-13 CARBOXYLATE
C0937775|T121|283682|RXNORM|PULSATILLA PRATENSIS EXTRACT|ANEMONE PRATENSIS EXTRACT
C1875404|T121|690702|RXNORM|ISOPROPYL ALCOHOL / SALICYLIC ACID / SODIUM THIOSULFATE|ISOPROPYL ALCOHOL / SALICYLIC ACID / SODIUM THIOSULFATE
C1875402|T121|690700|RXNORM|ISOPROPAMIDE / PROCHLORPERAZINE|ISOPROPAMIDE / PROCHLORPERAZINE
C0011796|T121|3275|RXNORM|DEXTRAN 75|DEXTRAN 75
C0011793|T121|3272|RXNORM|DEXTRAN 40|DEXTRAN 40
C0006720|T197|1925|RXNORM|CALCIUM SULFATE|CALCIUM SULFATE
C2928400|T121|1007478|RXNORM|BENZALKONIUM / LAURETH-9 / MEPIVACAINE|BENZALKONIUM / MEPIVACAINE / POLIDOCANOL
C0025629|T121|6825|RXNORM|METHARBITAL|METHARBITAL
C1874223|T121|692960|RXNORM|AMPHOTERICIN B / TETRACYCLINE|AMPHOTERICIN B / TETRACYCLINE
C1874719|T121|692969|RXNORM|CARBON DIOXIDE / NITROGEN|CARBON DIOXIDE / NITROGEN
C1532673|T121|484348|RXNORM|OMEGA-3 ACID ETHYL ESTERS (USP)|OMEGA-3 ACID ETHYL ESTERS (USP)
C2722034|T129|891721|RXNORM|COCOA BEAN ALLERGENIC EXTRACT|THEOBROMA CACAO ALLERGENIC EXTRACT
C0772172|T121|236850|RXNORM|ICTASOL|ICTASOL
C0075007|T121|36908|RXNORM|SPIRAPRIL|SPIRAPRIL
C0304631|T121|91326|RXNORM|HOMOSALATE|HOMOSALATE
C0053233|T121|18997|RXNORM|BENZOPHENONE|BENZOPHENONE
C0053230|T121|18994|RXNORM|BENZONIDAZOLE|BENZONIDAZOLE
C2929403|T121|1008499|RXNORM|CYSTEINE / VITAMIN B6|CYSTEINE / VITAMIN B6
C0053229|T121|18993|RXNORM|BENZONATATE|BENZONATATE
C0302961|T197|1311379|RXNORM|SULFUR IODIDE|SULFUR IODIDE
C0043367|T130|1311378|RXNORM|XYLENE|XYLENE
C0360518|T125|108074|RXNORM|CLOBETASONE|CLOBETASONE
C2929398|T121|1008494|RXNORM|BENZOATE / GUAIACOLSULFONATE|BENZOATE / GUAIACOLSULFONATE
C2929401|T121|1008497|RXNORM|DOCUSATE / FERROUS FUMARATE / FOLIC ACID|DOCUSATE / FERROUS FUMARATE / FOLIC ACID
C2348735|T121|1311374|RXNORM|GARDENIA JASMINOIDES FRUIT EXTRACT|GARDENIA JASMINOIDES FRUIT EXTRACT
C2929395|T121|1008491|RXNORM|ISOPROPYL ALCOHOL / METHYL SALICYLATE|ISOPROPYL ALCOHOL / METHYL SALICYLATE
C2929397|T121|1008493|RXNORM|BENZOATE / CODEINE|BENZOATE / CODEINE
C2929396|T121|1008492|RXNORM|CAFFEINE / PHENIRAMINE / PHENYLEPHRINE / SALICYLIC ACID|CAFFEINE / PHENIRAMINE / PHENYLEPHRINE / SALICYLIC ACID
C3527684|T121|1360726|RXNORM|PHENYLEPHRINE / THONZYLAMINE|PHENYLEPHRINE / THONZYLAMINE
C0068006|T121|1494066|RXNORM|MILTEFOSINE|MILTEFOSINE
C3273754|T121|1539753|RXNORM|EFINACONAZOLE|EFINACONAZOLE
C0020264|T121|5489|RXNORM|HYDROCODONE|HYDROCODONE
C0020261|T121|5487|RXNORM|HYDROCHLOROTHIAZIDE|HYDROCHLOROTHIAZIDE
C0020259|T197|5486|RXNORM|HYDROCHLORIC ACID|HYDROCHLORIC ACID
C0020259|T197|5486|RXNORM|HYDROCHLORIC ACID|HYDROCHLORIC ACID
C3255954|T121|1307828|RXNORM|MANGIFERA INDICA SEED BUTTER EXTRACT|MANGIFERA INDICA SEED BUTTER EXTRACT
C3256072|T121|1307829|RXNORM|PEG-4 RAPESEEDAMIDE|PEG-4 RAPESEEDAMIDE
C3486390|T121|1358956|RXNORM|ANACARDIUM OCCIDENTALE FRUIT EXTRACT|ANACARDIUM OCCIDENTALE FRUIT EXTRACT
C2697922|T168|1358957|RXNORM|LIME JUICE|LIME JUICE
C0026370|T168|1307820|RXNORM|MOLASSES|MOLASSES
C3256435|T109|1307822|RXNORM|PLUKENETIA VOLUBILIS SEED OIL|PLUKENETIA VOLUBILIS SEED OIL
C0064688|T121|1596928|RXNORM|DODECYL GALLATE|DODECYL GALLATE
C3256804|T121|1307824|RXNORM|SENNA ALATA LEAF EXTRACT|SENNA ALATA LEAF EXTRACT
C3486530|T109|1307825|RXNORM|OLEA EUROPAEA FRUIT VOLATILE OIL|OLEA EUROPAEA FRUIT VOLATILE OIL
C3256667|T121|1307826|RXNORM|CAMELLIA JAPONICA LEAF EXTRACT|CAMELLIA JAPONICA LEAF EXTRACT
C3256139|T121|1307827|RXNORM|COIX LACRYMA-JOBI VAR. MA-YUEN SEED EXTRACT|COIX LACRYMA-JOBI VAR. MA-YUEN SEED EXTRACT
C0982353|T121|314797|RXNORM|POTASSIUM LACTATE|POTASSIUM LACTATE
C0724624|T121|1310578|RXNORM|MEDIUM CHAIN TRIGLYCERIDES|MEDIUM CHAIN TRIGLYCERIDES
C0089147|T109|1310579|RXNORM|1-BUTANOL|1-BUTANOL
C0790024|T168|1310576|RXNORM|CORN SYRUP|CORN SYRUP
C0079594|T121|40138|RXNORM|ILOPROST|ILOPROST
C3484462|T121|1310574|RXNORM|CROSCARMELLOSE|CROSCARMELLOSE
C2986958|T130|1310575|RXNORM|FD&C RED NO. 4|FD&C RED NO. 4
C0060240|T197|1310572|RXNORM|FERRIC OXIDE|FERRIC OXIDE
C3255782|T109|1310570|RXNORM|LAURETH-3|LAURETH-3
C1366066|T121|1310571|RXNORM|SHEA BUTTER|SHEA BUTTER
C2724202|T129|892372|RXNORM|CELERY ALLERGENIC EXTRACT|APIUM GRAVEOLENS ALLERGENIC EXTRACT
C0004595|T007|1311119|RXNORM|BACILLUS SUBTILIS|BACILLUS SUBTILIS
C0060937|T196|1311118|RXNORM|GADOLINIUM OXIDE|GADOLINIUM OXIDE
C0004590|T007|1311112|RXNORM|BACILLUS CEREUS|BACILLUS CEREUS
C0065987|T197|1311110|RXNORM|MERCURIC CYANIDE|MERCURIC CYANIDE
C2604206|T121|840781|RXNORM|DROSPIRENONE / ETHINYL ESTRADIOL|DROSPIRENONE / ETHINYL ESTRADIOL
C3497902|T196|1311116|RXNORM|EUROPIUM OXIDE|EUROPIUM OXIDE
C0301318|T121|89736|RXNORM|PHTHALYLSULFACETAMIDE|PHTHALYLSULFACETAMIDE
C0534702|T197|1311114|RXNORM|LANTHANUM OXIDE|LANTHANUM OXIDE
C0000392|T123|61|RXNORM|BETA-ALANINE|BETA-ALANINE
C0008377|T123|2438|RXNORM|CHOLESTEROL|CHOLESTEROL
C0163518|T121|59247|RXNORM|DIPERODON|DIPERODON
C0304097|T168|1309373|RXNORM|CARAWAY OIL|CARAWAY OIL
C3700994|T121|1485741|RXNORM|CAMPHOR / CAPSAICIN|CAMPHOR / CAPSAICIN
C2929713|T121|1008814|RXNORM|DEHYDROCHOLATE / HOMATROPINE / PHENOBARBITAL|DEHYDROCHOLATE / HOMATROPINE / PHENOBARBITAL
C3485687|T121|1304558|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / BIOTIN / CHOLECALCIFEROL / DEXPANTHENOL / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN K 1|ALPHA TOCOPHEROL / ASCORBIC ACID / BIOTIN / CHOLECALCIFEROL / DEXPANTHENOL / FOLIC ACID / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN K 1
C3488955|T109|1309309|RXNORM|PINUS STROBUS BARK EXTRACT|PINUS STROBUS BARK EXTRACT
C1121849|T121|1098413|RXNORM|VANDETANIB|VANDETANIB
C3497397|T121|1309301|RXNORM|PYRIMETHAMINE / SULFADIAZINE|PYRIMETHAMINE / SULFADIAZINE
C0006882|T121|1982|RXNORM|CANRENONE|CANRENONE
C0065850|T121|29426|RXNORM|MECYSTEINE|MECYSTEINE
C0304145|T109|1309375|RXNORM|OIL OF NIAOULI|OIL OF NIAOULI
C0065844|T127|29421|RXNORM|MECOBALAMIN|METHYLCOBALAMIN
C0002475|T195|632|RXNORM|MITOMYCIN|MITOMYCIN
C0002475|T195|632|RXNORM|MITOMYCIN|MITOMYCIN
C0028923|T195|7629|RXNORM|LACTALBUMINS, HYDROLYZATES|OLEANDOMYCIN
C1950688|T121|705258|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / DOXYLAMINE|ACETAMINOPHEN / DEXTROMETHORPHAN / DOXYLAMINE
C1950688|T121|705258|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / DOXYLAMINE|ACETAMINOPHEN / DEXTROMETHORPHAN / DOXYLAMINE
C2075862|T121|812444|RXNORM|BENDROFLUMETHIAZIDE / CLONIDINE|BENDROFLUMETHIAZIDE / CLONIDINE
C0004234|T121|1218|RXNORM|ATRACURIUM|ATRACURIUM
C0877860|T121|262307|RXNORM|FELBINAC|FELBINAC
C1260235|T121||RXNORM|ETHINYL ESTRADIOL / NORETHINDRONE
C1260235|T121||RXNORM|ETHINYL ESTRADIOL / NORETHINDRONE
C2928140|T121|1007218|RXNORM|OUABAIN / PHENOBARBITAL|OUABAIN / PHENOBARBITAL
C2928141|T121|1007219|RXNORM|BLACK CURRANT PREPARATION / SODIUM CITRATE|BLACK CURRANT PREPARATION / SODIUM CITRATE
C2928138|T121|1007216|RXNORM|GLYCOL SALICYLATE / MENTHOL|GLYCOL SALICYLATE / MENTHOL
C2928139|T121|1007217|RXNORM|HOMATROPINE / SCOPOLAMINE|HOMATROPINE / SCOPOLAMINE
C2928136|T121|1007214|RXNORM|NIACINAMIDE / POTASSIUM|NIACINAMIDE / POTASSIUM
C2928137|T121|1007215|RXNORM|SHEEP SORREL POLLEN EXTRACT / YELLOW DOCK POLLEN EXTRACT|SHEEP SORREL POLLEN EXTRACT / YELLOW DOCK POLLEN EXTRACT
C2928134|T121|1007212|RXNORM|BENTONITE / SULFUR / TRICLOSAN|BENTONITE / SULFUR / TRICLOSAN
C2928135|T121|1007213|RXNORM|LACTOBACILLUS ACIDOPHILUS / PLANTAGO SEED|LACTOBACILLUS ACIDOPHILUS / PLANTAGO SEED
C2928132|T121|1007210|RXNORM|DIPYRONE / HOMATROPINE / PAPAVERINE|DIPYRONE / HOMATROPINE / PAPAVERINE
C2928133|T121|1007211|RXNORM|POLYOXYETHYLENE ETHER / SULFUR|POLYOXYETHYLENE ETHER / SULFUR
C3818811|T109|1489764|RXNORM|PEG-3 DISTEARATE|PEG-3 DISTEARATE
C3818810|T109|1489765|RXNORM|TERT-BUTYL METHACRYLATE|TERT-BUTYL METHACRYLATE
C3818814|T109|1489760|RXNORM|PAEONIA OFFICINALIS WHOLE EXTRACT|PAEONIA OFFICINALIS WHOLE EXTRACT
C3818813|T109|1489761|RXNORM|PEG-45 PALM KERNEL GLYCERIDES|PEG-45 PALM KERNEL GLYCERIDES
C1136262|T197|1489762|RXNORM|TECHNETIUM TC 99M PERTECHNETATE|TECHNETIUM TC 99M PERTECHNETATE
C3818812|T109|1489763|RXNORM|PADANG CASSIA OIL|PADANG CASSIA OIL
C3528229|T109|1362142|RXNORM|PROLINAMIDOETHYL IMIDAZOLE|PROLINAMIDOETHYL IMIDAZOLE
C0066101|T121|29648|RXNORM|METHDILAZINE|METHDILAZINE
C3528228|T109|1362141|RXNORM|PICEA MARIANA LEAF OIL|PICEA MARIANA LEAF OIL
C3528232|T109|1362146|RXNORM|LINALOOL, ()-|LINALOOL, ()-
C3464053|T121|1362147|RXNORM|HYDROXYETHYL CELLULOSE (100 MPA.S AT 2%)|HYDROXYETHYL CELLULOSE (100 MPA.S AT 2%)
C3528230|T109|1362144|RXNORM|C12-15 PARETH-9|C12-15 PARETH-9
C3528231|T109|1362145|RXNORM|PEG-120 STEARATE|PEG-120 STEARATE
C0072735|T121|35100|RXNORM|PYRITHIONE|PYRITHIONE
C0347993|T121|1232405|RXNORM|PYRETHRUM EXTRACT|PYRETHRUM
C3486633|T121|1337633|RXNORM|EUPHORBIA LATHYRIS EXTRACT|EUPHORBIA LATHYRIS EXTRACT
C0082608|T121|41127|RXNORM|FLUVASTATIN|FLUVASTATIN
C3488905|T121|1337637|RXNORM|HABANERO EXTRACT|HABANERO EXTRACT
C3486762|T121|1337634|RXNORM|LOMATIUM DISSECTUM ROOT EXTRACT|LOMATIUM DISSECTUM ROOT EXTRACT
C1134659|T129|1232150|RXNORM|AFLIBERCEPT|AFLIBERCEPT
C1134659|T129|1232150|RXNORM|AFLIBERCEPT|AFLIBERCEPT
C3249436|T121|1232409|RXNORM|PIPERONYL BUTOXIDE / PYRETHRUM EXTRACT|PIPERONYL BUTOXIDE / PYRETHRUM EXTRACT
C3539881|T129|1421648|RXNORM|GAMMA-INTERFERON|GAMMA-INTERFERON
C3256717|T109|1368192|RXNORM|PPG-14 BUTYL ETHER|PPG-14 BUTYL ETHER
C0677517|T196|196213|RXNORM|FLUORIDE ION|FLUORIDE ION
C0053782|T197|19469|RXNORM|BISMUTH CARBONATE|BISMUTH CARBONATE
C2918456|T121|995600|RXNORM|ROUGH COCKLEBUR POLLEN EXTRACT|ROUGH COCKLEBUR POLLEN EXTRACT
C3643660|T121|1421642|RXNORM|PHENOL / SCARLET RED|PHENOL / SCARLET RED
C3256541|T109|1368191|RXNORM|ISOCETYL ALCOHOL|ISOCETYL ALCOHOL
C0004749|T196|1311067|RXNORM|BARIUM|BARIUM
C3256455|T109|1368190|RXNORM|TRISILOXANE|TRISILOXANE
C0725101|T197|221456|RXNORM|ALUM, POTASSIUM|ALUM, POTASSIUM
C0040602|T123|1368197|RXNORM|TRAGACANTH|TRAGACANTH
C1832027|T129|712566|RXNORM|OFATUMUMAB|OFATUMUMAB
C0074002|T123|1311309|RXNORM|SALSOLINOL|SALSOLINOL
C2725885|T129|882469|RXNORM|PACIFIC HALIBUT ALLERGENIC EXTRACT|HIPPOGLOSSUS STENOLEPIS ALLERGENIC EXTRACT
C0717454|T121|594040|RXNORM|ATROPINE / DIPHENOXYLATE|ATROPINE / DIPHENOXYLATE
C3651792|T122|1428041|RXNORM|POLYQUATERNIUM-39 (22.5-51-26.5 ACRYLIC ACID-ACRYLAMIDE-DADMAC; 1600000 MW)|POLYQUATERNIUM-39 (22.5-51-26.5 ACRYLIC ACID-ACRYLAMIDE-DADMAC; 1600000 MW)
C3651791|T121|1428042|RXNORM|PANAX QUINQUEFOLIUS WHOLE EXTRACT|PANAX QUINQUEFOLIUS WHOLE EXTRACT
C3539111|T121|1428043|RXNORM|HYACINTHOIDES NON-SCRIPTA EXTRACT|HYACINTHOIDES NON-SCRIPTA EXTRACT
C1445424|T129|466195|RXNORM|BOTRYTIS CINEREA EXTRACT|BOTRYTIS CINEREA EXTRACT
C0023115|T122|1314891|RXNORM|LATEX|LATEX
C2073925|T121|813792|RXNORM|CHLORZOXAZONE / PIROXICAM|CHLORZOXAZONE / PIROXICAM
C2194203|T121|813791|RXNORM|ASCORBIC ACID / SODIUM FLUORIDE|ASCORBIC ACID / SODIUM FLUORIDE
C0995001|T121|318224|RXNORM|FLAXSEED EXTRACT|FLAXSEED EXTRACT
C0042971|T123|11274|RXNORM|VON WILLEBRAND FACTOR|VON WILLEBRAND FACTOR
C2725895|T129|882482|RXNORM|TROUT ALLERGENIC EXTRACT|TROUT ALLERGENIC EXTRACT
C0015091|T121|4158|RXNORM|ETHYLENEDIAMINE|ETHYLENEDIAMINE
C0168388|T121|60842|RXNORM|REBOXETINE|REBOXETINE
C0982443|T121|314881|RXNORM|UNDECYLENATE|UNDECYLENATE
C2723235|T121||RXNORM|MORPHINE / NALTREXONE
C3856128|T109|1549633|RXNORM|ABIES ALBA LEAF OIL|ABIES ALBA LEAF OIL
C3856127|T121|1549632|RXNORM|HYDROXYETHYL CETYLDIMONIUM PHOSPHATE|HYDROXYETHYL CETYLDIMONIUM PHOSPHATE
C2980896|T121|1094140|RXNORM|MELATONIN / TRYPTOPHAN|MELATONIN / TRYPTOPHAN
C1874989|T121|690492|RXNORM|DEXTROMETHORPHAN / TERPIN HYDRATE|DEXTROMETHORPHAN / TERPIN HYDRATE
C0875947|T121|261435|RXNORM|SODIUM FERRIC GLUCONATE COMPLEX|SODIUM FERRIC GLUCONATE COMPLEX
C0875944|T121|261432|RXNORM|PHENYLEPHRINE / PYRILAMINE|PHENYLEPHRINE / PYRILAMINE
C0875944|T121|261432|RXNORM|PHENYLEPHRINE / PYRILAMINE|PHENYLEPHRINE / PYRILAMINE
C0875944|T121|261432|RXNORM|PHENYLEPHRINE / PYRILAMINE|PHENYLEPHRINE / PYRILAMINE
C3818800|T121|1490684|RXNORM|LINDERA AGGREGATA WHOLE EXTRACT|LINDERA AGGREGATA WHOLE EXTRACT
C0285260|T121|82910|RXNORM|PIKETOPROFEN|PIKETOPROFEN
C0717579|T121|214382|RXNORM|CHLOROTHIAZIDE / METHYLDOPA|CHLOROTHIAZIDE / METHYLDOPA
C0717580|T121|214383|RXNORM|CHLOROTHIAZIDE / RESERPINE|CHLOROTHIAZIDE / RESERPINE
C3256381|T121|1313267|RXNORM|TRIDECETH-12|TRIDECETH-12
C3256559|T109|1313266|RXNORM|POLYETHYLENE GLYCOL 500|POLYETHYLENE GLYCOL 500
C3465014|T109|1313265|RXNORM|ETHYLHEXYL ETHYLHEXANOATE|ETHYLHEXYL ETHYLHEXANOATE
C3265832|T121|1313264|RXNORM|DIMETHICONE PEG-8 LAURATE|DIMETHICONE PEG-8 LAURATE
C0257715|T121|77674|RXNORM|OCTOCRYLENE|OCTOCRYLENE
C0048468|T121|1313261|RXNORM|4-METHYL ANISOLE|4-METHYL ANISOLE
C2728185|T129|1011027|RXNORM|PARSNIP ALLERGENIC EXTRACT|PARSNIP ALLERGENIC EXTRACT
C3818803|T121|1490681|RXNORM|ANGELICA PUBESCENS WHOLE EXTRACT|ANGELICA PUBESCENS WHOLE EXTRACT
C1113707|T121|324072|RXNORM|DIMETHICONE|DIMETICONE
C1113707|T121|324072|RXNORM|DIMETHICONE|DIMETICONE
C2940167|T129|1014707|RXNORM|REDWOOD POLLEN EXTRACT|SEQUOIA SEMPERVIRENS POLLEN EXTRACT
C3267310|T121|1313269|RXNORM|CITRONELLOL ACETATE, (S)-|CITRONELLOL ACETATE, (S)-
C2825626|T121|1313268|RXNORM|QUADROSILAN|QUADROSILAN
C1578246|T121|477468|RXNORM|MORPHINE LIPOSOMAL|MORPHINE LIPOSOMAL
C1530889|T121|1364468|RXNORM|TEDUGLUTIDE|TEDUGLUTIDE
C3818801|T121|1490683|RXNORM|CASTORYL MALEATE|CASTORYL MALEATE
C0982090|T121|1364462|RXNORM|COCOAMPHODIACETATE|COCOAMPHODIACETATE
C0018483|T007|1364467|RXNORM|HAEMOPHILUS INFLUENZAE|HAEMOPHILUS INFLUENZAE
C0069761|T121|32634|RXNORM|OXFENDAZOLE|OXFENDAZOLE
C0069760|T121|32633|RXNORM|OXETORONE|OXETORONE
C0052927|T121|1592893|RXNORM|BAICALEIN|BAICALEIN
C0068992|T125|31994|RXNORM|NORGESTIMATE|NORGESTIMATE
C0033405|T121|8745|RXNORM|PROMETHAZINE|PROMETHAZINE
C0069766|T121|32639|RXNORM|OXILOFRINE|OXILOFRINE
C0069765|T121|32638|RXNORM|OXICONAZOLE|OXICONAZOLE
C0012498|T121|3489|RXNORM|DIOSMIN|DIOSMIN
C0033401|T125|8744|RXNORM|PROMEGESTONE|PROMEGESTONE
C0003382|T121|981|RXNORM|ANTIMONY POTASSIUM TARTRATE|ANTIMONY POTASSIUM TARTRATE
C3818796|T121|1490689|RXNORM|SCROPHULARIA NINGPOENSIS WHOLE EXTRACT|SCROPHULARIA NINGPOENSIS WHOLE EXTRACT
C3696423|T121|1483193|RXNORM|BENZALKONIUM / BENZOCAINE / MENTHOL|BENZALKONIUM / BENZOCAINE / MENTHOL
C0031617|T123|8214|RXNORM|LECITHIN|PHOSPHATIDYL CHOLINE
C0031621|T123|8217|RXNORM|PHOSPHATIDYLINOSITOLS|PHOSPHATIDYLINOSITOLS
C3257044|T121|1241470|RXNORM|CARBOXYMETHYLCELLULOSE / GLYCERIN / POLYSORBATE 80|CARBOXYMETHYLCELLULOSE / GLYCERIN / POLYSORBATE 80
C0048318|T121|15080|RXNORM|MEQUINOL|MEQUINOL
C3256775|T109|1426558|RXNORM|LAMINARIA JAPONICA EXTRACT|LAMINARIA JAPONICA EXTRACT
C3256776|T121|1426559|RXNORM|LAMINARIA OCHROLEUCA EXTRACT|LAMINARIA OCHROLEUCA EXTRACT
C0037874|T123|1483263|RXNORM|SPERMINE|SPERMINE
C0037871|T123|1483262|RXNORM|SPERMIDINE|SPERMIDINE
C3665462|T122|1483267|RXNORM|RAW SUGAR|RAW SUGAR
C1188555|T007|1321355|RXNORM|ARTHROSPIRA PLATENSIS|ARTHROSPIRA PLATENSIS
C3667079|T109|1483230|RXNORM|HYDROGENATED JOJOBA OIL-JOJOBA OIL, RANDOMIZED (IODINE VALUE 57-61)|HYDROGENATED JOJOBA OIL-JOJOBA OIL, RANDOMIZED (IODINE VALUE 57-61)
C0872912|T123|579598|RXNORM|SOYBEAN LECITHIN|SOYBEAN LECITHIN
C3256335|T109|1307565|RXNORM|AMMONIUM LAURETH-2 SULFATE|AMMONIUM LAURETH-2 SULFATE
C3255667|T121|1307564|RXNORM|EPILOBIUM ANGUSTIFOLIUM FLOWERING TOP EXTRACT|EPILOBIUM ANGUSTIFOLIUM FLOWERING TOP EXTRACT
C0060246|T197|24913|RXNORM|FERRIC SULFATE|FERRIC SULFATE
C3256738|T121|1307566|RXNORM|URTICA URENS LEAF EXTRACT|URTICA URENS LEAF EXTRACT
C3256208|T121|1307561|RXNORM|CUCUMARIA SEA CUCUMBER EXTRACT|CUCUMARIA SEA CUCUMBER EXTRACT
C3154683|T121|1102200|RXNORM|ASCORBIC ACID / BIOTIN / CALCIUM CARBONATE / FOLIC ACID / NIACIN / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / SUCCINIC ACID / THIAMINE / VITAMIN B 12|ASCORBIC ACID / BIOTIN / CALCIUM CARBONATE / FOLIC ACID / NIACIN / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / SUCCINIC ACID / THIAMINE / VITAMIN B 12
C3256210|T168|1307563|RXNORM|CUCUMBER JUICE EXTRACT|CUCUMBER JUICE
C3256136|T109|1307562|RXNORM|COCONUT ACID|COCONUT ACID
C2825375|T130|1307569|RXNORM|BEHENETH-10|BEHENETH-10
C3256257|T121|1307568|RXNORM|ROSA DAMASCENA FLOWER EXTRACT|ROSA DAMASCENA FLOWER EXTRACT
C3668710|T121|1441298|RXNORM|AMANITA PANTHERINA WHOLE EXTRACT|AMANITA PANTHERINA WHOLE EXTRACT
C0036442|T121|9601|RXNORM|SCOPOLAMINE|SCOPOLAMINE
C0036442|T121|9601|RXNORM|SCOPOLAMINE|SCOPOLAMINE
C0036442|T121|9601|RXNORM|SCOPOLAMINE|SCOPOLAMINE
C0055147|T121|20610|RXNORM|CETIRIZINE|CETIRIZINE
C0058765|T121|23687|RXNORM|DROXICAM|DROXICAM
C3255938|T109|1306210|RXNORM|HYDROGENATED POLYBUTENE (370 MW)|HYDROGENATED POLYBUTENE (370 MW)
C3255994|T121|1306211|RXNORM|ARACHIDYL PROPIONATE|ARACHIDYL PROPIONATE
C3255995|T121|1306212|RXNORM|ARCTOSTAPHYLOS UVA-URSI LEAF EXTRACT|ARCTOSTAPHYLOS UVA-URSI LEAF EXTRACT
C3857952|T109|1552047|RXNORM|TRIETHANOLAMINE LAURATE|TRIETHANOLAMINE LAURATE
C0051716|T197|17784|RXNORM|AMMONIUM FERROUS SULFATE|AMMONIUM FERROUS SULFATE
C3668706|T121|1441294|RXNORM|ACALYPHA INDICA EXTRACT|ACALYPHA INDICA EXTRACT
C3668707|T121|1441295|RXNORM|ACONITUM LYCOCTONUM EXTRACT|ACONITUM LYCOCTONUM EXTRACT
C3668708|T121|1441296|RXNORM|AGAVE TEQUILANA TOP EXTRACT|AGAVE TEQUILANA TOP EXTRACT
C2936725|T121|1035579|RXNORM|TILETAMINE / ZOLAZEPAM|TILETAMINE / ZOLAZEPAM
C2194078|T121|817235|RXNORM|DOMPERIDONE / SIMETHICONE|DOMPERIDONE / SIMETHICONE
C0146337|T121|57330|RXNORM|TRANILAST|TRANILAST
C1720285|T121|644526|RXNORM|ACTIVATED CHARCOAL / MAGNESIUM HYDROXIDE|ACTIVATED CHARCOAL / MAGNESIUM HYDROXIDE
C2344275|T129|798230|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 6B CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 6B CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C1719978|T121|644529|RXNORM|FLUPHENAZINE / NORTRIPTYLINE|FLUPHENAZINE / NORTRIPTYLINE
C1370123|T121|618597|RXNORM|EICOSAPENTAENOATE|EICOSAPENTAENOATE
C0050521|T121|16784|RXNORM|ACETOXOLONE|ACETOXOLONE
C1579318|T129|845525|RXNORM|JAPANESE ENCEPHALITIS VIRUS VACCINE, INACTIVATED|JAPANESE ENCEPHALITIS VIRUS VACCINE, INACTIVATED
C2047875|T121|820465|RXNORM|CARISOPRODOL / DEXAMETHASONE / IBUPROFEN|CARISOPRODOL / DEXAMETHASONE / IBUPROFEN
C1301985|T121|392449|RXNORM|EPINEPHRINE / FLUOROURACIL|EPINEPHRINE / FLUOROURACIL
C2684354|T121|848929|RXNORM|ACAI BERRY EXTRACT|ACAI BERRY EXTRACT
C0022265|T121|6064|RXNORM|ISOTRETINOIN|ISOTRETINOIN
C0770986|T121|235808|RXNORM|PHENICARBAZIDE|PHENICARBAZIDE
C0022267|T121|6066|RXNORM|ISOXSUPRINE|ISOXSUPRINE
C2980839|T129|1426629|RXNORM|THERMOMYCES LANUGINOSUS ALLERGENIC EXTRACT|THERMOMYCES LANUGINOSUS ALLERGENIC EXTRACT
C0022322|T121|6069|RXNORM|IVERMECTIN|IVERMECTIN
C0022322|T121|6069|RXNORM|IVERMECTIN|IVERMECTIN
C3500692|T121|1315111|RXNORM|CASEIN, LACTOCOCCUS LACTIS CULTURED, AGED|CASEIN, LACTOCOCCUS LACTIS CULTURED, AGED
C2364481|T123|805452|RXNORM|ROMIPLOSTIM|ROMIPLOSTIM
C0009030|T121|2606|RXNORM|CLOPROSTENOL|CLOPROSTENOL
C3531206|T109|1366321|RXNORM|BAMBUSA TEXTILIS STEM EXTRACT|BAMBUSA TEXTILIS STEM EXTRACT
C0009018|T121|2601|RXNORM|CLONIXIN|CLONIXIN
C0031422|T121|8136|RXNORM|OXYPHENISATIN|OXYPHENISATIN
C0009025|T121|2603|RXNORM|CLOPAMIDE|CLOPAMIDE
C3531210|T121|1366326|RXNORM|GLYCINE MAX WHOLE EXTRACT|GLYCINE MAX WHOLE EXTRACT
C1576729|T121|594119|RXNORM|PEGAPTANIB SODIUM|PEGAPTANIB SODIUM
C3859422|T121|1592892|RXNORM|TETRAPEPTIDE-6|TETRAPEPTIDE-6
C3528227|T109|1362140|RXNORM|ASCORBYL TOCOPHERYL MALEATE|ASCORBYL TOCOPHERYL MALEATE
C3153176|T121|1098643|RXNORM|HYPROMELLOSE / TETRAHYDROZOLINE|HYPROMELLOSE / TETRAHYDROZOLINE
C3531211|T109|1366327|RXNORM|OCIMUM GRATISSIMUM LEAF OIL|OCIMUM GRATISSIMUM LEAF OIL
C3531208|T109|1366324|RXNORM|CITRUS JUNOS FRUIT EXTRACT|CITRUS JUNOS FRUIT EXTRACT
C3859817|T129|1594963|RXNORM|TURKEY FEATHER EXTRACT|MELEAGRIS GALLOPAVO FEATHER EXTRACT
C1569608|T121|591622|RXNORM|VARENICLINE|VARENICLINE
C0038143|T197|10030|RXNORM|STANNOUS FLUORIDE|STANNOUS FLUORIDE
C3859819|T129|1594965|RXNORM|SYRIAN HAMSTER HAIR EXTRACT|MESOCRICETUS AURATUS HAIR EXTRACT
C0038149|T125|10032|RXNORM|STANOZOLOL|STANOZOLOL
C2725008|T129|1427171|RXNORM|HEPATITIS B VIRUS SUBTYPE ADW2 HBSAG SURFACE PROTEIN ANTIGEN|HEPATITIS B VIRUS SUBTYPE ADW2 HBSAG SURFACE PROTEIN ANTIGEN
C3256839|T109|1427173|RXNORM|GLYCERYL 1-STEARATE|GLYCERYL 1-STEARATE
C1881354|T121|1427172|RXNORM|L-LACTATE|L-LACTATE
C0055897|T121|21247|RXNORM|CLOBUTINOL|CLOBUTINOL
C2316217|T121|1427179|RXNORM|ANTITHROMBIN ALFA|ANTITHROMBIN ALFA
C3645275|T129|1427178|RXNORM|THYMOCYTE IMMUNOGLOBULIN|THYMOCYTE IMMUNOGLOBULIN
C2980191|T121|1091891|RXNORM|CHLOROXYLENOL / KETOCONAZOLE|CHLOROXYLENOL / KETOCONAZOLE
C0771950|T125|236650|RXNORM|FLUPREDNIDENE|FLUPREDNIDENE
C0936182|T121|282470|RXNORM|DAMIANA LEAF PREPARATION|DAMIANA LEAF PREPARATION
C3486072|T121|1320405|RXNORM|HELIANTHEMUM CANADENSE EXTRACT|HELIANTHEMUM CANADENSE EXTRACT
C3486643|T121|1320407|RXNORM|ANISUM EXTRACT|ANISUM EXTRACT
C3486732|T121|1320409|RXNORM|SPIGELIA MARILANDICA ROOT EXTRACT|SPIGELIA MARILANDICA ROOT EXTRACT
C0001134|T197|236|RXNORM|BOTULISM ANTITOXIN B|ACIDULATED PHOSPHATE FLUORIDE
C0772201|T121|236876|RXNORM|THYMUS GLAND-CALF|THYMUS GLAND-CALF
C2702369|T129|892610|RXNORM|CRAB ALLERGENIC EXTRACT|CRAB ALLERGENIC EXTRACT
C0771562|T121|236303|RXNORM|ISOSPAGLUMIC ACID|ISOSPAGLUMIC ACID
C0771559|T121|236300|RXNORM|ACETIAMINE|ACETIAMINE
C0065086|T197|1310187|RXNORM|LITHIUM BROMIDE|LITHIUM BROMIDE
C3256706|T109|1426402|RXNORM|OCTYLDECANOL|OCTYLDECANOL
C2948243|T121|1043618|RXNORM|EUCALYPTOL / MENTHOL / METHYL SALICYLATE / THYMOL|EUCALYPTOL / MENTHOL / METHYL SALICYLATE / THYMOL
C3486684|T121|1310183|RXNORM|RUMEX CRISPUS TOP EXTRACT|RUMEX CRISPUS TOP EXTRACT
C0752344|T122|1426403|RXNORM|LOW-DENSITY POLYETHYLENE|LOW-DENSITY POLYETHYLENE
C0163272|T121|59161|RXNORM|BRIVUDINE|BRIVUDINE
C0982332|T129|798302|RXNORM|ACELLULAR PERTUSSIS VACCINE, INACTIVATED|ACELLULAR PERTUSSIS VACCINE, INACTIVATED
C2728179|T129|1012140|RXNORM|WHEAT BRAN ALLERGENIC EXTRACT|WHEAT BRAN ALLERGENIC EXTRACT
C2606286|T109|1426400|RXNORM|PONGAMOL|PONGAMOL
C3495122|T121|1310189|RXNORM|JUNIPERUS COMMUNIS FRUIT EXTRACT|JUNIPERUS COMMUNIS FRUIT EXTRACT
C0010637|T121|1426401|RXNORM|CYSTAMINE|CYSTAMINE
C0034330|T130|9036|RXNORM|PYRROLIDONECARBOXYLIC ACID|PYRROLIDONECARBOXYLIC ACID
C3486724|T121|1345679|RXNORM|CULEX PIPIENS PREPARATION|CULEX PIPIENS PREPARATION
C0026388|T121|7019|RXNORM|MOLINDONE|MOLINDONE
C3256177|T109|1426406|RXNORM|PENTAERYTHRITYL TETRAETHYLHEXANOATE|PENTAERYTHRITYL TETRAETHYLHEXANOATE
C0038878|T121|10255|RXNORM|SUPROFEN|SUPROFEN
C0038878|T121|10255|RXNORM|SUPROFEN|SUPROFEN
C0038880|T121|10256|RXNORM|SURAMIN|SURAMIN
C0043366|T121|1099660|RXNORM|XYLAZINE|XYLAZINE
C3255783|T109|1426404|RXNORM|LAUROYL LYSINE|LAUROYL LYSINE
C1966347|T121|746070|RXNORM|LITHIUM ASPARTATE|LITHIUM ASPARTATE
C2740700|T129|899550|RXNORM|YELLOW BIRCH POLLEN EXTRACT|BETULA ALLEGHANIENSIS POLLEN EXTRACT
C1533416|T122|1426405|RXNORM|POLYSORBATE 65|POLYSORBATE 65
C0085274|T005|1368364|RXNORM|HUMAN PARVOVIRUS B19 VIRUS|HUMAN PARVOVIRUS B19 VIRUS
C3256221|T121|1305549|RXNORM|CAMELLIA OLEIFERA LEAF EXTRACT|CAMELLIA OLEIFERA LEAF EXTRACT
C0062687|T130|1305548|RXNORM|HEXYLENE GLYCOL|HEXYLENE GLYCOL
C3485012|T121|1358959|RXNORM|LONICERA CONFUSA WHOLE EXTRACT|LONICERA CONFUSA WHOLE EXTRACT
C0718246|T121||RXNORM|ACTIVATED CHARCOAL / SORBITOL
C2756785|T121|1305545|RXNORM|EUCALYPTUS GLOBULUS LEAF EXTRACT|EUCALYPTUS GLOBULUS LEAF EXTRACT
C3256713|T109|1426408|RXNORM|OLETH-10|POLYOXYL-10 OLEYL ETHER
C0040302|T196|1305547|RXNORM|TITANIUM|TITANIUM
C3696416|T121|1484283|RXNORM|SUCROFERRIC OXYHYDROXIDE|SUCROFERRIC OXYHYDROXIDE
C0066409|T122|29897|RXNORM|METHYLMETHACRYLATE|METHYL METHACRYLATE
C0206816|T121|67182|RXNORM|DILOXANIDE|DILOXANIDE
C0206828|T127|67187|RXNORM|OXERUTINS|OXERUTINS
C2937409|T129|1368357|RXNORM|EMERICELLA NIDULANS ALLERGENIC EXTRACT|ASPERGILLUS NIDULANS ALLERGENIC EXTRACT
C0055152|T122|20615|RXNORM|CETYL ALCOHOL|CETYL ALCOHOL
C0066411|T121|29899|RXNORM|METHYLNALTREXONE|METHYLNALTREXONE
C0002699|T121|739|RXNORM|AMSACRINE|AMSACRINE
C3486728|T121|1310049|RXNORM|PEUMUS BOLDUS LEAF EXTRACT|PEUMUS BOLDUS LEAF EXTRACT
C2740631|T129|899434|RXNORM|HERRING ALLERGENIC EXTRACT|HERRING ALLERGENIC EXTRACT
C3692723|T121|1442508|RXNORM|DAUCUS CAROTA SUBSP. SATIVUS SEED EXTRACT|DAUCUS CAROTA SUBSP. SATIVUS SEED EXTRACT
C3651710|T121|1431226|RXNORM|POLYGLYCERYL-2 DIISOSTEARATE|POLYGLYCERYL-2 DIISOSTEARATE
C0770750|T197|1431227|RXNORM|ZINC PEROXIDE|ZINC PEROXIDE
C0452456|T168|1431224|RXNORM|GRAPEFRUIT JUICE|GRAPEFRUIT JUICE
C3651711|T121|1431225|RXNORM|CISTUS MONSPELIENSIS LEAF EXTRACT|CISTUS MONSPELIENSIS LEAF EXTRACT
C3695956|T109|1484498|RXNORM|ETHYLHEXYL COCOATE|ETHYLHEXYL COCOATE
C2741297|T129|900777|RXNORM|JAPANESE BLACK PINE POLLEN EXTRACT|PINUS THUNBERGII POLLEN EXTRACT
C0019602|T123|5340|RXNORM|HISTIDINE|HISTIDINE
C3282369|T121|1251201|RXNORM|CHLORHEXIDINE / GLYCERIN|CHLORHEXIDINE / GLYCERIN
C0669024|T121|1314374|RXNORM|OLETH-3-PHOSPHATE|OLETH-3-PHOSPHATE
C2979385|T197|1305899|RXNORM|ALUMINUM ZIRCONIUM PENTACHLOROHYDREX GLY|ALUMINUM ZIRCONIUM PENTACHLOROHYDREX GLY
C2242158|T129|763098|RXNORM|POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1)|POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1)
C0003524|T121|1029|RXNORM|APAZONE|APAZONE
C1384515|T121|1039062|RXNORM|CORNSTARCH|CORNSTARCH
C0669026|T121|1314375|RXNORM|OLETH-5|OLETH-5
C2928829|T121|1007915|RXNORM|DIHYDROXYBUTYL ETHER / PROPINOX|DIHYDROXYBUTYL ETHER / PROPINOX
C2928828|T121|1007914|RXNORM|AGAR / MINERAL OIL / PHENOLPHTHALEIN|AGAR / MINERAL OIL / PHENOLPHTHALEIN
C2928831|T121|1007917|RXNORM|HYDROXOCOBALAMIN / IBUPROFEN|HYDROXOCOBALAMIN / IBUPROFEN
C2928830|T121|1007916|RXNORM|ALUMINUM OXIDE / TRICLOSAN|ALUMINUM OXIDE / TRICLOSAN
C2928825|T121|1007911|RXNORM|ALUMINUM HYDROXIDE / ALUMINUM SUBACETATE|ALUMINUM HYDROXIDE / ALUMINUM SUBACETATE
C2928824|T121|1007910|RXNORM|METHACYCLINE / MURAMIDASE|METHACYCLINE / MURAMIDASE
C2928827|T121|1007913|RXNORM|AMYL SALICYLATE / HEXYLNICOTINATE|AMYL SALICYLATE / HEXYLNICOTINATE
C2928826|T121|1007912|RXNORM|BENZOCAINE / BENZYL BENZOATE|BENZOCAINE / BENZYL BENZOATE
C1875287|T121|690133|RXNORM|HYPROMELLOSE / NAPHAZOLINE|HYPROMELLOSE / NAPHAZOLINE
C2928833|T121|1007919|RXNORM|5-METHYL-8-HYDROXYQUINOLINE / TILBROQUINOL|5-METHYL-8-HYDROXYQUINOLINE / TILBROQUINOL
C2928832|T121|1007918|RXNORM|LACTATE / NONOXYNOL-9|LACTATE / NONOXYNOL-9
C3474130|T121|1310041|RXNORM|CITRUS JUNOS SEED EXTRACT|CITRUS JUNOS SEED EXTRACT
C0064725|T197|1593125|RXNORM|LEAD TETROXIDE|LEAD TETROXIDE
C3859491|T129|1593128|RXNORM|MENINGOCOCCAL GROUP B VACCINE|MENINGOCOCCAL GROUP B VACCINE
C0034257|T121|8997|RXNORM|PYRIDINOLCARBAMATE|PYRIDINOLCARBAMATE
C2929169|T121|1008262|RXNORM|ACETAMINOPHEN / DOXYLAMINE / SALICYLAMIDE|ACETAMINOPHEN / DOXYLAMINE / SALICYLAMIDE
C2929170|T121|1008263|RXNORM|ASCORBIC ACID / BIOTIN / FOLIC ACID / NIACIN / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|ASCORBIC ACID / BIOTIN / FOLIC ACID / NIACIN / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C2929167|T121|1008260|RXNORM|CHLORPHENIRAMINE / DIHYDROCODEINE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / DIHYDROCODEINE / PSEUDOEPHEDRINE
C0304936|T121|91498|RXNORM|LIVER,DESICCATED|LIVER,DESICCATED
C2929174|T121|1008267|RXNORM|DIMETHICONE / TRICLOSAN|DIMETHICONE / TRICLOSAN
C2929171|T121|1008264|RXNORM|CALCIUM CARBONATE / ERGOCALCIFEROL|CALCIUM CARBONATE / ERGOCALCIFEROL
C2929172|T121|1008265|RXNORM|DOCUSATE / SPERMACETI|DOCUSATE / SPERMACETI
C0360736|T121|108249|RXNORM|DILOXANIDE / METRONIDAZOLE|DILOXANIDE / METRONIDAZOLE
C2929176|T121|1008269|RXNORM|BAMETHAN / NIACIN|BAMETHAN / NIACIN
C0052820|T121|18651|RXNORM|AZOSEMIDE|AZOSEMIDE
C3282869|T168|1311589|RXNORM|EMPETRUM NIGRUM FRUIT JUICE|EMPETRUM NIGRUM FRUIT JUICE
C0301271|T121|89698|RXNORM|GAMBOGE|GAMBOGE
C0010980|T121|3108|RXNORM|DAPSONE|DAPSONE
C0010980|T121|3108|RXNORM|DAPSONE|DAPSONE
C0011015|T195|3109|RXNORM|DAUNORUBICIN|DAUNORUBICIN
C0010976|T121|3105|RXNORM|DANTROLENE|DANTROLENE
C0010934|T195|3100|RXNORM|DACTINOMYCIN|DACTINOMYCIN
C0010961|T125|3102|RXNORM|DANAZOL|DANAZOL
C0033056|T121|8673|RXNORM|FEPRAZONE|FEPRAZONE
C0937623|T121|283563|RXNORM|GAMMA LINOLEIC ACID|GAMMA LINOLEIC ACID
C0937620|T121|283560|RXNORM|ECHINACEA, AERIAL PARTS|ECHINACEA, AERIAL PARTS
C0937626|T121|283566|RXNORM|GRAPE SEED PROANTHOCYANIDINS|GRAPE SEED PROANTHOCYANIDINS
C3267333|T121|1312728|RXNORM|SCHINUS TEREBINTHIFOLIUS WHOLE EXTRACT|SCHINUS TEREBINTHIFOLIUS WHOLE EXTRACT
C0937624|T121|283564|RXNORM|GAMMA LINOLENIC OIL|GAMMA LINOLENIC OIL
C3496075|T121|1315118|RXNORM|GREEN BELL PEPPER EXTRACT|GREEN BELL PEPPER EXTRACT
C3256651|T121|1312724|RXNORM|TILIA CORDATA WOOD EXTRACT|TILIA CORDATA WOOD EXTRACT
C3267319|T121|1312727|RXNORM|PPG-2 METHYL ETHER|PPG-2 METHYL ETHER
C3500694|T121|1315114|RXNORM|DUNGENESS CRAB, COOKED PREPARATION|DUNGENESS CRAB, COOKED PREPARATION
C3488961|T121|1312721|RXNORM|POLYETHYLENE GLYCOL 700|POLYETHYLENE GLYCOL 700
C3256427|T121|1312720|RXNORM|PHYLLOSTACHYS RETICULATA RESIN|PHYLLOSTACHYS RETICULATA RESIN
C3256638|T121|1312723|RXNORM|POLYISOBUTYLENE (75000 MW)|POLYISOBUTYLENE (75000 MW)
C3256612|T121|1312722|RXNORM|DULSE EXTRACT|DULSE EXTRACT
C3714959|T121|1545038|RXNORM|ANAMIRTA COCCULUS WHOLE EXTRACT|ANAMIRTA COCCULUS WHOLE EXTRACT
C0014927|T125|4094|RXNORM|ESTRIOL|ESTRIOL
C0014938|T125|4099|RXNORM|ESTROGENS, CONJUGATED (USP)|ESTROGENS, CONJUGATED (USP)
C0014938|T125|4099|RXNORM|ESTROGENS, CONJUGATED (USP)|ESTROGENS, CONJUGATED (USP)
C0014938|T125|4099|RXNORM|ESTROGENS, CONJUGATED (USP)|ESTROGENS, CONJUGATED (USP)
C0887557|T127|267366|RXNORM|SODIUM ASCORBATE|SODIUM ASCORBATE
C3651746|T121|1429391|RXNORM|GLECHOMA LONGITUBA TOP EXTRACT|GLECHOMA LONGITUBA TOP EXTRACT
C0106940|T121|47295|RXNORM|BOVINE CARTILAGE EXTRACT|BOVINE CARTILAGE EXTRACT
C3256757|T121|1311638|RXNORM|CAPRYL METHICONE|CAPRYL METHICONE
C3256322|T109|1311639|RXNORM|ACETIC MONOETHANOLAMIDE|ACETIC MONOETHANOLAMIDE
C3255950|T121|1311636|RXNORM|MAHONIA AQUIFOLIUM FRUITING TOP EXTRACT|MAHONIA AQUIFOLIUM FRUITING TOP EXTRACT
C2983983|T121|1311637|RXNORM|ANISACRIL|ANISACRIL
C0025417|T197|1311634|RXNORM|MERCURIC CHLORIDE|MERCURIC CHLORIDE
C1135135|T121|337525|RXNORM|ERLOTINIB|ERLOTINIB
C3255774|T121|1311632|RXNORM|LYCIUM BARBARUM FRUIT EXTRACT|LYCIUM BARBARUM FRUIT EXTRACT
C1135132|T121|337523|RXNORM|IXABEPILONE|IXABEPILONE
C0529351|T121|136198|RXNORM|DARIFENACIN|DARIFENACIN
C0303540|T197|1311631|RXNORM|STRONTIUM BROMIDE|STRONTIUM BROMIDE
C2928582|T121|1007666|RXNORM|BROMELAINS / TRYPSIN|BROMELAINS / TRYPSIN
C2928581|T121|1007665|RXNORM|CARBOMER / MANNITOL|CARBOMER / MANNITOL
C2928580|T121|1007664|RXNORM|GLYCOL SALICYLATE / HISTAMINE / METHYLNICOTINATE|GLYCOL SALICYLATE / HISTAMINE / METHYLNICOTINATE
C2928579|T121|1007663|RXNORM|MAGNESIUM THIOSULFATE / SODIUM THIOSULFATE|MAGNESIUM THIOSULFATE / SODIUM THIOSULFATE
C2928578|T121|1007662|RXNORM|CHLOROXYLENOL / MENTHOL|CHLOROXYLENOL / MENTHOL
C2928577|T121|1007661|RXNORM|CAFFEINE / PHENYLTOLOXAMINE|CAFFEINE / PHENYLTOLOXAMINE
C2928576|T121|1007660|RXNORM|DOG HAIR EXTRACT / DOG SKIN EXTRACT|DOG HAIR EXTRACT / DOG SKIN EXTRACT
C3710012|T109|1488815|RXNORM|ISODON RUBESCENS TOP EXTRACT|ISODON RUBESCENS TOP EXTRACT
C3710011|T168|1488814|RXNORM|BLACK CURRANT JUICE EXTRACT|BLACK CURRANT JUICE
C3710014|T109|1488817|RXNORM|VERATRUM NIGRUM FLOWERING TOP EXTRACT|VERATRUM NIGRUM FLOWERING TOP EXTRACT
C3651744|T121|1429394|RXNORM|OCIMUM GRATISSIMUM WHOLE EXTRACT|OCIMUM GRATISSIMUM WHOLE EXTRACT
C2928277|T121|1007355|RXNORM|CALCIUM CARBONATE / MONOFLUOROPHOSPHATE|CALCIUM CARBONATE / MONOFLUOROPHOSPHATE
C2928585|T121|1007669|RXNORM|MOMETASONE / SALICYLIC ACID|MOMETASONE / SALICYLIC ACID
C2928584|T121|1007668|RXNORM|FLUOCINOLONE / LIDOCAINE|FLUOCINOLONE / LIDOCAINE
C0061377|T121|25834|RXNORM|GLUCAMETACIN|GLUCAMETACIN
C2928276|T121|1007354|RXNORM|CHLORPHENIRAMINE / DIHYDROCODEINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / DIHYDROCODEINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C2726168|T129|883414|RXNORM|TURNIP ALLERGENIC EXTRACT|BRASSICA RAPA ALLERGENIC EXTRACT
C0717808|T121|214603|RXNORM|GUAIFENESIN / HYDROCODONE / PHENYLEPHRINE|GUAIFENESIN / HYDROCODONE / PHENYLEPHRINE
C2928275|T121|1007353|RXNORM|ASPIRIN / CHLORPHENIRAMINE / DEXTROMETHORPHAN|ASPIRIN / CHLORPHENIRAMINE / DEXTROMETHORPHAN
C0717805|T121|214600|RXNORM|GUAIFENESIN / THEOPHYLLINE|GUAIFENESIN / THEOPHYLLINE
C0717811|T129|214606|RXNORM|HAEMOPHILUS B CONJUGATE VACCINE|HAEMOPHILUS B CONJUGATE VACCINE
C0717809|T121|214604|RXNORM|GUAIFENESIN / HYDROCODONE / PSEUDOEPHEDRINE|GUAIFENESIN / HYDROCODONE / PSEUDOEPHEDRINE
C3537211|T121|1432797|RXNORM|RICINUS COMMUNIS WHOLE EXTRACT|RICINUS COMMUNIS WHOLE EXTRACT
C0935989|T121|282388|RXNORM|IMATINIB|IMATINIB
C3663292|T121|1432794|RXNORM|OXYTROPIS LAMBERTII TOP EXTRACT|OXYTROPIS LAMBERTII TOP EXTRACT
C3645144|T121|1426701|RXNORM|SULFOOLEATE|SULFOOLEATE
C3265178|T109|1426703|RXNORM|PROSOLV SMCC 50|PROSOLV SMCC 50
C2928272|T121|1007350|RXNORM|CHROMOUS CHLORIDE / COPPER SULFATE / MANGANESE SULFATE / SELENIOUS ACID / ZINC SULFATE|CHROMOUS CHLORIDE / COPPER SULFATE / MANGANESE SULFATE / SELENIOUS ACID / ZINC SULFATE
C3486568|T121|1426705|RXNORM|MUCOR CIRCINELLOIDES F. LUSITANICUS PREPARATION|MUCOR CIRCINELLOIDES F. LUSITANICUS PREPARATION
C0166894|T121|1426704|RXNORM|NEUROTROPHIN 4|NEUROTROPHIN 4
C3539019|T121|1435389|RXNORM|ECKLONIA CAVA EXTRACT|ECKLONIA CAVA EXTRACT
C0251504|T121|74667|RXNORM|ZALEPLON|ZALEPLON
C1827962|T121|687096|RXNORM|BENZOCAINE / CHLOROXYLENOL|BENZOCAINE / CHLOROXYLENOL
C3255758|T121|1358486|RXNORM|ETHYL MENTHANE CARBOXAMIDE|ETHYL MENTHANE CARBOXAMIDE
C0069174|T109|1358484|RXNORM|NYLON 12|NYLON 12
C3505489|T109|1358485|RXNORM|LAURYL METHACRYLATE - GLYCOL DIMETHACRYLATE CROSSPOLYMER|LAURYL METHACRYLATE - GLYCOL DIMETHACRYLATE CROSSPOLYMER
C3505488|T121|1358482|RXNORM|CLEMATIS CHINENSIS ROOT EXTRACT|CLEMATIS CHINENSIS ROOT EXTRACT
C0043944|T121|1358483|RXNORM|1,3-DIMETHYLUREA|1,3-DIMETHYLUREA
C0031262|T122|8091|RXNORM|PETROLATUM|PETROLATUM
C0031262|T122|8091|RXNORM|PETROLATUM|PETROLATUM
C0048470|T121|15202|RXNORM|ARGATROBAN|ARGATROBAN
C3256039|T121|1307792|RXNORM|DIHYDROXYPROPYL PEG-5 LINOLEAMMONIUM CHLORIDE|DIHYDROXYPROPYL PEG-5 LINOLEAMMONIUM CHLORIDE
C3475263|T109|1307790|RXNORM|CALENDULA OFFICINALIS SEED OIL|CALENDULA OFFICINALIS SEED OIL
C3473227|T121|1307791|RXNORM|LITHOSPERMUM ERYTHRORHIZON ROOT EXTRACT|LITHOSPERMUM ERYTHRORHIZON ROOT EXTRACT
C1434716|T197|1307797|RXNORM|BARIUM CHROMATE|BARIUM CHROMATE
C3255860|T121|1307794|RXNORM|PANAX JAPONICUS ROOT EXTRACT|PANAX JAPONICUS ROOT EXTRACT
C3256178|T109|1358489|RXNORM|PENTAERYTHRITYL TETRAISOSTEARATE|PENTAERYTHRITYL TETRAISOSTEARATE
C3665151|T121|1435388|RXNORM|CHELIDONIUM MAJUS FLOWERING TOP EXTRACT|CHELIDONIUM MAJUS FLOWERING TOP EXTRACT
C2701227|T129|852011|RXNORM|COAST SAGE POLLEN EXTRACT|ARTEMISIA CALIFORNICA POLLEN EXTRACT
C2746078|T121|1100699|RXNORM|LINAGLIPTIN|LINAGLIPTIN
C2701231|T130|852015|RXNORM|CORN POLLEN EXTRACT|ZEA MAYS POLLEN EXTRACT
C2057755|T121|819684|RXNORM|GUAIFENESIN / PSEUDOEPHEDRINE / THEOPHYLLINE|GUAIFENESIN / PSEUDOEPHEDRINE / THEOPHYLLINE
C2242042|T129|762817|RXNORM|RUBELLA VIRUS VACCINE LIVE (WISTAR RA 27-3 STRAIN)|RUBELLA VIRUS VACCINE LIVE (WISTAR RA 27-3 STRAIN)
C3555517|T109|1374805|RXNORM|POLYISOBUTYLENE (800000 MW)|POLYISOBUTYLENE (800000 MW)
C2012664|T121|816111|RXNORM|AMMONIUM CHLORIDE / GUAIFENESIN|AMMONIUM CHLORIDE / GUAIFENESIN
C3700871|T197|1487155|RXNORM|MAGNESIUM PHOSPHATE, MONOBASIC, DIHYDRATE|MAGNESIUM PHOSPHATE, MONOBASIC, DIHYDRATE
C2756198|T129|967721|RXNORM|BREAD MOLD FUNGUS EXTRACT|BREAD MOLD FUNGUS EXTRACT
C3700870|T122|1487156|RXNORM|SODIUM LAUROYL METHYL ISETHIONATE|SODIUM LAUROYL METHYL ISETHIONATE
C1828451|T121|687225|RXNORM|ALBUTEROL / BECLOMETHASONE|ALBUTEROL / BECLOMETHASONE
C1828057|T121|687227|RXNORM|BISMUTH BISKALCITRATE|BISMUTH BISKALCITRATE
C0885849|T121|266364|RXNORM|BEARBERRY PREPARATION|UVA URSI
C0279218|T129|80726|RXNORM|EDRECOLOMAB|EDRECOLOMAB
C1874705|T121|691201|RXNORM|CANTHARIDIN / PODOPHYLLIN / SALICYLIC ACID|CANTHARIDIN / PODOPHYLLIN / SALICYLIC ACID
C3555538|T121|1373354|RXNORM|MYROTHAMNUS FLABELLIFOLIA LEAF EXTRACT|MYROTHAMNUS FLABELLIFOLIA LEAF EXTRACT
C2746107|T129|901624|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 19A CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 19A CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C0310589|T121|97016|RXNORM|VITAMIN A / VITAMIN D|VITAMIN A / VITAMIN D
C0034338|T130|1373350|RXNORM|PYRUVALDEHYDE|PYRUVALDEHYDE
C3555539|T109|1373353|RXNORM|CETYL DIMETHICONE 25|CETYL DIMETHICONE 25
C0054465|T197|1373352|RXNORM|CALCIUM BICARBONATE|CALCIUM BICARBONATE
C0075430|T122|1374803|RXNORM|SUCCINIC ANHYDRIDE|SUCCINIC ANHYDRIDE
C0608826|T121|161203|RXNORM|ACEPROMETAZINE|ACEPROMETAZINE
C2746111|T129|901628|RXNORM|STREPTOCOCCUS PNEUMONIAE SEROTYPE 3 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|STREPTOCOCCUS PNEUMONIAE SEROTYPE 3 CAPSULAR ANTIGEN DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C3256375|T121|1313186|RXNORM|MYRISTOYL-PALMITOYL OXOSTEARAMIDE-ARACHAMIDE MEA|MYRISTOYL-PALMITOYL OXOSTEARAMIDE-ARACHAMIDE MEA
C3256768|T109|1313187|RXNORM|GLUCAMINE|GLUCAMINE
C3256037|T121|1313184|RXNORM|DIHYDROGENATED TALLOW PHTHALIC ACID AMIDE|DIHYDROGENATED TALLOW PHTHALIC ACID AMIDE
C2827186|T121|1313185|RXNORM|HYPROMELLOSE ACETATE SUCCINATE 16070722 (3 MM2-S)|HYPROMELLOSE ACETATE SUCCINATE 16070722 (3 MM2-S)
C3486619|T121|1340183|RXNORM|CHONDRODENDRON TOMENTOSUM ROOT EXTRACT|CHONDRODENDRON TOMENTOSUM ROOT EXTRACT
C3255900|T121|1313183|RXNORM|MOTH BEAN EXTRACT|MOTH BEAN EXTRACT
C1095914|T121|1313180|RXNORM|REISHI MUSHROOM PREPARATION|REISHI MUSHROOM PREPARATION
C0040988|T121|10804|RXNORM|TRIFLUPERIDOL|TRIFLUPERIDOL
C0040989|T121|10805|RXNORM|TRIFLUPROMAZINE|TRIFLUPROMAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE|TRIFLUOPERAZINE
C3465012|T123|1313188|RXNORM|CYSTEINE, DL-|CYSTEINE, DL-
C0040987|T121|10803|RXNORM|TRIFLURIDINE|TRIFLURIDINE
C0044550|T121|1592897|RXNORM|1-OCTANESULFONIC ACID|1-OCTANESULFONIC ACID
C0023610|T125|6384|RXNORM|GONADORELIN|GONADORELIN
C0023610|T125|6384|RXNORM|GONADORELIN|GONADORELIN
C0023660|T121|6387|RXNORM|LIDOCAINE|LIDOCAINE
C0023660|T121|6387|RXNORM|LIDOCAINE|LIDOCAINE
C0023660|T121|6387|RXNORM|LIDOCAINE|LIDOCAINE
C0023660|T121|6387|RXNORM|LIDOCAINE|LIDOCAINE
C0023660|T121|6387|RXNORM|LIDOCAINE|LIDOCAINE
C0023660|T121|6387|RXNORM|LIDOCAINE|LIDOCAINE
C0771738|T121|236463|RXNORM|GLICOFOSFOPEPTICAL|GLICOFOSFOPEPTICAL
C2947856|T121|1042859|RXNORM|POTASSIUM BICARBONATE / SODIUM BICARBONATE / SODIUM CITRATE|POTASSIUM BICARBONATE / SODIUM BICARBONATE / SODIUM CITRATE
C0023607|T125|6383|RXNORM|LUTEINIZING HORMONE|LUTEINIZING HORMONE
C3475011|T121|1302454|RXNORM|OMEGA-3 ACID ETHYL ESTERS (USP) / SALMON OIL|OMEGA-3 ACID ETHYL ESTERS (USP) / SALMON OIL
C2929474|T121|1008571|RXNORM|POLYVINYL ALCOHOL / POVIDONE / TETRAHYDROZOLINE|POLYVINYL ALCOHOL / POVIDONE / TETRAHYDROZOLINE
C0054249|T121|19874|RXNORM|BUTOBARBITAL|BUTOBARBITONE
C0541155|T121|141626|RXNORM|COLESEVELAM|COLESEVELAM
C2203707|T121|818798|RXNORM|ASCORBIC ACID / ZINC GLUCONATE|ASCORBIC ACID / ZINC GLUCONATE
C2016181|T121|818791|RXNORM|ERGONOVINE / OXYTOCIN|ERGONOVINE / OXYTOCIN
C3505823|T121|1359426|RXNORM|GLYCYRRHIZINATE|GLYCYRRHIZINATE
C3505821|T121|1359424|RXNORM|BETA-BISABOLOL|BETA-BISABOLOL
C3505820|T121|1359423|RXNORM|PEG & PPG-17-6 COPOLYMER|PEG & PPG-17-6 COPOLYMER
C0051080|T121|1359422|RXNORM|ALANYLGLUTAMINE|ALANYL GLUTAMINE
C3555508|T109|1376095|RXNORM|DICETYLDIMONIUM CHLORIDE|DICETYLDIMONIUM CHLORIDE
C3858054|T121|1551467|RXNORM|BUPROPION / NALTREXONE|BUPROPION / NALTREXONE
C0065527|T197|29164|RXNORM|MAGNESIUM PHOSPHATE|MAGNESIUM PHOSPHATE
C3695957|T109|1484496|RXNORM|DIISOSTEAROYL POLYGLYCERYL-3 DIMER DILINOLEATE|DIISOSTEAROYL POLYGLYCERYL-3 DIMER DILINOLEATE
C0252643|T121|75207|RXNORM|BOSENTAN|BOSENTAN
C0108124|T121|47624|RXNORM|CALCIUM LEVULINATE|CALCIUM LAEVULATE
C0772108|T121|236795|RXNORM|DEMELVERIN|DEMELVERIN
C0060128|T121|24805|RXNORM|FEBANTEL|FEBANTEL
C0772110|T121|236797|RXNORM|ALPHA HYDROXY ACIDS|ALPHA HYDROXY ACIDS
C3555505|T109|1376098|RXNORM|CETYL PEG- PPG-10- 1 DIMETHICONE (HLB 3)|CETYL PEG- PPG-10- 1 DIMETHICONE (HLB 3)
C3666560|T121|1437307|RXNORM|ABELMOSCHUS ESCULENTUS SEED EXTRACT|ABELMOSCHUS ESCULENTUS SEED EXTRACT
C0525145|T109|1371054|RXNORM|METHYLDIETHANOLAMINE|METHYLDIETHANOLAMINE
C0163355|T197|1537801|RXNORM|AQUA REGIA|AQUA REGIA
C0006507|T121|1848|RXNORM|BUTYLATED HYDROXYTOLUENE|BUTYLATED HYDROXYTOLUENE
C0002707|T121|1371051|RXNORM|AMYGDALIN|AMYGDALIN
C3537592|T121|1371053|RXNORM|CASTOR CANADENSIS SCENT GLAND SECRETION PREPARATION|CASTOR CANADENSIS SCENT GLAND SECRETION PREPARATION
C0006491|T121|1841|RXNORM|BUTORPHANOL|BUTORPHANOL
C2929753|T121|1008855|RXNORM|AMPICILLIN / BROVANEXINE|AMPICILLIN / BROVANEXINE
C2929752|T121|1008854|RXNORM|CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE / PHENYLPROPANOLAMINE|CHLORPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C2929755|T121|1008857|RXNORM|PENTOSAN POLYSULFATE / UREA|PENTOSAN POLYSULFATE / UREA
C2929754|T121|1008856|RXNORM|ASCORBIC ACID / MAGNESIUM OXIDE|ASCORBIC ACID / MAGNESIUM OXIDE
C2929749|T121|1008851|RXNORM|INOSITOL / PHYTIC ACID|INOSITOL / PHYTIC ACID
C2929748|T121|1008850|RXNORM|ANISOTROPINE / DIPYRONE|ANISOTROPINE / DIPYRONE
C2929751|T121|1008853|RXNORM|DICHLORODIFLUOROMETHANE / TRICHLOROFLUOROMETHANE|DICHLORODIFLUOROMETHANE / TRICHLOROFLUOROMETHANE
C2929750|T121|1008852|RXNORM|HEMICELLULASE / OX BILE EXTRACT / PANCREATIN / SIMETHICONE|HEMICELLULASE / OX BILE EXTRACT / PANCREATIN / SIMETHICONE
C2587204|T125|4952|RXNORM|THYROTROPIN ALFA (USP)|THYROTROPIN ALFA
C2587204|T125|4952|RXNORM|THYROTROPIN ALFA (USP)|THYROTROPIN ALFA
C2929757|T121|1008859|RXNORM|AMMONIUM CHLORIDE / BETAINE|AMMONIUM CHLORIDE / BETAINE
C2929756|T121|1008858|RXNORM|CETYLPYRIDINIUM / TYROTHRICIN|CETYLPYRIDINIUM / TYROTHRICIN
C0017970|T121|4955|RXNORM|GLYCOPYRROLATE|GLYCOPYRROLATE
C2927904|T121|1006981|RXNORM|FRAMYCETIN / NAPHAZOLINE|FRAMYCETIN / NAPHAZOLINE
C2927903|T121|1006980|RXNORM|DIHYDROERGOTAMINE / PROPYPHENAZONE|DIHYDROERGOTAMINE / PROPYPHENAZONE
C2927906|T121|1006983|RXNORM|ALLANTOIN / THYMOL|ALLANTOIN / THYMOL
C2927905|T121|1006982|RXNORM|OROTIC ACID / VITAMIN E|OROTIC ACID / VITAMIN E
C2927908|T121|1006985|RXNORM|DEXTRAN / PHENYLBUTAZONE|DEXTRAN / PHENYLBUTAZONE
C2927907|T121|1006984|RXNORM|BROMHEXINE / CEFACLOR|BROMHEXINE / CEFACLOR
C2927910|T121|1006987|RXNORM|LINOLEATE / OMEGA-3 ACID ETHYL ESTERS (USP) / VITAMIN E|LINOLEATE / OMEGA-3 ACID ETHYL ESTERS (USP) / VITAMIN E
C2927909|T121|1006986|RXNORM|METOCLOPRAMIDE / PANCREATIN / PEPSIN A|METOCLOPRAMIDE / PANCREATIN / PEPSIN A
C2927912|T121|1006989|RXNORM|HEMATOPORPHYRIN / PROCAINE|HEMATOPORPHYRIN / PROCAINE
C2927911|T121|1006988|RXNORM|BRILLIANT GREEN / GENTIAN VIOLET|BRILLIANT GREEN / GENTIAN VIOLET
C3535680|T121|1368377|RXNORM|ILEX PARAGUARIENSIS WHOLE EXTRACT|ILEX PARAGUARIENSIS WHOLE EXTRACT
C3535920|T109|1368376|RXNORM|TRIS(TETRAMETHYLHYDROXYPIPERIDINOL)|TRIS(TETRAMETHYLHYDROXYPIPERIDINOL)
C0067067|T121|1368374|RXNORM|MYRICETIN|MYRICETIN
C0066372|T131|1368373|RXNORM|METHYLEUGENOL|METHYLEUGENOL
C2710463|T109|1368372|RXNORM|BENZOTRIAZOLYL DODECYL P-CRESOL|BENZOTRIAZOLYL DODECYL P-CRESOL
C0006699|T121|1908|RXNORM|CALCIUM GLUCONATE|CALCIUM GLUCONATE
C0006700|T121|1909|RXNORM|CALCIUM GLYCEROPHOSPHATE|CALCIUM GLYCEROPHOSPHATE
C0006698|T121|1907|RXNORM|CALCIUM GLUCARATE|CALCIUM GLUCARATE
C0007072|T126|1242127|RXNORM|GLUCARPIDASE|GLUCARPIDASE
C0006695|T197|1905|RXNORM|CALCIUM FLUORIDE|CALCIUM FLUORIDE
C1611088|T197|1902|RXNORM|CALCIUM CARBIMIDE|CALCIUM CARBIMIDE
C0011824|T125|3292|RXNORM|DEXTROTHYROXINE|DEXTROTHYROXINE
C0006686|T197|1901|RXNORM|CALCIUM CHLORIDE|CALCIUM CHLORIDE
C0301297|T121|1363702|RXNORM|CHLOROTHYMOL|CHLOROTHYMOL
C0286353|T121|1363701|RXNORM|SORBITAN MONOPALMITATE|SORBITAN MONOPALMITATE
C0285753|T121|1363700|RXNORM|DIBUTYL SEBACATE|DIBUTYL SEBACATE
C0063964|T109|1363706|RXNORM|ISOEUGENOL|ISOEUGENOL
C0526161|T121|1363705|RXNORM|LAURIC ACID DIETHANOLAMIDE|LAURIC ACID DIETHANOLAMIDE
C0303442|T197|1363704|RXNORM|MAGNESIUM CARBONATE HYDROXIDE|MAGNESIUM CARBONATE HYDROXIDE
C0000294|T121|44|RXNORM|MANGANESE HVP CHELATE|MESNA
C1875132|T121|692987|RXNORM|ESTRONE / PROGESTERONE|ESTRONE / PROGESTERONE
C0067309|T121|1363709|RXNORM|N,N'-DIPHENYL-4-PHENYLENEDIAMINE|N,N'-DIPHENYL-4-PHENYLENEDIAMINE
C0066367|T130|1363708|RXNORM|METHYLETHYL KETONE|METHYLETHYL KETONE
C0065555|T131|896038|RXNORM|MALACHITE GREEN|MALACHITE GREEN
C3489575|T121|36387|RXNORM|SENNOSIDES, USP|SENNA GLYCOSIDES
C3489575|T121|36387|RXNORM|SENNOSIDES, USP|SENNA GLYCOSIDES
C3489575|T121|36387|RXNORM|SENNOSIDES, USP|SENNA GLYCOSIDES
C0074391|T121|36435|RXNORM|SERTACONAZOLE|SERTACONAZOLE
C0074389|T126|36434|RXNORM|SERRATIOPEPTIDASE|SERRATIOPEPTIDASE
C0074393|T121|36437|RXNORM|SERTRALINE|SERTRALINE
C1302057|T121|392511|RXNORM|ACETAMINOPHEN / CHLORMEZANONE|ACETAMINOPHEN / CHLORMEZANONE
C3487963|T121|1311359|RXNORM|SUS SCROFA URINARY BLADDER PREPARATION|PORCINE URINARY BLADDER PREPARATION
C3487962|T121|1311358|RXNORM|SUS SCROFA URETHRA PREPARATION|PORCINE URETHRA PREPARATION
C2731378|T129|895070|RXNORM|MONGOLIAN GERBIL SKIN ALLERGENIC EXTRACT|MERIONES UNGUICULATUS ALLERGENIC EXTRACT
C3486844|T121|1311350|RXNORM|SUS SCROFA THALAMUS PREPARATION|PORCINE THALAMUS PREPARATION
C2073875|T121|816174|RXNORM|ASPIRIN / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE|ASPIRIN / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE
C3486847|T121|1311355|RXNORM|SUS SCROFA UMBILICAL CORD PREPARATION|PORCINE UMBILICAL CORD PREPARATION
C2955225|T121|1049912|RXNORM|ALUMINUM HYDROXIDE / DIMETHICONE / MAGNESIUM HYDROXIDE|ALUMINUM HYDROXIDE / DIMETHICONE / MAGNESIUM HYDROXIDE
C3486848|T121|1311356|RXNORM|SUS SCROFA URETER PREPARATION|PORCINE URETER PREPARATION
C3256150|T121|1307802|RXNORM|CORYDALIS BUNGEANA FLOWERING-FRUITING TOP EXTRACT|CORYDALIS BUNGEANA FLOWERING-FRUITING TOP EXTRACT
C3256514|T109|1307803|RXNORM|CLOVE STEM OIL|CLOVE STEM OIL
C3474977|T109|1307800|RXNORM|CAMELLIA KISSII SEED OIL|CAMELLIA KISSII SEED OIL
C0174148|T197|1307801|RXNORM|BARIUM OXIDE|BARIUM OXIDE
C3256658|T121|1307806|RXNORM|ARTEMISIA UMBELLIFORMIS FLOWER EXTRACT|ARTEMISIA UMBELLIFORMIS FLOWER EXTRACT
C3256796|T109|1307807|RXNORM|OPHIOPOGON JAPONICUS ROOT EXTRACT|OPHIOPOGON JAPONICUS ROOT EXTRACT
C3255673|T121|1307804|RXNORM|HEDYCHIUM CORONARIUM ROOT EXTRACT|HEDYCHIUM CORONARIUM ROOT EXTRACT
C3486293|T121|1307805|RXNORM|LITCHI CHINENSIS SEED EXTRACT|LITCHI CHINENSIS SEED EXTRACT
C3496398|T121|1367497|RXNORM|PLANTAGO ASIATICA EXTRACT|PLANTAGO ASIATICA EXTRACT
C3531672|T121|1367496|RXNORM|PINUS DENSIFLORA ROOT EXTRACT|PINUS DENSIFLORA ROOT EXTRACT
C3465258|T121|1307808|RXNORM|ISATIS TINCTORIA ROOT EXTRACT|ISATIS TINCTORIA ROOT EXTRACT
C3256043|T168|1307809|RXNORM|EUROPEAN HAZELNUT OIL|EUROPEAN HAZELNUT OIL
C3531669|T121|1367493|RXNORM|COCOS NUCIFERA WHOLE EXTRACT|COCOS NUCIFERA WHOLE EXTRACT
C3531668|T109|1367492|RXNORM|AMINOPROPYL DIHYDROGEN PHOSPHATE|AMINOPROPYL DIHYDROGEN PHOSPHATE
C3528057|T109|1361659|RXNORM|DIMETHICONE-VINYL DIMETHICONE CROSSPOLYMER|DIMETHICONE/VINYL DIMETHICONE CROSSPOLYMER (SOFT PARTICLE)
C3486397|T121|1353218|RXNORM|ARANEUS DIADEMATUS PREPARATION|ARANEUS DIADEMATUS PREPARATION
C3486565|T121|1353219|RXNORM|PSEUDOGNAPHALIUM LUTEOALBUM LEAF EXTRACT|PSEUDOGNAPHALIUM LUTEOALBUM LEAF EXTRACT
C1572601|T168|1358977|RXNORM|CRANBERRY JUICE|CRANBERRY JUICE
C1327962|T168|1358975|RXNORM|POMEGRANATE JUICE|POMEGRANATE JUICE
C0937766|T121|283674|RXNORM|ARNICA FLOWERS EXTRACT|ARNICA FLOWERS EXTRACT
C3255690|T121|1310519|RXNORM|LIMONIA ACIDISSIMA WOOD EXTRACT|LIMONIA ACIDISSIMA WOOD EXTRACT
C1879850|T121|1310510|RXNORM|BISOCTRIZOLE|BISOCTRIZOLE
C2962867|T121|1087297|RXNORM|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / NIACIN / POLYSACCHARIDE IRON COMPLEX|ASCORBIC ACID / FERROUS FUMARATE / FOLIC ACID / NIACIN / POLYSACCHARIDE IRON COMPLEX
C3256420|T168|1310512|RXNORM|MALTOSE SYRUP|MALTOSE SYRUP
C0079466|T121|40114|RXNORM|GUANFACINE|GUANFACINE
C0079466|T121|40114|RXNORM|GUANFACINE|GUANFACINE
C0022948|T126|1310514|RXNORM|LACTOPEROXIDASE|LACTOPEROXIDASE
C3465210|T121|1310517|RXNORM|ANCHOVY PREPARATION|ANCHOVY PREPARATION
C0772425|T121|237087|RXNORM|BISMUTH CAMPHOCARBONATE|BISMUTH CAMPHOCARBONATE
C0520472|T121|132889|RXNORM|LEVONORDEFRIN|LEVONORDEFRIN
C2928683|T121|1007768|RXNORM|CALCIUM LACTATE / ERGOCALCIFEROL|CALCIUM LACTATE / ERGOCALCIFEROL
C0107497|T121|47461|RXNORM|BUTENAFINE|BUTENAFINE
C0020406|T121|1426887|RXNORM|HYGROMYCIN B|HYGROMYCIN B
C0056036|T197|1426884|RXNORM|COBALTOUS CHLORIDE|COBALTOUS CHLORIDE
C0544348|T121|1426885|RXNORM|CHONDRUS PREPARATION|CHONDRUS PREPARATION
C2927981|T121|1007058|RXNORM|BUCLIZINE / VITAMIN B6|BUCLIZINE / VITAMIN B6
C2927982|T121|1007059|RXNORM|ACETAMINOPHEN / CAFFEINE / PAMABROM / VITAMIN B6|ACETAMINOPHEN / CAFFEINE / PAMABROM / VITAMIN B6
C3833357|T121|1541241|RXNORM|PETASITES HYBRIDUS ROOT EXTRACT|PETASITES HYBRIDUS ROOT EXTRACT
C2927977|T121|1007054|RXNORM|ALLANTOIN / CAMPHOR / MENTHOL|ALLANTOIN / CAMPHOR / MENTHOL
C2927978|T121|1007055|RXNORM|NIACIN / NIACINAMIDE|NIACIN / NIACINAMIDE
C2927979|T121|1007056|RXNORM|CETRIMIDE / DIMETHICONE|CETRIMIDE / DIMETHICONE
C2927980|T121|1007057|RXNORM|LYSINE / PROLINE|LYSINE / PROLINE
C2927973|T121|1007050|RXNORM|DEXTROMETHORPHAN / GUAIACOLSULFONATE / PHENYLEPHRINE|DEXTROMETHORPHAN / GUAIACOLSULFONATE / PHENYLEPHRINE
C2927975|T121|1007052|RXNORM|DEVIL'S CLAW PREPARATION / HAWTHORN FLOWER EXTRACT|DEVIL'S CLAW PREPARATION / HAWTHORN FLOWER EXTRACT
C2927976|T121|1007053|RXNORM|EPHEDRINE / PHOLCODINE|EPHEDRINE / PHOLCODINE
C3489001|T109|1309329|RXNORM|CRYPTOCARYA AGATHOPHYLLA LEAF OIL|CRYPTOCARYA AGATHOPHYLLA LEAF OIL
C3489002|T109|1309328|RXNORM|MELISSA OFFICINALIS LEAF OIL|MELISSA OFFICINALIS LEAF OIL
C0612505|T121|163426|RXNORM|TIOCLOMAROL|TIOCLOMAROL
C0292857|T197|1542454|RXNORM|CALCIUM CHLORATE DIHYDRATE|CALCIUM CHLORATE DIHYDRATE
C2353893|T129|819300|RXNORM|GOLIMUMAB|GOLIMUMAB
C3488914|T109|1309325|RXNORM|NOTOPTERYGIUM FRANHETII ROOT EXTRACT|NOTOPTERYGIUM FRANHETII ROOT EXTRACT
C2080611|T121|819306|RXNORM|GUAIFENESIN / HYDROCODONE / PHENIRAMINE / PHENYLPROPANOLAMINE / PYRILAMINE|GUAIFENESIN / HYDROCODONE / PHENIRAMINE / PHENYLPROPANOLAMINE / PYRILAMINE
C3488930|T109|1309327|RXNORM|MENTHA ARVENSIS FLOWERING TOP EXTRACT|MENTHA ARVENSIS FLOWERING TOP EXTRACT
C3488931|T109|1309326|RXNORM|MENTHA PIPERITA LEAF EXTRACT|PEPPERMINT LEAF EXTRACT
C1098320|T121|321064|RXNORM|OLMESARTAN|OLMESARTAN
C2928859|T121|1007946|RXNORM|ASCORBIC ACID / DOCUSATE / FOLIC ACID / IRON CARBONYL / VITAMIN B 12|ASCORBIC ACID / DOCUSATE / FOLIC ACID / IRON CARBONYL / VITAMIN B 12
C2928860|T121|1007947|RXNORM|ACETAMINOPHEN / RACEMETHIONINE|ACETAMINOPHEN / RACEMETHIONINE
C0981959|T129|314443|RXNORM|RHIZOPUS ORYZAE EXTRACT|RHIZOPUS ARRHIZUS VAR. ARRHIZUS EXTRACT
C2080565|T121|814304|RXNORM|AMMONIUM CHLORIDE / PHENYLPROPANOLAMINE|AMMONIUM CHLORIDE / PHENYLPROPANOLAMINE
C2928857|T121|1007944|RXNORM|DOBESILIC ACID / FLUNARIZINE|DOBESILIC ACID / FLUNARIZINE
C2193842|T121|1007586|RXNORM|AMPICILLIN / FLOXACILLIN|AMPICILLIN / FLOXACILLIN
C2928505|T121|1007587|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / DEXTROMETHORPHAN|ACETAMINOPHEN / CHLORPHENIRAMINE / DEXTROMETHORPHAN
C2928503|T121|1007584|RXNORM|ACELLULAR PERTUSSIS VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED|ACELLULAR PERTUSSIS VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED
C2928504|T121|1007585|RXNORM|PAPAVERETUM / SCOPOLAMINE|PAPAVERETUM / SCOPOLAMINE
C2928501|T121|1007582|RXNORM|CHLORPROPAMIDE / PHENFORMIN|CHLORPROPAMIDE / PHENFORMIN
C2928502|T121|1007583|RXNORM|CHLORDIAZEPOXIDE / ESTROGENS, ESTERIFIED (USP)|CHLORDIAZEPOXIDE / ESTROGENS, ESTERIFIED (USP)
C2025581|T121|1007580|RXNORM|AMBROXOL / CEFADROXIL|AMBROXOL / CEFADROXIL
C2928500|T121|1007581|RXNORM|CLOTRIMAZOLE / NIMORAZOLE|CLOTRIMAZOLE / NIMORAZOLE
C0002371|T197|612|RXNORM|ALUMINUM HYDROXIDE|ALUMINIUM HYDROXIDE
C2936691|T121|1007942|RXNORM|QUINIDINE / VERAPAMIL|QUINIDINE / VERAPAMIL
C0004521|T195|1272|RXNORM|AZTREONAM|AZTREONAM
C0004521|T195|1272|RXNORM|AZTREONAM|AZTREONAM
C0002370|T121|611|RXNORM|ALUMINUM ASPIRIN|ALUMINUM ASPIRIN
C2194236|T121|818876|RXNORM|DIETHYLAMINE SALICYLATE / MYRTECAINE|DIETHYLAMINE SALICYLATE / MYRTECAINE
C2928506|T121|1007588|RXNORM|EVENING PRIMROSE OIL / GAMMA-LINOLENATE|EVENING PRIMROSE OIL / GAMMA-LINOLENATE
C2928507|T121|1007589|RXNORM|DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED|DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED
C2928200|T121|1007278|RXNORM|ISOPROPYL ALCOHOL / SALICYLIC ACID|ISOPROPYL ALCOHOL / SALICYLIC ACID
C2928201|T121|1007279|RXNORM|INVERT SUGAR / SODIUM CHLORIDE|INVERT SUGAR / SODIUM CHLORIDE
C2928854|T121|1007940|RXNORM|LIDOCAINE / TYROTHRICIN|LIDOCAINE / TYROTHRICIN
C2928192|T121|1007270|RXNORM|INOSITOL / NIACIN|INOSITOL / NIACIN
C2928193|T121|1007271|RXNORM|CATALASE / ORGOTEIN|CATALASE / ORGOTEIN
C2928194|T121|1007272|RXNORM|ALANINE / ARGININE / ASPARTATE / GLUCOSE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / ASPARTATE / GLUCOSE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C0033509|T130|8793|RXNORM|PROPYLIODONE|PROPYLIODONE
C2928196|T121|1007274|RXNORM|GLUCOSE / POTASSIUM CHLORIDE / POTASSIUM LACTATE / SODIUM CHLORIDE / SODIUM PHOSPHATE, MONOBASIC|GLUCOSE / POTASSIUM CHLORIDE / POTASSIUM LACTATE / SODIUM CHLORIDE / SODIUM PHOSPHATE, MONOBASIC
C2928197|T121|1007275|RXNORM|ETHANOL / RESORCINOL|ETHANOL / RESORCINOL
C2928198|T121|1007276|RXNORM|CALCIUM PHOSPHATE / MELATONIN|CALCIUM PHOSPHATE / MELATONIN
C2928199|T121|1007277|RXNORM|BENZOCAINE / ETHANOL / TANNIC ACID|BENZOCAINE / ETHANOL / TANNIC ACID
C1271607|T125|388084|RXNORM|LUTROPIN ALFA|LUTROPIN ALFA
C1119842|T121|325524|RXNORM|GARLIC POWDER|GARLIC POWDER
C1119920|T121|325527|RXNORM|CORIANDER EXTRACT|CORIANDER EXTRACT
C3644741|T109|1425615|RXNORM|CITRUS LIMON SEED OIL|CITRUS LIMON SEED OIL
C1118156|T121|325521|RXNORM|THYROID (BEEF)|THYROID (BEEF)
C1117900|T121|325520|RXNORM|POTASSIUM OXYQUINOLONE|POTASSIUM OXYQUINOLONE
C1118917|T116|325523|RXNORM|LYMPHOCYTE IMMUNE GLOBULIN, RABBIT|LYMPHOCYTE IMMUNE GLOBULIN, RABBIT
C1118183|T121|325522|RXNORM|TISSUE RESPIRATORY FACTOR|TISSUE RESPIRATORY FACTOR
C0033501|T121|1311134|RXNORM|PROPYL GALLATE|PROPYL GALLATE
C0000966|T109|1311137|RXNORM|ACETALDEHYDE|ACETALDEHYDE
C3256644|T121|1314324|RXNORM|POLYQUATERNIUM-7 (76-24 ACRYLAMIDE-DADMAC; 120 KD)|POLYQUATERNIUM-7 (76-24 ACRYLAMIDE-DADMAC; 120 KD)
C0022071|T196|1311131|RXNORM|IRIDIUM|IRIDIUM
C0029383|T196|1311130|RXNORM|OSMIUM|OSMIUM
C3255781|T121|1311133|RXNORM|LARREA TRIDENTA TOP EXTRACT|LARREA TRIDENTA TOP EXTRACT
C3497608|T121|1314320|RXNORM|OREGANO LEAF OIL|OREGANO LEAF OIL
C0049865|T109|1362616|RXNORM|7-DEHYDROCHOLESTEROL|7-DEHYDROCHOLESTEROL
C0093558|T109|1362615|RXNORM|2-OCTANOL|2-OCTANOL
C0074730|T197|1311138|RXNORM|SODIUM BROMIDE|SODIUM BROMIDE
C3495674|T121|1314329|RXNORM|ACETYL HEXAPEPTIDE-8|ACETYL HEXAPEPTIDE-8
C0046202|T121|1314328|RXNORM|2-HYDROXYETHYL ACRYLATE|2-HYDROXYETHYL ACRYLATE
C1509576|T121|1421621|RXNORM|METHYL GLUCOSE DIOLEATE|METHYL GLUCOSE DIOLEATE
C3643362|T109|1421627|RXNORM|IPOMOEA PES-CAPRAE FLOWERING TOP EXTRACT|IPOMOEA PES-CAPRAE FLOWERING TOP EXTRACT
C3818752|T121|1493084|RXNORM|BOS TAURUS UTERUS PREPARATION|BOS TAURUS UTERUS PREPARATION
C3255769|T109|1368707|RXNORM|ETHYLHEXYL HYDROXYSTEARATE|ETHYLHEXYL HYDROXYSTEARATE
C3486598|T121|1313322|RXNORM|BEEF HEART PREPARATION|BEEF HEART PREPARATION
C3709437|T121|1487367|RXNORM|HYDROXYETHYL CELLULOSE (280 MPA.S AT 5%)|HYDROXYETHYL CELLULOSE (280 MPA.S AT 5%)
C0072186|T121|34658|RXNORM|PROPIONIC ACID|PROPIONIC ACID
C1725493|T121|1366627|RXNORM|STEARETH-30|STEARETH-30
C3538618|T121|1373160|RXNORM|RHUS CHINENSIS ROOT EXTRACT|RHUS CHINENSIS ROOT EXTRACT
C3538619|T121|1373161|RXNORM|SCROPHULARIA NODOSA ROOT EXTRACT|SCROPHULARIA NODOSA ROOT EXTRACT
C0771655|T121|236388|RXNORM|LEVOMENTHOL|LEVOMENTHOL
C0073085|T121|35382|RXNORM|RESORCINOL|RESORCINOL
C0028741|T195|7597|RXNORM|NYSTATIN|NYSTATIN
C0028741|T195|7597|RXNORM|NYSTATIN|NYSTATIN
C0028741|T195|7597|RXNORM|NYSTATIN|NYSTATIN
C0028741|T195|7597|RXNORM|NYSTATIN|NYSTATIN
C0040898|T131|1000581|RXNORM|TRICHLORFON|TRICHLORFON
C2356025|T121|802573|RXNORM|DEXTROMETHORPHAN / PSEUDOEPHEDRINE / PYRILAMINE|DEXTROMETHORPHAN / PSEUDOEPHEDRINE / PYRILAMINE
C1698003|T121|615170|RXNORM|ACETAMINOPHEN / CAFFEINE / PHENYLTOLOXAMINE|ACETAMINOPHEN / CAFFEINE / PHENYLTOLOXAMINE
C0037355|T129|9835|RXNORM|SMALLPOX VACCINE|SMALLPOX VACCINE
C2928794|T121|1251752|RXNORM|LINSEED OIL / SOY PROTEIN ISOLATE|LINSEED OIL / SOY PROTEIN ISOLATE
C2725898|T129|882488|RXNORM|VENISON ALLERGENIC EXTRACT|VENISON ALLERGENIC EXTRACT
C2725897|T129|882485|RXNORM|GOOSE ALLERGENIC EXTRACT|ANSER ANSER ALLERGENIC EXTRACT
C0018959|T123|5164|RXNORM|HEMATOPORPHYRIN|HEMATOPORPHYRIN
C0911837|T109|1426443|RXNORM|CALCIUM PEROXIDE|CALCIUM PEROXIDE
C2111788|T121|815308|RXNORM|POLYETHYLENE GLYCOL 3350 / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE|POLYETHYLENE GLYCOL 3350 / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE
C2111788|T121|815308|RXNORM|POLYETHYLENE GLYCOL 3350 / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE|POLYETHYLENE GLYCOL 3350 / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE
C2168871|T121|813223|RXNORM|PHENYLPROPANOLAMINE / PYRILAMINE|PHENYLPROPANOLAMINE / PYRILAMINE
C1875994|T109|692620|RXNORM|GADOBENATE|GADOBENATE
C3535659|T121|1369687|RXNORM|PETASITES HYBRIDUS LEAF EXTRACT|PETASITES HYBRIDUS LEAF EXTRACT
C3645181|T121|1426831|RXNORM|TRIMETHYLPENTANEDIOL-ADIPIC ACID-GLYCERIN CROSSPOLYMER (25000 MPA.S)|TRIMETHYLPENTANEDIOL-ADIPIC ACID-GLYCERIN CROSSPOLYMER (25000 MPA.S)
C3535658|T121|1369688|RXNORM|PROPYLENE GLYCOL DIOLEATE|PROPYLENE GLYCOL DIOLEATE
C3833343|T121|1541212|RXNORM|CHLORHEXIDINE / HYDROCORTISONE|CHLORHEXIDINE / HYDROCORTISONE
C0060156|T121|24830|RXNORM|FENBUFEN|FENBUFEN
C3486615|T121|1333265|RXNORM|CHELONE GLABRA EXTRACT|CHELONE GLABRA EXTRACT
C3486531|T121|1307848|RXNORM|OPUNTIA FICUS-INDICA FLOWER EXTRACT|OPUNTIA FICUS-INDICA FLOWER EXTRACT
C3488375|T121|1333267|RXNORM|LEMNA MINOR EXTRACT|LEMNA MINOR EXTRACT
C0015039|T121|4132|RXNORM|ETHOGLUCID|ETHOGLUCID
C3256670|T121|1307849|RXNORM|CAMELLIA OLEIFERA SEED EXTRACT|CAMELLIA OLEIFERA SEED EXTRACT
C0015042|T121|4134|RXNORM|PROFENAMINE|PROFENAMINE
C0015043|T121|4135|RXNORM|ETHOSUXIMIDE|ETHOSUXIMIDE
C0015046|T121|4136|RXNORM|ETHOTOIN|ETHOTOIN
C3256857|T121|1307846|RXNORM|LEVANT COTTON SEED EXTRACT|LEVANT COTTON SEED EXTRACT
C0020933|T195|5690|RXNORM|IMIPENEM|IMIPENEM
C0020934|T121|5691|RXNORM|IMIPRAMINE|IMIPRAMINE
C2193964|T121|815166|RXNORM|DEXTROMETHORPHAN / DOXYLAMINE|DEXTROMETHORPHAN / DOXYLAMINE
C3255694|T109|1307847|RXNORM|LIPPIA CITRIODORA FLOWERING TOP OIL|LIPPIA CITRIODORA FLOWERING TOP OIL
C0729681|T007|1544931|RXNORM|BARTONELLA CLARRIDGEIAE|BARTONELLA CLARRIDGEIAE
C0318324|T007|1544930|RXNORM|BARTONELLA BACILLIFORMIS|BARTONELLA BACILLIFORMIS
C0242631|T007|1544933|RXNORM|BARTONELLA HENSELAE|BARTONELLA HENSELAE
C3819178|T121|1494040|RXNORM|BENZALKONIUM / N-ALKYL ETHYLBENZYL DIMETHYL AMMONIUM (C12-C14)|BENZALKONIUM / N-ALKYL ETHYLBENZYL DIMETHYL AMMONIUM (C12-C14)
C3714984|T007|1544935|RXNORM|BARTONELLA VINSONII|BARTONELLA VINSONII
C0035791|T007|1544934|RXNORM|BARTONELLA QUINTANA|BARTONELLA QUINTANA
C0315218|T007|1544937|RXNORM|CITROBACTER KOSERI|CITROBACTER KOSERI
C2940176|T129|1014721|RXNORM|CALIFORNIA BLACK OAK POLLEN EXTRACT|QUERCUS KELLOGGII POLLEN EXTRACT
C2073868|T121|818496|RXNORM|ASPIRIN / CHLORPHENIRAMINE / PHENYLEPHRINE|ASPIRIN / CHLORPHENIRAMINE / PHENYLEPHRINE
C3488968|T121|1309428|RXNORM|GENTIANELLA AMARELLA FLOWER EXTRACT|GENTIANELLA AMARELLA FLOWER EXTRACT
C1177017|T121|358871|RXNORM|DEXTRAN 110|DEXTRAN 110
C0142046|T121|56188|RXNORM|SERMORELIN|SERMORELIN
C0142046|T121|56188|RXNORM|SERMORELIN|SERMORELIN
C0936148|T121|282446|RXNORM|POSACONAZOLE|POSACONAZOLE
C3474132|T121|1313240|RXNORM|ISOCETYL STEARATE|ISOCETYL STEARATE
C3475291|T109|1313243|RXNORM|MANGANESE VIOLET|MANGANESE VIOLET
C3153428|T121|1313242|RXNORM|LIQUIDAMBAR STYRACIFLUA RESIN|LIQUIDAMBAR STYRACIFLUA RESIN
C2825460|T121|1313245|RXNORM|METYRAPONE TARTRATE|METYRAPONE TARTRATE
C3464711|T121|1313244|RXNORM|METHYLSERINE|METHYLSERINE
C3465035|T121|1313247|RXNORM|MYRISTYL PROPIONATE|MYRISTYL PROPIONATE
C3256376|T109|1313246|RXNORM|MYRISTYL GLUCOSIDE|MYRISTYL GLUCOSIDE
C3256716|T121|1313249|RXNORM|POVIDONE K17|POVIDONE K17
C0046596|T131|1313248|RXNORM|O-XYLENE|O-XYLENE
C0982298|T121|1426398|RXNORM|OCTOXYNOL-5|OCTOXYNOL-5
C2744960|T121|1364449|RXNORM|CROFELEMER|CROFELEMER
C0936150|T121|282448|RXNORM|ARTEMETHER / LUMEFANTRINE|ARTEMETHER / LUMEFANTRINE
C3256036|T121|1313741|RXNORM|DIGLYCERIN|DIGLYCERIN
C1618782|T121|578635|RXNORM|CEREBRAL PHOSPHOLIPIDS|CEREBRAL PHOSPHOLIPIDS
C2929025|T121|1008118|RXNORM|BISACODYL / SIMETHICONE|BISACODYL / SIMETHICONE
C2929026|T121|1008119|RXNORM|CAPSAICIN / MENTHOL / METHYLNICOTINATE|CAPSAICIN / MENTHOL / METHYLNICOTINATE
C2929021|T121|1008114|RXNORM|HYDROCORTISONE / PRAMOXINE / ZINC SULFATE|HYDROCORTISONE / PRAMOXINE / ZINC SULFATE
C2929022|T121|1008115|RXNORM|COPPER GLUCONATE / ZINC PICOLINATE|COPPER GLUCONATE / ZINC PICOLINATE
C2929023|T121|1008116|RXNORM|BROMAZEPAM / TRIMEBUTINE|BROMAZEPAM / TRIMEBUTINE
C2929024|T121|1008117|RXNORM|WITCH HAZEL / ZINC OXIDE|WITCH HAZEL / ZINC OXIDE
C2929018|T121|1008110|RXNORM|CODEINE / DICLOFENAC|CODEINE / DICLOFENAC
C2193836|T121|1008111|RXNORM|AMOXICILLIN / FLOXACILLIN|AMOXICILLIN / FLOXACILLIN
C2929019|T121|1008112|RXNORM|CYCLOADIPHENINE / PROPYPHENAZONE|CYCLOADIPHENINE / PROPYPHENAZONE
C2929020|T121|1008113|RXNORM|ANGELICA SINENSIS PREPARATION / SOY GERM|ANGELICA SINENSIS PREPARATION / SOY GERM
C0022029|T130|5968|RXNORM|IOPHENDYLATE|IOPHENDYLATE
C0077047|T109|38585|RXNORM|TRICHLOROTRIFLUOROETHANE|TRICHLOROTRIFLUOROETHANE
C0054084|T121|19727|RXNORM|BRODIMOPRIM|BRODIMOPRIM
C0054015|T125|19666|RXNORM|NESIRITIDE|NESIRITIDE
C0069454|T121|32385|RXNORM|OLSALAZINE|OLSALAZINE
C3255852|T109|1426329|RXNORM|MAGNESIUM ALUMINOMETASILICATE TYPE I-A|MAGNESIUM ALUMINOMETASILICATE TYPE I-A
C0022026|T130|5966|RXNORM|IOPAMIDOL|IOPAMIDOL
C0022028|T130|5967|RXNORM|IOPANOIC ACID|IOPANOIC ACID
C3255659|T109|1306184|RXNORM|CETYL PHOSPHATE|CETYL PHOSPHATE
C3255660|T109|1306185|RXNORM|CETYLHYDROXYPROLINE PALMITAMIDE|CETYLHYDROXYPROLINE PALMITAMIDE
C3255653|T109|1306180|RXNORM|CETYL MYRISTATE|CETYL MYRISTATE
C3255654|T109|1306181|RXNORM|CETYL OCTANOATE|CETYL CAPRYLATE
C3255655|T109|1306182|RXNORM|CETYL OLEATE|CETYL OLEATE
C3255656|T109|1306183|RXNORM|CETYL PALMITOLEATE|CETYL PALMITOLEATE
C3265016|T109|1368144|RXNORM|C30-45 OLEFIN|C30-45 OLEFIN
C0054416|T197|1368145|RXNORM|CADMIUM SULFATE|CADMIUM SULFATE
C3475108|T109|1368146|RXNORM|CAPRYLYL-CAPRYL OLIGOGLUCOSIDE|CAPRYLYL-CAPRYL OLIGOGLUCOSIDE
C0006937|T131|1368147|RXNORM|CAPTAN|CAPTAN
C3255707|T109|1306188|RXNORM|NEOPENTYL GLYCOL DIHEPTANOATE|NEOPENTYL GLYCOL DIHEPTANOATE
C3255730|T109|1306189|RXNORM|HORDEUM VULGARE ROOT EXTRACT|HORDEUM VULGARE ROOT EXTRACT
C3256510|T109|1368142|RXNORM|C10-30 CHOLESTEROL-LANOSTEROL ESTERS|C10-30 CHOLESTEROL-LANOSTEROL ESTERS
C3256511|T109|1368143|RXNORM|C12-16 ALCOHOLS|C12-16 ALCOHOLS
C0304119|T168|90950|RXNORM|THYME OIL|THYME OIL
C1720421|T121|644895|RXNORM|DIPHENHYDRAMINE / IBUPROFEN|DIPHENHYDRAMINE / IBUPROFEN
C0016296|T131|4460|RXNORM|FLUNITRAZEPAM|FLUNITRAZEPAM
C0650160|T130|183830|RXNORM|IOCETAMIC ACID|IOCETAMIC ACID
C1576812|T121|1363567|RXNORM|HYPROMELLOSE 2910|HYPROMELLOSE 2910
C3162750|T121|1114846|RXNORM|CHOLECALCIFEROL / CHONDROITIN SULFATES / GLUCOSAMINE|CHOLECALCIFEROL / CHONDROITIN SULFATES / GLUCOSAMINE
C1533480|T121|1363566|RXNORM|LAURETH-7|LAURETH-7
C3256897|T121|1307589|RXNORM|CASSIA FISTULA FRUIT EXTRACT|CASSIA FISTULA FRUIT EXTRACT
C0282849|T123|82242|RXNORM|CHLOROPHYLLIN COPPER COMPLEX|CHLOROPHYLLIN COPPER COMPLEX
C3464954|T121|1307587|RXNORM|WITHANIA SOMNIFERA LEAF EXTRACT|WITHANIA SOMNIFERA LEAF EXTRACT
C3485013|T121|1307586|RXNORM|PARIS POLYPHYLLA ROOT EXTRACT|PARIS POLYPHYLLA ROOT EXTRACT
C3256566|T121|1307585|RXNORM|THUJA OCCIDENTALIS BARK EXTRACT|THUJA OCCIDENTALIS BARK EXTRACT
C3255953|T121|1307582|RXNORM|MALVA SYLVESTRIS LEAF EXTRACT|HIGH MALLOW LEAF EXTRACT
C3255946|T121|1307581|RXNORM|MAGNOLIA GRANDIFLORA BARK EXTRACT|MAGNOLIA GRANDIFLORA BARK EXTRACT
C3256720|T121|1307580|RXNORM|SALVIA MILTIORRHIZA ROOT EXTRACT|SALVIA MILTIORRHIZA ROOT EXTRACT
C0009002|T121|2594|RXNORM|CLOFIBRATE|CLOFIBRATE
C0982363|T121|1314411|RXNORM|PROPYLENE GLYCOL STEARATE|PROPYLENE GLYCOL MONOSTEARATE
C0009008|T121|2596|RXNORM|CLOMIPHENE|CLOMIPHENE
C0009010|T121|2597|RXNORM|CLOMIPRAMINE|CLOMIPRAMINE
C0008992|T121|2590|RXNORM|CLOBETASOL|CLOBETASOL
C3555460|T121|1421148|RXNORM|BOS TAURUS DUODENUM PREPARATION|BOVINE DUODENUM PREPARATION
C0008996|T130|2592|RXNORM|CLOFAZIMINE|CLOFAZIMINE
C3486578|T121|1314410|RXNORM|GERMANIUM SESQUIOXIDE|GERMANIUM SESQUIOXIDE
C2918653|T121|1306235|RXNORM|EQUISETUM ARVENSE TOP EXTRACT|EQUISETUM ARVENSE TOP EXTRACT
C0009011|T121|2598|RXNORM|CLONAZEPAM|CLONAZEPAM
C0009014|T121|2599|RXNORM|CLONIDINE|CLONIDINE
C0009014|T121|2599|RXNORM|CLONIDINE|CLONIDINE
C0015540|T123|1314412|RXNORM|FLAVIN-ADENINE DINUCLEOTIDE|FLAVIN-ADENINE DINUCLEOTIDE
C0032393|T121|1314414|RXNORM|POLOXALENE|POLOXALENE
C2746811|T121|903986|RXNORM|HYOSCYAMINE / PHENYLTOLOXAMINE|HYOSCYAMINE / PHENYLTOLOXAMINE
C0284711|T109|1314417|RXNORM|TRIBUTYL CITRATE|TRIBUTYL CITRATE
C0982050|T130|1364944|RXNORM|CALDIAMIDE|CALDIAMIDE
C0724614|T121|1314416|RXNORM|LEVO-METHAMPHETAMINE|LEVOMETAMFETAMINE
C3833081|T109|1540357|RXNORM|PEANUT OIL, HYDROGENATED|PEANUT OIL, HYDROGENATED
C3556196|T121|1375947|RXNORM|DOXYLAMINE / PYRIDOXINE|DOXYLAMINE / PYRIDOXINE
C0520520|T121|1314419|RXNORM|TRICAPRIN|TRICAPRIN
C3282133|T121|1250666|RXNORM|ACYCLOVIR / LIDOCAINE|ACYCLOVIR / LIDOCAINE
C0077021|T121|1314418|RXNORM|TRIBUTYL PHOSPHATE|TRIBUTYL PHOSPHATE
C0022230|T121|6048|RXNORM|INOSINE PRANOBEX|INOSINE PRANOBEX
C2933878|T121|1364947|RXNORM|5-BROMO-5-NITRO-1,3-DIOXANE|5-BROMO-5-NITRO-1,3-DIOXANE
C1589658|T121|544983|RXNORM|PROVIDONE-IODINE|PROVIDONE-IODINE
C0026202|T195|6985|RXNORM|MIOCAMYCIN|MIOCAMYCIN
C0009073|T121|2622|RXNORM|CLOTIAZEPAM|CLOTIAZEPAM
C0009074|T121|2623|RXNORM|CLOTRIMAZOLE|CLOTRIMAZOLE
C0009074|T121|2623|RXNORM|CLOTRIMAZOLE|CLOTRIMAZOLE
C0009074|T121|2623|RXNORM|CLOTRIMAZOLE|CLOTRIMAZOLE
C0009071|T121|2620|RXNORM|CLOTHIAPINE|CLOTHIAPINE
C0026196|T121|6984|RXNORM|MINOXIDIL|MINOXIDIL
C0026196|T121|6984|RXNORM|MINOXIDIL|MINOXIDIL
C0009079|T121|2626|RXNORM|CLOZAPINE|CLOZAPINE
C0009077|T195|2625|RXNORM|CLOXACILLIN|CLOXACILLIN
C2364500|T129|805471|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED, INFLUENZA B (B-FLORIDA-4-2006) STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED, INFLUENZA B (B-FLORIDA-4-2006) STRAIN
C2726999|T129|974140|RXNORM|ENGLISH SOLE ALLERGENIC EXTRACT|PAROPHRYS VETULUS ALLERGENIC EXTRACT
C3486675|T121|1313692|RXNORM|RED PEPPER EXTRACT|RED PEPPER EXTRACT
C0038071|T130|10014|RXNORM|SQUALENE|SQUALENE
C1713670|T121|636648|RXNORM|POTASSIUM BITARTRATE / SODIUM BICARBONATE|POTASSIUM BITARTRATE / SODIUM BICARBONATE
C3535851|T121|1370639|RXNORM|LAURYL SARCOSINATE|LAURYL SARCOSINATE
C3535852|T122|1370638|RXNORM|OLEANOLATE|OLEANOLATE
C3535853|T121|1370637|RXNORM|STARCH GLYCOLATE|STARCH GLYCOLATE
C3535854|T121|1370636|RXNORM|STARCH GLYCOLATE TYPE A POTATO|STARCH GLYCOLATE TYPE A POTATO
C3535855|T130|1370635|RXNORM|DEHYDROACETATE|DEHYDROACETATE
C3535856|T121|1370634|RXNORM|CUMENESULFONATE|CUMENESULFONATE
C2726191|T129|972365|RXNORM|PENICILLIUM ROQUEFORTII ALLERGENIC EXTRACT|PENICILLIUM ROQUEFORTII ALLERGENIC EXTRACT
C3535857|T121|1370631|RXNORM|COCOYL GLUTAMATE|COCOYL GLUTAMATE
C3535858|T109|1370630|RXNORM|AZELOYL DIGLYCINATE|AZELOYL DIGLYCINATE
C1874385|T121|689595|RXNORM|ATROPINE / CHLORPHENIRAMINE|ATROPINE / CHLORPHENIRAMINE
C0771584|T121|236324|RXNORM|MAGNESIUM GLUTAMATE|MAGNESIUM GLUTAMATE
C0763530|T121|232539|RXNORM|CALFACTANT|CALFACTANT
C2740713|T129|899576|RXNORM|PAPER BIRCH POLLEN EXTRACT|BETULA PAPYRIFERA POLLEN EXTRACT
C2726188|T129|883442|RXNORM|PASSALORA FULVA EXTRACT|PASSALORA FULVA EXTRACT
C3255762|T109|1313698|RXNORM|ETHYLCELLULOSE (4 MPA.S)|ETHYLCELLULOSE (4 MPA.S)
C2193874|T121|820916|RXNORM|MEBENDAZOLE / TINIDAZOLE|MEBENDAZOLE / TINIDAZOLE
C3537532|T109|1370989|RXNORM|MORUS ALBA EXTRACT|MORUS ALBA EXTRACT
C3537531|T121|1370988|RXNORM|TRIBULUS TERRESTRIS EXTRACT|TRIBULUS TERRESTRIS EXTRACT
C0070570|T121|33290|RXNORM|PHENOL|PHENOL
C0070570|T121|33290|RXNORM|PHENOL|PHENOL
C0070570|T121|33290|RXNORM|PHENOL|PHENOL
C0070570|T121|33290|RXNORM|PHENOL|PHENOL
C0070570|T121|33290|RXNORM|PHENOL|PHENOL
C0070570|T121|33290|RXNORM|PHENOL|PHENOL
C2014103|T121|814872|RXNORM|ACETAMINOPHEN / ORPHENADRINE|ACETAMINOPHEN / ORPHENADRINE
C3537526|T121|1370983|RXNORM|CHONDROITIN SULFATE (CHICKEN)|CHONDROITIN SULFATE (CHICKEN)
C2702402|T129|892499|RXNORM|TOMATO ALLERGENIC EXTRACT|TOMATO ALLERGENIC EXTRACT
C3537528|T121|1370985|RXNORM|TRAMETES VERSICOLOR FRUITING BODY EXTRACT|TRAMETES VERSICOLOR FRUITING BODY EXTRACT
C3537527|T121|1370984|RXNORM|LAGERSTROEMIA INDICA EXTRACT|LAGERSTROEMIA INDICA EXTRACT
C3537530|T109|1370987|RXNORM|MICROCITRUS AUSTRALIS FRUIT EXTRACT|MICROCITRUS AUSTRALIS FRUIT EXTRACT
C3500499|T121|1314665|RXNORM|ASCORBIC ACID / BIOTIN / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACIN / PANTOTHENATE / POLYSACCHARIDE IRON COMPLEX / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC SULFATE|ASCORBIC ACID / BIOTIN / COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACIN / PANTOTHENATE / POLYSACCHARIDE IRON COMPLEX / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC SULFATE
C0055014|T195|20492|RXNORM|CEFTIBUTEN|CEFTIBUTEN
C0057831|T121|22892|RXNORM|DICHLORALPHENAZONE|DICHLORALPHENAZONE
C0210630|T129|68442|RXNORM|FILGRASTIM|FILGRASTIM
C0055021|T121|20498|RXNORM|CELIPROLOL|CELIPROLOL
C0210657|T121|68446|RXNORM|PEMETREXED|PEMETREXED
C0064909|T125|1546435|RXNORM|SALMON GONADOTROPIN RELEASING HORMONE D-ARG6 ANALOG ETHYL AMIDE|SALMON GONADOTROPIN RELEASING HORMONE D-ARG6 ANALOG ETHYL AMIDE
C1166209|T121|350489|RXNORM|VISCUM ALBUM PREPARATION|VISCUM ALBUM PREPARATION
C0972314|T121|307296|RXNORM|ETORICOXIB|ETORICOXIB
C2929363|T121|1008459|RXNORM|ALPHA-D-GALACTOSIDASE ENZYME / BROMELAINS / PAPAIN|ALPHA-D-GALACTOSIDASE ENZYME / BROMELAINS / PAPAIN
C0062587|T195|26797|RXNORM|HETACILLIN|HETACILLIN
C0002823|T126|772|RXNORM|ANCROD|ANCROD
C0054560|T109|20129|RXNORM|CAMPESTEROL|CAMPESTEROL
C2726178|T129|1006510|RXNORM|BARLEY MALT ALLERGENIC EXTRACT|BARLEY MALT ALLERGENIC EXTRACT
C0000473|T127|74|RXNORM|4-AMINOBENZOIC ACID|AMINOBENZOIC ACID
C0000473|T127|74|RXNORM|4-AMINOBENZOIC ACID|AMINOBENZOIC ACID
C0000464|T123|73|RXNORM|DOCOSAHEXAENOATE|DOCOSAHEXAENOATE
C3540675|T109|1421644|RXNORM|BITTER ALMOND EXTRACT|BITTER ALMOND EXTRACT
C0010525|T121|2970|RXNORM|CYCLANDELATE|CYCLANDELATE
C0010547|T121|2977|RXNORM|CYCLIZINE|CYCLIZINE
C2740617|T129|899414|RXNORM|GARLIC ALLERGENIC EXTRACT|ALLIUM SATIVUM ALLERGENIC EXTRACT
C0003596|T121|1043|RXNORM|APOMORPHINE|APOMORPHINE
C0003596|T121|1043|RXNORM|APOMORPHINE|APOMORPHINE
C0019654|T129|5363|RXNORM|HISTOPLASMIN|HISTOPLASMIN
C0795635|T125|253182|RXNORM|REGULAR INSULIN, HUMAN|INSULIN (HUMAN)
C0109002|T121|47858|RXNORM|METHSUXIMIDE|MESUXIMIDE
C0051395|T121|17511|RXNORM|ALPHA-KETOGLUTARIC ACID|ALPHA-KETOGLUTARIC ACID
C0010560|T125|2983|RXNORM|CYCLOFENIL|CYCLOFENIL
C2709776|T129|854972|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 9N VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 9N VACCINE
C0066677|T121|30125|RXNORM|MODAFINIL|MODAFINIL
C2731373|T129|895062|RXNORM|HAMSTER SKIN EXTRACT|HAMSTER SKIN EXTRACT
C0005100|T121|1426|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, B-WISCONSIN-1-2010 STRAIN|BENZYL ALCOHOL
C0015689|T123|4301|RXNORM|OMEGA-3 FATTY ACIDS|OMEGA-3 FATTY ACIDS
C1667052|T121|620216|RXNORM|MARAVIROC|MARAVIROC
C2701580|T129|966925|RXNORM|COTTON FIBER ALLERGENIC EXTRACT|COTTON FIBER ALLERGENIC EXTRACT
C2740637|T129|899444|RXNORM|LENTIL ALLERGENIC EXTRACT|LENTIL ALLERGENIC EXTRACT
C0071214|T123|33835|RXNORM|PLASMA PROTEIN FRACTION|PLASMA PROTEIN FRACTION
C2929195|T121|1008288|RXNORM|BELLADONNA EXTRACT, USP / OPIUM|BELLADONNA EXTRACT, USP / OPIUM
C0042071|T126|11055|RXNORM|UROKINASE|UROKINASE
C3500826|T121|1356126|RXNORM|BRYONIA ALBA WHOLE EXTRACT|BRYONIA ALBA WHOLE EXTRACT
C2929192|T121|1008285|RXNORM|GLYCERIN / HYPROMELLOSE / PROPYLENE GLYCOL|GLYCERIN / HYPROMELLOSE / PROPYLENE GLYCOL
C2929193|T121|1008286|RXNORM|GLYCERIN / PHENOL|GLYCERIN / PHENOL
C2929194|T121|1008287|RXNORM|BELLADONNA EXTRACT, USP / CHARCOAL|BELLADONNA EXTRACT, USP / CHARCOAL
C2929188|T121|1008281|RXNORM|CHENODEOXYCHOLATE / URSODEOXYCHOLATE|CHENODEOXYCHOLATE / URSODEOXYCHOLATE
C2929189|T121|1008282|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / FOLIC ACID / PHYTOSTEROLS / VITAMIN B 12 / VITAMIN B6|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / FOLIC ACID / PHYTOSTEROLS / VITAMIN B 12 / VITAMIN B6
C2929190|T121|1008283|RXNORM|CALCIUM CHLORIDE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE|CALCIUM CHLORIDE / LACTATE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM ACETATE / SODIUM CHLORIDE
C0011134|T131|3129|RXNORM|DEET|DIETHYLTOLUAMIDE
C0002158|T125|525|RXNORM|ALLYLESTRENOL|ALLYLESTRENOL
C3696418|T121|1484957|RXNORM|FACTOR IX / FACTOR VII / FACTOR X / PROTEIN C / PROTHROMBIN / VITAMIN K-DEPENDENT PROTEIN S|FACTOR IX / FACTOR VII / FACTOR X / PROTEIN C / PROTEIN S / PROTHROMBIN
C0061932|T121|26290|RXNORM|GUAIAZULENE|GUAIAZULENE
C0939899|T121|285245|RXNORM|CINNAMON PREPARATION|CINNAMON PREPARATION
C0937604|T121|283545|RXNORM|BUSHMASTER VENOM|BUSHMASTER VENOM
C0049506|T121|15996|RXNORM|MIRTAZAPINE|MIRTAZAPINE
C0937598|T168|283540|RXNORM|APPLE PECTIN|APPLE PECTIN
C0937599|T121|283541|RXNORM|BARLEY GRAIN|BARLEY GRAIN
C0205705|T121|66870|RXNORM|CASANTHRANOL|CASANTHRANOL
C0068377|T121|31479|RXNORM|NALMEFENE|NALMEFENE
C0068366|T121|31475|RXNORM|NAFTAZONE|NAFTAZONE
C0068367|T121|31476|RXNORM|NAFTIFINE|NAFTIFINE
C3535666|T121|1369396|RXNORM|TROPAEOLUM MAJUS FLOWER EXTRACT|TROPAEOLUM MAJUS FLOWER EXTRACT
C0815310|T121|258439|RXNORM|HEAVY MINERAL OIL|HEAVY MINERAL OIL
C3535667|T121|1369395|RXNORM|APPLE SEED EXTRACT|APPLE SEED EXTRACT
C3489340|T121|1311658|RXNORM|POMEGRANATE FRUIT RIND EXTRACT|POMEGRANATE FRUIT RIND EXTRACT
C3488117|T121|1311659|RXNORM|PROPOLIS WAX|BEE PROPOLIS EXTACT
C3256734|T109|1311650|RXNORM|ULTRAMARINE BLUE|ULTRAMARINE BLUE
C3255962|T121|1311651|RXNORM|PASSIFLORA INCARNATA FRUIT EXTRACT|PASSIFLORA INCARNATA FRUIT EXTRACT
C3488939|T121|1311653|RXNORM|PERILLA FRUTESCENS FRUIT EXTRACT|PERILLA FRUTESCENS FRUIT EXTRACT
C3256426|T121|1311654|RXNORM|PHYLLANTHUS EMBLICA FRUIT EXTRACT|PHYLLANTHUS EMBLICA FRUIT EXTRACT
C3474469|T121|1311655|RXNORM|HYDROLYZED PLACENTAL PROTEIN (BOVINE)|HYDROLYZED PLACENTAL PROTEIN (BOVINE)
C3488953|T121|1311656|RXNORM|PHYLLANTHUS NIRURI TOP EXTRACT|PHYLLANTHUS NIRURI TOP EXTRACT
C2928557|T121|1007641|RXNORM|CAMPHOR / EUCALYPTUS OIL / MENTHOL / TURPENTINE|CAMPHOR / EUCALYPTUS OIL / MENTHOL / TURPENTINE
C2928556|T121|1007640|RXNORM|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G1 VACCINE / HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G2 VACCINE / HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G3 VACCINE / HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G4 VACCINE / HUMAN-BOVINE REASSORTANT ROTAVIRUS|HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G1 VACCINE / HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G2 VACCINE / HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G3 VACCINE / HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN G4 VACCINE / HUMAN-BOVINE REASSORTANT ROTAVIRUS STRAIN P1A[8] VACCINE
C3505266|T121|1358175|RXNORM|LEVULINATE|LEVULINATE
C2928561|T121|1007645|RXNORM|CALCIUM CHLORIDE / FIBRINOGEN / FIBRINOLYSIS INHIBITOR / THROMBIN|CALCIUM CHLORIDE / FIBRINOGEN / FIBRINOLYSIS INHIBITOR / THROMBIN
C2928560|T121|1007644|RXNORM|BELLADONNA ALKALOIDS / CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE|BELLADONNA ALKALOIDS / CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLPROPANOLAMINE
C2928562|T121|1007646|RXNORM|PHENYLEPHRINE / TRIPROLIDINE|PHENYLEPHRINE / TRIPROLIDINE
C2928565|T121|1007649|RXNORM|HYOSCYAMUS EXTRACT / PHENOBARBITAL|HYOSCYAMUS EXTRACT / PHENOBARBITAL
C2928564|T121|1007648|RXNORM|MANNITOL / PHENOBARBITAL|MANNITOL / PHENOBARBITAL
C0305048|T129|91596|RXNORM|POLYVALENT CROTALIDAE ANTIVENIN|POLYVALENT CROTALIDAE ANTIVENIN
C0530684|T121|1112990|RXNORM|EZOGABINE|RETIGABINE
C1961993|T121|725206|RXNORM|POMEGRANATE EXTRACT|POMEGRANATE EXTRACT
C1875118|T121|691245|RXNORM|EPINEPHRINE / PILOCARPINE|EPINEPHRINE / PILOCARPINE
C1875119|T121|691247|RXNORM|EPINEPHRINE / ZINC CHLORIDE|EPINEPHRINE / ZINC CHLORIDE
C2183347|T121|819516|RXNORM|ACETAMINOPHEN / DICLOFENAC|ACETAMINOPHEN / DICLOFENAC
C3265062|T121|1244014|RXNORM|VITAMIN D3|VITAMIN D3
C1364955|T121|435657|RXNORM|OLIVE LEAF EXTRACT|OLIVE LEAF EXTRACT
C1142738|T121|341018|RXNORM|ANIDULAFUNGIN|ANIDULAFUNGIN
C2194156|T121|817455|RXNORM|ASCORBIC ACID / ASPIRIN / CAFFEINE|ASCORBIC ACID / ASPIRIN / CAFFEINE
C1608295|T121|592464|RXNORM|ARTICAINE|ARTICAINE
C0076890|T121|38453|RXNORM|TRAMAZOLINE|TRAMAZOLINE
C3818717|T121|1535477|RXNORM|CYMBOPOGON MARTINI WHOLE EXTRACT|CYMBOPOGON MARTINI WHOLE EXTRACT
C3819173|T121|1534845|RXNORM|KETOCONAZOLE / PHYTOSPHINGOSINE|KETOCONAZOLE / PHYTOSPHINGOSINE
C0717685|T121|214485|RXNORM|DEXTRAN 1|DEXTRAN 1
C0048504|T121|15226|RXNORM|FOMEPIZOLE|FOMEPIZOLE
C0717690|T121|214489|RXNORM|DEXTROMETHORPHAN / PHENYLPROPANOLAMINE|DEXTROMETHORPHAN / PHENYLPROPANOLAMINE
C0717689|T121|214488|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN|DEXTROMETHORPHAN / GUAIFENESIN
C0717689|T121|214488|RXNORM|DEXTROMETHORPHAN / GUAIFENESIN|DEXTROMETHORPHAN / GUAIFENESIN
C0028116|T121|7435|RXNORM|NISOLDIPINE|NISOLDIPINE
C2075282|T121|813013|RXNORM|ANISE OIL / CITRIC ACID|ANISE OIL / CITRIC ACID
C2928788|T121|1007874|RXNORM|FOLIC ACID / LIVER EXTRACT / VITAMIN B 12|FOLIC ACID / LIVER EXTRACT / VITAMIN B 12
C3848615|T109|1544273|RXNORM|OCIMUM AFRICANUM LEAF EXTRACT|OCIMUM AFRICANUM LEAF EXTRACT
C2930043|T121|1009150|RXNORM|DEXAMETHASONE / SODIUM PHOSPHATE|DEXAMETHASONE / SODIUM PHOSPHATE
C0016865|T121|4604|RXNORM|FURSULTIAMIN|FURSULTIAMIN
C3500586|T121|1314843|RXNORM|CAPSICUM ANNUUM WHOLE EXTRACT|CAPSICUM ANNUUM WHOLE EXTRACT
C0025033|T131|6674|RXNORM|MECHLORETHAMINE|MECHLORETHAMINE
C0025033|T131|6674|RXNORM|MECHLORETHAMINE|MECHLORETHAMINE
C0025039|T121|6676|RXNORM|MECLIZINE|MECLIZINE
C3818751|T121|1493693|RXNORM|GYMNEMA SYLVESTRE LEAF EXTRACT|GYMNEMA SYLVESTRE LEAF EXTRACT
C3812144|T121|1493692|RXNORM|GELSEMIUM SEMPERVIRENS WHOLE EXTRACT|GELSEMIUM SEMPERVIRENS WHOLE EXTRACT
C0025029|T121|6673|RXNORM|MECAMYLAMINE|MECAMYLAMINE
C0025023|T121|6672|RXNORM|MEBENDAZOLE|MEBENDAZOLE
C3488430|T121|1330093|RXNORM|PACKERA AUREA EXTRACT|PACKERA AUREA EXTRACT
C3488254|T121|1330092|RXNORM|CIMEX LECTULARIUS PREPARATION|CIMEX LECTULARIUS PREPARATION
C3486811|T121|1330091|RXNORM|SEDUM ACRE EXTRACT|SEDUM ACRE EXTRACT
C3486810|T121|1330090|RXNORM|SCROPHULARIA NODOSA EXTRACT|SCROPHULARIA NODOSA EXTRACT
C2928463|T121|1007542|RXNORM|ERGOLOID MESYLATES, USP / NIFEDIPINE|ERGOLOID MESYLATES, USP / NIFEDIPINE
C0142915|T121|56512|RXNORM|SODIUM POLYSTYRENE SULFONATE|SODIUM POLYSTYRENE SULFONATE
C2928464|T121|1007543|RXNORM|GLYCERIN / PRAMOXINE|GLYCERIN / PRAMOXINE
C2727930|T129|889669|RXNORM|SMELT ALLERGENIC EXTRACT|SMELT ALLERGENIC EXTRACT
C2928461|T121|1007540|RXNORM|GLYCERIN / NAPHAZOLINE / ZINC SULFATE|GLYCERIN / NAPHAZOLINE / ZINC SULFATE
C1873948|T121|689558|RXNORM|ACETAMINOPHEN / BROMPHENIRAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / BROMPHENIRAMINE / PSEUDOEPHEDRINE
C2928159|T121|1007237|RXNORM|ANTIPYRINE / CAFFEINE|ANTIPYRINE / CAFFEINE
C0120107|T121|50610|RXNORM|GOSERELIN|GOSERELIN
C1873941|T121|689551|RXNORM|ACETAMINOPHEN / ASPIRIN / CAFFEINE / CALCIUM GLUCONATE|ACETAMINOPHEN / ASPIRIN / CAFFEINE / CALCIUM GLUCONATE
C2928152|T121|1007230|RXNORM|BROMHEXINE / SULFADIAZINE / TETROXOPRIM|BROMHEXINE / SULFADIAZINE / TETROXOPRIM
C1873943|T121|689553|RXNORM|ACETAMINOPHEN / ASPIRIN / CAFFEINE / HYDROCODONE|ACETAMINOPHEN / ASPIRIN / CAFFEINE / HYDROCODONE
C1873942|T121|689552|RXNORM|ACETAMINOPHEN / ASPIRIN / CAFFEINE / CODEINE / SALICYLAMIDE|ACETAMINOPHEN / ASPIRIN / CAFFEINE / CODEINE / SALICYLAMIDE
C1873945|T121|689555|RXNORM|ACETAMINOPHEN / ASPIRIN / CODEINE|ACETAMINOPHEN / ASPIRIN / CODEINE
C1873944|T121|689554|RXNORM|ACETAMINOPHEN / ASPIRIN / CAFFEINE / SALICYLAMIDE|ACETAMINOPHEN / ASPIRIN / CAFFEINE / SALICYLAMIDE
C1873947|T121|689557|RXNORM|ACETAMINOPHEN / ATROPINE / ETHAVERINE / SALICYLAMIDE|ACETAMINOPHEN / ATROPINE / ETHAVERINE / SALICYLAMIDE
C0041175|T121|10865|RXNORM|TROMETHAMINE|TROMETHAMINE
C0054222|T121|19850|RXNORM|BUNAZOSIN|BUNAZOSIN
C3488976|T121|1441658|RXNORM|SENNA OCCIDENTALIS EXTRACT|SENNA OCCIDENTALIS EXTRACT
C0657912|T121|187832|RXNORM|PREGABALIN|PREGABALIN
C2928154|T121|1007232|RXNORM|ALVERINE / SIMETHICONE|ALVERINE / SIMETHICONE
C2928155|T121|1007233|RXNORM|BUTAMBEN / TYROTHRICIN|BUTAMBEN / TYROTHRICIN
C0771669|T121|236401|RXNORM|MEGLUMINE BENZOATE|MEGLUMINE BENZOATE
C0717408|T121|214220|RXNORM|AMITRIPTYLINE / CHLORDIAZEPOXIDE|AMITRIPTYLINE / CHLORDIAZEPOXIDE
C0717411|T121|214223|RXNORM|AMLODIPINE / BENAZEPRIL|AMLODIPINE / BENAZEPRIL
C0015888|T121|4356|RXNORM|FERROUS ASCORBATE|FERROUS ASCORBATE
C2701741|T129|852693|RXNORM|HOUSE MOUSE SKIN EXTRACT|MUS MUSCULUS SKIN EXTRACT
C0063912|T121|27866|RXNORM|ISOAMINILE|ISOAMINILE
C2701745|T130|852697|RXNORM|CANARY GRASS POLLEN EXTRACT|PHALARIS ARUNDINACEA POLLEN EXTRACT
C3854861|T121|1546708|RXNORM|DISTEARETH-75 ISOPHORONE DIISOCYANATE|DISTEARETH-75 ISOPHORONE DIISOCYANATE
C0209137|T121|1546358|RXNORM|MOEXIPRILAT|MOEXIPRILAT
C0039947|T195|1365970|RXNORM|THIOSTREPTON|THIOSTREPTON
C1095913|T121|319834|RXNORM|ELDERBERRY PREPARATION|ELDERBERRY PREPARATION
C2006143|T121|821278|RXNORM|CALCIUM LACTATE / NIACIN|CALCIUM LACTATE / NIACIN
C3848561|T196|1546357|RXNORM|FERRIC CATION|FERRIC CATION
C2080478|T121|817911|RXNORM|ACETAMINOPHEN / CAFFEINE / PHENYLEPHRINE|ACETAMINOPHEN / CAFFEINE / PHENYLEPHRINE
C0299583|T125|1441651|RXNORM|LEPTIN|LEPTIN
C1628973|T121|608424|RXNORM|HYDRALAZINE / ISOSORBIDE DINITRATE|HYDRALAZINE / ISOSORBIDE DINITRATE
C0056739|T121|21954|RXNORM|CYCLOBUTYROL|CYCLOBUTYROL
C0206008|T121|1546354|RXNORM|2-MERCAPTOETHANESULFONIC ACID|2-MERCAPTOETHANESULFONIC ACID
C0055869|T121|21224|RXNORM|CLEBOPRIDE|CLEBOPRIDE
C0055871|T195|21226|RXNORM|CLEMIZOLPENICILLIN|CLEMIZOLPENICILLIN
C3667093|T130|1438510|RXNORM|PIGMENT YELLOW 138|PIGMENT YELLOW 138
C2740600|T129|899382|RXNORM|BLUEBERRY ALLERGENIC EXTRACT|BLUEBERRY ALLERGENIC EXTRACT
C2740603|T129|899386|RXNORM|BROCCOLI ALLERGENIC EXTRACT|BRASSICA BOTRYTIS ALLERGENIC EXTRACT
C3488989|T121|1441655|RXNORM|CERVUS ELAPHUS VELVET PREPARATION|CERVUS ELAPHUS VELVET PREPARATION
C3696061|T121|1484904|RXNORM|SAFFRON EXTRACT|SAFFRON EXTRACT
C2928785|T121|1007871|RXNORM|CHLORAMPHENICOL / NAPHAZOLINE|CHLORAMPHENICOL / NAPHAZOLINE
C3536903|T204|1441656|RXNORM|TRICHOMONAS VAGINALIS PREPARATION|TRICHOMONAS VAGINALIS PREPARATION
C3488945|T121|1441657|RXNORM|MIRABILIS JALAPA TOP EXTRACT|MIRABILIS JALAPA TOP EXTRACT
C2168866|T121|1241828|RXNORM|ACETAMINOPHEN / PHENYLEPHRINE / PYRILAMINE|ACETAMINOPHEN / PHENYLEPHRINE / PYRILAMINE
C3856260|T121|1549874|RXNORM|MYRISTIC DIISOPROPANOLAMIDE|MYRISTIC DIISOPROPANOLAMIDE
C3256949|T109|1309248|RXNORM|SORBITAN OLIVATE|SORBITAN OLIVATE
C2949338|T121|1046414|RXNORM|CALCIUM GLYCEROPHOSPHATE / MONOFLUOROPHOSPHATE|CALCIUM GLYCEROPHOSPHATE / MONOFLUOROPHOSPHATE
C1725664|T121|644718|RXNORM|FERROUS ASPARTO GLYCINATE|FERROUS ASPARTO GLYCINATE
C0007248|T121|2101|RXNORM|CARISOPRODOL|CARISOPRODOL
C0007258|T121|2106|RXNORM|CARNITINE|CARNITINE
C0007257|T121|2105|RXNORM|CARMUSTINE|CARMUSTINE
C1874519|T121|690268|RXNORM|BENZOCAINE / ISOPROPYL ALCOHOL / MENTHOL|BENZOCAINE / ISOPROPYL ALCOHOL / MENTHOL
C2025210|T121|816583|RXNORM|ACETAMINOPHEN / CARISOPRODOL|ACETAMINOPHEN / CARISOPRODOL
C1453933|T121|474128|RXNORM|TELBIVUDINE|TELBIVUDINE
C0010240|T007|1432987|RXNORM|COXIELLA BURNETII|COXIELLA BURNETII
C1509448|T121|1367127|RXNORM|PEGOXOL 7 STEARATE|PEGOXOL 7 STEARATE
C1509397|T121|1367126|RXNORM|HEXYL LAURATE|HEXYL LAURATE
C1509343|T121|1367125|RXNORM|PEAR PREPARATION|PEAR PREPARATION
C1136869|T109|1367124|RXNORM|OCTYL DODECANOL|OCTYL DODECANOL
C3531533|T109|1367123|RXNORM|BACKHOUSIA CITRIODORA LEAF EXTRACT|BACKHOUSIA CITRIODORA LEAF EXTRACT
C0982418|T121|1367122|RXNORM|STEARETH-21|STEARETH-21
C0982417|T109|1367121|RXNORM|STEARETH-20|STEARETH-20
C0982310|T121|1367120|RXNORM|PEG-100 STEARATE|PEG-100 STEARATE
C3487986|T121|1309754|RXNORM|THUJA OCCIDENTALIS LEAFY TWIG EXTRACT|THUJA OCCIDENTALIS LEAFY TWIG EXTRACT
C3488684|T121|1309757|RXNORM|CEANOTHUS AMERICANUS LEAF EXTRACT|CEANOTHUS AMERICANUS LEAF EXTRACT
C3488434|T121|1309750|RXNORM|JUGLANS CINEREA BRANCH BARK-ROOT BARK EXTRACT|JUGLANS CINEREA BRANCH BARK-ROOT BARK EXTRACT
C3488908|T121|1309751|RXNORM|PUERARIA MONTANA VAR. LOBATA ROOT EXTRACT|PUERARIA MONTANA VAR. LOBATA ROOT EXTRACT
C3488435|T121|1309752|RXNORM|IRIS GERMANICA ROOT EXTRACT|IRIS GERMANICA ROOT EXTRACT
C3486575|T121|1309753|RXNORM|QUERCUS ROBUR FLOWER EXTRACT|QUERCUS ROBUR FLOWER EXTRACT
C3486576|T121|1309758|RXNORM|TOXICODENDRON RADICANS LEAF EXTRACT|TOXICODENDRON RADICANS LEAF EXTRACT
C3488685|T121|1309759|RXNORM|CHIONANTHUS VIRGINICUS BARK EXTRACT|CHIONANTHUS VIRGINICUS BARK EXTRACT
C1110634|T121|324036|RXNORM|PODOPHYLLUM PELTATUM PREPARATION|PODOPHYLLUM PELTATUM PREPARATION
C0770623|T121|235534|RXNORM|POLYOXYETHYLENE ETHER|POLYOXYETHYLENE ETHER
C1958569|T121|1091643|RXNORM|AZILSARTAN|AZILSARTAN
C0132512|T121|53692|RXNORM|NILVADIPINE|NILVADIPINE
C0132515|T121|53694|RXNORM|NIMESULIDE|NIMESULIDE
C0039902|T121|10485|RXNORM|THIOGUANINE|THIOGUANINE
C2168878|T121|820059|RXNORM|PYRVINIUM / THIABENDAZOLE|PYRVINIUM / THIABENDAZOLE
C0054207|T121|19836|RXNORM|BUFLOMEDIL|BUFLOMEDIL
C1095918|T121|319839|RXNORM|MACA PREPARATION|MACA PREPARATION
C3864829|T129|1596933|RXNORM|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 52 VACCINE|L1 PROTEIN, HUMAN PAPILLOMAVIRUS TYPE 52 VACCINE
C3527644|T109|1360630|RXNORM|ARTEMISIA VULGARIS TOP OIL|ARTEMISIA VULGARIS TOP OIL
C0066969|T109|1360631|RXNORM|MUSTARD OIL|MUSTARD OIL
C0053570|T121|19295|RXNORM|BIFONAZOLE|BIFONAZOLE
C0302227|T168|1318515|RXNORM|APRICOT KERNEL OIL|APRICOT KERNEL OIL
C2701427|T129|852229|RXNORM|AUSTRALIAN PINE POLLEN EXTRACT|CASUARINA EQUISETIFOLIA POLLEN EXTRACT
C3256012|T121|1363589|RXNORM|HYPROMELLOSE 2910 3CP|HYPROMELLOSE 2910 3CP
C0074722|T121|36676|RXNORM|SODIUM BICARBONATE|SODIUM BICARBONATE
C0074722|T121|36676|RXNORM|SODIUM BICARBONATE|SODIUM BICARBONATE
C0074722|T121|36676|RXNORM|SODIUM BICARBONATE|SODIUM BICARBONATE
C3256736|T121|1310537|RXNORM|UNDECYL ALCOHOL|UNDECYL ALCOHOL
C0287041|T121|83515|RXNORM|EPROSARTAN|EPROSARTAN
C3256228|T109|1363580|RXNORM|DIPALMITOYL HYDROXYPROLINE|DIPALMITOYL HYDROXYPROLINE
C3256387|T121|1310538|RXNORM|TRIHYDROXYSTEARIN|TRIHYDROXYSTEARIN
C2827134|T130|1310539|RXNORM|DI-(4-TERT-BUTYLCYCLOHEXYL)PEROXYDICARBONATE|DI-(4-TERT-BUTYLCYCLOHEXYL)PEROXYDICARBONATE
C0982206|T121|1363585|RXNORM|HYDROXYPROPYL METHYLCELLULOSE 2208|HYDROXYPROPYL METHYLCELLULOSE 2208
C2825379|T130|1363584|RXNORM|HYDROXYPROPYL CELLULOSE, LOW SUBSTITUTED|LOW-SUBSTITUTED HYDROXYPROPYL CELLULOSE, UNSPECIFIED
C0122862|T130|1363587|RXNORM|HYDROXYPROPYL METHYLCELLULOSE PHTHALATE|HYDROXYPROPYL METHYLCELLULOSE PHTHALATE
C0982207|T121|1363586|RXNORM|HYDROXYPROPYL METHYLCELLULOSE 2910|HYDROXYPROPYL METHYLCELLULOSE 2910
C2186920|T121|820630|RXNORM|BENZTHIAZIDE / RESERPINE|BENZTHIAZIDE / RESERPINE
C0077373|T121|1537576|RXNORM|TROCLOSENE|TROCLOSENE
C2927999|T121|1007076|RXNORM|CHLORHEXIDINE / SODIUM NITRITE|CHLORHEXIDINE / SODIUM NITRITE
C2927998|T121|1007075|RXNORM|BEAN POD EXTRACT / GREEN TEA EXTRACT|BEAN POD EXTRACT / GREEN TEA EXTRACT
C2927996|T121|1007073|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / VITAMIN E|DOCOSAHEXAENOATE / EICOSAPENTAENOATE / VITAMIN E
C2927994|T121|1007071|RXNORM|CALCIUM CHLORIDE / GLUCOSE / GLUTATHIONE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC|CALCIUM CHLORIDE / GLUCOSE / GLUTATHIONE / MAGNESIUM CHLORIDE / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE / SODIUM PHOSPHATE, DIBASIC
C2756330|T129|967970|RXNORM|PYRETHRUM CINERARIIFOLIUM ALLERGENIC EXTRACT|TANACETUM CINERARIIFOLIUM ALLERGENIC EXTRACT
C2928001|T121|1007078|RXNORM|COMPOUND BENZOIN TINCTURE (USP) / PODOPHYLLUM PREPARATION|COMPOUND BENZOIN TINCTURE (USP) / PODOPHYLLUM PREPARATION
C2928002|T121|1007079|RXNORM|BELLADONNA EXTRACT, USP / CHLORPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE|BELLADONNA EXTRACT, USP / CHLORPHENIRAMINE / PHENYLEPHRINE / PYRILAMINE
C0770206|T125|1309342|RXNORM|INSULIN, PORK|INSULIN, PORK
C3488937|T109|1309347|RXNORM|GERANIUM OIL, ALGERIAN TYPE|GERANIUM OIL, ALGERIAN TYPE
C2740597|T129|899378|RXNORM|BLACKBERRY ALLERGENIC EXTRACT|RUBUS ALLEGHENIENSIS ALLERGENIC EXTRACT
C0025746|T130|6878|RXNORM|METHYLENE BLUE|METHYLENE BLUE
C0025746|T130|6878|RXNORM|METHYLENE BLUE|METHYLENE BLUE
C0025744|T121|6877|RXNORM|METHYLDOPATE|METHYLDOPATE
C0025741|T121|6876|RXNORM|METHYLDOPA|METHYLDOPA (LEVOROTATORY)
C0025729|T130|6873|RXNORM|METHYLCELLULOSE|METHYLCELLULOSE
C0025729|T130|6873|RXNORM|METHYLCELLULOSE|METHYLCELLULOSE
C0025729|T130|6873|RXNORM|METHYLCELLULOSE|METHYLCELLULOSE
C0051254|T121|17393|RXNORM|ALOXIPRIN|ALOXIPRIN
C1875173|T121|689313|RXNORM|FRUCTOSE / GLUCOSE / PHOSPHORIC ACID|FRUCTOSE / GLUCOSE / PHOSPHORIC ACID
C0057899|T121|1425983|RXNORM|DIDECYLDIMETHYLAMMONIUM|DIDECYLDIMETHYLAMMONIUM
C3486803|T121|1311332|RXNORM|SUS SCROFA MAMMARY GLAND PREPARATION|PORCINE MAMMARY GLAND PREPARATION
C3486801|T121|1311330|RXNORM|SUS SCROFA LUNG PREPARATION|PORCINE LUNG PREPARATION
C3486806|T121|1311337|RXNORM|SUS SCROFA PANCREAS PREPARATION|PORCINE PANCREAS PREPARATION
C3486805|T121|1311336|RXNORM|SUS SCROFA OVARY PREPARATION|PORCINE OVARY PREPARATION
C3486804|T121|1311334|RXNORM|SUS SCROFA NASAL MUCOSA PREPARATION|PORCINE NASAL MUCOSA PREPARATION
C2949004|T121|1045449|RXNORM|ETHANOL / MENTHOL|ETHANOL / MENTHOL
C3486827|T121|1311338|RXNORM|SUS SCROFA PLACENTA PREPARATION|PORCINE PLACENTA PREPARATION
C2928174|T121|1007252|RXNORM|CALCIUM ASCORBATE / CALCIUM THREONATE / FERROUS ASPARTO GLYCINATE / LIVER STOMACH CONCENTRATE / SUCCINIC ACID / VITAMIN B 12|CALCIUM ASCORBATE / CALCIUM THREONATE / FERROUS ASPARTO GLYCINATE / LIVER STOMACH CONCENTRATE / SUCCINIC ACID / VITAMIN B 12
C2928175|T121|1007253|RXNORM|CALCIUM CARBONATE / GELATIN / MAGNESIUM OXIDE|CALCIUM CARBONATE / GELATIN / MAGNESIUM OXIDE
C2928172|T121|1007250|RXNORM|ALANINE / ARGININE / DIBASIC POTASSIUM PHOSPHATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / PROLINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE|ALANINE / ARGININE / DIBASIC POTASSIUM PHOSPHATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / MAGNESIUM CHLORIDE / METHIONINE / PHENYLALANINE / PROLINE / SODIUM ACETATE / SODIUM CHLORIDE / THREONINE / TRYPTOPHAN / TYROSINE / VALINE
C2928173|T121|1007251|RXNORM|COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / SODIUM ASCORBATE / THIAMINE / VITAMIN B 12 / ZINC SULFATE|COPPER SULFATE / FERROUS FUMARATE / FOLIC ACID / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / SODIUM ASCORBATE / THIAMINE / VITAMIN B 12 / ZINC SULFATE
C2928178|T121|1007256|RXNORM|CLIOQUINOL / DEXAMETHASONE|CLIOQUINOL / DEXAMETHASONE
C2928179|T121|1007257|RXNORM|PHENYLEPHRINE / PREDNISOLONE|PHENYLEPHRINE / PREDNISOLONE
C2928176|T121|1007254|RXNORM|DEXPANTHENOL / NIACINAMIDE / RIBOFLAVIN / THIAMINE / VITAMIN B6|DEXPANTHENOL / NIACINAMIDE / RIBOFLAVIN / THIAMINE / VITAMIN B6
C2928177|T121|1007255|RXNORM|BENZYL ALCOHOL / LIDOCAINE|BENZYL ALCOHOL / LIDOCAINE
C2928180|T121|1007258|RXNORM|ISONIAZID / VITAMIN B6|ISONIAZID / VITAMIN B6
C2928181|T121|1007259|RXNORM|MUMPS VIRUS VACCINE LIVE, JERYL LYNN STRAIN / RUBELLA VIRUS VACCINE LIVE (WISTAR RA 27-3 STRAIN)|MUMPS VIRUS VACCINE LIVE, JERYL LYNN STRAIN / RUBELLA VIRUS VACCINE LIVE (WISTAR RA 27-3 STRAIN)
C2080627|T121|819182|RXNORM|MEPHOBARBITAL / PHENOBARBITAL / PHENYTOIN|MEPHOBARBITAL / PHENOBARBITAL / PHENYTOIN
C3256273|T109|1426343|RXNORM|SACCHAROMYCES LYSATE EXTRACT|SACCHAROMYCES LYSATE EXTRACT
C3474180|T168|1337618|RXNORM|WALNUT OIL|WALNUT OIL
C3254764|T121|1311606|RXNORM|AMYL CINNAMAL|AMYL CINNAMAL
C0772459|T129|237121|RXNORM|ESCHERICHIA COLI ANTIGEN|ESCHERICHIA COLI ANTIGEN
C0066139|T121|29682|RXNORM|METHIXENE|METIXENE
C0028752|T130|7602|RXNORM|O-PHTHALALDEHYDE|O-PHTHALALDEHYDE
C3256735|T121|1314301|RXNORM|ULVA COMPRESSA PROTEIN (ACID HYDROLYZED, 300-5000 MW)|ULVA COMPRESSA PROTEIN (ACID HYDROLYZED, 300-5000 MW)
C3256714|T121|1314300|RXNORM|OLETH-20|OLETH-20
C3256862|T121|1314303|RXNORM|PROPYLENE GLYCOL, (R)-|PROPYLENE GLYCOL, (R)-
C3255684|T168|1311604|RXNORM|HIPPOPHAE RHAMNOIDES FRUIT JUICE|HIPPOPHAE RHAMNOIDES FRUIT JUICE
C0035930|T196|1311489|RXNORM|RUBIDIUM|RUBIDIUM
C0910966|T121|1311488|RXNORM|POLY(VINYLPYRROLIDONE-CO-VINYL-ACETATE)|POLY(VINYLPYRROLIDONE-CO-VINYL-ACETATE)
C1608842|T121|1314307|RXNORM|CERAMIDE 6 II|CERAMIDE 6 II
C3282411|T121|1314306|RXNORM|ETHYLHEXYL LAURATE|ETHYLHEXYL LAURATE
C0282842|T123|1311485|RXNORM|CETYL PALMITATE|CETYL PALMITATE
C0015180|T196|1311484|RXNORM|EUROPIUM|EUROPIUM
C0765273|T121|233272|RXNORM|BEXAROTENE|BEXAROTENE
C0032904|T196|1311481|RXNORM|PRASEODYMIUM|PRASEODYMIUM
C1566537|T129|595060|RXNORM|RANIBIZUMAB|RANIBIZUMAB
C0014688|T196|1311483|RXNORM|ERBIUM|ERBIUM
C0013407|T196|1311482|RXNORM|DYSPROSIUM|DYSPROSIUM
C3465010|T121|1309966|RXNORM|CANANGA ODORATA FLOWER EXTRACT|CANANGA ODORATA FLOWER EXTRACT
C2948691|T121|1044578|RXNORM|CAMPHOR / CAPSAICIN / MENTHOL / METHYL SALICYLATE|CAMPHOR / CAPSAICIN / MENTHOL / METHYL SALICYLATE
C3486667|T121|1309961|RXNORM|ILEX AQUIFOLIUM FLOWERING TOP EXTRACT|ILEX AQUIFOLIUM FLOWERING TOP EXTRACT
C3486666|T121|1309960|RXNORM|IBERIS AMARA SEED EXTRACT|IBERIS AMARA SEED EXTRACT
C0756085|T195|229369|RXNORM|DALFOPRISTIN|DALFOPRISTIN
C3499594|T121|1312464|RXNORM|AMMONIUM CHLORIDE / POTASSIUM IODIDE|AMMONIUM CHLORIDE / POTASSIUM IODIDE
C1172637|T121|1311600|RXNORM|ABETIMUS|ABETIMUS
C2960912|T121|1043562|RXNORM|METFORMIN / SAXAGLIPTIN|METFORMIN / SAXAGLIPTIN
C3465016|T121|1309969|RXNORM|HEMIDESMUS INDICUS ROOT EXTRACT|HEMIDESMUS INDICUS ROOT EXTRACT
C3486670|T121|1309968|RXNORM|CARDIOSPERMUM HALICACABUM FLOWERING TOP EXTRACT|CARDIOSPERMUM HALICACABUM FLOWERING TOP EXTRACT
C0873126|T121|259460|RXNORM|BORAGE EXTRACT|BORAGE EXTRACT
C3859157|T109|1592258|RXNORM|METHYL GLUCOSE SESQUISTEARATE|METHYL GLUCOSE SESQUISTEARATE
C1873987|T121|689788|RXNORM|ACETAMINOPHEN / MEPERIDINE|ACETAMINOPHEN / MEPERIDINE
C0677666|T121|196238|RXNORM|SOY PROTEIN ISOLATE|SOY PROTEIN ISOLATE
C1873985|T121|689785|RXNORM|ACETAMINOPHEN / DIPHENHYDRAMINE / PHENYLEPHRINE|ACETAMINOPHEN / DIPHENHYDRAMINE / PHENYLEPHRINE
C1873986|T121|689786|RXNORM|ACETAMINOPHEN / DIPHENHYDRAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / DIPHENHYDRAMINE / PSEUDOEPHEDRINE
C1873986|T121|689786|RXNORM|ACETAMINOPHEN / DIPHENHYDRAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / DIPHENHYDRAMINE / PSEUDOEPHEDRINE
C1873983|T121|689780|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE|ACETAMINOPHEN / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE
C1873984|T121|689783|RXNORM|ACETAMINOPHEN / DIHYDROCODEINE / SALICYLAMIDE|ACETAMINOPHEN / DIHYDROCODEINE / SALICYLAMIDE
C2929450|T121|1008547|RXNORM|BELLADONNA EXTRACT, USP / BUTABARBITAL|BELLADONNA EXTRACT, USP / BUTABARBITAL
C2929449|T121|1008546|RXNORM|ALOE EXTRACT / SENNOSIDES, USP|ALOE EXTRACT / SENNOSIDES, USP
C2929448|T121|1008545|RXNORM|4-AMINOBENZOIC ACID / ARGININE|4-AMINOBENZOIC ACID / ARGININE
C2929447|T121|1008544|RXNORM|ECHINACEA PURPUREA EXTRACT / MENTHOL|ECHINACEA PURPUREA EXTRACT / MENTHOL
C2929446|T121|1008543|RXNORM|BUTHIAZIDE / RESERPINE|BUTHIAZIDE / RESERPINE
C2929445|T121|1008542|RXNORM|ACETIC ACID / ANTIPYRINE / BENZOCAINE|ACETIC ACID / ANTIPYRINE / BENZOCAINE
C2929443|T121|1008540|RXNORM|ASCORBIC ACID / NIACIN / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN D / VITAMIN E|ASCORBIC ACID / NIACIN / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN D / VITAMIN E
C0051724|T197|17792|RXNORM|AMMONIUM PHOSPHATE|AMMONIUM PHOSPHATE
C2929452|T121|1008549|RXNORM|METHENAMINE / PHENAZOPYRIDINE|METHENAMINE / PHENAZOPYRIDINE
C2929451|T121|1008548|RXNORM|ALLANTOIN / BENZOCAINE / CAMPHOR / PETROLATUM|ALLANTOIN / BENZOCAINE / CAMPHOR / PETROLATUM
C0004482|T131|1256|RXNORM|AZATHIOPRINE|AZATHIOPRINE
C0005330|T121|1525|RXNORM|BEZAFIBRATE|BEZAFIBRATE
C0108121|T121|47622|RXNORM|CALCIUM LACTATE|CALCIUM 2-HYDROXYPROPANOATE
C0005320|T121|1520|RXNORM|BETAXOLOL|BETAXOLOL
C0005320|T121|1520|RXNORM|BETAXOLOL|BETAXOLOL
C0064694|T109|28486|RXNORM|LAVENDER OIL|LAVENDER OIL
C1874936|T121|690300|RXNORM|CRYPTENAMINE / METHYCLOTHIAZIDE|CRYPTENAMINE / METHYCLOTHIAZIDE
C0108134|T197|47627|RXNORM|CALCIUM PHOSPHATE DIBASIC|CALCIUM PHOSPHATE DIBASIC
C0108136|T197|47628|RXNORM|TRICALCIUM PHOSPHATE|TRICALCIUM PHOSPHATE
C0301504|T129|89887|RXNORM|LATRODECTUS MACTANS ANTIVENIN|LATRODECTUS MACTANS ANTIVENIN
C0045287|T121|1368138|RXNORM|2,2-BIS(4-GLYCIDYLOXYPHENYL)PROPANE|2,2-BIS(4-GLYCIDYLOXYPHENYL)PROPANE
C2057748|T121|821526|RXNORM|ETOFYLLINE / THEOPHYLLINE|ETOFYLLINE / THEOPHYLLINE
C2939773|T121|1592257|RXNORM|LEVOMEFOLATE|L-METHYLFOLATE
C1875446|T121|690902|RXNORM|LITHIUM CARBONATE / SODIUM CHLORIDE|LITHIUM CARBONATE / SODIUM CHLORIDE
C0249529|T121|73689|RXNORM|FEBUXOSTAT|FEBUXOSTAT
C1720107|T121|1000705|RXNORM|BENZALKONIUM / TOLNAFTATE|BENZALKONIUM / TOLNAFTATE
C3833353|T109|1541234|RXNORM|AMMONIUM ACRYLOYLDIMETHYLTAURATE - BEHENETH-25 METHACRYLATE CROSSPOLYMER (52000 MPA.S)|AMMONIUM ACRYLOYLDIMETHYLTAURATE - BEHENETH-25 METHACRYLATE CROSSPOLYMER (52000 MPA.S)
C0014964|T121|4110|RXNORM|ETHAMBUTOL|ETHAMBUTOL
C1827585|T121|1000706|RXNORM|BENZOCAINE / SALICYLAMIDE|BENZOCAINE / SALICYLAMIDE
C3813322|T121|1541239|RXNORM|FRAGARIA VESCA WHOLE EXTRACT|FRAGARIA VESCA WHOLE EXTRACT
C0358967|T121|1000708|RXNORM|BETAMETHASONE / CLIOQUINOL|BETAMETHASONE / CLIOQUINOL
C2928719|T121|1007804|RXNORM|ACYCLOVIR / HYDROCORTISONE|ACYCLOVIR / HYDROCORTISONE
C0062106|T121|26422|RXNORM|HALOPROGIN|HALOPROGIN
C0014987|T121|4118|RXNORM|ETHCHLORVYNOL|ETHCHLORVYNOL
C3257442|T121|1368136|RXNORM|BETASIZOFIRAN|BETASIZOFIRAN
C3527806|T121|1361211|RXNORM|CHLOROXYLENOL / IODINE / MENTHOL|CHLOROXYLENOL / IODINE / MENTHOL
C1721377|T121|662281|RXNORM|NILOTINIB|NILOTINIB
C0051908|T121|17933|RXNORM|ANILERIDINE|ANILERIDINE
C3665584|T121|1487834|RXNORM|POGOSTEMON CABLIN WHOLE EXTRACT|POGOSTEMON CABLIN WHOLE EXTRACT
C3709598|T121|1487835|RXNORM|BUTYL LEVULINATE|BUTYL LEVULINATE
C3669110|T121|1487832|RXNORM|MELALEUCA ALTERNIFOLIA WHOLE EXTRACT|MELALEUCA ALTERNIFOLIA WHOLE EXTRACT
C0003781|T196|1368133|RXNORM|ARGON|ARGON
C3669245|T121|1487830|RXNORM|GERANIUM MACULATUM WHOLE EXTRACT|GERANIUM MACULATUM WHOLE EXTRACT
C3669383|T121|1487831|RXNORM|HYOSCYAMUS NIGER LEAF EXTRACT|HYOSCYAMUS NIGER LEAF EXTRACT
C2722035|T129|891611|RXNORM|COCONUT ALLERGENIC EXTRACT|COCOS NUCIFERA ALLERGENIC EXTRACT
C0069488|T121|32411|RXNORM|OMOCONAZOLE|OMOCONAZOLE
C2701778|T129|852750|RXNORM|WESTERN SYCAMORE POLLEN EXTRACT|PLATANUS RACEMOSA POLLEN EXTRACT
C2940192|T129|1014743|RXNORM|WHITE (MEXICAN) DOCK POLLEN EXTRACT|RUMEX SALICIFOLIUS VAR. MEXICANUS POLLEN EXTRACT
C1110649|T121|324039|RXNORM|FRANGULA PREPARATION|FRANGULA PREPARATION
C2701404|T129|852205|RXNORM|MUSTARD POLLEN EXTRACT|BRASSICA RAPA POLLEN EXTRACT
C3502823|T121|1368642|RXNORM|GENTISATE|GENTISATE
C2940196|T129|1014749|RXNORM|ABSIDIA RAMOSA EXTRACT|ABSIDIA RAMOSA EXTRACT
C0981993|T129|852209|RXNORM|YELLOW DOCK POLLEN EXTRACT|RUMEX CRISPUS POLLEN EXTRACT
C3848607|T121|1544485|RXNORM|FUMARYL DIKETOPIPERAZINE|FUMARYL DIKETOPIPERAZINE
C3848608|T121|1544484|RXNORM|EICHHORNIA CRASSIPES WHOLE EXTRACT|EICHHORNIA CRASSIPES WHOLE EXTRACT
C0360428|T121|107999|RXNORM|CETRIMIDE / CHLORHEXIDINE|CETRIMIDE / CHLORHEXIDINE
C2929043|T121|1008136|RXNORM|THIAMINE / VITAMIN B6|THIAMINE / VITAMIN B6
C2929044|T121|1008137|RXNORM|ASCORBIC ACID / MENTHOL|ASCORBIC ACID / MENTHOL
C2929041|T121|1008134|RXNORM|ECHINACEA PURPUREA EXTRACT / GOLDENSEAL EXTRACT|ECHINACEA PURPUREA EXTRACT / GOLDENSEAL EXTRACT
C2929042|T121|1008135|RXNORM|ASCORBIC ACID / FERROUS GLUCONATE / VITAMIN B 12|ASCORBIC ACID / FERROUS GLUCONATE / VITAMIN B 12
C2929039|T121|1008132|RXNORM|CLOBETASONE / NEOMYCIN|CLOBETASONE / NEOMYCIN
C2929040|T121|1008133|RXNORM|LYAPOLATE / NIACIN|LYAPOLATE / NIACIN
C2929037|T121|1008130|RXNORM|CHOLINE / GLUTAMINE / INOSITOL|CHOLINE / GLUTAMINE / INOSITOL
C2929038|T121|1008131|RXNORM|HYOSCYAMINE / PAPAVERINE|HYOSCYAMINE / PAPAVERINE
C3465209|T121|1313223|RXNORM|ACETYL TRIETHYLHEXYL CITRATE|ACETYL TRIETHYLHEXYL CITRATE
C3464314|T121|1313222|RXNORM|ACETYL CARBOXYMETHYL COCOYL GLYCINE|ACETYL CARBOXYMETHYL COCOYL GLYCINE
C3267308|T121|1313221|RXNORM|2-O-ETHYL ASCORBIC ACID|2-O-ETHYL ASCORBIC ACID
C3264671|T109|1313220|RXNORM|2-ETHYLAMINOETHANOL|2-ETHYLAMINOETHANOL
C3265015|T121|1313227|RXNORM|C30-45 ALKYL METHICONE|C30-45 ALKYL METHICONE
C3486286|T109|1313226|RXNORM|BIS-ETHYLHEXYL HYDROXYDIMETHOXY BENZYLMALONATE|BIS-ETHYLHEXYL HYDROXYDIMETHOXY BENZYLMALONATE
C2929045|T121|1008138|RXNORM|4-AMINOBENZOATE / SALICYLIC ACID|4-AMINOBENZOATE / SALICYLIC ACID
C2929046|T121|1008139|RXNORM|SODIUM FLUORIDE / SODIUM PHOSPHATE, MONOBASIC|SODIUM FLUORIDE / SODIUM PHOSPHATE, MONOBASIC
C3848591|T121|1545684|RXNORM|ONONIS REPENS ROOT EXTRACT|ONONIS REPENS ROOT EXTRACT
C3848590|T121|1545685|RXNORM|PHENYL BUTYRATE|PHENYL BUTYRATE
C0021978|T121|5942|RXNORM|CLIOQUINOL|CLIOQUINOL
C3848592|T121|1545681|RXNORM|CICHORIUM INTYBUS WHOLE EXTRACT|CICHORIUM INTYBUS WHOLE EXTRACT
C3714586|T121|1545682|RXNORM|COLCHICUM AUTUMNALE WHOLE EXTRACT|COLCHICUM AUTUMNALE WHOLE EXTRACT
C3812198|T121|1545683|RXNORM|KRAMERIA LAPPACEA WHOLE EXTRACT|KRAMERIA LAPPACEA WHOLE EXTRACT
C3535914|T130|1368644|RXNORM|CARMINATE|CARMINATE
C3255925|T121|1372007|RXNORM|CITRUS NOBILIS EXTRACT|CITRUS NOBILIS EXTRACT
C0062922|T121|27084|RXNORM|HOMATROPINE|HOMATROPINE
C0062922|T121|27084|RXNORM|HOMATROPINE|HOMATROPINE
C3256034|T121|1312551|RXNORM|DIETHYLHEXYL MALEATE|DIETHYLHEXYL MALEATE
C0071071|T121|1110783|RXNORM|PIMOBENDAN|PIMOBENDAN
C0064657|T122|28456|RXNORM|LAPYRIUM|LAPYRIUM
C1831731|T121|1307619|RXNORM|BOSUTINIB|BOSUTINIB
C3256782|T121|1307618|RXNORM|LARREA DIVARICATA LEAF EXTRACT|LARREA DIVARICATA LEAF EXTRACT
C3474582|T121|1307617|RXNORM|DUBOISIA LEICHHARDTII LEAF EXTRACT|DUBOISIA LEICHHARDTII LEAF EXTRACT
C3485016|T121|1307614|RXNORM|PLATYCODON GRANDIFLORUM ROOT EXTRACT|PLATYCODON GRANDIFLORUM ROOT EXTRACT
C3256709|T121|1307613|RXNORM|OENOTHERA BIENNIS FLOWERING TOP EXTRACT|OENOTHERA BIENNIS FLOWERING TOP EXTRACT
C3256252|T121|1307612|RXNORM|PHELLODENDRON CHINENSIS BARK EXTRACT|PHELLODENDRON CHINENSIS BARK EXTRACT
C3256226|T121|1307611|RXNORM|DIOSCOREA JAPONICA ROOT EXTRACT|DIOSCOREA JAPONICA ROOT EXTRACT
C3256327|T121|1307610|RXNORM|ACMELLA OLERACEA FLOWER EXTRACT|ACMELLA OLERACEA FLOWER EXTRACT
C3535912|T121|1368648|RXNORM|FERULATE|FERULATE
C3535849|T122|1370641|RXNORM|COCOAMPHODIPROPIONATE|COCOAMPHODIPROPIONATE
C3651950|T121|1429359|RXNORM|CHLOPHEDIANOL / PYRILAMINE|CHLOPHEDIANOL / PYRILAMINE
C3256264|T109|1309509|RXNORM|RUSCUS ACULEATUS ROOT EXTRACT|RUSCUS ACULEATUS ROOT EXTRACT
C3162766|T121|1114864|RXNORM|COCOA BUTTER / PHENYLEPHRINE|COCOA BUTTER / PHENYLEPHRINE
C3488152|T121|1309501|RXNORM|AGRIMONIA EUPATORIA FLOWER EXTRACT|AGRIMONIA EUPATORIA FLOWER EXTRACT
C3256270|T109|1309500|RXNORM|RORIPPA NASTURTIUM-AQUATICUM FLOWERING TOP EXTRACT|RORIPPA NASTURTIUM-AQUATICUM FLOWERING TOP EXTRACT
C2947473|T121|1309503|RXNORM|ALOE FEROX LEAF PREPARATION|ALOE FEROX LEAF PREPARATION
C0060389|T125|25025|RXNORM|FINASTERIDE|FINASTERIDE
C3256262|T109|1309505|RXNORM|ROSMARINUS OFFICINALIS FLOWER EXTRACT|ROSMARINUS OFFICINALIS FLOWER EXTRACT
C3489266|T121|1309504|RXNORM|AGRIMONIA EUPATORIA FLOWERING TOP EXTRACT|AGRIMONIA EUPATORIA FLOWERING TOP EXTRACT
C3256263|T121|1309507|RXNORM|RUBUS FRUTICOSUS LEAF EXTRACT|RUBUS FRUTICOSUS LEAF EXTRACT
C3488139|T121|1309506|RXNORM|APOCYNUM CANNABINUM ROOT EXTRACT|APOCYNUM CANNABINUM ROOT EXTRACT
C1875525|T121|693011|RXNORM|NEOMYCIN / PREDNISOLONE|NEOMYCIN / PREDNISOLONE
C1875523|T121|693010|RXNORM|NEOMYCIN / POLYMYXIN B / PREDNISOLONE|NEOMYCIN / POLYMYXIN B / PREDNISOLONE
C0063242|T121|27334|RXNORM|HYPROMELLOSE|HYPROMELLOSE
C0070276|T121|33055|RXNORM|PENTAERYTHRITOL|PENTAERYTHRITOL
C3854896|T121|1546887|RXNORM|ABACAVIR / DOLUTEGRAVIR / LAMIVUDINE|ABACAVIR / DOLUTEGRAVIR / LAMIVUDINE
C0795671|T121|253204|RXNORM|TRISODIUM CITRATE|TRISODIUM CITRATE
C2193876|T121|821514|RXNORM|IODOQUINOL / METRONIDAZOLE|IODOQUINOL / METRONIDAZOLE
C2740760|T129|899661|RXNORM|CAULIFLOWER ALLERGENIC EXTRACT|CAULIFLOWER ALLERGENIC EXTRACT
C2074989|T121|817588|RXNORM|CILAZAPRIL / HYDROCHLOROTHIAZIDE|CILAZAPRIL / HYDROCHLOROTHIAZIDE
C0034738|T121|9154|RXNORM|RAZOXANE|RAZOXANE
C2702222|T109|853406|RXNORM|COTTONSEED EXTRACT|COTTONSEED EXTRACT
C2080571|T121|817275|RXNORM|ASPIRIN / BROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE|ASPIRIN / BROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLPROPANOLAMINE
C0126948|T121|52403|RXNORM|MANGANESE GLUCONATE|MANGANESE GLUCONATE
C3256718|T121|1314209|RXNORM|PPG-2 ISOCETETH-20 ACETATE|PPG-2 ISOCETETH-20 ACETATE
C4048291|T123|1368166|RXNORM|HYDROXYLYSINE|5-HYDROXYLYSINE
C0031560|T109|1368167|RXNORM|PHLORETIN|PHLORETIN
C3256971|T109|1368164|RXNORM|TRIDECYL NEOPENTANOATE|TRIDECYL NEOPENTANOATE
C3256557|T109|1368165|RXNORM|POLYETHYLENE GLYCOL 350|POLYETHYLENE GLYCOL 350
C3256790|T121|1368162|RXNORM|NEOPENTYL GLYCOL|NEOPENTYL GLYCOL
C3257695|T121|1368163|RXNORM|COLLAGEN, SOLUBLE, FISH SKIN|MARINE COLLAGEN, SOLUBLE
C3474292|T121|1368160|RXNORM|PALMITOYL DIPEPTIDE-7|PALMITOYL LYSYLTHREONINE
C3257507|T109|1368161|RXNORM|POLYESTER-7|POLYESTER-7
C0022176|T121|6023|RXNORM|ISOETHARINE|ISOETARINE
C0022180|T121|6026|RXNORM|ISOFLURANE|ISOFLURANE
C0022181|T131|6027|RXNORM|ISOFLUROPHATE|ISOFLUROPHATE
C0770689|T129|235574|RXNORM|MEASLES VIRUS VACCINE,LIVE ATTENUATED|MEASLES, LIVE ATTENUATED
C0038329|T123|10079|RXNORM|STIGMASTEROL|STIGMASTEROL
C0178638|T127|62356|RXNORM|FOLATE|FOLATE
C3651748|T121|1429042|RXNORM|PORTULACA OLERACEA LEAF EXTRACT|PORTULACA OLERACEA LEAF EXTRACT
C3256552|T121|1314200|RXNORM|POLYESTER-10|POLYESTER-10
C0674428|T121|195085|RXNORM|EFAVIRENZ|EFAVIRENZ
C1739045|T121|1427136|RXNORM|N-CYCLOHEXYL-N'-PHENYL-1,4-PHENYLENEDIAMINE|N-CYCLOHEXYL-N'-PHENYL-1,4-PHENYLENEDIAMINE
C3256553|T121|1314201|RXNORM|POLYESTER-8 (1400 MW, CYANODIPHENYLPROPENOYL CAPPED)|POLYESTER-8 (1400 MW, CYANODIPHENYLPROPENOYL CAPPED)
C0982237|T130|314691|RXNORM|IODOHIPPURATE|IODOHIPPURATE
C3256795|T121|1427139|RXNORM|OPHIOCORDYCEPS SINENSIS EXTRACT|OPHIOCORDYCEPS SINENSIS EXTRACT
C3256912|T109|1305635|RXNORM|ECHIUM PLANTAGINEUM SEED OIL|ECHIUM PLANTAGINEUM SEED OIL
C0674432|T121|195088|RXNORM|LOPINAVIR|LOPINAVIR
C1445799|T121|466565|RXNORM|PRAMOXINE / ZINC OXIDE|PRAMOXINE / ZINC OXIDE
C3535867|T130|1370618|RXNORM|LAUROYL SARCOSINATE|LAUROYL SARCOSINATE
C0771603|T121|236340|RXNORM|ALEXITOL SODIUM|ALEXITOL SODIUM
C1445800|T121|466566|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / DIPHENHYDRAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / DEXTROMETHORPHAN / DIPHENHYDRAMINE / PSEUDOEPHEDRINE
C0771610|T121|236346|RXNORM|DIMECROTIC ACID|DIMECROTIC ACID
C0771607|T121|236344|RXNORM|SAW PALMETTO EXTRACT|SAW PALMETTO EXTRACT
C3535872|T123|1370611|RXNORM|SARCOSINATE|SARCOSINATE
C2827308|T121|1314204|RXNORM|POLYETHYLENE GLYCOL 900|POLYETHYLENE GLYCOL 900
C0771612|T121|236348|RXNORM|MORPHOLINE SALICYLATE|MORPHOLINE SALICYLATE
C3535871|T121|1370612|RXNORM|ETHYLENEDIAMINE DISUCCINATE|ETHYLENEDIAMINE DISUCCINATE
C1445803|T121|466569|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|ACETAMINOPHEN / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C1445803|T121|466569|RXNORM|ACETAMINOPHEN / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|ACETAMINOPHEN / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C1445802|T121|466568|RXNORM|CHLORPHENIRAMINE / CODEINE / PSEUDOEPHEDRINE|CHLORPHENIRAMINE / CODEINE / PSEUDOEPHEDRINE
C3535868|T121|1370617|RXNORM|LAURETH-2 SULFATE|LAURETH-2 SULFATE
C3535820|T121|1370616|RXNORM|ISOSTEAROYL LACTYLATE|ISOSTEAROYL LACTYLATE
C3256637|T121|1314206|RXNORM|POLYISOBUTYLENE (35000 MW)|POLYISOBUTYLENE (35000 MW)
C2146454|T121|817623|RXNORM|SULFAMETROLE / TRIMETHOPRIM|SULFAMETROLE / TRIMETHOPRIM
C3465269|T121|1305630|RXNORM|ZINGIBER CASSUMUNAR ROOT EXTRACT|ZINGIBER CASSUMUNAR ROOT EXTRACT
C0093437|T121|44281|RXNORM|CEVIMELINE|CEVIMELINE
C0034417|T121|9071|RXNORM|QUININE|QUININE
C3488280|T121|1309714|RXNORM|CROTON TIGLIUM SEED EXTRACT|CROTON TIGLIUM SEED EXTRACT
C2930696|T121|1357536|RXNORM|TOFACITINIB|TOFACITINIB
C3257524|T109|1311817|RXNORM|CULTIVATED MUSHROOM EXTRACT|CULTIVATED MUSHROOM EXTRACT
C2935868|T121|1311811|RXNORM|ALPHA-HEXYLCINNAMALDEHYDE|ALPHA-HEXYLCINNAMALDEHYDE
C3857942|T121|1552631|RXNORM|FERROUS PICRATE|FERROUS PICRATE
C3857941|T121|1552632|RXNORM|EQUUS CABALLUS WHOLE PREPARATION|EQUUS CABALLUS WHOLE PREPARATION
C2740722|T129|899593|RXNORM|MULBERRY POLLEN EXTRACT|BROUSSONETIA PAPYRIFERA POLLEN EXTRACT
C1719965|T121|645082|RXNORM|CHLORHEXIDINE / PHENOL|CHLORHEXIDINE / PHENOL
C1875020|T121|690681|RXNORM|DIETHYLSTILBESTROL / METHYLTESTOSTERONE|DIETHYLSTILBESTROL / METHYLTESTOSTERONE
C0012772|T121|3554|RXNORM|DISULFIRAM|DISULFIRAM
C1875023|T121|690685|RXNORM|DIMENHYDRINATE / NIACIN|DIMENHYDRINATE / NIACIN
C1875025|T121|690688|RXNORM|DIPERODON / HYDROCORTISONE / ZINC OXIDE|DIPERODON / HYDROCORTISONE / ZINC OXIDE
C3495095|T196|1546265|RXNORM|LITHIUM CATION|LITHIUM CATION
C1637395|T121|608531|RXNORM|CHLORHEXIDINE / CHLOROBUTANOL|CHLORHEXIDINE / CHLOROBUTANOL
C0010294|T123|2913|RXNORM|CREATININE|CREATININE
C0010303|T109|2915|RXNORM|CREOSOTE|CREOSOTE
C0002640|T121|719|RXNORM|AMOBARBITAL|AMOBARBITAL
C0002615|T197|712|RXNORM|AMMONIUM CHLORIDE|AMMONIUM CHLORIDE
C0772297|T121|236964|RXNORM|BISMUTH CHLORIDE OXIDE|BISMUTH CHLORIDE OXIDE
C1719859|T121|646063|RXNORM|DIPHENHYDRAMINE / LEVOMENTHOL|DIPHENHYDRAMINE / LEVOMENTHOL
C2929637|T121|1008738|RXNORM|ETHYLNICOTINATE / HEXYLNICOTINATE / THURFYL SALICYLATE|ETHYLNICOTINATE / HEXYLNICOTINATE / THURFYL SALICYLATE
C2929638|T121|1008739|RXNORM|DIHYDROXYALUMINUM SODIUM CARBONATE / DIMETHICONE|DIHYDROXYALUMINUM SODIUM CARBONATE / DIMETHICONE
C2929633|T121|1008734|RXNORM|ASCORBIC ACID / VITAMIN B6|ASCORBIC ACID / VITAMIN B6
C2929634|T121|1008735|RXNORM|NITROFURANTOIN / VITAMIN B6|NITROFURANTOIN / VITAMIN B6
C2929635|T121|1008736|RXNORM|DICYCLOMINE / DOXYLAMINE / VITAMIN B6|DICYCLOMINE / DOXYLAMINE / VITAMIN B6
C2929636|T121|1008737|RXNORM|GAMMA-AMINOBUTYRATE / VITAMIN B6|GAMMA-AMINOBUTYRATE / VITAMIN B6
C2929629|T121|1008730|RXNORM|OX BILE EXTRACT / PANCREATIN|OX BILE EXTRACT / PANCREATIN
C2929630|T121|1008731|RXNORM|ERGOCALCIFEROL / LECITHIN|ERGOCALCIFEROL / LECITHIN
C2929631|T121|1008732|RXNORM|CALCIUM CITRATE / ERGOCALCIFEROL / MAGNESIUM CITRATE|CALCIUM CITRATE / ERGOCALCIFEROL / MAGNESIUM CITRATE
C2929632|T121|1008733|RXNORM|ASCORBIC ACID / BETA CAROTENE / FOLIC ACID / IODINE / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENATE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN D / VITAMIN E / ZINC SULFATE|ASCORBIC ACID / BETA CAROTENE / FOLIC ACID / IODINE / MAGNESIUM SULFATE / MANGANESE SULFATE / NIACINAMIDE / PANTOTHENATE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN B6 / VITAMIN D / VITAMIN E / ZINC SULFATE
C2006118|T121|818119|RXNORM|CALCIUM CARBONATE / POTASSIUM TARTRATE|CALCIUM CARBONATE / POTASSIUM TARTRATE
C0077163|T121|38685|RXNORM|TRIMETHOBENZAMIDE|TRIMETHOBENZAMIDE
C2742503|T129|974779|RXNORM|OBINUTUZUMAB|OBINUTUZUMAB
C0019469|T121|5302|RXNORM|HEXOBARBITAL|HEXOBARBITAL
C0019471|T121|5303|RXNORM|HEXOBENDINE|HEXOBENDINE
C0019476|T121|5307|RXNORM|HEXOPRENALINE|HEXOPRENALINE
C0071021|T123|1363444|RXNORM|PHYTOSPHINGOSINE|PHYTOSPHINGOSINE
C3475292|T109|1363445|RXNORM|POLYGLYCERYL-2 DIPOLYHYDROXYSTEARATE|POLYGLYCERYL-2 DIPOLYHYDROXYSTEARATE
C1509789|T121|1363446|RXNORM|SOY STEROL|SOY STEROL
C1095801|T121|1372258|RXNORM|SPEARMINT EXTRACT|SPEARMINT EXTRACT
C3528821|T109|1363440|RXNORM|PASSIFLORA EDULIS SEED OIL|PASSIFLORA EDULIS SEED OIL
C3528822|T109|1363441|RXNORM|POLYETHYLENE GLYCOL 450|POLYETHYLENE GLYCOL 450
C3528823|T109|1363442|RXNORM|METHYL STEARIC ACID|METHYL STEARIC ACID
C3256372|T109|1363443|RXNORM|MUSKMELON EXTRACT|MUSKMELON EXTRACT
C3864837|T121|1596680|RXNORM|LINDEN LEAF EXTRACT|LINDEN LEAF EXTRACT
C2073805|T121|815833|RXNORM|CHLORAMPHENICOL / DEXAMETHASONE|CHLORAMPHENICOL / DEXAMETHASONE
C0015827|T121|4328|RXNORM|FENFLURAMINE|FENFLURAMINE
C3700891|T121|1486716|RXNORM|OPUNTIA STREPTACANTHA STEM EXTRACT|OPUNTIA STREPTACANTHA STEM EXTRACT
C3700890|T122|1486717|RXNORM|POLYQUATERNIUM-10 (1000 MPA.S AT 2%)|POLYQUATERNIUM-10 (1000 MPA.S AT 2%)
C3700889|T109|1486718|RXNORM|L-ERYTHRULOSE|L-ERYTHRULOSE
C3535923|T121|1369401|RXNORM|CHOLECALCIFEROL / LEVOCARNITINE|CHOLECALCIFEROL / LEVOCARNITINE
C2938093|T121|1011453|RXNORM|CHLORHEXIDINE / DIDECYLDIMETHYLAMMONIUM CHLORIDE|CHLORHEXIDINE / DIDECYLDIMETHYLAMMONIUM CHLORIDE
C0982401|T121|1364939|RXNORM|SODIUM TALLOWATE|SODIUM TALLOWATE
C0283828|T121|1011450|RXNORM|DIDECYLDIMETHYLAMMONIUM CHLORIDE|DIDECYLDIMETHYLAMMONIUM CHLORIDE
C2827592|T129|1484973|RXNORM|BLACK ALDER POLLEN EXTRACT|EUROPEAN ALDER POLLEN EXTRACT
C0082286|T121|3142|RXNORM|DEHYDROEMETINE|DEHYDROEMETINE
C0011185|T125|3143|RXNORM|DEHYDROEPIANDROSTERONE|PRASTERONE
C3695941|T129|1484976|RXNORM|MEADOW BROME POLLEN EXTRACT|BROMUS COMMUTATUS POLLEN EXTRACT
C3695940|T129|1484977|RXNORM|HEATHER POLLEN EXTRACT|COMMON HEATHER POLLEN EXTRACT
C3669203|T129|1484974|RXNORM|MEADOW FOXTAIL POLLEN EXTRACT|FIELD MEADOW FOXTAIL POLLEN EXTRACT
C3695942|T129|1484975|RXNORM|ARGENTINE CANOLA POLLEN EXTRACT|BRASSICA NAPUS SUBSP. NAPUS POLLEN EXTRACT
C3695939|T129|1484978|RXNORM|BLITUM BONUS-HENRICUS POLLEN EXTRACT|GOOD KING HENRY POLLEN EXTRACT
C1440492|T129|1484979|RXNORM|COMMON HAZEL POLLEN EXTRACT|CORYLUS AVELLANA POLLEN EXTRACT
C0916062|T121|280611|RXNORM|BEMIPARIN|BEMIPARIN
C1145759|T121|343047|RXNORM|ATAZANAVIR|ATAZANAVIR
C1302939|T121|392658|RXNORM|ACETAMINOPHEN / METOCLOPRAMIDE|ACETAMINOPHEN / METOCLOPRAMIDE
C1145760|T121|343048|RXNORM|TREPROSTINIL|TREPROSTINIL
C3488960|T109|1309288|RXNORM|ARNICA CHAMISSONIS FLOWER EXTRACT|ARNICA CHAMISSONIS FLOWER EXTRACT
C2911923|T121|1309289|RXNORM|CALENDULA OFFICINALIS FLOWER EXTRACT|CALENDULA OFFICINALIS FLOWER EXTRACT
C3488948|T109|1309286|RXNORM|ANGELICA ARCHANGELICA LEAF EXTRACT|ANGELICA ARCHANGELICA LEAF EXTRACT
C3488957|T109|1309287|RXNORM|TARAXACUM OFFICINALE LEAF EXTRACT|TARAXACUM OFFICINALE LEAF EXTRACT
C3488959|T121|1309284|RXNORM|ACTAEA CIMICIFUGA ROOT EXTRACT|ACTAEA CIMICIFUGA ROOT EXTRACT
C0952248|T121|289996|RXNORM|FORMALDEHYDESULFOXYLATE, MONOSODIUM SALT|FORMALDEHYDESULFOXYLATE, MONOSODIUM SALT
C3255816|T109|1309282|RXNORM|ACAI OIL|ACAI OIL
C3488972|T109|1309283|RXNORM|UNCARIA RHYNCHOPHYLLA STEM|UNCARIA RHYNCHOPHYLLA STEM
C3488958|T109|1309280|RXNORM|ABIES SACHALINENSIS VAR. SACHALINENSIS OIL|ABIES SACHALINENSIS VAR. SACHALINENSIS OIL
C3488973|T121|1309281|RXNORM|URTICA DIOICA LEAF EXTRACT|URTICA DIOICA LEAF EXTRACT
C0063456|T121|1311673|RXNORM|INDELOXAZINE|INDELOXAZINE
C0282774|T121|1311670|RXNORM|PIMAGEDINE|PIMAGEDINE
C3257033|T121|1311671|RXNORM|RUBUS CHAMAEMORUS FRUIT EXTRACT|RUBUS CHAMAEMORUS FRUIT EXTRACT
C0072954|T121|1311677|RXNORM|RACTOPAMINE|RACTOPAMINE
C3256724|T121|1311674|RXNORM|SAPINDUS MUKOROSSI FRUIT EXTRACT|SAPINDUS MUKOROSSI FRUIT EXTRACT
C3254748|T121|1311675|RXNORM|SCHISANDRA CHINENSIS FRUIT EXTRACT|SCHISANDRA CHINENSIS FRUIT EXTRACT
C0066771|T121|1311678|RXNORM|MONOOLEIN|GLYCERYL MONOOLEATE
C2979057|T121|1090016|RXNORM|ASCORBIC ACID / BUTCHER'S BROOM PREPARATION / DIOSMIN / HESPERIDIN|ASCORBIC ACID / BUTCHER'S BROOM PREPARATION / DIOSMIN / HESPERIDIN
C1704263|T121|659476|RXNORM|GREEN TEA EXTRACT|GREEN TEA EXTRACT
C0021234|T130|5775|RXNORM|INDOCYANINE GREEN|INDOCYANINE GREEN
C0062986|T195|27130|RXNORM|CEFPIROME|CEFPIROME
C2928546|T121|1007629|RXNORM|GARLIC PREPARATION / PARSLEY EXTRACT|GARLIC PREPARATION / PARSLEY EXTRACT
C2928545|T121|1007628|RXNORM|DEXAMETHASONE / DOBESILIC ACID / LIDOCAINE|DEXAMETHASONE / DOBESILIC ACID / LIDOCAINE
C3247610|T121|1192684|RXNORM|CHLOPHEDIANOL / PHENYLEPHRINE / PYRILAMINE|CHLOPHEDIANOL / PHENYLEPHRINE / PYRILAMINE
C2928540|T121|1007622|RXNORM|LIDOCAINE / TRIBENOSIDE|LIDOCAINE / TRIBENOSIDE
C2928539|T121|1007621|RXNORM|NIACINAMIDE / POTASSIUM IODIDE|NIACINAMIDE / POTASSIUM IODIDE
C2928538|T121|1007620|RXNORM|MICONAZOLE / TINIDAZOLE|MICONAZOLE / TINIDAZOLE
C2928544|T121|1007627|RXNORM|GARLIC PREPARATION / HAWTHORN PREPARATION|GARLIC PREPARATION / HAWTHORN PREPARATION
C2731508|T129|895495|RXNORM|DOG HAIR EXTRACT|DOG HAIR EXTRACT
C2928542|T121|1007625|RXNORM|BISMUTH SUBNITRATE / CERIUM OXALATE|BISMUTH SUBNITRATE / CERIUM OXALATE
C2193828|T121|1007624|RXNORM|AMOXICILLIN / BROVANEXINE|AMOXICILLIN / BROVANEXINE
C3505164|T109|1358002|RXNORM|SILYBUM MARIANUM SEED OIL|SILYBUM MARIANUM SEED OIL
C0971579|T121|306674|RXNORM|VARDENAFIL|VARDENAFIL
C0601893|T121|156075|RXNORM|VANILLYLAMINE|VANILLYLAMINE
C1875108|T121|691226|RXNORM|EPHEDRINE / GUAIFENESIN / PHENOBARBITAL / THEOPHYLLINE|EPHEDRINE / GUAIFENESIN / PHENOBARBITAL / THEOPHYLLINE
C2604572|T130|1428873|RXNORM|HC YELLOW NO. 5|HC YELLOW NO. 5
C3488428|T121|1426437|RXNORM|COD, UNSPECIFIED PREPARATION|COD, UNSPECIFIED PREPARATION
C3818730|T121|1534775|RXNORM|SIMMONDSIA CHINENSIS LEAF EXTRACT|SIMMONDSIA CHINENSIS LEAF EXTRACT
C0065093|T121|28817|RXNORM|LITHIUM SUCCINATE|LITHIUM SUCCINATE
C0065094|T197|28818|RXNORM|LITHIUM SULFATE|LITHIUM SULFATE
C3256673|T121|1307549|RXNORM|CYMBOPOGON CITRATUS LEAF EXTRACT|CYMBOPOGON CITRATUS LEAF EXTRACT
C2929347|T121|1008443|RXNORM|DEXTROMETHORPHAN / DIPHENHYDRAMINE / PHENYLEPHRINE|DEXTROMETHORPHAN / DIPHENHYDRAMINE / PHENYLEPHRINE
C3256490|T121|1307548|RXNORM|4-(P-HYDROXYPHENYL)-2-BUTANONE ACETATE|4-(P-HYDROXYPHENYL)-2-BUTANONE ACETATE
C0047821|T109|1546355|RXNORM|4,4'-DINITROCARBANILIDE|4,4'-DINITROCARBANILIDE
C3539986|T121|1428876|RXNORM|PETASITES FRAGRANS EXTRACT|PETASITES FRAGRANS EXTRACT
C1328071|T121|729596|RXNORM|METHOXY POLYETHYLENE GLYCOL-EPOETIN BETA|METHOXY POLYETHYLENE GLYCOL-EPOETIN BETA
C2183765|T121|817960|RXNORM|DIPYRONE / PRAMIVERINE|DIPYRONE / PRAMIVERINE
C0244104|T123|72031|RXNORM|PYRUVATE|PYRUVATE
C0914729|T121|279645|RXNORM|ALMOTRIPTAN|ALMOTRIPTAN
C3487967|T121|1342492|RXNORM|YUCCA FILAMENTOSA EXTRACT|YUCCA FILAMENTOSA EXTRACT
C0074770|T197|1293719|RXNORM|SODIUM SULFIDE|SODIUM SULFIDE
C0016945|T123|4626|RXNORM|GALACTOSE|GALACTOSE
C0000464|T123|73|RXNORM|SYNTHETIC LEVOTHYROXINE|DOCOSAHEXAENOATE
C0028066|T121|7417|RXNORM|NIFEDIPINE|NIFEDIPINE
C0028053|T121|7414|RXNORM|NICOTINYL ALCOHOL|NICOTINYL ALCOHOL (PYRIDYLCARBINOL)
C0028067|T121|7418|RXNORM|NIFLUMIC ACID|NIFLUMIC ACID
C0086728|T121|42826|RXNORM|OBIDOXIME|OBIDOXIME
C3645014|T121|1426286|RXNORM|AMYLASES / BROMELAINS / PAPAIN / PAPAYA PREPARATION|AMYLASES / BROMELAINS / PAPAIN / PAPAYA PREPARATION
C0526501|T121|135091|RXNORM|MOSAPRIDE|MOSAPRIDE
C3818696|T122|1536455|RXNORM|DECYL OLIVATE|DECYL OLIVATE
C0717565|T121|214368|RXNORM|CASCARA SAGRADA / MAGNESIUM HYDROXIDE|CASCARA SAGRADA / MAGNESIUM HYDROXIDE
C0717566|T121|214369|RXNORM|CASCARA SAGRADA / PHENOLPHTHALEIN|CASCARA SAGRADA / PHENOLPHTHALEIN
C3818823|T109|1489543|RXNORM|ANTIOXIDANT 119|ANTIOXIDANT 119
C3249516|T129|1232637|RXNORM|BROADLEAF CATTAIL POLLEN EXTRACT|TYPHA LATINFOLIA POLLEN EXTRACT
C3256124|T109|1307544|RXNORM|BLETILLA STRIATA BULB EXTRACT|BLETILLA STRIATA TUBER EXTRACT
C2727189|T129|1232630|RXNORM|TRAGACANTH ALLERGENIC EXTRACT|TRAGACANTH ALLERGENIC EXTRACT
C1873960|T121|689573|RXNORM|ACETAMINOPHEN / CAFFEINE / PHENYLPROPANOLAMINE / PYRILAMINE|ACETAMINOPHEN / CAFFEINE / PHENYLPROPANOLAMINE / PYRILAMINE
C1873959|T121|689572|RXNORM|ACETAMINOPHEN / CAFFEINE / ISOMETHEPTENE|ACETAMINOPHEN / CAFFEINE / ISOMETHEPTENE
C0143083|T125|56570|RXNORM|SOMATREM|SOMATREM
C1873957|T121|689570|RXNORM|ACETAMINOPHEN / CAFFEINE / GUAIFENESIN / PHENYLEPHRINE|ACETAMINOPHEN / CAFFEINE / GUAIFENESIN / PHENYLEPHRINE
C0041086|T121|10844|RXNORM|TRIOXSALEN|TRIOXSALEN
C1873962|T121|689576|RXNORM|ACETAMINOPHEN / CALCIUM CARBONATE|ACETAMINOPHEN / CALCIUM CARBONATE
C3205286|T121|1306883|RXNORM|BARLEY MALT SYRUP|BARLEY MALT SYRUP
C1873961|T121|689574|RXNORM|ACETAMINOPHEN / CAFFEINE / PHENYLPROPANOLAMINE / SALICYLAMIDE|ACETAMINOPHEN / CAFFEINE / PHENYLPROPANOLAMINE / SALICYLAMIDE
C3555537|T130|1373391|RXNORM|TECHNETIUM TC 99M TILMANOCEPT|TECHNETIUM TC 99M TILMANOCEPT
C0041098|T121|10849|RXNORM|TRIPROLIDINE|TRIPROLIDINE
C0041098|T121|10849|RXNORM|TRIPROLIDINE|TRIPROLIDINE
C1873964|T121|689579|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE|ACETAMINOPHEN / CHLORPHENIRAMINE / CODEINE / PHENYLEPHRINE
C0128811|T121|52853|RXNORM|MODIFIED FLUID GELATINS|MODIFIED FLUID GELATINS
C2369192|T130|1426748|RXNORM|IOBENGUANE I-123|IOBENGUANE I-123
C1720694|T121|645051|RXNORM|CALCIUM CARBONATE / SODIUM BICARBONATE|CALCIUM CARBONATE / SODIUM BICARBONATE
C3497859|T121|1426747|RXNORM|POLYGLYCERYL-10 LAURATE|POLYGLYCERYL-10 LAURATE
C0724613|T121|221113|RXNORM|LEVOROTATORY ALKALOIDS OF BELLADONNA|LEVOROTATORY ALKALOIDS OF BELLADONNA
C0754659|T121|228790|RXNORM|DUTASTERIDE|DUTASTERIDE
C0724603|T125|221110|RXNORM|ULTRALENTE INSULIN, HUMAN|ULTRALENTE INSULIN, HUMAN
C2722026|T129|891796|RXNORM|ASPARAGUS ALLERGENIC EXTRACT|ASPARAGUS OFFICINALIS ALLERGENIC EXTRACT
C1827476|T121|687089|RXNORM|ANTAZOLINE / XYLOMETAZOLINE|ANTAZOLINE / XYLOMETAZOLINE
C3472779|T109|1356144|RXNORM|ISOPROPYL TITANIUM TRIISOSTEARATE|ISOPROPYL TITANIUM TRIISOSTEARATE
C0207011|T121|67257|RXNORM|MYRRH EXTRACT|MYRRH EXTRACT
C2194108|T121|813567|RXNORM|FLAVOXATE / PROPYPHENAZONE|FLAVOXATE / PROPYPHENAZONE
C1095895|T121|319816|RXNORM|URTICA PREPARATION|URTICA PREPARATION
C3663711|T121|1433634|RXNORM|ADENOSINE / NIACINAMIDE|ADENOSINE / NIACINAMIDE
C0771693|T121|236421|RXNORM|MEFENIDRAMIUM|MEFENIDRAMIUM
C0018513|T121|5084|RXNORM|HALCINONIDE|HALCINONIDE
C1113412|T121|324054|RXNORM|MIXED VESPID VENOM PROTEIN|MIXED VESPID VENOM PROTEIN
C2740288|T129|898404|RXNORM|ANNUAL BLUEGRASS POLLEN EXTRACT|POA ANNUA POLLEN EXTRACT
C3486570|T121|1340182|RXNORM|TRIFOLIUM PRATENSE POLLEN EXTRACT|TRIFOLIUM PRATENSE POLLEN EXTRACT
C1875646|T121|689741|RXNORM|PHENIRAMINE / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE / PYRILAMINE|PHENIRAMINE / PHENYLPROPANOLAMINE / PHENYLTOLOXAMINE / PYRILAMINE
C0216231|T129|69634|RXNORM|SARGRAMOSTIM|SARGRAMOSTIM
C2697961|T121|1425099|RXNORM|TRAMETINIB|TRAMETINIB
C3488472|T121|1340185|RXNORM|LILIUM LANCIFOLIUM WHOLE FLOWERING EXTRACT|LILIUM LANCIFOLIUM WHOLE FLOWERING EXTRACT
C0008168|T195|2348|RXNORM|CHLORAMPHENICOL|CHLORAMPHENICOL
C0008168|T195|2348|RXNORM|CHLORAMPHENICOL|CHLORAMPHENICOL
C0008168|T195|2348|RXNORM|CHLORAMPHENICOL|CHLORAMPHENICOL
C0008168|T195|2348|RXNORM|CHLORAMPHENICOL|CHLORAMPHENICOL
C2701463|T129|852268|RXNORM|RED OAK POLLEN EXTRACT|QUERCUS RUBRA POLLEN EXTRACT
C2928999|T121|1008091|RXNORM|ASCORBIC ACID / HYALURONATE|ASCORBIC ACID / HYALURONATE
C2928998|T121|1008090|RXNORM|FERROUS FUMARATE / POLYSACCHARIDE IRON COMPLEX|FERROUS FUMARATE / POLYSACCHARIDE IRON COMPLEX
C2929001|T121|1008093|RXNORM|CARBOXYMETHYLCELLULOSE / HYPROMELLOSE|CARBOXYMETHYLCELLULOSE / HYPROMELLOSE
C2929000|T121|1008092|RXNORM|BROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE|BROMPHENIRAMINE / DEXTROMETHORPHAN / PHENYLEPHRINE
C2929003|T121|1008095|RXNORM|BACITRACIN / HYDROCORTISONE / NEOMYCIN|BACITRACIN / HYDROCORTISONE / NEOMYCIN
C2929002|T121|1008094|RXNORM|CLINDAMYCIN / GLUCOSE|CLINDAMYCIN / GLUCOSE
C1172566|T121|354606|RXNORM|EMODEPSIDE|EMODEPSIDE
C3856084|T197|1549555|RXNORM|BARIUM IODATE|BARIUM IODATE
C2929007|T121|1008099|RXNORM|BOVINE CARTILAGE EXTRACT / SHARK CARTILAGE EXTRACT|BOVINE CARTILAGE EXTRACT / SHARK CARTILAGE EXTRACT
C2929006|T121|1008098|RXNORM|DOXYLAMINE / PSEUDOEPHEDRINE|DOXYLAMINE / PSEUDOEPHEDRINE
C3818755|T109|1492942|RXNORM|TALL OIL ACID|TALL OIL ACID
C3818754|T121|1492943|RXNORM|BOLETUS LURIDUS FRUITING BODY EXTRACT|BOLETUS LURIDUS FRUITING BODY EXTRACT
C3818753|T109|1492944|RXNORM|CALCIUM-SODIUM MALEATE METHYL VINYL ETHER COPOLYMER (1000000 MW, 1900 MPA.S AT 11%)|CALCIUM-SODIUM MALEATE METHYL VINYL ETHER COPOLYMER (1000000 MW, 1900 MPA.S AT 11%)
C0303611|T130|90650|RXNORM|TECHNETIUM 99M|TECHNETIUM 99M
C1445716|T121|466482|RXNORM|PAPAIN / UREA|PAPAIN / UREA
C0066966|T121|1438530|RXNORM|MUSK KETONE|MUSK KETONE
C2586675|T121|1433887|RXNORM|CHOLINE FENOFIBRATE|CHOLINE FENOFIBRATE
C1445720|T121|466486|RXNORM|DEXTROMETHORPHAN / PHENYLEPHRINE|DEXTROMETHORPHAN / PHENYLEPHRINE
C1445721|T121|466487|RXNORM|PHENIRAMINE / PHENYLEPHRINE|PHENIRAMINE / PHENYLEPHRINE
C1445721|T121|466487|RXNORM|PHENIRAMINE / PHENYLEPHRINE|PHENIRAMINE / PHENYLEPHRINE
C1445721|T121|466487|RXNORM|PHENIRAMINE / PHENYLEPHRINE|PHENIRAMINE / PHENYLEPHRINE
C1445723|T121|466489|RXNORM|CODEINE / GUAIFENESIN / PSEUDOEPHEDRINE|CODEINE / GUAIFENESIN / PSEUDOEPHEDRINE
C1446539|T121||RXNORM|TEGAFUR / URACIL
C0981883|T129|901299|RXNORM|WHOLE WHEAT ALLERGENIC EXTRACT|WHOLE WHEAT ALLERGENIC EXTRACT
C0002406|T131|1433189|RXNORM|AMARANTH DYE|AMARANTH DYE
C2016762|T121|818288|RXNORM|SODIUM BICARBONATE / SODIUM PHOSPHATE|SODIUM BICARBONATE / SODIUM PHOSPHATE
C0006657|T127|1889|RXNORM|CALCIFEDIOL|CALCIFEDIOL
C0051570|T121|17665|RXNORM|AMEZINIUM|AMEZINIUM
C0006644|T121|1886|RXNORM|CAFFEINE|CAFFEINE
C2741480|T129|901291|RXNORM|VANILLA BEAN ALLERGENIC EXTRACT|VANILLA BEAN ALLERGENIC EXTRACT
C0013340|T125|3706|RXNORM|DYDROGESTERONE|DYDROGESTERONE
C3495102|T121|1330284|RXNORM|ACONITUM NAPELLUS ROOT EXTRACT|ACONITUM NAPELLUS ROOT EXTRACT
C0981840|T129|314324|RXNORM|ASPERGILLUS TERREUS ALLERGENIC EXTRACT|ASPERGILLUS TERREUS ALLERGENIC EXTRACT
C2701576|T129|852419|RXNORM|BEECH POLLEN EXTRACT|FAGUS GRANDIFOLIA POLLEN EXTRACT
C3268278|T121|1306882|RXNORM|REDROOT PIGWEED WHOLE ALLERGENIC EXTRACT|AMARANTHUS RETROFLEXUS WHOLE ALLERGENIC EXTRACT
C0007710|T121|2228|RXNORM|MECLOFENOXATE|MECLOFENOXATE
C0017890|T123|4919|RXNORM|GLYCINE|GLYCINE
C0007343|T121|2129|RXNORM|CASTOR OIL|CASTOR OIL
C0017887|T121|4917|RXNORM|NITROGLYCERIN|NITROGLYCERIN
C0017887|T121|4917|RXNORM|NITROGLYCERIN|NITROGLYCERIN
C3530452|T109|1364406|RXNORM|MALPIGHIA GLABRA FRUIT EXTRACT|MALPIGHIA GLABRA FRUIT EXTRACT
C3152868|T129|1098232|RXNORM|LITTLESEED CANARY GRASS POLLEN EXTRACT|PHALARIS MINOR POLLEN EXTRACT
C0017861|T123|4910|RXNORM|GLYCERIN|GLYCERIN
C0017861|T123|4910|RXNORM|GLYCERIN|GLYCERIN
C0017861|T123|4910|RXNORM|GLYCERIN|GLYCERIN
C0017861|T123|4910|RXNORM|GLYCERIN|GLYCERIN
C0017861|T123|4910|RXNORM|GLYCERIN|GLYCERIN
C0017861|T123|4910|RXNORM|GLYCERIN|GLYCERIN
C2927846|T121|1006922|RXNORM|LIDOCAINE / PHENOL|LIDOCAINE / PHENOL
C2929796|T121|1008899|RXNORM|MALACHITE GREEN / METRONIDAZOLE / MICROCRYSTALLINE CELLULOSE / TRICHLORFON|MALACHITE GREEN / METRONIDAZOLE / MICROCRYSTALLINE CELLULOSE / TRICHLORFON
C2929795|T121|1008898|RXNORM|POLYETHYLENE GLYCOL 400 / TETRAHYDROZOLINE|POLYETHYLENE GLYCOL 400 / TETRAHYDROZOLINE
C0004924|T122|1356|RXNORM|BEESWAX|BEESWAX
C2929788|T121|1008891|RXNORM|DAPSONE / ISONIAZID / PROTHIONAMIDE|DAPSONE / ISONIAZID / PROTHIONAMIDE
C0071972|T121|34482|RXNORM|CILASTATIN / IMIPENEM|CILASTATIN / IMIPENEM
C2929790|T121|1008893|RXNORM|ACETAMINOPHEN / CHLORPHENIRAMINE / DIPHENHYDRAMINE / PSEUDOEPHEDRINE|ACETAMINOPHEN / CHLORPHENIRAMINE / DIPHENHYDRAMINE / PSEUDOEPHEDRINE
C2929789|T121|1008892|RXNORM|CHONDROITIN SULFATES / HYALURONATE|CHONDROITIN SULFATES / HYALURONATE
C2929792|T121|1008895|RXNORM|DEXCHLORPHENIRAMINE / GUAIFENESIN / HYDROCODONE / PHENYLEPHRINE|DEXCHLORPHENIRAMINE / GUAIFENESIN / HYDROCODONE / PHENYLEPHRINE
C2929791|T121|1008894|RXNORM|OXYQUINOLINE / TETRACAINE|OXYQUINOLINE / TETRACAINE
C2929794|T121|1008897|RXNORM|BENDROFLUMETHIAZIDE / RAUWOLFIA PREPARATION|BENDROFLUMETHIAZIDE / RAUWOLFIA PREPARATION
C3538506|T121|1372932|RXNORM|RHODIOLA CRENULATA ROOT EXTRACT|RHODIOLA CRENULATA ROOT EXTRACT
C3538507|T121|1372933|RXNORM|PEG-20 SORBITAN ISOSTEARATE|PEG-20 SORBITAN ISOSTEARATE
C3538505|T109|1372930|RXNORM|CATALINA PREPARATION|CATALINA PREPARATION
C1509773|T121|1372931|RXNORM|STEARALKONIUM HECTORITE|STEARALKONIUM HECTORITE
C0357084|T197|105673|RXNORM|SODIUM IRONEDETATE|SODIUM FEREDETATE
C3538509|T121|1372935|RXNORM|SODIUM TRIDECETH SULFATE|SODIUM TRIDECETH SULFATE
C0085845|T123|42543|RXNORM|ASPARTATE|ASPARTATE
C0772389|T121|1367109|RXNORM|STARCH, WHEAT|STARCH, WHEAT
C3535684|T109|1368339|RXNORM|PHRAGMITES AUSTRALIS WHOLE EXTRACT|PHRAGMITES AUSTRALIS WHOLE EXTRACT
C3535685|T109|1368338|RXNORM|PHOENIX DACTYLIFERA SEED EXTRACT|PHOENIX DACTYLIFERA SEED EXTRACT
C3535670|T109|1368621|RXNORM|HUMAN ADIPOSE PREPARATION|HUMAN ADIPOSE PREPARATION
C3535687|T109|1368332|RXNORM|HELIANTHUS ANNUUS SPROUT EXTRACT|HELIANTHUS ANNUUS SPROUT EXTRACT
C3535688|T109|1368331|RXNORM|COMMIPHORA MADAGASCARIENSIS RESIN EXTRACT|COMMIPHORA MADAGASCARIENSIS RESIN
C3651699|T121|1431993|RXNORM|METHYL LACTATE, L-|METHYL LACTATE, L-
C3535686|T109|1368337|RXNORM|PETASITES JAPONICUS ROOT EXTRACT|PETASITES JAPONICUS ROOT EXTRACT
C3692546|T121|1442198|RXNORM|CAMELLIA SINENSIS VAR. ASSAMICA WHOLE EXTRACT|CAMELLIA SINENSIS VAR. ASSAMICA WHOLE EXTRACT
C1874359|T121|689507|RXNORM|ASPIRIN / BUTALBITAL / CAFFEINE / PHENACETIN|ASPIRIN / BUTALBITAL / CAFFEINE / PHENACETIN
C3486591|T121|1309776|RXNORM|CLEMATIS VIRGINIANA TOP|CLEMATIS VIRGINIANA TOP
C2928405|T121|1007483|RXNORM|DEXAMETHASONE / HYPROMELLOSE|DEXAMETHASONE / HYPROMELLOSE
C3486590|T121|1309774|RXNORM|CLEMATIS RECTA FLOWERING TOP EXTRACT|CLEMATIS RECTA FLOWERING TOP EXTRACT
C3489212|T121|1309775|RXNORM|CALENDULA OFFICINALIS FLOWERING TOP EXTRACT|CALENDULA OFFICINALIS FLOWERING TOP EXTRACT
C3486857|T121|1309772|RXNORM|CITRULLUS COLOCYNTHIS FRUIT PULP EXTRACT|CITRULLUS COLOCYNTHIS FRUIT PULP EXTRACT
C3486588|T121|1309770|RXNORM|AESCULUS CARNEA FLOWER EXTRACT|AESCULUS CARNEA FLOWER EXTRACT
C3489011|T121|1309771|RXNORM|CINCHONA OFFICINALIS BARK EXTRACT|CINCHONA OFFICINALIS BARK EXTRACT
C0393022|T129|121191|RXNORM|RITUXIMAB|RITUXIMAB
C0023870|T196|6448|RXNORM|LITHIUM|LITHIUM
C1874357|T121|689502|RXNORM|ALUMINUM HYDROXIDE / ASPIRIN / CALCIUM CARBONATE / MAGNESIUM HYDROXIDE|ALUMINUM HYDROXIDE / ASPIRIN / CALCIUM CARBONATE / MAGNESIUM HYDROXIDE
C3474174|T121|1300367|RXNORM|BORDETELLA PERTUSSIS FILAMENTOUS HEMAGGLUTININ VACCINE, INACTIVATED / BORDETELLA PERTUSSIS PERTACTIN VACCINE, INACTIVATED / BORDETELLA PERTUSSIS TOXOID VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED|BORDETELLA PERTUSSIS FILAMENTOUS HEMAGGLUTININ VACCINE, INACTIVATED / BORDETELLA PERTUSSIS PERTACTIN VACCINE, INACTIVATED / BORDETELLA PERTUSSIS TOXOID VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / TETANUS TOXOID VACCINE, INACTIVATED
C3256126|T196|1424875|RXNORM|BORATE ION|BORATE ION
C3256801|T109|1424874|RXNORM|PPG-5-CETETH-20|PPG-5-CETETH-20
C3256207|T109|1424877|RXNORM|CUCUMARIA FRONDOSA PREPARATION|CUCUMARIA FRONDOSA PREPARATION
C0665917|T109|1424876|RXNORM|CITRONELLAL|CITRONELLAL
C3486551|T121|1344641|RXNORM|CONVALLARIA MAJALIS EXTRACT|CONVALLARIA MAJALIS EXTRACT
C3695954|T109|1484500|RXNORM|C11-13 PARETH-6|C11-13 PARETH-6
C0358787|T121|619749|RXNORM|BENSERAZIDE / LEVODOPA|BENSERAZIDE / LEVODOPA
C3255932|T109|1424878|RXNORM|DIAMOND TURBOT EXTRACT|DIAMOND FLOUNDER EXTRACT
C3486741|T121|1344643|RXNORM|SAMBUCUS NIGRA FLOWER EXTRACT|SAMBUCUS NIGRA FLOWER EXTRACT
C3486555|T129|1344642|RXNORM|INFLUENZA A-B VIRUS IMMUNOSERUM RABBIT|INFLUENZA A-B VIRUS IMMUNOSERUM RABBIT
C0083183|T126|41397|RXNORM|LACTASE|TILACTASE
C3700869|T121|1487162|RXNORM|ALPHA-BISABOLOL, (+)-|ALPHA-BISABOLOL, (+)-
C0074747|T197|36699|RXNORM|SODIUM MOLYBDATE(VI)|SODIUM MOLYBDATE(VI)
C0874067|T121|260040|RXNORM|EVENING PRIMROSE EXTRACT|OENOTHERA BIENNIS
C0074744|T197|36696|RXNORM|SODIUM METABISULFITE|SODIUM METABISULFITE
C0027396|T121|7258|RXNORM|NAPROXEN|NAPROXEN
C0027396|T121|7258|RXNORM|NAPROXEN|NAPROXEN
C0699817|T121|202912|RXNORM|INTERFERON ALFA-N1|INTERFERON ALFA-N1
C2927933|T121|1007010|RXNORM|METHYCLOTHIAZIDE / TRIAMTERENE|METHYCLOTHIAZIDE / TRIAMTERENE
C0025684|T123|6854|RXNORM|METHOXSALEN|METHOXSALEN
C0025684|T123|6854|RXNORM|METHOXSALEN|METHOXSALEN
C2927935|T121|1007012|RXNORM|PANTOTHENATE / RIBOFLAVIN / VITAMIN B6|PANTOTHENATE / RIBOFLAVIN / VITAMIN B6
C2927936|T121|1007013|RXNORM|CHLORHEXIDINE / MURAMIDASE / TETRACAINE|CHLORHEXIDINE / MURAMIDASE / TETRACAINE
C2927937|T121|1007014|RXNORM|MAGNESIUM CITRATE / MAGNESIUM GLUCONATE|MAGNESIUM CITRATE / MAGNESIUM GLUCONATE
C2927938|T121|1007015|RXNORM|ESTROPIPATE / MEDROXYPROGESTERONE|ESTROPIPATE / MEDROXYPROGESTERONE
C0025681|T121|6853|RXNORM|METHOXAMINE|METHOXAMINE
C0025678|T121|6852|RXNORM|METHOTRIMEPRAZINE|METHOTRIMEPRAZINE
C2927941|T121|1007018|RXNORM|CLORAZEPIC ACID / DOMPERIDONE|CLORAZEPIC ACID / DOMPERIDONE
C2927942|T121|1007019|RXNORM|CINNARIZINE / XANTHINOL|CINNARIZINE / XANTHINOL
C3864838|T121|1596141|RXNORM|HYDROXYPROPYL CELLULOSE (TYPE G)|HYDROXYPROPYL CELLULOSE (TYPE G)
C2701419|T129|852221|RXNORM|SHAGBARK HICKORY POLLEN EXTRACT|SHAGBARK HICKORY POLLEN EXTRACT
C3257522|T121|1309369|RXNORM|COTTON SEED EXTRACT|COTTON SEED EXTRACT
C2827306|T121|1309368|RXNORM|POLYETHYELENE GLYCOL 7000|POLYETHYELENE GLYCOL 7000
C3488932|T109|1309365|RXNORM|PEG-20 GLYCERYL STEARATE|PEG-20 GLYCERYL STEARATE
C3488974|T109|1309364|RXNORM|KUKUI NUT OIL|KUKUI NUT OIL
C3488933|T121|1309367|RXNORM|PEG-6 STEARATE|PEG-6 STEARATE
C3281577|T121|1309366|RXNORM|PEG-32 STEARATE|PEG-32 STEARATE
C3256025|T121|1309361|RXNORM|CNIDIUM SEED EXTRACT|CNIDIUM SEED EXTRACT
C3265865|T109|1309360|RXNORM|HYDROGENATED PALM KERNEL OIL|HYDROGENATED PALM KERNEL OIL
C0982311|T109|1309363|RXNORM|PEG-120 METHYL GLUCOSE DIOLEATE|PEG-120 METHYL GLUCOSE DIOLEATE
C2343923|T121|797426|RXNORM|NAPROXEN / SUMATRIPTAN|NAPROXEN / SUMATRIPTAN
C1874805|T121|689379|RXNORM|CHLORPHENIRAMINE / CODEINE / IODINATED GLYCEROL|CHLORPHENIRAMINE / CODEINE / IODINATED GLYCEROL
C0982005|T129|314488|RXNORM|CORN SMUT ALLERGENIC EXTRACT|USTILAGO MAYDIS ALLERGENIC EXTRACT
C0068334|T121|31448|RXNORM|ALLERGENIC EXTRACT,LYCOPERDON PYRIFORME|NABUMETONE
C0068334|T121|31448|RXNORM|ALLERGENIC EXTRACT,PENICILLIUM FREQUENTANS|NABUMETONE
C1874638|T121|690837|RXNORM|CALAMINE / DIPHENHYDRAMINE|CALAMINE / DIPHENHYDRAMINE
C0068334|T121|31448|RXNORM|ALLERGENIC EXTRACT,COPRINUS MICACEUS|NABUMETONE
C1874801|T121|689374|RXNORM|CHLOROXYLENOL / PRAMOXINE|CHLOROXYLENOL / PRAMOXINE
C0068334|T121|31448|RXNORM|ALLERGENIC EXTRACT,CALVATIA CYATHIFORMIS|NABUMETONE
C3486131|T121|1311319|RXNORM|PORK COLLAGEN PREPARATION|PORCINE COLLAGEN PREPARATION
C3486763|T121|1311318|RXNORM|LONICERA XYLOSTEUM FRUIT EXTRACT|LONICERA XYLOSTEUM FRUIT EXTRACT
C3486782|T121|1311315|RXNORM|SUS SCROFA CAPILLARY TISSUE PREPARATION|PORCINE CAPILLARY TISSUE PREPARATION
C3486630|T197|1311314|RXNORM|FERRIC PICRATE PREPARATION|FERRIC PICRATE PREPARATION
C3486785|T121|1311317|RXNORM|SUS SCROFA CEREBRAL CORTEX PREPARATION|PORCINE CEREBRAL CORTEX PREPARATION
C3486784|T121|1311316|RXNORM|SUS SCROFA CEREBELLUM PREPARATION|PORCINE CEREBELLUM PREPARATION
C2347679|T121|1311310|RXNORM|PRIMULA VERIS EXTRACT|PRIMULA VERIS EXTRACT
C0074741|T197|1311313|RXNORM|SODIUM HYPOPHOSPHITE|SODIUM HYPOPHOSPHITE
C0024477|T197|6582|RXNORM|MAGNESIUM OXIDE|MAGNESIUM OXIDE
C0024476|T197|6581|RXNORM|MAGNESIUM HYDROXIDE|MAGNESIUM HYDROXIDE
C0024476|T197|6581|RXNORM|MAGNESIUM HYDROXIDE|MAGNESIUM HYDROXIDE
C0078811|T121|39969|RXNORM|ZIPEPROL|ZIPEPROL
C0033439|T121|8758|RXNORM|PROPANIDID|PROPANIDID
C0024480|T197|6585|RXNORM|MAGNESIUM SULFATE|MAGNESIUM SULFATE
C0024480|T197|6585|RXNORM|MAGNESIUM SULFATE|MAGNESIUM SULFATE
C0024480|T197|6585|RXNORM|MAGNESIUM SULFATE|MAGNESIUM SULFATE
C0071808|T121|34345|RXNORM|PRALIDOXIME|PRALIDOXIME
C0071810|T121|34347|RXNORM|PRAMOXINE|PRAMOXINE
C0071810|T121|34347|RXNORM|PRAMOXINE|PRAMOXINE
C0071810|T121|34347|RXNORM|PRAMOXINE|PRAMOXINE
C0028906|T168|7624|RXNORM|CLOVE OIL|CLOVE OIL
C0028902|T195|7623|RXNORM|OFLOXACIN|OFLOXACIN
C0028902|T195|7623|RXNORM|OFLOXACIN|OFLOXACIN
C0028902|T195|7623|RXNORM|OFLOXACIN|OFLOXACIN
C2726203|T129|971198|RXNORM|PLEOSPORA HERBARUM EXTRACT|PLEOSPORA HERBARUM EXTRACT
C0028923|T195|7629|RXNORM|OLEANDOMYCIN|OLEANDOMYCIN
C0077138|T109|1426368|RXNORM|TRIISOPROPANOLAMINE|TRIISOPROPANOLAMINE
C2927648|T129|1006495|RXNORM|INDIAN WORMWOOD SAGE POLLEN EXTRACT|ARTEMISIA DRACUNCULUS POLLEN EXTRACT
C0993223|T125|317598|RXNORM|NPH INSULIN, BEEF-PORK|INSULIN BEEF-PORK, ISOPHANE
C1874906|T121|690096|RXNORM|CODEINE / POTASSIUM CITRATE|CODEINE / POTASSIUM CITRATE
C3834170|T121|1543095|RXNORM|FACTOR VIII (B-DOMAIN DELETED RECOMBINANT) FC FUSION PROTEIN|(1-743)-(1638-2332)-BLOOD-COAGULATION FACTOR VIII (SYNTHETIC HUMAN) FUSION PROTEIN WITH IMMUNOGLOBULIN G1 (SYNTHETIC HUMAN FC DOMAIN FRAGMENT), (1444-6'),(1447-9')-BIS(DISULFIDE) WITH IMMUNOGLOBULIN G1 (SYNTHETIC HUMAN FC DOMAIN FRAGMENT)
C1874905|T121|690095|RXNORM|CODEINE / PHENYLPROPANOLAMINE / PROMETHAZINE|CODEINE / PHENYLPROPANOLAMINE / PROMETHAZINE
C1874904|T121|690093|RXNORM|CODEINE / PHENYLEPHRINE / PSEUDOEPHEDRINE|CODEINE / PHENYLEPHRINE / PSEUDOEPHEDRINE
C1656322|T121|1314363|RXNORM|ETHYLENE BRASSYLATE|ETHYLENE BRASSYLATE
C0015075|T121|1314362|RXNORM|ETHYLENE|ETHYLENE
C0059779|T121|1314361|RXNORM|ETHYL OLEATE|ETHYL OLEATE
C0732093|T121|226623|RXNORM|FACTOR VIII / VON WILLEBRAND FACTOR|FACTOR VIII / VON WILLEBRAND FACTOR
C0732093|T121|226623|RXNORM|FACTOR VIII / VON WILLEBRAND FACTOR|FACTOR VIII / VON WILLEBRAND FACTOR
C0069963|T109|1314367|RXNORM|PALMATINE|PALMATINE
C0065641|T197|1314366|RXNORM|MANGANESE CARBONATE|MANGANESE CARBONATE
C0046088|T130|1314365|RXNORM|2-ETHOXYETHANOL|2-ETHOXYETHANOL
C0015083|T131|1314364|RXNORM|ETHYLENE GLYCOL|ETHYLENE GLYCOL
C3486637|T121|1309940|RXNORM|FALLOPIA MULTIFLORA ROOT EXTRACT|REYNOUTRIA MULTIFLORA ROOT EXTRACT
C3486639|T121|1309943|RXNORM|ARNICA ANGUSTIFOLIA FLOWER EXTRACT|ARNICA ANGUSTIFOLIA FLOWER EXTRACT
C3282119|T121|1309942|RXNORM|PLANTAGO OVATA SEED EXTRACT|PLANTAGO OVATA SEED EXTRACT
C3486645|T121|1309947|RXNORM|ARNICA MONTANA ROOT EXTRACT|ARNICA MONTANA ROOT EXTRACT
C3486640|T121|1309946|RXNORM|MIMULUS GUTTATUS FLOWERING TOP EXTRACT|MIMULUS GUTTATUS FLOWERING TOP EXTRACT
C0072225|T121|34693|RXNORM|PROPYLENE GLYCOL|PROPYLENE GLYCOL
C0072225|T121|34693|RXNORM|PROPYLENE GLYCOL|PROPYLENE GLYCOL
C3486649|T121|1309948|RXNORM|QUILLAJA SAPONARIA BARK EXTRACT|QUILLAJA SAPONARIA BARK EXTRACT
C0001480|T123|318|RXNORM|ADENOSINE TRIPHOSPHATE|ADENOSINE TRIPHOSPHATE
C0077126|T121|38655|RXNORM|TRIFLUSAL|TRIFLUSAL
C0037512|T197|9876|RXNORM|GOLD SODIUM THIOSULFATE|SODIUM AUROTIOSULFATE
C3541373|T123|9152|RXNORM|RAUWOLFIA ALKALOIDS|RAUWOLFIA ALKALOIDS
C0037508|T197|9873|RXNORM|SODIUM FLUORIDE|SODIUM FLUORIDE
C0037508|T197|9873|RXNORM|SODIUM FLUORIDE|SODIUM FLUORIDE
C0037508|T197|9873|RXNORM|SODIUM FLUORIDE|SODIUM FLUORIDE
C2929464|T121|1008561|RXNORM|ACETAMINOPHEN / NAPROXEN|ACETAMINOPHEN / NAPROXEN
C2929463|T121|1008560|RXNORM|BISMUTH CAMPHOCARBONATE / GUAIFENESIN|BISMUTH CAMPHOCARBONATE / GUAIFENESIN
C2929466|T121|1008563|RXNORM|ASAFETIDA EXTRACT / CASCARA SAGRADA|ASAFETIDA EXTRACT / CASCARA SAGRADA
C2929465|T121|1008562|RXNORM|ALLANTOIN / SULFADIAZINE|ALLANTOIN / SULFADIAZINE
C2929468|T121|1008565|RXNORM|LACTATE / SALICYLIC ACID|LACTATE / SALICYLIC ACID
C2929467|T121|1008564|RXNORM|METHYLENE BLUE / NAPHAZOLINE|METHYLENE BLUE / NAPHAZOLINE
C2929470|T121|1008567|RXNORM|CHONDROITIN SULFATES / GLUCOSAMINE|CHONDROITIN SULFATES / GLUCOSAMINE
C2929469|T121|1008566|RXNORM|BENZOCAINE / EPHEDRINE|BENZOCAINE / EPHEDRINE
C2929472|T121|1008569|RXNORM|LIDOCAINE / RIFAMYCIN SV|LIDOCAINE / RIFAMYCIN SV
C2929471|T121|1008568|RXNORM|BENZOCAINE / MAGNESIUM SULFATE|BENZOCAINE / MAGNESIUM SULFATE
C0059760|T121|24513|RXNORM|ETHYL CYSTEINE|ETHYL CYSTEINE
C1572766|T121|1368185|RXNORM|OCTOXYNOL-1|OCTOXYNOL-1
C1827175|T121|687113|RXNORM|CAFFEINE / GLUCOSE|CAFFEINE / GLUCOSE
C1533505|T121|477379|RXNORM|ECHINACEA ROOT EXTRACT|ECHINACEA ROOT EXTRACT
C1720719|T121|690329|RXNORM|RESORCINOL / SULFUR|RESORCINOL / SULFUR
C2073917|T121|815347|RXNORM|CHLORPROMAZINE / DIPYRONE|CHLORPROMAZINE / DIPYRONE
C3537698|T109|1371320|RXNORM|MENTHOL 1-PROPYLENE GLYCOL CARBONATE, (-)-|MENTHOL 1-PROPYLENE GLYCOL CARBONATE, (-)-
C3857936|T121|1591919|RXNORM|TURNERA DIFFUSA LEAF EXTRACT|TURNERA DIFFUSA LEAF EXTRACT
C3537699|T121|1371321|RXNORM|POLYQUATERNIUM-16 (N-VINYLPYRROLIDINONE:3-METHYL-1-VINYLIMIDAZOLIUM CHLORIDE (5:5))|POLYQUATERNIUM-16 (N-VINYLPYRROLIDINONE:3-METHYL-1-VINYLIMIDAZOLIUM CHLORIDE (5:5))
C3857474|T121|1591911|RXNORM|CHLORELLA PYRENOIDOSA EXTRACT|CHLORELLA PYRENOIDOSA EXTRACT
C3864966|T121|1591913|RXNORM|RICINOLEAMIDOPROPYLTRIMONIUM|RICINOLEAMIDOPROPYLTRIMONIUM
C2725894|T129|895542|RXNORM|HOG HAIR EXTRACT|SUS SCROFA HAIR EXTRACT
C3854017|T121|1591914|RXNORM|SPANISH SARDINE PREPARATION|SPANISH SARDINE PREPARATION
C0079349|T123|1591916|RXNORM|FIBROBLAST GROWTH FACTOR-1|FIBROBLAST GROWTH FACTOR-1
C1966117|T121|745526|RXNORM|CHLOROPHYLLIN COPPER COMPLEX / PAPAIN / UREA|CHLOROPHYLLIN COPPER COMPLEX / PAPAIN / UREA
C3856158|T121|1549697|RXNORM|RIBES NIGRUM FLOWER BUD EXTRACT|RIBES NIGRUM FLOWER BUD EXTRACT
C0612303|T109|1442197|RXNORM|OCTENYL SUCCINATE|OCTENYL SUCCINATE
C3855137|T109|1547469|RXNORM|SPARGANIUM STOLONIFERIUM WHOLE EXTRACT|SPARGANIUM STOLONIFERIUM WHOLE EXTRACT
C0076733|T197|38323|RXNORM|TITANIUM DIOXIDE|TITANIUM DIOXIDE
C0075504|T195|37320|RXNORM|SULFABENZAMIDE|SULFABENZAMIDE
C3535695|T109|1367687|RXNORM|ZANTHOXYLUM BUNGEANUM FRUIT RIND EXTRACT|ZANTHOXYLUM BUNGEANUM FRUIT RIND EXTRACT
C3281530|T121|1322526|RXNORM|PERSIMMON EXTRACT|PERSIMMON EXTRACT
C0042682|T121|11204|RXNORM|VINDESINE|VINDESINE
C0009979|T130|1366888|RXNORM|COPPER EDTA|COPPER EDTA
C0991877|T121|1426352|RXNORM|STEARETH-2|STEARETH-2
C3256438|T109|1426353|RXNORM|STEARIC MONOETHANOLAMIDE|STEARIC MONOETHANOLAMIDE
C3486705|T121|1313750|RXNORM|GERANIUM ROBERTIANUM EXTRACT|GERANIUM ROBERTIANUM EXTRACT
C2940204|T129|1014762|RXNORM|BALSAM POPLAR POLLEN EXTRACT|BALSAM POPLAR POLLEN EXTRACT
C0248347|T121|73409|RXNORM|CALCIUM CITRATE MALATE|CALCIUM CITRATE MALATE
C2940207|T129|1014766|RXNORM|JERUSALEM OAK POLLEN EXTRACT|CHENOPODIUM BOTRYS POLLEN EXTRACT
C3669001|T121|1485120|RXNORM|SENECIO VULGARIS EXTRACT|SENECIO VULGARIS EXTRACT
C2929057|T121|1008150|RXNORM|BENZYL ALCOHOL / CAMPHOR / MENTHOL|BENZYL ALCOHOL / CAMPHOR / MENTHOL
C1874010|T121|690204|RXNORM|ACETIC ACID / OXYQUINOLINE|ACETIC ACID / OXYQUINOLINE
C2929059|T121|1008152|RXNORM|TRICLOSAN / UNDECYLENATE|TRICLOSAN / UNDECYLENATE
C2929060|T121|1008153|RXNORM|BIOTIN / FOLIC ACID / MAGNESIUM OXIDE / PANTOTHENATE / VITAMIN A / VITAMIN E|BIOTIN / FOLIC ACID / MAGNESIUM OXIDE / PANTOTHENATE / VITAMIN A / VITAMIN E
C2929061|T121|1008154|RXNORM|BENZETHONIUM / EPINEPHRINE|BENZETHONIUM / EPINEPHRINE
C0060462|T121|25082|RXNORM|FLOPROPIONE|FLOPROPIONE
C2929063|T121|1008156|RXNORM|LYSINE / NIACINAMIDE / THIAMINE|LYSINE / NIACINAMIDE / THIAMINE
C2929064|T121|1008157|RXNORM|ACETAMINOPHEN / ALUMINUM ACETATE / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE|ACETAMINOPHEN / ALUMINUM ACETATE / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE
C2929065|T121|1008158|RXNORM|CARBON DIOXIDE / HELIUM / HYDROGEN / NITROGEN / OXYGEN|CARBON DIOXIDE / HELIUM / HYDROGEN / NITROGEN / OXYGEN
C3530614|T121|1364950|RXNORM|MEADOWFOAMAMIDOPROPYL BETAINE|MEADOWFOAMAMIDOPROPYL BETAINE
C2825689|T121|1420978|RXNORM|PYRITIDIUM|PYRITIDIUM
C3555465|T197|1420979|RXNORM|SCHORL TOURMALINE|SCHORL TOURMALINE
C0676547|T197|195983|RXNORM|CALCIUM BROMIDE|CALCIUM BROMIDE
C2756533|T129|968475|RXNORM|OAT LOOSE SMUT EXTRACT|OAT LOOSE SMUT EXTRACT
C3555472|T121|1420970|RXNORM|INGA EDULIS SEED EXTRACT|INGA EDULIS SEED EXTRACT
C0069833|T121|32698|RXNORM|OXYPHENCYCLIMINE|OXYPHENCYCLIMINE
C3555470|T121|1420972|RXNORM|LIQUIDAMBAR ORIENTALIS RESIN|LIQUIDAMBAR ORIENTALIS RESIN
C3555469|T121|1420973|RXNORM|MOMORDICA COCHINCHINENSIS SEED EXTRACT|MOMORDICA COCHINCHINENSIS SEED EXTRACT
C3555468|T121|1420974|RXNORM|MORUS AUSTRALIS LEAF EXTRACT|MORUS AUSTRALIS LEAF EXTRACT
C3555467|T121|1420975|RXNORM|NELUMBO NUCIFERA STAMEN EXTRACT|NELUMBO NUCIFERA STAMEN EXTRACT
C3555466|T121|1420976|RXNORM|PAEONIA VEITCHII ROOT EXTRACT|PAEONIA VEITCHII ROOT EXTRACT
C3538842|T121|1420977|RXNORM|POLYGONUM CUSPIDATUM WHOLE EXTRACT|POLYGONUM CUSPIDATUM WHOLE EXTRACT
C2699277|T121|1307639|RXNORM|SCHIZONEPETA TENUIFOLIA FLOWERING TOP EXTRACT|NEPETA TENUIFOLIA FLOWERING TOP EXTRACT
C3264705|T121|1307638|RXNORM|LEPIDIUM MEYENII ROOT EXTRACT|LEPIDIUM MEYENII ROOT EXTRACT
C0795661|T121|253199|RXNORM|ROTAVIRUS VACCINE, LIVE|ROTAVIRUS VACCINE, LIVE
C3668772|T121|1441399|RXNORM|RUSSULA EMETICA PREPARATION|RUSSULA EMETICA PREPARATION
C3505519|T121|1358700|RXNORM|BENZOTRIAZOLYL BUTYLPHENOL SULFONATE|BENZOTRIAZOLYL BUTYLPHENOL SULFONATE
C1874194|T121|690788|RXNORM|AMINOPHYLLINE / EPHEDRINE / GUAIFENESIN / PHENOBARBITAL|AMINOPHYLLINE / EPHEDRINE / GUAIFENESIN / PHENOBARBITAL
C3256099|T121|1307631|RXNORM|BAMBUSA ARUNDINACEA LEAF EXTRACT|BAMBUSA ARUNDINACEA LEAF EXTRACT
C0795652|T121|253193|RXNORM|PASSIFLORA INCARNATA EXTRACT|PASSIFLORA INCARNATA EXTRACT
C0795649|T121|253190|RXNORM|OAT BRAN|OAT BRAN
C0795658|T121|253196|RXNORM|RESPIRATORY VACCINE|RESPIRATORY VACCINE
C3255841|T121|1307637|RXNORM|ECHINACEA PURPUREA FLOWERING TOP EXTRACT|ECHINACEA PURPUREA FLOWERING TOP EXTRACT
C3474162|T121|1307636|RXNORM|HAMAMELIS VIRGINIANA FLOWER WATER EXTRACT|HAMAMELIS VIRGINIANA FLOWER WATER EXTRACT
C3255226|T121|1236445|RXNORM|CHLOPHEDIANOL / CHLORCYCLIZINE / PSEUDOEPHEDRINE|CHLOPHEDIANOL / CHLORCYCLIZINE / PSEUDOEPHEDRINE
C0650235|T121|183875|RXNORM|FOMINOBEN|FOMINOBEN
C0650237|T121|183877|RXNORM|CLOFEZONE|CLOFEZONE
C0440015|T121|124150|RXNORM|DANDELION EXTRACT|DANDELION EXTRACT
C2740952|T129|900025|RXNORM|ATLANTIC COD ALLERGENIC EXTRACT|ATLANTIC COD ALLERGENIC EXTRACT
C0314974|T007|285148|RXNORM|BIFIDOBACTERIUM BIFIDUM|BIFIDOBACTERIUM BIFIDUM
C0939797|T121|285149|RXNORM|BANANA EXTRACT|BANANA EXTRACT
C3692931|T121|1442882|RXNORM|CERVUS NIPPON VELVET PREPARATION|CERVUS NIPPON VELVET PREPARATION
C0077524|T121|1114883|RXNORM|TURMERIC EXTRACT|TURMERIC EXTRACT
C0873055|T121|259393|RXNORM|SIBERIAN GINSENG ROOT|SIBERIAN GINSENG ROOT
C1524076|T122|259399|RXNORM|AMILOMER|AMILOMER
C3256554|T121|1314202|RXNORM|POLYETHYLENE GLYCOL 1000000|POLYETHYLENE GLYCOL 1000000
C0254215|T121|75960|RXNORM|REVIPARIN|REVIPARIN
C2987716|T121|1242987|RXNORM|VISMODEGIB|VISMODEGIB
C3555497|T121|1376154|RXNORM|TETRAHYDRODEMETHOXYDIFERULOYLMETHANE|TETRAHYDRODEMETHOXYDIFERULOYLMETHANE
C0028978|T121|7646|RXNORM|OMEPRAZOLE|OMEPRAZOLE
C1719971|T121|644580|RXNORM|LITHIUM SUCCINATE / ZINC SULFATE|LITHIUM SUCCINATE / ZINC SULFATE
C2193899|T121|817255|RXNORM|CAFFEINE / NITROGLYCERIN|CAFFEINE / NITROGLYCERIN
C3488927|T121|1309466|RXNORM|FAGUS SYLVATICA FLOWERING TOP|FAGUS SYLVATICA FLOWERING TOP
C3245306|T121|1190930|RXNORM|ACETAMINOPHEN / DEXBROMPHENIRAMINE|ACETAMINOPHEN / DEXBROMPHENIRAMINE
C3256560|T109|1314203|RXNORM|POLYETHYLENE GLYCOL 600000|POLYETHYLENE GLYCOL 600000
C2928890|T121|1007977|RXNORM|RESORCINOL / SALICYLIC ACID / SODIUM THIOSULFATE|RESORCINOL / SALICYLIC ACID / SODIUM THIOSULFATE
C2727876|T129|975996|RXNORM|PHOMA GLOMERATA ALLERGENIC EXTRACT|PHOMA GLOMERATA ALLERGENIC EXTRACT
C2918532|T129|995754|RXNORM|AMERICAN BASSWOOD POLLEN EXTRACT|TILIA AMERICANA POLLEN EXTRACT
C0054340|T121|19959|RXNORM|ACRIVASTINE|ACRIVASTINE
C0085057|T197|42279|RXNORM|ZINC HYDROXIDE|ZINC HYDROXIDE
C0618388|T121|166718|RXNORM|TILBROQUINOL|TILBROQUINOL
C3555526|T121|1374398|RXNORM|BROSIMUM ACUTIFOLIUM BARK EXTRACT|BROSIMUM ACUTIFOLIUM BARK EXTRACT
C2348390|T121|1374399|RXNORM|EICOSENOIC ACID|GONDOIC ACID
C0011122|T121|1314345|RXNORM|DECOQUINATE|DECOQUINATE
C0028005|T121|7396|RXNORM|NICARDIPINE|NICARDIPINE
C0078569|T121|39786|RXNORM|VENLAFAXINE|VENLAFAXINE
C0771144|T121|235940|RXNORM|CYNARA PREPARATION|CYNARA PREPARATION
C0027996|T127|7393|RXNORM|NIACIN|NIACIN
C0009226|T123|1314344|RXNORM|COENZYME A|COENZYME A
C0028008|T121|7398|RXNORM|NICERGOLINE|NICERGOLINE
C3535822|T130|1370673|RXNORM|SESQUICARBONATE|SESQUICARBONATE
C3535823|T122|1370672|RXNORM|HYDROXYMETHYLGLYCINATE|HYDROXYMETHYLGLYCINATE
C3535824|T122|1370671|RXNORM|STEAROYL LACTYLATE|STEAROYL LACTYLATE
C0057827|T121|1314346|RXNORM|DICETYLPHOSPHATE|DICETYLPHOSPHATE
C0626252|T121|1370677|RXNORM|RETINYL LINOLEATE|RETINYL LINOLEATE
C3535629|T109|1370676|RXNORM|THYMUS CITRIODORUS LEAF EXTRACT|THYMUS CITRIODORUS LEAF EXTRACT
C3535821|T121|1370674|RXNORM|DIHYDROXYBENZOATE|DIHYDROXYBENZOATE
C1725639|T109|1314341|RXNORM|CETETH-10|CETETH-10
C0205951|T197|1370679|RXNORM|SODIUM CHLORIDE, (22)NA|SODIUM CHLORIDE, (22)NA
C3535628|T121|1370678|RXNORM|POLYQUATERNIUM-37 (10000 MPA.S)|POLYQUATERNIUM-37 (10000 MPA.S)
C1875765|T121|690527|RXNORM|SODIUM BICARBONATE / TARTARIC ACID|SODIUM BICARBONATE / TARTARIC ACID
C0771635|T121|236368|RXNORM|SARSAPARILLA PREPARATION|SARSAPARILLA PREPARATION
C1445783|T121|466549|RXNORM|ASPIRIN / CAFFEINE / ORPHENADRINE|ASPIRIN / CAFFEINE / ORPHENADRINE
C0041980|T123|1427088|RXNORM|URIC ACID|URIC ACID
C1445780|T121|466546|RXNORM|ETHINYL ESTRADIOL / FERROUS FUMARATE / NORETHINDRONE|ETHINYL ESTRADIOL / FERROUS FUMARATE / NORETHINDRONE
C0771627|T121|236361|RXNORM|TILIA EXTRACT|TILIA EXTRACT
C1445775|T121|466541|RXNORM|NEOMYCIN / POLYMYXIN B|NEOMYCIN / POLYMYXIN B
C1445775|T121|466541|RXNORM|NEOMYCIN / POLYMYXIN B|NEOMYCIN / POLYMYXIN B
C1445775|T121|466541|RXNORM|NEOMYCIN / POLYMYXIN B|NEOMYCIN / POLYMYXIN B
C1445774|T121|466540|RXNORM|BACITRACIN / NEOMYCIN / POLYMYXIN B / PRAMOXINE|BACITRACIN / NEOMYCIN / POLYMYXIN B / PRAMOXINE
C2146605|T121|814657|RXNORM|ACETAMINOPHEN / CAFFEINE / CODEINE|ACETAMINOPHEN / CAFFEINE / CODEINE
C3256692|T109|1314207|RXNORM|KOJIC DIPALMITATE|KOJIC DIPALMITATE
C3645269|T122|1427125|RXNORM|DIISOCETYL DODECANEDIOATE|DIISOCETYL DODECANEDIOATE
C0368663|T121|113374|RXNORM|AMINOSALICYLATE|AMINOSALICYLATE
C0368663|T121|113374|RXNORM|AMINOSALICYLATE|AMINOSALICYLATE
C0368662|T121|113373|RXNORM|AMINOCAPROATE|AMINOCAPROATE
C2183865|T121|820778|RXNORM|GLUCOSE / LIDOCAINE|GLUCOSE / LIDOCAINE
C3848600|T121|1545040|RXNORM|CONIUM MACULATUM ROOT EXTRACT|CONIUM MACULATUM ROOT EXTRACT
C3855230|T109|1547578|RXNORM|CURCUMA AMADA WHOLE EXTRACT|CURCUMA AMADA WHOLE EXTRACT
C3484528|T121|1342487|RXNORM|CAULOPHYLLUM THALICTROIDES ROOT EXTRACT|CAULOPHYLLUM THALICTROIDES ROOT EXTRACT
C0377349|T121|1595589|RXNORM|SODIUM GLYCEROPHOSPHATE|SODIUM GLYCEROPHOSPHATE
C3486610|T121|1342489|RXNORM|FUCUS SERRATUS EXTRACT|FUCUS SERRATUS EXTRACT
C3486389|T121|1342488|RXNORM|LYCOSA TARANTULA PREPARATION|LYCOSA TARANTULA PREPARATION
C3864846|T121|1595584|RXNORM|LEPIDIUM MEYENII WHOLE EXTRACT|LEPIDIUM MEYENII WHOLE EXTRACT
C3855229|T109|1547577|RXNORM|LACTARIUS INDIGO WHOLE EXTRACT|LACTARIUS INDIGO WHOLE EXTRACT
C0537551|T125|139953|RXNORM|PRAMLINTIDE|PRAMLINTIDE
C3855223|T109|1547571|RXNORM|PIELLIA TERNATA WHOLE EXTRACT|PIELLIA TERNATA WHOLE EXTRACT
C3864850|T121|1595580|RXNORM|OENANTHE CROCATA ROOT EXTRACT|OENANTHE CROCATA ROOT EXTRACT
C3256500|T109|1309405|RXNORM|ARDISIA JAPONICA STEM EXTRACT|ARDISIA JAPONICA STEM EXTRACT
C2702395|T129|895488|RXNORM|DOMESTIC COW HAIR EXTRACT|DOMESTIC COW HAIR EXTRACT
C2979512|T121|1090967|RXNORM|ASCORBIC ACID / CHOLECALCIFEROL / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E|ASCORBIC ACID / CHOLECALCIFEROL / NIACINAMIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E
C1570906|T121|596554|RXNORM|VILDAGLIPTIN|VILDAGLIPTIN
C3264738|T121|1427085|RXNORM|PEPPER EXTRACT|PEPPER EXTRACT
C0018546|T121|5093|RXNORM|HALOPERIDOL|HALOPERIDOL
C1720463|T121|645061|RXNORM|CAMPHOR / CHLOROXYLENOL|CAMPHOR / CHLOROXYLENOL
C0018549|T121|5095|RXNORM|HALOTHANE|HALOTHANE
C3486283|T121|1427084|RXNORM|7-OXO-PRASTERONE|7-KETO-DEHYDROEPIANDROSTERONE
C2719430|T131|860178|RXNORM|RIMABOTULINUMTOXINB|RIMABOTULINUMTOXINB
C0016368|T121|4496|RXNORM|FLUPHENAZINE|FLUPHENAZINE
C0016367|T121|4495|RXNORM|FLUPENTHIXOL|FLUPENTHIXOL
C0016366|T125|4494|RXNORM|FLUOXYMESTERONE|FLUOXYMESTERONE
C0907850|T123|274964|RXNORM|CICLESONIDE|CICLESONIDE
C0907850|T123|274964|RXNORM|CICLESONIDE|CICLESONIDE
C0016360|T121|4492|RXNORM|FLUOROURACIL|FLUOROURACIL
C0016360|T121|4492|RXNORM|FLUOROURACIL|FLUOROURACIL
C0220839|T123|70602|RXNORM|GLUTAMATE|GLUTAMATE
C0220840|T109|70603|RXNORM|GLYCOLATE|GLYCOLATE
C0220840|T109|70603|RXNORM|GLYCOLATE|GLYCOLATE
C2344072|T129|797635|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP Y CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE|NEISSERIA MENINGITIDIS SEROGROUP Y CAPSULAR POLYSACCHARIDE DIPHTHERIA TOXOID PROTEIN CONJUGATE VACCINE
C0907410|T195|274786|RXNORM|TELITHROMYCIN|TELITHROMYCIN
C1656690|T121|605572|RXNORM|CARBINOXAMINE / HYDROCODONE / PHENYLEPHRINE|CARBINOXAMINE / HYDROCODONE / PHENYLEPHRINE
C0009213|T168|2669|RXNORM|COD LIVER OIL|COD LIVER OIL
C2929615|T121|1008716|RXNORM|BENZOCAINE / CHLOROXYLENOL / ISOPROPYL ALCOHOL / RESORCINOL / SALICYLIC ACID|BENZOCAINE / CHLOROXYLENOL / ISOPROPYL ALCOHOL / RESORCINOL / SALICYLIC ACID
C2929616|T121|1008717|RXNORM|ALANINE / ARGININE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE|ALANINE / ARGININE / CYSTEINE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / PHENYLALANINE / PHOSPHORIC ACID / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE
C2929613|T121|1008714|RXNORM|COCOA BUTTER / SHARK LIVER OIL|COCOA BUTTER / SHARK LIVER OIL
C2929614|T121|1008715|RXNORM|COCOA BUTTER / PHENYLEPHRINE / SHARK LIVER OIL|COCOA BUTTER / PHENYLEPHRINE / SHARK LIVER OIL
C2929612|T121|1008713|RXNORM|ALANINE / ARGININE / ASPARTATE / GLUCOSE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / N-ACETYLTYROSINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE|ALANINE / ARGININE / ASPARTATE / GLUCOSE / GLUTAMATE / GLYCINE / HISTIDINE / ISOLEUCINE / LEUCINE / LYSINE / METHIONINE / N-ACETYLTYROSINE / PHENYLALANINE / PROLINE / SERINE / THREONINE / TRYPTOPHAN / VALINE
C2929609|T121|1008710|RXNORM|LACTASE / LACTOBACILLUS ACIDOPHILUS|LACTASE / LACTOBACILLUS ACIDOPHILUS
C2929610|T121|1008711|RXNORM|BENZOCAINE / OXYQUINOLINE|BENZOCAINE / OXYQUINOLINE
C3651709|T121|1431284|RXNORM|GLECHOMA HEDERACEA FLOWERING TOP EXTRACT|GLECHOMA HEDERACEA FLOWERING TOP EXTRACT
C3651708|T109|1431285|RXNORM|TOMATO SEED OIL|TOMATO SEED OIL
C2929617|T121|1008718|RXNORM|DOCOSAHEXAENOATE / EICOSAPENTAENOATE|DOCOSAHEXAENOATE / EICOSAPENTAENOATE
C2929618|T121|1008719|RXNORM|ETHANOL / SALICYLIC ACID|ETHANOL / SALICYLIC ACID
C2929618|T121|1008719|RXNORM|ETHANOL / SALICYLIC ACID|ETHANOL / SALICYLIC ACID
C3486349|T109|1305715|RXNORM|ROSA CANINA FRUIT OIL|ROSA CANINA FRUIT OIL
C2183068|T121|818139|RXNORM|DEXAMETHASONE / TERFENADINE|DEXAMETHASONE / TERFENADINE
C0071145|T121|33783|RXNORM|PIROCTONE OLAMINE|PIROCTONE OLAMINE
C0051242|T121|1318494|RXNORM|ALLYLTHIOUREA|ALLYLTHIOUREA
C2722689|T129|864701|RXNORM|INFLUENZA A-CALIFORNIA-7-2009-(H1N1)V-LIKE VIRUS VACCINE|INFLUENZA A-CALIFORNIA-7-2009-(H1N1)V-LIKE VIRUS VACCINE
C0077144|T121|38668|RXNORM|TRILOSTANE|TRILOSTANE
C3643657|T121|1423306|RXNORM|DEXTROMETHORPHAN / PYRILAMINE|DEXTROMETHORPHAN / PYRILAMINE
C3643341|T121|1424462|RXNORM|THAUMATOCOCCUS DANIELLII FRUIT EXTRACT|THAUMATOCOCCUS DANIELLII FRUIT EXTRACT
C3643651|T121|1424461|RXNORM|COCOYL GLYCINATE|COCOYL GLYCINATE
C3528829|T121|1363468|RXNORM|RHODOMYRTUS TOMENTOSA FRUIT EXTRACT|RHODOMYRTUS TOMENTOSA FRUIT EXTRACT
C3528830|T121|1363469|RXNORM|VACHELLIA FARNESIANA FLOWER EXTRACT|VACHELLIA FARNESIANA FLOWER EXTRACT
C2938378|T121|1012123|RXNORM|CHLORCYCLIZINE / CODEINE / PSEUDOEPHEDRINE|CHLORCYCLIZINE / CODEINE / PSEUDOEPHEDRINE
C3812628|T121|1490685|RXNORM|MENTHA ARVENSIS WHOLE EXTRACT|MENTHA ARVENSIS WHOLE EXTRACT
C0076115|T121|37806|RXNORM|TERCONAZOLE|TERCONAZOLE
C3818798|T121|1490687|RXNORM|PAEONIA LACTIFLORA WHOLE EXTRACT|PAEONIA LACTIFLORA WHOLE EXTRACT
C3818799|T121|1490686|RXNORM|NOTOPTERYGIUM INCISUM WHOLE EXTRACT|NOTOPTERYGIUM INCISUM WHOLE EXTRACT
C3464429|T121|1292029|RXNORM|CHOLECALCIFEROL / DOCOSAHEXAENOATE / EICOSAPENTAENOATE|CHOLECALCIFEROL / DOCOSAHEXAENOATE / EICOSAPENTAENOATE
C0720955|T121||RXNORM|HYDROCORTISONE / IODOQUINOL
C0076110|T121|37801|RXNORM|TERBINAFINE|TERBINAFINE
C0076110|T121|37801|RXNORM|TERBINAFINE|TERBINAFINE
C3818802|T121|1490682|RXNORM|BLETILLA STRIATA WHOLE EXTRACT|BLETILLA STRIATA WHOLE EXTRACT
C0068742|T121|31782|RXNORM|NIFUROXAZIDE|NIFUROXAZIDE
C0720956|T121|217627|RXNORM|HYDROCORTISONE / NEOMYCIN / POLYMYXIN B|HYDROCORTISONE / NEOMYCIN / POLYMYXIN B
C0720956|T121|217627|RXNORM|HYDROCORTISONE / NEOMYCIN / POLYMYXIN B|HYDROCORTISONE / NEOMYCIN / POLYMYXIN B
C0720956|T121|217627|RXNORM|HYDROCORTISONE / NEOMYCIN / POLYMYXIN B|HYDROCORTISONE / NEOMYCIN / POLYMYXIN B
C2962068|T129|1427044|RXNORM|PENICILLIUM DIGITATUM ALLERGENIC EXTRACT|PENICILLIUM DIGITATUM ALLERGENIC EXTRACT
C3818797|T121|1490688|RXNORM|REHMANNIA GLUTINOSA WHOLE EXTRACT|REHMANNIA GLUTINOSA WHOLE EXTRACT
C0051736|T121|17804|RXNORM|AMOROLFINE|AMOROLFINE
C2947886|T121|1042981|RXNORM|CATALASE / CYSTEINE / LYSINE / METHIONINE / SUPEROXIDE DISMUTASE|CATALASE / CYSTEINE / LYSINE / METHIONINE / SUPEROXIDE DISMUTASE
C3486648|T121|1353883|RXNORM|PRUNUS CERASIFERA FLOWER EXTRACT|PRUNUS CERASIFERA FLOWER EXTRACT
C0063479|T121|27518|RXNORM|INDOBUFEN|INDOBUFEN
C0772488|T121|237148|RXNORM|BISMUTH-FORMIC-IODIDE|BISMUTH-FORMIC-IODIDE
C0008292|T121|2407|RXNORM|CHLORQUINALDOL|CHLORQUINALDOL
C3484465|T121|1353881|RXNORM|HEDEOMA PULEGIOIDES EXTRACT|HEDEOMA PULEGIOIDES EXTRACT
C0066282|T121|29787|RXNORM|METHYL SALICYLATE|METHYL SALICYLATE
C0002680|T195|733|RXNORM|AMPICILLIN|AMPICILLIN
C0002679|T195|732|RXNORM|AMPHOTERICIN B|AMPHOTERICIN B
C0002679|T195|732|RXNORM|AMPHOTERICIN B|AMPHOTERICIN B
C3692720|T121|1442505|RXNORM|CUPRESSUS SEMPERVIRENS LEAFY TWIG EXTRACT|CUPRESSUS SEMPERVIRENS LEAFY TWIG EXTRACT
C3692719|T121|1442504|RXNORM|AZADIRACHTA INDICA SEED EXTRACT|AZADIRACHTA INDICA SEED EXTRACT
C3692722|T121|1442507|RXNORM|CYMBOPOGON MARTINI TOP EXTRACT|CYMBOPOGON MARTINI TOP EXTRACT
C3692721|T121|1442506|RXNORM|CYMBOPOGON FLEXUOSUS WHOLE EXTRACT|CYMBOPOGON FLEXUOSUS WHOLE EXTRACT
C3692724|T121|1442509|RXNORM|LITSEA CUBEBA FRUIT EXTRACT|LITSEA CUBEBA FRUIT EXTRACT
C0002697|T121|738|RXNORM|INAMRINONE|INAMRINONE
C3486729|T121|1353886|RXNORM|PETROSELINUM CRISPUM EXTRACT|PETROSELINUM CRISPUM EXTRACT
C3848602|T121|1545037|RXNORM|ABIES ALBA LEAFY TWIG EXTRACT|ABIES ALBA LEAFY TWIG EXTRACT
C3486701|T121|1353885|RXNORM|EUPHRASIA STRICTA EXTRACT|EUPHRASIA STRICTA EXTRACT
C3255591|T121|1311694|RXNORM|GLYCERYL COCOATE|GLYCERYL COCOATE
C1576815|T122|1311695|RXNORM|GLYCERYL ISOSTEARATE|GLYCERYL ISOSTEARATE
C3848601|T121|1545039|RXNORM|BOS TAURUS COLON PREPARATION|BOS TAURUS COLON PREPARATION
C1531654|T121|484139|RXNORM|CHLORHEXIDINE / ISOPROPYL ALCOHOL|CHLORHEXIDINE / ISOPROPYL ALCOHOL
C1962788|T121|1311690|RXNORM|GLYCERYL DISTEARATE|GLYCERYL DISTEARATE
C3256841|T121|1311691|RXNORM|GLYCERYL DILAURATE|GLYCERYL DILAURATE
C3267302|T121|1311692|RXNORM|GLYCERYL MYRISTATE|GLYCERYL MYRISTATE
C1509379|T121|1311693|RXNORM|GLYCERYL LAURATE|GLYCERYL LAURATE
C2928523|T121|1007605|RXNORM|PHENYLEPHRINE / POLYVINYL ALCOHOL|PHENYLEPHRINE / POLYVINYL ALCOHOL
C2928522|T121|1007604|RXNORM|BACITRACIN / DIPERODON / NEOMYCIN|BACITRACIN / DIPERODON / NEOMYCIN
C2928525|T121|1007607|RXNORM|MAGNESIUM HYDROXIDE / MALIC ACID|MAGNESIUM HYDROXIDE / MALIC ACID
C2928524|T121|1007606|RXNORM|CHROMOUS CHLORIDE / COPPER SULFATE / MANGANESE CHLORIDE / MOLYBDENUM / SELENIOUS ACID / SODIUM IODIDE / ZINC SULFATE|CHROMOUS CHLORIDE / COPPER SULFATE / MANGANESE CHLORIDE / MOLYBDENUM / SELENIOUS ACID / SODIUM IODIDE / ZINC SULFATE
C2928519|T121|1007601|RXNORM|BRILLIANT GREEN / LACTATE|BRILLIANT GREEN / LACTATE
C2928274|T121|1007352|RXNORM|BROMELAINS / PAPAIN|BROMELAINS / PAPAIN
C2928273|T121|1007351|RXNORM|GLYCOLATE / HYDROQUINONE|GLYCOLATE / HYDROQUINONE
C2928520|T121|1007602|RXNORM|COAL TAR / PINE TAR|COAL TAR / PINE TAR
C2928527|T121|1007609|RXNORM|MERCURY, AMMONIATED / SALICYLIC ACID|MERCURY, AMMONIATED / SALICYLIC ACID
C2928526|T121|1007608|RXNORM|BELLADONNA ALKALOIDS / PHENOBARBITAL|BELLADONNA ALKALOIDS / PHENOBARBITAL
C2928280|T121|1007358|RXNORM|GLYCERIN / HYPROMELLOSE / NAPHAZOLINE|GLYCERIN / HYPROMELLOSE / NAPHAZOLINE
C3555518|T122|1374804|RXNORM|C12-15 PARETH-12|C12-15 PARETH-12
C1874708|T121|691205|RXNORM|CARAMIPHEN / CHLORPHENIRAMINE / ISOPROPAMIDE / PHENYLPROPANOLAMINE|CARAMIPHEN / CHLORPHENIRAMINE / ISOPROPAMIDE / PHENYLPROPANOLAMINE
C3152587|T121|1095603|RXNORM|ASCORBIC ACID / BIOTIN / CHOLECALCIFEROL / FOLIC ACID / NIACIN / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12|ASCORBIC ACID / BIOTIN / CHOLECALCIFEROL / FOLIC ACID / NIACIN / PANTOTHENIC ACID / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C0886631|T121|1374802|RXNORM|POTASSIUM CITRATE ANHYDROUS|POTASSIUM CITRATE ANHYDROUS
C2928267|T121|1007345|RXNORM|DOXYLAMINE / VITAMIN B6|DOXYLAMINE / VITAMIN B6
C2928268|T121|1007346|RXNORM|ALLANTOIN / HEXACHLOROPHENE / SQUALENE|ALLANTOIN / HEXACHLOROPHENE / SQUALENE
C2928529|T121|1007611|RXNORM|BACITRACIN / LIDOCAINE / NEOMYCIN / POLYMYXIN B|BACITRACIN / LIDOCAINE / NEOMYCIN / POLYMYXIN B
C1176020|T121|357977|RXNORM|SUNITINIB|SUNITINIB
C3555506|T109|1376097|RXNORM|TRIMETHYLBENZENEPROPANOL|TRIMETHYLBENZENEPROPANOL
C3555507|T109|1376096|RXNORM|ETHYL LINALOOL|ETHYL LINALOOL
C3555504|T109|1376099|RXNORM|GLYCERYL TRIBEHENATE- ISOSTEARATE- EICOSANDIOATE|GLYCERYL TRIBEHENATE- ISOSTEARATE- EICOSANDIOATE
C2928262|T121|1007340|RXNORM|CHLORTHALIDONE / METOPROLOL|CHLORTHALIDONE / METOPROLOL
C2928263|T121|1007341|RXNORM|VITAMIN B6 / ZINC PICOLINATE|VITAMIN B6 / ZINC PICOLINATE
C2720503|T129|862460|RXNORM|CASEIN ALLERGENIC EXTRACT|CASEIN ALLERGENIC EXTRACT
C2722031|T129|862461|RXNORM|CHERRY ALLERGENIC EXTRACT|CHERRY ALLERGENIC EXTRACT
C2928264|T121|1007342|RXNORM|LINOLEATE / RICINOLEATE|LINOLEATE / RICINOLEATE
C2928265|T121|1007343|RXNORM|FLUOROMETHOLONE / NEOMYCIN|FLUOROMETHOLONE / NEOMYCIN
C0106556|T121|47181|RXNORM|BISMUTH SUBCITRATE|BISMUTH SUBCITRATE
C0106555|T121|47180|RXNORM|BISMUTH TRIBROMOPHENATE|BISMUTH TRIBROMOPHENATE
C0937769|T121|283677|RXNORM|CORN SILK PREPARATION|CORN SILK PREPARATION
C0032613|T121|8565|RXNORM|POLYTHIAZIDE|POLYTHIAZIDE
C0937767|T121|283675|RXNORM|CINA ARTEMISIA PREPARATION|CINA ARTEMISIA PREPARATION
C0032602|T122|8561|RXNORM|POLYSORBATES|POLYSORBATES
C0032601|T122|8560|RXNORM|POLYSORBATE 80|POLYSORBATE 80
C1966712|T121|747890|RXNORM|CITRIC ACID / POTASSIUM BICARBONATE|CITRIC ACID / POTASSIUM BICARBONATE
C0072826|T122|283678|RXNORM|QUATERNIUM-15|QUATERNIUM-15
C0937771|T121|283679|RXNORM|EUPHRASIA OFFICINALIS PREPARATION|EUPHRASIA OFFICINALIS PREPARATION
C2718386|T129|857921|RXNORM|INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN|INFLUENZA VIRUS VACCINE, INACTIVATED B-BRISBANE-60-2008 STRAIN
C3465069|T121|1293735|RXNORM|CHROMIC CHLORIDE / COPPER SULFATE / MANGANESE SULFATE / SELENIOUS ACID / ZINC SULFATE|CHROMIC CHLORIDE / COPPER SULFATE / MANGANESE SULFATE / SELENIOUS ACID / ZINC SULFATE
C2934193|T121|1546059|RXNORM|OLODATEROL|OLODATEROL
C3255770|T109|1369682|RXNORM|ETHYLHEXYL STEARATE|ETHYLHEXYL STEARATE
C3535662|T121|1369683|RXNORM|ISOCETETH-10|ISOCETETH-10
C2827093|T121|1085787|RXNORM|BUTYLSCOPOLAMINE|BUTYLSCOPOLAMINE
C3535660|T121|1369686|RXNORM|LONICERA JAPONICA TOP EXTRACT|LONICERA JAPONICA TOP EXTRACT
C1876200|T125|1044584|RXNORM|TESAMORELIN|TESAMORELIN
C3500171|T121|1313924|RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / BETA CAROTENE / CALCIUM CARBONATE / CHOLECALCIFEROL / DOCUSATE / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC OXIDE|ALPHA TOCOPHEROL / ASCORBIC ACID / BETA CAROTENE / CALCIUM CARBONATE / CHOLECALCIFEROL / DOCUSATE / FERROUS FUMARATE / FOLIC ACID / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12 / ZINC OXIDE
C3535657|T121|1369689|RXNORM|SIMMONDSIA CHINENSIS WHOLE EXTRACT|SIMMONDSIA CHINENSIS WHOLE EXTRACT
C0028193|T197|7476|RXNORM|NITROPRUSSIDE|NITROPRUSSIDE
C3255108|T127|1236136|RXNORM|TOCOPHEROL|TOCOPHEROL
C2684342|T129|851898|RXNORM|SWEET VERNAL GRASS POLLEN EXTRACT|ANTHOXANTHUM ODORATUM POLLEN EXTRACT
C0054086|T121|19729|RXNORM|IDROCILAMIDE|IDROCILAMIDE
C0723505|T121||RXNORM|SULFABENZAMIDE / SULFACETAMIDE / SULFATHIAZOLE
C0042523|T121|11170|RXNORM|VERAPAMIL|VERAPAMIL
C0042523|T121|11170|RXNORM|VERAPAMIL|VERAPAMIL
C3499523|T121|1312391|RXNORM|GLYCERETH-17 COCOATE|GLYCERETH-17 COCOATE
C2183746|T121|816286|RXNORM|DIPHENYLPYRALINE / PHENYLPROPANOLAMINE|DIPHENYLPYRALINE / PHENYLPROPANOLAMINE
C0057605|T121|22696|RXNORM|DEXBROMPHENIRAMINE|DEXBROMPHENIRAMINE
C0057606|T121|22697|RXNORM|DEXCHLORPHENIRAMINE|DEXCHLORPHENIRAMINE
C3555462|T121|1421146|RXNORM|PIKEA ROBUSTA EXTRACT|PIKEA ROBUSTA EXTRACT
C3555461|T121|1421147|RXNORM|BOS TAURUS BONE PREPARATION|BOVINE BONE PREPARATION
C0024742|T121|6633|RXNORM|MANNOSE|MANNOSE
C3255761|T121|1313697|RXNORM|ETHYLCELLULOSE (20 MPA.S)|ETHYLCELLULOSE (20 MPA.S)
C0718050|T121|214824|RXNORM|SEVELAMER|SEVELAMER
C1874389|T121|689599|RXNORM|ATROPINE / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE|ATROPINE / CHLORPHENIRAMINE / PHENYLPROPANOLAMINE
C1874388|T121|689598|RXNORM|ATROPINE / CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLTOLOXAMINE|ATROPINE / CHLORPHENIRAMINE / PHENYLEPHRINE / PHENYLTOLOXAMINE
C3485009|T121|1313690|RXNORM|EUPATORIUM JAPONICUM WHOLE EXTRACT|EUPATORIUM JAPONICUM WHOLE EXTRACT
C3486529|T121|1313691|RXNORM|NASTURTIUM OFFICIENALE WHOLE EXTRACT|NASTURTIUM OFFICIENALE WHOLE EXTRACT
C1533126|T121|588250|RXNORM|MILNACIPRAN|MILNACIPRAN
C1874387|T121|689597|RXNORM|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PHENYLEPHRINE / SCOPOLAMINE|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PHENYLEPHRINE / SCOPOLAMINE
C1874386|T121|689596|RXNORM|ATROPINE / CHLORPHENIRAMINE / EPHEDRINE|ATROPINE / CHLORPHENIRAMINE / EPHEDRINE
C1874383|T121|689593|RXNORM|ATROPINE / BROMPHENIRAMINE / PHENYLTOLOXAMINE / PSEUDOEPHEDRINE|ATROPINE / BROMPHENIRAMINE / PHENYLTOLOXAMINE / PSEUDOEPHEDRINE
C3255822|T109|1313699|RXNORM|METHYLCELLULOSE (15 CPS)|METHYLCELLULOSE (15 CPS)
C3848626|T121|1544128|RXNORM|SUS SCROFA MENISCUS PREPARATION|SUS SCROFA MENISCUS PREPARATION
C3834045|T109|1543773|RXNORM|PEG-8 CAPRYLIC-CAPRIC GLYCERIDES|PEG-8 CAPRYLIC-CAPRIC GLYCERIDES
C0055617|T197|21009|RXNORM|CHROMIC CHLORIDE|CHROMIC CHLORIDE
C2193906|T121|818351|RXNORM|AMILORIDE / FUROSEMIDE|AMILORIDE / FUROSEMIDE
C3666698|T121|1437505|RXNORM|STYPHNOLOBIUM JAPONICUM LEAF EXTRACT|STYPHNOLOBIUM JAPONICUM LEAF EXTRACT
C2347739|T168|1437504|RXNORM|QUINOA OIL|QUINOA OIL
C2000261|T121|1307404|RXNORM|LINACLOTIDE|LINACLOTIDE
C0054654|T121|20206|RXNORM|CARBARSON|CARBARSON
C3666697|T121|1437503|RXNORM|OENOTHERA BIENNIS SEED EXTRACT|OENOTHERA BIENNIS SEED EXTRACT
C0459821|T121|126291|RXNORM|PUMPKIN SEED EXTRACT|PUMPKIN SEED EXTRACT
C2741588|T129|901509|RXNORM|NEISSERIA MENINGITIDIS SEROGROUP W-135 OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE|NEISSERIA MENINGITIDIS SEROGROUP W-135 OLIGOSACCHARIDE DIPHTHERIA CRM197 PROTEIN CONJUGATE VACCINE
C0717453|T121|214261|RXNORM|ATROPINE / DIFENOXIN|ATROPINE / DIFENOXIN
C0717456|T121|214263|RXNORM|ATROPINE / PHENOBARBITAL|ATROPINE / PHENOBARBITAL
C0717455|T121|214262|RXNORM|ATROPINE / EDROPHONIUM|ATROPINE / EDROPHONIUM
C0717459|T121|214265|RXNORM|AZATADINE / PSEUDOEPHEDRINE|AZATADINE / PSEUDOEPHEDRINE
C0717444|T121|669119|RXNORM|ASPIRIN / DIPHENHYDRAMINE|ASPIRIN / DIPHENHYDRAMINE
C3486065|T109|1312646|RXNORM|PEG-150 PENTAERYTHRITYL TETRASTEARATE|PEG-150 PENTAERYTHRITYL TETRASTEARATE
C0377223|T121|114464|RXNORM|ARGININE GLUTAMATE|ARGININE GLUTAMATE
C3667883|T109|1440250|RXNORM|HYDROGENATED DIDECENE|HYDROGENATED DIDECENE
C2928219|T121|1007297|RXNORM|GUAIACOLSULFONATE / GUAIFENESIN|GUAIACOLSULFONATE / GUAIFENESIN
C3832606|T109|1539193|RXNORM|STYPHNOLOBIUM JAPONICUM FLOWER EXTRACT|STYPHNOLOBIUM JAPONICUM FLOWER EXTRACT
C0719064|T121|215799|RXNORM|CHOLINE MAGNESIUM TRISALICYCLATE|CHOLINE MAGNESIUM TRISALICYCLATE
C1443114|T129|465168|RXNORM|ANTHOXANTHUM ODORATUM ANTIGEN|ANTHOXANTHUM ODORATUM ANTIGEN
C2368977|T121|824547|RXNORM|ACAI EXTRACT|ACAI EXTRACT
C2073872|T121|814767|RXNORM|CHLORPHENIRAMINE / PHENYLEPHRINE / SALICYLAMIDE|CHLORPHENIRAMINE / PHENYLEPHRINE / SALICYLAMIDE
C0304933|T121|91495|RXNORM|SOY PROTEIN-IRON COMPLEX|SOY PROTEIN-IRON COMPLEX
C3832605|T109|1539192|RXNORM|TILIA PLATYPHYLLOS FLOWER EXTRACT|TILIA PLATYPHYLLOS FLOWER EXTRACT
C2928213|T121|1007291|RXNORM|POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, DIBASIC|POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, DIBASIC
C0056686|T121|21914|RXNORM|CICLETANINE|CICLETANINE
C1698215|T121|640062|RXNORM|REGADENOSON|REGADENOSON
C2364537|T129|805537|RXNORM|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-SOUTH DAKOTA-6-2007 (H1N1) (A-BRISBANE-59-2007-LIKE) STRAIN|INFLUENZA VIRUS VACCINE, LIVE ATTENUATED, A-SOUTH DAKOTA-6-2007 (H1N1) (A-BRISBANE-59-2007-LIKE) STRAIN
C3537577|T121|1371037|RXNORM|LIPPIA CITRIODORA LEAF EXTRACT|LIPPIA CITRIODORA LEAF EXTRACT
C3537575|T121|1371034|RXNORM|CRAMBE MARITIMA LEAF EXTRACT|CRAMBE MARITIMA LEAF EXTRACT
C3555510|T109|1376087|RXNORM|CESTRUM LATIFOLIUM LEAF EXTRACT|CESTRUM LATIFOLIUM LEAF EXTRACT
C3537578|T123|1371038|RXNORM|CROTON LECHLERI RESIN|CROTON LECHLERI RESIN
C0051252|T121|17392|RXNORM|ALOGLUTAMOL|ALOGLUTAMOL
C0016986|T121|4648|RXNORM|GALLOPAMIL|GALLOPAMIL
C2222729|T121|814770|RXNORM|BENZOCAINE / TETRACAINE|BENZOCAINE / TETRACAINE
C3832604|T109|1539191|RXNORM|UNCARIA GAMBIR WHOLE EXTRACT|UNCARIA GAMBIR WHOLE EXTRACT
C2080439|T121|814467|RXNORM|PHENAZOPYRIDINE / TERIZIDONE|PHENAZOPYRIDINE / TERIZIDONE
C0085250|T197|1488368|RXNORM|TECHNETIUM TC-99M PYROPHOSPHATE|TECHNETIUM TC-99M PYROPHOSPHATE
C0303381|T197|90521|RXNORM|CALCIUM SULFIDE|CALCIUM SULFIDE
C0008574|T196|2496|RXNORM|CHROMIUM|CHROMIUM
C0054270|T121|19895|RXNORM|BUTRIPTYLINE|BUTRIPTYLINE
C2000128|T197|1483618|RXNORM|SODIUM HYDRIDE|SODIUM HYDRIDE
C1165664|T129|852363|RXNORM|EASTERN COTTONWOOD POLLEN EXTRACT|POPULUS DELTOIDES POLLEN EXTRACT
C0004599|T195|1291|RXNORM|OMEGA-3 ACID ETHYL ESTERS (USP) / PHYTOSTEROLS|BACITRACIN
C0030349|T121|7894|RXNORM|PAPAVERETUM|PAPAVERETUM
C0030350|T121|7895|RXNORM|PAPAVERINE|PAPAVERINE
C0030346|T126|7892|RXNORM|PAPAIN|PAPAIN
C0030342|T127|7891|RXNORM|PANTOTHENIC ACID|PANTOTHENIC ACID
C0243417|T197|1367162|RXNORM|HECTORITE|HECTORITE
C0073102|T121|1367161|RXNORM|RETINAMIDE|RETINAMIDE
C0072227|T109|1367160|RXNORM|PROPYLENE GLYCOL METHYL ETHER|PROPYLENE GLYCOL METHYL ETHER
C2725366|T122|1367167|RXNORM|ISONONYL ISONONANOATE|ISONONYL ISONONANOATE
C0046343|T121|1367166|RXNORM|2-METHYL-4-ISOTHIAZOLIN-3-ONE|METHYLISOTHIAZOLINONE
C0982254|T121|1367165|RXNORM|LAURETH-23|LAURETH-23
C0772204|T121|1367164|RXNORM|PURSLANE OIL|PURSLANE OIL
C3245388|T121|1191209|RXNORM|DOG HAIR EXTRACT / SHORT RAGWEED POLLEN EXTRACT|DOG HAIR EXTRACT / SHORT RAGWEED POLLEN EXTRACT
C3486553|T129|1367192|RXNORM|HAEMOPHILUS INFLUENZAE IMMUNOSERUM RABBIT|HAEMOPHILUS INFLUENZAE IMMUNOSERUM RABBIT
C0357059|T121|105655|RXNORM|FERROUS GLYCINE SULFATE|FERROUS GLYCINE SULFATE
C3255825|T121|1367168|RXNORM|METHYLPROPANEDIOL|METHYLPROPANEDIOL
C0000665|T130|110|RXNORM|OXYQUINOLINE|OXYQUINOLINE
C2827263|T122|1309718|RXNORM|METHACRYLIC ACID - ETHYL ACRYLATE COPOLYMER (1:1) TYPE A|METHACRYLIC ACID - ETHYL ACRYLATE COPOLYMER (1:1) TYPE A
C3488291|T121|1309719|RXNORM|JUNIPERUS SABINA LEAFY TWIG EXTRACT|JUNIPERUS SABINA LEAFY TWIG EXTRACT
C3489245|T121|1309710|RXNORM|NEOPICRORHIZA SCROPHULARIIFLORA ROOT EXTRACT|NEOPICRORHIZA SCROPHULARIIFLORA ROOT EXTRACT
C3486866|T121|1309711|RXNORM|PHYTOLACCA AMERICANA ROOT EXTRACT|PHYTOLACCA AMERICANA ROOT EXTRACT
C3489246|T121|1309713|RXNORM|PTELEA TRIFOLIATA BARK EXTRACT|PTELEA TRIFOLIATA BARK EXTRACT
C0074414|T121|36453|RXNORM|SEVOFLURANE|SEVOFLURANE
C3485059|T121|1309716|RXNORM|VERBASCUM PHLOMOIDES FLOWER EXTRACT|VERBASCUM PHLOMOIDES FLOWER EXTRACT
C3486867|T121|1309717|RXNORM|RHODODENDRON AUREUM LEAF EXTRACT|RHODODENDRON CHRYSANTHUM LEAF EXTRACT
C0054053|T130|19698|RXNORM|BRILLIANT GREEN|BRILLIANT GREEN
C0314881|T007|1316426|RXNORM|BACILLUS FIRMUS|BACILLUS FIRMUS
C0314840|T007|1316425|RXNORM|ALCALIGENES FAECALIS|ALCALIGENES FAECALIS
C2005695|T121|820541|RXNORM|ACETAMINOPHEN / BUTABARBITAL|ACETAMINOPHEN / BUTABARBITAL
C2722038|T129|862475|RXNORM|GOAT MILK ALLERGENIC EXTRACT|GOAT MILK ALLERGENIC EXTRACT
C0772179|T121|236857|RXNORM|VALEPOTRIATE|VALEPOTRIATE
C0050953|T121|1441428|RXNORM|AGARIC ACID|AGARIC ACID
C3536783|T121|1424898|RXNORM|LOCUST BEAN GUM EXTRACT|LOCUST BEAN GUM EXTRACT
C0873014|T121|1424897|RXNORM|JUJUBE FRUIT EXTRACT|JUJUBE FRUIT EXTRACT
C1712062|T121|637205|RXNORM|PHYTOSTEROL ESTERS|PHYTOSTEROL ESTERS
C3832608|T109|1539195|RXNORM|BABASSU SEED EXTRACT|BABASSU SEED EXTRACT
C2698896|T121|1356149|RXNORM|PROPYLENE GLYCOL MONOLAURATE|PROPYLENE GLYCOL MONOLAURATE
C1136868|T109|1356148|RXNORM|OCTYLDODECYL STEAROYL STEARATE|OCTYLDODECYL STEAROYL STEARATE
C1302895|T121|392617|RXNORM|IBUPROFEN / MENTHOL|IBUPROFEN / MENTHOL
C0982266|T121|314718|RXNORM|MAGNESIUM ACETATE|MAGNESIUM ACETATE
C3500840|T121|1356141|RXNORM|UNDECETH-7|UNDECETH-7
C3500839|T168|1356140|RXNORM|PHYLLANTHUS EMBLICA FRUIT JUICE EXTRACT|PHYLLANTHUS EMBLICA FRUIT JUICE
C3256777|T204|1356143|RXNORM|SACCHARINA LATISSIMA EXTRACT|SACCHARINA LATISSIMA EXTRACT
C0536786|T197|1356142|RXNORM|STRONTIUM NITRATE|STRONTIUM NITRATE
C0982259|T121|314712|RXNORM|LILIUM LONGIFLORIUM|LILIUM LONGIFLORIUM
C0672708|T121|194337|RXNORM|VORINOSTAT|VORINOSTAT
C0605820|T109|1356147|RXNORM|STEARYL GLYCYRRHETINATE|STEARYL GLYCYRRHETINATE
C3500841|T121|1356146|RXNORM|ERYTHORBATE|ERYTHORBATE
C2929929|T121|1009034|RXNORM|ASCORBIC ACID / FERROUS FUMARATE / VITAMIN B 12|ASCORBIC ACID / FERROUS FUMARATE / VITAMIN B 12
C0003438|T121|1009|RXNORM|BILBERRY EXTRACT / BIOFLAVONOIDS / QUERCETIN / RUTIN|ANTITHROMBIN III
C2929931|T121|1009036|RXNORM|AMBROXOL / AMPICILLIN|AMBROXOL / AMPICILLIN
C2929932|T121|1009037|RXNORM|IBUPROFEN / METHOCARBAMOL|IBUPROFEN / METHOCARBAMOL
C2929925|T121|1009030|RXNORM|CAMPHOR / CAPSICUM EXTRACT / MENTHOL|CAMPHOR / CAPSICUM EXTRACT / MENTHOL
C2929926|T121|1009031|RXNORM|ASTEMIZOLE / PSEUDOEPHEDRINE|ASTEMIZOLE / PSEUDOEPHEDRINE
C2927852|T121|1006929|RXNORM|AMYLASES / CELLULASE / ENDOPEPTIDASES / HYOSCYAMINE / LIPASE / PHENYLTOLOXAMINE|AMYLASES / CELLULASE / ENDOPEPTIDASES / HYOSCYAMINE / LIPASE / PHENYLTOLOXAMINE
C2927851|T121|1006928|RXNORM|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PHENYLEPHRINE|ATROPINE / CHLORPHENIRAMINE / HYOSCYAMINE / PHENYLEPHRINE
C2927850|T121|1006927|RXNORM|DIFLUCORTOLONE / SALICYLIC ACID|DIFLUCORTOLONE / SALICYLIC ACID
C2927849|T121|1006926|RXNORM|BISACODYL / CASANTHRANOL|BISACODYL / CASANTHRANOL
C2927848|T121|1006925|RXNORM|MONOFLUOROPHOSPHATE / SODIUM FLUORIDE|MONOFLUOROPHOSPHATE / SODIUM FLUORIDE
C2927847|T121|1006924|RXNORM|CHLORQUINALDOL / DIFLUCORTOLONE|CHLORQUINALDOL / DIFLUCORTOLONE
C2929933|T121|1009038|RXNORM|ASPIRIN / PAPAVERINE / PHENOBARBITAL|ASPIRIN / PAPAVERINE / PHENOBARBITAL
C2929934|T121|1009039|RXNORM|ADENOSINE TRIPHOSPHATE / VITAMIN B6|ADENOSINE TRIPHOSPHATE / VITAMIN B6
C2927845|T121|1006921|RXNORM|CLIOQUINOL / TRIAMCINOLONE|CLIOQUINOL / TRIAMCINOLONE
C2927844|T121|1006920|RXNORM|MICONAZOLE / ZINC OXIDE|MICONAZOLE / ZINC OXIDE
C0025639|T121|6833|RXNORM|METHENOLONE|METHENOLONE
C0025638|T121|6832|RXNORM|METHENAMINE|METHENAMINE
C2927961|T121|1007038|RXNORM|AFRICAN PYGEUM EXTRACT / STINGING NETTLE EXTRACT|AFRICAN PYGEUM EXTRACT / STINGING NETTLE EXTRACT
C2927962|T121|1007039|RXNORM|BETAMETHASONE / BETAMETHASONE ACETATE|BETAMETHASONE / BETAMETHASONE ACETATE
C0025646|T123|6837|RXNORM|METHIONINE|METHIONINE
C0025644|T121|6835|RXNORM|METHIMAZOLE|METHIMAZOLE
C0025641|T121|6834|RXNORM|METERGOLINE|METERGOLINE
C2927955|T121|1007032|RXNORM|BENTONITE / GOLDENSEAL EXTRACT / SYMPHYTUM UPLANDICUM LEAF EXTRACT|BENTONITE / GOLDENSEAL EXTRACT / SYMPHYTUM UPLANDICUM LEAF EXTRACT
C3486823|T121|1344644|RXNORM|ELYMUS REPENS TOP EXTRACT|ELYMUS REPENS TOP EXTRACT
C2927953|T121|1007030|RXNORM|ACETAMINOPHEN / TOLPERISONE|ACETAMINOPHEN / TOLPERISONE
C2927954|T121|1007031|RXNORM|CALCIUM LACTATE / MAGNESIUM SULFATE|CALCIUM LACTATE / MAGNESIUM SULFATE
C2927959|T121|1007036|RXNORM|CARBAMIDE PEROXIDE / EDETIC ACID|CARBAMIDE PEROXIDE / EDETIC ACID
C2927957|T121|1007034|RXNORM|ECHINACEA PURPUREA AERIAL PARTS EXTRACT / GOLDEN SEAL ROOT|ECHINACEA PURPUREA AERIAL PARTS EXTRACT / GOLDEN SEAL ROOT
C2927958|T121|1007035|RXNORM|DEQUALINIUM / LAURETH-9 / PREDNISOLONE|DEQUALINIUM / POLIDOCANOL / PREDNISOLONE
C1875662|T121|689760|RXNORM|PHOSPHORUS / POTASSIUM|PHOSPHORUS / POTASSIUM
C0040096|T121|10553|RXNORM|THYMOL|THYMOL
C1875520|T121|691433|RXNORM|NAPHAZOLINE / ZINC SULFATE|NAPHAZOLINE / ZINC SULFATE
C1875519|T121|691432|RXNORM|NAPHAZOLINE / PHENYLEPHRINE / PYRILAMINE|NAPHAZOLINE / PHENYLEPHRINE / PYRILAMINE
C2189662|T121|814044|RXNORM|ASCORBIC ACID / VINCAMINE|ASCORBIC ACID / VINCAMINE
C3818704|T122|1535631|RXNORM|GLYCERETH-7 TRIACETATE|GLYCERETH-7 TRIACETATE
C0602107|T121|156240|RXNORM|ETHYLNOREPINEPHRINE|ETHYLNOREPINEPHRINE
C1609686|T109|1293254|RXNORM|LUCINACTANT|LUCINACTANT
C3855135|T109|1547467|RXNORM|ARTEMISIA PRINCEPS LEAF OIL|ARTEMISIA PRINCEPS LEAF OIL
C3528058|T121|1361660|RXNORM|PICRASMA QUASSIOIDES WOOD EXTRACT|PICRASMA QUASSIOIDES WOOD EXTRACT
C0036113|T007|1329877|RXNORM|SALMONELLA ENTERICA SUBSP. ENTERICA SEROVAR ENTERITIDIS|SALMONELLA ENTERICA SUBSP. ENTERICA SEROVAR ENTERITIDIS
C3855133|T109|1547465|RXNORM|ACACIA CATECHU BARK EXTRACT|ACACIA CATECHU BARK EXTRACT
C0033603|T123|8826|RXNORM|PROTAMINES|PROTAMINES
C0075512|T195|37328|RXNORM|SULFAMETROLE|SULFAMETROLE
C0033602|T130|8825|RXNORM|PROTAMINE SULFATE (USP)|PROTAMINE SULFATE (USP)
C0075508|T121|37324|RXNORM|SULFAETHIDOLE|SULFAETHIDOLE
C3855136|T109|1547468|RXNORM|RUBIA CORDIFOLIA ROOT EXTRACT|RUBIA CORDIFOLIA ROOT EXTRACT
C0772056|T121|236749|RXNORM|BENPROPERINE|BENPROPERINE
C0543464|T121|142141|RXNORM|POTASSIUM AMINOBENZOATE|POTASSIUM AMINOBENZOATE
C0071836|T121|34369|RXNORM|PREDNICARBATE|PREDNICARBATE
C3695930|T109|1485121|RXNORM|BUTYL ACRYLATE - C16-C20 ALKYL METHACRYLATE - METHACRYLIC ACID - METHYL METHACRYLATE COPOLYMER|BUTYL ACRYLATE - C16-C20 ALKYL METHACRYLATE - METHACRYLIC ACID - METHYL METHACRYLATE COPOLYMER
C2948128|T121|1043468|RXNORM|DOCOSAHEXAENOATE / OMEGA-3 ACID ETHYL ESTERS (USP)|DOCOSAHEXAENOATE / OMEGA-3 ACID ETHYL ESTERS (USP)
C2709734|T129|854930|RXNORM|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 1 VACCINE|PNEUMOCOCCAL CAPSULAR POLYSACCHARIDE TYPE 1 VACCINE
C3464737|T121|1293032|RXNORM|LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS BULGARICUS|LACTOBACILLUS ACIDOPHILUS / LACTOBACILLUS BULGARICUS
C0969677|T127|237099|RXNORM|ALPHA TOCOPHEROL|ALPHA TOCOPHEROL
C0033473|T121|8770|RXNORM|PROPIOMAZINE|PROPIOMAZINE
C3555501|T121|1376150|RXNORM|HYDROXYETHYL CELLULOSE (40 MPA.S AT 2%)|HYDROXYETHYL CELLULOSE (40 MPA.S AT 2%)
C3555500|T109|1376151|RXNORM|LINGONBERRY SEED OIL|LINGONBERRY SEED OIL
C3555499|T122|1376152|RXNORM|PHENYLISOHEXANOL|PHENYLISOHEXANOL
C3555498|T121|1376153|RXNORM|TETRAHYDROBISDEMETHOXYDIFERULOYLMETHANE|TETRAHYDROBISDEMETHOXYDIFERULOYLMETHANE
C0961209|T121|298665|RXNORM|NEPAFENAC|NEPAFENAC
C2928849|T121|1007935|RXNORM|BENZOCAINE / LAPYRIUM / TYROTHRICIN|BENZOCAINE / LAPYRIUM / TYROTHRICIN
C3555495|T121|1376156|RXNORM|RIBOPRINE|RIBOPRINE
C3486566|T121|1311193|RXNORM|CORALLIUM RUBRUM EXOSKELETON PREPARATION|CORALLIUM RUBRUM EXOSKELETON PREPARATION
C3497911|T121|1311192|RXNORM|BOS TAURUS JOINT CAPSULE PREPARATION|BOVINE JOINT CAPSULE PREPARATION
C0114217|T121|1314347|RXNORM|DIOSMETIN|DIOSMETIN
C0018026|T196|1311190|RXNORM|GOLD|GOLD
C3256780|T121|1311197|RXNORM|LARICIFOMES OFFICINALIS FRUITING BODY EXTRACT|LARICIFOMES OFFICINALIS FRUITING BODY EXTRACT
C1816312|T121|1314340|RXNORM|CETEARYL ETHYLHEXANOATE|CETEARYL ETHYLHEXANOATE
C0255574|T121|1314343|RXNORM|CETYL MYRISTOLEATE|CETYL MYRISTOLEATE
C1576852|T109|1314342|RXNORM|CETETH-10 PHOSPHATE|CETETH-10 PHOSPHATE
C3489016|T121|1311199|RXNORM|SUS SCROFA PEYER'S PATCH PREPARATION|PORCINE SMALL INTESTINE MUCOSA LYMPH FOLLICLE PREPARATION
C0043684|T121|1314349|RXNORM|EDETOL|EDETOL
C3257293|T109|1314348|RXNORM|DIPROPYLENE GLYCOL DIBENZOATE|DIPROPYLENE GLYCOL DIBENZOATE
C3665091|T121|1435280|RXNORM|UNCARIA TOMENTOSA ROOT EXTRACT|UNCARIA TOMENTOSA ROOT EXTRACT
C3665092|T121|1435281|RXNORM|3-IODO-1-PROPANOL|3-IODO-1-PROPANOL
C0055444|T131|1435282|RXNORM|CHLOROPROPYLATE|CHLOROPROPYLATE
C3665093|T121|1435283|RXNORM|COCO MONOISOPROPANOLAMIDE|COCO MONOISOPROPANOLAMIDE
C2930097|T121|596050|RXNORM|CHOLINE / MAGNESIUM SALICYLATE|CHOLINE / MAGNESIUM SALICYLATE
C0047693|T121|1435286|RXNORM|M-PHENYLENEDIAMINE|M-PHENYLENEDIAMINE
C3665094|T121|1435288|RXNORM|CITRACONATE|CITRACONATE
C0038792|T121|10237|RXNORM|SULINDAC|SULINDAC
C2365882|T109|1305716|RXNORM|MANDARIN OIL|MANDARIN OIL
C0614705|T109|1426380|RXNORM|ETHYLHEXYL PALMITATE|ETHYLHEXYL PALMITATE
C0034616|T130|9133|RXNORM|SELENOMETHIONINE SE 75|SELENOMETHIONINE SE 75
C3489270|T121|1309929|RXNORM|TRIFOLIUM REPENS FLOWER EXTRACT|TRIFOLIUM REPENS FLOWER EXTRACT
C3489269|T121|1309928|RXNORM|SOLIDAGO CANADENSIS FLOWERING TOP EXTRACT|SOLIDAGO CANADENSIS FLOWERING TOP EXTRACT
C0073709|T123|35890|RXNORM|RUSCOGENIN|RUSCOGENIN
C2740751|T129|899645|RXNORM|BITTERNUT HICKORY POLLEN EXTRACT|CARYA CORDIFORMIS POLLEN EXTRACT
C0081408|T121|40575|RXNORM|ZILEUTON|ZILEUTON
C0011892|T131|3304|RXNORM|HEROIN|HEROIN
C2825368|T121|1145945|RXNORM|TOCERANIB|TOCERANIB
C2929413|T121|1008509|RXNORM|INSULIN, REGULAR, PORK / NPH INSULIN, PORK|INSULIN, ISOPHANE / INSULIN, REGULAR, PORK
C2929412|T121|1008508|RXNORM|ASCORBIC ACID / CALCIUM CITRATE / CHOLECALCIFEROL / CUPRIC OXIDE / DOCUSATE / FOLIC ACID / IRON CARBONYL / NIACINAMIDE / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC OXIDE|ASCORBIC ACID / CALCIUM CITRATE / CHOLECALCIFEROL / CUPRIC OXIDE / DOCUSATE / FOLIC ACID / IRON CARBONYL / NIACINAMIDE / POTASSIUM IODIDE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN A / VITAMIN B 12 / VITAMIN E / ZINC OXIDE
C3537764|T121|1371445|RXNORM|DODECAMETHYLPENTASILOXANE|DODECAMETHYLPENTASILOXANE
C2929407|T121|1008503|RXNORM|ASCORBIC ACID / FOLIC ACID / VITAMIN D|ASCORBIC ACID / FOLIC ACID / VITAMIN D
C2929406|T121|1008502|RXNORM|IBUPROFEN / PSEUDOISOCYTIDINE|IBUPROFEN / PSEUDOISOCYTIDINE
C2929405|T121|1008501|RXNORM|NPH INSULIN, HUMAN / REGULAR INSULIN, HUMAN|INSULIN, ISOPHANE / REGULAR INSULIN, HUMAN
C2929404|T121|1008500|RXNORM|ACETAMINOPHEN / BROMPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE|ACETAMINOPHEN / BROMPHENIRAMINE / DEXTROMETHORPHAN / PSEUDOEPHEDRINE
C2929411|T121|1008507|RXNORM|AGKISTRODON PISCIVORUS ANTIVENIN / CROTALUS ADAMANTEUS ANTIVENIN / CROTALUS ATROX ANTIVENIN / CROTALUS SCUTULATUS ANTIVENIN|AGKISTRODON PISCIVORUS ANTIVENIN / CROTALUS ADAMANTEUS ANTIVENIN / CROTALUS ATROX ANTIVENIN / CROTALUS SCUTULATUS ANTIVENIN
C2929410|T121|1008506|RXNORM|LINCOMYCIN / NIACIN|LINCOMYCIN / NIACIN
C2929408|T121|1008504|RXNORM|NIACIN / PENTIFYLLINE|NIACIN / PENTIFYLLINE
C2928218|T121|1007296|RXNORM|HISTAMINE / MENTHOL|HISTAMINE / MENTHOL
C3247723|T121|1192832|RXNORM|CAT HAIR EXTRACT / DOG HAIR EXTRACT|CAT HAIR EXTRACT / DOG HAIR EXTRACT
C2928216|T121|1007294|RXNORM|DEXCHLORPHENIRAMINE / METHSCOPOLAMINE / PHENYLEPHRINE|DEXCHLORPHENIRAMINE / METHSCOPOLAMINE / PHENYLEPHRINE
C3255960|T168|1312645|RXNORM|PAPAYA JUICE|PAPAYA JUICE
C2928214|T121|1007292|RXNORM|DIPHENHYDRAMINE / NIACIN|DIPHENHYDRAMINE / NIACIN
C2928215|T121|1007293|RXNORM|CODEINE / POTASSIUM|CODEINE / POTASSIUM
C2928212|T121|1007290|RXNORM|ACELLULAR PERTUSSIS VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY) / POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1) / POLIOVIRUS VACCINE INACTIVATED, TYPE 3 (SAUKETT) / TETANUS TOXOID VACCI|ACELLULAR PERTUSSIS VACCINE, INACTIVATED / DIPHTHERIA TOXOID VACCINE, INACTIVATED / POLIOVIRUS VACCINE INACTIVATED, TYPE 1 (MAHONEY) / POLIOVIRUS VACCINE INACTIVATED, TYPE 2 (MEF-1) / POLIOVIRUS VACCINE INACTIVATED, TYPE 3 (SAUKETT) / TETANUS TOXOID VACCINE, INACTIVATED
C2929839|T121|1008942|RXNORM|CHLORAMPHENICOL / PREDNISONE|CHLORAMPHENICOL / PREDNISONE
C0004609|T121|1292|RXNORM|BACLOFEN|BACLOFEN
C0004599|T195|1291|RXNORM|BACITRACIN|BACITRACIN
C0004599|T195|1291|RXNORM|BACITRACIN|BACITRACIN
C0004599|T195|1291|RXNORM|BACITRACIN|BACITRACIN
C2928220|T121|1007298|RXNORM|THIOCTATE / VITAMIN E|THIOCTATE / VITAMIN E
C2928221|T121|1007299|RXNORM|GLYCERYL MONOLAURATE / OLIVE LEAF EXTRACT|GLYCERYL MONOLAURATE / OLIVE LEAF EXTRACT
C3537763|T121|1371444|RXNORM|BOSWELLIA SACRA BARK EXTRACT|BOSWELLIA SACRA BARK EXTRACT
C3857953|T197|1552046|RXNORM|LEAD MONOSILICATE|LEAD MONOSILICATE
C0249458|T121|73645|RXNORM|VALACYCLOVIR|VALACYCLOVIR
C3473979|T121|1299865|RXNORM|CAMPHOR / TURPENTINE|CAMPHOR / TURPENTINE
C0063322|T121|27392|RXNORM|TROPISETRON|TROPISETRON
C1443691|T121||RXNORM|CIPROFLOXACIN / DEXAMETHASONE
C0072732|T121|35097|RXNORM|PYRISUCCIDEANOL|PIRISUDANOL
C0064324|T121|28198|RXNORM|KEBUZONE|KEBUZONE
C1995590|T121|751543|RXNORM|COLLAGEN,ACTIVATED|COLLAGEN,ACTIVATED
C2718454|T121|858027|RXNORM|GLYCERIN / NAPHAZOLINE|GLYCERIN / NAPHAZOLINE
C0002520|T123||RXNORM|AMINO ACIDS
C0002520|T121||RXNORM|AMINO ACIDS
C0002520|T116||RXNORM|AMINO ACIDS
C0005492|T127||RXNORM|BIOFLAVONOIDS
C0005492|T121||RXNORM|BIOFLAVONOIDS
C0005492|T109||RXNORM|BIOFLAVONOIDS
C0016388|T127|1925821|RXNORM|FLAVIN MONONUCLEOTIDE|RIBOFLAVIN 5'-PHOSPHATE
C0016388|T121|1925821|RXNORM|FLAVIN MONONUCLEOTIDE|RIBOFLAVIN 5'-PHOSPHATE
C0016388|T114|1925821|RXNORM|FLAVIN MONONUCLEOTIDE|RIBOFLAVIN 5'-PHOSPHATE
C0072733|T197|1544140|RXNORM|PYRITE|FERROUS DISULFIDE
C0075629|T195||RXNORM|SULTAMICILLIN
C0075629|T109||RXNORM|SULTAMICILLIN
C0145918|T121||RXNORM|CLAVULANIC ACID / TICARCILLIN
C0717902|T121||RXNORM|MALT SOUP EXTRACT / PSYLLIUM
C0873197|T116|285170|RXNORM|YELLOW JACKET VEN PROTEIN|YELLOW JACKET VENOM PROTEIN
C0873197|T121|285170|RXNORM|YELLOW JACKET VEN PROTEIN|YELLOW JACKET VENOM PROTEIN
C0982043|T121||RXNORM|CITRUS BIOFLAVONOIDS
C0982043|T109||RXNORM|CITRUS BIOFLAVONOIDS
C1273035|T109||RXNORM|CARBOMER-980
C1273035|T121||RXNORM|CARBOMER-980
C1329980|T121||RXNORM|ASPIRIN / PRAVASTATIN
C1329986|T121||RXNORM|BUPIVACAINE / FENTANYL
C1329986|T121||RXNORM|BUPIVACAINE / FENTANYL
C1337136|T121||RXNORM|L-METHYLFOLATE
C1337136|T127||RXNORM|L-METHYLFOLATE
C1337136|T109||RXNORM|L-METHYLFOLATE
C0981839|T129|1742530|RXNORM|ASPERGILLUS NIGER EXTRACT|ASPERGILLUS NIGER ALLERGENIC EXTRACT
C0981839|T121|1742530|RXNORM|ASPERGILLUS NIGER EXTRACT|ASPERGILLUS NIGER ALLERGENIC EXTRACT
C0872901|T007||RXNORM|LACTOBACILLUS SPOROGENES
C1602511|T109||RXNORM|IBADRONATE
C1602511|T121||RXNORM|IBADRONATE
C1875386|T121||RXNORM|IODINE / POTASSIUM IODIDE / ZINC PHENOLSULFONATE
C0303918|T109||RXNORM|INSOLUBLE BERLIN BLUE STAIN
C0303918|T130||RXNORM|INSOLUBLE BERLIN BLUE STAIN
C1950494|T121||RXNORM|BUPIVACAINE / HYDROMORPHONE
C1950494|T121||RXNORM|BUPIVACAINE / HYDROMORPHONE
C2112883|T121||RXNORM|ASCORBIC ACID / POTASSIUM CHLORIDE
C1110640|T121||RXNORM|HOUSE DUST MITE EXTRACT, DERMATOPHAGOIDES FARINAE
C1110640|T129||RXNORM|HOUSE DUST MITE EXTRACT, DERMATOPHAGOIDES FARINAE
C0446330|T121||RXNORM|HOUSE DUST MITE EXTRACT, DERMATOPHAGOIDES PTERONYSSINUS
C0446330|T129||RXNORM|HOUSE DUST MITE EXTRACT, DERMATOPHAGOIDES PTERONYSSINUS
C2702308|T129||RXNORM|ACACIA LONGIFOLIA POLLEN EXTRACT
C2702308|T121||RXNORM|ACACIA LONGIFOLIA POLLEN EXTRACT
C2756337|T121||RXNORM|BAKER'S YEAST (SACCHAROMYCES CEREVISIAE) ALLERGENIC EXTRACT
C2756337|T129||RXNORM|BAKER'S YEAST (SACCHAROMYCES CEREVISIAE) ALLERGENIC EXTRACT
C2930257|T025||RXNORM|AUTOLOGOUS CULTURED CHONDROCYTES
C2927943|T121||RXNORM|BIOFLAVONOIDS / HORSE CHESTNUT PREPARATION
C2927945|T121||RXNORM|BIOFLAVONOIDS / PENTOXIFYLLINE
C2927947|T121||RXNORM|ASCORBIC ACID / CITRUS BIOFLAVONOIDS
C2927963|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / HESPERIDIN
C2927964|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / HESPERIDIN / RUTIN
C2927989|T121||RXNORM|BIOFLAVONOIDS / QUERCETIN / VITIS EXTRACT
C2927993|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / CALCIUM ASCORBATE
C2927995|T121||RXNORM|ACEXAMIC ACID / GENTAMICIN SULFATE (USP)
C2928114|T121||RXNORM|SODIUM PHOSPHATE, DIBASIC, ANHYDROUS / SODIUM PHOSPHATE,MONOBASIC,MONOHYDRATE / TRIBASIC POTASSIUM PHOSPHATE
C2928167|T121||RXNORM|THYROXINE / TRIIODOTHYRONINE
C2928228|T121||RXNORM|BIOFLAVONOIDS / GRAPE SEED EXTRACT
C2928283|T121||RXNORM|PAPAVERINE / PHENTOLAMINE
C2928549|T121||RXNORM|DIETHYLSTILBESTROL / LACTATE
C2928596|T121||RXNORM|BUPIVACAINE / MEPERIDINE
C2928646|T121||RXNORM|GENTAMICIN SULFATE (USP) / PREDNISOLONE
C2928646|T121||RXNORM|GENTAMICIN SULFATE (USP) / PREDNISOLONE
C2928668|T121||RXNORM|RACEPINEPHRINE / ZINC PHENOLSULFONATE
C2928741|T121||RXNORM|AMINOPHYLLINE / GUAIFENESIN / PHENOBARBITAL
C2928741|T121||RXNORM|AMINOPHYLLINE / GUAIFENESIN / PHENOBARBITAL
C2928753|T121||RXNORM|SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE,MONOBASIC,MONOHYDRATE
C2928930|T121||RXNORM|BETAMETHASONE / GENTAMICIN SULFATE (USP) / TOLNAFTATE
C2928983|T121||RXNORM|HEPARIN / ZINC SULFATE
C2929033|T121||RXNORM|FRUIT EXTRACTS / LUTEIN / LYCOPENE
C2929173|T121||RXNORM|ERGOCALCIFEROL / GENTAMICIN SULFATE (USP)
C2929183|T121||RXNORM|CITRIC ACID / MAGNESIUM CARBONATE / POTASSIUM CITRATE
C2929242|T121||RXNORM|AMMONIUM PHOSPHATE / DISODIUM PYROPHOSPHATE / SODIUM PHOSPHATE, MONOBASIC
C2929266|T121||RXNORM|BETAMETHASONE / VITAMIN B 12
C2929292|T121||RXNORM|CALCIUM CHLORIDE / GLUCOSE / MAGNESIUM SULFATE / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE / SODIUM PHOSPHATE
C2929298|T121||RXNORM|POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC, ANHYDROUS
C2929409|T121||RXNORM|GENTAMICIN SULFATE (USP) / HYDROCORTISONE
C2929422|T121||RXNORM|DIBASIC POTASSIUM PHOSPHATE / SODIUM PHOSPHATE,MONOBASIC,MONOHYDRATE
C2929587|T121||RXNORM|BETAMETHASONE / GENTAMICIN SULFATE (USP)
C2929611|T121||RXNORM|GLUCOSE / HEPARIN
C2929626|T121||RXNORM|DIFLORASONE / GENTAMICIN SULFATE (USP)
C2929641|T121||RXNORM|FLUOROMETHOLONE / GENTAMICIN SULFATE (USP)
C2929642|T121||RXNORM|BETAMETHASONE / GENTAMICIN SULFATE (USP) / MICONAZOLE
C2929661|T121||RXNORM|BIOFLAVONOIDS / GRAPE SEED PROANTHOCYANIDINS
C2929697|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / GRAPE SEED EXTRACT
C2929704|T121||RXNORM|OMEGA-3 ACID ETHYL ESTERS (USP) / VITAMIN E
C2929741|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / ECHINACEA PREPARATION
C2929785|T121||RXNORM|FLUPREDNIDENE / GENTAMICIN SULFATE (USP)
C2929825|T121||RXNORM|GENTAMICIN SULFATE (USP) / HYDROCORTISONE / KETOCONAZOLE
C2929866|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOID, LEMON / ECHINACEA PREPARATION
C2978449|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / CHOLINE / INOSITOL / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C3160611|T121||RXNORM|GLYCERIN / PANTHENOL / VITAMIN E
C3190699|T121||RXNORM|ACETYLCYSTEINE / L-METHYLFOLATE / MECOBALAMIN
C3204800|T121||RXNORM|DEXTRANOMER / HYALURONATE
C3244536|T121||RXNORM|DIPHENHYDRAMINE / HYDROCORTISONE / NYSTATIN / TETRACYCLINE
C3244536|T121||RXNORM|DIPHENHYDRAMINE / HYDROCORTISONE / NYSTATIN / TETRACYCLINE
C3244757|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / BROMELAINS / QUERCETIN
C3247717|T121||RXNORM|BUPIVACAINE / SUFENTANIL
C3247717|T121||RXNORM|BUPIVACAINE / SUFENTANIL
C3248019|T121||RXNORM|MAGNESIUM CITRATE / SIMETHICONE
C3249779|T121||RXNORM|BUPIVACAINE / EPINEPHRINE / FENTANYL
C3249779|T121||RXNORM|BUPIVACAINE / EPINEPHRINE / FENTANYL
C3265664|T121||RXNORM|GENTAMICIN SULFATE (USP) / HYDROCORTISONE / MICONAZOLE
C3268132|T121||RXNORM|ALUMINUM HYDROXIDE / DIPHENHYDRAMINE / LIDOCAINE / MAGNESIUM HYDROXIDE / SIMETHICONE
C3268132|T121||RXNORM|ALUMINUM HYDROXIDE / DIPHENHYDRAMINE / LIDOCAINE / MAGNESIUM HYDROXIDE / SIMETHICONE
C3268139|T121||RXNORM|DIPHENHYDRAMINE / HYDROCORTISONE / NYSTATIN
C3268139|T121||RXNORM|DIPHENHYDRAMINE / HYDROCORTISONE / NYSTATIN
C0002520|T123||RXNORM|AMINO ACIDS
C0002520|T121||RXNORM|AMINO ACIDS
C0002520|T116||RXNORM|AMINO ACIDS
C0005492|T127||RXNORM|BIOFLAVONOIDS
C0005492|T121||RXNORM|BIOFLAVONOIDS
C0005492|T109||RXNORM|BIOFLAVONOIDS
C0016388|T127|1925821|RXNORM|FLAVIN MONONUCLEOTIDE|RIBOFLAVIN 5'-PHOSPHATE
C0016388|T121|1925821|RXNORM|FLAVIN MONONUCLEOTIDE|RIBOFLAVIN 5'-PHOSPHATE
C0016388|T114|1925821|RXNORM|FLAVIN MONONUCLEOTIDE|RIBOFLAVIN 5'-PHOSPHATE
C0072733|T197|1544140|RXNORM|PYRITE|FERROUS DISULFIDE
C0075629|T195||RXNORM|SULTAMICILLIN
C0075629|T109||RXNORM|SULTAMICILLIN
C0145918|T121||RXNORM|CLAVULANIC ACID / TICARCILLIN
C0717902|T121||RXNORM|MALT SOUP EXTRACT / PSYLLIUM
C0873197|T116|285170|RXNORM|YELLOW JACKET VEN PROTEIN|YELLOW JACKET VENOM PROTEIN
C0873197|T121|285170|RXNORM|YELLOW JACKET VEN PROTEIN|YELLOW JACKET VENOM PROTEIN
C0982043|T121||RXNORM|CITRUS BIOFLAVONOIDS
C0982043|T109||RXNORM|CITRUS BIOFLAVONOIDS
C1273035|T109||RXNORM|CARBOMER-980
C1273035|T121||RXNORM|CARBOMER-980
C1329980|T121||RXNORM|ASPIRIN / PRAVASTATIN
C1329986|T121||RXNORM|BUPIVACAINE / FENTANYL
C1329986|T121||RXNORM|BUPIVACAINE / FENTANYL
C1337136|T121||RXNORM|L-METHYLFOLATE
C1337136|T127||RXNORM|L-METHYLFOLATE
C1337136|T109||RXNORM|L-METHYLFOLATE
C0981839|T129|1742530|RXNORM|ASPERGILLUS NIGER EXTRACT|ASPERGILLUS NIGER ALLERGENIC EXTRACT
C0981839|T121|1742530|RXNORM|ASPERGILLUS NIGER EXTRACT|ASPERGILLUS NIGER ALLERGENIC EXTRACT
C0872901|T007||RXNORM|LACTOBACILLUS SPOROGENES
C1602511|T109||RXNORM|IBADRONATE
C1602511|T121||RXNORM|IBADRONATE
C1875386|T121||RXNORM|IODINE / POTASSIUM IODIDE / ZINC PHENOLSULFONATE
C0303918|T109||RXNORM|INSOLUBLE BERLIN BLUE STAIN
C0303918|T130||RXNORM|INSOLUBLE BERLIN BLUE STAIN
C1950494|T121||RXNORM|BUPIVACAINE / HYDROMORPHONE
C1950494|T121||RXNORM|BUPIVACAINE / HYDROMORPHONE
C2112883|T121||RXNORM|ASCORBIC ACID / POTASSIUM CHLORIDE
C1110640|T121||RXNORM|HOUSE DUST MITE EXTRACT, DERMATOPHAGOIDES FARINAE
C1110640|T129||RXNORM|HOUSE DUST MITE EXTRACT, DERMATOPHAGOIDES FARINAE
C0446330|T121||RXNORM|HOUSE DUST MITE EXTRACT, DERMATOPHAGOIDES PTERONYSSINUS
C0446330|T129||RXNORM|HOUSE DUST MITE EXTRACT, DERMATOPHAGOIDES PTERONYSSINUS
C2702308|T129||RXNORM|ACACIA LONGIFOLIA POLLEN EXTRACT
C2702308|T121||RXNORM|ACACIA LONGIFOLIA POLLEN EXTRACT
C2756337|T121||RXNORM|BAKER'S YEAST (SACCHAROMYCES CEREVISIAE) ALLERGENIC EXTRACT
C2756337|T129||RXNORM|BAKER'S YEAST (SACCHAROMYCES CEREVISIAE) ALLERGENIC EXTRACT
C2930257|T025||RXNORM|AUTOLOGOUS CULTURED CHONDROCYTES
C2927943|T121||RXNORM|BIOFLAVONOIDS / HORSE CHESTNUT PREPARATION
C2927945|T121||RXNORM|BIOFLAVONOIDS / PENTOXIFYLLINE
C2927947|T121||RXNORM|ASCORBIC ACID / CITRUS BIOFLAVONOIDS
C2927963|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / HESPERIDIN
C2927964|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / HESPERIDIN / RUTIN
C2927989|T121||RXNORM|BIOFLAVONOIDS / QUERCETIN / VITIS EXTRACT
C2927993|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / CALCIUM ASCORBATE
C2927995|T121||RXNORM|ACEXAMIC ACID / GENTAMICIN SULFATE (USP)
C2928114|T121||RXNORM|SODIUM PHOSPHATE, DIBASIC, ANHYDROUS / SODIUM PHOSPHATE,MONOBASIC,MONOHYDRATE / TRIBASIC POTASSIUM PHOSPHATE
C2928167|T121||RXNORM|THYROXINE / TRIIODOTHYRONINE
C2928228|T121||RXNORM|BIOFLAVONOIDS / GRAPE SEED EXTRACT
C2928283|T121||RXNORM|PAPAVERINE / PHENTOLAMINE
C2928549|T121||RXNORM|DIETHYLSTILBESTROL / LACTATE
C2928596|T121||RXNORM|BUPIVACAINE / MEPERIDINE
C2928646|T121||RXNORM|GENTAMICIN SULFATE (USP) / PREDNISOLONE
C2928646|T121||RXNORM|GENTAMICIN SULFATE (USP) / PREDNISOLONE
C2928668|T121||RXNORM|RACEPINEPHRINE / ZINC PHENOLSULFONATE
C2928741|T121||RXNORM|AMINOPHYLLINE / GUAIFENESIN / PHENOBARBITAL
C2928741|T121||RXNORM|AMINOPHYLLINE / GUAIFENESIN / PHENOBARBITAL
C2928753|T121||RXNORM|SODIUM PHOSPHATE, DIBASIC / SODIUM PHOSPHATE,MONOBASIC,MONOHYDRATE
C2928930|T121||RXNORM|BETAMETHASONE / GENTAMICIN SULFATE (USP) / TOLNAFTATE
C2928983|T121||RXNORM|HEPARIN / ZINC SULFATE
C2929033|T121||RXNORM|FRUIT EXTRACTS / LUTEIN / LYCOPENE
C2929173|T121||RXNORM|ERGOCALCIFEROL / GENTAMICIN SULFATE (USP)
C2929183|T121||RXNORM|CITRIC ACID / MAGNESIUM CARBONATE / POTASSIUM CITRATE
C2929242|T121||RXNORM|AMMONIUM PHOSPHATE / DISODIUM PYROPHOSPHATE / SODIUM PHOSPHATE, MONOBASIC
C2929266|T121||RXNORM|BETAMETHASONE / VITAMIN B 12
C2929292|T121||RXNORM|CALCIUM CHLORIDE / GLUCOSE / MAGNESIUM SULFATE / POTASSIUM CHLORIDE / SODIUM BICARBONATE / SODIUM CHLORIDE / SODIUM PHOSPHATE
C2929298|T121||RXNORM|POTASSIUM PHOSPHATE / SODIUM PHOSPHATE, MONOBASIC, ANHYDROUS
C2929409|T121||RXNORM|GENTAMICIN SULFATE (USP) / HYDROCORTISONE
C2929422|T121||RXNORM|DIBASIC POTASSIUM PHOSPHATE / SODIUM PHOSPHATE,MONOBASIC,MONOHYDRATE
C2929587|T121||RXNORM|BETAMETHASONE / GENTAMICIN SULFATE (USP)
C2929611|T121||RXNORM|GLUCOSE / HEPARIN
C2929626|T121||RXNORM|DIFLORASONE / GENTAMICIN SULFATE (USP)
C2929641|T121||RXNORM|FLUOROMETHOLONE / GENTAMICIN SULFATE (USP)
C2929642|T121||RXNORM|BETAMETHASONE / GENTAMICIN SULFATE (USP) / MICONAZOLE
C2929661|T121||RXNORM|BIOFLAVONOIDS / GRAPE SEED PROANTHOCYANIDINS
C2929697|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / GRAPE SEED EXTRACT
C2929704|T121||RXNORM|OMEGA-3 ACID ETHYL ESTERS (USP) / VITAMIN E
C2929741|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / ECHINACEA PREPARATION
C2929785|T121||RXNORM|FLUPREDNIDENE / GENTAMICIN SULFATE (USP)
C2929825|T121||RXNORM|GENTAMICIN SULFATE (USP) / HYDROCORTISONE / KETOCONAZOLE
C2929866|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOID, LEMON / ECHINACEA PREPARATION
C2978449|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / CHOLINE / INOSITOL / NIACINAMIDE / PANTOTHENATE / PYRIDOXINE / RIBOFLAVIN / THIAMINE / VITAMIN B 12
C3160611|T121||RXNORM|GLYCERIN / PANTHENOL / VITAMIN E
C3190699|T121||RXNORM|ACETYLCYSTEINE / L-METHYLFOLATE / MECOBALAMIN
C3204800|T121||RXNORM|DEXTRANOMER / HYALURONATE
C3244536|T121||RXNORM|DIPHENHYDRAMINE / HYDROCORTISONE / NYSTATIN / TETRACYCLINE
C3244536|T121||RXNORM|DIPHENHYDRAMINE / HYDROCORTISONE / NYSTATIN / TETRACYCLINE
C3244757|T121||RXNORM|ASCORBIC ACID / BIOFLAVONOIDS / BROMELAINS / QUERCETIN
C3247717|T121||RXNORM|BUPIVACAINE / SUFENTANIL
C3247717|T121||RXNORM|BUPIVACAINE / SUFENTANIL
C3248019|T121||RXNORM|MAGNESIUM CITRATE / SIMETHICONE
C3249779|T121||RXNORM|BUPIVACAINE / EPINEPHRINE / FENTANYL
C3249779|T121||RXNORM|BUPIVACAINE / EPINEPHRINE / FENTANYL
C3265664|T121||RXNORM|GENTAMICIN SULFATE (USP) / HYDROCORTISONE / MICONAZOLE
C0043393|T004||RXNORM|YEASTS
C0074071|T121|1364901|RXNORM|SARKOSYL|SODIUM LAUROYL SARCOSINATE
C0873035|T121||RXNORM|ENZYMES,DIGESTIVE (PLANT)
C0981923|T121||RXNORM|ALLERGENIC EXTRACT, MAPLE
C0981929|T121||RXNORM|ALLERGENIC EXTRACT, MOUNTAIN CEDAR
C0981932|T121||RXNORM|ALLERGENIC EXTRACT, MUCOR RACEMOSUS MOLD
C0981933|T121||RXNORM|ALLERGENIC EXTRACT, OAK
C0981935|T121||RXNORM|ALLERGENIC EXTRACT, OLIVE
C0981938|T121||RXNORM|ALLERGENIC EXTRACT, PENICILLIN
C0981941|T121||RXNORM|ALLERGENIC EXTRACT, PHOMA BETAE MOLD
C0981942|T121||RXNORM|ALLERGENIC EXTRACT, PIGWEED, ROUGH
C0981945|T121||RXNORM|ALLERGENIC EXTRACT, PLANTAIN, ENGLISH
C0981948|T121||RXNORM|ALLERGENIC EXTRACT, POPLAR
C0981949|T121||RXNORM|ALLERGENIC EXTRACT, POPULUS ALBA, P. DELTOIDES
C0981966|T121||RXNORM|ALLERGENIC EXTRACT, SCALE MIX
C0981967|T121||RXNORM|ALLERGENIC EXTRACT, SHEEP SORREL
C0981968|T121||RXNORM|ALLERGENIC EXTRACT, SHEEP WOOL
C0981973|T121||RXNORM|ALLERGENIC EXTRACT, STEMPHYLLUM BOTRYOSUM MOLD
C0981974|T121||RXNORM|ALLERGENIC EXTRACT, STINGING INSECT
C0981979|T121||RXNORM|ALLERGENIC EXTRACT, SYCAMORE
C0991781|T121||RXNORM|ALLERGENIC EXTRACT, LAMB QUARTERS
C0991782|T121||RXNORM|ALLERGENIC EXTRACT, MESQUITE
C0991788|T121||RXNORM|ALLERGENIC EXTRACT, THISTLE, RUSSIAN
C0991790|T121||RXNORM|ALLERGENIC EXTRACT, WEED, CARELESS
C0991792|T121||RXNORM|ALLERGENIC EXTRACT,AGARICUS CAMPESTRIS
C0993207|T121||RXNORM|ALLERGENIC EXTRACT, RAGWEED STOCK POLLEN
C2017850|T121||RXNORM|SAFFLOWER OIL / SOYBEAN OIL
C2138494|T121||RXNORM|CROMOLYN / NAPHAZOLINE
C2193935|T121||RXNORM|NAPHAZOLINE / PREDNISOLONE
C2347615|T121|1999323|RXNORM|PLUMERIA EXTRACT|PLUMERIA ALBA FLOWER EXTRACT
C3256328|T121||RXNORM|AMINO ACIDS, WHEAT
C3256597|T121|1307719|RXNORM|ATRACTYLODES JAPONICA ROOT|ATRACTYLODES JAPONICA ROOT EXTRACT
C3538555|T109|1373037|RXNORM|TUMERIC OIL|TURMERIC OIL
C3864844|T109|1747570|RXNORM|ALLYL METHACRYLATE/GLYCOL DIMETHACRYLATE CROSSPOLYMER|ALLYL METHACRYLATE-GLYCOL DIMETHACRYLATE CROSSPOLYMER
C0108406|T109||RXNORM|CARBOMER HOMOPOLYMER TYPE B
C0991774|T121||RXNORM|ALLERGENIC EXTRACT, COMMON MUGWORT
C1703487|T121||RXNORM|HYALURONIDASE, HUMAN
C2927885|T121||RXNORM|HYALURONIDASE / LIDOCAINE
C2927902|T121||RXNORM|CAMPHOR / GLYCOL SALICYLATE / MENTHOL
C2928028|T121||RXNORM|NITROFURAZONE / XYLOMETAZOLINE
C2928115|T121||RXNORM|PHOSPHOLIPIDS / SOYBEAN OIL
C2928385|T121||RXNORM|CHOLINE / YEASTS
C2928462|T121||RXNORM|EGG YOLK PHOSPHATIDES / GLYCERIN / SAFFLOWER OIL / SOYBEAN PREPARATION
C2928705|T121||RXNORM|BEESWAX / BOSWELLIA PREPARATION / MOMORDICAE / MYRRH EXTRACT
C2928737|T121||RXNORM|TINIDAZOLE / TIOCONAZOLE
C2928997|T121||RXNORM|LAUROMACROGOLS / SOYBEAN OIL
C2929191|T121||RXNORM|EGG YOLK PHOSPHOLIPIDS / GLYCERIN / SAFFLOWER OIL / SOYBEAN OIL
C2929300|T121||RXNORM|ALBUMIN,AGGREGATED / STANNOUS CHLORIDE / TIN
C2929431|T121||RXNORM|EGG YOLK PHOSPHOLIPIDS / GLYCERIN / SOYBEAN OIL
C2929538|T121||RXNORM|PHOSPHOLIPIDS / SOYBEAN PREPARATION
C2929676|T121||RXNORM|EGG YOLK PHOSPHATIDES / GLYCERIN / SOYBEAN PREPARATION
C2929693|T121||RXNORM|CYCLOBENZAPRINE / METHYLSULFONYLMETHANE
C3265067|T121||RXNORM|CALCIUM CARBONATE / VITAMIN D3
C3267609|T121||RXNORM|LACTOSE / SACCHAROMYCES BOULARDII LYO
C3281532|T121||RXNORM|STEMMACANTHA CARTHAMOIDES ROOT EXTRACT
C3472881|T121||RXNORM|BALD-FACED HORNET VENOM PROTEIN / COMMON WASP VENOM PROTEIN / EASTERN YELLOWJACKET VENOM PROTEIN / GERMAN WASP VENOM PROTEIN / SOUTHERN YELLOWJACKET VENOM PROTEIN / WESTERN YELLOWJACKET VENOM PROTEIN / YELLOW HORNET VENOM PROTEIN
C3472899|T121||RXNORM|COMMON WASP VENOM PROTEIN / EASTERN YELLOWJACKET VENOM PROTEIN / GERMAN WASP VENOM PROTEIN / SOUTHERN YELLOWJACKET VENOM PROTEIN / WESTERN YELLOWJACKET VENOM PROTEIN
C3651742|T121||RXNORM|KONJAC MANNAN
C3651793|T121||RXNORM|STYRAX BENZOIN RESIN
C3693129|T121||RXNORM|ALPHA TOCOPHEROL / GLYCOL SALICYLATE / MENTHOL / NONIVAMIDE
C3700995|T121||RXNORM|ALPHA TOCOPHEROL / ASCORBIC ACID / DOCONEXENT / DOCUSATE / FERROUS FUMARATE / FOLIC ACID / PYRIDOXINE / TRICALCIUM PHOSPHATE
C3819184|T121||RXNORM|BORNEOL / MENTHOL
