67162-8|T077|strict|67162-8|LNC|PATIENT DISPOSITION|PATIENT DISPOSITION
67162-8|T077|strict|67162-8|LNC|DISPOSITION|DISPOSITION
67162-8|T077|strict|67162-8|LNC|PATIENT DISPOSITION|PATIENT DISPOSITION
67162-8|T077|strict|67162-8|LNC|DISPOSITION ON DISCHARGE|DISPOSITION ON DISCHARGE
67162-8|T077|strict|67162-8|LNC|DISCHARGE DISPOSITION|DISCHARGE DISPOSITION
67162-8|T077|strict|67162-8|LNC|POSTPARTUM DISPOSITION|POSTPARTUM DISPOSITION
67162-8|T077|strict|67162-8|LNC|PROCEDURE DISPOSITION|PROCEDURE DISPOSITION
78033-8|T077|strict|78033-8|LNC|HOSPITAL STAY DURATION|HOSPITAL STAY DURATION
78033-8|T077|multi|78033-8|LNC|LOS|LOS
78033-8|T077|strict|78033-8|LNC|LENGTH OF STAY|LENGTH OF STAY
78033-8|T077|strict|78033-8|LNC|HOSPITALIZATION STAY|HOSPITALIZATION STAY
46240-8|T077|strict|46240-8|LNC|HISTORY OF HOSPITALIZATION|HISTORY OF HOSPITALIZATION
46240-8|T077|strict|46240-8|LNC|HISTORY OF HOSPITALIZATIONS|HISTORY OF HOSPITALIZATIONS
46240-8|T077|strict|46240-8|LNC|HX OF HOSPITALIZATION|HX OF HOSPITALIZATION
46240-8|T077|strict|46240-8|LNC|HOSPITALIZATION/MAJOR|HOSPITALIZATION/MAJOR
46240-8|T077|strict|46240-8|LNC|HOSPITALIZATIONS|HOSPITALIZATIONS
46240-8|T077|multi|46240-8|LNC|HOSPITALIZATION|HOSPITALIZATION
46240-8|T077|strict|46240-8|LNC|HISTORY OF ENCOUNTERS|HISTORY OF ENCOUNTERS
46240-8|T077|multi|46240-8|LNC|EPISODES|EPISODES
11347-2|T077|strict|11347-2|LNC|HISTORY OF OUTPATIENT VISITS|HISTORY OF OUTPATIENT VISITS
11347-2|T077|strict|11347-2|LNC|OUTPATIENT VISITS|OUTPATIENT VISITS
11347-2|T077|strict|11347-2|LNC|OUTPATIENT VISIT|OUTPATIENT VISIT
11347-2|T077|multi|11347-2|LNC|OUTPATIENT|OUTPATIENT
52536-0|T077|strict|52536-0|LNC|ADMISSION INFORMATION|ADMISSION INFORMATION
34111-5|T077|strict|34111-5|LNC|EMERGENCY DEPARTMENT|EMERGENCY DEPARTMENT
34111-5|T077|strict|34111-5|LNC|EMERGENCY VISITS|EMERGENCY VISITS
34111-5|T077|strict|34111-5|LNC|EMERGENCY VISIT|EMERGENCY VISIT
34111-5|T077|strict|34111-5|LNC|ED VISITS|ED VISITS
34111-5|T077|strict|34111-5|LNC|ED VISIT|ED VISIT
34111-5|T077|strict|34111-5|LNC|ER VISIT|ER VISIT
75504-1|T077|strict|75504-1|LNC|URGENT CARE CENTER|URGENT CARE CENTER
75504-1|T077|strict|75504-1|LNC|URGENT CARE VISIT|URGENT CARE VISIT
75504-1|T077|strict|75504-1|LNC|URGENT CARE ENCOUNTER|URGENT CARE ENCOUNTER
85208-7|T077|strict|85208-7|LNC|TELEHEALTH CONSULT|TELEHEALTH CONSULT
85208-7|T077|strict|85208-7|LNC|TELEMEDECINE|TELEMEDECINE
85208-7|T077|strict|85208-7|LNC|VIRTUAL|VIRTUAL
76427-4|T077|strict|76427-4|LNC|VISIT DATE|VISIT DATE
76427-4|T077|strict|76427-4|LNC|DATE OF VISIT|DATE OF VISIT
76427-4|T077|strict|76427-4|LNC|ENCOUNTER DATE|ENCOUNTER DATE
76427-4|T077|strict|76427-4|LNC|ENC DATE|ENC DATE
76427-4|T077|strict|76427-4|LNC|REGISTRATION DATE|REGISTRATION DATE
76427-4|T077|strict|76427-4|LNC|SERVICE DATE|SERVICE DATE
76427-4|T077|strict|76427-4|LNC|DATE ISSUED|DATE ISSUED
76427-4|T077|strict|76427-4|LNC|REPORT DATE|REPORT DATE
76427-4|T077|strict|76427-4|LNC|RECORD DATE|RECORD DATE
76427-4|T077|strict|76427-4|LNC|STUDY DATE|STUDY DATE
76427-4|T077|strict|76427-4|LNC|EPISODE DATE|EPISODE DATE
76427-4|T077|strict|76427-4|LNC|TODAY IS|TODAY IS
76427-4|T077|strict|76427-4|LNC|DATE TIME|DATE TIME
76427-4|T077|strict|76427-4|LNC|DATE|DATE
91582-7|T077|strict|91582-7|LNC|REPORT STATUS|REPORT STATUS
91582-7|T077|strict|91582-7|LNC|REPORT STAGE|REPORT STAGE
91582-7|T077|strict|91582-7|LNC|DOCUMENT STATUS|DOCUMENT STATUS
52455-3|T077|strict|52455-3|LNC|ADMISSION DATE|ADMISSION DATE
52455-3|T077|strict|52455-3|LNC|ADMISSION DATA|ADMISSION DATA
52525-3|T077|strict|52525-3|LNC|DISCHARGE DATE|DISCHARGE DATE
52525-3|T077|strict|52525-3|LNC|DISCHARGE DATE/TIME|DISCHARGE DATE/TIME
52525-3|T077|strict|52525-3|LNC|DISCHARGE TIME|DISCHARGE TIME
52525-3|T077|strict|52525-3|LNC|DISCHARGE DATE TIME|DISCHARGE DATE TIME
52525-3|T077|strict|52525-3|LNC|DISCHARGE DATETIME|DISCHARGE DATETIME
52525-3|T077|strict|52525-3|LNC|DATE OF DISCHARGE|DATE OF DISCHARGE
92707-9|T077|strict|92707-9|LNC|CARE TEAM|CARE TEAM
92707-9|T077|strict|92707-9|LNC|TREATMENT TEAM|TREATMENT TEAM
92707-9|T077|strict|92707-9|LNC|CARE PROVIDER|CARE PROVIDER
92707-9|T077|multi|92707-9|LNC|PROVIDER|PROVIDER
92707-9|T077|strict|92707-9|LNC|PHYSICIAN|PHYSICIAN
92707-9|T077|strict|92707-9|LNC|DOCTOR|DOCTOR
92707-9|T077|strict|92707-9|LNC|NURSE|NURSE
92707-9|T077|strict|92707-9|LNC|ORDERING PHYSICIAN|ORDERING PHYSICIAN
92707-9|T077|strict|92707-9|LNC|TESTING PERFORMED BY|TESTING PERFORMED BY
92707-9|T077|strict|92707-9|LNC|PCP|PCP
92707-9|T077|strict|92707-9|LNC|OBSTETRICIAN|OBSTETRICIAN
92707-9|T077|strict|92707-9|LNC|PATHOLOGIST|PATHOLOGIST
92707-9|T077|strict|92707-9|LNC|RADIOLOGIST|RADIOLOGIST
92707-9|T077|strict|92707-9|LNC|SURGEON|SURGEON
92707-9|T077|multi|92707-9|LNC|ATTENDING|ATTENDING
92707-9|T077|multi|92707-9|LNC|ADMITTING|ADMITTING
92707-9|T077|multi|92707-9|LNC|RESIDENT|RESIDENT
92707-9|T077|multi|92707-9|LNC|SUPERVISING|SUPERVISING
44951-2|T077|strict|44951-2|LNC|PHYSICIAN NPI|PHYSICIAN NPI
44951-2|T077|strict|44951-2|LNC|NPI|NPI
44951-2|T077|strict|44951-2|LNC|PHYSICIAN DETAILS|PHYSICIAN DETAILS
44951-2|T077|strict|44951-2|LNC|NATIONAL PROVIDER IDENTIFIER|NATIONAL PROVIDER IDENTIFIER
44951-2|T077|strict|44951-2|LNC|PROVIDER INFORMATION|PROVIDER INFORMATION
44951-2|T077|strict|44951-2|LNC|PROVIDER ID|PROVIDER ID
44951-2|T077|strict|44951-2|LNC|PROVIDER NUMBER|PROVIDER NUMBER
46209-3|T077|multi|46209-3|LNC|PROVIDER ORDERS|PROVIDER ORDERS
46209-3|T077|multi|46209-3|LNC|ORDERING PROVIDER|ORDERING PROVIDER
46209-3|T077|multi|46209-3|LNC|CPOE|CPOE
46209-3|T077|multi|46209-3|LNC|COMPUTERIZED PHYSICIAN ORDER ENTRY|COMPUTERIZED PHYSICIAN ORDER ENTRY
46209-3|T077|multi|46209-3|LNC|ORDERS|ORDERS
46209-3|T077|multi|46209-3|LNC|ORDER|ORDER
46209-3|T077|multi|46209-3|LNC|ORDER DATE|ORDER DATE
46209-3|T077|multi|46209-3|LNC|ORDERED|ORDERED
46209-3|T077|multi|46209-3|LNC|ORDER DETAILS|ORDER DETAILS
46209-3|T077|multi|46209-3|LNC|ORDER STATUS|ORDER STATUS
18770-8|T077|strict|18770-8|LNC|DICTATION|DICTATION
18770-8|T077|strict|18770-8|LNC|DICTATED BY|DICTATED BY
18770-8|T077|strict|18770-8|LNC|DICTATED ON|DICTATED ON
18770-8|T077|strict|18770-8|LNC|DICTATED DATE|DICTATED DATE
18770-8|T077|strict|18770-8|LNC|DICTATED|DICTATED
18770-8|T077|strict|18770-8|LNC|TRANSCRIBED DOCUMENT PRINT|TRANSCRIBED DOCUMENT PRINT
18770-8|T077|strict|18770-8|LNC|TRANSCRIBED BY|TRANSCRIBED BY
18770-8|T077|strict|18770-8|LNC|TRANSCRIBED DATE|TRANSCRIBED DATE
18770-8|T077|strict|18770-8|LNC|TRANSCRIBED DOCUMENT|TRANSCRIBED DOCUMENT
18770-8|T077|strict|18770-8|LNC|PRINTED FROM|PRINTED FROM
18770-8|T077|strict|18770-8|LNC|PRINTED BY|PRINTED BY
18770-8|T077|strict|18770-8|LNC|PRINTED|PRINTED
18770-8|T077|strict|18770-8|LNC|PRINTED ON|PRINTED ON
18770-8|T077|strict|18770-8|LNC|DATE PRINTED|DATE PRINTED
18770-8|T077|strict|18770-8|LNC|AUTHOR|AUTHOR
18770-8|T077|strict|18770-8|LNC|AUTHORED BY|AUTHORED BY
18770-8|T077|multi|18770-8|LNC|REQUESTED BY|REQUESTED BY
18770-8|T077|strict|18770-8|LNC|GENERATED ON|GENERATED ON
18770-8|T077|strict|18770-8|LNC|GENERATED BY|GENERATED BY
18770-8|T077|strict|18770-8|LNC|LAST UPDATED|LAST UPDATED
18770-8|T077|strict|18770-8|LNC|LAST UPDATED BY|LAST UPDATED BY
18770-8|T077|strict|18770-8|LNC|MODIFIED REPORT|MODIFIED REPORT
18770-8|T077|strict|18770-8|LNC|COMPLETED BY|COMPLETED BY
18770-8|T077|strict|18770-8|LNC|ENTERED BY|ENTERED BY
18770-8|T077|strict|18770-8|LNC|SEEN BY|SEEN BY
18770-8|T077|multi|18770-8|LNC|FINAL REPORT|FINAL REPORT
18770-8|T077|strict|18770-8|LNC|END OF REPORT|END OF REPORT
76696-4|T077|multi|76696-4|LNC|FACILITY NAME|FACILITY NAME
76696-4|T077|multi|76696-4|LNC|FACILITY|FACILITY
76696-4|T077|multi|76696-4|LNC|SERVICE|SERVICE
76696-4|T077|multi|76696-4|LNC|BUILDING|BUILDING
76696-4|T077|multi|76696-4|LNC|CAMPUS|CAMPUS
76696-4|T077|multi|76696-4|LNC|DEPARTMENT|DEPARTMENT
76696-4|T077|multi|76696-4|LNC|LABCORP|LABCORP
80412-0|T077|strict|80412-0|LNC|ENCOUNTER LOCATION|ENCOUNTER LOCATION
80412-0|T077|strict|80412-0|LNC|VISIT LOCATION|VISIT LOCATION
80412-0|T077|strict|80412-0|LNC|LOCATION OF VISIT|LOCATION OF VISIT
80412-0|T077|multi|80412-0|LNC|LOCATION|LOCATION
80412-0|T077|multi|80412-0|LNC|ROOM|ROOM
18841-7|T077|multi|18841-7|LNC|HOSPITAL CONSULTATIONS|HOSPITAL CONSULTATIONS
18841-7|T077|multi|18841-7|LNC|CONSULT|CONSULT
18841-7|T077|multi|18841-7|LNC|CONSULTATION|CONSULTATION
48768-6|T077|strict|48768-6|LNC|PAYMENT SOURCES|PAYMENT SOURCES
48768-6|T077|strict|48768-6|LNC|BILLING INFORMATION|BILLING INFORMATION
48768-6|T077|strict|48768-6|LNC|INSURANCE GROUP NUMBER|INSURANCE GROUP NUMBER
48768-6|T077|strict|48768-6|LNC|INSURANCE NUMBER|INSURANCE NUMBER
48768-6|T077|strict|48768-6|LNC|MEDICARE|MEDICARE
48768-6|T077|strict|48768-6|LNC|MEDICARE PPO|MEDICARE PPO
48768-6|T077|strict|48768-6|LNC|MEDICAID|MEDICAID
48768-6|T077|strict|48768-6|LNC|GROUP #|GROUP #
48768-6|T077|multi|48768-6|LNC|INS|INS
76428-2|T077|strict|76428-2|LNC|VISIT CHARGE|VISIT CHARGE
76428-2|T077|strict|76428-2|LNC|ENCOUNTER CHARGE|ENCOUNTER CHARGE
76428-2|T077|strict|76428-2|LNC|CHARGES|CHARGES
76428-2|T077|strict|76428-2|LNC|CHARGE FOR|CHARGE FOR
75519-9|T077|strict|75519-9|LNC|ENCOUNTER IDENTIFIER|ENCOUNTER IDENTIFIER
75519-9|T077|strict|75519-9|LNC|ENCOUNTER ID|ENCOUNTER ID
75519-9|T077|strict|75519-9|LNC|ENCOUNTER NUM|ENCOUNTER NUM
75519-9|T077|strict|75519-9|LNC|ENCOUNTER #|ENCOUNTER #
75519-9|T077|strict|75519-9|LNC|ACCESSION|ACCESSION
75519-9|T077|strict|75519-9|LNC|VISIT ID|VISIT ID
75519-9|T077|strict|75519-9|LNC|CASE NUM|CASE NUM
75519-9|T077|strict|75519-9|LNC|CASE #|CASE #
75519-9|T077|strict|75519-9|LNC|CASE#|CASE#
75519-9|T077|strict|75519-9|LNC|REQUISITION|REQUISITION
57122-4|T077|strict|57122-4|LNC|TYPE OF ENCOUNTER|TYPE OF ENCOUNTER
57122-4|T077|strict|57122-4|LNC|ENCOUNTER INFORMATION|ENCOUNTER INFORMATION
57122-4|T077|strict|57122-4|LNC|ENCOUNTER INFO|ENCOUNTER INFO
57122-4|T077|strict|57122-4|LNC|ENCOUNTER|ENCOUNTER
57122-4|T077|strict|57122-4|LNC|APPOINTMENT|APPOINTMENT
57122-4|T077|strict|57122-4|LNC|APPOINTMENTS|APPOINTMENTS
57122-4|T077|strict|57122-4|LNC|APPOINTMENT INFORMATION|APPOINTMENT INFORMATION
11293-8|T077|strict|11293-8|LNC|REFERRAL SOURCE|REFERRAL SOURCE
11293-8|T077|strict|11293-8|LNC|REFERRED BY|REFERRED BY
11293-8|T077|strict|11293-8|LNC|REFERRAL|REFERRAL
11293-8|T077|strict|11293-8|LNC|REFERRING PROVIDER|REFERRING PROVIDER
11293-8|T077|strict|11293-8|LNC|ADMIT PROVIDER|ADMIT PROVIDER
39289-4|T077|strict|39289-4|LNC|FOLLOW-UP|FOLLOW-UP
39289-4|T077|strict|39289-4|LNC|FOLLOW UP|FOLLOW UP
39289-4|T077|strict|39289-4|LNC|FOLLOW UP APPOINTMENT|FOLLOW UP APPOINTMENT
39289-4|T077|strict|39289-4|LNC|FOLLOW UP APPOINTMENTS|FOLLOW UP APPOINTMENTS
85647-6|T077|strict|85647-6|LNC|SIGNATURE|SIGNATURE
85647-6|T077|strict|85647-6|LNC|SIGNATURE LINE|SIGNATURE LINE
85647-6|T077|strict|85647-6|LNC|ELECTRONICALLY SIGNED|ELECTRONICALLY SIGNED
85647-6|T077|strict|85647-6|LNC|SIGNED|SIGNED
85647-6|T077|strict|85647-6|LNC|SIGNED BY|SIGNED BY
85647-6|T077|strict|85647-6|LNC|SIGNED OFF BY|SIGNED OFF BY
85647-6|T077|strict|85647-6|LNC|SIGNED ELECTRONICALLY BY|SIGNED ELECTRONICALLY BY
85647-6|T077|strict|85647-6|LNC|SIGNATURE ON FILE|SIGNATURE ON FILE
80567-1|T077|strict|80567-1|LNC|FLOWSHEET|FLOWSHEET
80567-1|T077|strict|80567-1|LNC|FLOW SHEET|FLOW SHEET
80567-1|T077|multi|80567-1|LNC|FLOW|FLOW
89442-8|T077|multi|89442-8|LNC|OBSTETRICS ADMINISTRATIVE|OBSTETRICS ADMINISTRATIVE
89442-8|T077|multi|89442-8|LNC|PAST GYNECOLOGICAL HISTORY|PAST GYNECOLOGICAL HISTORY
89442-8|T077|multi|89442-8|LNC|NSVD|NSVD
89442-8|T077|multi|89442-8|LNC|CESAREAN STATUS|CESAREAN STATUS
89442-8|T077|multi|89442-8|LNC|DELIVERY DATE|DELIVERY DATE
89442-8|T077|multi|89442-8|LNC|MATERNAL TRANSFER|MATERNAL TRANSFER
89442-8|T077|multi|89442-8|LNC|POSTPARTUM MEASLES MUMPS RUBELLA VACCINE|POSTPARTUM MEASLES MUMPS RUBELLA VACCINE
89442-8|T077|multi|89442-8|LNC|POSTPARTUM CARE SITE|POSTPARTUM CARE SITE
89442-8|T077|multi|89442-8|LNC|PRIMARY PEDIATRIC CARE|PRIMARY PEDIATRIC CARE
89442-8|T077|multi|89442-8|LNC|PRIMARY PEDIATRICIAN|PRIMARY PEDIATRICIAN
89442-8|T077|multi|89442-8|LNC|CESAREAN STATUS|CESAREAN STATUS
89442-8|T077|multi|89442-8|LNC|BREAST FEEDING AT DISCHARGE|BREAST FEEDING AT DISCHARGE
89442-8|T077|multi|89442-8|LNC|DELIVERY|DELIVERY
89442-8|T077|multi|89442-8|LNC|PRENATAL SCREENS|PRENATAL SCREENS
89442-8|T077|multi|89442-8|LNC|EPIDURAL VAGINAL DELIVERY|EPIDURAL VAGINAL DELIVERY
89442-8|T077|multi|89442-8|LNC|UTERINE INCISION TYPE|UTERINE INCISION TYPE
89442-8|T077|multi|89442-8|LNC|NURSERY RECORDS|NURSERY RECORDS
89442-8|T077|multi|89442-8|LNC|VAGINAL DELIVERY|VAGINAL DELIVERY
79191-3|T077|strict|79191-3|LNC|PATIENT DEMOGRAPHICS|PATIENT DEMOGRAPHICS
79191-3|T077|strict|79191-3|LNC|DEMOGRAPHICS|DEMOGRAPHICS
79191-3|T077|multi|79191-3|LNC|PATIENT|PATIENT
79191-3|T077|multi|79191-3|LNC|SUBJECT|SUBJECT
79191-3|T077|multi|79191-3|LNC|PATIENT INFORMATION|PATIENT INFORMATION
79191-3|T077|multi|79191-3|LNC|PATIENT INFO|PATIENT INFO
45392-8|T077|strict|45392-8|LNC|FIRST NAME|FIRST NAME
45392-8|T077|strict|45392-8|LNC|GIVEN NAME|GIVEN NAME
45394-4|T077|strict|45394-4|LNC|LAST NAME|LAST NAME
45394-4|T077|strict|45394-4|LNC|FAMILY NAME|FAMILY NAME
87226-7|T077|strict|87226-7|LNC|PATIENT NAME|PATIENT NAME
87226-7|T077|strict|87226-7|LNC|LEGAL NAME|LEGAL NAME
87226-7|T077|strict|87226-7|LNC|FULL NAME|FULL NAME
87226-7|T077|strict|87226-7|LNC|NICK NAME|NICK NAME
87226-7|T077|strict|87226-7|LNC|SUBSCRIBER|SUBSCRIBER
87226-7|T077|strict|87226-7|LNC|SUBSCRIBER NAME|SUBSCRIBER NAME
87226-7|T077|strict|87226-7|LNC|INSURANCE SUBSCRIBER NAME|INSURANCE SUBSCRIBER NAME
72143-1|T077|strict|72143-1|LNC|ADMINISTRATIVE GENDER|ADMINISTRATIVE GENDER
72143-1|T077|strict|72143-1|LNC|PATIENT GENDER|PATIENT GENDER
72143-1|T077|strict|72143-1|LNC|GENDER|GENDER
72143-1|T077|strict|72143-1|LNC|PATIENT SEX|PATIENT SEX
72143-1|T077|multi|72143-1|LNC|SEX|SEX
21112-8|T077|strict|21112-8|LNC|BIRTH DATE|BIRTH DATE
21112-8|T077|strict|21112-8|LNC|DATE OF BIRTH|DATE OF BIRTH
21112-8|T077|strict|21112-8|LNC|DOB|DOB
21112-8|T077|strict|21112-8|LNC|PATIENT DATE OF BIRTH|PATIENT DATE OF BIRTH
21112-8|T077|strict|21112-8|LNC|SUBSCRIBER DATE OF BIRTH|SUBSCRIBER DATE OF BIRTH
81954-0|T077|strict|81954-0|LNC|DATE OF DEATH|DATE OF DEATH
81954-0|T077|multi|81954-0|LNC|DEATH|DEATH
21612-7|T077|strict|21612-7|LNC|PATIENT AGE|PATIENT AGE
21612-7|T077|strict|21612-7|LNC|AGE|AGE
80977-2|T077|strict|80977-2|LNC|PATIENT RACE|PATIENT RACE
80977-2|T077|multi|80977-2|LNC|RACE|RACE
80977-2|T077|strict|80977-2|LNC|TABULATED RACE|TABULATED RACE
80977-2|T077|strict|80977-2|LNC|CDC RACE|CDC RACE
80978-0|T077|strict|80978-0|LNC|PATIENT ETHNICITY|PATIENT ETHNICITY
80978-0|T077|strict|80978-0|LNC|ETHNICITY|ETHNICITY
80978-0|T077|strict|80978-0|LNC|CDC ETHNICITY|CDC ETHNICITY
80978-0|T077|strict|80978-0|LNC|TABULATED ETHNICITY|TABULATED ETHNICITY
54899-0|T077|strict|54899-0|LNC|PREFERRED LANGUAGE|PREFERRED LANGUAGE
54899-0|T077|strict|54899-0|LNC|PREF LANGUAGE|PREF LANGUAGE
54899-0|T077|strict|54899-0|LNC|PATIENT LANGUAGE|PATIENT LANGUAGE
54899-0|T077|strict|54899-0|LNC|LANGUAGE|LANGUAGE
42078-6|T077|strict|42078-6|LNC|FOLLOW-UP CONTACT|FOLLOW-UP CONTACT
42078-6|T077|strict|42078-6|LNC|EMERGENCY CONTACT|EMERGENCY CONTACT
42078-6|T077|multi|42078-6|LNC|CONTACT|CONTACT
42078-6|T077|strict|42078-6|LNC|CONTACT BY|CONTACT BY
76458-9|T077|strict|76458-9|LNC|PATIENT EMAIL ADDRESS|PATIENT EMAIL ADDRESS
76458-9|T077|strict|76458-9|LNC|EMAIL ADDRESS|EMAIL ADDRESS
76458-9|T077|strict|76458-9|LNC|TRUSTED EMAIL|TRUSTED EMAIL
76458-9|T077|multi|76458-9|LNC|EMAIL|EMAIL
76458-9|T077|multi|76458-9|LNC|E-MAIL|E-MAIL
92634-5|T077|multi|92634-5|LNC|ADDRESS TYPE|ADDRESS TYPE
92634-5|T077|multi|92634-5|LNC|CITY/ST|CITY/ST
92634-5|T077|multi|92634-5|LNC|CITY,ST|CITY,ST
92634-5|T077|multi|92634-5|LNC|CITY|CITY
92634-5|T077|multi|92634-5|LNC|STATE|STATE
56799-0|T077|strict|56799-0|LNC|PATIENT ADDRESS|PATIENT ADDRESS
56799-0|T077|strict|56799-0|LNC|HOME ADDRESS|HOME ADDRESS
56799-0|T077|multi|56799-0|LNC|ADDRESS|ADDRESS
56799-0|T077|strict|56799-0|LNC|WORK ADDRESS|WORK ADDRESS
56799-0|T077|strict|56799-0|LNC|ADDRESS LINE 1|ADDRESS LINE 1
56799-0|T077|strict|56799-0|LNC|ADDRESS LINE 2|ADDRESS LINE 2
56799-0|T077|strict|56799-0|LNC|STREET ADDRESS|STREET ADDRESS
56799-0|T077|multi|56799-0|LNC|STREET|STREET
42077-8|T077|strict|42077-8|LNC|PATIENT PHONE NUMBER|PATIENT PHONE NUMBER
42077-8|T077|strict|42077-8|LNC|CELL PHONE|CELL PHONE
42077-8|T077|strict|42077-8|LNC|HOME PHONE|HOME PHONE
42077-8|T077|multi|42077-8|LNC|PHONE NUMBER|PHONE NUMBER
42077-8|T077|strict|42077-8|LNC|PHONE|PHONE
42077-8|T077|strict|42077-8|LNC|WORK PHONE|WORK PHONE
42077-8|T077|strict|42077-8|LNC|PHONE EXTENSION|PHONE EXTENSION
42077-8|T077|strict|42077-8|LNC|WORK PHONE EXTENSION|WORK PHONE EXTENSION
42077-8|T077|multi|42077-8|LNC|EXTENSION|EXTENSION
42077-8|T077|strict|42077-8|LNC|MOBILE PHONE|MOBILE PHONE
42077-8|T077|strict|42077-8|LNC|MOBILE|MOBILE
68997-6|T077|strict|68997-6|LNC|PATIENT CITY|PATIENT CITY
68997-6|T077|multi|68997-6|LNC|CITY|CITY
46499-0|T077|strict|46499-0|LNC|PATIENT STATE|PATIENT STATE
46499-0|T077|strict|46499-0|LNC|PATIENT HOME STATE|PATIENT HOME STATE
46499-0|T077|strict|46499-0|LNC|STATE OF RESIDENCE|STATE OF RESIDENCE
46499-0|T077|multi|46499-0|LNC|STATE|STATE
45401-7|T077|strict|45401-7|LNC|POSTAL CODE|POSTAL CODE
45401-7|T077|strict|45401-7|LNC|PATIENT ZIP|PATIENT ZIP
45401-7|T077|strict|45401-7|LNC|ZIP CODE|ZIP CODE
45401-7|T077|multi|45401-7|LNC|ZIP|ZIP
45401-7|T077|strict|45401-7|LNC|POSTAL|POSTAL
87721-7|T077|strict|87721-7|LNC|COUNTY OF RESIDENCE|COUNTY OF RESIDENCE
87721-7|T077|multi|87721-7|LNC|COUNTY|COUNTY
66477-1|T077|strict|66477-1|LNC|COUNTRY OF CURRENT RESIDENCE|COUNTRY OF CURRENT RESIDENCE
66477-1|T077|multi|66477-1|LNC|COUNTRY|COUNTRY
81365-9|T077|strict|81365-9|LNC|RELIGIOUS AFFILIATION|RELIGIOUS AFFILIATION
81365-9|T077|strict|81365-9|LNC|PATIENT RELIGION|PATIENT RELIGION
81365-9|T077|strict|81365-9|LNC|RELIGION|RELIGION
85658-3|T077|strict|85658-3|LNC|PROFESSION|PROFESSION
85658-3|T077|strict|85658-3|LNC|OCCUPATION|OCCUPATION
85658-3|T077|strict|85658-3|LNC|OCCUPATION TYPE|OCCUPATION TYPE
85658-3|T077|strict|85658-3|LNC|EMPLOYER NAME|EMPLOYER NAME
85658-3|T077|strict|85658-3|LNC|EMPLOYER ADDRESS|EMPLOYER ADDRESS
85658-3|T077|strict|85658-3|LNC|JOB|JOB
46106-1|T077|strict|46106-1|LNC|MEDICAL RECORD NUMBER|MEDICAL RECORD NUMBER
46106-1|T077|strict|46106-1|LNC|MEDICAL RECORD #|MEDICAL RECORD #
46106-1|T077|strict|46106-1|LNC|CHART NUMBER|CHART NUMBER
46106-1|T077|strict|46106-1|LNC|MRN|MRN
45396-9|T077|strict|45396-9|LNC|SSN|SSN
45396-9|T077|strict|45396-9|LNC|SOCIAL SECURITY NUMBER|SOCIAL SECURITY NUMBER
45396-9|T077|strict|45396-9|LNC|INSURANCE SUBSCRIBER SSN|INSURANCE SUBSCRIBER SSN
45396-9|T077|strict|45396-9|LNC|SOCIAL SECURITY NO|SOCIAL SECURITY NO
45396-9|T077|strict|45396-9|LNC|SOCIAL SECURITY NUM|SOCIAL SECURITY NUM
45396-9|T077|strict|45396-9|LNC|SOCIAL SEC NO|SOCIAL SEC NO
45396-9|T077|strict|45396-9|LNC|SOC SEC NO|SOC SEC NO
45396-9|T077|strict|45396-9|LNC|SOC. SEC. NO|SOC. SEC. NO
45396-9|T077|strict|45396-9|LNC|SOCIAL SECURITY #|SOCIAL SECURITY #
76435-7|T077|strict|76435-7|LNC|PATIENT ID|PATIENT ID
76435-7|T077|strict|76435-7|LNC|PATIENT IDENTIFIER|PATIENT IDENTIFIER
76435-7|T077|multi|76435-7|LNC|ACC|ACC
76435-7|T077|strict|76435-7|LNC|ACCOUNT|ACCOUNT
76435-7|T077|strict|76435-7|LNC|PATIENT NUMBER|PATIENT NUMBER
76435-7|T077|strict|76435-7|LNC|IDENTIFICATION DATA|IDENTIFICATION DATA
76435-7|T077|strict|76435-7|LNC|IDENTIFYING DATA|IDENTIFYING DATA
76435-7|T077|multi|76435-7|LNC|IDENTIFICATION|IDENTIFICATION
76435-7|T077|strict|76435-7|LNC|INSURANCE ID NUMBER|INSURANCE ID NUMBER
76435-7|T077|strict|76435-7|LNC|EXTERNAL ID|EXTERNAL ID
76437-3|T077|strict|76437-3|LNC|PRIMARY INSURANCE DATA|PRIMARY INSURANCE DATA
76437-3|T077|strict|76437-3|LNC|PRIMARY INSURANCE|PRIMARY INSURANCE
76437-3|T077|strict|76437-3|LNC|ACTIVE PRIMARY INSURANCE|ACTIVE PRIMARY INSURANCE
76437-3|T077|strict|76437-3|LNC|PAYOR SOURCE|PAYOR SOURCE
76437-3|T077|strict|76437-3|LNC|PAYERS|PAYERS
76437-3|T077|strict|76437-3|LNC|PAYORS|PAYORS
76437-3|T077|strict|76437-3|LNC|INSURANCE|INSURANCE
76437-3|T077|strict|76437-3|LNC|SECONDARY INSURANCE|SECONDARY INSURANCE
76437-3|T077|strict|76437-3|LNC|INSURANCE COMPANY|INSURANCE COMPANY
76437-3|T077|strict|76437-3|LNC|INSURANCE DATA|INSURANCE DATA
76437-3|T077|strict|76437-3|LNC|INSURANCE PROVIDERS|INSURANCE PROVIDERS
76437-3|T077|strict|76437-3|LNC|HEALTH INSURANCE|HEALTH INSURANCE
76437-3|T077|strict|76437-3|LNC|BENEFITS ASSIGNED|BENEFITS ASSIGNED
76437-3|T077|strict|76437-3|LNC|INSURANCE|INSURANCE
11366-2|T077|strict|11366-2|LNC|SMOKING STATUS|SMOKING STATUS
11366-2|T077|strict|11366-2|LNC|HISTORY OF TOBACCO USE|HISTORY OF TOBACCO USE
11366-2|T077|strict|11366-2|LNC|TOBACCO USE STATUS|TOBACCO USE STATUS
11366-2|T077|strict|11366-2|LNC|SMOKING HISTORY|SMOKING HISTORY
11366-2|T077|strict|11366-2|LNC|SMOKING EXPOSURE|SMOKING EXPOSURE
11366-2|T077|strict|11366-2|LNC|SMOKING EXPOSURE|SMOKING EXPOSURE
11366-2|T077|strict|11366-2|LNC|TOBACCO USE|TOBACCO USE
11366-2|T077|strict|11366-2|LNC|SMOKING|SMOKING
11366-2|T077|strict|11366-2|LNC|TOBACCO|TOBACCO
11366-2|T077|multi|11366-2|LNC|DATE QUIT|DATE QUIT
11366-2|T077|multi|11366-2|LNC|QUIT DATE|QUIT DATE
29762-2|T077|strict|29762-2|LNC|SOCIAL HISTORY|SOCIAL HISTORY
29762-2|T077|strict|29762-2|LNC|SOCIAL HX|SOCIAL HX
29762-2|T077|strict|29762-2|LNC|POVERTY STATUS|POVERTY STATUS
29762-2|T077|multi|29762-2|LNC|DRINKING|DRINKING
29762-2|T077|strict|29762-2|LNC|PHYSICAL EXERCISE|PHYSICAL EXERCISE
29762-2|T077|multi|29762-2|LNC|EXERCISE|EXERCISE
29762-2|T077|multi|29762-2|LNC|SOCIAL|SOCIAL
29762-2|T077|strict|29762-2|LNC|HABITS|HABITS
29762-2|T077|strict|29762-2|LNC|POVERTY|POVERTY
29762-2|T077|strict|29762-2|LNC|HOMELESS|HOMELESS
29762-2|T077|strict|29762-2|LNC|SHX|SHX
29762-2|T077|strict|29762-2|LNC|PSH|PSH
47420-5|T077|strict|47420-5|LNC|FUNCTIONAL STATUS ASSESSMENT NOTE|FUNCTIONAL STATUS ASSESSMENT NOTE
47420-5|T077|strict|47420-5|LNC|FUNCTIONAL STATUS ASSESSMENT|FUNCTIONAL STATUS ASSESSMENT
47420-5|T077|strict|47420-5|LNC|FUNCTIONAL STATUS|FUNCTIONAL STATUS
47420-5|T077|strict|47420-5|LNC|FUNCTIONAL ABILITIES|FUNCTIONAL ABILITIES
47420-5|T077|strict|47420-5|LNC|CURRENT HEALTH STATUS|CURRENT HEALTH STATUS
47420-5|T077|strict|47420-5|LNC|PREVENTIVE|PREVENTIVE
47420-5|T077|multi|47420-5|LNC|IMPAIRMENTS|IMPAIRMENTS
47420-5|T077|strict|47420-5|LNC|DISCHARGE CONDITION|DISCHARGE CONDITION
47420-5|T077|strict|47420-5|LNC|DISCHARGED CONDITION ON DISCHARGE|DISCHARGED CONDITION ON DISCHARGE
47420-5|T077|strict|47420-5|LNC|DISCHARGE STATUS|DISCHARGE STATUS
47420-5|T077|strict|47420-5|LNC|CONDITION ON DISCHARGE|CONDITION ON DISCHARGE
47420-5|T077|strict|47420-5|LNC|CONDITION ON TRANSFER|CONDITION ON TRANSFER
10160-0|T077|strict|10160-0|LNC|MEDICATION LIST|MEDICATION LIST
10160-0|T077|strict|10160-0|LNC|FINAL MEDICATIONS|FINAL MEDICATIONS
10160-0|T077|strict|10160-0|LNC|HISTORY OF MEDICATION USE|HISTORY OF MEDICATION USE
10160-0|T077|strict|10160-0|LNC|LIST MEDICATIONS|LIST MEDICATIONS
10160-0|T077|strict|10160-0|LNC|CONDITION MEDICATIONS|CONDITION MEDICATIONS
10160-0|T077|strict|10160-0|LNC|CURRENT MEDICATIONS|CURRENT MEDICATIONS
10160-0|T077|strict|10160-0|LNC|AS NEEDED MEDICATIONS|AS NEEDED MEDICATIONS
10160-0|T077|strict|10160-0|LNC|THE FOLLOWING MEDICATIONS|THE FOLLOWING MEDICATIONS
10160-0|T077|strict|10160-0|LNC|FOLLOWING MEDICATIONS|FOLLOWING MEDICATIONS
10160-0|T077|strict|10160-0|LNC|FOLLOWING MEDICATIONS|FOLLOWING MEDICATIONS
10160-0|T077|strict|10160-0|LNC|DRUG HISTORY|DRUG HISTORY
10160-0|T077|strict|10160-0|LNC|HOME MEDICATIONS|HOME MEDICATIONS
10160-0|T077|strict|10160-0|LNC|MEDICATIONS AT HOME|MEDICATIONS AT HOME
10160-0|T077|strict|10160-0|LNC|INHOSPITAL MEDICATIONS|INHOSPITAL MEDICATIONS
10160-0|T077|strict|10160-0|LNC|MOST RECENT MEDICATIONS|MOST RECENT MEDICATIONS
10160-0|T077|strict|10160-0|LNC|NEW MEDICATIONS|NEW MEDICATIONS
10160-0|T077|strict|10160-0|LNC|MEDICATION CHANGES|MEDICATION CHANGES
10160-0|T077|strict|10160-0|LNC|MEDICATIONS AT REHAB|MEDICATIONS AT REHAB
10160-0|T077|strict|10160-0|LNC|MEDICATIONS AT REHABILITATION|MEDICATIONS AT REHABILITATION
10160-0|T077|strict|10160-0|LNC|MEDICATIONS ON PRESENTATION|MEDICATIONS ON PRESENTATION
10160-0|T077|strict|10160-0|LNC|OUTPATIENT MEDICATIONS|OUTPATIENT MEDICATIONS
10160-0|T077|strict|10160-0|LNC|NUMBER OF DOSES REQUIRED APPROXIMATE|NUMBER OF DOSES REQUIRED APPROXIMATE
10160-0|T077|strict|10160-0|LNC|MEDS AT HOME|MEDS AT HOME
10160-0|T077|strict|10160-0|LNC|MEDS|MEDS
10160-0|T077|strict|10160-0|LNC|PRESCRIPTIONS|PRESCRIPTIONS
10160-0|T077|strict|10160-0|LNC|PRN MEDICATIONS|PRN MEDICATIONS
10160-0|T077|strict|10160-0|LNC|MEDICATIONS|MEDICATIONS
10160-0|T077|strict|10160-0|LNC|MEDICATION|MEDICATION
42346-7|T077|strict|42346-7|LNC|MEDICATIONS ON ADMISSION|MEDICATIONS ON ADMISSION
42346-7|T077|strict|42346-7|LNC|ADMISSION MEDICATIONS|ADMISSION MEDICATIONS
42346-7|T077|strict|42346-7|LNC|MEDICATIONS AT ADMISSION|MEDICATIONS AT ADMISSION
42346-7|T077|strict|42346-7|LNC|MEDICATIONS UPON ADMISSION|MEDICATIONS UPON ADMISSION
42346-7|T077|strict|42346-7|LNC|MEDICATIONS AT THE TIME OF ADMISSION|MEDICATIONS AT THE TIME OF ADMISSION
42346-7|T077|strict|42346-7|LNC|MEDICATIONS AT TIME OF ADMISSION|MEDICATIONS AT TIME OF ADMISSION
42346-7|T077|strict|42346-7|LNC|MEDICATION CHANGES MADE DURING THIS ADMISSION|MEDICATION CHANGES MADE DURING THIS ADMISSION
42346-7|T077|strict|42346-7|LNC|RX ON ADMIT|RX ON ADMIT
42346-7|T077|strict|42346-7|LNC|MEDICATIONS PRIOR TO ADMISSION|MEDICATIONS PRIOR TO ADMISSION
42346-7|T077|strict|42346-7|LNC|PREADMISSION MEDICATIONS|PREADMISSION MEDICATIONS
42346-7|T077|strict|42346-7|LNC|PREOP MEDICATIONS|PREOP MEDICATIONS
42346-7|T077|strict|42346-7|LNC|PREOPERATIVE MEDICATIONS|PREOPERATIVE MEDICATIONS
42346-7|T077|strict|42346-7|LNC|HOME MEDICATIONS ON ADMISSION|HOME MEDICATIONS ON ADMISSION
42346-7|T077|strict|42346-7|LNC|BLOCK MEDICATIONS ON ADMISSION|BLOCK MEDICATIONS ON ADMISSION
29549-3|T077|multi|29549-3|LNC|MEDICATION ADMINISTERED|MEDICATION ADMINISTERED
29549-3|T077|strict|29549-3|LNC|MEDICATION ADMINISTERED|MEDICATION ADMINISTERED
29549-3|T077|strict|29549-3|LNC|FLUIDS RECEIVED|FLUIDS RECEIVED
29549-3|T077|strict|29549-3|LNC|IV FLUIDS|IV FLUIDS
29549-3|T077|strict|29549-3|LNC|FLUIDS|FLUIDS
10183-2|T077|strict|10183-2|LNC|HOSPITAL DISCHARGE MEDICATIONS|HOSPITAL DISCHARGE MEDICATIONS
10183-2|T077|strict|10183-2|LNC|DISCHARGE MEDICATIONS|DISCHARGE MEDICATIONS
10183-2|T077|strict|10183-2|LNC|DISCHARGE MEDICATIONS INCLUDE|DISCHARGE MEDICATIONS INCLUDE
10183-2|T077|strict|10183-2|LNC|DISCHARGE MEDICATION|DISCHARGE MEDICATION
10183-2|T077|strict|10183-2|LNC|DISCHARGED TO HOME ON THE FOLLOWING MEDICATIONS|DISCHARGED TO HOME ON THE FOLLOWING MEDICATIONS
10183-2|T077|strict|10183-2|LNC|ADDENDUM TO MEDICATIONS ON DISCHARGE|ADDENDUM TO MEDICATIONS ON DISCHARGE
10183-2|T077|strict|10183-2|LNC|REHABILITATION HOSPITAL DISCHARGE MEDICATIONS|REHABILITATION HOSPITAL DISCHARGE MEDICATIONS
10183-2|T077|strict|10183-2|LNC|MEDICATIONS UPON DISCHARGE|MEDICATIONS UPON DISCHARGE
10183-2|T077|strict|10183-2|LNC|MEDICATION AT THE TIME OF DISCHARGE|MEDICATION AT THE TIME OF DISCHARGE
10183-2|T077|strict|10183-2|LNC|MEDICATION AT TIME OF DISCHARGE|MEDICATION AT TIME OF DISCHARGE
10183-2|T077|strict|10183-2|LNC|MEDICATIONS AT THAT TIME OF DISCHARGE|MEDICATIONS AT THAT TIME OF DISCHARGE
10183-2|T077|strict|10183-2|LNC|MEDICATIONS AT THE TIME OF DISCHARGE|MEDICATIONS AT THE TIME OF DISCHARGE
10183-2|T077|strict|10183-2|LNC|MEDICATIONS AT TIME OF DISCHARGE|MEDICATIONS AT TIME OF DISCHARGE
10183-2|T077|strict|10183-2|LNC|MEDICATIONS ON DISCHARGE|MEDICATIONS ON DISCHARGE
10183-2|T077|strict|10183-2|LNC|MEDICATION ON DISCHARGE|MEDICATION ON DISCHARGE
10183-2|T077|strict|10183-2|LNC|MEDICATIONS AT DISCHARGE|MEDICATIONS AT DISCHARGE
10183-2|T077|strict|10183-2|LNC|MEDICATIONS UPON TRANSFER|MEDICATIONS UPON TRANSFER
10183-2|T077|strict|10183-2|LNC|MEDICATIONS ON TRANSFER|MEDICATIONS ON TRANSFER
10183-2|T077|strict|10183-2|LNC|TRANSFER MEDICATIONS|TRANSFER MEDICATIONS
10183-2|T077|strict|10183-2|LNC|MEDICATIONS AT THE TIME OF TRANSFER|MEDICATIONS AT THE TIME OF TRANSFER
10183-2|T077|strict|10183-2|LNC|MEDICATIONS AT THE TIME OF TRANSFER TO THE CCU|MEDICATIONS AT THE TIME OF TRANSFER TO THE CCU
10183-2|T077|strict|10183-2|LNC|MEDICATIONS AT THE TIME OF TRANSFER TO THE ICU|MEDICATIONS AT THE TIME OF TRANSFER TO THE ICU
10183-2|T077|strict|10183-2|LNC|MEDS ON TRANSFER|MEDS ON TRANSFER
45841-4|T077|strict|45841-4|LNC|CHEMOTHERAPY|CHEMOTHERAPY
45841-4|T077|strict|45841-4|LNC|CHEMO|CHEMO
45851-3|T077|strict|45851-3|LNC|TRANSFUSIONS|TRANSFUSIONS
45843-0|T077|strict|45843-0|LNC|IV MEDICATION|IV MEDICATION
45843-0|T077|strict|45843-0|LNC|IV MEDICATIONS|IV MEDICATIONS
45843-0|T077|strict|45843-0|LNC|IV|IV
48765-2|T077|strict|48765-2|LNC|ALLERGY LIST|ALLERGY LIST
48765-2|T077|strict|48765-2|LNC|ALLERGIES, ADVERSE REACTIONS, ALERTS|ALLERGIES, ADVERSE REACTIONS, ALERTS
48765-2|T077|strict|48765-2|LNC|ALLERGIES & ADVERSE REACTIONS|ALLERGIES & ADVERSE REACTIONS
48765-2|T077|strict|48765-2|LNC|ALLERGIES AND ADVERSE REACTIONS|ALLERGIES AND ADVERSE REACTIONS
48765-2|T077|strict|48765-2|LNC|ADVERSE DRUG REACTIONS|ADVERSE DRUG REACTIONS
48765-2|T077|strict|48765-2|LNC|ADVERSE REACTIONS|ADVERSE REACTIONS
48765-2|T077|strict|48765-2|LNC|DRUG ALLERGIES|DRUG ALLERGIES
48765-2|T077|strict|48765-2|LNC|POTENTIALLY SERIOUS INTERACTION|POTENTIALLY SERIOUS INTERACTION
48765-2|T077|strict|48765-2|LNC|SERIOUS INTERACTION|SERIOUS INTERACTION
48765-2|T077|strict|48765-2|LNC|ALLERGIES LIST|ALLERGIES LIST
48765-2|T077|multi|48765-2|LNC|ALERTS|ALERTS
48765-2|T077|strict|48765-2|LNC|MEDICATION ALLERGIES|MEDICATION ALLERGIES
48765-2|T077|strict|48765-2|LNC|MEDICATION ALLERGY|MEDICATION ALLERGY
48765-2|T077|strict|48765-2|LNC|ALLERGIES|ALLERGIES
48765-2|T077|strict|48765-2|LNC|ALLERGY|ALLERGY
48765-2|T077|multi|48765-2|LNC|REACTIONS|REACTIONS
48765-2|T077|multi|48765-2|LNC|REACTION|REACTION
48765-2|T077|strict|48765-2|LNC|ENVIRONMENTAL ALLERGIES|ENVIRONMENTAL ALLERGIES
48765-2|T077|strict|48765-2|LNC|FOOD ALLERGIES|FOOD ALLERGIES
48765-2|T077|strict|48765-2|LNC|NO KNOWN ALLERGIES|NO KNOWN ALLERGIES
48765-2|T077|strict|48765-2|LNC|NO KNOWN DRUG ALLERGIES|NO KNOWN DRUG ALLERGIES
48765-2|T077|strict|48765-2|LNC|NKA|NKA
48765-2|T077|strict|48765-2|LNC|N.K.A.|N.K.A.
48765-2|T077|strict|48765-2|LNC|NKDA|NKDA
48765-2|T077|strict|48765-2|LNC|N.K.D.A.|N.K.D.A.
11369-6|T077|multi|11369-6|LNC|HISTORY OF IMMUNIZATION|HISTORY OF IMMUNIZATION
11369-6|T077|strict|11369-6|LNC|HISTORY OF IMMUNIZATIONS|HISTORY OF IMMUNIZATIONS
11369-6|T077|strict|11369-6|LNC|IMMUNIZATION HISTORY|IMMUNIZATION HISTORY
11369-6|T077|strict|11369-6|LNC|IMMUNIZATIONS AND VACCINES|IMMUNIZATIONS AND VACCINES
11369-6|T077|strict|11369-6|LNC|LIST OF VACCINES|LIST OF VACCINES
11369-6|T077|strict|11369-6|LNC|VACCINES LIST|VACCINES LIST
11369-6|T077|strict|11369-6|LNC|IMMUNIZATIONS LIST|IMMUNIZATIONS LIST
11369-6|T077|strict|11369-6|LNC|IMMUNIZATIONS PROVIDED|IMMUNIZATIONS PROVIDED
11369-6|T077|strict|11369-6|LNC|IMMUNIZATION|IMMUNIZATION
11369-6|T077|strict|11369-6|LNC|IMMUNIZATIONS|IMMUNIZATIONS
11369-6|T077|strict|11369-6|LNC|VACCINE|VACCINE
11369-6|T077|strict|11369-6|LNC|VACCINES|VACCINES
11369-6|T077|strict|11369-6|LNC|IMMUNIZATIONS RECOMMENDED|IMMUNIZATIONS RECOMMENDED
8716-3|T077|strict|8716-3|LNC|VITAL SIGNS|VITAL SIGNS
8716-3|T077|strict|8716-3|LNC|VITAL SIGNS PANEL|VITAL SIGNS PANEL
8716-3|T077|strict|8716-3|LNC|VITALS ON ADMISSION|VITALS ON ADMISSION
8716-3|T077|strict|8716-3|LNC|VS/MEASUREMENTS|VS/MEASUREMENTS
8716-3|T077|strict|8716-3|LNC|FILED VITALS|FILED VITALS
8716-3|T077|strict|8716-3|LNC|VS|VS
8716-3|T077|multi|8716-3|LNC|VITALS|VITALS
8716-3|T077|multi|8716-3|LNC|PULSE|PULSE
8716-3|T077|strict|8716-3|LNC|BODY TEMPERATURE|BODY TEMPERATURE
8716-3|T077|strict|8716-3|LNC|TEMPERATURE CHART|TEMPERATURE CHART
8716-3|T077|strict|8716-3|LNC|TEMPERATURE CHARTS|TEMPERATURE CHARTS
8716-3|T077|multi|8716-3|LNC|TEMPERATURE|TEMPERATURE
8716-3|T077|multi|8716-3|LNC|TEMP|TEMP
8716-3|T077|multi|8716-3|LNC|HEART RATE|HEART RATE
8716-3|T077|multi|8716-3|LNC|RESPIRATORY RATE|RESPIRATORY RATE
8716-3|T077|multi|8716-3|LNC|BLOOD PRESSURE|BLOOD PRESSURE
8716-3|T077|multi|8716-3|LNC|RATE|RATE
30954-2|T077|strict|30954-2|LNC|RELEVANT DIAGNOSTIC TESTS/LABORATORY DATA|RELEVANT DIAGNOSTIC TESTS/LABORATORY DATA
30954-2|T077|strict|30954-2|LNC|RELEVANT DIAGNOSTIC TESTS LABORATORY DATA|RELEVANT DIAGNOSTIC TESTS LABORATORY DATA
30954-2|T077|strict|30954-2|LNC|RELEVANT DIAGNOSTIC TESTS OR LABORATORY DATA|RELEVANT DIAGNOSTIC TESTS OR LABORATORY DATA
30954-2|T077|strict|30954-2|LNC|NOTABLE LABS|NOTABLE LABS
30954-2|T077|strict|30954-2|LNC|PERTINENT LAB VALUES|PERTINENT LAB VALUES
30954-2|T077|strict|30954-2|LNC|PERTINENT LABORATORY RESULTS|PERTINENT LABORATORY RESULTS
30954-2|T077|strict|30954-2|LNC|PERTINENT LABORATORY TESTS AND RESULTS|PERTINENT LABORATORY TESTS AND RESULTS
30954-2|T077|strict|30954-2|LNC|PERTINENT LABORATORY TESTS AND STUDIES|PERTINENT LABORATORY TESTS AND STUDIES
30954-2|T077|strict|30954-2|LNC|PERTINENT LABS UPON PRESENTATION|PERTINENT LABS UPON PRESENTATION
30954-2|T077|strict|30954-2|LNC|PERTINENT LABS|PERTINENT LABS
30954-2|T077|strict|30954-2|LNC|RELEVANT LABS|RELEVANT LABS
30954-2|T077|strict|30954-2|LNC|NOTABLE LABORATORY VALUES ON ADMISSION|NOTABLE LABORATORY VALUES ON ADMISSION
30954-2|T077|strict|30954-2|LNC|PERTINENT LABORATORY DATA ON ADMISSION|PERTINENT LABORATORY DATA ON ADMISSION
30954-2|T077|strict|30954-2|LNC|PERTINENT LABS ON ADMISSION|PERTINENT LABS ON ADMISSION
30954-2|T077|strict|30954-2|LNC|RELEVANT ADMISSION LABS|RELEVANT ADMISSION LABS
30954-2|T077|strict|30954-2|LNC|SIGNIFICANT LABS ON ADMISSION|SIGNIFICANT LABS ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORIES OF NOTE|LABORATORIES OF NOTE
30954-2|T077|strict|30954-2|LNC|ADMISSION LAB|ADMISSION LAB
30954-2|T077|strict|30954-2|LNC|ADMISSION LABS|ADMISSION LABS
30954-2|T077|strict|30954-2|LNC|ADMISSION LABS AND STUDIES|ADMISSION LABS AND STUDIES
30954-2|T077|strict|30954-2|LNC|ADMISSION LABORATORY|ADMISSION LABORATORY
30954-2|T077|strict|30954-2|LNC|ADMISSION LABORATORIES|ADMISSION LABORATORIES
30954-2|T077|strict|30954-2|LNC|ADMISSION LABORATORY DATA|ADMISSION LABORATORY DATA
30954-2|T077|strict|30954-2|LNC|ADMISSION LABORATORY STUDIES|ADMISSION LABORATORY STUDIES
30954-2|T077|strict|30954-2|LNC|ADMISSION LABORATORY RESULTS|ADMISSION LABORATORY RESULTS
30954-2|T077|strict|30954-2|LNC|ADMISSION LABORATORY VALUES|ADMISSION LABORATORY VALUES
30954-2|T077|strict|30954-2|LNC|ADMISSIONS LABORATORIES|ADMISSIONS LABORATORIES
30954-2|T077|strict|30954-2|LNC|ADMITTING LABORATORY|ADMITTING LABORATORY
30954-2|T077|multi|30954-2|LNC|LABORATORY FINDINGS ON ADMISSION|LABORATORY FINDINGS ON ADMISSION
30954-2|T077|strict|30954-2|LNC|PREOPERATIVE LAB|PREOPERATIVE LAB
30954-2|T077|strict|30954-2|LNC|PREOPERATIVE LABS|PREOPERATIVE LABS
30954-2|T077|strict|30954-2|LNC|PREOPERATIVE LABORATORY DATA|PREOPERATIVE LABORATORY DATA
30954-2|T077|strict|30954-2|LNC|PREOPERATIVE LABORATORY RESULTS|PREOPERATIVE LABORATORY RESULTS
30954-2|T077|strict|30954-2|LNC|PREOPERATIVE LABORATORY VALUES|PREOPERATIVE LABORATORY VALUES
30954-2|T077|strict|30954-2|LNC|PREOP LABS|PREOP LABS
30954-2|T077|strict|30954-2|LNC|ADMIT LABS|ADMIT LABS
30954-2|T077|strict|30954-2|LNC|LAB STUDIES ON ADMISSION|LAB STUDIES ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORIES ON ADMISSION|LABORATORIES ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORY DATA AT ADMISSION|LABORATORY DATA AT ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORY DATA ON ADMISSION|LABORATORY DATA ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORY DATA UPON ADMISSION|LABORATORY DATA UPON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORY EXAM ON ADMISSION|LABORATORY EXAM ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORY EXAMS UPON ADMISSION|LABORATORY EXAMS UPON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORY ON ADMISSION|LABORATORY ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORY STUDIES ON ADMISSION|LABORATORY STUDIES ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORY STUDIES UPON ADMISSION|LABORATORY STUDIES UPON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABORATORY VALUES ON ADMISSION|LABORATORY VALUES ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABS AND STUDIES ON ADMISSION|LABS AND STUDIES ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABS AT ADMISSION|LABS AT ADMISSION
30954-2|T077|strict|30954-2|LNC|LABS ON ADMISSION|LABS ON ADMISSION
30954-2|T077|strict|30954-2|LNC|LABS ON ADMIT|LABS ON ADMIT
30954-2|T077|strict|30954-2|LNC|LABS UPON ADMISSION|LABS UPON ADMISSION
30954-2|T077|multi|30954-2|LNC|RESULTS DIAGNOSTIC FINDINGS|RESULTS DIAGNOSTIC FINDINGS
30954-2|T077|strict|30954-2|LNC|INITIAL LABORATORY DATA|INITIAL LABORATORY DATA
30954-2|T077|strict|30954-2|LNC|INITIAL LABORATORY STUDIES|INITIAL LABORATORY STUDIES
30954-2|T077|strict|30954-2|LNC|LABORATORY DATA|LABORATORY DATA
30954-2|T077|strict|30954-2|LNC|LAB RESULTS|LAB RESULTS
30954-2|T077|strict|30954-2|LNC|LABORATORY EXAM|LABORATORY EXAM
30954-2|T077|strict|30954-2|LNC|LABORATORY EXAMS|LABORATORY EXAMS
30954-2|T077|strict|30954-2|LNC|LABORATORY EVALUATION|LABORATORY EVALUATION
30954-2|T077|strict|30954-2|LNC|LABORATORY EXAMINATION|LABORATORY EXAMINATION
30954-2|T077|strict|30954-2|LNC|LABORATORY TESTS|LABORATORY TESTS
30954-2|T077|strict|30954-2|LNC|LAB VALUES|LAB VALUES
30954-2|T077|strict|30954-2|LNC|CHEMISTRY STUDIES|CHEMISTRY STUDIES
30954-2|T077|multi|30954-2|LNC|STUDIES|STUDIES
30954-2|T077|multi|30954-2|LNC|LABORATORY INFORMATION|LABORATORY INFORMATION
30954-2|T077|strict|30954-2|LNC|LABORATORY RESULTS|LABORATORY RESULTS
30954-2|T077|strict|30954-2|LNC|LABORATORY STUDIES|LABORATORY STUDIES
30954-2|T077|strict|30954-2|LNC|LABORATORY VALUES|LABORATORY VALUES
30954-2|T077|strict|30954-2|LNC|BENIGN LABS|BENIGN LABS
30954-2|T077|strict|30954-2|LNC|NORMAL LABS|NORMAL LABS
30954-2|T077|multi|30954-2|LNC|RESULTS DIAGNOSTIC FINDINGS|RESULTS DIAGNOSTIC FINDINGS
30954-2|T077|multi|30954-2|LNC|LABS AND DIAGNOSTIC STUDIES|LABS AND DIAGNOSTIC STUDIES
30954-2|T077|multi|30954-2|LNC|DIAGNOSTIC STUDIES|DIAGNOSTIC STUDIES
30954-2|T077|multi|30954-2|LNC|DIAGNOSTIC DATA|DIAGNOSTIC DATA
30954-2|T077|multi|30954-2|LNC|DIAGNOSTIC TESTS|DIAGNOSTIC TESTS
30954-2|T077|multi|30954-2|LNC|SHOWED THE FOLLOWING RESULTS|SHOWED THE FOLLOWING RESULTS
30954-2|T077|multi|30954-2|LNC|RESULTS SUMMARY|RESULTS SUMMARY
30954-2|T077|multi|30954-2|LNC|TESTS|TESTS
30954-2|T077|multi|30954-2|LNC|RESULTS|RESULTS
30954-2|T077|multi|30954-2|LNC|OBSERVATIONS|OBSERVATIONS
30954-2|T077|multi|30954-2|LNC|PERTINENT RESULTS|PERTINENT RESULTS
30954-2|T077|multi|30954-2|LNC|TEST NAME|TEST NAME
30954-2|T077|multi|30954-2|LNC|RESULTS/INTERPRETATION|RESULTS/INTERPRETATION
30954-2|T077|strict|30954-2|LNC|LAB DATA|LAB DATA
30954-2|T077|strict|30954-2|LNC|LABORATORIES|LABORATORIES
30954-2|T077|strict|30954-2|LNC|LABORATORY|LABORATORY
30954-2|T077|strict|30954-2|LNC|CHEMISTRIES|CHEMISTRIES
30954-2|T077|strict|30954-2|LNC|LABORATORY STUDIES WERE SENT OFF INCLUDING|LABORATORY STUDIES WERE SENT OFF INCLUDING
30954-2|T077|strict|30954-2|LNC|FOLLOW-UP LABORATORY TESTING|FOLLOW-UP LABORATORY TESTING
30954-2|T077|strict|30954-2|LNC|FOLLOW UP LABORATORY TESTING|FOLLOW UP LABORATORY TESTING
30954-2|T077|strict|30954-2|LNC|FOLLOW UP LABS|FOLLOW UP LABS
30954-2|T077|strict|30954-2|LNC|LABS TO FU|LABS TO FU
30954-2|T077|multi|30954-2|LNC|LABS|LABS
30954-2|T077|multi|30954-2|LNC|LAB|LAB
30954-2|T077|strict|30954-2|LNC|LAB NO|LAB NO
30954-2|T077|strict|30954-2|LNC|LAB NO.|LAB NO.
82159-5|T077|strict|82159-5|LNC|RESPIRATORY PATHOGEN PROFILE, PCR|RESPIRATORY PATHOGEN PROFILE, PCR
82159-5|T077|strict|82159-5|LNC|ADENOVIRUS|ADENOVIRUS
82159-5|T077|strict|82159-5|LNC|CORONAVIRUS HKU1|CORONAVIRUS HKU1
82159-5|T077|strict|82159-5|LNC|HKU1|HKU1
82159-5|T077|strict|82159-5|LNC|CORONAVIRUS NL63|CORONAVIRUS NL63
82159-5|T077|strict|82159-5|LNC|NL63|NL63
82159-5|T077|strict|82159-5|LNC|CORONAVIRUS 229E|CORONAVIRUS 229E
82159-5|T077|strict|82159-5|LNC|229E|229E
82159-5|T077|strict|82159-5|LNC|CORONAVIRUS OC43|CORONAVIRUS OC43
82159-5|T077|strict|82159-5|LNC|OC43|OC43
82159-5|T077|strict|82159-5|LNC|HUMAN METAPNEUMOVIRUS|HUMAN METAPNEUMOVIRUS
82159-5|T077|strict|82159-5|LNC|HUMAN RHINOVIRUS/ENTEROVIRUS|HUMAN RHINOVIRUS/ENTEROVIRUS
82159-5|T077|strict|82159-5|LNC|RHINOVIRUS|RHINOVIRUS
82159-5|T077|strict|82159-5|LNC|ENTEROVIRUS|ENTEROVIRUS
82159-5|T077|strict|82159-5|LNC|INFLUENZA A|INFLUENZA A
82159-5|T077|strict|82159-5|LNC|INFLUENZA A/H1|INFLUENZA A/H1
82159-5|T077|strict|82159-5|LNC|INFLUENZA A/H1-2009|INFLUENZA A/H1-2009
82159-5|T077|strict|82159-5|LNC|INFLUENZA A/H3|INFLUENZA A/H3
82159-5|T077|strict|82159-5|LNC|INFLUENZA B|INFLUENZA B
82159-5|T077|strict|82159-5|LNC|PARAINFLUENZA 1|PARAINFLUENZA 1
82159-5|T077|strict|82159-5|LNC|PIVI|PIVI
82159-5|T077|strict|82159-5|LNC|PARAINFLUENZA 2|PARAINFLUENZA 2
82159-5|T077|strict|82159-5|LNC|PIV2|PIV2
82159-5|T077|strict|82159-5|LNC|PARAINFLUENZA 3|PARAINFLUENZA 3
82159-5|T077|strict|82159-5|LNC|PIV3|PIV3
82159-5|T077|strict|82159-5|LNC|PARAINFLUENZA 4|PARAINFLUENZA 4
82159-5|T077|strict|82159-5|LNC|PIV4|PIV4
82159-5|T077|strict|82159-5|LNC|RESPIRATORY SYNCYTIAL VIRUS|RESPIRATORY SYNCYTIAL VIRUS
82159-5|T077|strict|82159-5|LNC|RESP SYNCYTIAL VIRUS|RESP SYNCYTIAL VIRUS
82159-5|T077|strict|82159-5|LNC|BORDETELLA PERTUSSIS|BORDETELLA PERTUSSIS
82159-5|T077|strict|82159-5|LNC|BORDETELLA PARAPERTUSSIS|BORDETELLA PARAPERTUSSIS
82159-5|T077|strict|82159-5|LNC|CHLAMYDOPHILA PNEUMONIAE|CHLAMYDOPHILA PNEUMONIAE
82159-5|T077|strict|82159-5|LNC|MYCOPLASMA PNEUMONIAE|MYCOPLASMA PNEUMONIAE
77029-7|T077|strict|77029-7|LNC|RESPIRATORY PATHOGENS DNA AND RNA 14 PANEL|RESPIRATORY PATHOGENS DNA AND RNA 14 PANEL
50023-1|T077|strict|50023-1|LNC|HEPATITIS C VIRUS RNA PANEL|HEPATITIS C VIRUS RNA PANEL
50023-1|T077|strict|50023-1|LNC|VIRAL SCREENS AND IMMUNIZATIONS|VIRAL SCREENS AND IMMUNIZATIONS
664-3|T077|strict|664-3|LNC|GRAM STAIN FINAL|GRAM STAIN FINAL
664-3|T077|strict|664-3|LNC|GRAM STAIN|GRAM STAIN
11493-4|T077|strict|11493-4|LNC|HOSPITAL DISCHARGE STUDIES SUMMARY|HOSPITAL DISCHARGE STUDIES SUMMARY
11493-4|T077|strict|11493-4|LNC|DISCHARGE LAB DATA|DISCHARGE LAB DATA
11493-4|T077|strict|11493-4|LNC|DISCHARGE LABORATORIES|DISCHARGE LABORATORIES
11493-4|T077|strict|11493-4|LNC|DISCHARGE LABORATORY DATA|DISCHARGE LABORATORY DATA
11493-4|T077|strict|11493-4|LNC|DISCHARGE LABORATORY VALUES|DISCHARGE LABORATORY VALUES
11493-4|T077|strict|11493-4|LNC|DISCHARGE LABS|DISCHARGE LABS
11493-4|T077|strict|11493-4|LNC|LAB VALUES ON DAY OF DISCHARGE|LAB VALUES ON DAY OF DISCHARGE
11493-4|T077|strict|11493-4|LNC|LABORATORY DATA AT DISCHARGE|LABORATORY DATA AT DISCHARGE
11493-4|T077|strict|11493-4|LNC|LABORATORY DATA ON DISCHARGE|LABORATORY DATA ON DISCHARGE
11493-4|T077|strict|11493-4|LNC|LABORATORY VALUES ON DISCHARGE|LABORATORY VALUES ON DISCHARGE
11493-4|T077|strict|11493-4|LNC|LABORATORY STUDIES ON DISCHARGE|LABORATORY STUDIES ON DISCHARGE
11493-4|T077|strict|11493-4|LNC|LABORATORY STUDIES UPON DISCHARGE|LABORATORY STUDIES UPON DISCHARGE
11493-4|T077|strict|11493-4|LNC|LABS AT DISCHARGE|LABS AT DISCHARGE
11493-4|T077|strict|11493-4|LNC|LABS AT TIME OF DISCHARGE|LABS AT TIME OF DISCHARGE
11493-4|T077|strict|11493-4|LNC|LABS ON DAY OF DISCHARGE|LABS ON DAY OF DISCHARGE
11493-4|T077|strict|11493-4|LNC|LABS ON TRANSFER|LABS ON TRANSFER
11493-4|T077|strict|11493-4|LNC|LABORATORY PENDING ON DISCHARGE|LABORATORY PENDING ON DISCHARGE
61149-1|T077|multi|61149-1|LNC|OBJECTIVE|OBJECTIVE
61149-1|T077|multi|61149-1|LNC|OBJECTIVE DATA|OBJECTIVE DATA
18723-7|T077|strict|18723-7|LNC|HEMATOLOGY STUDIES|HEMATOLOGY STUDIES
18723-7|T077|strict|18723-7|LNC|HEMATOLOGY|HEMATOLOGY
18723-7|T077|strict|18723-7|LNC|HEMATOLOGIC|HEMATOLOGIC
18723-7|T077|strict|18723-7|LNC|COAGULATION STUDIES|COAGULATION STUDIES
18723-7|T077|multi|18723-7|LNC|HEME|HEME
56846-9|T077|multi|56846-9|LNC|CARDIAC BIOMARKERS|CARDIAC BIOMARKERS
56846-9|T077|multi|56846-9|LNC|LIPID PANEL|LIPID PANEL
56846-9|T077|multi|56846-9|LNC|METABOLIC PANEL|METABOLIC PANEL
56846-9|T077|multi|56846-9|LNC|CHOLESTEROL|CHOLESTEROL
18729-4|T077|strict|18729-4|LNC|URINALYSIS STUDIES|URINALYSIS STUDIES
18729-4|T077|strict|18729-4|LNC|URINALYSIS|URINALYSIS
18729-4|T077|strict|18729-4|LNC|UA ANALYSIS|UA ANALYSIS
18729-4|T077|strict|18729-4|LNC|URINE OUTPUT|URINE OUTPUT
18728-6|T077|strict|18728-6|LNC|TOXICOLOGY STUDIES|TOXICOLOGY STUDIES
18728-6|T077|strict|18728-6|LNC|TOXICOLOGY|TOXICOLOGY
56874-1|T077|multi|56874-1|LNC|SEROLOGY AND BLOOD BANK STUDIES|SEROLOGY AND BLOOD BANK STUDIES
56874-1|T077|multi|56874-1|LNC|SEROLOGY|SEROLOGY
56874-1|T077|multi|56874-1|LNC|IGG|IGG
56874-1|T077|multi|56874-1|LNC|IGM|IGM
56874-1|T077|multi|56874-1|LNC|IGG/IGM|IGG/IGM
56874-1|T077|multi|56874-1|LNC|IGG+IGM|IGG+IGM
56874-1|T077|multi|56874-1|LNC|ANTIBODIES|ANTIBODIES
18725-2|T077|strict|18725-2|LNC|MICROBIOLOGY STUDIES|MICROBIOLOGY STUDIES
18725-2|T077|multi|18725-2|LNC|MICROBIOLOGY|MICROBIOLOGY
56847-7|T077|strict|56847-7|LNC|CALCULATED AND DERIVED VALUES|CALCULATED AND DERIVED VALUES
56847-7|T077|strict|56847-7|LNC|DERIVED VALUES|DERIVED VALUES
19147-8|T077|strict|19147-8|LNC|REFERENCE LAB TEST REFERENCE RANGE|REFERENCE LAB TEST REFERENCE RANGE
19147-8|T077|strict|19147-8|LNC|REFERENCE RANGE|REFERENCE RANGE
19147-8|T077|strict|19147-8|LNC|REFERENCE|REFERENCE
19147-8|T077|strict|19147-8|LNC|RANGE|RANGE
94531-1|T077|strict|94531-1|LNC|SARS CORONAVIRUS 2 RNA PANEL|SARS CORONAVIRUS 2 RNA PANEL
94531-1|T077|strict|94531-1|LNC|2019 NOVEL CORONAVIRUS|2019 NOVEL CORONAVIRUS
94531-1|T077|strict|94531-1|LNC|SARS-COV-2 RNA|SARS-COV-2 RNA
94531-1|T077|multi|94531-1|LNC|RTPCR|RTPCR
94531-1|T077|strict|94531-1|LNC|PCR|PCR
94531-1|T077|strict|94531-1|LNC|NAA|NAA
94531-1|T077|multi|94531-1|LNC|COVID-19|COVID-19
94531-1|T077|multi|94531-1|LNC|COVID19|COVID19
94531-1|T077|strict|94531-1|LNC|COVID19|COVID19
94531-1|T077|strict|94531-1|LNC|COVID+|COVID+
94531-1|T077|strict|94531-1|LNC|COVID|COVID
94531-1|T077|multi|94531-1|LNC|SARS-COV|SARS-COV
94531-1|T077|multi|94531-1|LNC|SARS-COV-2|SARS-COV-2
94531-1|T077|strict|94531-1|LNC|MERS-COV|MERS-COV
94531-1|T077|strict|94531-1|LNC|SARS-COV|SARS-COV
94531-1|T077|strict|94531-1|LNC|CORONAVIRUS|CORONAVIRUS
94531-1|T077|strict|94531-1|LNC|HKU1|HKU1
94531-1|T077|strict|94531-1|LNC|NL63|NL63
94531-1|T077|strict|94531-1|LNC|229E|229E
94531-1|T077|strict|94531-1|LNC|OC43|OC43
11502-2|T077|multi|11502-2|LNC|LABORATORY REPORT (COLUMNS)|LABORATORY REPORT (COLUMNS)
11502-2|T077|multi|11502-2|LNC|REFERENCE RANGE|REFERENCE RANGE
11502-2|T077|multi|11502-2|LNC|COMPONENT|COMPONENT
11502-2|T077|multi|11502-2|LNC|RANGE|RANGE
11502-2|T077|multi|11502-2|LNC|FLAG|FLAG
92236-9|T077|multi|92236-9|LNC|RESULT STATUS|RESULT STATUS
92236-9|T077|multi|92236-9|LNC|RESULT TYPE|RESULT TYPE
92236-9|T077|multi|92236-9|LNC|RESULT DATE|RESULT DATE
92236-9|T077|multi|92236-9|LNC|RESULT STATUS|RESULT STATUS
92236-9|T077|multi|92236-9|LNC|RESULTED|RESULTED
92236-9|T077|multi|92236-9|LNC|RESULT TITLE|RESULT TITLE
19005-8|T077|strict|19005-8|LNC|RADIOLOGY IMAGING STUDY IMPRESSION|RADIOLOGY IMAGING STUDY IMPRESSION
18783-1|T077|strict|18783-1|LNC|RADIOLOGY STUDY RECOMMENDATION|RADIOLOGY STUDY RECOMMENDATION
18834-2|T077|strict|18834-2|LNC|RADIOLOGY COMPARISON STUDY OBSERVATION|RADIOLOGY COMPARISON STUDY OBSERVATION
18834-2|T077|strict|18834-2|LNC|COMPARISON|COMPARISON
55111-9|T077|multi|55111-9|LNC|CURRENT IMAGING PROCEDURE DESCRIPTIONS|CURRENT IMAGING PROCEDURE DESCRIPTIONS
55111-9|T077|multi|55111-9|LNC|CURRENT IMAGING PROCEDURE|CURRENT IMAGING PROCEDURE
55111-9|T077|multi|55111-9|LNC|DIAGNOSTIC PROCEDURE|DIAGNOSTIC PROCEDURE
55115-0|T077|strict|55115-0|LNC|REQUESTED IMAGING STUDIES INFORMATION|REQUESTED IMAGING STUDIES INFORMATION
55115-0|T077|strict|55115-0|LNC|REQUESTED IMAGING STUDIES|REQUESTED IMAGING STUDIES
55115-0|T077|strict|55115-0|LNC|IMAGING STUDIES|IMAGING STUDIES
55115-0|T077|strict|55115-0|LNC|RADIOGRAPHIC STUDIES|RADIOGRAPHIC STUDIES
55115-0|T077|strict|55115-0|LNC|RADIOLOGIC STUDIES|RADIOLOGIC STUDIES
55115-0|T077|strict|55115-0|LNC|RADIOLOGY IMAGING|RADIOLOGY IMAGING
55115-0|T077|strict|55115-0|LNC|IMAGING RESULTS|IMAGING RESULTS
55115-0|T077|strict|55115-0|LNC|RELEVANT IMAGING|RELEVANT IMAGING
55115-0|T077|strict|55115-0|LNC|RADIOGRAPHIC|RADIOGRAPHIC
55115-0|T077|multi|55115-0|LNC|RADIOLOGY|RADIOLOGY
55115-0|T077|multi|55115-0|LNC|IMAGING|IMAGING
55115-0|T077|strict|55115-0|LNC|ECG|ECG
55115-0|T077|strict|55115-0|LNC|EKG|EKG
55115-0|T077|strict|55115-0|LNC|ECHO|ECHO
55115-0|T077|strict|55115-0|LNC|ELECTROCARDIOGRAM|ELECTROCARDIOGRAM
55115-0|T077|strict|55115-0|LNC|CXR|CXR
55115-0|T077|strict|55115-0|LNC|CHEST XRAY|CHEST XRAY
55115-0|T077|strict|55115-0|LNC|X-RAY|X-RAY
55115-0|T077|strict|55115-0|LNC|XRAY|XRAY
55115-0|T077|strict|55115-0|LNC|XR|XR
55115-0|T077|strict|55115-0|LNC|KUB|KUB
55115-0|T077|strict|55115-0|LNC|MRA KIDNEY|MRA KIDNEY
55115-0|T077|strict|55115-0|LNC|MRI|MRI
55115-0|T077|strict|55115-0|LNC|MRI HEAD|MRI HEAD
55113-5|T077|strict|55113-5|LNC|KEY IMAGES|KEY IMAGES
75321-0|T077|multi|75321-0|LNC|CLINICAL FINDING|CLINICAL FINDING
75321-0|T077|multi|75321-0|LNC|FINDINGS|FINDINGS
59776-5|T077|multi|59776-5|LNC|PROCEDURE FINDINGS|PROCEDURE FINDINGS
59776-5|T077|strict|59776-5|LNC|OPERATIVE FINDINGS|OPERATIVE FINDINGS
18782-3|T077|strict|18782-3|LNC|RADIOLOGY STUDY OBSERVATION FINDINGS|RADIOLOGY STUDY OBSERVATION FINDINGS
22029-3|T077|strict|22029-3|LNC|PHYSICAL EXAM|PHYSICAL EXAM
22029-3|T077|strict|22029-3|LNC|HEAD EYES EARS NOSE THROAT|HEAD EYES EARS NOSE THROAT
22029-3|T077|strict|22029-3|LNC|ADMISSION PHYSICAL EXAMINATION|ADMISSION PHYSICAL EXAMINATION
22029-3|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION|PHYSICAL EXAMINATION
22029-3|T077|strict|22029-3|LNC|PHYSICAL EXAM ON ADMISSION|PHYSICAL EXAM ON ADMISSION
22029-3|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION ON ADMISSION|PHYSICAL EXAMINATION ON ADMISSION
22029-3|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION UPON ADMISSION|PHYSICAL EXAMINATION UPON ADMISSION
22029-3|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION ON DISCHARGE|PHYSICAL EXAMINATION ON DISCHARGE
22029-3|T077|strict|22029-3|LNC|HOSPITAL DISCHARGE PHYSICAL|HOSPITAL DISCHARGE PHYSICAL
22029-3|T077|strict|22029-3|LNC|PHYSICAL EXAMINATION ON PRESENTATION|PHYSICAL EXAMINATION ON PRESENTATION
10184-0|T077|strict|10184-0|LNC|HOSPITAL DISCHARGE PHYSICAL FINDINGS|HOSPITAL DISCHARGE PHYSICAL FINDINGS
10210-3|T077|strict|10210-3|LNC|PHYSICAL FINDINGS OF GENERAL STATUS|PHYSICAL FINDINGS OF GENERAL STATUS
10210-3|T077|multi|10210-3|LNC|GENERAL STATUS|GENERAL STATUS
10187-3|T077|strict|10187-3|LNC|REVIEW OF SYSTEMS|REVIEW OF SYSTEMS
10187-3|T077|strict|10187-3|LNC|GENERAL ROS|GENERAL ROS
10187-3|T077|strict|10187-3|LNC|ROS|ROS
10190-7|T077|strict|10190-7|LNC|MENTAL STATUS|MENTAL STATUS
29545-1|T077|strict|29545-1|LNC|PHYSICAL FINDINGS|PHYSICAL FINDINGS
29545-1|T077|strict|29545-1|LNC|PHYS FIND|PHYS FIND
11384-5|T077|multi|11384-5|LNC|EXAM|EXAM
11384-5|T077|multi|11384-5|LNC|EXAMINATION|EXAMINATION
11384-5|T077|multi|11384-5|LNC|ABD|ABD
11384-5|T077|multi|11384-5|LNC|ABDOMEN|ABDOMEN
11384-5|T077|multi|11384-5|LNC|ADNEXA|ADNEXA
11384-5|T077|multi|11384-5|LNC|APPEARANCE|APPEARANCE
11384-5|T077|multi|11384-5|LNC|BACK|BACK
11384-5|T077|multi|11384-5|LNC|BMI|BMI
11384-5|T077|multi|11384-5|LNC|BODY MASS INDEX|BODY MASS INDEX
11384-5|T077|multi|11384-5|LNC|BREASTS|BREASTS
11384-5|T077|multi|11384-5|LNC|CHEST|CHEST
11384-5|T077|multi|11384-5|LNC|CARDIAC|CARDIAC
11384-5|T077|multi|11384-5|LNC|CARDIAC EXAMINATION|CARDIAC EXAMINATION
11384-5|T077|multi|11384-5|LNC|CARDS|CARDS
11384-5|T077|multi|11384-5|LNC|CVS|CVS
11384-5|T077|multi|11384-5|LNC|CARDIOVASCULAR|CARDIOVASCULAR
11384-5|T077|multi|11384-5|LNC|CARDIOVASCULAR EXAM|CARDIOVASCULAR EXAM
11384-5|T077|multi|11384-5|LNC|CARDIOVASCULAR STATUS|CARDIOVASCULAR STATUS
11384-5|T077|multi|11384-5|LNC|CAROTIDS|CAROTIDS
11384-5|T077|multi|11384-5|LNC|CEREBELLAR EXAM|CEREBELLAR EXAM
11384-5|T077|multi|11384-5|LNC|COORDINATION|COORDINATION
11384-5|T077|multi|11384-5|LNC|CRANIAL|CRANIAL
11384-5|T077|multi|11384-5|LNC|CRANIAL NERVES|CRANIAL NERVES
11384-5|T077|multi|11384-5|LNC|EAR/NOSE/THROAT|EAR/NOSE/THROAT
11384-5|T077|multi|11384-5|LNC|ENDO|ENDO
11384-5|T077|multi|11384-5|LNC|ENDOCRINE|ENDOCRINE
11384-5|T077|multi|11384-5|LNC|EXTREMITIES|EXTREMITIES
11384-5|T077|multi|11384-5|LNC|EXTREMITY EXAM|EXTREMITY EXAM
11384-5|T077|multi|11384-5|LNC|EYE EXAM|EYE EXAM
11384-5|T077|multi|11384-5|LNC|EYES|EYES
11384-5|T077|multi|11384-5|LNC|FOOT EXAM|FOOT EXAM
11384-5|T077|multi|11384-5|LNC|FUNCTIONAL AND COGNITIVE STATUS|FUNCTIONAL AND COGNITIVE STATUS
11384-5|T077|multi|11384-5|LNC|COGNITION|COGNITION
11384-5|T077|multi|11384-5|LNC|GAIT|GAIT
11384-5|T077|multi|11384-5|LNC|GEN|GEN
11384-5|T077|multi|11384-5|LNC|GENERAL|GENERAL
11384-5|T077|multi|11384-5|LNC|GENITOURINARY|GENITOURINARY
11384-5|T077|multi|11384-5|LNC|GI|GI
11384-5|T077|multi|11384-5|LNC|GASTROINTESTINAL|GASTROINTESTINAL
11384-5|T077|multi|11384-5|LNC|GU|GU
11384-5|T077|multi|11384-5|LNC|HEAD EYES EARS NOSE AND THROAT|HEAD EYES EARS NOSE AND THROAT
11384-5|T077|multi|11384-5|LNC|HEAD EYES EARS NOSE AND THROAT EXAM|HEAD EYES EARS NOSE AND THROAT EXAM
11384-5|T077|multi|11384-5|LNC|HEENT|HEENT
11384-5|T077|multi|11384-5|LNC|HENT|HENT
11384-5|T077|multi|11384-5|LNC|EARS|EARS
11384-5|T077|multi|11384-5|LNC|LEFT EAR|LEFT EAR
11384-5|T077|multi|11384-5|LNC|RIGHT EAR|RIGHT EAR
11384-5|T077|multi|11384-5|LNC|HEART|HEART
11384-5|T077|multi|11384-5|LNC|HEMODYNAMICS|HEMODYNAMICS
11384-5|T077|multi|11384-5|LNC|INITIAL NEWBORN EXAM|INITIAL NEWBORN EXAM
11384-5|T077|multi|11384-5|LNC|LUNGS|LUNGS
11384-5|T077|multi|11384-5|LNC|LYMPH|LYMPH
11384-5|T077|multi|11384-5|LNC|LYMPH NODES|LYMPH NODES
11384-5|T077|multi|11384-5|LNC|NODES|NODES
11384-5|T077|multi|11384-5|LNC|MENTAL STATUS EXAMINATION|MENTAL STATUS EXAMINATION
11384-5|T077|multi|11384-5|LNC|MSK|MSK
11384-5|T077|multi|11384-5|LNC|MUSCULOSKELETAL|MUSCULOSKELETAL
11384-5|T077|multi|11384-5|LNC|NECK|NECK
11384-5|T077|multi|11384-5|LNC|NEUROLOGICAL EXAMINATION|NEUROLOGICAL EXAMINATION
11384-5|T077|multi|11384-5|LNC|NEURO|NEURO
11384-5|T077|multi|11384-5|LNC|NEUROLOGICAL|NEUROLOGICAL
11384-5|T077|multi|11384-5|LNC|NEUROLOGIC|NEUROLOGIC
11384-5|T077|multi|11384-5|LNC|NEUROLOGIC EXAM|NEUROLOGIC EXAM
11384-5|T077|multi|11384-5|LNC|NEUROLOGY|NEUROLOGY
11384-5|T077|multi|11384-5|LNC|OPHTHALMOLOGY|OPHTHALMOLOGY
11384-5|T077|multi|11384-5|LNC|PE|PE
11384-5|T077|multi|11384-5|LNC|PELVIC|PELVIC
11384-5|T077|multi|11384-5|LNC|PSYCH|PSYCH
11384-5|T077|multi|11384-5|LNC|PSYCHOSOCIAL|PSYCHOSOCIAL
11384-5|T077|multi|11384-5|LNC|PULM|PULM
11384-5|T077|multi|11384-5|LNC|PULMONARY|PULMONARY
11384-5|T077|multi|11384-5|LNC|PULSE|PULSE
11384-5|T077|multi|11384-5|LNC|PUPILS|PUPILS
11384-5|T077|multi|11384-5|LNC|RECTAL|RECTAL
11384-5|T077|multi|11384-5|LNC|REFLEXES|REFLEXES
11384-5|T077|multi|11384-5|LNC|RENAL|RENAL
11384-5|T077|multi|11384-5|LNC|RESP|RESP
11384-5|T077|multi|11384-5|LNC|RESPIRATORY|RESPIRATORY
11384-5|T077|multi|11384-5|LNC|SENSORY|SENSORY
11384-5|T077|multi|11384-5|LNC|SENSORY EXAMINATION|SENSORY EXAMINATION
11384-5|T077|multi|11384-5|LNC|SKIN|SKIN
11384-5|T077|multi|11384-5|LNC|SPINE|SPINE
10154-3|T077|strict|10154-3|LNC|CHIEF COMPLAINT|CHIEF COMPLAINT
10154-3|T077|strict|10154-3|LNC|PATIENT COMPLAINT|PATIENT COMPLAINT
10154-3|T077|strict|10154-3|LNC|PATIENT STATES COMPLAINT|PATIENT STATES COMPLAINT
10154-3|T077|strict|10154-3|LNC|COMPLAINTS|COMPLAINTS
10154-3|T077|multi|10154-3|LNC|CC|CC
46239-0|T077|strict|46239-0|LNC|REASON FOR VISIT AND CHIEF COMPLAINT|REASON FOR VISIT AND CHIEF COMPLAINT
46239-0|T077|strict|46239-0|LNC|REASON FOR VISIT/CHIEF COMPLAINT|REASON FOR VISIT/CHIEF COMPLAINT
46239-0|T077|strict|46239-0|LNC|CHIEF COMPLAINT AND REASON FOR VISIT|CHIEF COMPLAINT AND REASON FOR VISIT
46239-0|T077|strict|46239-0|LNC|CHIEF COMPLAINT REASON FOR VISIT|CHIEF COMPLAINT REASON FOR VISIT
75325-1|T077|strict|75325-1|LNC|SYMPTOM|SYMPTOM
75325-1|T077|strict|75325-1|LNC|SYMPTOMS|SYMPTOMS
75325-1|T077|strict|75325-1|LNC|PATIENT SYMPTOMS|PATIENT SYMPTOMS
29299-5|T077|strict|29299-5|LNC|REASON FOR VISIT|REASON FOR VISIT
29299-5|T077|strict|29299-5|LNC|REASON FOR ADMISSION|REASON FOR ADMISSION
29299-5|T077|strict|29299-5|LNC|HISTORY AND REASON FOR HOSPITALIZATION|HISTORY AND REASON FOR HOSPITALIZATION
29299-5|T077|strict|29299-5|LNC|REASON FOR HOSPITALIZATION|REASON FOR HOSPITALIZATION
29299-5|T077|strict|29299-5|LNC|HISTORY AND REASON FOR ADMISSION|HISTORY AND REASON FOR ADMISSION
29299-5|T077|strict|29299-5|LNC|HISTORY REASON FOR HOSPITALIZATION|HISTORY REASON FOR HOSPITALIZATION
42349-1|T077|strict|42349-1|LNC|REASON FOR CONSULT|REASON FOR CONSULT
42349-1|T077|strict|42349-1|LNC|REASON FOR CONSULTATION|REASON FOR CONSULTATION
42349-1|T077|strict|42349-1|LNC|REASON FOR REFERRAL|REASON FOR REFERRAL
42349-1|T077|strict|42349-1|LNC|REASON FOR CLINIC VISIT|REASON FOR CLINIC VISIT
42349-1|T077|strict|42349-1|LNC|REASON FOR APPOINTMENT|REASON FOR APPOINTMENT
42349-1|T077|strict|42349-1|LNC|REASON FOR EXAM|REASON FOR EXAM
42349-1|T077|strict|42349-1|LNC|REASON FOR THIS EXAMINATION|REASON FOR THIS EXAMINATION
59768-2|T077|strict|59768-2|LNC|PROCEDURE INDICATION|PROCEDURE INDICATION
59768-2|T077|strict|59768-2|LNC|PROCEDURE INDICATIONS|PROCEDURE INDICATIONS
59768-2|T077|strict|59768-2|LNC|INDICATION FOR PROCEDURE|INDICATION FOR PROCEDURE
59768-2|T077|strict|59768-2|LNC|INDICATION FOR SURGERY|INDICATION FOR SURGERY
59768-2|T077|strict|59768-2|LNC|INDICATION FOR INDUCTION|INDICATION FOR INDUCTION
59768-2|T077|strict|59768-2|LNC|INDICATION FOR OPERATION|INDICATION FOR OPERATION
59768-2|T077|strict|59768-2|LNC|INDICATION FOR TESTING|INDICATION FOR TESTING
59768-2|T077|strict|59768-2|LNC|INDICATION FOR TEST|INDICATION FOR TEST
59768-2|T077|strict|59768-2|LNC|TEST INDICATION|TEST INDICATION
59768-2|T077|multi|59768-2|LNC|INDICATION|INDICATION
59768-2|T077|multi|59768-2|LNC|INDICATION|INDICATION
59768-2|T077|strict|59768-2|LNC|PROCEDURE INDICATIONS INTERPRETATION|PROCEDURE INDICATIONS INTERPRETATION
18785-6|T077|strict|18785-6|LNC|RADIOLOGY REASON FOR STUDY|RADIOLOGY REASON FOR STUDY
11450-4|T077|strict|11450-4|LNC|PROBLEM LIST|PROBLEM LIST
11450-4|T077|strict|11450-4|LNC|LIST OF PROBLEM|LIST OF PROBLEM
11450-4|T077|strict|11450-4|LNC|LIST OF PROBLEMS|LIST OF PROBLEMS
11450-4|T077|strict|11450-4|LNC|PROBLEMS BY SYSTEMS|PROBLEMS BY SYSTEMS
11450-4|T077|strict|11450-4|LNC|PROBLEMS BY SYSTEM|PROBLEMS BY SYSTEM
11450-4|T077|strict|11450-4|LNC|PROBLEM LIST AND DIAGNOSIS|PROBLEM LIST AND DIAGNOSIS
11450-4|T077|strict|11450-4|LNC|PROBLEMS AND DIAGNOSIS|PROBLEMS AND DIAGNOSIS
11450-4|T077|strict|11450-4|LNC|LIST OF PROBLEMS DURING ADMISSION|LIST OF PROBLEMS DURING ADMISSION
11450-4|T077|strict|11450-4|LNC|LIST OF PROBLEMS DURING HOSPITALIZATION|LIST OF PROBLEMS DURING HOSPITALIZATION
11450-4|T077|strict|11450-4|LNC|HOSPITAL PROBLEM LIST|HOSPITAL PROBLEM LIST
11450-4|T077|strict|11450-4|LNC|ACTIVE PROBLEMS LIST|ACTIVE PROBLEMS LIST
11450-4|T077|strict|11450-4|LNC|ACTIVE PROBLEMS|ACTIVE PROBLEMS
11450-4|T077|strict|11450-4|LNC|PRINCIPAL PROBLEM|PRINCIPAL PROBLEM
11450-4|T077|strict|11450-4|LNC|SIGNIFICANT PROBLEMS|SIGNIFICANT PROBLEMS
11450-4|T077|strict|11450-4|LNC|OTHER SIGNIFICANT PROBLEMS|OTHER SIGNIFICANT PROBLEMS
11450-4|T077|strict|11450-4|LNC|OTHER PROBLEMS|OTHER PROBLEMS
11450-4|T077|strict|11450-4|LNC|OTHER ASSOCIATED PROBLEMS|OTHER ASSOCIATED PROBLEMS
11450-4|T077|strict|11450-4|LNC|PROBLEM CARDIOVASCULAR|PROBLEM CARDIOVASCULAR
11450-4|T077|strict|11450-4|LNC|NEW PROBLEMS|NEW PROBLEMS
11450-4|T077|strict|11450-4|LNC|SPONTANEOUS CONDITION|SPONTANEOUS CONDITION
11450-4|T077|strict|11450-4|LNC|UNDERLYING MEDICAL CONDITION|UNDERLYING MEDICAL CONDITION
11450-4|T077|strict|11450-4|LNC|MEDICAL PROBLEMS|MEDICAL PROBLEMS
11450-4|T077|strict|11450-4|LNC|PROBLEM|PROBLEM
11450-4|T077|strict|11450-4|LNC|PROBLEMS|PROBLEMS
11450-4|T077|strict|11450-4|LNC|CONDITIONS|CONDITIONS
61133-5|T077|strict|61133-5|LNC|PRIMARY PROBLEM INTERPRETATION|PRIMARY PROBLEM INTERPRETATION
61133-5|T077|strict|61133-5|LNC|IMPRESSION ON ADMISSION|IMPRESSION ON ADMISSION
61133-5|T077|strict|61133-5|LNC|CLINICAL IMPRESSION|CLINICAL IMPRESSION
61133-5|T077|strict|61133-5|LNC|IMPRESSION|IMPRESSION
51898-5|T077|strict|51898-5|LNC|RISK FACTORS|RISK FACTORS
51898-5|T077|strict|51898-5|LNC|CARDIAC RISK FACTORS|CARDIAC RISK FACTORS
51898-5|T077|strict|51898-5|LNC|CORONARY RISK FACTORS|CORONARY RISK FACTORS
51898-5|T077|strict|51898-5|LNC|HYPERTENSIVE URGENCY|HYPERTENSIVE URGENCY
51898-5|T077|strict|51898-5|LNC|HYPERGLYCEMIC SYMPTOMS|HYPERGLYCEMIC SYMPTOMS
10157-6|T077|strict|10157-6|LNC|HISTORY OF FAMILY MEMBER DISEASES|HISTORY OF FAMILY MEMBER DISEASES
10157-6|T077|strict|10157-6|LNC|FAMILY HISTORY|FAMILY HISTORY
10157-6|T077|strict|10157-6|LNC|FHX|FHX
10157-6|T077|strict|10157-6|LNC|FATHER|FATHER
10157-6|T077|strict|10157-6|LNC|MOTHER|MOTHER
10157-6|T077|strict|10157-6|LNC|SIBLINGS|SIBLINGS
10157-6|T077|strict|10157-6|LNC|SPOUSE|SPOUSE
10157-6|T077|strict|10157-6|LNC|OFFSPRING|OFFSPRING
10157-6|T077|strict|10157-6|LNC|PEDIGREE|PEDIGREE
32435-0|T077|multi|32435-0|LNC|HISTORY OF HEREDITARY DISORDERS|HISTORY OF HEREDITARY DISORDERS
32435-0|T077|multi|32435-0|LNC|HEREDITARY|HEREDITARY
32435-0|T077|multi|32435-0|LNC|ANCESTRAL|ANCESTRAL
32435-0|T077|multi|32435-0|LNC|ANCESTRY|ANCESTRY
32435-0|T077|multi|32435-0|LNC|HEREDITARY|HEREDITARY
32435-0|T077|multi|32435-0|LNC|INHERITANCE|INHERITANCE
10164-2|T077|strict|10164-2|LNC|HISTORY OF PRESENT ILLNESS|HISTORY OF PRESENT ILLNESS
10164-2|T077|strict|10164-2|LNC|HPI|HPI
10164-2|T077|strict|10164-2|LNC|HX PRESENT ILLNESS|HX PRESENT ILLNESS
10164-2|T077|strict|10164-2|LNC|HX OF PRES ILLNESS|HX OF PRES ILLNESS
10164-2|T077|strict|10164-2|LNC|HX OF PRESENT ILLNESS|HX OF PRESENT ILLNESS
10164-2|T077|strict|10164-2|LNC|HISTORY PRESENT ILLNESS|HISTORY PRESENT ILLNESS
10164-2|T077|strict|10164-2|LNC|BRIEF HISTORY OF PHYSICAL ILLNESS|BRIEF HISTORY OF PHYSICAL ILLNESS
10164-2|T077|strict|10164-2|LNC|BRIEF ADMISSION HISTORY OF PRESENT ILLNESS|BRIEF ADMISSION HISTORY OF PRESENT ILLNESS
10164-2|T077|strict|10164-2|LNC|BRIEF HISTORY OF PRESENT ILLNESS|BRIEF HISTORY OF PRESENT ILLNESS
10164-2|T077|multi|10164-2|LNC|HISTORY OF PRESENT ILLNESS AND HOSPITAL COURSE|HISTORY OF PRESENT ILLNESS AND HOSPITAL COURSE
10164-2|T077|strict|10164-2|LNC|HISTORY OF PRESENT ILLNESS AND REASON FOR HOSPITALIZATION|HISTORY OF PRESENT ILLNESS AND REASON FOR HOSPITALIZATION
10164-2|T077|strict|10164-2|LNC|HISTORY OF PRESENTING ILLNESS|HISTORY OF PRESENTING ILLNESS
10164-2|T077|strict|10164-2|LNC|HISTORY OF THE PRESENT ILLNESS|HISTORY OF THE PRESENT ILLNESS
10164-2|T077|strict|10164-2|LNC|HISTORY AND PHYSICAL HISTORY OF PRESENT ILLNESS|HISTORY AND PHYSICAL HISTORY OF PRESENT ILLNESS
10164-2|T077|strict|10164-2|LNC|HEALTH CONCERNS|HEALTH CONCERNS
10164-2|T077|strict|10164-2|LNC|HISTORY AND PHYSICAL|HISTORY AND PHYSICAL
10164-2|T077|strict|10164-2|LNC|HISTORY AND PHYSICALS|HISTORY AND PHYSICALS
10164-2|T077|strict|10164-2|LNC|H&P|H&P
10164-2|T077|strict|10164-2|LNC|H&P BY|H&P BY
10164-2|T077|strict|10164-2|LNC|BRIEF HISTORY|BRIEF HISTORY
10164-2|T077|strict|10164-2|LNC|PRESENT ILLNESS|PRESENT ILLNESS
61150-9|T077|multi|61150-9|LNC|SUBJECTIVE DATA|SUBJECTIVE DATA
61150-9|T077|multi|61150-9|LNC|SUBJECTIVE|SUBJECTIVE
51848-0|T077|multi|51848-0|LNC|EVALUATION NOTE|EVALUATION NOTE
51848-0|T077|strict|51848-0|LNC|EVALUATION|EVALUATION
51848-0|T077|multi|51848-0|LNC|EVAL NOTE|EVAL NOTE
51848-0|T077|multi|51848-0|LNC|ASSESSMENT/PLAN|ASSESSMENT/PLAN
51848-0|T077|strict|51848-0|LNC|ASSESSMENT|ASSESSMENT
51848-0|T077|multi|51848-0|LNC|ASSESSMENTS|ASSESSMENTS
61146-7|T077|strict|61146-7|LNC|GOALS|GOALS
61146-7|T077|strict|61146-7|LNC|SHORT TERM GOAL|SHORT TERM GOAL
61146-7|T077|strict|61146-7|LNC|LONG TERM GOAL|LONG TERM GOAL
61146-7|T077|strict|61146-7|LNC|GOAL|GOAL
61146-7|T077|strict|61146-7|LNC|GOALS|GOALS
61146-7|T077|strict|61146-7|LNC|GOAL DATE|GOAL DATE
55108-5|T077|multi|55108-5|LNC|CLINICAL PRESENTATIONS|CLINICAL PRESENTATIONS
55108-5|T077|multi|55108-5|LNC|CLINICAL PRESENTATION|CLINICAL PRESENTATION
55109-3|T077|strict|55109-3|LNC|COMPLICATIONS DOCUMENT|COMPLICATIONS DOCUMENT
55109-3|T077|strict|55109-3|LNC|COMPLICATIONS|COMPLICATIONS
55109-3|T077|strict|55109-3|LNC|CONCERNS|CONCERNS
55752-0|T077|multi|55752-0|LNC|CLINICAL INFORMATION|CLINICAL INFORMATION
55752-0|T077|multi|55752-0|LNC|CLINICAL DATA|CLINICAL DATA
11329-0|T077|multi|11329-0|LNC|HISTORY GENERAL|HISTORY GENERAL
11329-0|T077|multi|11329-0|LNC|MEDICAL GENERAL HISTORY|MEDICAL GENERAL HISTORY
11329-0|T077|multi|11329-0|LNC|GENERAL HISTORY|GENERAL HISTORY
11329-0|T077|multi|11329-0|LNC|BRIEF HISTORY|BRIEF HISTORY
8648-8|T077|strict|8648-8|LNC|HOSPITAL COURSE|HOSPITAL COURSE
8648-8|T077|strict|8648-8|LNC|HOSPITAL COURSE BY SYSTEM|HOSPITAL COURSE BY SYSTEM
8648-8|T077|strict|8648-8|LNC|HOSPITAL COURSE BY SYSTEMS|HOSPITAL COURSE BY SYSTEMS
8648-8|T077|strict|8648-8|LNC|SUMMARY OF HOSPITAL COURSE|SUMMARY OF HOSPITAL COURSE
8648-8|T077|strict|8648-8|LNC|COURSE BY PROBLEM|COURSE BY PROBLEM
8648-8|T077|strict|8648-8|LNC|BRIEF HOSPITAL COURSE|BRIEF HOSPITAL COURSE
8648-8|T077|strict|8648-8|LNC|EMERGENCY DEPARTMENT COURSE|EMERGENCY DEPARTMENT COURSE
8648-8|T077|strict|8648-8|LNC|HOSPITAL COURSE BY PROBLEM|HOSPITAL COURSE BY PROBLEM
8648-8|T077|strict|8648-8|LNC|HOSPITAL COURSE BY PROBLEMS|HOSPITAL COURSE BY PROBLEMS
8648-8|T077|strict|8648-8|LNC|HOSPITAL COURSE BY SYSTEM AND PROBLEM|HOSPITAL COURSE BY SYSTEM AND PROBLEM
8648-8|T077|strict|8648-8|LNC|HOSPITAL COURSE AND TREATMENT|HOSPITAL COURSE AND TREATMENT
55112-7|T077|strict|55112-7|LNC|DOCUMENT SUMMARY|DOCUMENT SUMMARY
55112-7|T077|strict|55112-7|LNC|DISCUSSION|DISCUSSION
55112-7|T077|strict|55112-7|LNC|SUMMARY|SUMMARY
46241-6|T077|strict|46241-6|LNC|HOSPITAL ADMISSION DIAGNOSIS|HOSPITAL ADMISSION DIAGNOSIS
46241-6|T077|strict|46241-6|LNC|HOSPITAL ADMISSION DX|HOSPITAL ADMISSION DX
11535-2|T077|strict|11535-2|LNC|HOSPITAL DISCHARGE DX|HOSPITAL DISCHARGE DX
11535-2|T077|strict|11535-2|LNC|HOSPITAL DISCHARGE DIAGNOSIS|HOSPITAL DISCHARGE DIAGNOSIS
42347-5|T077|strict|42347-5|LNC|ADMISSION DIAGNOSIS|ADMISSION DIAGNOSIS
42347-5|T077|strict|42347-5|LNC|ADMISSION DIAGNOSES|ADMISSION DIAGNOSES
42347-5|T077|strict|42347-5|LNC|ADMIT DIAGNOSIS|ADMIT DIAGNOSIS
42347-5|T077|strict|42347-5|LNC|ADMIT DIAGNOSES|ADMIT DIAGNOSES
42347-5|T077|strict|42347-5|LNC|ADMITTING DIAGNOSIS|ADMITTING DIAGNOSIS
42347-5|T077|strict|42347-5|LNC|ADMITTING DIAGNOSES|ADMITTING DIAGNOSES
42347-5|T077|strict|42347-5|LNC|LIST OF DIAGNOSIS DURING ADMISSION|LIST OF DIAGNOSIS DURING ADMISSION
42347-5|T077|strict|42347-5|LNC|PRINCIPAL ADMISSION DIAGNOSIS|PRINCIPAL ADMISSION DIAGNOSIS
42347-5|T077|strict|42347-5|LNC|PRINCIPAL DIAGNOSIS FOR ADMISSION|PRINCIPAL DIAGNOSIS FOR ADMISSION
42347-5|T077|strict|42347-5|LNC|PRINCIPAL DIAGNOSIS ON ADMISSION|PRINCIPAL DIAGNOSIS ON ADMISSION
42347-5|T077|strict|42347-5|LNC|PRIMARY ADMISSION DIAGNOSIS|PRIMARY ADMISSION DIAGNOSIS
42347-5|T077|strict|42347-5|LNC|PRIMARY ADMITTING DIAGNOSIS|PRIMARY ADMITTING DIAGNOSIS
42347-5|T077|strict|42347-5|LNC|PRIMARY DIAGNOSIS DURING THIS ADMISSION|PRIMARY DIAGNOSIS DURING THIS ADMISSION
42347-5|T077|strict|42347-5|LNC|PRIMARY DIAGNOSIS ON ADMISSION|PRIMARY DIAGNOSIS ON ADMISSION
42347-5|T077|strict|42347-5|LNC|PRINCIPLE ADMISSION DIAGNOSIS|PRINCIPLE ADMISSION DIAGNOSIS
42347-5|T077|strict|42347-5|LNC|ADDITIONAL ADMITTING DIAGNOSIS|ADDITIONAL ADMITTING DIAGNOSIS
42347-5|T077|strict|42347-5|LNC|PRELIMINARY DIAGNOSIS|PRELIMINARY DIAGNOSIS
78375-3|T077|strict|78375-3|LNC|DISCHARGE DIAGNOSIS|DISCHARGE DIAGNOSIS
78375-3|T077|strict|78375-3|LNC|PRINCIPLE DISCHARGE DIAGNOSIS|PRINCIPLE DISCHARGE DIAGNOSIS
78375-3|T077|strict|78375-3|LNC|DISCHARGE DIAGNOSES|DISCHARGE DIAGNOSES
78375-3|T077|strict|78375-3|LNC|ASSOCIATE DISCHARGE DIAGNOSIS|ASSOCIATE DISCHARGE DIAGNOSIS
78375-3|T077|strict|78375-3|LNC|PRINCIPAL DIAGNOSIS ON DISCHARGE|PRINCIPAL DIAGNOSIS ON DISCHARGE
78375-3|T077|strict|78375-3|LNC|PRINCIPAL DIAGNOSIS ON THIS PATIENT|PRINCIPAL DIAGNOSIS ON THIS PATIENT
78375-3|T077|strict|78375-3|LNC|PRIMARY DISCHARGE DIAGNOSIS|PRIMARY DISCHARGE DIAGNOSIS
78375-3|T077|strict|78375-3|LNC|PRINCIPAL DISCHARGE DIAGNOSIS|PRINCIPAL DISCHARGE DIAGNOSIS
78375-3|T077|strict|78375-3|LNC|PRINCIPAL DISCHARGE DIAGNOSES|PRINCIPAL DISCHARGE DIAGNOSES
78375-3|T077|strict|78375-3|LNC|DIAGNOSIS AT DISCHARGE|DIAGNOSIS AT DISCHARGE
78375-3|T077|strict|78375-3|LNC|ASSOCIATED DISCHARGE DIAGNOSES|ASSOCIATED DISCHARGE DIAGNOSES
78375-3|T077|strict|78375-3|LNC|OTHER DIAGNOSES ON DISCHARGE|OTHER DIAGNOSES ON DISCHARGE
78375-3|T077|strict|78375-3|LNC|OTHER DIAGNOSIS AT DISCHARGE|OTHER DIAGNOSIS AT DISCHARGE
78375-3|T077|strict|78375-3|LNC|OTHER DISCHARGE DIAGNOSES|OTHER DISCHARGE DIAGNOSES
78375-3|T077|strict|78375-3|LNC|OTHER MEDICAL DIAGNOSIS|OTHER MEDICAL DIAGNOSIS
78375-3|T077|strict|78375-3|LNC|SECONDARY DISCHARGE DIAGNOSES|SECONDARY DISCHARGE DIAGNOSES
78375-3|T077|strict|78375-3|LNC|OTHER DIAGNOSES AND CONDITIONS AFFECTING TREATMENT OR STAY|OTHER DIAGNOSES AND CONDITIONS AFFECTING TREATMENT OR STAY
78375-3|T077|strict|78375-3|LNC|CONDITION AT DISCHARGE|CONDITION AT DISCHARGE
52534-5|T077|strict|52534-5|LNC|PRINCIPAL DIAGNOSIS|PRINCIPAL DIAGNOSIS
52534-5|T077|strict|52534-5|LNC|PRINCIPLE DIAGNOSIS|PRINCIPLE DIAGNOSIS
52534-5|T077|strict|52534-5|LNC|PRIMARY DIAGNOSIS|PRIMARY DIAGNOSIS
52534-5|T077|strict|52534-5|LNC|PRIMARY DX|PRIMARY DX
52534-5|T077|strict|52534-5|LNC|PRIMARY DIAGNOSES|PRIMARY DIAGNOSES
52534-5|T077|strict|52534-5|LNC|PRIMARY MEDICAL DIAGNOSIS|PRIMARY MEDICAL DIAGNOSIS
52534-5|T077|strict|52534-5|LNC|CURRENT DIAGNOSIS|CURRENT DIAGNOSIS
54531-9|T077|strict|54531-9|LNC|ACTIVE DISEASE DIAGNOSIS|ACTIVE DISEASE DIAGNOSIS
54531-9|T077|strict|54531-9|LNC|ACTIVE DISEASE DIAGNOSES|ACTIVE DISEASE DIAGNOSES
54531-9|T077|strict|54531-9|LNC|ACTIVE DIAGNOSES|ACTIVE DIAGNOSES
54531-9|T077|strict|54531-9|LNC|ACUTE DIAGNOSES|ACUTE DIAGNOSES
54531-9|T077|strict|54531-9|LNC|CHRONIC DIAGNOSES|CHRONIC DIAGNOSES
54531-9|T077|strict|54531-9|LNC|HOME CARE DIAGNOSIS|HOME CARE DIAGNOSIS
54531-9|T077|strict|54531-9|LNC|CLINICAL DIAGNOSIS|CLINICAL DIAGNOSIS
54531-9|T077|strict|54531-9|LNC|ACTIVE DIAGNOSIS|ACTIVE DIAGNOSIS
54545-9|T077|strict|54545-9|LNC|ADDITIONAL DIAGNOSES|ADDITIONAL DIAGNOSES
54545-9|T077|strict|54545-9|LNC|SECONDARY DIAGNOSIS|SECONDARY DIAGNOSIS
54545-9|T077|strict|54545-9|LNC|SECONDARY DIAGNOSES|SECONDARY DIAGNOSES
54545-9|T077|strict|54545-9|LNC|RELATED DIAGNOSES|RELATED DIAGNOSES
54545-9|T077|strict|54545-9|LNC|LIST OF OTHER DIAGNOSES|LIST OF OTHER DIAGNOSES
54545-9|T077|strict|54545-9|LNC|LIST OF OTHER PROBLEMS AND DIAGNOSES|LIST OF OTHER PROBLEMS AND DIAGNOSES
54545-9|T077|strict|54545-9|LNC|LIST OF PROBLEMS AND OTHER DIAGNOSES|LIST OF PROBLEMS AND OTHER DIAGNOSES
54545-9|T077|strict|54545-9|LNC|LISTS OF PROBLEMS AND DIAGNOSES|LISTS OF PROBLEMS AND DIAGNOSES
54545-9|T077|strict|54545-9|LNC|OTHER SIGNIFICANT DIAGNOSES|OTHER SIGNIFICANT DIAGNOSES
54545-9|T077|strict|54545-9|LNC|OTHER MEDICAL DIAGNOSIS|OTHER MEDICAL DIAGNOSIS
54545-9|T077|strict|54545-9|LNC|OTHER MEDICAL DIAGNOSES|OTHER MEDICAL DIAGNOSES
54545-9|T077|strict|54545-9|LNC|OTHER PROBLEMS AND DIAGNOSES|OTHER PROBLEMS AND DIAGNOSES
54545-9|T077|strict|54545-9|LNC|OTHER PROBLEMS AND DIAGNOSIS|OTHER PROBLEMS AND DIAGNOSIS
54545-9|T077|strict|54545-9|LNC|OTHER DIAGNOSES|OTHER DIAGNOSES
54545-9|T077|strict|54545-9|LNC|OTHER DIAGNOSIS|OTHER DIAGNOSIS
54545-9|T077|strict|54545-9|LNC|ADDITIONAL DIAGNOSES|ADDITIONAL DIAGNOSES
54545-9|T077|strict|54545-9|LNC|ADDITIONAL DIAGNOSIS|ADDITIONAL DIAGNOSIS
54545-9|T077|strict|54545-9|LNC|ASSOCIATED DIAGNOSES|ASSOCIATED DIAGNOSES
54545-9|T077|strict|54545-9|LNC|ASSOCIATED DIAGNOSIS|ASSOCIATED DIAGNOSIS
29308-4|T077|strict|29308-4|LNC|DIAGNOSIS|DIAGNOSIS
29308-4|T077|strict|29308-4|LNC|DIAGNOSES|DIAGNOSES
29308-4|T077|strict|29308-4|LNC|DIAGNOSES|DIAGNOSES
29308-4|T077|strict|29308-4|LNC|CONDITION|CONDITION
29308-4|T077|strict|29308-4|LNC|VISIT DIAGNOSIS|VISIT DIAGNOSIS
29308-4|T077|strict|29308-4|LNC|VISIT DIAGNOSES|VISIT DIAGNOSES
29308-4|T077|strict|29308-4|LNC|ENCOUNTER DIAGNOSIS|ENCOUNTER DIAGNOSIS
29308-4|T077|strict|29308-4|LNC|ENCOUNTER DIAGNOSES|ENCOUNTER DIAGNOSES
29308-4|T077|strict|29308-4|LNC|DIAGNOSIS LIST|DIAGNOSIS LIST
29308-4|T077|strict|29308-4|LNC|DIAGNOSES LIST|DIAGNOSES LIST
29308-4|T077|strict|29308-4|LNC|LIST OF PROBLEMS AND DIAGNOSES|LIST OF PROBLEMS AND DIAGNOSES
29308-4|T077|strict|29308-4|LNC|LIST OF DIAGNOSES|LIST OF DIAGNOSES
29308-4|T077|strict|29308-4|LNC|PROBLEMS AND DIAGNOSIS|PROBLEMS AND DIAGNOSIS
29308-4|T077|strict|29308-4|LNC|ADDITIONAL DIAGNOSES INCLUDE|ADDITIONAL DIAGNOSES INCLUDE
55110-1|T077|multi|55110-1|LNC|CONCLUSIONS DOCUMENT|CONCLUSIONS DOCUMENT
55110-1|T077|multi|55110-1|LNC|INTERPRETATION DOCUMENT|INTERPRETATION DOCUMENT
55110-1|T077|multi|55110-1|LNC|CONCLUSIONS INTERPRETATION|CONCLUSIONS INTERPRETATION
55110-1|T077|multi|55110-1|LNC|DIAGNOSTIC IMPRESSION|DIAGNOSTIC IMPRESSION
55110-1|T077|multi|55110-1|LNC|INTERPRETATION|INTERPRETATION
55110-1|T077|multi|55110-1|LNC|CONCLUSION|CONCLUSION
55110-1|T077|multi|55110-1|LNC|CONCLUSIONS|CONCLUSIONS
11348-0|T077|strict|11348-0|LNC|PAST MEDICAL HISTORY|PAST MEDICAL HISTORY
11348-0|T077|strict|11348-0|LNC|PMH|PMH
11348-0|T077|strict|11348-0|LNC|PMHX|PMHX
11348-0|T077|strict|11348-0|LNC|CLINICAL HISTORY|CLINICAL HISTORY
11348-0|T077|strict|11348-0|LNC|PERSONAL HISTORY|PERSONAL HISTORY
11348-0|T077|strict|11348-0|LNC|PAST HISTORY|PAST HISTORY
11348-0|T077|strict|11348-0|LNC|HISTORY OF PAST ILLNESS|HISTORY OF PAST ILLNESS
11348-0|T077|strict|11348-0|LNC|PAST GYN HISTORY|PAST GYN HISTORY
11348-0|T077|strict|11348-0|LNC|PAST GYNECOLOGIC HISTORY|PAST GYNECOLOGIC HISTORY
11348-0|T077|strict|11348-0|LNC|PAST PSYCHIATRIC HISTORY|PAST PSYCHIATRIC HISTORY
11348-0|T077|multi|11348-0|LNC|PSYCHIATRIC|PSYCHIATRIC
10219-4|T077|strict|10219-4|LNC|SURGICAL OPERATION NOTE PREOPERATIVE DIAGNOSIS|SURGICAL OPERATION NOTE PREOPERATIVE DIAGNOSIS
10219-4|T077|strict|10219-4|LNC|SURGICAL OPERATION NOTE PREOPERATIVE DX|SURGICAL OPERATION NOTE PREOPERATIVE DX
10219-4|T077|strict|10219-4|LNC|PREOPERATIVE DX|PREOPERATIVE DX
10219-4|T077|strict|10219-4|LNC|OPERATIVE NOTE PRE-OP DX|OPERATIVE NOTE PRE-OP DX
10219-4|T077|strict|10219-4|LNC|PREOPERATIVE DIAGNOSES|PREOPERATIVE DIAGNOSES
10219-4|T077|strict|10219-4|LNC|PREOPERATIVE DIAGNOSIS|PREOPERATIVE DIAGNOSIS
10218-6|T077|strict|10218-6|LNC|SURGICAL OPERATION NOTE POSTOPERATIVE DIAGNOSIS|SURGICAL OPERATION NOTE POSTOPERATIVE DIAGNOSIS
10218-6|T077|multi|10218-6|LNC|POSTPROCEDURE DIAGNOSIS|POSTPROCEDURE DIAGNOSIS
10218-6|T077|strict|10218-6|LNC|POSTOPERATIVE DIAGNOSES|POSTOPERATIVE DIAGNOSES
10218-6|T077|strict|10218-6|LNC|POSTOPERATIVE DIAGNOSIS|POSTOPERATIVE DIAGNOSIS
93127-9|T077|strict|93127-9|LNC|RISK ADJUSTMENT FACTOR|RISK ADJUSTMENT FACTOR
93127-9|T077|strict|93127-9|LNC|RISK SCORE|RISK SCORE
93127-9|T077|strict|93127-9|LNC|RISK ADJUSTMENT|RISK ADJUSTMENT
93127-9|T077|strict|93127-9|LNC|RISK FACTOR|RISK FACTOR
93127-9|T077|strict|93127-9|LNC|RISK|RISK
93127-9|T077|multi|93127-9|LNC|DRG|DRG
93127-9|T077|multi|93127-9|LNC|HCC|HCC
93127-9|T077|multi|93127-9|LNC|HCC/CMS|HCC/CMS
22637-3|T077|strict|22637-3|LNC|PATHOLOGY REPORT FINAL DIAGNOSIS|PATHOLOGY REPORT FINAL DIAGNOSIS
22637-3|T077|strict|22637-3|LNC|HISTOPATHOLOGICAL DIAGNOSIS|HISTOPATHOLOGICAL DIAGNOSIS
22637-3|T077|strict|22637-3|LNC|PATHOLOGIC DIAGNOSIS|PATHOLOGIC DIAGNOSIS
22637-3|T077|multi|22637-3|LNC|FINAL DIAGNOSES|FINAL DIAGNOSES
22637-3|T077|multi|22637-3|LNC|FINAL DIAGNOSIS|FINAL DIAGNOSIS
52797-8|T077|multi|52797-8|LNC|ICD-10-CM|ICD-10-CM
52797-8|T077|multi|52797-8|LNC|ICD-9-CM|ICD-9-CM
52797-8|T077|multi|52797-8|LNC|ICD-10|ICD-10
52797-8|T077|multi|52797-8|LNC|ICD-9|ICD-9
52797-8|T077|multi|52797-8|LNC|ICD10|ICD10
52797-8|T077|multi|52797-8|LNC|ICD9|ICD9
47519-4|T077|strict|47519-4|LNC|HISTORY OF PROCEDURES|HISTORY OF PROCEDURES
47519-4|T077|strict|47519-4|LNC|PROCEDURES HX DOC|PROCEDURES HX DOC
47519-4|T077|strict|47519-4|LNC|PROCEDURES HX|PROCEDURES HX
47519-4|T077|strict|47519-4|LNC|PROCEDURE LIST|PROCEDURE LIST
47519-4|T077|strict|47519-4|LNC|PROCEDURES|PROCEDURES
59772-4|T077|strict|59772-4|LNC|PLANNED PROCEDURE|PLANNED PROCEDURE
55114-3|T077|strict|55114-3|LNC|PRIOR PROCEDURE DESCRIPTIONS|PRIOR PROCEDURE DESCRIPTIONS
55114-3|T077|strict|55114-3|LNC|PRIOR PROCEDURE HISTORY|PRIOR PROCEDURE HISTORY
55114-3|T077|strict|55114-3|LNC|PROCEDURE HISTORY|PROCEDURE HISTORY
55114-3|T077|strict|55114-3|LNC|PROCEDURES HISTORY|PROCEDURES HISTORY
29554-3|T077|multi|29554-3|LNC|PROCEDURE NARRATIVE|PROCEDURE NARRATIVE
29554-3|T077|multi|29554-3|LNC|PRINCIPAL PROCEDURE|PRINCIPAL PROCEDURE
29554-3|T077|multi|29554-3|LNC|PROCEDURE DESCRIPTION|PROCEDURE DESCRIPTION
29554-3|T077|multi|29554-3|LNC|TITLE OF OPERATION|TITLE OF OPERATION
29554-3|T077|multi|29554-3|LNC|PROCEDURES AND SURGICAL/MEDICAL HISTORY|PROCEDURES AND SURGICAL/MEDICAL HISTORY
29554-3|T077|multi|29554-3|LNC|PROCEDURE|PROCEDURE
59773-2|T077|strict|59773-2|LNC|PROCEDURE SPECIMENS TAKEN|PROCEDURE SPECIMENS TAKEN
59773-2|T077|strict|59773-2|LNC|SPECIMENS TAKEN|SPECIMENS TAKEN
46062-6|T077|strict|46062-6|LNC|TREATMENTS SET|TREATMENTS SET
46062-6|T077|strict|46062-6|LNC|TREATMENTS|TREATMENTS
46062-6|T077|strict|46062-6|LNC|CURRENT TREATMENT|CURRENT TREATMENT
46062-6|T077|strict|46062-6|LNC|DIALYSIS|DIALYSIS
46062-6|T077|strict|46062-6|LNC|OSTOMY|OSTOMY
46062-6|T077|strict|46062-6|LNC|RADIATION|RADIATION
46062-6|T077|strict|46062-6|LNC|SUCTIONING|SUCTIONING
46062-6|T077|strict|46062-6|LNC|TRACHEOSTOMY|TRACHEOSTOMY
46062-6|T077|strict|46062-6|LNC|STRESS TEST|STRESS TEST
69967-8|T077|strict|69967-8|LNC|PROCEDURE CODE|PROCEDURE CODE
69967-8|T077|strict|69967-8|LNC|PROCEDURE CODES|PROCEDURE CODES
69967-8|T077|strict|69967-8|LNC|ICD PROCEDURES|ICD PROCEDURES
69967-8|T077|multi|69967-8|LNC|ICD|ICD
69967-8|T077|strict|69967-8|LNC|ICD-10-PCS|ICD-10-PCS
69967-8|T077|strict|69967-8|LNC|CPT|CPT
69967-8|T077|strict|69967-8|LNC|CURRENT PROCEDURAL TERMINOLOGY|CURRENT PROCEDURAL TERMINOLOGY
69967-8|T077|strict|69967-8|LNC|HCPCS|HCPCS
69967-8|T077|strict|69967-8|LNC|HEALTHCARE COMMON PROCEDURE CODING SYSTEM|HEALTHCARE COMMON PROCEDURE CODING SYSTEM
70949-3|T077|strict|70949-3|LNC|PATHOLOGY REPORT|PATHOLOGY REPORT
70949-3|T077|strict|70949-3|LNC|FORMATTED PATH REPORT|FORMATTED PATH REPORT
70949-3|T077|strict|70949-3|LNC|SURGICAL PATHOLOGY STUDY|SURGICAL PATHOLOGY STUDY
70949-3|T077|strict|70949-3|LNC|SURGICAL PATHOLOGY CONSULTATION REPORT|SURGICAL PATHOLOGY CONSULTATION REPORT
70949-3|T077|strict|70949-3|LNC|SURGICAL PATHOLOGY CONSULT|SURGICAL PATHOLOGY CONSULT
70949-3|T077|strict|70949-3|LNC|PATHOLOGY SYNOPTIC REPORT|PATHOLOGY SYNOPTIC REPORT
70949-3|T077|strict|70949-3|LNC|PATHOLOGY CONSULT NOTE|PATHOLOGY CONSULT NOTE
70949-3|T077|strict|70949-3|LNC|DEPARTMENT OF CANCER PATHOLOGY|DEPARTMENT OF CANCER PATHOLOGY
70949-3|T077|strict|70949-3|LNC|PATHOLOGY DEPARTMENT|PATHOLOGY DEPARTMENT
70949-3|T077|strict|70949-3|LNC|COPATH CYTOLOGY REPORT|COPATH CYTOLOGY REPORT
70949-3|T077|strict|70949-3|LNC|DEPARTMENT OF PATHOLOGY|DEPARTMENT OF PATHOLOGY
70949-3|T077|strict|70949-3|LNC|PATHOLOGY ADDENDUM|PATHOLOGY ADDENDUM
70949-3|T077|strict|70949-3|LNC|TAMTRON PRINT|TAMTRON PRINT
70949-3|T077|strict|70949-3|LNC|POWERPATH|POWERPATH
70949-3|T077|strict|70949-3|LNC|CYTOLOGY REQUEST|CYTOLOGY REQUEST
70949-3|T077|strict|70949-3|LNC|PATH REPORT|PATH REPORT
70949-3|T077|multi|70949-3|LNC|PATHOLOGY|PATHOLOGY
22635-7|T077|strict|22635-7|LNC|PATHOLOGY REPORT MICROSCOPIC OBSERVATION|PATHOLOGY REPORT MICROSCOPIC OBSERVATION
22635-7|T077|strict|22635-7|LNC|MICROSCOPIC OBSERVATION|MICROSCOPIC OBSERVATION
22635-7|T077|strict|22635-7|LNC|MICROSCOPIC DESCRIPTION|MICROSCOPIC DESCRIPTION
22635-7|T077|strict|22635-7|LNC|MICROSCOPIC EXAMINATION|MICROSCOPIC EXAMINATION
22635-7|T077|strict|22635-7|LNC|MICROSCOPIC|MICROSCOPIC
33732-9|T077|strict|33732-9|LNC|HISTOLOGY GRADE|HISTOLOGY GRADE
33732-9|T077|strict|33732-9|LNC|HISTOLOGIC GRADE|HISTOLOGIC GRADE
33732-9|T077|strict|33732-9|LNC|HISTOLOGIC|HISTOLOGIC
33732-9|T077|strict|33732-9|LNC|HISTOLOGY|HISTOLOGY
21859-4|T077|strict|21859-4|LNC|PRIMARY CANCER SITE|PRIMARY CANCER SITE
21859-4|T077|strict|21859-4|LNC|ANATOMIC SITE|ANATOMIC SITE
21859-4|T077|strict|21859-4|LNC|SITE OF TISSUE|SITE OF TISSUE
21859-4|T077|strict|21859-4|LNC|TISSUE SITE|TISSUE SITE
21859-4|T077|strict|21859-4|LNC|TUMOR LOCATION|TUMOR LOCATION
21859-4|T077|strict|21859-4|LNC|TUMOR SITE|TUMOR SITE
21939-4|T077|strict|21939-4|LNC|SURGICAL MARGINS|SURGICAL MARGINS
21939-4|T077|strict|21939-4|LNC|MARGINS|MARGINS
92833-3|T077|strict|92833-3|LNC|LYMPH NODES|LYMPH NODES
42186-7|T077|strict|42186-7|LNC|SPECIMENS RECEIVED|SPECIMENS RECEIVED
42186-7|T077|strict|42186-7|LNC|RECEIVED SPECIMEN|RECEIVED SPECIMEN
42186-7|T077|strict|42186-7|LNC|SPECIMEN DETAILS|SPECIMEN DETAILS
42186-7|T077|strict|42186-7|LNC|SPECIMEN ID|SPECIMEN ID
42186-7|T077|strict|42186-7|LNC|MATERIAL COLLECTED ON|MATERIAL COLLECTED ON
42186-7|T077|strict|42186-7|LNC|MATERIAL RECEIVED ON|MATERIAL RECEIVED ON
42186-7|T077|strict|42186-7|LNC|MATERIAL RECEIVED|MATERIAL RECEIVED
66746-9|T077|strict|66746-9|LNC|SPECIMEN TYPE|SPECIMEN TYPE
66746-9|T077|strict|66746-9|LNC|SPECIMEN|SPECIMEN
66746-9|T077|strict|66746-9|LNC|SPECIMENS|SPECIMENS
66746-9|T077|strict|66746-9|LNC|SPECIMEN SOURCE|SPECIMEN SOURCE
66746-9|T077|strict|66746-9|LNC|TISSUE SPECIFICATION|TISSUE SPECIFICATION
90041-5|T077|strict|90041-5|LNC|SPECIMEN COLLECTION|SPECIMEN COLLECTION
90041-5|T077|strict|90041-5|LNC|MATERIAL COLLECTED|MATERIAL COLLECTED
90041-5|T077|strict|90041-5|LNC|SPECIMEN SUBMITTED|SPECIMEN SUBMITTED
90041-5|T077|strict|90041-5|LNC|SPECIMENS SUBMITTED|SPECIMENS SUBMITTED
90041-5|T077|strict|90041-5|LNC|TISSUE SUBMITTED|TISSUE SUBMITTED
90041-5|T077|multi|90041-5|LNC|DATE COLLECTED|DATE COLLECTED
90041-5|T077|multi|90041-5|LNC|COLLECTION DATE|COLLECTION DATE
90041-5|T077|multi|90041-5|LNC|DATE RECEIVED|DATE RECEIVED
90041-5|T077|multi|90041-5|LNC|DATE ENTERED|DATE ENTERED
90041-5|T077|multi|90041-5|LNC|DATE REPORTED|DATE REPORTED
67203-0|T077|strict|67203-0|LNC|AJCC CANCER STAGING|AJCC CANCER STAGING
67203-0|T077|strict|67203-0|LNC|AJCC STAGING|AJCC STAGING
67203-0|T077|strict|67203-0|LNC|AJCC CLASSIFICATION|AJCC CLASSIFICATION
67203-0|T077|strict|67203-0|LNC|AJCC|AJCC
75621-3|T077|strict|75621-3|LNC|TNM PATHOLOGIC STAGING|TNM PATHOLOGIC STAGING
75621-3|T077|strict|75621-3|LNC|TNM PATHOLOGIC STAGING AFTER SURGERY PANEL|TNM PATHOLOGIC STAGING AFTER SURGERY PANEL
75621-3|T077|strict|75621-3|LNC|TNM PATHOLOGIC STAGING|TNM PATHOLOGIC STAGING
75621-3|T077|strict|75621-3|LNC|TNM STAGING|TNM STAGING
75621-3|T077|strict|75621-3|LNC|PATHOLOGIC STAGE|PATHOLOGIC STAGE
75621-3|T077|strict|75621-3|LNC|PATHOLOGY STAGE|PATHOLOGY STAGE
75621-3|T077|strict|75621-3|LNC|NOTTINGHAM HISTOLOGIC SCORE|NOTTINGHAM HISTOLOGIC SCORE
75621-3|T077|strict|75621-3|LNC|TNM STAGE|TNM STAGE
75621-3|T077|strict|75621-3|LNC|STAGING|STAGING
51960-3|T077|strict|51960-3|LNC|MOLECULAR RESULTS|MOLECULAR RESULTS
51960-3|T077|strict|51960-3|LNC|BIOMARKER TESTING|BIOMARKER TESTING
51960-3|T077|strict|51960-3|LNC|MUTATION SCREENING|MUTATION SCREENING
51960-3|T077|strict|51960-3|LNC|MUTATIONAL ANALYSIS|MUTATIONAL ANALYSIS
51960-3|T077|strict|51960-3|LNC|MUTATION ANALYSIS PANEL REPORT|MUTATION ANALYSIS PANEL REPORT
51960-3|T077|strict|51960-3|LNC|DNA MARKER RESULTS PANEL|DNA MARKER RESULTS PANEL
51960-3|T077|strict|51960-3|LNC|DNA TESTING RESULT|DNA TESTING RESULT
51960-3|T077|strict|51960-3|LNC|GENOMIC REFERENCE SEQUENCE|GENOMIC REFERENCE SEQUENCE
51960-3|T077|strict|51960-3|LNC|TRANSCRIPT REFERENCE SEQUENCE|TRANSCRIPT REFERENCE SEQUENCE
51960-3|T077|strict|51960-3|LNC|GENETIC VARIATION CLINICAL SIGNIFICANCE|GENETIC VARIATION CLINICAL SIGNIFICANCE
51960-3|T077|strict|51960-3|LNC|GENE SYMBOL|GENE SYMBOL
51960-3|T077|strict|51960-3|LNC|HGNC|HGNC
51960-3|T077|strict|51960-3|LNC|HUGO|HUGO
51960-3|T077|strict|51960-3|LNC|EXON|EXON
51960-3|T077|strict|51960-3|LNC|EXONS|EXONS
51960-3|T077|strict|51960-3|LNC|INTRON|INTRON
51960-3|T077|strict|51960-3|LNC|INTRONS|INTRONS
51960-3|T077|strict|51960-3|LNC|CODON|CODON
51960-3|T077|strict|51960-3|LNC|CODONS|CODONS
51960-3|T077|strict|51960-3|LNC|GENETIC VARIATION|GENETIC VARIATION
51960-3|T077|strict|51960-3|LNC|GENETIC VARIANT|GENETIC VARIANT
51960-3|T077|strict|51960-3|LNC|DNA TEST RESULT|DNA TEST RESULT
51960-3|T077|strict|51960-3|LNC|DNA CHANGE|DNA CHANGE
51960-3|T077|strict|51960-3|LNC|AMINO ACID CHANGE|AMINO ACID CHANGE
51960-3|T077|strict|51960-3|LNC|PHGVS|PHGVS
51960-3|T077|strict|51960-3|LNC|C.HGVS|C.HGVS
51960-3|T077|strict|51960-3|LNC|HGVS|HGVS
33746-9|T077|strict|33746-9|LNC|PATHOLOGIC FINDINGS|PATHOLOGIC FINDINGS
33746-9|T077|strict|33746-9|LNC|ADDITIONAL PATHOLOGIC FINDINGS|ADDITIONAL PATHOLOGIC FINDINGS
22634-0|T077|strict|22634-0|LNC|PATHOLOGY REPORT GROSS OBSERVATION|PATHOLOGY REPORT GROSS OBSERVATION
22634-0|T077|strict|22634-0|LNC|PATHOLOGY REPORT GROSS OBSERVATION|PATHOLOGY REPORT GROSS OBSERVATION
22634-0|T077|strict|22634-0|LNC|PATHOLOGY REPORT GROSS DESCRIPTION|PATHOLOGY REPORT GROSS DESCRIPTION
22634-0|T077|strict|22634-0|LNC|MACROSCOPIC ANATOMIC OBSERVATIONS|MACROSCOPIC ANATOMIC OBSERVATIONS
22634-0|T077|strict|22634-0|LNC|MACROSCOPIC OBSERVATIONS|MACROSCOPIC OBSERVATIONS
22634-0|T077|strict|22634-0|LNC|MACROSCOPIC DESCRIPTIONS|MACROSCOPIC DESCRIPTIONS
22634-0|T077|strict|22634-0|LNC|MACROSCOPIC EXAMINATION|MACROSCOPIC EXAMINATION
22634-0|T077|strict|22634-0|LNC|MACROSCOPY|MACROSCOPY
22634-0|T077|strict|22634-0|LNC|SPECIMEN INFORMATION|SPECIMEN INFORMATION
22634-0|T077|strict|22634-0|LNC|SPECIMEN INFO|SPECIMEN INFO
22634-0|T077|strict|22634-0|LNC|SPECIMEN|SPECIMEN
22634-0|T077|strict|22634-0|LNC|TISSUE|TISSUE
22634-0|T077|strict|22634-0|LNC|TUMOR SIZE|TUMOR SIZE
22634-0|T077|strict|22634-0|LNC|TUMOR EXTENT|TUMOR EXTENT
22634-0|T077|strict|22634-0|LNC|TUMOR|TUMOR
22634-0|T077|strict|22634-0|LNC|GROSS DESCRIPTION TEXT|GROSS DESCRIPTION TEXT
22634-0|T077|strict|22634-0|LNC|GROSS DESCRIPTION TEXT|GROSS DESCRIPTION TEXT
22634-0|T077|strict|22634-0|LNC|GROSS OBSERVATION|GROSS OBSERVATION
22634-0|T077|strict|22634-0|LNC|GROSS TEXT|GROSS TEXT
22634-0|T077|strict|22634-0|LNC|GROSS FINDINGS|GROSS FINDINGS
2638-1|T077|strict|2638-1|LNC|INTERPRETATION|INTERPRETATION
2638-1|T077|strict|2638-1|LNC|RESULTS|RESULTS
2638-1|T077|strict|2638-1|LNC|RESULT|RESULT
2638-1|T077|strict|2638-1|LNC|CONCLUSION|CONCLUSION
2638-1|T077|strict|2638-1|LNC|COMMENTS|COMMENTS
21902-2|T077|strict|21902-2|LNC|STAGE GROUP|STAGE GROUP
21902-2|T077|strict|21902-2|LNC|CLINICAL STAGE|CLINICAL STAGE
21902-2|T077|strict|21902-2|LNC|CANCER STAGE|CANCER STAGE
21902-2|T077|strict|21902-2|LNC|STAGE IVB|STAGE IVB
21902-2|T077|strict|21902-2|LNC|STAGE IVA|STAGE IVA
21902-2|T077|strict|21902-2|LNC|STAGE IV|STAGE IV
21902-2|T077|strict|21902-2|LNC|STAGE IIIC|STAGE IIIC
21902-2|T077|strict|21902-2|LNC|STAGE IIIB|STAGE IIIB
21902-2|T077|strict|21902-2|LNC|STAGE IIIA|STAGE IIIA
21902-2|T077|strict|21902-2|LNC|STAGE III|STAGE III
21902-2|T077|strict|21902-2|LNC|STAGE IIC|STAGE IIC
21902-2|T077|strict|21902-2|LNC|STAGE IIB|STAGE IIB
21902-2|T077|strict|21902-2|LNC|STAGE IIA|STAGE IIA
21902-2|T077|strict|21902-2|LNC|STAGE II|STAGE II
21902-2|T077|strict|21902-2|LNC|STAGE IB|STAGE IB
21902-2|T077|strict|21902-2|LNC|STAGE IA|STAGE IA
21902-2|T077|strict|21902-2|LNC|STAGE I|STAGE I
21902-2|T077|strict|21902-2|LNC|STAGE IVC|STAGE IVC
21902-2|T077|strict|21902-2|LNC|STAGE IS|STAGE IS
21902-2|T077|strict|21902-2|LNC|STAGE IB2|STAGE IB2
21902-2|T077|strict|21902-2|LNC|STAGE IB1|STAGE IB1
21902-2|T077|strict|21902-2|LNC|STAGE IA2|STAGE IA2
21902-2|T077|strict|21902-2|LNC|STAGE IA1|STAGE IA1
21902-2|T077|strict|21902-2|LNC|STAGE 0IS|STAGE 0IS
21902-2|T077|strict|21902-2|LNC|STAGE 0A|STAGE 0A
21902-2|T077|strict|21902-2|LNC|STAGE 0|STAGE 0
21902-2|T077|strict|21902-2|LNC|STAGE IC|STAGE IC
21902-2|T077|strict|21902-2|LNC|STAGE IE|STAGE IE
21902-2|T077|strict|21902-2|LNC|STAGE 2A1|STAGE 2A1
21902-2|T077|strict|21902-2|LNC|STAGE 2A2|STAGE 2A2
21902-2|T077|strict|21902-2|LNC|STAGE IIE|STAGE IIE
21902-2|T077|strict|21902-2|LNC|STAGE IIS|STAGE IIS
21902-2|T077|strict|21902-2|LNC|STAGE 3C1|STAGE 3C1
21902-2|T077|strict|21902-2|LNC|STAGE 3C2|STAGE 3C2
21902-2|T077|strict|21902-2|LNC|STAGE IIIE|STAGE IIIE
21902-2|T077|strict|21902-2|LNC|STAGE IIIS|STAGE IIIS
21902-2|T077|strict|21902-2|LNC|STAGE IVE|STAGE IVE
21902-2|T077|strict|21902-2|LNC|STAGE IVS|STAGE IVS
59774-0|T077|strict|59774-0|LNC|PROCEDURE ANESTHESIA|PROCEDURE ANESTHESIA
59774-0|T077|strict|59774-0|LNC|ANESTHESIA SECTION|ANESTHESIA SECTION
59774-0|T077|strict|59774-0|LNC|PRIMARY ANESTHESIA|PRIMARY ANESTHESIA
59774-0|T077|strict|59774-0|LNC|ANESTHESIA|ANESTHESIA
83321-0|T077|strict|83321-0|LNC|PATHOLOGY REPORT INTRAOPERATIVE OBSERVATION IN SPECIMEN|PATHOLOGY REPORT INTRAOPERATIVE OBSERVATION IN SPECIMEN
83321-0|T077|strict|83321-0|LNC|INTRAOPERATIVE DIAGNOSIS|INTRAOPERATIVE DIAGNOSIS
8724-7|T077|strict|8724-7|LNC|SURGICAL OPERATION NOTE DESCRIPTION|SURGICAL OPERATION NOTE DESCRIPTION
8724-7|T077|strict|8724-7|LNC|DESCRIPTION OF OPERATION|DESCRIPTION OF OPERATION
8724-7|T077|strict|8724-7|LNC|OPERATION DESCRIPTION|OPERATION DESCRIPTION
8724-7|T077|strict|8724-7|LNC|DESCRIPTION OF THE OPERATION|DESCRIPTION OF THE OPERATION
8724-7|T077|strict|8724-7|LNC|TITLE OF OPERATION|TITLE OF OPERATION
8724-7|T077|strict|8724-7|LNC|OPERATION PERFORMED|OPERATION PERFORMED
8724-7|T077|strict|8724-7|LNC|NAME OF OPERATION|NAME OF OPERATION
59770-8|T077|strict|59770-8|LNC|PROCEDURE ESTIMATED BLOOD LOSS |PROCEDURE ESTIMATED BLOOD LOSS 
59770-8|T077|multi|59770-8|LNC|BLOOD LOSS|BLOOD LOSS
59770-8|T077|strict|59770-8|LNC|ESTIMATED BLOOD LOSS|ESTIMATED BLOOD LOSS
8690-0|T077|strict|8690-0|LNC|HISTORY OF SURGICAL PROCEDURES|HISTORY OF SURGICAL PROCEDURES
8690-0|T077|strict|8690-0|LNC|PAST SURGICAL HISTORY|PAST SURGICAL HISTORY
8690-0|T077|strict|8690-0|LNC|SURGICAL HISTORY|SURGICAL HISTORY
8690-0|T077|strict|8690-0|LNC|OPERATIONS|OPERATIONS
8690-0|T077|strict|8690-0|LNC|OPERATIONS PERFORMED|OPERATIONS PERFORMED
8690-0|T077|strict|8690-0|LNC|OPERATION|OPERATION
8690-0|T077|strict|8690-0|LNC|SURGERIES|SURGERIES
11537-8|T077|strict|11537-8|LNC|SURGICAL DRAINS|SURGICAL DRAINS
11537-8|T077|strict|11537-8|LNC|SURGICAL DRAINS NOTE|SURGICAL DRAINS NOTE
59771-6|T077|strict|59771-6|LNC|PROCEDURE IMPLANTS|PROCEDURE IMPLANTS
59771-6|T077|strict|59771-6|LNC|IMPLANTS|IMPLANTS
10216-0|T077|strict|10216-0|LNC|SURGICAL OPERATION NOTE FLUIDS|SURGICAL OPERATION NOTE FLUIDS
10216-0|T077|strict|10216-0|LNC|OPERATIVE NOTE FLUIDS|OPERATIVE NOTE FLUIDS
10223-6|T077|strict|10223-6|LNC|SURGICAL OPERATION NOTE SURGICAL PROCEDURE|SURGICAL OPERATION NOTE SURGICAL PROCEDURE
10223-6|T077|strict|10223-6|LNC|OPERATIVE NOTE SURGICAL|OPERATIVE NOTE SURGICAL
10223-6|T077|strict|10223-6|LNC|SURGICAL PROCEDURE|SURGICAL PROCEDURE
62387-6|T077|strict|62387-6|LNC|INTERVENTIONS|INTERVENTIONS
62387-6|T077|strict|62387-6|LNC|INTERVENTIONS PROVIDED|INTERVENTIONS PROVIDED
46264-8|T077|strict|46264-8|LNC|HISTORY OF MEDICAL DEVICE USE|HISTORY OF MEDICAL DEVICE USE
46264-8|T077|strict|46264-8|LNC|MEDICAL DEVICE|MEDICAL DEVICE
46264-8|T077|strict|46264-8|LNC|MEDICAL DEVICES|MEDICAL DEVICES
45752-3|T077|strict|45752-3|LNC|VENTILATOR OR RESPIRATOR|VENTILATOR OR RESPIRATOR
45752-3|T077|strict|45752-3|LNC|VENTILATOR|VENTILATOR
45752-3|T077|strict|45752-3|LNC|RESPIRATOR|RESPIRATOR
45752-3|T077|multi|45752-3|LNC|VENT|VENT
8653-8|T077|strict|8653-8|LNC|HOSPITAL DISCHARGE INSTRUCTIONS|HOSPITAL DISCHARGE INSTRUCTIONS
8653-8|T077|strict|8653-8|LNC|DISCHARGE INSTRUCTIONS|DISCHARGE INSTRUCTIONS
69730-0|T077|strict|69730-0|LNC|INSTRUCTIONS|INSTRUCTIONS
69730-0|T077|strict|69730-0|LNC|CARE AND RECOMMENDATIONS|CARE AND RECOMMENDATIONS
69730-0|T077|strict|69730-0|LNC|INSTRUCTIONS|INSTRUCTIONS
69730-0|T077|strict|69730-0|LNC|PATIENT EDUCATION|PATIENT EDUCATION
69730-0|T077|multi|69730-0|LNC|EDUCATION|EDUCATION
18776-5|T077|strict|18776-5|LNC|PLAN OF CARE NOTE|PLAN OF CARE NOTE
18776-5|T077|strict|18776-5|LNC|PLAN OF TREATMENT|PLAN OF TREATMENT
18776-5|T077|strict|18776-5|LNC|CARE PLAN|CARE PLAN
18776-5|T077|strict|18776-5|LNC|CARE RECOMMENDATIONS|CARE RECOMMENDATIONS
18776-5|T077|multi|18776-5|LNC|PLAN|PLAN
51847-2|T077|multi|51847-2|LNC|EVALUATION + PLAN|EVALUATION + PLAN
51847-2|T077|multi|51847-2|LNC|EVALUATION+PLAN|EVALUATION+PLAN
51847-2|T077|multi|51847-2|LNC|EVALUATION AND PLAN|EVALUATION AND PLAN
51847-2|T077|multi|51847-2|LNC|ASSESSMENT AND PLAN|ASSESSMENT AND PLAN
51847-2|T077|multi|51847-2|LNC|ASSESSMENT & PLAN|ASSESSMENT & PLAN
51847-2|T077|multi|51847-2|LNC|ASSESSMENT/PLAN|ASSESSMENT/PLAN
51847-2|T077|multi|51847-2|LNC|IMPRESSION AND PLAN|IMPRESSION AND PLAN
51847-2|T077|multi|51847-2|LNC|A+P|A+P
51847-2|T077|multi|51847-2|LNC|A&P|A&P
61144-2|T077|strict|61144-2|LNC|DIET AND NUTRITION|DIET AND NUTRITION
61144-2|T077|strict|61144-2|LNC|DIET+NUTRITION|DIET+NUTRITION
61144-2|T077|strict|61144-2|LNC|DIET|DIET
61144-2|T077|strict|61144-2|LNC|NUTRITION|NUTRITION
42344-2|T077|strict|42344-2|LNC|DISCHARGE DIET|DISCHARGE DIET
42348-3|T077|strict|42348-3|LNC|ADVANCED DIRECTIVES|ADVANCED DIRECTIVES
42348-3|T077|strict|42348-3|LNC|ADVANCE DIRECTIVES|ADVANCE DIRECTIVES
42348-3|T077|strict|42348-3|LNC|DIRECTIVES|DIRECTIVES
45474-4|T077|strict|45474-4|LNC|ADVANCE DIRECTIVE - DO NOT RESUSCITATE|ADVANCE DIRECTIVE - DO NOT RESUSCITATE
45474-4|T077|strict|45474-4|LNC|DO NOT RESUSCITATE|DO NOT RESUSCITATE
45474-4|T077|strict|45474-4|LNC|DNR|DNR
64289-2|T077|strict|64289-2|LNC|FAX COVER SHEET|FAX COVER SHEET
64289-2|T077|strict|64289-2|LNC|COVER SHEET|COVER SHEET
64289-2|T077|strict|64289-2|LNC|COVER PAGE|COVER PAGE
64289-2|T077|strict|64289-2|LNC|MEDICAL RECORDS REQUEST|MEDICAL RECORDS REQUEST
64289-2|T077|strict|64289-2|LNC|RECORD PULL LIST|RECORD PULL LIST
71727-2|T077|strict|71727-2|LNC|FAX NUMBER|FAX NUMBER
71727-2|T077|strict|71727-2|LNC|FAX|FAX
71727-2|T077|strict|71727-2|LNC|EFAX|EFAX
71727-2|T077|strict|71727-2|LNC|E-FAX|E-FAX
71727-2|T077|strict|71727-2|LNC|SECURE FAX|SECURE FAX
71727-2|T077|strict|71727-2|LNC|HEALTHPORT|HEALTHPORT
71727-2|T077|strict|71727-2|LNC|HEALTH PORT|HEALTH PORT
71727-2|T077|strict|71727-2|LNC|FACESHEET|FACESHEET
71727-2|T077|strict|71727-2|LNC|FACSIMILE TRANSMITTAL SHEET|FACSIMILE TRANSMITTAL SHEET
71727-2|T077|strict|71727-2|LNC|FAX FROM|FAX FROM
71727-2|T077|strict|71727-2|LNC|FAX TO|FAX TO
71727-2|T077|strict|71727-2|LNC|FAX #|FAX #
71727-2|T077|strict|71727-2|LNC|FAXPHONE|FAXPHONE
19826-7|T077|strict|19826-7|LNC|INFORMED CONSENT OBTAINED|INFORMED CONSENT OBTAINED
19826-7|T077|strict|19826-7|LNC|INSTITUTIONAL REVIEW BOARD|INSTITUTIONAL REVIEW BOARD
19826-7|T077|strict|19826-7|LNC|IRB|IRB
19826-7|T077|strict|19826-7|LNC|IRB APPROVAL|IRB APPROVAL
19826-7|T077|strict|19826-7|LNC|IRB APPROVALS|IRB APPROVALS
19826-7|T077|strict|19826-7|LNC|IRB APPROVED|IRB APPROVED
19826-7|T077|strict|19826-7|LNC|WIRB|WIRB
19826-7|T077|strict|19826-7|LNC|WESTERN IRB|WESTERN IRB
19826-7|T077|strict|19826-7|LNC|EXEMPTION REQUEST|EXEMPTION REQUEST
19826-7|T077|strict|19826-7|LNC|INFORMED CONSENT|INFORMED CONSENT
19826-7|T077|strict|19826-7|LNC|PATIENT CONSENT|PATIENT CONSENT
19826-7|T077|strict|19826-7|LNC|CONSENT|CONSENT
55277-8|T077|multi|55277-8|LNC|HIV STATUS|HIV STATUS
55277-8|T077|multi|55277-8|LNC|HIV|HIV
55277-8|T077|multi|55277-8|LNC|HUMAN IMMUNODEFICIENCY VIRUS|HUMAN IMMUNODEFICIENCY VIRUS
76469-6|T077|strict|76469-6|LNC|FEDERAL AGENCY|FEDERAL AGENCY
76469-6|T077|strict|76469-6|LNC|CDC|CDC
76469-6|T077|strict|76469-6|LNC|CENTERS FOR DISEASE CONTROL|CENTERS FOR DISEASE CONTROL
76469-6|T077|strict|76469-6|LNC|DPH|DPH
76469-6|T077|strict|76469-6|LNC|DEPARTMENT OF PUBLIC HEALTH|DEPARTMENT OF PUBLIC HEALTH
76469-6|T077|strict|76469-6|LNC|FDA|FDA
76469-6|T077|strict|76469-6|LNC|FEDERAL DRUG ADMINISTRATION|FEDERAL DRUG ADMINISTRATION
76469-6|T077|strict|76469-6|LNC|SSA|SSA
76469-6|T077|strict|76469-6|LNC|SOCIAL SECURITY ADMINISTRATION|SOCIAL SECURITY ADMINISTRATION
76469-6|T077|strict|76469-6|LNC|SSA-827|SSA-827
76469-6|T077|strict|76469-6|LNC|DISABILITY DETERMINATION|DISABILITY DETERMINATION
76469-6|T077|strict|76469-6|LNC|HIPAA|HIPAA
76469-6|T077|strict|76469-6|LNC|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT|HEALTH INSURANCE PORTABILITY AND ACCOUNTABILITY ACT
76469-6|T077|strict|76469-6|LNC|45 CFR|45 CFR
76469-6|T077|strict|76469-6|LNC|45CFR|45CFR
94137-7|T077|strict|94137-7|LNC|STARS AND HEDIS MEASURE GUIDELINES AND CHECKLIST|STARS AND HEDIS MEASURE GUIDELINES AND CHECKLIST
94137-7|T077|strict|94137-7|LNC|STARS AND HEDIS® MEASURE GUIDELINES AND CHECKLIST|STARS AND HEDIS® MEASURE GUIDELINES AND CHECKLIST
94137-7|T077|strict|94137-7|LNC|HEDIS®|HEDIS®
94137-7|T077|strict|94137-7|LNC|HEDIS|HEDIS
94137-7|T077|strict|94137-7|LNC|HEDIS MEASURE GUIDELINES AND CHECKLIST|HEDIS MEASURE GUIDELINES AND CHECKLIST
94137-7|T077|strict|94137-7|LNC|HEDIS GUIDELINES|HEDIS GUIDELINES
94137-7|T077|strict|94137-7|LNC|HEDIS MEASURE|HEDIS MEASURE
94137-7|T077|strict|94137-7|LNC|HEDIS MEASURES|HEDIS MEASURES