C0011849|T047|73211009|SNOMEDCT_US|DIABETES MELLITUS|DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|ACIDOSES, DIABETIC|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC ACIDOSES|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC KETOACIDOSES|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC KETOACIDOSIS|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|KETOACIDOSES, DIABETIC|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|KETOSIS, DIABETIC|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC ACIDOSIS|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETES MELLITUS WITH KETOACIDOSIS|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|KETOACIDOSIS IN DIABETES MELLITUS |KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|KETOACIDOSIS IN DIABETES MELLITUS|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETES WITH KETOACIDOSIS|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETES MELLITUS WITH KETOACIDOSIS |KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|ACIDOSIS, DIABETIC|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC KETOSIS|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|KETOACIDOSIS, DIABETIC|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC KETOACIDOSIS [DISEASE/FINDING]|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETES MELLITUS NOS WITH KETOACIDOSIS |KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|KETOACIDOSIS - DIABETIC|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETES MELLITUS NOS WITH KETOACIDOSIS|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETES MELLITUS (& [KETOACIDOSIS]) |KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETES MELLITUS (& [KETOACIDOSIS])|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETES WITH KETOACIDOSIS |KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DKA - DIABETIC KETOACIDOSIS|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DKA|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|KETOACIDOSIS (DIABETIC)|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|ACIDOSIS DIABETIC|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC ACIDOSIS WITHOUT COMA|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC KETOSIS WITHOUT COMA|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC ACIDOSIS, NOS|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|DIABETIC KETOSES|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011880|T047|420422005|SNOMEDCT_US|KETOSES, DIABETIC|KETOACIDOSIS IN DIABETES MELLITUS (DISORDER)
C0011875|T047||SNOMEDCT_US|ANGIOPATHIES, DIABETIC
C0011875|T047||SNOMEDCT_US|DIABETIC ANGIOPATHIES
C0011875|T047||SNOMEDCT_US|ANGIOPATHY, DIABETIC
C0011875|T047||SNOMEDCT_US|DIABETIC ANGIOPATHY
C0011875|T047||SNOMEDCT_US|DIABETIC ANGIOPATHIES [DISEASE/FINDING]
C0011875|T047||SNOMEDCT_US|DIABETIC VASCULAR DISEASES
C0011875|T047||SNOMEDCT_US|DIABETIC VASCULAR COMPLICATIONS
C0011875|T047||SNOMEDCT_US|DIABETIC VASCULAR DISORDER
C0011875|T047||SNOMEDCT_US|DIABETIC VASCULAR DISORDER NOS
C0011875|T047||SNOMEDCT_US|DIABETES; ANGIOPATHY (MANIFESTATION)
C0011875|T047||SNOMEDCT_US|ANGIOPATHY; DIABETES (MANIFESTATION)
C0011875|T047||SNOMEDCT_US|DIABETIC VASCULAR COMPLICATION
C0011875|T047||SNOMEDCT_US|DIABETIC VASCULAR DISEASE
C0011875|T047||SNOMEDCT_US|VASCULAR COMPLICATION, DIABETIC
C0011875|T047||SNOMEDCT_US|VASCULAR COMPLICATIONS, DIABETIC
C0011875|T047||SNOMEDCT_US|VASCULAR DISEASE, DIABETIC
C0011875|T047||SNOMEDCT_US|VASCULAR DISEASES, DIABETIC
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC NEPHROPATHIES|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|NEPHROPATHIES, DIABETIC|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETES WITH RENAL MANIFESTATIONS|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|NEPHROPATHY, DIABETIC|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC NEPHROPATHY|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC NEPHROPATHY |RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC KIDNEY DISEASE|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC NEPHROPATHIES [DISEASE/FINDING]|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|NEPHROPATHY;DIABETIC|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETES WITH RENAL MANIFESTATIONS |RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC KIDNEY PROBLEMS|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETES + NEPHROPATHY|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETES WITH RENAL MANIFESTATIONS |RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|NEPHROPATHY - DIABETIC|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|-- DIABETIC KIDNEY DISEASE|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC NEPHROPATHY NOS|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC RENAL DISEASE|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC RENAL DISEASE |RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETES; NEPHROPATHY (MANIFESTATION)|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|NEPHROPATHY; DIABETES (MANIFESTATION)|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|DIABETIC KIDNEY DISEASES|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|KIDNEY DISEASE, DIABETIC|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011881|T047|127013003|SNOMEDCT_US|KIDNEY DISEASES, DIABETIC|RENAL DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHIES|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHIES, DIABETIC|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES WITH NEUROLOGICAL MANIFESTATIONS|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHY|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHY, DIABETIC|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHIES [DISEASE/FINDING]|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHY;DIABETIC|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHY - DIABETIC|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES + NEUROPATHY|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHY |DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES MELLITUS WITH NEUROPATHY|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES MELLITUS NOS WITH NEUROLOGICAL MANIFESTATION |DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETES MELLITUS NOS WITH NEUROLOGICAL MANIFESTATION|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|NEUROPATHY; DIABETES (MANIFESTATION)|DIABETIC NEUROPATHY (DISORDER)
C0011882|T047|230572002|SNOMEDCT_US|DIABETIC NEUROPATHY  [AMBIGUOUS]|DIABETIC NEUROPATHY (DISORDER)
C0085207|T047|11687002|SNOMEDCT_US|DIABETES, GESTATIONAL|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES, PREGNANCY INDUCED|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|GESTATIONAL DIABETES MELLITUS|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|PREGNANCY-INDUCED DIABETES|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|GDM|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES MELLITUS ARISING IN PREGNANCY|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|GESTATIONAL DIABETES|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES IN PREGNANCY|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES PREGN IND|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|GESTATIONAL DIABETES MELLITUS |MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|GESTATIONAL DIABETES MELLITUS NOS|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES, PREGNANCY-INDUCED|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES, GESTATIONAL [DISEASE/FINDING]|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES MELLITUS, GESTATIONAL|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES;DURING PREGNANCY|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES AND PREGNANCY|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|GESTATIONAL DIABETES MELLITUS |MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|MATERNAL GESTATIONAL DIABETES MELLITUS|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|MATERNAL GESTATIONAL DIABETES MELLITUS |MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|-- GESTATIONAL DIABETES|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|MATERNAL DIABETES|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|DIABETES MELLITUS GESTATIONAL|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|GDM - GESTATIONAL DIABETES MELLITUS|MATERNAL GESTATIONAL DIABETES MELLITUS
C0085207|T047|11687002|SNOMEDCT_US|GESTATIONAL DIABETES MELLITUS, NOS|MATERNAL GESTATIONAL DIABETES MELLITUS
C0011854|T047|190362004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, INSULIN-DEPENDENT|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, JUVENILE ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, KETOSIS PRONE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|IDDM|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN-DEPENDENT DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE-ONSET DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KETOSIS-PRONE DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, INSULIN DEPENDENT|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN DEPENDENT DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, SUDDEN ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|MELLITUS, SUDDEN-ONSET DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|SUDDEN-ONSET DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JOD|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|IDDM1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN-DEPENDENT DIABETES MELLITUS 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN-DEPENDENT DIABETES MELLITUS (TYPE I)|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, INSULIN-DEPENDENT, 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS TYPE 01|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN DEPENDENT DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE I DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KETOSIS PRONE DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|IDD|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE 1 DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE 1 DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE I DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, KETOSIS-PRONE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KPD|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|BRITTLE DIABETES (MELLITUS)|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE ONSET DIABETES (MELLITUS)|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KETOSIS-PRONE DIABETES (MELLITUS)|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, TYPE 1 [DISEASE/FINDING]|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, BRITTLE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, JUVENILE-ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, SUDDEN-ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS, TYPE I|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES;TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES;INSULIN DEPENDENT|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES;JUVENILE ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN DEPENDENT DIABETES MELLITUS 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE ONSET DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES, JUVENILE-ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE-ONSET DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN-DEPENDENT DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS: [JUVENILE] OR [INSULIN DEPENDENT]|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS - JUVENILE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS: [JUVENILE] OR [INSULIN DEPENDENT] |TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE ONSET DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE I DIABETES MELLITUS |TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|IDDM - INSULIN-DEPENDENT DIABETES MELLITUS|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN DEPENDENT DIABETES MEL|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|-- DIABETES TYPE 1|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS TYPE I|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE 1 DIABETES MELLITUS |TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS JUVENILE ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS INSULIN-DEPENDENT|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN DEPENDENT DIABETIC|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES MELLITUS TYPE 1 |TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES; INSULIN-DEPENDENT|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES; JUVENILE-ONSET|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES; KETOSIS-PRONE|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|DIABETES; TYPE I|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|INSULIN-DEPENDENT; DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE-ONSET; DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|KETOSIS, PRONE; DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|TYPE I; DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011854|T047|190362004|SNOMEDCT_US|JUVENILE ONSET OF DIABETES|TYPE I DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|ADULT-ONSET DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, ADULT ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, KETOSIS RESISTANT|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, NON-INSULIN-DEPENDENT|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|KETOSIS-RESISTANT DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NIDDM|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NON-INSULIN-DEPENDENT DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|STABLE DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, MATURITY ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|MATURITY ONSET DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NONINSULIN DEPENDENT DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, SLOW ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|SLOW-ONSET DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NONINSULIN-DEPENDENT DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, NONINSULIN-DEPENDENT|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS TYPE 02|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|ADULT ONSET DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|TYPE II DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|KETOSIS RESISTANT DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS NON INSULIN-DEP|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|TYPE 2 DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|AODM|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|TYPE 2 DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NON-INSULIN DEPENDENT DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|ADULT-ONSET DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|TYPE 2 DIABETES MELLITUS NON-INSULIN DEPENDENT|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|TYPE II DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|T2D|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|T2DM - TYPE 2 DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES, TYPE 2|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, STABLE|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|MODY|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, TYPE 2|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, KETOSIS-RESISTANT|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, NON INSULIN DEPENDENT|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, SLOW-ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, NONINSULIN DEPENDENT|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, TYPE 2 [DISEASE/FINDING]|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|MATURITY-ONSET DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, MATURITY-ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, ADULT-ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS, TYPE II|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES;TYPE 2|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES;ADULT ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES;NON INSULIN DEPEND|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS (NIDDM)|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|MATURITY-ONSET DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES TYPE 2|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS TYPE 2|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS - ADULT ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS: [ADULT ONSET] OR [NONINSULIN DEPENDENT]|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS: [ADULT ONSET] OR [NONINSULIN DEPENDENT] |TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS -ADULT ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NIDDM - NON-INSULIN DEPENDENT DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|TYPE II DIABETES MELLITUS |TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|MATURITY ONSET DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NONINSULIN DEPENDENT DIAB.MELL|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NON-INSULIN-DEPENDENT DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|-- DIABETES TYPE 2|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NONINSULIN DEPENDENT DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|TYPE I I DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|ADULT ONSET DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NONINSULIN DEPENDENT DIABETES MELLITUS (NIDDM)|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NONINSULIN-DEPENDENT DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS TYPE II|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NIDDM DIABETES MELLITUS|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|TYPE 2 DIABETES MELLITUS |TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS MATURITY ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS NON-INSULIN-DEPENDENT|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES MELLITUS TYPE 2 |TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NIDDM; DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES; NIDDM|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES; ADULT-ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES; MATURITY-ONSET|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES; NON-INSULIN-DEPENDENT|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES; NONKETOTIC|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|DIABETES; TYPE II|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|MATURITY-ONSET; DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NON-INSULIN-DEPENDENT; DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NONKETOTIC; DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|ADULT-ONSET; DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|TYPE II; DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NCDMM|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NON-INSULIN DEPENDENT DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0011860|T047|190384004|SNOMEDCT_US|NON INSULIN DEPENDENT DIABETES|TYPE II DIABETES MELLITUS (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PREDIABETIC STATE|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PREDIABETIC STATES|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|STATE, PREDIABETIC|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|STATES, PREDIABETIC|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PREDIABETES|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PREDIABETIC STATE [DISEASE/FINDING]|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PRE DIABETES|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PREDIABETES |PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PRE-DIABETIC|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|BORDERLINE DIABETES|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PRE-DIABETES|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PREDIABETES |PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PREDIABETES SYNDROME|PREDIABETES (DISORDER)
C0362046|T047|15777000|SNOMEDCT_US|PRE-DIABETES NOS|PREDIABETES (DISORDER)
C0271646|T047|5368009|SNOMEDCT_US|DRUG RELATED DIABETES MELLITUS|DRUG-INDUCED DIABETES MELLITUS (DISORDER)
C0271646|T047|5368009|SNOMEDCT_US|DRUG-INDUCED DIABETES MELLITUS |DRUG-INDUCED DIABETES MELLITUS (DISORDER)
C0271646|T047|5368009|SNOMEDCT_US|DRUG-INDUCED DIABETES MELLITUS|DRUG-INDUCED DIABETES MELLITUS (DISORDER)
C0597655|T047||SNOMEDCT_US|VIRUS RELATED DIABETES MELLITUS
C0920358|T047||SNOMEDCT_US|DIABETIC OPHTHALMOPATHY
C0853897|T047||SNOMEDCT_US|DIABETIC CARDIOMYOPATHY
C0853897|T047||SNOMEDCT_US|DIABETIC CARDIOMYOPATHIES
C0853897|T047||SNOMEDCT_US|CARDIOMYOPATHY, DIABETIC
C0853897|T047||SNOMEDCT_US|CARDIOMYOPATHIES, DIABETIC
C0853897|T047||SNOMEDCT_US|DIABETIC CARDIOMYOPATHIES [DISEASE/FINDING]
C0348447|T047|191045007|SNOMEDCT_US|OTHER SPECIFIED DIABETES MELLITUS|[X]OTHER SPECIFIED DIABETES MELLITUS (DISORDER)
C0348447|T047|191045007|SNOMEDCT_US|[X]OTHER SPECIFIED DIABETES MELLITUS|[X]OTHER SPECIFIED DIABETES MELLITUS (DISORDER)
C0348447|T047|191045007|SNOMEDCT_US|[X]OTHER SPECIFIED DIABETES MELLITUS |[X]OTHER SPECIFIED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|MALNUTRITION-RELATED DIABETES MELLITUS|MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|DIABETES MELLITUS MALNUTRITION-RELATED|MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|MALNUTRITION-RELATED DIABETES MELLITUS |MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|MALNUTRITION-RELATED DIABETES MELLITUS |MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|DIABETES MELLITUS SECONDARY MALNUTRITION-RELATED|MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|MRDM|MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|MALNUTRITION RELATED DIABETES MELLITUS|MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|MALNUTRITION RELATED DIABETES MELLITUS |MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|DIABETES; MALNUTRITION-RELATED|MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0271641|T047|75524006|SNOMEDCT_US|MALNUTRITION; DIABETES|MALNUTRITION RELATED DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES MELLITUS|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES MELLITUS |DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DM|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES NOS|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES MELLITUS [DISEASE/FINDING]|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES MELLITUS (E08-E13)|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES MELLITUS |DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES MELLITUS NOS|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES MELLLITUS|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|MED: DIABETES MELLITUS|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DM - DIABETES MELLITUS|DIABETES MELLITUS (DISORDER)
C0011849|T047|73211009|SNOMEDCT_US|DIABETES MELLITUS, NOS|DIABETES MELLITUS (DISORDER)
C0348939|T047|190383005|SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH MULTIPLE COMPLICATIONS|UNSPECIFIED DIABETES MELLITUS WITH MULTIPLE COMPLICATIONS (DISORDER)
C0348939|T047|190383005|SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH MULTIPLE COMPLICATIONS |UNSPECIFIED DIABETES MELLITUS WITH MULTIPLE COMPLICATIONS (DISORDER)
C0348450|T047|191048009|SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH RENAL COMPLICATIONS|[X]UNSPECIFIED DIABETES MELLITUS WITH RENAL COMPLICATIONS (DISORDER)
C0348450|T047|191048009|SNOMEDCT_US|[X]UNSPECIFIED DIABETES MELLITUS WITH RENAL COMPLICATIONS |[X]UNSPECIFIED DIABETES MELLITUS WITH RENAL COMPLICATIONS (DISORDER)
C0348450|T047|191048009|SNOMEDCT_US|[X]UNSPECIFIED DIABETES MELLITUS WITH RENAL COMPLICATIONS|[X]UNSPECIFIED DIABETES MELLITUS WITH RENAL COMPLICATIONS (DISORDER)
C0494295|T047||SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH COMA
C0494296|T047||SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH KETOACIDOSIS
C2362567|T047||SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH NEUROLOGICAL COMPLICATIONS
C1744704|T047||SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH OPHTHALMIC COMPLICATIONS
C0494300|T047||SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS
C0011871|T047|982001|SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH PERIPHERAL CIRCULATORY COMPLICATIONS|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETIC PERIPHERAL ANGIOPATHY|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETES MELLITUS WITH PERIPHERAL CIRCULATORY DISORDER|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETES MELLITUS WITH PERIPHERAL CIRCULATORY DISORDER |DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETES WITH PERIPHERAL CIRCULATORY DISORDER|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETES MELLITUS WITH PERIPHERAL CIRCULATORY DISORDER |DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS |DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETES MELLITUS NOS WITH PERIPHERAL CIRCULATORY DISORDER |DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETES MELLITUS NOS WITH PERIPHERAL CIRCULATORY DISORDER|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETES + PERIPH.CIRCULAT.DIS|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETIC PERIPHERAL VASCULAR DISEASE|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETIC PERIPHERAL ANGIOPATHY |DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0011871|T047|982001|SNOMEDCT_US|DIABETIC PERIPHERAL VASCULAR DISORDER|DIABETES WITH PERIPHERAL CIRCULATORY DISORDERS (DISORDER)
C0342257|T047|74627003|SNOMEDCT_US|DISORDER ASSOCIATED WITH DIABETES MELLITUS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITH UNSPECIFIED COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES COMPL|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|COMPL DIABETES MELLITUS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES RELAT COMPL|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETIC COML|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS WITH COMPLICATION |DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS WITH COMPLICATION|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES WITH UNSPECIFIED COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETIC COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS WITH COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES COMPLICATION|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES-RELATED COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES COMPLICATIONS [DISEASE/FINDING]|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|COMPLICATIONS OF DIABETES MELLITUS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES;COMPLICATED|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS NOS WITH UNSPECIFIED COMPLICATION|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS WITH UNSPECIFIED COMPLICATION|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES WITH DIABETIC COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS WITH UNSPECIFIED COMPLICATION |DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS WITH COMPLICATION |DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS NOS WITH UNSPECIFIED COMPLICATION |DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES--COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES WITH UNSPECIFIED COMPLICATION|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETIC COMPLICATION|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETIC COMPLICATION NOS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETIC COMPLICATION |DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETIC COMPLICATION, NOS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES MELLITUS COMPLICATION|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES RELATED COMPLICATIONS|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|DIABETES-RELATED COMPLICATION|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0342257|T047|74627003|SNOMEDCT_US|COMPLICATED DIABETES|DISORDER ASSOCIATED WITH DIABETES MELLITUS
C0271635|T047|111552007|SNOMEDCT_US|DIABETES MELLITUS WITHOUT COMPLICATION|DIABETES MELLITUS WITHOUT COMPLICATION (DISORDER)
C0271635|T047|111552007|SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS WITHOUT COMPLICATIONS|DIABETES MELLITUS WITHOUT COMPLICATION (DISORDER)
C0271635|T047|111552007|SNOMEDCT_US|DIABETES MELLITUS WITHOUT COMPLICATION |DIABETES MELLITUS WITHOUT COMPLICATION (DISORDER)
C0271635|T047|111552007|SNOMEDCT_US|DIABETES MELLITUS NOS WITH NO MENTION OF COMPLICATION|DIABETES MELLITUS WITHOUT COMPLICATION (DISORDER)
C0271635|T047|111552007|SNOMEDCT_US|DIABETES MELLITUS WITH NO MENTION OF COMPLICATION |DIABETES MELLITUS WITHOUT COMPLICATION (DISORDER)
C0271635|T047|111552007|SNOMEDCT_US|DIABETES MELLITUS WITH NO MENTION OF COMPLICATION|DIABETES MELLITUS WITHOUT COMPLICATION (DISORDER)
C0271635|T047|111552007|SNOMEDCT_US|DIABETES MELLITUS NOS WITH NO MENTION OF COMPLICATION |DIABETES MELLITUS WITHOUT COMPLICATION (DISORDER)
C0271635|T047|111552007|SNOMEDCT_US|DIABETES MELLITUS WITHOUT MENTION OF COMPLICATION|DIABETES MELLITUS WITHOUT COMPLICATION (DISORDER)
C0271635|T047|111552007|SNOMEDCT_US|DIABETES MELLITUS WITHOUT COMPLICATION |DIABETES MELLITUS WITHOUT COMPLICATION (DISORDER)
C2711205|T047|441628001|SNOMEDCT_US|MULTIPLE COMPLICATIONS DUE TO DIABETES MELLITUS |MULTIPLE COMPLICATIONS DUE TO DIABETES MELLITUS (DISORDER)
C2711205|T047|441628001|SNOMEDCT_US|MULTIPLE COMPLICATIONS DUE TO DIABETES MELLITUS|MULTIPLE COMPLICATIONS DUE TO DIABETES MELLITUS (DISORDER)
C0265344|T047|111307005|SNOMEDCT_US|DONOHUE SYNDROME}CONGENITAL CONDITION, INSULIN RECEPTOR IMPAIRED|LEPRECHAUNISM SYNDROME (DISORDER)
C0265344|T047|111307005|SNOMEDCT_US|LEPRECHAUNISMS|LEPRECHAUNISM SYNDROME (DISORDER)
C0265344|T047|111307005|SNOMEDCT_US|SYNDROME, DONOHUE|LEPRECHAUNISM SYNDROME (DISORDER)
C0265344|T047|111307005|SNOMEDCT_US|DONOHUE SYNDROME [DISEASE/FINDING]|LEPRECHAUNISM SYNDROME (DISORDER)
C0265344|T047|111307005|SNOMEDCT_US|LEPRECHAUNISM|LEPRECHAUNISM SYNDROME (DISORDER)
C0265344|T047|111307005|SNOMEDCT_US|LEPRECHAUNISM SYNDROME|LEPRECHAUNISM SYNDROME (DISORDER)
C0265344|T047|111307005|SNOMEDCT_US|DONOHUE'S SYNDROME|LEPRECHAUNISM SYNDROME (DISORDER)
C0265344|T047|111307005|SNOMEDCT_US|LEPRECHAUNISM SYNDROME |LEPRECHAUNISM SYNDROME (DISORDER)
C0265344|T047|111307005|SNOMEDCT_US|DONOHUE|LEPRECHAUNISM SYNDROME (DISORDER)
C2827448|T047||SNOMEDCT_US|CHILDHOOD DIABETES MELLITUS
C2873880|T047||SNOMEDCT_US|DIABETES MELLITUS DUE TO UNDERLYING CONDITION
C2873948|T047||SNOMEDCT_US|DRUG OR CHEMICAL INDUCED DIABETES MELLITUS
C2919615|T047|445260006|SNOMEDCT_US|POSTTRANSPLANT DIABETES MELLITUS |POSTTRANSPLANT DIABETES MELLITUS (DISORDER)
C2919615|T047|445260006|SNOMEDCT_US|POSTTRANSPLANT DIABETES MELLITUS|POSTTRANSPLANT DIABETES MELLITUS (DISORDER)
C0554876|T047||SNOMEDCT_US|POORLY CONTROLLED DIABETES MELLITUS 
C0554876|T047||SNOMEDCT_US|DIABETES MELLITUS POORLY CONTROLLED
C0554876|T047||SNOMEDCT_US|POORLY CONTROLLED DIABETES MELLITUS
C1720078|T047|422088007|SNOMEDCT_US|DIABETIC NEUROLOGIC DISEASE|DIABETIC NEUROLOGIC DISEASE
C1720078|T047|422088007|SNOMEDCT_US|NEUROLOGIC COMPLICATION OF DIABETES MELLITUS|DIABETIC NEUROLOGIC DISEASE
C1720078|T047|422088007|SNOMEDCT_US|NEUROLOGIC DISORDER ASSOCIATED WITH DIABETES MELLITUS |DIABETIC NEUROLOGIC DISEASE
C1720078|T047|422088007|SNOMEDCT_US|NEUROLOGIC DISORDER ASSOCIATED WITH DIABETES MELLITUS|DIABETIC NEUROLOGIC DISEASE
C1720078|T047|422088007|SNOMEDCT_US|DIABETES MELLITUS WITH NEUROLOGICAL COMPLICATIONS |DIABETIC NEUROLOGIC DISEASE
C1720078|T047|422088007|SNOMEDCT_US|DIABETES WITH NEUROLOGICAL COMPLICATIONS|DIABETIC NEUROLOGIC DISEASE
C1720078|T047|422088007|SNOMEDCT_US|DIABETES MELLITUS WITH NEUROLOGICAL COMPLICATIONS|DIABETIC NEUROLOGIC DISEASE
C0342245|T047|25093002|SNOMEDCT_US|DIABETES WITH OPHTHALMIC MANIFESTATIONS|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETES MELLITUS WITH OPHTHALMIC MANIFESTATIONS |DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETES MELLITUS WITH OPHTHALMIC MANIFESTATIONS|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETIC EYE DISEASE|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETIC EYE PROBLEMS|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETES MELLITUS NOS WITH OPHTHALMIC MANIFESTATION|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETES MELLITUS WITH OPHTHALMIC MANIFESTATION |DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETES MELLITUS WITH OPHTHALMIC MANIFESTATION|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETES + EYE MANIFESTATION|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETES MELLITUS NOS WITH OPHTHALMIC MANIFESTATION |DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETIC EYE DISEASE NOS|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|OPHTHALMIC MANIFESTATIONS OF DIABETES|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETIC OCULOPATHY |DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETIC OCULOPATHY|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETIC OCULOPATHY, NOS|DIABETIC OCULOPATHY (DISORDER)
C0342245|T047|25093002|SNOMEDCT_US|DIABETIC EYE DISEASE, NOS|DIABETIC OCULOPATHY (DISORDER)
C2062378|T047||SNOMEDCT_US|DIABETES MELLITUS UNDER CONTROL
C2062378|T047||SNOMEDCT_US|DIABETES MELLITUS UNDER CONTROL 
C0553772|T047|310505005|SNOMEDCT_US|DIABETES MELLITUS WITH HYPEROSMOLAR NONKETOTIC STATE |DIABETIC HYPEROSMOLAR NON-KETOTIC STATE (DISORDER)
C0553772|T047|310505005|SNOMEDCT_US|DIABETES MELLITUS WITH HYPEROSMOLAR NONKETOTIC STATE|DIABETIC HYPEROSMOLAR NON-KETOTIC STATE (DISORDER)
C0553772|T047|310505005|SNOMEDCT_US|HYPERGLYCEMIC HYPEROSMOLAR NONKETOTIC STATE|DIABETIC HYPEROSMOLAR NON-KETOTIC STATE (DISORDER)
C0553772|T047|310505005|SNOMEDCT_US|DIABETIC HYPEROSMOLAR NON-KETOTIC STATE|DIABETIC HYPEROSMOLAR NON-KETOTIC STATE (DISORDER)
C0553772|T047|310505005|SNOMEDCT_US|HONKS - DIABETIC HYPEROSMOLAR NON-KETOTIC STATE|DIABETIC HYPEROSMOLAR NON-KETOTIC STATE (DISORDER)
C0553772|T047|310505005|SNOMEDCT_US|DIABETIC HYPEROSMOLAR NON-KETOTIC STATE |DIABETIC HYPEROSMOLAR NON-KETOTIC STATE (DISORDER)
C0860163|T047||SNOMEDCT_US|DIABETIC GASTROPATHY
C0860163|T047||SNOMEDCT_US|DIABETES MELLITUS WITH GASTROPATHY 
C0860163|T047||SNOMEDCT_US|DIABETES MELLITUS WITH GASTROPATHY
C0271640|T047|8801005|SNOMEDCT_US|SECONDARY DIABETES MELLITUS|SECONDARY DIABETES MELLITUS (DISORDER)
C0271640|T047|8801005|SNOMEDCT_US|SECONDARY DIABETES MELLITUS NOS|SECONDARY DIABETES MELLITUS (DISORDER)
C0271640|T047|8801005|SNOMEDCT_US|SECONDARY DIABETES MELLITUS |SECONDARY DIABETES MELLITUS (DISORDER)
C0271640|T047|8801005|SNOMEDCT_US|SECONDARY DIABETES MELLITUS |SECONDARY DIABETES MELLITUS (DISORDER)
C0271640|T047|8801005|SNOMEDCT_US|SECONDARY DIABETES MELLITUS, NOS|SECONDARY DIABETES MELLITUS (DISORDER)
C0158981|T047|49817004|SNOMEDCT_US|NEONATAL DIABETES MELLITUS|NEONATAL DIABETES MELLITUS (DISORDER)
C0158981|T047|49817004|SNOMEDCT_US|NEONATAL DIABETES MELLITUS |NEONATAL DIABETES MELLITUS (DISORDER)
C0158981|T047|49817004|SNOMEDCT_US|NEONATAL DIABETES|NEONATAL DIABETES MELLITUS (DISORDER)
C0158981|T047|49817004|SNOMEDCT_US|NEONAT DIABETES MELLITUS|NEONATAL DIABETES MELLITUS (DISORDER)
C0158981|T047|49817004|SNOMEDCT_US|DIABETES MELLITUS SYNDROME IN NEWBORN INFANT|NEONATAL DIABETES MELLITUS (DISORDER)
C0158981|T047|49817004|SNOMEDCT_US|CONGENITAL DIABETES MELLITUS|NEONATAL DIABETES MELLITUS (DISORDER)
C0158981|T047|49817004|SNOMEDCT_US|NEONATAL DIABETES MELLITUS |NEONATAL DIABETES MELLITUS (DISORDER)
C0158981|T047|49817004|SNOMEDCT_US|DIABETES; NEONATAL|NEONATAL DIABETES MELLITUS (DISORDER)
C0158981|T047|49817004|SNOMEDCT_US|NEONATAL; DIABETES|NEONATAL DIABETES MELLITUS (DISORDER)
C0865166|T047||SNOMEDCT_US|DIABETIC HYPOGLYCEMIA NOS
C0865166|T047||SNOMEDCT_US|DIABETES MELLITUS WITH HYPOGLYCEMIA
C0865166|T047||SNOMEDCT_US|DIABETIC HYPOGLYCEMIA
C0865166|T047||SNOMEDCT_US|DIABETIC HYPOGLYCEMIA 
C2930860|T047||SNOMEDCT_US|PREMATURE AGING, OKAMOTO TYPE
C2931057|T047||SNOMEDCT_US|LIPOATROPHY WITH DIABETES, HEPATIC STEATOSIS, CARDIOMYOPATHY, AND LEUKOMELANODERMIC PAPULES
C2931125|T047|720519003|SNOMEDCT_US|FEIGENBAUM BERGERON RICHARDSON SYNDROME|ATHEROSCLEROSIS, DEAFNESS, DIABETES, EPILEPSY, NEPHROPATHY SYNDROME (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|CHARACTERIZED BY DM ALONG WITH OTHER THINGS|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|THIAMINE-RESPONSIVE MEGALOBLASTIC ANEMIA SYNDROME|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|THIAMINE RESPONSIVE MYELODYSPLASIA|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|THIAMINE RESPONSIVE MEGALOBLASTIC ANEMIA SYNDROME|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|ABBOUD SYNDROME|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|ROGERS SYNDROME|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|THMD1|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|THIAMINE-RESPONSIVE MYELODYSPLASIA|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|THIAMINE-RESPONSIVE ANEMIA SYNDROME|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|THIAMINE METABOLISM DYSFUNCTION SYNDROME 1 (MEGALOBLASTIC ANEMIA, DIABETES MELLITUS, AND DEAFNESS TYPE)|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|MEGALOBLASTIC ANAEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C0342287|T047|237617006|SNOMEDCT_US|MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS |MEGALOBLASTIC ANEMIA, THIAMINE-RESPONSIVE, WITH DIABETES MELLITUS AND SENSORINEURAL DEAFNESS (DISORDER)
C2931296|T047|722206009|SNOMEDCT_US|PANCREATIC HYPOPLASIA DIABETES HEART DISEASE|PANCREATIC HYPOPLASIA, DIABETES MELLITUS, CONGENITAL HEART DISEASE SYNDROME (DISORDER)
C2931296|T047|722206009|SNOMEDCT_US|YORIFUJI OKUNO SYNDROME|PANCREATIC HYPOPLASIA, DIABETES MELLITUS, CONGENITAL HEART DISEASE SYNDROME (DISORDER)
C0342286|T047|237616002|SNOMEDCT_US|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA ,MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES (DISORDER)
C0342286|T047|237616002|SNOMEDCT_US|WOODHOUSE SAKATI SYNDROME|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES (DISORDER)
C0342286|T047|237616002|SNOMEDCT_US|EXTRAPYRAMIDAL DISORDER, PROGRESSIVE, WITH PRIMARY HYPOGONADISM, MENTAL RETARDATION, AND ALOPECIA|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES (DISORDER)
C0342286|T047|237616002|SNOMEDCT_US|HYPOGONADISM, ALOPECIA, DIABETES MELLITUS, MENTAL RETARDATION, AND EXTRAPYRAMIDAL SYNDROME|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES (DISORDER)
C0342286|T047|237616002|SNOMEDCT_US|WOODHOUSE-SAKATI SYNDROME|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES (DISORDER)
C0342286|T047|237616002|SNOMEDCT_US|HYPOGONADISM, ALOPECIA, DIABETES MELLITUS, MENTAL RETARDATION, DEAFNESS, AND EXTRAPYRAMIDAL SYNDROME|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES (DISORDER)
C0342286|T047|237616002|SNOMEDCT_US|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES |HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES (DISORDER)
C0342286|T047|237616002|SNOMEDCT_US|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES (DISORDER)
C0342286|T047|237616002|SNOMEDCT_US|HYPOGONADISM, DIABETES MELLITUS, ALOPECIA ,MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES |HYPOGONADISM, DIABETES MELLITUS, ALOPECIA, MENTAL RETARDATION AND ELECTROCARDIOGRAPHIC ABNORMALITIES (DISORDER)
C1838655|T047||SNOMEDCT_US|PANCREATIC BETA CELL AGENESIS WITH NEONATAL DIABETES MELLITUS
C1838655|T047||SNOMEDCT_US|CONGENITAL ABSENCE OF INSULIN-PRODUCING BETA CELLS WITH DIABETES MELLITUS
C1809475|T047|237612000|SNOMEDCT_US|PHOTOMYOCLONUS, DIABETES MELLITUS, DEAFNESS, NEPHROPATHY, AND CEREBRAL DYSFUNCTION|PHOTOMYOCLONUS, DIABETES MELLITUS, DEAFNESS, NEPHROPATHY AND CEREBRAL DYSFUNCTION (DISORDER)
C1809475|T047|237612000|SNOMEDCT_US|HERRMANN SYNDROME|PHOTOMYOCLONUS, DIABETES MELLITUS, DEAFNESS, NEPHROPATHY AND CEREBRAL DYSFUNCTION (DISORDER)
C1809475|T047|237612000|SNOMEDCT_US|PHOTOMYOCLONUS, DIABETES MELLITUS, DEAFNESS, NEPHROPATHY AND CEREBRAL DYSFUNCTION|PHOTOMYOCLONUS, DIABETES MELLITUS, DEAFNESS, NEPHROPATHY AND CEREBRAL DYSFUNCTION (DISORDER)
C1809475|T047|237612000|SNOMEDCT_US|PHOTOMYOCLONUS, DIABETES MELLITUS, DEAFNESS, NEPHROPATHY AND CEREBRAL DYSFUNCTION |PHOTOMYOCLONUS, DIABETES MELLITUS, DEAFNESS, NEPHROPATHY AND CEREBRAL DYSFUNCTION (DISORDER)
C2931765|T047||SNOMEDCT_US|FURUKAWA TAKAGI NAKAO SYNDROME
C0431693|T047|446641003|SNOMEDCT_US|RENAL CYSTS AND DIABETES SYNDROME|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|MODY5|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|HYPERURICEMIC NEPHROPATHY, FAMILIAL JUVENILE, ATYPICAL|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|GLOMERULOCYSTIC KIDNEY DISEASE, HYPOPLASTIC TYPE|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|GLOMERULOCYSTIC KIDNEY, FAMILIAL HYPOPLASTIC|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG, TYPE 5|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|RENAL CYSTS AND DIABETES SYNDROME |RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG, TYPE 5 |RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|FAMILIAL HYPOPLASTIC, GLOMERULOCYSTIC KIDNEY|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|FAMILIAL HYPOPLASTIC, GLOMERULOCYSTIC KIDNEY |RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|RCAD|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG - TYPE 5 |RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG - TYPE 5|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|FJHN, ATYPICAL|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|CONGENITAL ANOMALIES OF THE KIDNEY AND URINARY TRACT WITH DIABETES|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|CAKUT WITH DIABETES|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|RCAD SYNDROME|RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0431693|T047|446641003|SNOMEDCT_US|FAMILIAL HYPOPLASTIC, GLOMERULOCYSTIC KIDNEY |RENAL CYSTS AND DIABETES SYNDROME (DISORDER)
C0406682|T047|238982009|SNOMEDCT_US|DIABETIC DERMOPATHY|DIABETIC DERMOPATHY (DISORDER)
C0406682|T047|238982009|SNOMEDCT_US|DIABETES MELLITUS WITH DERMATOLOGICAL MANIFESTATIONS|DIABETIC DERMOPATHY (DISORDER)
C0406682|T047|238982009|SNOMEDCT_US|DIABETES MELLITUS WITH DERMATOLOGICAL MANIFESTATIONS |DIABETIC DERMOPATHY (DISORDER)
C0406682|T047|238982009|SNOMEDCT_US|DIABETES MELLITUS WITH DIABETIC DERMATITIS|DIABETIC DERMOPATHY (DISORDER)
C0406682|T047|238982009|SNOMEDCT_US|DIABETES MELLITUS WITH DIABETIC DERMATITIS |DIABETIC DERMOPATHY (DISORDER)
C0406682|T047|238982009|SNOMEDCT_US|DIABETIC DERMATITIS|DIABETIC DERMOPATHY (DISORDER)
C0406682|T047|238982009|SNOMEDCT_US|DIABETIC DERMOPATHY |DIABETIC DERMOPATHY (DISORDER)
C3250577|T047||SNOMEDCT_US|DIABETES MELLITUS WITH ORAL CAVITY MANIFESTATIONS 
C3250577|T047||SNOMEDCT_US|DIABETES MELLITUS WITH ORAL CAVITY MANIFESTATIONS
C0375121|T047||SNOMEDCT_US|DIABETES MELLITUS WITH HYPEROSMOLARITY
C0375121|T047||SNOMEDCT_US|DIABETES MELLITUS WITH HYPEROSMOLARITY 
C3534592|T047||SNOMEDCT_US|DIABETES IN CHILDREN AND TEENS
C0524620|T047|237602007|SNOMEDCT_US|SYNDROME X, REAVEN|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|DYSMETABOLIC SYNDROME X|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|DYSMETABOLIC SYNDROME X |METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|INSULIN RESISTANCE SYNDROME|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|METABOLIC SYNDROME|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|METABOLIC SYNDROME X|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|INSULIN RESISTANCE SYNDROME X|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|METABOLIC X SYNDROME|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|SYNDROME X, INSULIN RESISTANCE|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|METABOLIC SYNDROME X [DISEASE/FINDING]|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|METABOLIC CARDIOVASCULAR SYNDROME|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|REAVEN SYNDROME X|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|SYNDROME X, METABOLIC|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|CARDIOVASCULAR SYNDROME, METABOLIC|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|CARDIOVASCULAR SYNDROMES, METABOLIC|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|SYNDROME, METABOLIC CARDIOVASCULAR|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|SYNDROME X (METABOLIC)|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|METABOLIC SYNDROME X |METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|EQUINE METABOLIC SYNDROME|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|SYNDROME X, DYSMETABOLIC|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|SYNDROME, METABOLIC X|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|X SYNDROME, METABOLIC|METABOLIC SYNDROME X (DISORDER)
C0524620|T047|237602007|SNOMEDCT_US|REAVEN'S SYNDROME|METABOLIC SYNDROME X (DISORDER)
C0206172|T047|280137006|SNOMEDCT_US|DIABETIC FOOT|DIABETIC FOOT (DISORDER)
C0206172|T047|280137006|SNOMEDCT_US|FEET, DIABETIC|DIABETIC FOOT (DISORDER)
C0206172|T047|280137006|SNOMEDCT_US|FOOT, DIABETIC|DIABETIC FOOT (DISORDER)
C0206172|T047|280137006|SNOMEDCT_US|DIABETIC FEET|DIABETIC FOOT (DISORDER)
C0206172|T047|280137006|SNOMEDCT_US|DIABETIC FOOT [DISEASE/FINDING]|DIABETIC FOOT (DISORDER)
C0206172|T047|280137006|SNOMEDCT_US|DIABETIC FOOT |DIABETIC FOOT (DISORDER)
C3534591|T047||SNOMEDCT_US|DIABETIC HEART DISEASE
C0020616|T047|9356005|SNOMEDCT_US|AGENTS, HYPOGLYCEMIC|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC AGENTS|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC AGENT|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|DRUGS, HYPOGLYCEMIC|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|ANTIHYPERGLYCEMIC|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCAEMIC DRUG|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC DRUG|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|ANTI-HYPERGLYCEMICS|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|AGENTS, ANTIHYPERGLYCEMIC|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC MEDICINES|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|DIABETES MEDICINES|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|DRUGS FOR HYPOGLYCEMIA|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|DRUGS FOR HYPOGLYCAEMIA|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC PRODUCT |HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCAEMIC PRODUCT|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC PRODUCT|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|DRUGS FOR HYPOGLYCEMIA |HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC AGENT |HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCAEMIC|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|ANTIHYPERGLYCEMICS|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMICS|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|ANTIHYPERGLYCEMIC AGENTS|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC DRUGS|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCAEMIC AGENT|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC AGENT |HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC DRUG, NOS|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCAEMIC DRUG, NOS|HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|DRUGS FOR HYPOGLYCEMIA |HYPOGLYCEMIC PRODUCT (PRODUCT)
C0020616|T047|9356005|SNOMEDCT_US|HYPOGLYCEMIC DRUG |HYPOGLYCEMIC PRODUCT (PRODUCT)
C1456657|T047||SNOMEDCT_US|DIABETIC NERVE PROBLEMS
C0559093|T047|154689003|SNOMEDCT_US|DIABETES WITH OTHER COMPLICATIONS |DIABETES WITH OTHER COMPLICATIONS (DISORDER)
C0559093|T047|154689003|SNOMEDCT_US|DIABETES WITH OTHER COMPLICATIONS|DIABETES WITH OTHER COMPLICATIONS (DISORDER)
C0011870|T047|33248009|SNOMEDCT_US|DIABETES WITH OTHER COMA|DIABETES WITH NON-KETOTIC NON-HYPEROSMOLAR COMA
C0011870|T047|33248009|SNOMEDCT_US|DIABETES WITH NON-KETOTIC NON-HYPEROSMOLAR COMA |DIABETES WITH NON-KETOTIC NON-HYPEROSMOLAR COMA
C0011870|T047|33248009|SNOMEDCT_US|DIABETES WITH NON-KETOTIC NON-HYPEROSMOLAR COMA|DIABETES WITH NON-KETOTIC NON-HYPEROSMOLAR COMA
C1275078|T047|205813009|SNOMEDCT_US|CARPENTER SYNDROME|CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|TYPE II ACROCEPHALOPOLYSYNDACTYLY|CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|ACROCEPHALOPOLYSYNDACTYLY TYPE II|CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|ACPS II|CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|CARPENTER SYNDROME 1|CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|CRPT1|CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|CARPENTER SYNDROME |CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|CARPENTER 'S SYNDROME|CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|CARPENTER'S SYNDROME|CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|CARPENTER'S SYNDROME |CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|ACROCEPHALOPOLYSYNDACTYLY TYPE II |CARPENTER'S SYNDROME (DISORDER)
C1275078|T047|205813009|SNOMEDCT_US|ACROCEPHALOPOLYSYNDACTYLY TYPE 2|CARPENTER'S SYNDROME (DISORDER)
C0342254|T047|190342007|SNOMEDCT_US|DIABETES MELLITIS WITH NEPHROPATHY NOS |DIABETES MELLITIS WITH NEPHROPATHY NOS (DISORDER)
C0342254|T047|190342007|SNOMEDCT_US|DIABETES MELLITUS WITH RENAL MANIFESTATION|DIABETES MELLITIS WITH NEPHROPATHY NOS (DISORDER)
C0342254|T047|190342007|SNOMEDCT_US|DIABETES MELLITUS WITH RENAL MANIFESTATION |DIABETES MELLITIS WITH NEPHROPATHY NOS (DISORDER)
C0342254|T047|190342007|SNOMEDCT_US|DIABETES MELLITIS WITH NEPHROPATHY NOS|DIABETES MELLITIS WITH NEPHROPATHY NOS (DISORDER)
C0342290|T047|237620003|SNOMEDCT_US|ABNORMAL METABOLIC STATE IN DIABETES MELLITUS|ABNORMAL METABOLIC STATE IN DIABETES MELLITUS (DISORDER)
C0342290|T047|237620003|SNOMEDCT_US|ABNORMAL METABOLIC STATE IN DIABETES MELLITUS |ABNORMAL METABOLIC STATE IN DIABETES MELLITUS (DISORDER)
C0342264|T047|267379000|SNOMEDCT_US|DIABETES MELLITUS, JUVENILE TYPE, WITH NO MENTION OF COMPLICATION|DIABETES MELLITUS, JUVENILE TYPE, WITH NO MENTION OF COMPLICATION (DISORDER)
C0342264|T047|267379000|SNOMEDCT_US|DIABETES MELLITUS, JUVENILE TYPE, WITH NO MENTION OF COMPLICATION |DIABETES MELLITUS, JUVENILE TYPE, WITH NO MENTION OF COMPLICATION (DISORDER)
C1282941|T047|267382005|SNOMEDCT_US|DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION |DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION (DISORDER)
C1282941|T047|267382005|SNOMEDCT_US|DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION|DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION (DISORDER)
C1282941|T047|267382005|SNOMEDCT_US|DIABETIC NEUROPATHY WITH NEUROLOGICAL COMPLICATION |DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION (DISORDER)
C1282941|T047|267382005|SNOMEDCT_US|DIABETIC NEUROPATHY WITH NEUROLOGICAL COMPLICATION|DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION (DISORDER)
C1282941|T047|267382005|SNOMEDCT_US|DIABETES WITH NEUROLOGICAL MANIFESTATIONS|DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION (DISORDER)
C1282941|T047|267382005|SNOMEDCT_US|DIABETIC NEUROPATHY WITH NEUROLOGIC COMPLICATION|DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION (DISORDER)
C1282941|T047|267382005|SNOMEDCT_US|DIABETIC NEUROPATHY WITH NEUROLOGIC COMPLICATION |DIABETES MELLITUS WITH NEUROLOGICAL MANIFESTATION (DISORDER)
C0342265|T047|267380002|SNOMEDCT_US|DIABETES MELLITUS, ADULT ONSET, WITH NO MENTION OF COMPLICATION |DIABETES MELLITUS, ADULT ONSET, WITH NO MENTION OF COMPLICATION (DISORDER)
C0342265|T047|267380002|SNOMEDCT_US|DIABETES MELLITUS, ADULT ONSET, WITH NO MENTION OF COMPLICATION|DIABETES MELLITUS, ADULT ONSET, WITH NO MENTION OF COMPLICATION (DISORDER)
C0554436|T047|422275004|SNOMEDCT_US|DIABETIC GANGRENE|GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0554436|T047|422275004|SNOMEDCT_US|GANGRENE ASSOCIATED WITH DIABETES MELLITUS |GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0554436|T047|422275004|SNOMEDCT_US|GANGRENE ASSOCIATED WITH DIABETES MELLITUS|GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0554436|T047|422275004|SNOMEDCT_US|GANGRENE - DIABETIC|GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0554436|T047|422275004|SNOMEDCT_US|DIABETES MELLITUS WITH GANGRENE|GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0554436|T047|422275004|SNOMEDCT_US|DIABETES MELLITUS WITH GANGRENE |GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0554436|T047|422275004|SNOMEDCT_US|DIABETES WITH GANGRENE|GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0554436|T047|422275004|SNOMEDCT_US|DIABETIC GANGRENE |GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0554436|T047|422275004|SNOMEDCT_US|GANGRENE ASSOCIATED WITH DIABETES MELLITUS |GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0554436|T047|422275004|SNOMEDCT_US|DIABETIC GANGRENE |GANGRENE ASSOCIATED WITH DIABETES MELLITUS
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS COMPLICATING PREGNANCY, CHILDBIRTH, OR THE PUERPERIUM|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS OF MOTHER, COMP PREGNANCY,CHILDBIRTH, OR THE PUERP, UNSPEC AS TO EOC|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS OF MOTHER, COMPLICATING PREGNANCY, CHILDBIRTH, OR THE PUERPERIUM, UNSPECIFIED AS T|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES IN PREG-UNSPEC|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS IN PREGNANCY, CHILDBIRTH, AND THE PUERPERIUM|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|UNSPECIFIED DIABETES MELLITUS IN PREGNANCY, CHILDBIRTH AND THE PUERPERIUM|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS OF MOTHER, COMPLICATING PREGNANCY, CHILDBIRTH, OR THE PUERPERIUM, UNSPECIFIED AS TO EPISODE OF CARE|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS OF MOTHER, COMPLICATING PREGNANCY, CHILDBIRTH, OR THE PUERPERIUM, UNSPECIFIED AS TO EPISODE OF CARE OR NOT APPLICABLE|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS IN PREGNANCY, CHILDBIRTH, AND PUERPERIUM |DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS IN PREGNANCY, CHILDBIRTH, AND PUERPERIUM|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM |DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH OR THE PUERPERIUM NOS |DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH OR THE PUERPERIUM NOS|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS IN MOTHER COMPLICATING PREGNANCY, CHILDBIRTH, AND PUERPERIUM|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS IN MOTHER COMPLICATING PREGNANCY, CHILDBIRTH, AND PUERPERIUM |DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS IN MOTHER COMPLICATING PREGNANCY, CHILDBIRTH AND/OR PUERPERIUM |DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS IN MOTHER COMPLICATING PREGNANCY, CHILDBIRTH AND/OR PUERPERIUM|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|DIABETES MELLITUS IN MOTHER COMPLICATING PREGNANCY, CHILDBIRTH OR PUERPERIUM|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0341893|T047|199223000|SNOMEDCT_US|GESTATIONAL DIABETES COMPLICATING PREGNANCY, CHILDBIRTH, OR THE PUERPERIUM|DIABETES MELLITUS DURING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM (DISORDER)
C0348933|T047|190336008|SNOMEDCT_US|OTHER SPECIFIED DIABETES MELLITUS WITH COMA|OTHER SPECIFIED DIABETES MELLITUS WITH COMA (DISORDER)
C0348933|T047|190336008|SNOMEDCT_US|OTHER SPECIFIED DIABETES MELLITUS WITH COMA |OTHER SPECIFIED DIABETES MELLITUS WITH COMA (DISORDER)
C0342260|T047|190417004|SNOMEDCT_US|DIABETES MELLITUS NOS WITH OTHER SPECIFIED MANIFESTATION |DIABETES MELLITUS WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342260|T047|190417004|SNOMEDCT_US|DIABETES MELLITUS WITH OTHER SPECIFIED MANIFESTATION |DIABETES MELLITUS WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342260|T047|190417004|SNOMEDCT_US|DIABETES MELLITUS NOS WITH OTHER SPECIFIED MANIFESTATION|DIABETES MELLITUS WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342260|T047|190417004|SNOMEDCT_US|DIABETES MELLITUS WITH OTHER SPECIFIED MANIFESTATION|DIABETES MELLITUS WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0348931|T047|190420007|SNOMEDCT_US|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS (DISORDER)
C0348931|T047|190420007|SNOMEDCT_US|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS (DISORDER)
C0348931|T047|190420007|SNOMEDCT_US|OTH DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS (DISORDER)
C0348931|T047|190420007|SNOMEDCT_US|OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS |OTHER SPECIFIED DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS (DISORDER)
C0342261|T047|190418009|SNOMEDCT_US|TYPE I DIABETES MELLITUS WITH OTHER SPECIFIED MANIFESTATIONS|DIABETES MELLITUS, JUVENILE TYPE, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342261|T047|190418009|SNOMEDCT_US|INSULIN-DEPENDENT DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS|DIABETES MELLITUS, JUVENILE TYPE, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342261|T047|190418009|SNOMEDCT_US|TYPE 1 DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS|DIABETES MELLITUS, JUVENILE TYPE, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342261|T047|190418009|SNOMEDCT_US|TYPE 1 DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION|DIABETES MELLITUS, JUVENILE TYPE, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342261|T047|190418009|SNOMEDCT_US|DIABETES MELLITUS, JUVENILE TYPE, WITH OTHER SPECIFIED MANIFESTATION|DIABETES MELLITUS, JUVENILE TYPE, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342261|T047|190418009|SNOMEDCT_US|DIABETES MELLITUS, JUVENILE TYPE, WITH OTHER SPECIFIED MANIFESTATION |DIABETES MELLITUS, JUVENILE TYPE, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0348938|T047|190382000|SNOMEDCT_US|OTHER SPECIFIED DIABETES MELLITUS WITH MULTIPLE COMPLICATIONS|OTHER SPECIFIED DIABETES MELLITUS WITH MULTIPLE COMPLICATIONS (DISORDER)
C0348938|T047|190382000|SNOMEDCT_US|OTHER SPECIFIED DIABETES MELLITUS WITH MULTIPLE COMPLICATIONS |OTHER SPECIFIED DIABETES MELLITUS WITH MULTIPLE COMPLICATIONS (DISORDER)
C0342262|T047|190419001|SNOMEDCT_US|TYPE II DIABETES MELLITUS WITH OTHER SPECIFIED MANIFESTATIONS|DIABETES MELLITUS, ADULT ONSET, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342262|T047|190419001|SNOMEDCT_US|NON-INSULIN-DEPENDENT DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS|DIABETES MELLITUS, ADULT ONSET, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342262|T047|190419001|SNOMEDCT_US|TYPE 2 DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATIONS|DIABETES MELLITUS, ADULT ONSET, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342262|T047|190419001|SNOMEDCT_US|TYPE 2 DIABETES MELLITUS WITH OTHER SPECIFIED COMPLICATION|DIABETES MELLITUS, ADULT ONSET, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342262|T047|190419001|SNOMEDCT_US|DIABETES MELLITUS, ADULT ONSET, WITH OTHER SPECIFIED MANIFESTATION |DIABETES MELLITUS, ADULT ONSET, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C0342262|T047|190419001|SNOMEDCT_US|DIABETES MELLITUS, ADULT ONSET, WITH OTHER SPECIFIED MANIFESTATION|DIABETES MELLITUS, ADULT ONSET, WITH OTHER SPECIFIED MANIFESTATION (DISORDER)
C3646651|T047||SNOMEDCT_US|PREGNANCY COMPLICATIONS: CHRONIC DIABETES MELLITUS
C3646651|T047||SNOMEDCT_US|PREGNANCY COMPLICATED BY CHRONIC DIABETES MELLITUS 
C3646651|T047||SNOMEDCT_US|PREGNANCY COMPLICATIONS: DIABETES MELLITUS CHRONIC
C3646651|T047||SNOMEDCT_US|PREGNANCY COMPLICATED BY CHRONIC DIABETES MELLITUS
C2874125|T047|609568004|SNOMEDCT_US|DIABETES MELLITUS DUE TO GENETIC DEFECTS OF BETA-CELL FUNCTION|DIABETES MELLITUS DUE TO GENETIC DEFECT IN BETA CELL FUNCTION (DISORDER)
C2874125|T047|609568004|SNOMEDCT_US|DIABETES MELLITUS DUE TO GENETIC DEFECT IN BETA CELL FUNCTION|DIABETES MELLITUS DUE TO GENETIC DEFECT IN BETA CELL FUNCTION (DISORDER)
C2874125|T047|609568004|SNOMEDCT_US|DIABETES MELLITUS DUE TO GENETIC DEFECT IN BETA CELL FUNCTION |DIABETES MELLITUS DUE TO GENETIC DEFECT IN BETA CELL FUNCTION (DISORDER)
C2874124|T047|609569007|SNOMEDCT_US|DIABETES MELLITUS DUE TO GENETIC DEFECTS IN INSULIN ACTION|DIABETES MELLITUS DUE TO GENETIC DEFECT IN INSULIN ACTION (DISORDER)
C2874124|T047|609569007|SNOMEDCT_US|DIABETES MELLITUS DUE TO GENETIC DEFECT IN INSULIN ACTION |DIABETES MELLITUS DUE TO GENETIC DEFECT IN INSULIN ACTION (DISORDER)
C2874124|T047|609569007|SNOMEDCT_US|DIABETES MELLITUS DUE TO GENETIC DEFECT IN INSULIN ACTION|DIABETES MELLITUS DUE TO GENETIC DEFECT IN INSULIN ACTION (DISORDER)
C0271687|T047|91352004|SNOMEDCT_US|DIABETES MELLITUS DUE TO STRUCTURALLY ABNORMAL INSULIN |DIABETES MELLITUS DUE TO STRUCTURALLY ABNORMAL INSULIN (DISORDER)
C0271687|T047|91352004|SNOMEDCT_US|DIABETES MELLITUS DUE TO STRUCTURALLY ABNORMAL INSULIN|DIABETES MELLITUS DUE TO STRUCTURALLY ABNORMAL INSULIN (DISORDER)
C0271687|T047|91352004|SNOMEDCT_US|DIABETES MELLITUS DUE TO STRUCTURALLY ABNORMAL INSULIN |DIABETES MELLITUS DUE TO STRUCTURALLY ABNORMAL INSULIN (DISORDER)
C0271687|T047|91352004|SNOMEDCT_US|INSULINOPATHY|DIABETES MELLITUS DUE TO STRUCTURALLY ABNORMAL INSULIN (DISORDER)
C0271687|T047|91352004|SNOMEDCT_US|DIABETES MELLITUS DUE TO ABNORMAL INSULIN|DIABETES MELLITUS DUE TO STRUCTURALLY ABNORMAL INSULIN (DISORDER)
C0271687|T047|91352004|SNOMEDCT_US|INSULINOPATHY, NOS|DIABETES MELLITUS DUE TO STRUCTURALLY ABNORMAL INSULIN (DISORDER)
C0342274|T047|5969009|SNOMEDCT_US|DIABETES MELLITUS ASSOCIATED WITH GENETIC SYNDROME |DIABETES MELLITUS ASSOCIATED WITH GENETIC SYNDROME (DISORDER)
C0342274|T047|5969009|SNOMEDCT_US|DIABETES MELLITUS ASSOCIATED WITH GENETIC SYNDROME|DIABETES MELLITUS ASSOCIATED WITH GENETIC SYNDROME (DISORDER)
C0342274|T047|5969009|SNOMEDCT_US|GENETIC SYNDROMES OF DIABETES MELLITUS|DIABETES MELLITUS ASSOCIATED WITH GENETIC SYNDROME (DISORDER)
C0342274|T047|5969009|SNOMEDCT_US|DIABETES MELLITUS ASSOCIATED WITH GENETIC SYNDROME |DIABETES MELLITUS ASSOCIATED WITH GENETIC SYNDROME (DISORDER)
C0342283|T047|237613005|SNOMEDCT_US|HYPERPROINSULINEMIA|HYPERPROINSULINEMIA (DISORDER)
C0342283|T047|237613005|SNOMEDCT_US|HYPERPROINSULINEMIA |HYPERPROINSULINEMIA (DISORDER)
C0342283|T047|237613005|SNOMEDCT_US|DIABETES MELLITUS HYPERPROINSULINEMIA|HYPERPROINSULINEMIA (DISORDER)
C0342283|T047|237613005|SNOMEDCT_US|HYPERPROINSULINAEMIA|HYPERPROINSULINEMIA (DISORDER)
C0342283|T047|237613005|SNOMEDCT_US|HYPERPROINSULINEMIA |HYPERPROINSULINEMIA (DISORDER)
C1263962|T047|123763000|SNOMEDCT_US|HOUSSAY SYNDROME|HOUSSAY'S SYNDROME (DISORDER)
C1263962|T047|123763000|SNOMEDCT_US|HOUSSAY'S SYNDROME|HOUSSAY'S SYNDROME (DISORDER)
C1263962|T047|123763000|SNOMEDCT_US|HOUSSAY'S SYNDROME |HOUSSAY'S SYNDROME (DISORDER)
C1263962|T047|123763000|SNOMEDCT_US|HOUSSAY'S SYNDROME |HOUSSAY'S SYNDROME (DISORDER)
C1960272|T047|426875007|SNOMEDCT_US|LATENT AUTOIMMUNE DIABETES MELLITUS IN ADULT |LATENT AUTOIMMUNE DIABETES MELLITUS IN ADULT (DISORDER)
C1960272|T047|426875007|SNOMEDCT_US|LATENT AUTOIMMUNE DIABETES MELLITUS IN ADULT|LATENT AUTOIMMUNE DIABETES MELLITUS IN ADULT (DISORDER)
C1960272|T047|426875007|SNOMEDCT_US|LATENT AUTOIMMUNE DIABETES MELLITUS IN ADULT (LADA)|LATENT AUTOIMMUNE DIABETES MELLITUS IN ADULT (DISORDER)
C1960272|T047|426875007|SNOMEDCT_US|DIABETES MELLITUS LATENT AUTOIMMUNE IN ADULT|LATENT AUTOIMMUNE DIABETES MELLITUS IN ADULT (DISORDER)
C1960272|T047|426875007|SNOMEDCT_US|LATENT AUTOIMMUNE DIABETES MELLITUS IN ADULT |LATENT AUTOIMMUNE DIABETES MELLITUS IN ADULT (DISORDER)
C1960626|T047|426705001|SNOMEDCT_US|DIABETES MELLITUS ASSOCIATED WITH CYSTIC FIBROSIS|DIABETES MELLITUS ASSOCIATED WITH CYSTIC FIBROSIS (DISORDER)
C1960626|T047|426705001|SNOMEDCT_US|DIABETES MELLITUS ASSOCIATED WITH CYSTIC FIBROSIS |DIABETES MELLITUS ASSOCIATED WITH CYSTIC FIBROSIS (DISORDER)
C1960626|T047|426705001|SNOMEDCT_US|DIABETES MELLITUS ASSOCIATED WITH CYSTIC FIBROSIS |DIABETES MELLITUS ASSOCIATED WITH CYSTIC FIBROSIS (DISORDER)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE DIABETES MELLITUS|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE DIABETES MELLITUS |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES MELLITUS |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|DIABETES BRITTLE|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|LABILE DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE; DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|DIABETES; BRITTLE|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|DIABETES; UNSTABLE|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE; DIABETES|BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|BRITTLE DIABETES |BRITTLE DIABETES MELLITUS (FINDING)
C0342302|T047|11530004|SNOMEDCT_US|UNSTABLE DIABETES |BRITTLE DIABETES MELLITUS (FINDING)
C0271701|T047|75682002|SNOMEDCT_US|DM DUE TO INSULIN RECEPTOR AB|DM DUE TO INSULIN RECEPTOR AB
C0271701|T047|75682002|SNOMEDCT_US|DIABETES MELLITUS DUE TO INSULIN RECEPTOR ANTIBODIES |DM DUE TO INSULIN RECEPTOR AB
C0271701|T047|75682002|SNOMEDCT_US|DIABETES MELLITUS DUE TO INSULIN RECEPTOR ANTIBODIES|DM DUE TO INSULIN RECEPTOR AB
C0271701|T047|75682002|SNOMEDCT_US|DIABETES MELLITUS DUE TO INSULIN RECEPTOR ANTIBODIES |DM DUE TO INSULIN RECEPTOR AB
C0271701|T047|75682002|SNOMEDCT_US|DIABETES MELLITUS CAUSED BY INSULIN RECEPTOR ANTIBODIES|DM DUE TO INSULIN RECEPTOR AB
C0271701|T047|75682002|SNOMEDCT_US|DM CAUSED BY INSULIN RECEPTOR AB|DM DUE TO INSULIN RECEPTOR AB
C0271701|T047|75682002|SNOMEDCT_US|DIABETES MELLITUS CAUSED BY INSULIN RECEPTOR ANTIBODIES |DM DUE TO INSULIN RECEPTOR AB
C1720029|T047|420662003|SNOMEDCT_US|COMA ASSOCIATED WITH DIABETES MELLITUS |COMA ASSOCIATED WITH DIABETES MELLITUS (DISORDER)
C1720029|T047|420662003|SNOMEDCT_US|COMA ASSOCIATED WITH DIABETES MELLITUS|COMA ASSOCIATED WITH DIABETES MELLITUS (DISORDER)
C1720029|T047|420662003|SNOMEDCT_US|COMA ASSOCIATED WITH DIABETES MELLITUS |COMA ASSOCIATED WITH DIABETES MELLITUS (DISORDER)
C1857775|T047||SNOMEDCT_US|DIABETES MELLITUS, NEONATAL, WITH CONGENITAL HYPOTHYROIDISM
C1857775|T047||SNOMEDCT_US|NDH SYNDROME
C1835887|T047|609580007|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL, 2|TNDM2
C1835887|T047|609580007|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL, 2 |TNDM2
C1835887|T047|609580007|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL 2 |TNDM2
C1835887|T047|609580007|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL 2|TNDM2
C1835887|T047|609580007|SNOMEDCT_US|TNDM2|TNDM2
C1853564|T047||SNOMEDCT_US|DEND
C1853564|T047||SNOMEDCT_US|DEVELOPMENTAL DELAY, EPILEPSY, AND NEONATAL DIABETES
C1839028|T047||SNOMEDCT_US|MITOCHONDRIAL MYOPATHY WITH DIABETES
C1839028|T047||SNOMEDCT_US|MITOCHONDRIAL MYOPATHY, LIPID TYPE
C1864623|T047|609581006|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL, 3|TNDM3
C1864623|T047|609581006|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL, 3 |TNDM3
C1864623|T047|609581006|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL 3|TNDM3
C1864623|T047|609581006|SNOMEDCT_US|TNDM3|TNDM3
C1864623|T047|609581006|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL 3 |TNDM3
C0342278|T047|237606005|SNOMEDCT_US|DIABETES MELLITUS, INSULIN-RESISTANT, WITH ACANTHOSIS NIGRICANS|HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE (DISORDER)
C0342278|T047|237606005|SNOMEDCT_US|INSULIN RECEPTOR DEFECT WITH INSULIN-RESISTANT DIABETES MELLITUS AND ACANTHOSIS NIGRICANS|HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE (DISORDER)
C0342278|T047|237606005|SNOMEDCT_US|IRAN, TYPE A|HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE (DISORDER)
C0342278|T047|237606005|SNOMEDCT_US|DIABETES MELLITUS, INSULIN-RESISTANT, WITH ACANTHOSIS NIGRICANS, TYPE A|HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE (DISORDER)
C0342278|T047|237606005|SNOMEDCT_US|INSULIN RECEPTOR, DEFECT IN, WITH INSULIN-RESISTANT DIABETES MELLITUS AND ACANTHOSIS NIGRICANS|HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE (DISORDER)
C0342278|T047|237606005|SNOMEDCT_US|HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE|HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE (DISORDER)
C0342278|T047|237606005|SNOMEDCT_US|INSULIN-RESISTANT ACANTHOSIS NIGRICANS TYPE A|HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE (DISORDER)
C0342278|T047|237606005|SNOMEDCT_US|HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE |HEREDITARY BENIGN ACANTHOSIS NIGRICANS WITH INSULIN RESISTANCE (DISORDER)
C1864839|T047|609574004|SNOMEDCT_US|MODY7|MODY7
C1864839|T047|609574004|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG, TYPE 7|MODY7
C1864839|T047|609574004|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG, TYPE 7 |MODY7
C1864839|T047|609574004|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG - TYPE 7|MODY7
C1864839|T047|609574004|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG - TYPE 7 |MODY7
C2748662|T047||SNOMEDCT_US|MITCHELL-RILEY SYNDROME
C2748662|T047||SNOMEDCT_US|MTCHRS
C2748662|T047||SNOMEDCT_US|DIABETES, NEONATAL, WITH PANCREATIC HYPOPLASIA, INTESTINAL ATRESIA, AND GALLBLADDER APLASIA OR HYPOPLASIA
C0342281|T047|237611007|SNOMEDCT_US|MUSCULAR ATROPHY, ATAXIA, RETINITIS PIGMENTOSA, AND DIABETES MELLITUS|MUSCULAR ATROPHY, ATAXIA, RETINITIS PIGMENTOSA, AND DIABETES MELLITUS (DISORDER)
C0342281|T047|237611007|SNOMEDCT_US|MUSCULAR ATROPHY, ATAXIA, RETINITIS PIGMENTOSA, AND DIABETES MELLITUS |MUSCULAR ATROPHY, ATAXIA, RETINITIS PIGMENTOSA, AND DIABETES MELLITUS (DISORDER)
C3711391|T047||SNOMEDCT_US|TNDM TYPE 1
C3711391|T047||SNOMEDCT_US|6Q24-RELATED TRANSIENT NEONATAL DIABETES MELLITUS
C3711391|T047||SNOMEDCT_US|6Q24-TNDM
C1857958|T047||SNOMEDCT_US|DIABETES MELLITUS, CONGENITAL AUTOIMMUNE
C1836780|T047||SNOMEDCT_US|PANCREATIC AND CEREBELLAR AGENESIS
C1836780|T047||SNOMEDCT_US|PACA
C1836780|T047||SNOMEDCT_US|DIABETES MELLITUS, PERMANENT NEONATAL, WITH CEREBELLAR AGENESIS
C1859965|T047|733072002|SNOMEDCT_US|ALANINURIA WITH MICROCEPHALY, DWARFISM, ENAMEL HYPOPLASIA, AND DIABETES MELLITUS|STIMMLER SYNDROME
C1859965|T047|733072002|SNOMEDCT_US|STIMMLER SYNDROME|STIMMLER SYNDROME
C1859596|T047||SNOMEDCT_US|ATHEROSCLEROSIS, PREMATURE, WITH DEAFNESS, NEPHROPATHY, DIABETES MELLITUS, PHOTOMYOCLONUS, AND DEGENERATIVE NEUROLOGIC DISEASE
C1838782|T047||SNOMEDCT_US|WOLFRAM SYNDROME, MITOCHONDRIAL FORM
C1838782|T047||SNOMEDCT_US|DIDMOAD SYNDROME, MITOCHONDRIAL FORM
C1838782|T047||SNOMEDCT_US|DIABETES INSIPIDUS AND MELLITUS WITH OPTIC ATROPHY AND DEAFNESS, MITOCHONDRIAL FORM
C1832386|T047|609579009|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL, 1|TNDM1
C1832386|T047|609579009|SNOMEDCT_US|TNDM1|TNDM1
C1832386|T047|609579009|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL 1|TNDM1
C1832386|T047|609579009|SNOMEDCT_US|DIABETES MELLITUS, TRANSIENT NEONATAL 1 |TNDM1
C1832386|T047|609579009|SNOMEDCT_US|TNDM|TNDM1
C1832386|T047|609579009|SNOMEDCT_US|DMTN|TNDM1
C1838780|T047||SNOMEDCT_US|PANCREATIC HYPOPLASIA, CONGENITAL, WITH DIABETES MELLITUS AND CONGENITAL HEART DISEASE
C2675066|T047||SNOMEDCT_US|LYMPHEDEMA-DISTICHIASIS SYNDROME WITH RENAL DISEASE AND DIABETES MELLITUS
C1833102|T047||SNOMEDCT_US|DIABETES MELLITUS, PERMANENT NEONATAL, WITH NEUROLOGIC FEATURES
C1833104|T047|609565001|SNOMEDCT_US|DIABETES MELLITUS, PERMANENT NEONATAL|PERMANENT DIABETES MELLITUS OF INFANCY
C1833104|T047|609565001|SNOMEDCT_US|PNDM|PERMANENT DIABETES MELLITUS OF INFANCY
C1833104|T047|609565001|SNOMEDCT_US|PDMI|PERMANENT DIABETES MELLITUS OF INFANCY
C1833104|T047|609565001|SNOMEDCT_US|DIABETES MELLITUS, PERMANENT, OF INFANCY|PERMANENT DIABETES MELLITUS OF INFANCY
C1833104|T047|609565001|SNOMEDCT_US|PERMANENT DIABETES MELLITUS OF INFANCY|PERMANENT DIABETES MELLITUS OF INFANCY
C1833104|T047|609565001|SNOMEDCT_US|PERMANENT NEONATAL DIABETES MELLITUS |PERMANENT DIABETES MELLITUS OF INFANCY
C1833104|T047|609565001|SNOMEDCT_US|PERMANENT NEONATAL DIABETES MELLITUS|PERMANENT DIABETES MELLITUS OF INFANCY
C1832443|T047||SNOMEDCT_US|MARTINEZ FRIAS SYNDROME
C1832443|T047||SNOMEDCT_US|DIABETES, NEONATAL, WITH PANCREATIC HYPOPLASIA, INTESTINAL ATRESIA, AND GALLBLADDER APLASIA OR HYPOPLASIA
C1832443|T047||SNOMEDCT_US|MARTINEZ-FRIAS SYNDROME
C1832443|T047||SNOMEDCT_US|PANCREATIC HYPOPLASIA, INTESTINAL ATRESIA, AND GALLBLADDER APLASIA OR HYPOPLASIA, WITH OR WITHOUT TRACHEOESOPHAGEAL FISTULA
C3828492|T047||SNOMEDCT_US|PRE-GESTATIONAL DIABETES
C3828492|T047||SNOMEDCT_US|PREGESTATIONAL DIABETES
C3837964|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD3
C3837964|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD3 
C3837962|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD5
C3837962|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD5 
C3837966|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD1
C3837966|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD1 
C3837963|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD4
C3837963|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD4 
C3837965|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD2 
C3837965|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD2
C3837960|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD7
C3837960|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD7 
C3837961|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD6
C3837961|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS - MVCD6 
C3837959|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS
C3837959|T047||SNOMEDCT_US|DIABETES MELLITUS WITH MICROVASCULAR COMPLICATIONS 
C0021655|T047|48606007|SNOMEDCT_US|INSULIN RESISTANCE|DRUG RESISTANCE TO INSULIN (DISORDER)
C0021655|T047|48606007|SNOMEDCT_US|RESISTANCE, INSULIN|DRUG RESISTANCE TO INSULIN (DISORDER)
C0021655|T047|48606007|SNOMEDCT_US|INSULIN RESISTANCE [DISEASE/FINDING]|DRUG RESISTANCE TO INSULIN (DISORDER)
C0021655|T047|48606007|SNOMEDCT_US|INSULIN RESISTANCE |DRUG RESISTANCE TO INSULIN (DISORDER)
C0021655|T047|48606007|SNOMEDCT_US|DRUG RESISTANCE TO INSULIN|DRUG RESISTANCE TO INSULIN (DISORDER)
C0021655|T047|48606007|SNOMEDCT_US|DRUG RESISTANCE TO INSULIN |DRUG RESISTANCE TO INSULIN (DISORDER)
C3839440|T047|703136005|SNOMEDCT_US|DIABETES MELLITUS IN REMISSION |DIABETES MELLITUS IN REMISSION (DISORDER)
C3839440|T047|703136005|SNOMEDCT_US|DIABETES MELLITUS IN REMISSION|DIABETES MELLITUS IN REMISSION (DISORDER)
C3875503|T047|105401000119101|SNOMEDCT_US|DIABETES MELLITUS DUE TO PANCREATIC INJURY|DIABETES MELLITUS DUE TO PANCREATIC INJURY (DISORDER)
C3875503|T047|105401000119101|SNOMEDCT_US|DIABETES MELLITUS DUE TO PANCREATIC INJURY |DIABETES MELLITUS DUE TO PANCREATIC INJURY (DISORDER)
C3896643|T047||SNOMEDCT_US|NODAT
C3896643|T047||SNOMEDCT_US|NEW ONSET DIABETES AFTER TRANSPLANT
C0342276|T047|390715006|SNOMEDCT_US|MATURITY ONSET DIABETES MELLITUS IN YOUNG|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MODY|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MASON-TYPE DIABETES|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|DIABETES, MATURITY-ONSET, OF THE YOUNG (MODY)|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MATURITY ONSET DIABETES IN YOUTH TYPE 1|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG |DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MATURITY ONSET DIABETES MELLITUS IN YOUNG |DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MODY - MATURITY ONSET DIABETES IN YOUTH TYPE 1|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|DIABETES MELLITUS AUTOSOMAL DOMINANT |DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|DIABETES MELLITUS AUTOSOMAL DOMINANT|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|AUTOSOMAL DOMINANT DIABETES MELLITUS|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MODY - MATURITY ONSET DIABETES IN YOUTH TYPE I|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MATURITY ONSET DIABETES IN YOUTH|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|NIDDY|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MATURITY-ONSET DIABETES OF THE YOUNG |DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0342276|T047|390715006|SNOMEDCT_US|MATURITY ONSET DIABETES OF THE YOUNG|DIABETES MELLITUS AUTOSOMAL DOMINANT (DISORDER)
C0854110|T047||SNOMEDCT_US|INSULIN-RESISTANT DIABETES MELLITUS
C0854110|T047||SNOMEDCT_US|INSULIN RESISTANT DIABETES
C0854110|T047||SNOMEDCT_US|INSULIN-RESISTANT DIABETES
C0854110|T047||SNOMEDCT_US|INSULIN RESISTANT DIABETES MELLITUS
C0854110|T047||SNOMEDCT_US|INSULIN RESISTANT DIABETES (MELLITUS)
C0854110|T047||SNOMEDCT_US|DIABETES MELLITUS, INSULIN-RESISTANT
C4039625|T047|709147009|SNOMEDCT_US|GINGIVITIS CO-OCCURRENT WITH DIABETES MELLITUS|GINGIVITIS CO-OCCURRENT WITH DIABETES MELLITUS (DISORDER)
C4039625|T047|709147009|SNOMEDCT_US|GINGIVITIS CO-OCCURRENT WITH DIABETES MELLITUS |GINGIVITIS CO-OCCURRENT WITH DIABETES MELLITUS (DISORDER)
C0477821|T047|200505002|SNOMEDCT_US|PRE-EXISTING DIABETES MELLITUS, UNSPECIFIED|[X]PRE-EXISTING DIABETES MELLITUS, UNSPECIFIED (DISORDER)
C0477821|T047|200505002|SNOMEDCT_US|[X]PRE-EXISTING DIABETES MELLITUS, UNSPECIFIED |[X]PRE-EXISTING DIABETES MELLITUS, UNSPECIFIED (DISORDER)
C0477821|T047|200505002|SNOMEDCT_US|[X]PRE-EXISTING DIABETES MELLITUS, UNSPECIFIED|[X]PRE-EXISTING DIABETES MELLITUS, UNSPECIFIED (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|SYNDROME, WOLFRAM|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|WOLFRAM SYNDROME|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIDMOAD|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|WOLFRAM SYNDROME 1|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|WFS1|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|WOLFRAM SYNDROME [DISEASE/FINDING]|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIDMOAD SYNDROME|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIABETES INSIPIDUS AND MELLITUS WITH OPTIC ATROPHY AND DEAFNESS|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS |DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIABETES INSIPIDUS, DIABETES MELLITUS, OPTIC ATROPHY, AND DEAFNESS|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIDMOADUD|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIABETES INSIPIDUS,DIABETES MELLITUS, OPTIC ATROPHY AND DEAFNESS|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIABETES INSIPIDUS, DIABETES MELLITUS, OPTIC ATROPHY AND DEAFNESS|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIDMOAD - DIABETES INSIPIDUS, DIABETES MELLITUS, OPTIC ATROPHY AND DEAFNESS|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIDMOAD - DIABETES INSIPIDUS,DIABETES MELLITUS, OPTIC ATROPHY AND DEAFNESS|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|WFS|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|MARQUARDT-LORIAUX SYNDROME|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS |DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C0043207|T047|70694009|SNOMEDCT_US|DIABETES INSIPIDUS,DIABETES MELLITUS, OPTIC ATROPHY AND DEAFNESS |DIABETES MELLITUS AND INSIPIDUS WITH OPTIC ATROPHY AND DEAFNESS (DISORDER)
C1283034|T047|359939009|SNOMEDCT_US|MATERNAL DIABETES MELLITUS|MATERNAL DIABETES MELLITUS (DISORDER)
C1283034|T047|359939009|SNOMEDCT_US|MATERNAL DIABETES MELLITUS |MATERNAL DIABETES MELLITUS (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|PINEAL HYPERPLASIA, INSULIN-RESISTANT DIABETES MELLITUS, AND SOMATIC ABNORMALITIES|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|RABSON-MENDENHALL SYNDROME|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|RABSON MENDENHALL SYNDROME|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|SYNDROME, MENDENHALL|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|SYNDROME, RABSON-MENDENHALL|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME |PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|DIABETES MELLITUS ASSOCIATED WITH GENETIC SYNDROME PINEAL HYPERPLASIA|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|MENDENHALL SYNDROME|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|PINEAL HYPERPLASIA, INSULIN-RESISTANT DIABETES MELLITUS AND SOMATIC ABNORMALITIES|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME |PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271695|T047|33559001|SNOMEDCT_US|PINEAL HYPERPLASIA, INSULIN-RESISTANT DIABETES MELLITUS AND SOMATIC ABNORMALITIES |PINEAL HYPERPLASIA AND DIABETES MELLITUS SYNDROME (DISORDER)
C0271670|T047|82260000|SNOMEDCT_US|PREGESTATIONAL DIABETES MELLITUS AND/OR IMPAIRED GLUCOSE TOLERANCE, MODIFIED WHITE CLASS R |PREGESTATIONAL DIABETES MELLITUS AND/OR IMPAIRED GLUCOSE TOLERANCE, MODIFIED WHITE CLASS R (DISORDER)
C0271670|T047|82260000|SNOMEDCT_US|PREGESTATIONAL DIABETES MELLITUS AND/OR IMPAIRED GLUCOSE TOLERANCE, MODIFIED WHITE CLASS R|PREGESTATIONAL DIABETES MELLITUS AND/OR IMPAIRED GLUCOSE TOLERANCE, MODIFIED WHITE CLASS R (DISORDER)
C0271670|T047|82260000|SNOMEDCT_US|PREGESTATIONAL DIABETES MELLITUS OR IMPAIRED GLUCOSE TOLERANCE, MODIFIED WHITE CLASS R|PREGESTATIONAL DIABETES MELLITUS AND/OR IMPAIRED GLUCOSE TOLERANCE, MODIFIED WHITE CLASS R (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|INSULIN AUTOIMMUNE SYNDROME|INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|AUTOIMMUNE ENDOCRINE DISEASE INSULIN SYNDROME|INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|AUTOIMMUNE INSULIN SYNDROME|INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|AUTOIMMUNE INSULIN SYNDROME |INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0854359|T047|408539000|SNOMEDCT_US|INSULIN AUTOIMMUNE SYNDROME |INSULIN AUTOIMMUNE SYNDROME (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|DIABETES MELLITUS, LIPOATROPHIC|LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|LIPOATROPHIC DIABETES MELLITUS|LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|LIPOATROPHIC DIABETES|LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|DIABETES MELLITUS, LIPOATROPHIC [DISEASE/FINDING]|LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|DIABETES, LIPOATROPHIC|LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|LIPOATROPHIC DIABETE|LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|DIABETE, LIPOATROPHIC|LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|LIPOATROPHIC DIABETES |LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|LIPODYSTROPHIC DIABETES|LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|LIPOATROPHIC DIABETES, NOS|LIPOATROPHIC DIABETES (DISORDER)
C0011859|T047|127012008|SNOMEDCT_US|LIPODYSTROPHIC DIABETES, NOS|LIPOATROPHIC DIABETES (DISORDER)
C0154183|T047||SNOMEDCT_US|DIABETES WITH OTHER SPECIFIED MANIFESTATIONS
C0154172|T047||SNOMEDCT_US|TYPE I DIABETES MELLITUS WITH HYPEROSMOLAR COMA
C0235397|T047||SNOMEDCT_US|DIABETES MELLITUS PRECIPITATED
C0235398|T047||SNOMEDCT_US|DIABETES MELLITUS AGGRAVATED
C0235398|T047||SNOMEDCT_US|DIABETES MELLITUS EXACERBATED
C0235399|T047||SNOMEDCT_US|DIABETES MELLITUS REACTIVATED
C0241861|T047||SNOMEDCT_US|DIABETES; STABLE
C0241861|T047||SNOMEDCT_US|STABLE; DIABETES
C0342297|T047|190331003|SNOMEDCT_US|DIABETES MELLITUS, ADULT ONSET, WITH HYPEROSMOLAR COMA |DIABETES MELLITUS, ADULT ONSET, WITH HYPEROSMOLAR COMA (DISORDER)
C0342297|T047|190331003|SNOMEDCT_US|TYPE 2 DIABETES MELLITUS WITH HYPEROSMOLAR COMA|DIABETES MELLITUS, ADULT ONSET, WITH HYPEROSMOLAR COMA (DISORDER)
C0342297|T047|190331003|SNOMEDCT_US|TYPE 2 DIABETES MELLITUS WITH HYPEROSMOLAR COMA |DIABETES MELLITUS, ADULT ONSET, WITH HYPEROSMOLAR COMA (DISORDER)
C0342297|T047|190331003|SNOMEDCT_US|DIABETES MELLITUS, ADULT ONSET, WITH HYPEROSMOLAR COMA|DIABETES MELLITUS, ADULT ONSET, WITH HYPEROSMOLAR COMA (DISORDER)
C0342297|T047|190331003|SNOMEDCT_US|TYPE II DIABETES MELLITUS WITH HYPEROSMOLAR COMA|DIABETES MELLITUS, ADULT ONSET, WITH HYPEROSMOLAR COMA (DISORDER)
C0494293|T047||SNOMEDCT_US|OTHER SPECIFIED DIABETES MELLITUS WITHOUT COMPLICATIONS
C0342269|T047|190447002|SNOMEDCT_US|STEROID-INDUCED DIABETES|STEROID-INDUCED DIABETES (DISORDER)
C0342269|T047|190447002|SNOMEDCT_US|STEROID-INDUCED DIABETES |STEROID-INDUCED DIABETES (DISORDER)
C0342269|T047|190447002|SNOMEDCT_US|DIABETES STEROID-INDUCED|STEROID-INDUCED DIABETES (DISORDER)
C0546950|T047||SNOMEDCT_US|TYPE II DIABETES MELLITUS WITHOUT MENTION OF COMPLICATION
C0011884|T047|4855003|SNOMEDCT_US|DIABETIC RETINOPATHIES|DR
C0011884|T047|4855003|SNOMEDCT_US|DIABETIC RETINOPATHY|DR
C0011884|T047|4855003|SNOMEDCT_US|RETINOPATHIES, DIABETIC|DR
C0011884|T047|4855003|SNOMEDCT_US|RETINOPATHY, DIABETIC|DR
C0011884|T047|4855003|SNOMEDCT_US|DR - DIABETIC RETINOPATHY|DR
C0011884|T047|4855003|SNOMEDCT_US|DIABETIC RETINOPATHY [DISEASE/FINDING]|DR
C0011884|T047|4855003|SNOMEDCT_US|RETINOPATHY;DIABETIC|DR
C0011884|T047|4855003|SNOMEDCT_US|RETINOPATHY - DIABETIC|DR
C0011884|T047|4855003|SNOMEDCT_US|RETINAL ABNORMALITY - DIABETES-RELATED |DR
C0011884|T047|4855003|SNOMEDCT_US|RETINAL ABNORMALITY - DIABETES-RELATED|DR
C0011884|T047|4855003|SNOMEDCT_US|DIABETIC RETINOPATHY NOS |DR
C0011884|T047|4855003|SNOMEDCT_US|DIABETIC RETINOPATHY |DR
C0011884|T047|4855003|SNOMEDCT_US|DIABETIC RETINOPATHY NOS|DR
C0011884|T047|4855003|SNOMEDCT_US|DIABETES WITH DIABETIC RETINOPATHY|DR
C0011884|T047|4855003|SNOMEDCT_US|DIABETES WITH DIABETIC RETINOPATHY |DR
C0011884|T047|4855003|SNOMEDCT_US|DIABETES MELLITUS WITH DIABETIC RETINOPATHY|DR
C0011884|T047|4855003|SNOMEDCT_US|RETINOPATHY DIABETIC|DR
C0011884|T047|4855003|SNOMEDCT_US|DIABETIC RETINOPATHY, NOS|DR
C0865162|T047||SNOMEDCT_US|DIABETES MELLITUS WITHOUT MENTION OF COMPLICATION OR MANIFESTATION
