// CUI|TUI|TTY|CODE|VOCAB|TXT|PREF TEXT
C000001|T109|UNK|1|CUSTOM|aspirin|aspirin
C000002|T019|UNK|2|CUSTOM|heart attack|heart attack
C000003|T109|UNK|3|CUSTOM|COPD|COPD