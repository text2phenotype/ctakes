C0412621|T060|241549007|SNOMEDCT_US|COMPUTED TOMOGRAPHY (CT) OF LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0882012|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:LIVER:NARRATIVE:COMPUTERIZED TOMOGRAPHY
C2317166|T060|429862006|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER WITH CONTRAST |COMPUTED TOMOGRAPHY OF LIVER WITH CONTRAST
C2317166|T060|429862006|SNOMEDCT_US|COMPUTED TOMOGRAPHY (CT) OF LIVER WITH CONTRAST|COMPUTED TOMOGRAPHY OF LIVER WITH CONTRAST
C2317166|T060|429862006|SNOMEDCT_US|CT SCAN OF LIVER WITH CONTRAST|COMPUTED TOMOGRAPHY OF LIVER WITH CONTRAST
C2317166|T060|429862006|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER WITH CONTRAST|COMPUTED TOMOGRAPHY OF LIVER WITH CONTRAST
C2317166|T060|429862006|SNOMEDCT_US|CT OF LIVER WITH CONTRAST|COMPUTED TOMOGRAPHY OF LIVER WITH CONTRAST
C2315699|T060|432905004|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER AND PORTAL VEIN |COMPUTED TOMOGRAPHY (CT) OF LIVER AND PORTAL VEIN
C2315699|T060|432905004|SNOMEDCT_US|COMPUTED TOMOGRAPHY (CT) OF LIVER AND PORTAL VEIN|COMPUTED TOMOGRAPHY (CT) OF LIVER AND PORTAL VEIN
C2315699|T060|432905004|SNOMEDCT_US|CT OF LIVER AND PORTAL VEIN|COMPUTED TOMOGRAPHY (CT) OF LIVER AND PORTAL VEIN
C2315699|T060|432905004|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER AND PORTAL VEIN|COMPUTED TOMOGRAPHY (CT) OF LIVER AND PORTAL VEIN
C2585273|T060|438305004|SNOMEDCT_US|COMPUTED TOMOGRAPHY DUAL PHASE STUDY OF LIVER |COMPUTED TOMOGRAPHY DUAL PHASE STUDY OF LIVER
C2585273|T060|438305004|SNOMEDCT_US|COMPUTED TOMOGRAPHY DUAL PHASE STUDY OF LIVER|COMPUTED TOMOGRAPHY DUAL PHASE STUDY OF LIVER
C2585273|T060|438305004|SNOMEDCT_US|CT DUAL PHASE STUDY OF LIVER|COMPUTED TOMOGRAPHY DUAL PHASE STUDY OF LIVER
C2585560|T060|438591004|SNOMEDCT_US|COMPUTED TOMOGRAPHY TRIPLE PHASE STUDY OF LIVER |COMPUTED TOMOGRAPHY TRIPLE PHASE STUDY OF LIVER (PROCEDURE)
C2585560|T060|438591004|SNOMEDCT_US|COMPUTED TOMOGRAPHY TRIPLE PHASE STUDY OF LIVER|COMPUTED TOMOGRAPHY TRIPLE PHASE STUDY OF LIVER (PROCEDURE)
C2585560|T060|438591004|SNOMEDCT_US|CT TRIPLE PHASE STUDY OF LIVER|COMPUTED TOMOGRAPHY TRIPLE PHASE STUDY OF LIVER (PROCEDURE)
C2321544|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER FIRST WITHOUT, THEN WITH CONTRAST
C2321544|T060||SNOMEDCT_US|CT SCAN OF LIVER FIRST WITHOUT, THEN WITH CONTRAST
C2321544|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER FIRST WITHOUT, THEN WITH CONTRAST 
C0412621|T060|241549007|SNOMEDCT_US|CT OF LIVER |COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER |COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|ABDOMINAL COMPUTED TOMOGRAPHY LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|COMPUTED TOMOGRAPHY (CT) OF LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|CT SCAN OF LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|CT OF LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|CT SCAN OF LIVER |COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|COMPUTERISED TOMOGRAM LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|CT SCAN LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|COMPUTERIZED TOMOGRAM LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|CT SCAN;LIVER|COMPUTED TOMOGRAPHY OF LIVER
C0412621|T060|241549007|SNOMEDCT_US|CT SCAN OF THE LIVER|COMPUTED TOMOGRAPHY OF LIVER
C2321546|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER WITHOUT CONTRAST
C2321546|T060||SNOMEDCT_US|CT SCAN OF LIVER WITHOUT CONTRAST
C2321546|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF LIVER WITHOUT CONTRAST 
C3697202|T060|699586000|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF LIVER USING YTTRIUM 90 MICROSPHERES|POSITRON EMISSION TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF LIVER USING YTTRIUM 90 MICROSPHERES (PROCEDURE)
C3697202|T060|699586000|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF LIVER USING YTTRIUM 90 MICROSPHERES |POSITRON EMISSION TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF LIVER USING YTTRIUM 90 MICROSPHERES (PROCEDURE)
C1636186|T060|418158005|SNOMEDCT_US|CT AND DRAINAGE OF LIVER|COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER
C1636186|T060|418158005|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER |COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER
C1636186|T060|418158005|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER|COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER
C1640379|T060|418458003|SNOMEDCT_US|CT AND ASPIRATION OF LIVER|COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER
C1640379|T060|418458003|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER |COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER
C1640379|T060|418458003|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER|COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER
C1628488|T060|418749009|SNOMEDCT_US|CT AND BIOPSY OF LIVER|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER
C1628488|T060|418749009|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER |COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER
C1628488|T060|418749009|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER
C0882012|T060||SNOMEDCT_US|LIVER CT
C0882012|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:LIVER:NARRATIVE:COMPUTERIZED TOMOGRAPHY
C0882012|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMEN>LIVER:DOC:CT
C0882012|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1652991|T060||SNOMEDCT_US|CHEST AND ABDOMEN CT W CONTRAST IV
C1652991|T060||SNOMEDCT_US|CHEST+ABD CT W CONTR IV
C1652991|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:CHEST+ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1652991|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:CHEST+ABDOMEN:DOC:CT
C3533360|T060||SNOMEDCT_US|ABDOMEN AND PELVIS MRI W CONTRAST PO AND WO AND W CONTRAST IV
C3533360|T060||SNOMEDCT_US|ABD+PELVIS MRI W CONTR PO+WO+W IV
C3533360|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST ORAL+WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN+PELVIS:DOCUMENT:MRI
C3533360|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST PO+WO & W CONTRAST IV:FIND:PT:ABDOMEN+PELVIS:DOC:MRI
C1524450|T060||SNOMEDCT_US|ABD CT LTD W CONTR IV
C1524450|T060||SNOMEDCT_US|ABDOMEN CT LIMITED W CONTRAST IV
C1524450|T060||SNOMEDCT_US|MULTISECTION LIMITED^W CONTRAST IV:FIND:PT:ABDOMEN:DOC:CT
C1524450|T060||SNOMEDCT_US|MULTISECTION LIMITED^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1524458|T060||SNOMEDCT_US|ABDOMEN CT LIMITED WO CONTRAST
C1524458|T060||SNOMEDCT_US|ABD CT LTD WO CONTR
C1524458|T060||SNOMEDCT_US|MULTISECTION LIMITED^WO CONTRAST:FIND:PT:ABDOMEN:DOC:CT
C1524458|T060||SNOMEDCT_US|MULTISECTION LIMITED^WO CONTRAST:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1524809|T060||SNOMEDCT_US|ABDOMEN CT WO CONTRAST
C1524809|T060||SNOMEDCT_US|ABD CT WO CONTR
C1524809|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FIND:PT:ABDOMEN:DOC:CT
C1524809|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1830219|T060||SNOMEDCT_US|ABD CT WO+W RED CONTR VOL IV
C1830219|T060||SNOMEDCT_US|MULTISECTION^WO & W REDUCED CONTRAST VOLUME IV:FIND:PT:ABDOMEN:DOC:CT
C1830219|T060||SNOMEDCT_US|ABDOMEN CT WO AND W REDUCED CONTRAST VOLUME IV
C1830219|T060||SNOMEDCT_US|MULTISECTION^WO & W REDUCED CONTRAST VOLUME INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1525189|T060||SNOMEDCT_US|ABD+PELVIS CT W CONTR IV
C1525189|T060||SNOMEDCT_US|ABDOMEN AND PELVIS CT W CONTRAST IV
C1525189|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:ABDOMEN+PELVIS:DOC:CT
C1525189|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN+PELVIS:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1644645|T060||SNOMEDCT_US|ABDOMEN CT
C1644645|T060||SNOMEDCT_US|ABD CT
C1644645|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:COMPUTERIZED TOMOGRAPHY
C1644645|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1644645|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMEN:DOC:CT
C1114439|T060||SNOMEDCT_US|LIVER CT WO CONTRAST
C1114439|T060||SNOMEDCT_US|LIVER CT WO CONTR
C1114439|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1114439|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FIND:PT:ABDOMEN>LIVER:DOC:CT
C1715387|T060||SNOMEDCT_US|ABD+PELVIS CT
C1715387|T060||SNOMEDCT_US|ABDOMEN AND PELVIS CT
C1715387|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMEN+PELVIS:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1715387|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMEN+PELVIS:DOC:CT
C1715410|T060||SNOMEDCT_US|ABD+PELVIS RI FOR TUMOR
C1715410|T060||SNOMEDCT_US|ABDOMEN AND PELVIS SCAN FOR TUMOR
C1715410|T060||SNOMEDCT_US|VIEWS FOR TUMOR:FINDING:POINT IN TIME:ABDOMEN+PELVIS:DOCUMENT:RADNUC
C1715410|T060||SNOMEDCT_US|VIEWS FOR TUMOR:FIND:PT:ABDOMEN+PELVIS:DOC:RADNUC
C1114428|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST:FIND:PT:ABDOMEN:DOC:CT
C1114428|T060||SNOMEDCT_US|DEPRECATED ABD CT W CONTR
C1114428|T060||SNOMEDCT_US|DEPRECATED ABDOMEN CT W CONTRAST
C1114428|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1525284|T060||SNOMEDCT_US|ABD+PELVIS CT WO CONTR
C1525284|T060||SNOMEDCT_US|ABDOMEN AND PELVIS CT WO CONTRAST
C1525284|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FIND:PT:ABDOMEN+PELVIS:DOC:CT
C1525284|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FINDING:POINT IN TIME:ABDOMEN+PELVIS:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1630749|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:ABDOMEN+PELVIS:DOC:CT
C1630749|T060||SNOMEDCT_US|ABDOMEN AND PELVIS CT WO AND W CONTRAST IV
C1630749|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN+PELVIS:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1630749|T060||SNOMEDCT_US|ABD+PELVIS CT WO+W CONTR IV
C1631257|T060||SNOMEDCT_US|CHEST AND ABDOMEN CT WO CONTRAST
C1631257|T060||SNOMEDCT_US|CHEST+ABD CT WO CONTR
C1524601|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:ABDOMEN:DOC:CT
C1524601|T060||SNOMEDCT_US|ABDOMEN CT WO AND W CONTRAST IV
C1524601|T060||SNOMEDCT_US|ABD CT WO+W CONTR IV
C1524601|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C0882540|T060||SNOMEDCT_US|LIVER CT W CONTR IV
C0882540|T060||SNOMEDCT_US|LIVER CT W CONTRAST IV
C0882540|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C0882540|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:ABDOMEN>LIVER:DOC:CT
C1114440|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:ABDOMEN>LIVER:DOC:CT
C1114440|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1114440|T060||SNOMEDCT_US|LIVER CT WO+W CONTR IV
C1114440|T060||SNOMEDCT_US|LIVER CT WO AND W CONTRAST IV
C1631258|T060||SNOMEDCT_US|CHEST+ABD CT WO+W CONTR IV
C1631258|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:CHEST+ABDOMEN:DOC:CT
C1631258|T060||SNOMEDCT_US|CHEST AND ABDOMEN CT WO AND W CONTRAST IV
C1631258|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:CHEST+ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C4070458|T060||SNOMEDCT_US|CHEST AND ABDOMEN CT 3D POST PROCESSING WO CONTRAST
C4070458|T060||SNOMEDCT_US|CHEST+ABD CT P 3D PROC WO CONTR
C4070458|T060||SNOMEDCT_US|MULTISECTION 3D POST PROCESSING^WO CONTRAST:FIND:PT:CHEST+ABDOMEN:DOC:CT
C4070458|T060||SNOMEDCT_US|MULTISECTION 3D POST PROCESSING^WO CONTRAST:FINDING:POINT IN TIME:CHEST+ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C4070453|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:ABDOMEN:DOC:CT
C4070453|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C4070453|T060||SNOMEDCT_US|ABD CT W CONTR IV
C4070453|T060||SNOMEDCT_US|ABDOMEN CT W CONTRAST IV
C4070490|T060||SNOMEDCT_US|ABD+PELVIS CT P 3D PROC WO CONTR
C4070490|T060||SNOMEDCT_US|MULTISECTION 3D POST PROCESSING^WO CONTRAST:FINDING:POINT IN TIME:ABDOMEN+PELVIS:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C4070490|T060||SNOMEDCT_US|ABDOMEN AND PELVIS CT 3D POST PROCESSING WO CONTRAST
C4070490|T060||SNOMEDCT_US|MULTISECTION 3D POST PROCESSING^WO CONTRAST:FIND:PT:ABDOMEN+PELVIS:DOC:CT
C4070489|T060||SNOMEDCT_US|ABDOMEN CT 3D POST PROCESSING WO CONTRAST
C4070489|T060||SNOMEDCT_US|MULTISECTION 3D POST PROCESSING^WO CONTRAST:FIND:PT:ABDOMEN:DOC:CT
C4070489|T060||SNOMEDCT_US|MULTISECTION 3D POST PROCESSING^WO CONTRAST:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C4070489|T060||SNOMEDCT_US|ABD CT P 3D PROC WO CONTR
C0412620|T060|303670004|SNOMEDCT_US|CT OF ABDOMEN |COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|CT OF ABDOMINAL ORGANS |COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN |COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|CT OF ABDOMEN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|CT SCAN OF ABDOMEN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|ABDOMINAL CT SCAN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|C.A.T. SCAN OF ABDOMEN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|CT SCAN ABDOMEN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS |COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|CT OF ABDOMINAL ORGANS|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|COMPUTED TOMOGRAPHY, ABDOMEN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|CT SCAN - ABDOMINAL|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|COMPUTERIZED AXIAL TOMOGRAPHY OF ABDOMEN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|CT SCAN;ABDOMEN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412620|T060|303670004|SNOMEDCT_US|CT SCAN OF THE ABDOMEN|COMPUTED TOMOGRAPHY OF ABDOMINAL ORGANS
C0412694|T060|241622002|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING (MRI) OF LIVER|MAGNETIC RESONANCE IMAGING OF LIVER (PROCEDURE)
C1644183|T060|418234000|SNOMEDCT_US|RADIONUCLIDE LIVER AND SPLEEN STUDY|RADIONUCLIDE LIVER AND SPLEEN IMAGING PROCEDURE
C2314954|T060|431839003|SNOMEDCT_US|MRI OF LIVER WITH CONTRAST|MAGNETIC RESONANCE IMAGING OF LIVER WITH CONTRAST (PROCEDURE)
C2315791|T060|432633002|SNOMEDCT_US|MRI OF LIVER AND BILIARY TRACT WITH CONTRAST|MAGNETIC RESONANCE IMAGING (MRI) OF LIVER AND BILIARY TRACT WITH CONTRAST
C2318037|T060|409901000119107|SNOMEDCT_US|MRI OF LIVER WITHOUT CONTRAST|MAGNETIC RESONANCE IMAGING OF LIVER WITHOUT CONTRAST
C1524478|T060||SNOMEDCT_US|ABD MRI W CONTR IV
C1524478|T060||SNOMEDCT_US|ABDOMEN MRI W CONTRAST IV
C1524478|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:MRI
C1524478|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:ABDOMEN:DOC:MRI
C1527050|T060||SNOMEDCT_US|LIVER MRI
C1527050|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:LIVER:NARRATIVE:MRI
C1527050|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:LIVER:DOC:MRI
C1527050|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:LIVER:DOCUMENT:MRI
C0881795|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:MRI
C0881795|T060||SNOMEDCT_US|ABDOMEN MRI
C0881795|T060||SNOMEDCT_US|ABD MRI
C0881795|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMEN:DOC:MRI
C0881795|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:MRI
C1524565|T060||SNOMEDCT_US|LIVER MRI W CONTR IV
C1524565|T060||SNOMEDCT_US|LIVER MRI W CONTRAST IV
C1524565|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:LIVER:DOC:MRI
C1524565|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:MRI
C1114492|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:MRI
C1114492|T060||SNOMEDCT_US|LIVER MRI WO+W CONTR IV
C1114492|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:LIVER:DOC:MRI
C1114492|T060||SNOMEDCT_US|LIVER MRI WO AND W CONTRAST IV
C1525274|T060||SNOMEDCT_US|CHEST AND ABDOMEN MRI W CONTRAST IV
C1525274|T060||SNOMEDCT_US|CHEST+ABD MRI W CONTR IV
C1525274|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:CHEST+ABDOMEN:DOCUMENT:MRI
C1525274|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:CHEST+ABDOMEN:DOC:MRI
C1714786|T060||SNOMEDCT_US|LIVER MRI WO+W FERUMOXIDES IV
C1714786|T060||SNOMEDCT_US|LIVER MRI WO AND W FERUMOXIDES IV
C1714786|T060||SNOMEDCT_US|MULTISECTION^WO & W FERUMOXIDES INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:MRI
C1714786|T060||SNOMEDCT_US|MULTISECTION^WO & W FERUMOXIDES IV:FIND:PT:LIVER:DOC:MRI
C3533799|T060||SNOMEDCT_US|ABDOMEN AND PELVIS MRI W CONTRAST PO AND WO CONTRAST IV
C3533799|T060||SNOMEDCT_US|ABD+PELVIS MRI W CONTR PO+WO IV
C3533799|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST PO+WO CONTRAST IV:FIND:PT:ABDOMEN+PELVIS:DOC:MRI
C3533799|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST ORAL+WO CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN+PELVIS:DOCUMENT:MRI
C1114491|T060||SNOMEDCT_US|LIVER MRI WO CONTRAST
C1114491|T060||SNOMEDCT_US|LIVER MRI WO CONTR
C1114491|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FIND:PT:LIVER:DOC:MRI
C1114491|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FINDING:POINT IN TIME:LIVER:DOCUMENT:MRI
C0412694|T060|241622002|SNOMEDCT_US|MRI OF LIVER |MAGNETIC RESONANCE IMAGING OF LIVER (PROCEDURE)
C0412694|T060|241622002|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER |MAGNETIC RESONANCE IMAGING OF LIVER (PROCEDURE)
C0412694|T060|241622002|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING (MRI) OF LIVER|MAGNETIC RESONANCE IMAGING OF LIVER (PROCEDURE)
C0412694|T060|241622002|SNOMEDCT_US|MRI OF LIVER|MAGNETIC RESONANCE IMAGING OF LIVER (PROCEDURE)
C0412694|T060|241622002|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER|MAGNETIC RESONANCE IMAGING OF LIVER (PROCEDURE)
C2317182|T060|432551009|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING (MRI) OF LIVER AND SPLEEN|MAGNETIC RESONANCE IMAGING OF LIVER AND SPLEEN
C2317182|T060|432551009|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER AND SPLEEN |MAGNETIC RESONANCE IMAGING OF LIVER AND SPLEEN
C2317182|T060|432551009|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER AND SPLEEN|MAGNETIC RESONANCE IMAGING OF LIVER AND SPLEEN
C2317182|T060|432551009|SNOMEDCT_US|MRI OF LIVER AND SPLEEN|MAGNETIC RESONANCE IMAGING OF LIVER AND SPLEEN
C2314954|T060|431839003|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER WITH CONTRAST |MAGNETIC RESONANCE IMAGING OF LIVER WITH CONTRAST (PROCEDURE)
C2314954|T060|431839003|SNOMEDCT_US|ABDOMINAL MRI LIVER WITH CONTRAST|MAGNETIC RESONANCE IMAGING OF LIVER WITH CONTRAST (PROCEDURE)
C2314954|T060|431839003|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER WITH CONTRAST|MAGNETIC RESONANCE IMAGING OF LIVER WITH CONTRAST (PROCEDURE)
C2314954|T060|431839003|SNOMEDCT_US|MRI OF LIVER WITH CONTRAST|MAGNETIC RESONANCE IMAGING OF LIVER WITH CONTRAST (PROCEDURE)
C2318037|T060|409901000119107|SNOMEDCT_US|ABDOMINAL MRI LIVER WITHOUT CONTRAST|MAGNETIC RESONANCE IMAGING OF LIVER WITHOUT CONTRAST
C2318037|T060|409901000119107|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER WITHOUT CONTRAST |MAGNETIC RESONANCE IMAGING OF LIVER WITHOUT CONTRAST
C2318037|T060|409901000119107|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER WITHOUT CONTRAST|MAGNETIC RESONANCE IMAGING OF LIVER WITHOUT CONTRAST
C2318039|T060||SNOMEDCT_US|ABDOMINAL MRI LIVER WITHOUT, THEN WITH CONTRAST
C2318039|T060||SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER WITHOUT, THEN WITH CONTRAST 
C2318039|T060||SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER WITHOUT, THEN WITH CONTRAST
C2315791|T060|432633002|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING (MRI) OF LIVER AND BILIARY TRACT WITH CONTRAST|MAGNETIC RESONANCE IMAGING (MRI) OF LIVER AND BILIARY TRACT WITH CONTRAST
C2315791|T060|432633002|SNOMEDCT_US|HEPATOBILIARY MAGNETIC RESONANCE IMAGING (MRI) WITH CONTRAST|MAGNETIC RESONANCE IMAGING (MRI) OF LIVER AND BILIARY TRACT WITH CONTRAST
C2315791|T060|432633002|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER AND BILIARY TRACT WITH CONTRAST |MAGNETIC RESONANCE IMAGING (MRI) OF LIVER AND BILIARY TRACT WITH CONTRAST
C2315791|T060|432633002|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF LIVER AND BILIARY TRACT WITH CONTRAST|MAGNETIC RESONANCE IMAGING (MRI) OF LIVER AND BILIARY TRACT WITH CONTRAST
C2315791|T060|432633002|SNOMEDCT_US|MRI OF LIVER AND BILIARY TRACT WITH CONTRAST|MAGNETIC RESONANCE IMAGING (MRI) OF LIVER AND BILIARY TRACT WITH CONTRAST
C0882015|T060||SNOMEDCT_US|LIVER+DIAPHRAGM US
C0882015|T060||SNOMEDCT_US|LIVER AND DIAPHRAGM US
C0882015|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:LIVER+DIAPHRAGM:DOC:US
C0882015|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:LIVER+DIAPHRAGM:DOCUMENT:ULTRASOUND
C0881774|T060||SNOMEDCT_US|ABDOMEN RUQ US
C0881774|T060||SNOMEDCT_US|ABD.RUQ US
C0881774|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMEN.RUQ:DOC:US
C0881774|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMEN.RUQ:DOCUMENT:ULTRASOUND
C0881797|T060||SNOMEDCT_US|ABDOMEN US
C0881797|T060||SNOMEDCT_US|ABD US
C0881797|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMEN:DOC:US
C0881797|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:ULTRASOUND
C1543530|T060||SNOMEDCT_US|LIVER TRANSPLANT US
C1543530|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:LIVER TRANSPLANT:DOCUMENT:ULTRASOUND
C1543530|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:LIVER TRANSPLANT:DOC:US
C0944197|T060||SNOMEDCT_US|LIVER US
C0944197|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:LIVER:DOC:US
C0944197|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:LIVER:DOCUMENT:ULTRASOUND
C1543491|T060||SNOMEDCT_US|GASTROINTESTINE US
C1543491|T060||SNOMEDCT_US|GI US
C1543491|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:GASTROINTESTINE:DOC:US
C1543491|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:GASTROINTESTINE:DOCUMENT:ULTRASOUND
C1114937|T060||SNOMEDCT_US|LIVER US DURING SURGERY
C1114937|T060||SNOMEDCT_US|LIVER US IN SURG
C1114937|T060||SNOMEDCT_US|MULTISECTION^DURING SURGERY:FIND:PT:LIVER:DOC:US
C1114937|T060||SNOMEDCT_US|MULTISECTION^DURING SURGERY:FINDING:POINT IN TIME:LIVER:DOCUMENT:ULTRASOUND
C1114520|T060||SNOMEDCT_US|ABD US LTD
C1114520|T060||SNOMEDCT_US|ABDOMEN US LIMITED
C1114520|T060||SNOMEDCT_US|MULTISECTION LIMITED:FIND:PT:ABDOMEN:DOC:US
C1114520|T060||SNOMEDCT_US|MULTISECTION LIMITED:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:ULTRASOUND
C0412534|T060|241470004|SNOMEDCT_US|ULTRASOUND ABDOMINAL LIVER|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|ABDOMINAL ULTRASOUND LIVER|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|ULTRASOUND LIVER|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|HEPATIC ULTRASOUND|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|LIVER ULTRASOUND|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|ULTRASOUND OF ABDOMEN: APPEARANCE OF LIVER |US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|ULTRASOUND OF ABDOMEN: APPEARANCE OF LIVER|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|US SCAN OF LIVER|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|US SCAN OF LIVER |US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|LUSS - ULTRASOUND SCAN OF LIVER|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|ULTRASONOGRAPHY OF LIVER|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|LIVER US SCAN|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|ULTRASONOGRAPHY OF LIVER |US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|ULTRASOUND OF THE LIVER|US SCAN OF LIVER (PROCEDURE)
C0412534|T060|241470004|SNOMEDCT_US|ULTRASOUND;LIVER|US SCAN OF LIVER (PROCEDURE)
C0411889|T060|168766006|SNOMEDCT_US|LIVER SOFT TISSUE X-RAY|LIVER SOFT TISSUE X-RAY (PROCEDURE)
C0411889|T060|168766006|SNOMEDCT_US|LIVER SOFT TISSUE X-RAY |LIVER SOFT TISSUE X-RAY (PROCEDURE)
C2923070|T060||SNOMEDCT_US|ABDOMEN MRCP WO CONTRAST
C2923070|T060||SNOMEDCT_US|ABD MRCP WO CONTR
C2923070|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^WO CONTRAST:FIND:PT:LIVER+BILIARY DUCTS+PANCREAS:DOC:MRI
C2923070|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^WO CONTRAST:FINDING:POINT IN TIME:LIVER+BILIARY DUCTS+PANCREAS:DOCUMENT:MRI
C3533798|T060||SNOMEDCT_US|ABDOMEN MRCP WITH AND WITHOUT CONTRAST IV
C3533798|T060||SNOMEDCT_US|ABD MRCP W+WO CONTR IV
C3533798|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^WO & W CONTRAST IV:FIND:PT:LIVER+BILIARY DUCTS+PANCREAS:DOC:MRI
C3533798|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:LIVER+BILIARY DUCTS+PANCREAS:DOCUMENT:MRI
C0203761|T060|54780008|SNOMEDCT_US|LIVER IMAGING WITH VASCULAR FLOW|LIVER IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203767|T060|81391006|SNOMEDCT_US|LIVER AND SPLEEN IMAGING WITH VASCULAR FLOW|LIVER AND SPLEEN IMAGING WITH VASCULAR FLOW (PROCEDURE)
C2123630|T060||SNOMEDCT_US|ABDOMINAL CT LIVER NONSPECIFIC ABNORMALITY
C2123630|T060||SNOMEDCT_US|CT OF ABDOMEN NONSPECIFIC ABNORMALITY OF LIVER
C2123630|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: APPEARANCE OF NONSPECIFIC ABNORMALITY OF LIVER
C2123630|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: APPEARANCE OF NONSPECIFIC ABNORMALITY OF LIVER 
C2220596|T060||SNOMEDCT_US|ABDOMINAL COMPUTED TOMOGRAPHY LIVER MASS LESION
C2220596|T060||SNOMEDCT_US|CT SCAN OF LIVER: MASS LESION
C2220596|T060||SNOMEDCT_US|ABDOMINAL CT LIVER MASS LESION
C2220596|T060||SNOMEDCT_US|CT SCAN OF LIVER MASS LESION
C2220596|T060||SNOMEDCT_US|CT SCAN OF LIVER: MASS LESION 
C2220584|T060||SNOMEDCT_US|CT OF ABDOMEN LIVER CYST
C2220584|T060||SNOMEDCT_US|ABDOMINAL CT LIVER CYST
C2220584|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: LIVER CYST
C2220584|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: LIVER CYST 
C2220588|T060||SNOMEDCT_US|CT OF ABDOMEN DIFFUSE ENLARGEMENT OF LIVER
C2220588|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: DIFFUSE ENLARGEMENT OF LIVER
C2220588|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: DIFFUSE ENLARGEMENT OF LIVER 
C2220590|T060||SNOMEDCT_US|CT OF ABDOMEN FOCAL ENLARGEMENT OF LIVER
C2220590|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: FOCAL ENLARGEMENT OF LIVER 
C2220590|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: FOCAL ENLARGEMENT OF LIVER
C2220583|T060||SNOMEDCT_US|CT OF ABDOMEN CALCIFICATION OF LIVER
C2220583|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: CALCIFICATION OF LIVER 
C2220583|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: CALCIFICATION OF LIVER
C2021976|T060||SNOMEDCT_US|ABDOMINAL COMPUTED TOMOGRAPHY SCAN LIVER FIBROTIC CHANGES
C2021976|T060||SNOMEDCT_US|ABDOMINAL CT FIBROTIC CHANGES IN LIVER
C2021976|T060||SNOMEDCT_US|CT OF ABDOMEN FIBROTIC CHANGES IN LIVER
C2021976|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: FIBROTIC CHANGES IN LIVER 
C2021976|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: FIBROTIC CHANGES IN LIVER
C2021977|T060||SNOMEDCT_US|ABDOMINAL CT LIVER REGENERATING NODULES
C2021977|T060||SNOMEDCT_US|CT OF ABDOMEN REGENERATING NODULES OF LIVER
C2021977|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: REGENERATING NODULES OF LIVER
C2021977|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: REGENERATING NODULES OF LIVER 
C2021978|T060||SNOMEDCT_US|CT OF ABDOMEN SHRUNKEN LIVER
C2021978|T060||SNOMEDCT_US|ABDOMINAL CT SHRUNKEN LIVER
C2021978|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: SHRUNKEN LIVER
C0476419|T060|158663005|SNOMEDCT_US|[D]ABNORMAL LIVER SCAN (CONTEXT-DEPENDENT CATEGORY)|[D]ABNORMAL LIVER SCAN (SITUATION)
C0476419|T060|158663005|SNOMEDCT_US|[D]ABNORMAL LIVER SCAN |[D]ABNORMAL LIVER SCAN (SITUATION)
C0476419|T060|158663005|SNOMEDCT_US|[D]ABNORMAL LIVER SCAN|[D]ABNORMAL LIVER SCAN (SITUATION)
C0476419|T060|158663005|SNOMEDCT_US|SCAN LIVER NOS ABNORMAL|[D]ABNORMAL LIVER SCAN (SITUATION)
C0476419|T060|158663005|SNOMEDCT_US|LIVER SCAN ABNORMAL|[D]ABNORMAL LIVER SCAN (SITUATION)
C0476419|T060|158663005|SNOMEDCT_US|LIVER SCAN NOS ABNORMAL|[D]ABNORMAL LIVER SCAN (SITUATION)
C0476419|T060|158663005|SNOMEDCT_US|ABNORMAL LIVER SCAN|[D]ABNORMAL LIVER SCAN (SITUATION)
C3648818|T060||SNOMEDCT_US|IMAGING STUDIES NONSPECIFIC ABNORMAL FINDINGS LIVER
C3648818|T060||SNOMEDCT_US|IMAGING STUDIES: NONSPECIFIC ABNORMAL FINDINGS OF LIVER
C3648818|T060||SNOMEDCT_US|NONSPECIFIC ABNORMAL IMAGING FINDINGS OF LIVER
C3648818|T060||SNOMEDCT_US|IMAGING STUDIES: NONSPECIFIC ABNORMAL FINDINGS OF LIVER 
C4076645|T060|15633881000119102|SNOMEDCT_US|ULTRASONOGRAPHY OF LIVER ABNORMAL |ULTRASONOGRAPHY OF LIVER ABNORMAL (FINDING)
C4076645|T060|15633881000119102|SNOMEDCT_US|ULTRASONOGRAPHY OF LIVER ABNORMAL|ULTRASONOGRAPHY OF LIVER ABNORMAL (FINDING)
C2227710|T060||SNOMEDCT_US|ABDOMINAL X-RAY, AP VIEW: BILIARY CALCIFICATION
C2227710|T060||SNOMEDCT_US|ABDOMINAL X-RAY, AP VIEW: BILIARY CALCIFICATION 
C0495790|T060|274527008|SNOMEDCT_US|ABNORMAL FINDINGS ON DIAGNOSTIC IMAGING OF LIVER AND BILIARY TRACT|ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER+BILIARY TRACT (FINDING)
C0495790|T060|274527008|SNOMEDCT_US|ABNORMAL FINDINGS ON DX IMAGING OF LIVER AND BILIARY TRACT|ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER+BILIARY TRACT (FINDING)
C0495790|T060|274527008|SNOMEDCT_US|ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER AND BILIARY TRACT|ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER+BILIARY TRACT (FINDING)
C0495790|T060|274527008|SNOMEDCT_US|ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER+BILIARY TRACT|ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER+BILIARY TRACT (FINDING)
C0495790|T060|274527008|SNOMEDCT_US|ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER+BILIARY TRACT |ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER+BILIARY TRACT (FINDING)
C0495790|T060|274527008|SNOMEDCT_US|ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER AND BILIARY TRACT |ABNORMAL FINDINGS DIAGNOSTIC IMAGING OF LIVER+BILIARY TRACT (FINDING)
C1385723|T060||SNOMEDCT_US|DIAGNOSTIC IMAGING; ABNORMAL, BILE DUCTS (COMMON) (HEPATIC)
C1385723|T060||SNOMEDCT_US|ABNORMAL; DIAGNOSTIC IMAGING, BILE DUCTS (COMMON) (HEPATIC)
C1385728|T060||SNOMEDCT_US|DIAGNOSTIC IMAGING; ABNORMAL, LIVER
C1385728|T060||SNOMEDCT_US|ABNORMAL; DIAGNOSTIC IMAGING, LIVER
C2047961|T060||SNOMEDCT_US|IMAGING STUDIES: NONSPECIFIC ABNORMAL FINDING OF BILIARY TRACT 
C2047961|T060||SNOMEDCT_US|IMAGING STUDIES: NONSPECIFIC ABNORMAL FINDING OF BILIARY TRACT
C2711639|T060|442086001|SNOMEDCT_US|MRI OF HEART AND LIVER FOR ASSESSMENT OF CARDIAC AND HEPATIC IRON LOAD|MAGNETIC RESONANCE IMAGING OF HEART AND LIVER FOR ASSESSMENT OF CARDIAC AND HEPATIC IRON LOAD (PROCEDURE)
C2733010|T060|443637005|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF HAEMANGIOMA OF LIVER|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER (PROCEDURE)
C2733010|T060|443637005|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER |SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER (PROCEDURE)
C2733010|T060|443637005|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER (PROCEDURE)
C2733442|T060|443638000|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF LIVER AND SPLEEN|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF LIVER AND SPLEEN (PROCEDURE)
C2733442|T060|443638000|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF LIVER AND SPLEEN |SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY WITH COMPUTED TOMOGRAPHY OF LIVER AND SPLEEN (PROCEDURE)
C2220587|T060||SNOMEDCT_US|ABDOMINAL CT LIVER DENSITY (HU)
C2220587|T060||SNOMEDCT_US|CT OF ABDOMEN LIVER DENSITY (HU)
C2220587|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: LIVER DENSITY (HU) 
C2220587|T060||SNOMEDCT_US|COMPUTED TOMOGRAPHY OF ABDOMEN: LIVER DENSITY (HU)
C1830072|T060||SNOMEDCT_US|LIVER SPECT BLOOD POOL
C1830072|T060||SNOMEDCT_US|LIVER SPECT BP W RNC IV
C1830072|T060||SNOMEDCT_US|MULTISECTION BLOOD POOL^W RADIONUCLIDE IV:FIND:PT:LIVER:DOC:RADNUC.SPECT
C1830072|T060||SNOMEDCT_US|MULTISECTION BLOOD POOL^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC.SPECT
C0882014|T060||SNOMEDCT_US|LIVER SPECT W TC99MIV
C0882014|T060||SNOMEDCT_US|LIVER SPECT W TC-99M IV
C0882014|T060||SNOMEDCT_US|MULTISECTION^W TC-99M IV:FIND:PT:LIVER:DOC:RADNUC.SPECT
C0882014|T060||SNOMEDCT_US|MULTISECTION^W TC-99M INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC.SPECT
C0203758|T060|386552000|SNOMEDCT_US|RADIOISOTOPE FUNCTION STUDY OF LIVER|RADIOISOTOPE STUDY OF LIVER
C0203759|T060|169147005|SNOMEDCT_US|ISOTOPE STATIC SCAN LIVE|ISOTOPE STATIC SCAN LIVER (PROCEDURE)
C0589338|T060|271460007|SNOMEDCT_US|DYNAMIC NON-IMAGING ISOTOPE STUDY: LIVER|DYNAMIC NON-IMAGING ISOTOPE STUDY: LIVER (PROCEDURE)
C1543919|T060||SNOMEDCT_US|LIVER+LUNG RI W RNC IV
C1543919|T060||SNOMEDCT_US|LIVER AND LUNG SCAN
C1543919|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE IV:FIND:PT:LIVER+LUNG:DOC:RADNUC
C1543919|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER+LUNG:DOCUMENT:RADNUC
C1715023|T060||SNOMEDCT_US|LIVER+BDS+GB RI W SINC+RNC IV
C1715023|T060||SNOMEDCT_US|LIVER AND BILIARY DUCTS AND GALLBLADDER SCAN W SINCALIDE AND W RADIONUCLIDE IV
C1715023|T060||SNOMEDCT_US|VIEWS^W SINCALIDE & W RADIONUCLIDE IV:FIND:PT:LIVER+BILIARY DUCTS+GALLBLADDER:DOC:RADNUC
C1715023|T060||SNOMEDCT_US|VIEWS^W SINCALIDE & W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER+BILIARY DUCTS+GALLBLADDER:DOCUMENT:RADNUC
C1543899|T060||SNOMEDCT_US|LIVER+SPLEEN RI W RNC IV
C1543899|T060||SNOMEDCT_US|LIVER AND SPLEEN SCAN
C1543899|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE IV:FIND:PT:LIVER+SPLEEN:DOC:RADNUC
C1543899|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER+SPLEEN:DOCUMENT:RADNUC
C1543900|T060||SNOMEDCT_US|LIVER+SPLEEN RI STATIC W RNC IV
C1543900|T060||SNOMEDCT_US|LIVER AND SPLEEN SCAN STATIC
C1543900|T060||SNOMEDCT_US|VIEWS STATIC^W RADIONUCLIDE IV:FIND:PT:LIVER+SPLEEN:DOC:RADNUC
C1543900|T060||SNOMEDCT_US|VIEWS STATIC^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER+SPLEEN:DOCUMENT:RADNUC
C1717314|T060||SNOMEDCT_US|LIVER RI W 133XE IH
C1717314|T060||SNOMEDCT_US|VIEWS^W XE-133 IH:FIND:PT:LIVER:DOC:RADNUC
C1717314|T060||SNOMEDCT_US|VIEWS^W XE-133 INHALATION:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC
C1717314|T060||SNOMEDCT_US|LIVER SCAN W XE-133 IH
C1715027|T060||SNOMEDCT_US|LIVER SPECT FLOW W RNC IV
C1715027|T060||SNOMEDCT_US|LIVER SPECT FLOW
C1715027|T060||SNOMEDCT_US|MULTISECTION FLOW^W RADIONUCLIDE IV:FIND:PT:LIVER:DOC:RADNUC.SPECT
C1715027|T060||SNOMEDCT_US|MULTISECTION FLOW^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC.SPECT
C1652987|T060||SNOMEDCT_US|LIVER SCAN BLOOD POOL
C1652987|T060||SNOMEDCT_US|LIVER RI BP W RNC IV
C1652987|T060||SNOMEDCT_US|VIEWS BLOOD POOL^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC
C1652987|T060||SNOMEDCT_US|VIEWS BLOOD POOL^W RADIONUCLIDE IV:FIND:PT:LIVER:DOC:RADNUC
C0882016|T060||SNOMEDCT_US|LIVER+SPLEEN RI W TC99MCA COLLOID IV
C0882016|T060||SNOMEDCT_US|LIVER AND SPLEEN SCAN W TC-99M CALCIUM COLLOID IV
C0882016|T060||SNOMEDCT_US|VIEWS^W TC-99M CALCIUM COLLOID IV:FIND:PT:LIVER+SPLEEN:DOC:RADNUC
C0882016|T060||SNOMEDCT_US|VIEWS^W TC-99M CALCIUM COLLOID INTRAVENOUS:FINDING:POINT IN TIME:LIVER+SPLEEN:DOCUMENT:RADNUC
C1765325|T060||SNOMEDCT_US|LIVER RI W TC99MRBC IV
C1765325|T060||SNOMEDCT_US|LIVER SCAN W TC-99M TAGGED RBC IV
C1765325|T060||SNOMEDCT_US|VIEWS^W TC-99M TAGGED RBC IV:FIND:PT:LIVER:DOC:RADNUC
C1765325|T060||SNOMEDCT_US|VIEWS^W TC-99M TAGGED RBC INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC
C1543744|T060||SNOMEDCT_US|LIVER SPECT
C1543744|T060||SNOMEDCT_US|LIVER SPECT W RNC IV
C1543744|T060||SNOMEDCT_US|MULTISECTION^W RADIONUCLIDE IV:FIND:PT:LIVER:DOC:RADNUC.SPECT
C1543744|T060||SNOMEDCT_US|MULTISECTION^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC.SPECT
C1543790|T060||SNOMEDCT_US|ABD RI W IN-111 SATMB IV
C1543790|T060||SNOMEDCT_US|ABDOMEN SCAN W IN-111 SATUMOMAB IV
C1543790|T060||SNOMEDCT_US|VIEWS^W IN-111 SATUMOMAB INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:RADNUC
C1543790|T060||SNOMEDCT_US|VIEWS^W IN-111 SATUMOMAB IV:FIND:PT:ABDOMEN:DOC:RADNUC
C1543876|T060||SNOMEDCT_US|RI W IN-111 SATMB IV
C1543876|T060||SNOMEDCT_US|SCAN W IN-111 SATUMOMAB IV
C1543876|T060||SNOMEDCT_US|VIEWS^W IN-111 SATUMOMAB INTRAVENOUS:FINDING:POINT IN TIME:^PATIENT:DOCUMENT:RADNUC
C1543876|T060||SNOMEDCT_US|VIEWS^W IN-111 SATUMOMAB IV:FIND:PT:^PATIENT:DOC:RADNUC
C1715024|T060||SNOMEDCT_US|LIVER+SPLEEN SPECT FLOW W RNC IV
C1715024|T060||SNOMEDCT_US|LIVER AND SPLEEN SPECT FLOW
C1715024|T060||SNOMEDCT_US|MULTISECTION FLOW^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER+SPLEEN:DOCUMENT:RADNUC.SPECT
C1715024|T060||SNOMEDCT_US|MULTISECTION FLOW^W RADIONUCLIDE IV:FIND:PT:LIVER+SPLEEN:DOC:RADNUC.SPECT
C1543743|T060||SNOMEDCT_US|LIVER SPECT W TC99MRBC IV
C1543743|T060||SNOMEDCT_US|LIVER SPECT W TC-99M TAGGED RBC IV
C1543743|T060||SNOMEDCT_US|MULTISECTION^W TC-99M TAGGED RBC IV:FIND:PT:LIVER:DOC:RADNUC.SPECT
C1543743|T060||SNOMEDCT_US|MULTISECTION^W TC-99M TAGGED RBC INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC.SPECT
C1543745|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER:NARRATIVE:RADNUC
C1543745|T060||SNOMEDCT_US|LIVER RI W RNC IV
C1543745|T060||SNOMEDCT_US|LIVER SCAN
C1543745|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE IV:FIND:PT:LIVER:DOC:RADNUC
C1543745|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC
C1543874|T060||SNOMEDCT_US|LIVER SCAN STATIC
C1543874|T060||SNOMEDCT_US|LIVER RI STATIC W RNC IV
C1543874|T060||SNOMEDCT_US|VIEWS STATIC^W RADIONUCLIDE IV:FIND:PT:LIVER:DOC:RADNUC
C1543874|T060||SNOMEDCT_US|VIEWS STATIC^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC
C1543746|T060||SNOMEDCT_US|LIVER TRANSPLANT SCAN
C1543746|T060||SNOMEDCT_US|LIVER TRANSPLANT RI W RNC IV
C1543746|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER TRANSPLANT:DOCUMENT:RADNUC
C1543746|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE IV:FIND:PT:LIVER TRANSPLANT:DOC:RADNUC
C1543898|T060||SNOMEDCT_US|LIVER+SPLEEN SPECT W RNC IV
C1543898|T060||SNOMEDCT_US|LIVER AND SPLEEN SPECT
C1543898|T060||SNOMEDCT_US|MULTISECTION^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER+SPLEEN:DOCUMENT:RADNUC.SPECT
C1543898|T060||SNOMEDCT_US|MULTISECTION^W RADIONUCLIDE IV:FIND:PT:LIVER+SPLEEN:DOC:RADNUC.SPECT
C1715025|T060||SNOMEDCT_US|LIVER+SPLEEN RI FLOW W RNC IV
C1715025|T060||SNOMEDCT_US|LIVER AND SPLEEN SCAN FLOW
C1715025|T060||SNOMEDCT_US|VIEWS FLOW^W RADIONUCLIDE IV:FIND:PT:LIVER+SPLEEN:DOC:RADNUC
C1715025|T060||SNOMEDCT_US|VIEWS FLOW^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER+SPLEEN:DOCUMENT:RADNUC
C3263042|T060||SNOMEDCT_US|LIVER SPECT W TC99MSC IV
C3263042|T060||SNOMEDCT_US|LIVER SPECT W TC-99M SC IV
C3263042|T060||SNOMEDCT_US|MULTISECTION^W TC-99M SUBCUTANEOUS INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC.SPECT
C3263042|T060||SNOMEDCT_US|MULTISECTION^W TC-99M SC IV:FIND:PT:LIVER:DOC:RADNUC.SPECT
C1715411|T060||SNOMEDCT_US|LIVER+SPLEEN RI W TC99MMAA IV
C1715411|T060||SNOMEDCT_US|LIVER AND SPLEEN SCAN W TC-99M MAA IV
C1715411|T060||SNOMEDCT_US|VIEWS^W TC-99M MAA INTRAVENOUS:FINDING:POINT IN TIME:LIVER+SPLEEN:DOCUMENT:RADNUC
C1715411|T060||SNOMEDCT_US|VIEWS^W TC-99M MAA IV:FIND:PT:LIVER+SPLEEN:DOC:RADNUC
C1714946|T060||SNOMEDCT_US|LIVER+BDS+GB RI W RNC IV
C1714946|T060||SNOMEDCT_US|LIVER AND BILIARY DUCTS AND GALLBLADDER SCAN
C1714946|T060||SNOMEDCT_US|VIEWS^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER+BILIARY DUCTS+GALLBLADDER:DOCUMENT:RADNUC
C3263043|T060||SNOMEDCT_US|LIVER SCAN W TC-99M SC IV
C3263043|T060||SNOMEDCT_US|LIVER RI W TC99MSC IV
C3263043|T060||SNOMEDCT_US|VIEWS^W TC-99M SUBCUTANEOUS INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC
C3263043|T060||SNOMEDCT_US|VIEWS^W TC-99M SC IV:FIND:PT:LIVER:DOC:RADNUC
C4036766|T060||SNOMEDCT_US|LIVER STIFFNESS BY US.TRANSIENT ELASTOGRAPHY
C4036766|T060||SNOMEDCT_US|LIVER STIFFNESS:PRESSURE:POINT IN TIME:LIVER:QUANTITATIVE:ULTRASOUND.TRANSIENT ELASTOGRAPHY
C4036766|T060||SNOMEDCT_US|LIVER STIFFNESS US.TE
C4036766|T060||SNOMEDCT_US|LIVER STIFFNESS:PRES:PT:LIVER:QN:US.TRANSIENT ELASTOGRAPHY
C0412760|T060|169258005|SNOMEDCT_US|THERMOGRAPHY - HEPATIC REGION |THERMOGRAPHY - HEPATIC REGION (PROCEDURE)
C0412760|T060|169258005|SNOMEDCT_US|THERMOGRAPHY - HEPATIC REGION|THERMOGRAPHY - HEPATIC REGION (PROCEDURE)
C0203758|T060|386552000|SNOMEDCT_US|RADIOISOTOPE FUNCTION STUDY OF LIVER|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|LIVER SCAN/ISOTOPE FUNCT|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|LIVER IMAGING|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|RADIOISOTOPE FUNCTION STUDY OF LIVER |RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|RADIONUCLIDE HEPATIC FUNCTION STUDY|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|LIVER SCAN|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|RADIONUCLIDE LIVER STUDIES|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|LIVER ISOTOPE STUDIES|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|LIVER SCAN NOS|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|SCAN LIVER NOS|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|RADIOISOTOPE STUDY OF LIVER |RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|RADIOISOTOPE STUDY OF LIVER|RADIOISOTOPE STUDY OF LIVER
C0203758|T060|386552000|SNOMEDCT_US|LIVER SCAN AND RADIOISOTOPE FUNCTION STUDY|RADIOISOTOPE STUDY OF LIVER
C2316126|T060|431948007|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY (SPECT) OF HEMANGIOMA OF LIVER|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER (PROCEDURE)
C2316126|T060|431948007|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER (PROCEDURE)
C2316126|T060|431948007|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF HAEMANGIOMA OF LIVER|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER (PROCEDURE)
C2316126|T060|431948007|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER |SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER (PROCEDURE)
C2316126|T060|431948007|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY (SPECT) OF HAEMANGIOMA OF LIVER|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF HEMANGIOMA OF LIVER (PROCEDURE)
C0203759|T060|169147005|SNOMEDCT_US|ISOTOPE STATIC SCAN LIVER |ISOTOPE STATIC SCAN LIVER (PROCEDURE)
C2315171|T060|429791001|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF LIVER AND SPLEEN|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY (SPECT) OF LIVER AND SPLEEN
C2315171|T060|429791001|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY OF LIVER AND SPLEEN |SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY (SPECT) OF LIVER AND SPLEEN
C2315171|T060|429791001|SNOMEDCT_US|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY (SPECT) OF LIVER AND SPLEEN|SINGLE PHOTON EMISSION COMPUTED TOMOGRAPHY (SPECT) OF LIVER AND SPLEEN
C0473930|T060|241346004|SNOMEDCT_US|TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - DYNAMIC |TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - DYNAMIC (PROCEDURE)
C0473930|T060|241346004|SNOMEDCT_US|TC99M-LABELLED COLLOID LIVER AND SPLEEN STUDY - DYNAMIC |TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - DYNAMIC (PROCEDURE)
C0473930|T060|241346004|SNOMEDCT_US|TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - DYNAMIC|TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - DYNAMIC (PROCEDURE)
C0473930|T060|241346004|SNOMEDCT_US|TC99M-LABELLED COLLOID LIVER AND SPLEEN STUDY - DYNAMIC|TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - DYNAMIC (PROCEDURE)
C0412394|T060|241341009|SNOMEDCT_US|RADIONUCLIDE STUDY OF LIVER, SPLEEN AND BILIARY TRACT|RADIONUCLIDE STUDY OF LIVER, SPLEEN AND BILIARY TRACT (PROCEDURE)
C0412394|T060|241341009|SNOMEDCT_US|RADIONUCLIDE STUDY OF LIVER, SPLEEN AND BILIARY TRACT |RADIONUCLIDE STUDY OF LIVER, SPLEEN AND BILIARY TRACT (PROCEDURE)
C0473931|T060|241350006|SNOMEDCT_US|TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - STATIC |TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - STATIC (PROCEDURE)
C0473931|T060|241350006|SNOMEDCT_US|TC99M-LABELLED COLLOID LIVER AND SPLEEN STUDY - STATIC|TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - STATIC (PROCEDURE)
C0473931|T060|241350006|SNOMEDCT_US|TC99M-LABELLED COLLOID LIVER AND SPLEEN STUDY - STATIC |TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - STATIC (PROCEDURE)
C0473931|T060|241350006|SNOMEDCT_US|TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - STATIC|TC99M-LABELED COLLOID LIVER AND SPLEEN STUDY - STATIC (PROCEDURE)
C1644183|T060|418234000|SNOMEDCT_US|RADIONUCLIDE LIVER AND SPLEEN IMAGING PROCEDURE |RADIONUCLIDE LIVER AND SPLEEN IMAGING PROCEDURE
C1644183|T060|418234000|SNOMEDCT_US|RADIONUCLIDE LIVER AND SPLEEN IMAGING PROCEDURE|RADIONUCLIDE LIVER AND SPLEEN IMAGING PROCEDURE
C1644183|T060|418234000|SNOMEDCT_US|RADIONUCLIDE LIVER AND SPLEEN STUDY|RADIONUCLIDE LIVER AND SPLEEN IMAGING PROCEDURE
C2585276|T060|440204002|SNOMEDCT_US|RADIONUCLIDE STUDY OF PERFUSION OF LIVER|RADIONUCLIDE STUDY OF PERFUSION OF LIVER (PROCEDURE)
C2585276|T060|440204002|SNOMEDCT_US|RADIONUCLIDE STUDY OF PERFUSION OF LIVER |RADIONUCLIDE STUDY OF PERFUSION OF LIVER (PROCEDURE)
C2108323|T060||SNOMEDCT_US|RADIOISOTOPE SCAN OF LIVER 
C2108323|T060||SNOMEDCT_US|RADIOISOTOPE SCAN OF LIVER
C2054285|T060||SNOMEDCT_US|TECHNETIUM SCAN OF LIVER 
C2054285|T060||SNOMEDCT_US|TECHNETIUM SCAN OF LIVER
C0412396|T060|169164008|SNOMEDCT_US|ISOTOPE DYNAMIC LIVER SCAN |ISOTOPE DYNAMIC LIVER SCAN (PROCEDURE)
C0412396|T060|169164008|SNOMEDCT_US|ISOTOPE DYNAMIC LIVER SCAN|ISOTOPE DYNAMIC LIVER SCAN (PROCEDURE)
C0203760|T060|45588000|SNOMEDCT_US|LIVER FUNCTION STUDY WITH SERIAL IMAGES|LIVER FUNCTION STUDY WITH SERIAL IMAGES (PROCEDURE)
C0203760|T060|45588000|SNOMEDCT_US|LIVER FUNCTION STUDY WITH SERIAL IMAGES |LIVER FUNCTION STUDY WITH SERIAL IMAGES (PROCEDURE)
C0589338|T060|271460007|SNOMEDCT_US|DYNAMIC NON-IMAGING ISOTOPE: LIVER (& [STUDY]) |DYNAMIC NON-IMAGING ISOTOPE STUDY: LIVER (PROCEDURE)
C0589338|T060|271460007|SNOMEDCT_US|DYNAMIC NON-IMAGING ISOTOPE: LIVER (& [STUDY])|DYNAMIC NON-IMAGING ISOTOPE STUDY: LIVER (PROCEDURE)
C0589338|T060|271460007|SNOMEDCT_US|DYNAMIC NON-IMAGING ISOTOPE STUDY: LIVER |DYNAMIC NON-IMAGING ISOTOPE STUDY: LIVER (PROCEDURE)
C0589338|T060|271460007|SNOMEDCT_US|DYNAMIC NON-IMAGING ISOTOPE STUDY: LIVER|DYNAMIC NON-IMAGING ISOTOPE STUDY: LIVER (PROCEDURE)
C0589338|T060|271460007|SNOMEDCT_US|DYNAM.NON-IM.ISOTOPE: LIVER|DYNAMIC NON-IMAGING ISOTOPE STUDY: LIVER (PROCEDURE)
C0581583|T060|303866009|SNOMEDCT_US|TC99M-LABELLED COLLOID LIVER STUDY - DYNAMIC|TC99M-LABELED COLLOID LIVER STUDY - DYNAMIC (PROCEDURE)
C0581583|T060|303866009|SNOMEDCT_US|TC99M-LABELED COLLOID LIVER STUDY - DYNAMIC|TC99M-LABELED COLLOID LIVER STUDY - DYNAMIC (PROCEDURE)
C0581583|T060|303866009|SNOMEDCT_US|TC99M-LABELED COLLOID LIVER STUDY - DYNAMIC |TC99M-LABELED COLLOID LIVER STUDY - DYNAMIC (PROCEDURE)
C0581583|T060|303866009|SNOMEDCT_US|TC99M-LABELLED COLLOID LIVER STUDY - DYNAMIC |TC99M-LABELED COLLOID LIVER STUDY - DYNAMIC (PROCEDURE)
C0581584|T060|303867000|SNOMEDCT_US|TC99M-LABELED COLLOID LIVER STUDY - STATIC|TC99M-LABELED COLLOID LIVER STUDY - STATIC (PROCEDURE)
C0581584|T060|303867000|SNOMEDCT_US|TC99M-LABELLED COLLOID LIVER STUDY - STATIC|TC99M-LABELED COLLOID LIVER STUDY - STATIC (PROCEDURE)
C0581584|T060|303867000|SNOMEDCT_US|TC99M-LABELLED COLLOID LIVER STUDY - STATIC |TC99M-LABELED COLLOID LIVER STUDY - STATIC (PROCEDURE)
C0581584|T060|303867000|SNOMEDCT_US|TC99M-LABELED COLLOID LIVER STUDY - STATIC |TC99M-LABELED COLLOID LIVER STUDY - STATIC (PROCEDURE)
C0203764|T060|113125002|SNOMEDCT_US|RADIOLABELED ROSE BENGAL STUDY|RADIOIODINATED ROSE BENGAL STUDY OF LIVER (PROCEDURE)
C0203764|T060|113125002|SNOMEDCT_US|RADIOIODINATED ROSE BENGAL STUDY OF LIVER|RADIOIODINATED ROSE BENGAL STUDY OF LIVER (PROCEDURE)
C0203764|T060|113125002|SNOMEDCT_US|RADIOLABELLED ROSE BENGAL STUDY|RADIOIODINATED ROSE BENGAL STUDY OF LIVER (PROCEDURE)
C0203764|T060|113125002|SNOMEDCT_US|RADIOIODINATED ROSE BENGAL STUDY OF LIVER |RADIOIODINATED ROSE BENGAL STUDY OF LIVER (PROCEDURE)
C2094547|T060||SNOMEDCT_US|RADIONUCLIDE SCAN OF LIVER AND SPLEEN WITH VASCULAR FLOW 
C2094547|T060||SNOMEDCT_US|RADIONUCLIDE SCAN OF LIVER AND SPLEEN WITH VASCULAR FLOW
C2711639|T060|442086001|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF HEART AND LIVER FOR ASSESSMENT OF CARDIAC AND HEPATIC IRON LOAD |MAGNETIC RESONANCE IMAGING OF HEART AND LIVER FOR ASSESSMENT OF CARDIAC AND HEPATIC IRON LOAD (PROCEDURE)
C2711639|T060|442086001|SNOMEDCT_US|MAGNETIC RESONANCE IMAGING OF HEART AND LIVER FOR ASSESSMENT OF CARDIAC AND HEPATIC IRON LOAD|MAGNETIC RESONANCE IMAGING OF HEART AND LIVER FOR ASSESSMENT OF CARDIAC AND HEPATIC IRON LOAD (PROCEDURE)
C2711639|T060|442086001|SNOMEDCT_US|MRI OF HEART AND LIVER FOR ASSESSMENT OF CARDIAC AND HEPATIC IRON LOAD|MAGNETIC RESONANCE IMAGING OF HEART AND LIVER FOR ASSESSMENT OF CARDIAC AND HEPATIC IRON LOAD (PROCEDURE)
C2094545|T060||SNOMEDCT_US|RADIONUCLIDE SCAN OF LIVER AND SPLEEN 
C2094545|T060||SNOMEDCT_US|RADIONUCLIDE SCAN OF LIVER AND SPLEEN
C2094546|T060||SNOMEDCT_US|STATIC RADIONUCLIDE SCAN OF LIVER AND SPLEEN 
C2094546|T060||SNOMEDCT_US|STATIC RADIONUCLIDE SCAN OF LIVER AND SPLEEN
C0881804|T060||SNOMEDCT_US|VIEWS AP (KUB & UPRIGHT) & UPRIGHT CHEST:FINDING:POINT IN TIME:CHEST+ABDOMEN:NARRATIVE:XR
C0881804|T060||SNOMEDCT_US|DEPRECATED CHEST+ABD XR
C0881804|T060||SNOMEDCT_US|VIEWS AP (KUB & UPRIGHT) & UPRIGHT CHEST:FIND:PT:CHEST+ABDOMEN:NAR:XR
C0881804|T060||SNOMEDCT_US|DEPRECATED CHEST AND ABDOMEN NARRATIVE X-RAY
C1978440|T060||SNOMEDCT_US|DEPRECATED VIEWS AP & LATERAL:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C1978440|T060||SNOMEDCT_US|DEPRECATED ABD XR AP+LAT
C1978440|T060||SNOMEDCT_US|DEPRECATED ABDOMEN X-RAY AP & LATERAL
C1978440|T060||SNOMEDCT_US|VIEWS AP & LATERAL:FIND:PT:ABDOMEN:NAR:XR
C1978440|T060||SNOMEDCT_US|VIEWS AP & LATERAL:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C0881998|T060||SNOMEDCT_US|ABD XR AP (SUP+UPR)
C0881998|T060||SNOMEDCT_US|ABDOMEN X-RAY AP (SUPINE AND UPRIGHT)
C0881998|T060||SNOMEDCT_US|VIEWS AP (SUPINE & UPRIGHT):FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881998|T060||SNOMEDCT_US|VIEWS AP (SUPINE & UPRIGHT):FIND:PT:ABDOMEN:DOC:XR
C1624698|T060||SNOMEDCT_US|CHEST AND ABDOMEN X-RAY SINGLE VIEW
C1624698|T060||SNOMEDCT_US|CHEST+ABD XR 1V
C1624698|T060||SNOMEDCT_US|VIEW 1:FIND:PT:CHEST+ABDOMEN:DOC:XR
C1624698|T060||SNOMEDCT_US|VIEW 1:FINDING:POINT IN TIME:CHEST+ABDOMEN:DOCUMENT:XR
C1626841|T060||SNOMEDCT_US|DEPRECATED VIEW AP:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C1626841|T060||SNOMEDCT_US|DEPRECATED ABD XR AP 1V
C1626841|T060||SNOMEDCT_US|VIEW AP:FIND:PT:ABDOMEN:NAR:XR
C1626841|T060||SNOMEDCT_US|DEPRECATED ABDOMEN X-RAY AP
C0881997|T060||SNOMEDCT_US|ABD XR AP+OBL PRONE
C0881997|T060||SNOMEDCT_US|ABDOMEN X-RAY AP AND OBLIQUE PRONE
C0881997|T060||SNOMEDCT_US|VIEWS AP & OBLIQUE PRONE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881997|T060||SNOMEDCT_US|VIEWS AP & OBLIQUE PRONE:FIND:PT:ABDOMEN:DOC:XR
C1525954|T060||SNOMEDCT_US|ABDOMEN X-RAY
C1525954|T060||SNOMEDCT_US|ABD XR
C1525954|T060||SNOMEDCT_US|VIEWS:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C1525954|T060||SNOMEDCT_US|VIEWS:FIND:PT:ABDOMEN:DOC:XR
C1525954|T060||SNOMEDCT_US|VIEWS:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1644644|T060||SNOMEDCT_US|ABDOMEN X-RAY DURING SURGERY
C1644644|T060||SNOMEDCT_US|ABD XR IN SURG
C1644644|T060||SNOMEDCT_US|VIEW^DURING SURGERY:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1644644|T060||SNOMEDCT_US|VIEW^DURING SURGERY:FIND:PT:ABDOMEN:DOC:XR
C0881801|T060||SNOMEDCT_US|ABD XR AP (L+R LAT DECUB)
C0881801|T060||SNOMEDCT_US|ABDOMEN X-RAY AP (LEFT LATERAL-DECUBITUS AND RIGHT LATERAL-DECUBITUS)
C0881801|T060||SNOMEDCT_US|VIEWS AP (L-LATERAL-DECUBITUS & R-LATERAL-DECUBITUS):FIND:PT:ABDOMEN:DOC:XR
C0881801|T060||SNOMEDCT_US|VIEWS AP (L-LATERAL-DECUBITUS & R-LATERAL-DECUBITUS):FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C3262888|T060||SNOMEDCT_US|ABD XR AP+LAT XTABLE
C3262888|T060||SNOMEDCT_US|ABDOMEN X-RAY AP AND LATERAL CROSSTABLE
C3262888|T060||SNOMEDCT_US|VIEWS AP & LATERAL CROSSTABLE:FIND:PT:ABDOMEN:DOC:XR
C3262888|T060||SNOMEDCT_US|VIEWS AP & LATERAL CROSSTABLE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881803|T060||SNOMEDCT_US|ABDOMEN X-RAY AP UPRIGHT PORTABLE
C0881803|T060||SNOMEDCT_US|ABD XR AP UPR PORT
C0881803|T060||SNOMEDCT_US|VIEW AP UPRIGHT PORTABLE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881803|T060||SNOMEDCT_US|VIEW AP UPRIGHT PORTABLE:FIND:PT:ABDOMEN:DOC:XR
C1648947|T060||SNOMEDCT_US|DEPRECATED VIEW AP PORTABLE:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C1648947|T060||SNOMEDCT_US|DEPRECATED ABDOMEN X-RAY AP PORTABLE
C1648947|T060||SNOMEDCT_US|VIEW AP PORTABLE:FIND:PT:ABDOMEN:NAR:XR
C1648947|T060||SNOMEDCT_US|DEPRECATED ABD XR AP PORT
C1648947|T060||SNOMEDCT_US|VIEW AP PORTABLE:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C0881992|T060||SNOMEDCT_US|ABD XR AP+AP L-LAT DECUB PORT
C0881992|T060||SNOMEDCT_US|ABDOMEN X-RAY AP AND AP LEFT LATERAL-DECUBITUS PORTABLE
C0881992|T060||SNOMEDCT_US|VIEWS AP & AP L-LATERAL-DECUBITUS PORTABLE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881992|T060||SNOMEDCT_US|VIEWS AP & AP L-LATERAL-DECUBITUS PORTABLE:FIND:PT:ABDOMEN:DOC:XR
C1524218|T060||SNOMEDCT_US|VIEW AP PORTABLE:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C1524218|T060||SNOMEDCT_US|ABDOMEN X-RAY AP PORTABLE SINGLE VIEW
C1524218|T060||SNOMEDCT_US|ABD XR AP V1 PORT
C1524218|T060||SNOMEDCT_US|VIEW AP PORTABLE:FIND:PT:ABDOMEN:DOC:XR
C1524218|T060||SNOMEDCT_US|VIEW AP PORTABLE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1525327|T060||SNOMEDCT_US|ABDOMEN X-RAY LEFT LATERAL
C1525327|T060||SNOMEDCT_US|ABD XR L-LAT
C1525327|T060||SNOMEDCT_US|VIEW L-LATERAL:FIND:PT:ABDOMEN:DOC:XR
C1525327|T060||SNOMEDCT_US|VIEW L-LATERAL:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1508084|T060||SNOMEDCT_US|ABD XR AP+L-POST OBL
C1508084|T060||SNOMEDCT_US|ABDOMEN X-RAY AP AND LEFT POSTERIOR OBLIQUE
C1508084|T060||SNOMEDCT_US|VIEWS AP & L-POSTERIOR OBLIQUE:FIND:PT:ABDOMEN:DOC:XR
C1508084|T060||SNOMEDCT_US|VIEWS AP & L-POSTERIOR OBLIQUE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1525301|T060||SNOMEDCT_US|DEPRECATED VIEW DECUBITUS:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C1525301|T060||SNOMEDCT_US|VIEW DECUBITUS:FIND:PT:ABDOMEN:NAR:XR
C1525301|T060||SNOMEDCT_US|DEPRECATED ABD XR DECUBITUS
C1525301|T060||SNOMEDCT_US|VIEW DECUBITUS:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C0881799|T060||SNOMEDCT_US|ABD XR AP L-LAT DECUB PORT
C0881799|T060||SNOMEDCT_US|ABDOMEN X-RAY AP LEFT LATERAL-DECUBITUS PORTABLE
C0881799|T060||SNOMEDCT_US|VIEW AP L-LATERAL-DECUBITUS PORTABLE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881799|T060||SNOMEDCT_US|VIEW AP L-LATERAL-DECUBITUS PORTABLE:FIND:PT:ABDOMEN:DOC:XR
C1114571|T060||SNOMEDCT_US|ABD XR AP+LAT XTABLE PORT
C1114571|T060||SNOMEDCT_US|ABDOMEN X-RAY AP AND LATERAL CROSSTABLE PORTABLE
C1114571|T060||SNOMEDCT_US|VIEWS AP & LATERAL CROSSTABLE PORTABLE:FIND:PT:ABDOMEN:DOC:XR
C1114571|T060||SNOMEDCT_US|VIEWS AP & LATERAL CROSSTABLE PORTABLE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1524221|T060||SNOMEDCT_US|ABDOMEN X-RAY UPRIGHT
C1524221|T060||SNOMEDCT_US|ABD XR UPR
C1524221|T060||SNOMEDCT_US|VIEW UPRIGHT:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1524221|T060||SNOMEDCT_US|VIEW UPRIGHT:FIND:PT:ABDOMEN:DOC:XR
C1524955|T060||SNOMEDCT_US|ABD XR OBL 1V
C1524955|T060||SNOMEDCT_US|ABDOMEN X-RAY OBLIQUE SINGLE VIEW
C1524955|T060||SNOMEDCT_US|VIEW OBLIQUE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1524955|T060||SNOMEDCT_US|VIEW OBLIQUE:FIND:PT:ABDOMEN:DOC:XR
C1632257|T060||SNOMEDCT_US|ABD XR AP (UPR+L LAT DECUB)
C1632257|T060||SNOMEDCT_US|ABDOMEN X-RAY AP (UPRIGHT AND LEFT LATERAL DECUBITUS)
C1632257|T060||SNOMEDCT_US|VIEWS AP (UPRIGHT & L-LATERAL DECUBITUS):FIND:PT:ABDOMEN:DOC:XR
C1632257|T060||SNOMEDCT_US|VIEWS AP (UPRIGHT & L-LATERAL DECUBITUS):FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881999|T060||SNOMEDCT_US|VIEW AP:FINDING:POINT IN TIME:ABDOMEN:NARRATIVE:XR
C0881999|T060||SNOMEDCT_US|ABDOMEN X-RAY AP SINGLE VIEW
C0881999|T060||SNOMEDCT_US|ABD XR AP 1V
C0881999|T060||SNOMEDCT_US|VIEW AP:FIND:PT:ABDOMEN:DOC:XR
C0881999|T060||SNOMEDCT_US|VIEW AP:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1525316|T060||SNOMEDCT_US|ABD XR LAT XTABLE
C1525316|T060||SNOMEDCT_US|ABDOMEN X-RAY LATERAL CROSSTABLE
C1525316|T060||SNOMEDCT_US|VIEW LATERAL CROSSTABLE:FIND:PT:ABDOMEN:DOC:XR
C1525316|T060||SNOMEDCT_US|VIEW LATERAL CROSSTABLE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1524683|T060||SNOMEDCT_US|ABDOMEN X-RAY PA PRONE
C1524683|T060||SNOMEDCT_US|ABD XR PA PRONE
C1524683|T060||SNOMEDCT_US|VIEW PA PRONE:FIND:PT:ABDOMEN:DOC:XR
C1524683|T060||SNOMEDCT_US|VIEW PA PRONE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1525530|T060||SNOMEDCT_US|ABD XR R-LAT+L-LAT
C1525530|T060||SNOMEDCT_US|ABDOMEN X-RAY RIGHT LATERAL AND LEFT LATERAL
C1525530|T060||SNOMEDCT_US|VIEWS R-LATERAL & L-LATERAL:FIND:PT:ABDOMEN:DOC:XR
C1525530|T060||SNOMEDCT_US|VIEWS R-LATERAL & L-LATERAL:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1714950|T060||SNOMEDCT_US|CHEST AND ABDOMEN X-RAY AP UPRIGHT AND AP CHEST
C1714950|T060||SNOMEDCT_US|CHEST+ABD XR AP UPR+AP CHST
C1714950|T060||SNOMEDCT_US|VIEWS AP UPRIGHT & AP CHEST:FIND:PT:CHEST+ABDOMEN:DOC:XR
C1714950|T060||SNOMEDCT_US|VIEWS AP UPRIGHT & AP CHEST:FINDING:POINT IN TIME:CHEST+ABDOMEN:DOCUMENT:XR
C1525496|T060||SNOMEDCT_US|ABD XR AP(SUP+LAT DECUB)
C1525496|T060||SNOMEDCT_US|ABDOMEN X-RAY AP (SUPINE AND LATERAL-DECUBITUS)
C1525496|T060||SNOMEDCT_US|VIEWS AP (SUPINE & LATERAL-DECUBITUS):FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1525496|T060||SNOMEDCT_US|VIEWS AP (SUPINE & LATERAL-DECUBITUS):FIND:PT:ABDOMEN:DOC:XR
C1525519|T060||SNOMEDCT_US|ABD XR AP+OBL
C1525519|T060||SNOMEDCT_US|ABDOMEN X-RAY AP AND OBLIQUE
C1525519|T060||SNOMEDCT_US|VIEWS AP & OBLIQUE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1525519|T060||SNOMEDCT_US|VIEWS AP & OBLIQUE:FIND:PT:ABDOMEN:DOC:XR
C1524619|T060||SNOMEDCT_US|ABDOMEN X-RAY 3 VIEWS
C1524619|T060||SNOMEDCT_US|ABD XR 3V
C1524619|T060||SNOMEDCT_US|VIEWS 3:FIND:PT:ABDOMEN:DOC:XR
C1524619|T060||SNOMEDCT_US|VIEWS 3:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881996|T060||SNOMEDCT_US|ABD XR AP+AP L-LAT DECUB
C0881996|T060||SNOMEDCT_US|ABDOMEN X-RAY AP AND AP LEFT LATERAL-DECUBITUS
C0881996|T060||SNOMEDCT_US|VIEWS AP & AP L-LATERAL-DECUBITUS:FIND:PT:ABDOMEN:DOC:XR
C0881996|T060||SNOMEDCT_US|VIEWS AP & AP L-LATERAL-DECUBITUS:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881994|T060||SNOMEDCT_US|ABD XR AP+LAT
C0881994|T060||SNOMEDCT_US|ABDOMEN X-RAY AP AND LATERAL
C0881994|T060||SNOMEDCT_US|VIEWS AP & LATERAL:FIND:PT:ABDOMEN:DOC:XR
C0881994|T060||SNOMEDCT_US|VIEWS AP & LATERAL:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881995|T060||SNOMEDCT_US|ABD XR AP (SUPINE+UPR) PORT
C0881995|T060||SNOMEDCT_US|ABDOMEN X-RAY AP (SUPINE AND UPRIGHT) PORTABLE
C0881995|T060||SNOMEDCT_US|VIEWS AP (SUPINE & UPRIGHT) PORTABLE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0881995|T060||SNOMEDCT_US|VIEWS AP (SUPINE & UPRIGHT) PORTABLE:FIND:PT:ABDOMEN:DOC:XR
C0881802|T060||SNOMEDCT_US|ABD XR AP R-LAT DECUB
C0881802|T060||SNOMEDCT_US|ABDOMEN X-RAY AP RIGHT LATERAL-DECUBITUS
C0881802|T060||SNOMEDCT_US|VIEW AP R-LATERAL-DECUBITUS:FIND:PT:ABDOMEN:DOC:XR
C0881802|T060||SNOMEDCT_US|VIEW AP R-LATERAL-DECUBITUS:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1543409|T060||SNOMEDCT_US|ABD XR R-POST OBL
C1543409|T060||SNOMEDCT_US|ABDOMEN X-RAY RIGHT POSTERIOR OBLIQUE
C1543409|T060||SNOMEDCT_US|VIEW R-POSTERIOR OBLIQUE:FIND:PT:ABDOMEN:DOC:XR
C1543409|T060||SNOMEDCT_US|VIEW R-POSTERIOR OBLIQUE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1524939|T060||SNOMEDCT_US|ABDOMEN X-RAY LATERAL
C1524939|T060||SNOMEDCT_US|ABD XR LAT
C1524939|T060||SNOMEDCT_US|VIEW LATERAL:FIND:PT:ABDOMEN:DOC:XR
C1524939|T060||SNOMEDCT_US|VIEW LATERAL:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C1624108|T060||SNOMEDCT_US|CHEST+ABD XR AP+PA CHST
C1624108|T060||SNOMEDCT_US|CHEST AND ABDOMEN X-RAY AP AND PA CHEST
C1624108|T060||SNOMEDCT_US|VIEWS AP & PA CHEST:FIND:PT:CHEST+ABDOMEN:DOC:XR
C1624108|T060||SNOMEDCT_US|VIEWS AP & PA CHEST:FINDING:POINT IN TIME:CHEST+ABDOMEN:DOCUMENT:XR
C4070261|T060||SNOMEDCT_US|ABD XR GE 3V
C4070261|T060||SNOMEDCT_US|VIEWS GE 3:FIND:PT:ABDOMEN:DOC:XR
C4070261|T060||SNOMEDCT_US|ABDOMEN X-RAY GE 3 VIEWS
C4070261|T060||SNOMEDCT_US|VIEWS GE 3:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR
C0034573|T060|145931009|SNOMEDCT_US|RADIOGRAPHY, ABDOMINAL|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|ABDOMINAL RADIOGRAPHIES|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|RADIOGRAPHIES, ABDOMINAL|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|ABDOMINAL X-RAY|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|RADIOGR ABDOMINAL|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|ABDOMINAL RADIOGR|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|X-RAY OF ABDOMEN |ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|X-RAY OF ABDOMEN|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|X-RAY;ABDOMEN|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|ABDOMINAL X-RAY |ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|RADIOLOGIC EXAMINATION, ABDOMEN|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|ABDOMEN--RADIOGRAPHY|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|ABDOMINAL X-RAY NOS|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|ABDOMINAL RADIOGRAPHY|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|AXR - ABDOMINAL X-RAY|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|DIAGNOSTIC RADIOGRAPHY OF ABDOMEN |ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|DIAGNOSTIC RADIOGRAPHY OF ABDOMEN|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|RADIOLOGIC EXAMINATION OF ABDOMEN|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|RADIOLOGIC PROCEDURE ON ABDOMEN|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|RADIOLOGIC EXAMINATION OF ABDOMEN, NOS|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|X-RAY OF ABDOMEN, NOS|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|RADIOLOGIC PROCEDURE ON ABDOMEN, NOS|ABDOMINAL X-RAY (PROCEDURE)
C0034573|T060|145931009|SNOMEDCT_US|X-RAY OF THE ABDOMEN|ABDOMINAL X-RAY (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|GASTROINTESTINAL TRACT X-RAY NOS|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|DIGESTIVE TRACT X-RAY|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|GI TRACT X-RAY NOS|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|X-RAY GASTROINTESTINAL TRACT|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|X-RAY NOS GASTROINTESTINAL TRACT|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|DIGESTIVE TRACT X-RAY NOS|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|RADIOGRAPHY OF GASTROINTESTINAL TRACT|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|GASTROINTESTINAL TRACT X-RAY|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|RADIOGRAPHY OF GASTROINTESTINAL TRACT |RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|RADIOGRAPHY OF DIGESTIVE TRACT, NOS|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|GASTROINTESTINAL TRACT X-RAY, NOS|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203054|T060|75679007|SNOMEDCT_US|X-RAY OF THE DIGESTIVE TRACT|RADIOGRAPHY OF GASTROINTESTINAL TRACT (PROCEDURE)
C0203102|T060|31911002|SNOMEDCT_US|X-RAY OF KIDNEY, URETER & BLADDER|RADIOGRAPHY OF KIDNEY-URETER-BLADDER (PROCEDURE)
C0203102|T060|31911002|SNOMEDCT_US|KUB X-RAY|RADIOGRAPHY OF KIDNEY-URETER-BLADDER (PROCEDURE)
C0203102|T060|31911002|SNOMEDCT_US|RADIOGRAPHY OF KIDNEY-URETER-BLADDER|RADIOGRAPHY OF KIDNEY-URETER-BLADDER (PROCEDURE)
C0203102|T060|31911002|SNOMEDCT_US|KIDNEYS, URETER, BLADDER X-RAY|RADIOGRAPHY OF KIDNEY-URETER-BLADDER (PROCEDURE)
C0203102|T060|31911002|SNOMEDCT_US|RADIOGRAPHY OF KIDNEY-URETER-BLADDER |RADIOGRAPHY OF KIDNEY-URETER-BLADDER (PROCEDURE)
C0203102|T060|31911002|SNOMEDCT_US|X-RAY OF THE KIDNEY/URETER/BLADDER|RADIOGRAPHY OF KIDNEY-URETER-BLADDER (PROCEDURE)
C0203102|T060|31911002|SNOMEDCT_US|X-RAY;KIDNEY/URETER/BLADDER|RADIOGRAPHY OF KIDNEY-URETER-BLADDER (PROCEDURE)
C2711860|T060|441802002|SNOMEDCT_US|IMAGING OF LIVER|IMAGING OF LIVER (PROCEDURE)
C0203765|T060|37537004|SNOMEDCT_US|LIVER AND SPLEEN IMAGING|LIVER AND SPLEEN IMAGING (PROCEDURE)
C2711446|T060|442684004|SNOMEDCT_US|IMAGING OF LIVER ABNORMAL|IMAGING OF LIVER ABNORMAL (FINDING)
C0203765|T060|37537004|SNOMEDCT_US|LIVER AND SPLEEN IMAGING|LIVER AND SPLEEN IMAGING (PROCEDURE)
C0203765|T060|37537004|SNOMEDCT_US|IMAGING OF LIVER AND SPLEEN|LIVER AND SPLEEN IMAGING (PROCEDURE)
C0203765|T060|37537004|SNOMEDCT_US|LIVER AND SPLEEN IMAGING |LIVER AND SPLEEN IMAGING (PROCEDURE)
C0203758|T060|386552000|SNOMEDCT_US|LIVER SCANNING|RADIOISOTOPE STUDY OF LIVER
C0203761|T060|54780008|SNOMEDCT_US|LIVER IMAGING; WITH VASCULAR FLOW|LIVER IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203761|T060|54780008|SNOMEDCT_US|LIVER IMAGING W/VASCULAR FLOW|LIVER IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203761|T060|54780008|SNOMEDCT_US|IMAGING OF LIVER BLOOD FLOW|LIVER IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203761|T060|54780008|SNOMEDCT_US|LIVER IMAGING WITH VASCULAR FLOW|LIVER IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203761|T060|54780008|SNOMEDCT_US|LIVER IMAGING WITH VASCULAR FLOW |LIVER IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203761|T060|54780008|SNOMEDCT_US|LIVER IMAGING WITH FLOW|LIVER IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203759|T060|169147005|SNOMEDCT_US|LIVER IMAGING; STATIC ONLY|ISOTOPE STATIC SCAN LIVER (PROCEDURE)
C0203759|T060|169147005|SNOMEDCT_US|ISOTOPE STATIC SCAN LIVER|ISOTOPE STATIC SCAN LIVER (PROCEDURE)
C0203759|T060|169147005|SNOMEDCT_US|LIVER IMAGING STATIC ONLY|ISOTOPE STATIC SCAN LIVER (PROCEDURE)
C0203767|T060|81391006|SNOMEDCT_US|LIVER AND SPLEEN IMAGING; WITH VASCULAR FLOW|LIVER AND SPLEEN IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203767|T060|81391006|SNOMEDCT_US|LIVER & SPLEEN IMAGING W/VASCULAR FLOW|LIVER AND SPLEEN IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203767|T060|81391006|SNOMEDCT_US|LIVER AND SPLEEN IMAGING WITH VASCULAR FLOW|LIVER AND SPLEEN IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203767|T060|81391006|SNOMEDCT_US|LIVER AND SPLEEN IMAGING WITH VASCULAR FLOW |LIVER AND SPLEEN IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203767|T060|81391006|SNOMEDCT_US|LIVER & SPLEEN IMAGE/FLOW|LIVER AND SPLEEN IMAGING WITH VASCULAR FLOW (PROCEDURE)
C0203766|T060|13307003|SNOMEDCT_US|LIVER AND SPLEEN IMAGING; STATIC ONLY|RETIRED PROCEDURE [13307003]
C0203766|T060|13307003|SNOMEDCT_US|LIVER & SPLEEN IMAGING STATIC ONLY|RETIRED PROCEDURE [13307003]
C0203766|T060|13307003|SNOMEDCT_US|LIVER AND SPLEEN IMAGING|RETIRED PROCEDURE [13307003]
C1715022|T060||SNOMEDCT_US|LIVER+BDS+GB RI W CCK+RNC IV
C1715022|T060||SNOMEDCT_US|LIVER AND BILIARY DUCTS AND GALLBLADDER SCAN W CHOLECYSTOKININ AND W RADIONUCLIDE IV
C1715022|T060||SNOMEDCT_US|VIEWS^W CHOLECYSTOKININ & W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER+BILIARY DUCTS+GALLBLADDER:DOCUMENT:RADNUC
C1715022|T060||SNOMEDCT_US|VIEWS^W CHOLECYSTOKININ & W RADIONUCLIDE IV:FIND:PT:LIVER+BILIARY DUCTS+GALLBLADDER:DOC:RADNUC
C1715394|T060||SNOMEDCT_US|BD+PDS MRI WO CONTR
C1715394|T060||SNOMEDCT_US|BILIARY DUCTS AND PANCREATIC DUCT MRI WO CONTRAST
C1715394|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:MRI
C1715394|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:MRI
C1525616|T060||SNOMEDCT_US|BD+PDS MRI
C1525616|T060||SNOMEDCT_US|BILIARY DUCTS AND PANCREATIC DUCT MRI
C1525616|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:MRI
C1525616|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:MRI
C0881812|T060||SNOMEDCT_US|BDS+GB FLR IN SURG W CONTR BD
C0881812|T060||SNOMEDCT_US|BILIARY DUCTS AND GALLBLADDER FLUOROSCOPY DURING SURGERY W CONTRAST BILIARY DUCT
C0881812|T060||SNOMEDCT_US|VIEWS^DURING SURGERY W CONTRAST BILIARY DUCT:FINDING:POINT IN TIME:BILIARY DUCTS+GALLBLADDER:DOCUMENT:XR.FLUOR
C0881812|T060||SNOMEDCT_US|VIEWS^DURING SURGERY W CONTRAST BILIARY DUCT:FIND:PT:BILIARY DUCTS+GALLBLADDER:DOC:XR.FLUOR
C0881811|T060||SNOMEDCT_US|BDS+GB XR W CONTR IV
C0881811|T060||SNOMEDCT_US|BILIARY DUCTS AND GALLBLADDER X-RAY W CONTRAST IV
C0881811|T060||SNOMEDCT_US|VIEWS^W CONTRAST IV:FIND:PT:BILIARY DUCTS+GALLBLADDER:DOC:XR
C0881811|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:BILIARY DUCTS+GALLBLADDER:DOCUMENT:XR
C1114931|T060||SNOMEDCT_US|BDS+GB FLR W CONTR VIA T-TB
C1114931|T060||SNOMEDCT_US|BILIARY DUCTS AND GALLBLADDER FLUOROSCOPY W CONTRAST VIA T-TUBE
C1114931|T060||SNOMEDCT_US|VIEWS^W CONTRAST VIA T-TUBE:FIND:PT:BILIARY DUCTS+GALLBLADDER:DOC:XR.FLUOR
C1114931|T060||SNOMEDCT_US|VIEWS^W CONTRAST VIA T-TUBE:FINDING:POINT IN TIME:BILIARY DUCTS+GALLBLADDER:DOCUMENT:XR.FLUOR
C0882518|T060||SNOMEDCT_US|BDS+GB RI FOR BIL PAT+EF W SINC+RNC IV
C0882518|T060||SNOMEDCT_US|BILIARY DUCTS AND GALLBLADDER SCAN FOR PATENCY OF BILIARY STRUCTURES AND EJECTION FRACTION W SINCALIDE AND W RADIONUCLIDE IV
C0882518|T060||SNOMEDCT_US|VIEWS FOR PATENCY OF BILIARY STRUCTURES & EJECTION FRACTION^W SINCALIDE & W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:BILIARY DUCTS+GALLBLADDER:DOCUMENT:RADNUC
C0882518|T060||SNOMEDCT_US|VIEWS FOR PATENCY OF BILIARY STRUCTURES & EJECTION FRACTION^W SINCALIDE & W RADIONUCLIDE IV:FIND:PT:BILIARY DUCTS+GALLBLADDER:DOC:RADNUC
C1715395|T060||SNOMEDCT_US|BD+PDS MRI W CONTR IV
C1715395|T060||SNOMEDCT_US|BILIARY DUCTS AND PANCREATIC DUCT MRI W CONTRAST IV
C1715395|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:MRI
C1715395|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:MRI
C1525615|T060||SNOMEDCT_US|BILIARY DUCTS MRI
C1525615|T060||SNOMEDCT_US|BDS MRI
C1525615|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:BILIARY DUCTS:DOCUMENT:MRI
C1525615|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:BILIARY DUCTS:DOC:MRI
C1525276|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:MRI
C1525276|T060||SNOMEDCT_US|BILIARY DUCTS AND PANCREATIC DUCT MRI WO AND W CONTRAST IV
C1525276|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:MRI
C1525276|T060||SNOMEDCT_US|BD+PDS MRI WO+W CONTR IV
C1715115|T060||SNOMEDCT_US|LIVER+BDS+GB RI FOR PAT W TC99MIV
C1715115|T060||SNOMEDCT_US|LIVER AND BILIARY DUCTS AND GALLBLADDER SCAN FOR PATENCY W TC-99M IV
C1715115|T060||SNOMEDCT_US|VIEWS FOR PATENCY^W TC-99M INTRAVENOUS:FINDING:POINT IN TIME:LIVER+BILIARY DUCTS+GALLBLADDER:DOCUMENT:RADNUC
C1715115|T060||SNOMEDCT_US|VIEWS FOR PATENCY^W TC-99M IV:FIND:PT:LIVER+BILIARY DUCTS+GALLBLADDER:DOC:RADNUC
C4070470|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:ABDOMEN>BILIARY DUCTS:DOC:CT
C4070470|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN>BILIARY DUCTS:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C4070470|T060||SNOMEDCT_US|BILIARY DUCTS CT WO AND W CONTRAST IV
C4070470|T060||SNOMEDCT_US|BD CT WO+W CONTR IV
C0008307|T060|28367004|SNOMEDCT_US|CHOLANGIOGRAPHIES|CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|CHOLANGIOGRAPHY|CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|CHOLANGIOGRAM|CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|CHOLANGIOGR|CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|BILIARY CONTRAST RADIOGRAPHY|CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|BILIARY CONTRAST RADIOGRAPHY NOS|CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|BILIARY CONTRAST RADIOG|CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|BILIARY CONTRAST RADIOGRAPHY NOS |CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|CHOLANGIOGRAM |CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|CONTRAST RADIOGRAPHY OF BILE DUCTS|CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|BILIARY CONTRAST RADIOGRAPHY |CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|CHOLANGIOGRAM, NOS|CHOLANGIOGRAM (PROCEDURE)
C0008307|T060|28367004|SNOMEDCT_US|CONTRAST RADIOGRAPHY OF BILE DUCTS, NOS|CHOLANGIOGRAM (PROCEDURE)
C0008327|T060|241175004|SNOMEDCT_US|CHOLECYSTOGRAPHIES|CHOLECYSTOGRAM (PROCEDURE)
C0008327|T060|241175004|SNOMEDCT_US|CHOLECYSTOGRAPHY|CHOLECYSTOGRAM (PROCEDURE)
C0008327|T060|241175004|SNOMEDCT_US|CHOLECYSTOGR|CHOLECYSTOGRAM (PROCEDURE)
C0008327|T060|241175004|SNOMEDCT_US|CHOLECYSTOGRAM|CHOLECYSTOGRAM (PROCEDURE)
C0008327|T060|241175004|SNOMEDCT_US|CG - CHOLECYSTOGRAM|CHOLECYSTOGRAM (PROCEDURE)
C0008327|T060|241175004|SNOMEDCT_US|CHOLECYSTOGRAM |CHOLECYSTOGRAM (PROCEDURE)
C0203082|T060|81618005|SNOMEDCT_US|INTRAVENOUS CHOLANGIOGRAPHY|INTRAVENOUS CHOLANGIOGRAM (PROCEDURE)
C0203082|T060|81618005|SNOMEDCT_US|INTRAVENOUS CHOLANGIOGRAPHY |INTRAVENOUS CHOLANGIOGRAM (PROCEDURE)
C0203082|T060|81618005|SNOMEDCT_US|X-RAY IV. CHOLANGIOGRAPHY (IVC)|INTRAVENOUS CHOLANGIOGRAM (PROCEDURE)
C0203082|T060|81618005|SNOMEDCT_US|INTRAVEN CHOLANGIOGRAM|INTRAVENOUS CHOLANGIOGRAM (PROCEDURE)
C0203082|T060|81618005|SNOMEDCT_US|INTRAVENOUS CHOLANGIOGRAM|INTRAVENOUS CHOLANGIOGRAM (PROCEDURE)
C0203082|T060|81618005|SNOMEDCT_US|INTRAVENOUS CHOLANGIOGRAM |INTRAVENOUS CHOLANGIOGRAM (PROCEDURE)
C0203082|T060|81618005|SNOMEDCT_US|IVC - INTRAVENOUS CHOLANGIOGRAM|INTRAVENOUS CHOLANGIOGRAM (PROCEDURE)
C0203082|T060|81618005|SNOMEDCT_US|INFUSION CHOLANGIOGRAM|INTRAVENOUS CHOLANGIOGRAM (PROCEDURE)
C0029538|T060||SNOMEDCT_US|CHOLANGIOGRAM NEC
C0029538|T060||SNOMEDCT_US|OTHER CHOLANGIOGRAM
C0177740|T060||SNOMEDCT_US|BILIARY TRACT X-RAY NEC
C0177740|T060||SNOMEDCT_US|OTHER BILIARY TRACT X-RAY
C0881931|T060||SNOMEDCT_US|GALLBLADDER US
C0881931|T060||SNOMEDCT_US|GB US
C0881931|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:GALLBLADDER:DOC:US
C0881931|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:GALLBLADDER:DOCUMENT:ULTRASOUND
C1543917|T060||SNOMEDCT_US|GB RI EF W TC99MDISIDA IV
C1543917|T060||SNOMEDCT_US|GALLBLADDER SCAN EJECTION FRACTION W TC-99M DISIDA IV
C1543917|T060||SNOMEDCT_US|VIEWS EJECTION FRACTION^W TC-99M DISIDA IV:FIND:PT:GALLBLADDER:DOC:RADNUC
C1543917|T060||SNOMEDCT_US|VIEWS EJECTION FRACTION^W TC-99M DISIDA INTRAVENOUS:FINDING:POINT IN TIME:GALLBLADDER:DOCUMENT:RADNUC
C1526261|T060||SNOMEDCT_US|GALLBLADDER US LIMITED
C1526261|T060||SNOMEDCT_US|GB US LTD
C1526261|T060||SNOMEDCT_US|MULTISECTION LIMITED:FIND:PT:GALLBLADDER:DOC:US
C1526261|T060||SNOMEDCT_US|MULTISECTION LIMITED:FINDING:POINT IN TIME:GALLBLADDER:DOCUMENT:ULTRASOUND
C1526263|T060||SNOMEDCT_US|GB US W CCK
C1526263|T060||SNOMEDCT_US|GALLBLADDER US W CHOLECYSTOKININ
C1526263|T060||SNOMEDCT_US|MULTISECTION^W CHOLECYSTOKININ:FIND:PT:GALLBLADDER:DOC:US
C1526263|T060||SNOMEDCT_US|MULTISECTION^W CHOLECYSTOKININ:FINDING:POINT IN TIME:GALLBLADDER:DOCUMENT:ULTRASOUND
C1542969|T060||SNOMEDCT_US|GB RI W TC99MDISIDA IV
C1542969|T060||SNOMEDCT_US|GALLBLADDER SCAN W TC-99M DISIDA IV
C1542969|T060||SNOMEDCT_US|VIEWS^W TC-99M DISIDA INTRAVENOUS:FINDING:POINT IN TIME:GALLBLADDER:DOCUMENT:RADNUC
C1542969|T060||SNOMEDCT_US|VIEWS^W TC-99M DISIDA IV:FIND:PT:GALLBLADDER:DOC:RADNUC
C2608012|T060||SNOMEDCT_US|VIEWS^W CONTRAST TRANSHEPATIC:FINDING:POINT IN TIME:PORTAL VEIN:NARRATIVE:XR.FLUOR.ANGIO
C2608012|T060||SNOMEDCT_US|PORTAL VEIN FLUOROSCOPIC ANGIOGRAM W CONTRAST TRANSHEPATIC
C2608012|T060||SNOMEDCT_US|PORTAL V XRA W CONTR TH
C2608012|T060||SNOMEDCT_US|VIEWS^W CONTRAST TRANSHEPATIC:FINDING:POINT IN TIME:PORTAL VEIN:DOCUMENT:XR.FLUOR.ANGIO
C2608012|T060||SNOMEDCT_US|VIEWS^W CONTRAST TRANSHEPATIC:FIND:PT:PORTAL VEIN:DOC:XR.FLUOR.ANGIO
C0882151|T060||SNOMEDCT_US|SPLENIC V+PORTAL V XRA W CONTR IA
C0882151|T060||SNOMEDCT_US|SPLENIC VEIN AND PORTAL VEIN FLUOROSCOPIC ANGIOGRAM W CONTRAST IA
C0882151|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRA-ARTERIAL:FINDING:POINT IN TIME:SPLENIC VEIN+PORTAL VEIN:DOCUMENT:XR.FLUOR.ANGIO
C0882151|T060||SNOMEDCT_US|VIEWS^W CONTRAST IA:FIND:PT:SPLENIC VEIN+PORTAL VEIN:DOC:XR.FLUOR.ANGIO
C1114641|T060||SNOMEDCT_US|VIEWS^W CONTRAST TRANSHEPATIC & W HEMODYNAMICS:FINDING:POINT IN TIME:PORTAL VEIN:NARRATIVE:XR.FLUOR.ANGIO
C1114641|T060||SNOMEDCT_US|PORTAL V XRA W CONTR TH+HEMODYN
C1114641|T060||SNOMEDCT_US|PORTAL VEIN FLUOROSCOPIC ANGIOGRAM W CONTRAST TRANSHEPATIC AND W HEMODYNAMICS
C1114641|T060||SNOMEDCT_US|VIEWS^W CONTRAST TRANSHEPATIC & W HEMODYNAMICS:FINDING:POINT IN TIME:PORTAL VEIN:DOCUMENT:XR.FLUOR.ANGIO
C1114641|T060||SNOMEDCT_US|VIEWS^W CONTRAST TRANSHEPATIC & W HEMODYNAMICS:FIND:PT:PORTAL VEIN:DOC:XR.FLUOR.ANGIO
C3263063|T060||SNOMEDCT_US|PORTAL V XRA W CONTR IV
C3263063|T060||SNOMEDCT_US|PORTAL VEIN FLUOROSCOPIC ANGIOGRAM W CONTRAST IV
C3263063|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:PORTAL VEIN:DOCUMENT:XR.FLUOR.ANGIO
C1524919|T060||SNOMEDCT_US|PORTAL VEIN MRI ANGIOGRAM WO CONTRAST
C1524919|T060||SNOMEDCT_US|PORTAL V MRI.ANGIO WO CONTR
C1524919|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FINDING:POINT IN TIME:PORTAL VEIN:DOCUMENT:MRI.ANGIO
C1524919|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FIND:PT:PORTAL VEIN:DOC:MRI.ANGIO
C1524189|T060||SNOMEDCT_US|PORTAL V MRI.ANGIO
C1524189|T060||SNOMEDCT_US|PORTAL VEIN MRI ANGIOGRAM
C1524189|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:PORTAL VEIN:DOC:MRI.ANGIO
C1524189|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:PORTAL VEIN:DOCUMENT:MRI.ANGIO
C0202977|T060|55612007|SNOMEDCT_US|VENOGRAPHY OF LIVER |HEPATIC VENOGRAPHY (PROCEDURE)
C0202977|T060|55612007|SNOMEDCT_US|VENOGRAPHY OF LIVER|HEPATIC VENOGRAPHY (PROCEDURE)
C0202977|T060|55612007|SNOMEDCT_US|HEPATIC VENOGRAPHY|HEPATIC VENOGRAPHY (PROCEDURE)
C0202977|T060|55612007|SNOMEDCT_US|HEPATIC VENOGRAM|HEPATIC VENOGRAPHY (PROCEDURE)
C0202977|T060|55612007|SNOMEDCT_US|HEPATIC VENOGRAPHY |HEPATIC VENOGRAPHY (PROCEDURE)
C0202977|T060|55612007|SNOMEDCT_US|HEPATIC PHLEBOGRAPHY|HEPATIC VENOGRAPHY (PROCEDURE)
C0412627|T060|241554003|SNOMEDCT_US|CT ARTERIOPORTOGRAPHY |COMPUTED TOMOGRAPHY ARTERIOPORTOGRAPHY
C0412627|T060|241554003|SNOMEDCT_US|COMPUTED TOMOGRAPHY ARTERIOPORTOGRAPHY |COMPUTED TOMOGRAPHY ARTERIOPORTOGRAPHY
C0412627|T060|241554003|SNOMEDCT_US|COMPUTED TOMOGRAPHY ARTERIOPORTOGRAPHY|COMPUTED TOMOGRAPHY ARTERIOPORTOGRAPHY
C0412627|T060|241554003|SNOMEDCT_US|CT ARTERIOPORTOGRAPHY|COMPUTED TOMOGRAPHY ARTERIOPORTOGRAPHY
C1525185|T060||SNOMEDCT_US|HEPATIC ARTERY CT ANGIOGRAM W CONTRAST IA
C1525185|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IA:FIND:PT:ABDOMEN>HEPATIC ARTERY:DOC:CT.ANGIO
C1525185|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRA-ARTERIAL:FINDING:POINT IN TIME:ABDOMEN>HEPATIC ARTERY:DOCUMENT:COMPUTERIZED TOMOGRAPHY.ANGIO
C1525185|T060||SNOMEDCT_US|ABD>HEP A CT.ANGIO W CONTR IA
C4039140|T060|708733006|SNOMEDCT_US|LIVER ANGIOGRAPHY|ANGIOGRAPHY OF LIVER (PROCEDURE)
C4039140|T060|708733006|SNOMEDCT_US|ANGIOGRAPHY OF LIVER |ANGIOGRAPHY OF LIVER (PROCEDURE)
C4039140|T060|708733006|SNOMEDCT_US|ANGIOGRAPHY OF LIVER|ANGIOGRAPHY OF LIVER (PROCEDURE)
C1114644|T060||SNOMEDCT_US|IVC XRA W CONTR IV
C1114644|T060||SNOMEDCT_US|INFERIOR VENA CAVA FLUOROSCOPIC ANGIOGRAM W CONTRAST IV
C1114644|T060||SNOMEDCT_US|VIEWS^W CONTRAST IV:FIND:PT:VENA CAVA.INFERIOR:DOC:XR.FLUOR.ANGIO
C1114644|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:VENA CAVA.INFERIOR:DOCUMENT:XR.FLUOR.ANGIO
C1114661|T060||SNOMEDCT_US|ABD VV+IVC MRI.ANGIO
C1114661|T060||SNOMEDCT_US|ABDOMINAL VEINS AND IVC MRI ANGIOGRAM
C1114661|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMINAL VEINS+VENA CAVA.INFERIOR:DOC:MRI.ANGIO
C1114661|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMINAL VEINS+VENA CAVA.INFERIOR:DOCUMENT:MRI.ANGIO
C1525107|T060||SNOMEDCT_US|ABD VV MRI.ANGIO
C1525107|T060||SNOMEDCT_US|ABDOMINAL VEINS MRI ANGIOGRAM
C1525107|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMINAL VEINS:DOC:MRI.ANGIO
C1525107|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMINAL VEINS:DOCUMENT:MRI.ANGIO
C1524195|T060||SNOMEDCT_US|IVC MRI
C1524195|T060||SNOMEDCT_US|INFERIOR VENA CAVA MRI
C1524195|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:VENA CAVA.INFERIOR:DOCUMENT:MRI
C1524195|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:VENA CAVA.INFERIOR:DOC:MRI
C0882181|T060||SNOMEDCT_US|VC XRA W CONTR IV
C0882181|T060||SNOMEDCT_US|VENA CAVA FLUOROSCOPIC ANGIOGRAM W CONTRAST IV
C0882181|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:VENA CAVA:DOCUMENT:XR.FLUOR.ANGIO
C0882181|T060||SNOMEDCT_US|VIEWS^W CONTRAST IV:FIND:PT:VENA CAVA:DOC:XR.FLUOR.ANGIO
C1543874|T060||SNOMEDCT_US|LIVER SCAN STATIC
C1543874|T060||SNOMEDCT_US|LIVER RI STATIC W RNC IV
C1543874|T060||SNOMEDCT_US|VIEWS STATIC^W RADIONUCLIDE IV:FIND:PT:LIVER:DOC:RADNUC
C1543874|T060||SNOMEDCT_US|VIEWS STATIC^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:RADNUC
C1524194|T060||SNOMEDCT_US|IVC MRI.ANGIO
C1524194|T060||SNOMEDCT_US|INFERIOR VENA CAVA MRI ANGIOGRAM
C1524194|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:VENA CAVA.INFERIOR:DOCUMENT:MRI.ANGIO
C1524194|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:VENA CAVA.INFERIOR:DOC:MRI.ANGIO
C1543214|T060||SNOMEDCT_US|HEP VS XRA W CONTR IV
C1543214|T060||SNOMEDCT_US|HEPATIC VEINS FLUOROSCOPIC ANGIOGRAM W CONTRAST IV
C1543214|T060||SNOMEDCT_US|VIEWS^W CONTRAST IV:FIND:PT:HEPATIC VEINS:DOC:XR.FLUOR.ANGIO
C1543214|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:HEPATIC VEINS:DOCUMENT:XR.FLUOR.ANGIO
C1525728|T060||SNOMEDCT_US|CELIAC A+GASTRIC A-L+SMA XRA W CONTR IA
C1525728|T060||SNOMEDCT_US|CELIAC ARTERY AND GASTRIC ARTERY - LEFT AND SUPERIOR MESENTERIC ARTERY FLUOROSCOPIC ANGIOGRAM W CONTRAST IA
C1525728|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRA-ARTERIAL:FINDING:POINT IN TIME:CELIAC ARTERY+GASTRIC ARTERY.LEFT+SUPERIOR MESENTERIC ARTERY:DOCUMENT:XR.FLUOR.ANGIO
C1525728|T060||SNOMEDCT_US|VIEWS^W CONTRAST IA:FIND:PT:CELIAC ARTERY+GASTRIC ARTERY.LEFT+SUPERIOR MESENTERIC ARTERY:DOC:XR.FLUOR.ANGIO
C1525229|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:ABDOMINAL VESSELS:DOC:MRI.ANGIO
C1525229|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:MRI.ANGIO
C1525229|T060||SNOMEDCT_US|ABD VES MRI.ANGIO WO+W CONTR IV
C1525229|T060||SNOMEDCT_US|ABDOMINAL VESSELS MRI ANGIOGRAM WO AND W CONTRAST IV
C1525203|T060||SNOMEDCT_US|ABD VES CT.ANGIO W CONTR IV
C1525203|T060||SNOMEDCT_US|ABDOMINAL VESSELS CT ANGIOGRAM W CONTRAST IV
C1525203|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:ABDOMEN>VESSELS:DOC:CT.ANGIO
C1525203|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN>VESSELS:DOCUMENT:COMPUTERIZED TOMOGRAPHY.ANGIO
C3262889|T060||SNOMEDCT_US|ABD VES XRA W CONTR IV
C3262889|T060||SNOMEDCT_US|ABDOMINAL VESSELS FLUOROSCOPIC ANGIOGRAM W CONTRAST IV
C3262889|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:XR.FLUOR.ANGIO
C3262889|T060||SNOMEDCT_US|VIEWS^W CONTRAST IV:FIND:PT:ABDOMINAL VESSELS:DOC:XR.FLUOR.ANGIO
C1525117|T060||SNOMEDCT_US|ABDOMINAL VESSELS MRI ANGIOGRAM
C1525117|T060||SNOMEDCT_US|ABD VES MRI.ANGIO
C1525117|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMINAL VESSELS:DOC:MRI.ANGIO
C1525117|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:MRI.A
C0881776|T060||SNOMEDCT_US|ABDOMINAL VESSELS US.DOPPLER
C0881776|T060||SNOMEDCT_US|ABD VES DOP
C0881776|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:ULTRASOUND.DOPPLER
C0881776|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMINAL VESSELS:DOC:US.DOPPLER
C0881775|T060||SNOMEDCT_US|ABD VES MRI.ANGIO W CONTR IV
C0881775|T060||SNOMEDCT_US|ABDOMINAL VESSELS MRI ANGIOGRAM W CONTRAST IV
C0881775|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:MRI.ANGIO
C0881775|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:ABDOMINAL VESSELS:DOC:MRI.ANGIO
C1525251|T060||SNOMEDCT_US|ABD VES MRI.ANGIO WO CONTR
C1525251|T060||SNOMEDCT_US|ABDOMINAL VESSELS MRI ANGIOGRAM WO CONTRAST
C1525251|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:MRI.ANGIO
C1525251|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FIND:PT:ABDOMINAL VESSELS:DOC:MRI.ANGIO
C0882186|T060||SNOMEDCT_US|ABD AA XRA W CONTR IA
C0882186|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRA-ARTERIAL:FINDING:POINT IN TIME:ABDOMINAL ARTERIES:DOCUMENT:XR.FLUOR.ANGIO
C0882186|T060||SNOMEDCT_US|VIEWS^W CONTRAST IA:FIND:PT:ABDOMINAL ARTERIES:DOC:XR.FLUOR.ANGIO
C0882186|T060||SNOMEDCT_US|ABDOMINAL ARTERIES FLUOROSCOPIC ANGIOGRAM W CONTRAST IA
C1114660|T060||SNOMEDCT_US|AORTA+ABD AA MRI.ANGIO
C1114660|T060||SNOMEDCT_US|ABDOMINAL AORTA AND ARTERIES MRI ANGIOGRAM
C1114660|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:AORTA+ABDOMINAL ARTERIES:DOC:MRI.ANGIO
C1114660|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:AORTA+ABDOMINAL ARTERIES:DOCUMENT:MRI.ANGIO
C1114662|T060||SNOMEDCT_US|CELIAC VES+SM VES MRI.ANGIO
C1114662|T060||SNOMEDCT_US|CELIAC VESSELS AND SUPERIOR MESENTERIC VESSELS MRI ANGIOGRAM
C1114662|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:CELIAC VESSELS+SUPERIOR MESENTERIC VESSELS:DOCUMENT:MRI.ANGIO
C1114662|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:CELIAC VESSELS+SUPERIOR MESENTERIC VESSELS:DOC:MRI.ANGIO
C1525229|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:ABDOMINAL VESSELS:DOC:MRI.ANGIO
C1525229|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:MRI.ANGIO
C1525229|T060||SNOMEDCT_US|ABD VES MRI.ANGIO WO+W CONTR IV
C1525229|T060||SNOMEDCT_US|ABDOMINAL VESSELS MRI ANGIOGRAM WO AND W CONTRAST IV
C1525203|T060||SNOMEDCT_US|ABD VES CT.ANGIO W CONTR IV
C1525203|T060||SNOMEDCT_US|ABDOMINAL VESSELS CT ANGIOGRAM W CONTRAST IV
C1525203|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:ABDOMEN>VESSELS:DOC:CT.ANGIO
C1525203|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN>VESSELS:DOCUMENT:COMPUTERIZED TOMOGRAPHY.ANGIO
C3262889|T060||SNOMEDCT_US|ABD VES XRA W CONTR IV
C3262889|T060||SNOMEDCT_US|ABDOMINAL VESSELS FLUOROSCOPIC ANGIOGRAM W CONTRAST IV
C3262889|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:XR.FLUOR.ANGIO
C3262889|T060||SNOMEDCT_US|VIEWS^W CONTRAST IV:FIND:PT:ABDOMINAL VESSELS:DOC:XR.FLUOR.ANGIO
C1525117|T060||SNOMEDCT_US|ABDOMINAL VESSELS MRI ANGIOGRAM
C1525117|T060||SNOMEDCT_US|ABD VES MRI.ANGIO
C1525117|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMINAL VESSELS:DOC:MRI.ANGIO
C1525117|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:MRI.A
C0881776|T060||SNOMEDCT_US|ABDOMINAL VESSELS US.DOPPLER
C0881776|T060||SNOMEDCT_US|ABD VES DOP
C0881776|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:ULTRASOUND.DOPPLER
C0881776|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:ABDOMINAL VESSELS:DOC:US.DOPPLER
C0881775|T060||SNOMEDCT_US|ABD VES MRI.ANGIO W CONTR IV
C0881775|T060||SNOMEDCT_US|ABDOMINAL VESSELS MRI ANGIOGRAM W CONTRAST IV
C0881775|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:MRI.ANGIO
C0881775|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:ABDOMINAL VESSELS:DOC:MRI.ANGIO
C1525251|T060||SNOMEDCT_US|ABD VES MRI.ANGIO WO CONTR
C1525251|T060||SNOMEDCT_US|ABDOMINAL VESSELS MRI ANGIOGRAM WO CONTRAST
C1525251|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FINDING:POINT IN TIME:ABDOMINAL VESSELS:DOCUMENT:MRI.ANGIO
C1525251|T060||SNOMEDCT_US|MULTISECTION^WO CONTRAST:FIND:PT:ABDOMINAL VESSELS:DOC:MRI.ANGIO
C0882186|T060||SNOMEDCT_US|ABD AA XRA W CONTR IA
C0882186|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRA-ARTERIAL:FINDING:POINT IN TIME:ABDOMINAL ARTERIES:DOCUMENT:XR.FLUOR.ANGIO
C0882186|T060||SNOMEDCT_US|VIEWS^W CONTRAST IA:FIND:PT:ABDOMINAL ARTERIES:DOC:XR.FLUOR.ANGIO
C0882186|T060||SNOMEDCT_US|ABDOMINAL ARTERIES FLUOROSCOPIC ANGIOGRAM W CONTRAST IA
C1114660|T060||SNOMEDCT_US|AORTA+ABD AA MRI.ANGIO
C1114660|T060||SNOMEDCT_US|ABDOMINAL AORTA AND ARTERIES MRI ANGIOGRAM
C1114660|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:AORTA+ABDOMINAL ARTERIES:DOC:MRI.ANGIO
C1114660|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:AORTA+ABDOMINAL ARTERIES:DOCUMENT:MRI.ANGIO
C1114662|T060||SNOMEDCT_US|CELIAC VES+SM VES MRI.ANGIO
C1114662|T060||SNOMEDCT_US|CELIAC VESSELS AND SUPERIOR MESENTERIC VESSELS MRI ANGIOGRAM
C1114662|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:CELIAC VESSELS+SUPERIOR MESENTERIC VESSELS:DOCUMENT:MRI.ANGIO
C1114662|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:CELIAC VESSELS+SUPERIOR MESENTERIC VESSELS:DOC:MRI.ANGIO
C2713072|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:VESSELS.ABDOMEN:NAR:US.DOPPLER
C2713072|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:VESSELS.ABDOMEN:NARRATIVE:ULTRASOUND.DOPPLER
C1525720|T060||SNOMEDCT_US|CELIAC A+SMA+IMA XRA W CONTR IA
C1525720|T060||SNOMEDCT_US|CELIAC ARTERY AND SUPERIOR MESENTERIC ARTERY AND INFERIOR MESENTERIC ARTERY FLUOROSCOPIC ANGIOGRAM W CONTRAST IA
C1525720|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRA-ARTERIAL:FINDING:POINT IN TIME:CELIAC ARTERY+SUPERIOR MESENTERIC ARTERY+INFERIOR MESENTERIC ARTERY:DOCUMENT:XR.FLUOR.ANGIO
C1525720|T060||SNOMEDCT_US|VIEWS^W CONTRAST IA:FIND:PT:CELIAC ARTERY+SUPERIOR MESENTERIC ARTERY+INFERIOR MESENTERIC ARTERY:DOC:XR.FLUOR.ANGIO
C0881854|T060||SNOMEDCT_US|CELIAC A XRA W CONTR IA
C0881854|T060||SNOMEDCT_US|CELIAC ARTERY FLUOROSCOPIC ANGIOGRAM W CONTRAST IA
C0881854|T060||SNOMEDCT_US|VIEWS^W CONTRAST IA:FIND:PT:CELIAC ARTERY:DOC:XR.FLUOR.ANGIO
C0881854|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRA-ARTERIAL:FINDING:POINT IN TIME:CELIAC ARTERY:DOCUMENT:XR.FLUOR.ANGIO
C4036483|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:CHEST+ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.THORACIC+AORTA.ABDOMINAL+RO VESSELS.BILATERAL:DOCUMENT:COMPUTERIZED TOMOGRAPHY.ANGIO
C4036483|T060||SNOMEDCT_US|T+A.AO+RO V-BL CT.ANGIO WO+W CONTR IV
C4036483|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:CHEST+ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.THORACIC+AORTA.ABDOMINAL+RO VESSELS.BILATERAL:DOC:CT.ANGIO
C4036483|T060||SNOMEDCT_US|THORACIC AND ABDOMINAL AORTA AND BILATERAL RUNOFF VESSELS CT ANGIOGRAM WO AND W CONTRAST IV
C4036886|T060||SNOMEDCT_US|MULTISECTION FOR ENDOGRAFT:FIND:PT:CHEST+ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.THORACIC+AORTA.ABDOMINAL+VESSELS.BILATERAL:DOC:CT.ANGIO
C4036886|T060||SNOMEDCT_US|THORACIC AND ABDOMINAL AORTA AND BILATERAL VESSELS CT ANGIOGRAM FOR ENDOGRAFT
C4036886|T060||SNOMEDCT_US|T AO+ABD AO+VES-BL CT.ANGIO FOR ENDOGRAF
C4036886|T060||SNOMEDCT_US|MULTISECTION FOR ENDOGRAFT:FINDING:POINT IN TIME:CHEST+ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.THORACIC+AORTA.ABDOMINAL+VESSELS.BILATERAL:DOCUMENT:COMPUTERIZED TOMOGRAPHY.ANGIO
C4036484|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.ABDOMINAL+RO VESSELS.BILATERAL:DOCUMENT:COMPUTERIZED TOMOGRAPHY.ANGIO
C4036484|T060||SNOMEDCT_US|MULTISECTION^WO & W CONTRAST IV:FIND:PT:ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.ABDOMINAL+RO VESSELS.BILATERAL:DOC:CT.ANGIO
C4036484|T060||SNOMEDCT_US|ABDOMINAL AORTA AND BILATERAL RUNOFF VESSELS CT ANGIOGRAM WO AND W CONTRAST IV
C4036484|T060||SNOMEDCT_US|ABD AORTA+ROVES-BL CT.ANGIO WO+WCONTRIV
C4036480|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.ABDOMINAL+RO VESSELS.BILATERAL:DOCUMENT:COMPUTERIZED TOMOGRAPHY.ANGIO
C4036480|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.ABDOMINAL+RO VESSELS.BILATERAL:DOC:CT.ANGIO
C4036480|T060||SNOMEDCT_US|ABDOMINAL AORTA AND BILATERAL RUNOFF VESSELS CT ANGIOGRAM W CONTRAST IV
C4036480|T060||SNOMEDCT_US|ABD AORTA+RO VES-BL CT.ANGIO W CONTR IV
C4036887|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:CHEST+ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.THORACIC+AORTA.ABDOMINAL+VESSELS.BILATERAL:DOC:CT.ANGIO
C4036887|T060||SNOMEDCT_US|DEPRECATED CHEST+ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.THORACIC+AORTA.ABDOMINAL+VESSELS CT ANGIOGRAM W CONTRAST IV
C4036887|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:CHEST+ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.THORACIC+AORTA.ABDOMINAL+VESSELS.BILATERAL:DOCUMENT:COMPUTERIZED TOMOGRAPHY.ANGIO
C4036887|T060||SNOMEDCT_US|DEPRECATED C+A+P+LXB>A.TH+A CT.ANGIO W C
C4036479|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:CHEST+ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.THORACIC+AORTA.ABDOMINAL+RO VESSELS.BILATERAL:DOCUMENT:COMPUTERIZED TOMOGRAPHY.ANGIO
C4036479|T060||SNOMEDCT_US|THORACIC AND ABDOMINAL AORTA AND BILATERAL RUNOFF VESSELS CT ANGIOGRAM W CONTRAST IV
C4036479|T060||SNOMEDCT_US|T+A.AO+RO V-BL CT.ANGIO W CONTR IV
C4036479|T060||SNOMEDCT_US|MULTISECTION^W CONTRAST IV:FIND:PT:CHEST+ABDOMEN+PELVIS+LOWER EXTREMITY.BILATERAL>AORTA.THORACIC+AORTA.ABDOMINAL+RO VESSELS.BILATERAL:DOC:CT.ANGIO
C1524140|T060||SNOMEDCT_US|LYMPH ABD+PELVIC FLR W CONTR IL
C1524140|T060||SNOMEDCT_US|LYMPHATICS ABDOMINAL AND LYMPHATICS PELVIC FLUOROSCOPY W CONTRAST INTRA LYMPHATIC
C1524140|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRA LYMPHATIC:FIND:PT:LYMPHATICS.ABDOMINAL+LYMPHATICS.PELVIC:DOC:XR.FLUOR
C1524140|T060||SNOMEDCT_US|VIEWS^W CONTRAST INTRA LYMPHATIC:FINDING:POINT IN TIME:LYMPHATICS.ABDOMINAL+LYMPHATICS.PELVIC:DOCUMENT:XR.FLUOR
C0202991|T060|91119001|SNOMEDCT_US|ABDOMINAL LYMPHANGIOGRAM|ABDOMINAL LYMPHANGIOGRAM (PROCEDURE)
C0202991|T060|91119001|SNOMEDCT_US|ABDOMINAL LYMPHANGIOGRAM |ABDOMINAL LYMPHANGIOGRAM (PROCEDURE)
C0202991|T060|91119001|SNOMEDCT_US|LYMPHANGIOGRAPHY ABDOMEN|ABDOMINAL LYMPHANGIOGRAM (PROCEDURE)
C0202991|T060|91119001|SNOMEDCT_US|ABDOMINAL LYMPHANGIOGRAM, NOS|ABDOMINAL LYMPHANGIOGRAM (PROCEDURE)
C2584955|T060|438529005|SNOMEDCT_US|MRI GUIDED ABLATION OF LIVER|ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE
C4039879|T060|708697000|SNOMEDCT_US|IMAGING GUIDED PERCUTANEOUS FINE NEEDLE ASPIRATION BIOPSY OF LIVER|PERCUTANEOUS FINE NEEDLE ASPIRATION BIOPSY OF LIVER USING IMAGING GUIDANCE
C2584862|T060|441138007|SNOMEDCT_US|MRI GUIDED FOCUSED ULTRASOUND ABLATION OF LIVER|FOCUSED ULTRASOUND ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE (PROCEDURE)
C2317407|T060|432226009|SNOMEDCT_US|ABLATION OF LESION OF LIVER USING COMPUTED TOMOGRAPHY (CT) GUIDANCE|ABLATION OF LESION OF LIVER USING COMPUTED TOMOGRAPHY (CT) GUIDANCE
C2317407|T060|432226009|SNOMEDCT_US|ABLATION OF LESION OF LIVER USING COMPUTED TOMOGRAPHY GUIDANCE |ABLATION OF LESION OF LIVER USING COMPUTED TOMOGRAPHY (CT) GUIDANCE
C2317407|T060|432226009|SNOMEDCT_US|ABLATION OF LESION OF LIVER USING COMPUTED TOMOGRAPHY GUIDANCE|ABLATION OF LESION OF LIVER USING COMPUTED TOMOGRAPHY (CT) GUIDANCE
C2317407|T060|432226009|SNOMEDCT_US|CT GUIDED ABLATION OF LESION OF LIVER|ABLATION OF LESION OF LIVER USING COMPUTED TOMOGRAPHY (CT) GUIDANCE
C1636186|T060|418158005|SNOMEDCT_US|CT AND DRAINAGE OF LIVER|COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER
C1636186|T060|418158005|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER |COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER
C1636186|T060|418158005|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER|COMPUTED TOMOGRAPHY AND DRAINAGE OF LIVER
C1640379|T060|418458003|SNOMEDCT_US|CT AND ASPIRATION OF LIVER|COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER
C1640379|T060|418458003|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER |COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER
C1640379|T060|418458003|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER|COMPUTED TOMOGRAPHY AND ASPIRATION OF LIVER
C1628488|T060|418749009|SNOMEDCT_US|CT AND BIOPSY OF LIVER|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER
C1628488|T060|418749009|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER |COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER
C1628488|T060|418749009|SNOMEDCT_US|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER|COMPUTED TOMOGRAPHY AND BIOPSY OF LIVER
C1715485|T060||SNOMEDCT_US|LIVER FLR BX NEEDLE GUID W CONTR IV
C1715485|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR NEEDLE BIOPSY OF LIVER-- W CONTRAST IV
C1715485|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.NEEDLE^W CONTRAST IV:FIND:PT:LIVER:DOC:XR.FLUOR
C1715485|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.NEEDLE^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:XR.FLUOR
C3262915|T060||SNOMEDCT_US|CT GUIDANCE FOR BIOPSY OF LIVER-- WO CONTRAST
C3262915|T060||SNOMEDCT_US|LIVER CT BX GUID WO CONTR
C3262915|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY^WO CONTRAST:FIND:PT:ABDOMEN>LIVER:DOC:CT
C3262915|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY^WO CONTRAST:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C3262920|T060||SNOMEDCT_US|CT GUIDANCE FOR NEEDLE BIOPSY OF LIVER
C3262920|T060||SNOMEDCT_US|LIVER CT BX NEEDLE GUID
C3262920|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.NEEDLE:FIND:PT:ABDOMEN>LIVER:DOC:CT
C3262920|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.NEEDLE:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C3263059|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR PERCUTANEOUS NEEDLE BIOPSY OF LIVER
C3263059|T060||SNOMEDCT_US|LIVER FLR PC BX NEEDLE GUID
C3263059|T060||SNOMEDCT_US|GUIDANCE FOR PERCUTANEOUS BIOPSY.NEEDLE:FINDING:POINT IN TIME:LIVER:DOCUMENT:XR.FLUOR
C3263059|T060||SNOMEDCT_US|GUIDANCE FOR PERCUTANEOUS BIOPSY.NEEDLE:FIND:PT:LIVER:DOC:XR.FLUOR
C0882010|T060||SNOMEDCT_US|CT GUIDANCE FOR BIOPSY OF LIVER
C0882010|T060||SNOMEDCT_US|LIVER CT BX GUID
C0882010|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FIND:PT:ABDOMEN>LIVER:DOC:CT
C0882010|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1524318|T060||SNOMEDCT_US|CT GUIDANCE FOR DRAINAGE OF LIVER
C1524318|T060||SNOMEDCT_US|LIVER CT DRAIN GUID
C1524318|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1524318|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE:FIND:PT:ABDOMEN>LIVER:DOC:CT
C1525161|T060||SNOMEDCT_US|US GUIDANCE FOR BIOPSY OF LIVER TRANSPLANT
C1525161|T060||SNOMEDCT_US|LIVER TRANSPLANT US BX GUID
C1525161|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FIND:PT:LIVER TRANSPLANT:DOC:US
C1525161|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FINDING:POINT IN TIME:LIVER TRANSPLANT:DOCUMENT:ULTRASOUND
C1524299|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR BIOPSY OF LIVER
C1524299|T060||SNOMEDCT_US|LIVER FLR BX GUID
C1524299|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FINDING:POINT IN TIME:LIVER:DOCUMENT:XR.FLUOR
C1524299|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FIND:PT:LIVER:DOC:XR.FLUOR
C1633403|T060||SNOMEDCT_US|LIVER FLR TUBE PLAC GUID
C1633403|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR PLACEMENT OF TUBE IN LIVER
C1633403|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF TUBE:FINDING:POINT IN TIME:LIVER:DOCUMENT:XR.FLUOR
C1633403|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF TUBE:FIND:PT:LIVER:DOC:XR.FLUOR
C0882009|T060||SNOMEDCT_US|LIVER CT ASP GUID
C0882009|T060||SNOMEDCT_US|CT GUIDANCE FOR ASPIRATION OF LIVER
C0882009|T060||SNOMEDCT_US|GUIDANCE FOR ASPIRATION:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C0882009|T060||SNOMEDCT_US|GUIDANCE FOR ASPIRATION:FIND:PT:ABDOMEN>LIVER:DOC:CT
C1114431|T060||SNOMEDCT_US|CT GUIDANCE FOR FINE NEEDLE ASPIRATION OF LIVER
C1114431|T060||SNOMEDCT_US|LIVER CT FNA ASP
C1114431|T060||SNOMEDCT_US|GUIDANCE FOR ASPIRATION.FINE NEEDLE:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1114431|T060||SNOMEDCT_US|GUIDANCE FOR ASPIRATION.FINE NEEDLE:FIND:PT:ABDOMEN>LIVER:DOC:CT
C3262948|T060||SNOMEDCT_US|LIVER FLR BX NEEDLE GUID
C3262948|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR NEEDLE BIOPSY OF LIVER
C3262948|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.NEEDLE:FINDING:POINT IN TIME:LIVER:DOCUMENT:XR.FLUOR
C3262948|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.NEEDLE:FIND:PT:LIVER:DOC:XR.FLUOR
C1715480|T060||SNOMEDCT_US|LIVER FLR FNA ASP
C1715480|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR FINE NEEDLE ASPIRATION OF LIVER
C1715480|T060||SNOMEDCT_US|GUIDANCE FOR ASPIRATION.FINE NEEDLE:FIND:PT:LIVER:DOC:XR.FLUOR
C1715480|T060||SNOMEDCT_US|GUIDANCE FOR ASPIRATION.FINE NEEDLE:FINDING:POINT IN TIME:LIVER:DOCUMENT:XR.FLUOR
C0882011|T060||SNOMEDCT_US|LIVER CT BX CN GUID
C0882011|T060||SNOMEDCT_US|CT GUIDANCE FOR CORE NEEDLE BIOPSY OF LIVER
C0882011|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.CORE NEEDLE:FIND:PT:ABDOMEN>LIVER:DOC:CT
C0882011|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.CORE NEEDLE:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C3262906|T060||SNOMEDCT_US|ABD CT BX GUID WO CONTR
C3262906|T060||SNOMEDCT_US|CT GUIDANCE FOR BIOPSY OF ABDOMEN-- WO CONTRAST
C3262906|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY^WO CONTRAST:FIND:PT:ABDOMEN:DOC:CT
C3262906|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY^WO CONTRAST:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C0881937|T060||SNOMEDCT_US|LIVER FLR TJ BX GUID W CONTR IV
C0881937|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR TRANSJUGULAR BIOPSY OF LIVER-- W CONTRAST IV
C0881937|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.TRANSJUGULAR ^W CONTRAST IV:FIND:PT:LIVER:DOC:XR.FLUOR
C0881937|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.TRANSJUGULAR^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:LIVER:DOCUMENT:XR.FLUOR
C0882013|T060||SNOMEDCT_US|US GUIDANCE FOR BIOPSY OF LIVER
C0882013|T060||SNOMEDCT_US|LIVER US BX GUID
C0882013|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FINDING:POINT IN TIME:LIVER:DOCUMENT:ULTRASOUND
C0882013|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FIND:PT:LIVER:DOC:US
C1543445|T060||SNOMEDCT_US|LIVER FLR ABSCESS DRAIN GUID
C1543445|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR DRAINAGE OF ABSCESS OF LIVER
C1543445|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE OF ABSCESS:FIND:PT:LIVER:DOC:XR.FLUOR
C1543445|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE OF ABSCESS:FINDING:POINT IN TIME:LIVER:DOCUMENT:XR.FLUOR
C1631786|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE OF ABSCESS:FINDING:POINT IN TIME:ABDOMEN>LIVER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1631786|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE OF ABSCESS:FIND:PT:ABDOMEN>LIVER:DOC:CT
C1631786|T060||SNOMEDCT_US|CT GUIDANCE FOR DRAINAGE OF ABSCESS OF LIVER
C1631786|T060||SNOMEDCT_US|LIVER CT ABSCESS DRAIN GUID
C4039879|T060|708697000|SNOMEDCT_US|PERCUTANEOUS FINE NEEDLE ASPIRATION BIOPSY OF LIVER USING IMAGING GUIDANCE |PERCUTANEOUS FINE NEEDLE ASPIRATION BIOPSY OF LIVER USING IMAGING GUIDANCE
C4039879|T060|708697000|SNOMEDCT_US|PERCUTANEOUS FINE NEEDLE ASPIRATION BIOPSY OF LIVER USING IMAGING GUIDANCE|PERCUTANEOUS FINE NEEDLE ASPIRATION BIOPSY OF LIVER USING IMAGING GUIDANCE
C2584955|T060|438529005|SNOMEDCT_US|ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE |ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE
C2584955|T060|438529005|SNOMEDCT_US|MRI GUIDED ABLATION OF LIVER|ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE
C2584955|T060|438529005|SNOMEDCT_US|ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE|ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE
C2584862|T060|441138007|SNOMEDCT_US|FOCUSED ULTRASOUND ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE |FOCUSED ULTRASOUND ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE (PROCEDURE)
C2584862|T060|441138007|SNOMEDCT_US|FOCUSED ULTRASOUND ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE|FOCUSED ULTRASOUND ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE (PROCEDURE)
C2584862|T060|441138007|SNOMEDCT_US|MRI GUIDED FOCUSED ULTRASOUND ABLATION OF LIVER|FOCUSED ULTRASOUND ABLATION OF LIVER USING MAGNETIC RESONANCE IMAGING GUIDANCE (PROCEDURE)
C1715475|T060||SNOMEDCT_US|BDS FLR ENDO GUID W CONTR RETRO
C1715475|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR ENDOSCOPY OF BILIARY DUCTS-- W CONTRAST RETROGRADE
C1715475|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^W CONTRAST RETROGRADE:FINDING:POINT IN TIME:BILIARY DUCTS:DOCUMENT:XR.FLUOR
C1715475|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^W CONTRAST RETROGRADE:FIND:PT:BILIARY DUCTS:DOC:XR.FLUOR
C1714814|T060||SNOMEDCT_US|BD+PDS FLR ENDO GUID 1H P CONTR RETRO
C1714814|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR ENDOSCOPY OF BILIARY DUCTS AND PANCREATIC DUCT-- 1 HOUR POST CONTRAST RETROGRADE
C1714814|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^1 HOUR POST CONTRAST RETROGRADE:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:XR.FLUOR
C1714814|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^1H POST CONTRAST RETROGRADE:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:XR.FLUOR
C1714813|T060||SNOMEDCT_US|BD+PDS FLR ENDO GUID 45M P CONTR RETRO
C1714813|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR ENDOSCOPY OF BILIARY DUCTS AND PANCREATIC DUCT-- 45 MINUTES POST CONTRAST RETROGRADE
C1714813|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^45M POST CONTRAST RETROGRADE:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:XR.FLUOR
C1714813|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^45M POST CONTRAST RETROGRADE:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:XR.FLUOR
C1714815|T060||SNOMEDCT_US|BD+PDS FLR ENDO GUID 1.5H P CONTR RETRO
C1714815|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR ENDOSCOPY OF BILIARY DUCTS AND PANCREATIC DUCT-- 1.5 HOURS POST CONTRAST RETROGRADE
C1714815|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^1 1/2 HOUR POST CONTRAST RETROGRADE:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:XR.FLUOR
C1714815|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^1.5H POST CONTRAST RETROGRADE:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:XR.FLUOR
C1114616|T060||SNOMEDCT_US|BD+PDS FLR ENDO GUID W CONTR RETRO
C1114616|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR ENDOSCOPY OF BILIARY DUCTS AND PANCREATIC DUCT-- W CONTRAST RETROGRADE
C1114616|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^W CONTRAST RETROGRADE:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:XR.FLUOR
C1114616|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^W CONTRAST RETROGRADE:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:XR.FLUOR
C1830086|T060||SNOMEDCT_US|BDS FLR PC DRAIN GUID
C1830086|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR PERCUTANEOUS DRAINAGE OF BILIARY DUCTS
C1830086|T060||SNOMEDCT_US|GUIDANCE FOR PERCUTANEOUS DRAINAGE:FINDING:POINT IN TIME:BILIARY DUCTS:DOCUMENT:XR.FLUOR
C1830086|T060||SNOMEDCT_US|GUIDANCE FOR PERCUTANEOUS DRAINAGE:FIND:PT:BILIARY DUCTS:DOC:XR.FLUOR
C1525098|T060||SNOMEDCT_US|BDS+GB CT DRAIN GUID
C1525098|T060||SNOMEDCT_US|CT GUIDANCE FOR DRAINAGE OF BILIARY DUCTS AND GALLBLADDER
C1525098|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE:FIND:PT:ABDOMEN>BILIARY DUCTS+GALLBLADDER:DOC:CT
C1525098|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE:FINDING:POINT IN TIME:ABDOMEN>BILIARY DUCTS+GALLBLADDER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1714811|T060||SNOMEDCT_US|BD+PDS FLR ENDO GUID 15M P CONTR RETRO
C1714811|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR ENDOSCOPY OF BILIARY DUCTS AND PANCREATIC DUCT-- 15 MINUTES POST CONTRAST RETROGRADE
C1714811|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^15 MINUTES POST CONTRAST RETROGRADE:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:XR.FLUOR
C1714811|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^15M POST CONTRAST RETROGRADE:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:XR.FLUOR
C1714812|T060||SNOMEDCT_US|BD+PDS FLR ENDO GUID 30M P CONTR RETRO
C1714812|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR ENDOSCOPY OF BILIARY DUCTS AND PANCREATIC DUCT-- 30 MINUTES POST CONTRAST RETROGRADE
C1714812|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^30 MINUTES POST CONTRAST RETROGRADE:FINDING:POINT IN TIME:BILIARY DUCTS+PANCREATIC DUCT:DOCUMENT:XR.FLUOR
C1714812|T060||SNOMEDCT_US|GUIDANCE FOR ENDOSCOPY^30M POST CONTRAST RETROGRADE:FIND:PT:BILIARY DUCTS+PANCREATIC DUCT:DOC:XR.FLUOR
C0881809|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR STONE REMOVAL OF BILIARY DUCT COMMON-- W CONTRAST INTRA BILIARY DUCT
C0881809|T060||SNOMEDCT_US|CBD FLR STONE REM GUID W CONTR INTRA BD
C0881809|T060||SNOMEDCT_US|GUIDANCE FOR STONE REMOVAL^W CONTRAST INTRA BILIARY DUCT:FIND:PT:BILIARY DUCT.COMMON:DOC:XR.FLUOR
C0881809|T060||SNOMEDCT_US|GUIDANCE FOR STONE REMOVAL^W CONTRAST INTRA BILIARY DUCT:FINDING:POINT IN TIME:BILIARY DUCT.COMMON:DOCUMENT:XR.FLUOR
C0881810|T060||SNOMEDCT_US|BDS+GB RI FOR BIL PAT W TC99MIV
C0881810|T060||SNOMEDCT_US|BILIARY DUCTS AND GALLBLADDER SCAN FOR PATENCY OF BILIARY STRUCTURES W TC-99M IV
C0881810|T060||SNOMEDCT_US|VIEWS FOR PATENCY OF BILIARY STRUCTURES^W TC-99M IV:FIND:PT:BILIARY DUCTS+GALLBLADDER:DOC:RADNUC
C0881810|T060||SNOMEDCT_US|VIEWS FOR PATENCY OF BILIARY STRUCTURES^W TC-99M INTRAVENOUS:FINDING:POINT IN TIME:BILIARY DUCTS+GALLBLADDER:DOCUMENT:RADNUC
C0881813|T060||SNOMEDCT_US|BDS+GB FLR W CONTR PC TRANSHEPATIC
C0881813|T060||SNOMEDCT_US|BILIARY DUCTS AND GALLBLADDER FLUOROSCOPY W CONTRAST PERCUTANEOUS TRANSHEPATIC
C0881813|T060||SNOMEDCT_US|VIEWS^W CONTRAST PERCUTANEOUS TRANSHEPATIC:FINDING:POINT IN TIME:BILIARY DUCTS+GALLBLADDER:DOCUMENT:XR.FLUOR
C0881813|T060||SNOMEDCT_US|VIEWS^W CONTRAST PERCUTANEOUS TRANSHEPATIC:FIND:PT:BILIARY DUCTS+GALLBLADDER:DOC:XR.FLUOR
C3533557|T060||SNOMEDCT_US|GUIDANCE FOR REPLACEMENT OF PERCUTANEOUS DRAINAGE TUBE:FINDING:POINT IN TIME:BILIARY DUCTS+GALLBLADDER:DOCUMENT:XR.FLUOR
C3533557|T060||SNOMEDCT_US|GUIDANCE FOR REPLACEMENT OF PERCUTANEOUS DRAINAGE TUBE:FIND:PT:BILIARY DUCTS+GALLBLADDER:DOC:XR.FLUOR
C3533557|T060||SNOMEDCT_US|BDS+GB FLR REPLAC OF PC DRAIN TUBE GUID
C3533557|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR REPLACEMENT OF PERCUTANEOUS DRAINAGE TUBE IN BILIARY DUCTS AND GALLBLADDER
C0400529|T060|174653005|SNOMEDCT_US|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY AND COLLECTION OF PANCREATIC JUICE|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY AND COLLECTION OF PANCREATIC JUICE (PROCEDURE)
C0400529|T060|174653005|SNOMEDCT_US|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY AND COLLECTION OF PANCREATIC JUICE |ENDOSCOPIC RETROGRADE PANCREATOGRAPHY AND COLLECTION OF PANCREATIC JUICE (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|X-RAY GASTROINTESTINAL EPR|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY |ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|ENDOSC RETRO PANCREATOG|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF PANCREATIC DUCT NOS |ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF PANCREATIC DUCT NOS|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|ERP|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|ERP - ENDOSCOPIC RETROGRADE PANCREATOGRAPHY|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF PANCREATIC DUCT|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0337380|T060|174651007|SNOMEDCT_US|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY [ERP]|ENDOSCOPIC RETROGRADE PANCREATOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|ENDOSC RETRO CHOLANGIO|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|ERC|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF BILE DUCT NOS|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF BILE DUCT NOS |ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|ERC - ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY |ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF BILE DUCT|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF BILE DUCT |ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|ERC, NOS|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193504|T060|386722005|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY [ERC]|ENDOSCOPIC RETROGRADE CHOLANGIOGRAPHY (PROCEDURE)
C0193505|T060|6157006|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP); WITH BIOPSY, SINGLE OR MULTIPLE|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY (PROCEDURE)
C0193505|T060|6157006|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP) WITH BIOPSY|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY (PROCEDURE)
C0193505|T060|6157006|SNOMEDCT_US|ERCP W/BIOPSY SINGLE/MULTIPLE|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY (PROCEDURE)
C0193505|T060|6157006|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY (PROCEDURE)
C0193505|T060|6157006|SNOMEDCT_US|ERCP WITH BIOPSY|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY (PROCEDURE)
C0193505|T060|6157006|SNOMEDCT_US|ERCP WITH BIOPSY |ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY (PROCEDURE)
C0193505|T060|6157006|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY |ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY (PROCEDURE)
C0193505|T060|6157006|SNOMEDCT_US|ENDO CHOLANGIOPANCREATOGRAPH|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY WITH BIOPSY (PROCEDURE)
C0193527|T060|53054006|SNOMEDCT_US|LAPAROSCOPY WITH GUIDED TRANSHEPATIC CHOLANGIOGRAPHY|LAPAROSCOPY WITH GUIDED TRANSHEPATIC CHOLANGIOGRAPHY (PROCEDURE)
C0193527|T060|53054006|SNOMEDCT_US|LAPAROSCOPY WITH GUIDED TRANSHEPATIC CHOLANGIOGRAPHY |LAPAROSCOPY WITH GUIDED TRANSHEPATIC CHOLANGIOGRAPHY (PROCEDURE)
C0008310|T060|386718000|SNOMEDCT_US|CHOLANGIOPANCREATOGRAPHIES, ENDOSCOPIC RETROGRADE|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|CHOLANGIOPANCREATOGRAPHY, ENDOSCOPIC RETROGRADE|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHIES|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|RETROGRADE CHOLANGIOPANCREATOGRAPHIES, ENDOSCOPIC|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|CHOLANGIOPANCREATOGR ENDOSCOPIC RETROGRADE|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGR|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|RETROGRADE CHOLANGIOPANCREATOGR ENDOSCOPIC|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ERCP (ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY)|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY -RETIRED-|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSC RETRO CHOLANGIOPA|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY |ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY |ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ERCP|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF BILE DUCT AND PANCREATIC DUCT NOS|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF BILE DUCT AND PANCREATIC DUCT|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ERCP - ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF BILE DUCT AND PANCREATIC DUCT NOS |ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP)|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|RETROGRADE CHOLANGIOPANCREATOGRAPHY, ENDOSCOPIC|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC CATHETERIZATION OF PANCREATIC DUCT AND BILE DUCT SYSTEMS|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|DIAGNOSTIC ENDOSCOPIC RETROGRADE EXAMINATION OF BILE DUCT AND PANCREATIC DUCT |ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC CATHETERISATION OF PANCREATIC DUCT AND BILE DUCT SYSTEMS|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC CATHETERIZATION OF PANCREATIC DUCT AND BILE DUCT SYSTEMS |ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY, NOS|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ERCP, NOS|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY  [AMBIGUOUS]|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0008310|T060|386718000|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY [ERCP]|ENDOSCOPIC RETROGRADE CHOLEDOCHOPANCREATOGRAPHY
C0177739|T060||SNOMEDCT_US|PERC HEPAT CHOLANGIOGRAM
C0177739|T060||SNOMEDCT_US|PERCUTANEOUS HEPATIC CHOLANGIOGRAM
C0400786|T060|235583009|SNOMEDCT_US|ERCP SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL |ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP) SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL
C0400786|T060|235583009|SNOMEDCT_US|ERCP SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP) SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL
C0400786|T060|235583009|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL |ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP) SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL
C0400786|T060|235583009|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP) SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL
C0400786|T060|235583009|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP) SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP) SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL
C0400786|T060|235583009|SNOMEDCT_US|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP) SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL |ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGRAPHY (ERCP) SPHINCTEROTOMY SPHINCTER OF ODDI AND CALCULUS REMOVAL
C1633404|T060||SNOMEDCT_US|PORTAL V XRA CATH PLAC GUID W CONTR IV
C1633404|T060||SNOMEDCT_US|FLUOROSCOPIC ANGIOGRAM GUIDANCE FOR PLACEMENT OF CATHETER IN PORTAL VEIN-- W CONTRAST IV
C1633404|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF CATHETER^W CONTRAST IV:FIND:PT:PORTAL VEIN:DOC:XR.FLUOR.ANGIO
C1633404|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF CATHETER^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:PORTAL VEIN:DOCUMENT:XR.FLUOR.ANGIO
C1632228|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF INFUSION PORT:FIND:PT:HEPATIC ARTERY:NAR:RADNUC
C1632228|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF INFUSION PORT:FINDING:POINT IN TIME:HEPATIC ARTERY:NARRATIVE:RADNUC
C1632228|T060||SNOMEDCT_US|DEPRECATED SCAN GUIDANCE FOR PLACEMENT OF INFUSION PORT IN HEPATIC ARTERY
C1632228|T060||SNOMEDCT_US|DEPRECATED HEP A RI INFUSION PORT PLAC G
C0884114|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR PLACEMENT OF STENT IN INTRAHEPATIC PORTAL SYSTEM
C0884114|T060||SNOMEDCT_US|IHP FLR STENT PLAC GUID
C0884114|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF STENT:FIND:PT:INTRAHEPATIC PORTAL SYSTEM:DOC:XR.FLUOR
C0884114|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF STENT:FINDING:POINT IN TIME:INTRAHEPATIC PORTAL SYSTEM:DOCUMENT:XR.FLUOR
C1978441|T060||SNOMEDCT_US|PORTAL+HEPATIC V XRA TIPS PLAC GUID
C1978441|T060||SNOMEDCT_US|FLUOROSCOPIC ANGIOGRAM GUIDANCE FOR PLACEMENT OF TRANSJUGULAR INTRAHEPATIC PORTOSYSTEMIC SHUNT IN PORTAL VEIN AND HEPATIC VEIN
C1978441|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF TRANSJUGULAR INTRAHEPATIC PORTOSYSTEMIC SHUNT:FIND:PT:PORTAL VEIN+HEPATIC VEIN:DOC:XR.FLUOR.ANGIO
C1978441|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF TRANSJUGULAR INTRAHEPATIC PORTOSYSTEMIC SHUNT:FINDING:POINT IN TIME:PORTAL VEIN+HEPATIC VEIN:DOCUMENT:XR.FLUOR.ANGIO
C0882225|T060||SNOMEDCT_US|HEP A XRA CATH PLAC GUID W CONTR IA
C0882225|T060||SNOMEDCT_US|FLUOROSCOPIC ANGIOGRAM GUIDANCE FOR PLACEMENT OF CATHETER IN HEPATIC ARTERY-- W CONTRAST IA
C0882225|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF CATHETER^W CONTRAST INTRA-ARTERIAL:FINDING:POINT IN TIME:HEPATIC ARTERY:DOCUMENT:XR.FLUOR.ANGIO
C0882225|T060||SNOMEDCT_US|GUIDANCE FOR PLACEMENT OF CATHETER^W CONTRAST IA:FIND:PT:HEPATIC ARTERY:DOC:XR.FLUOR.ANGIO
C1524281|T060||SNOMEDCT_US|IVC XRA ANGPSTY W CONTR IV
C1524281|T060||SNOMEDCT_US|INFERIOR VENA CAVA FLUOROSCOPIC ANGIOGRAM ANGIOPLASTY W CONTRAST IV
C1524281|T060||SNOMEDCT_US|ANGIOPLASTY^W CONTRAST INTRAVENOUS:FINDING:POINT IN TIME:VENA CAVA.INFERIOR:DOCUMENT:XR.FLUOR.ANGIO
C1524281|T060||SNOMEDCT_US|ANGIOPLASTY^W CONTRAST IV:FIND:PT:VENA CAVA.INFERIOR:DOC:XR.FLUOR.ANGIO
C1715409|T060||SNOMEDCT_US|PET WB
C1715409|T060||SNOMEDCT_US|PET WHOLE BODY
C1715409|T060||SNOMEDCT_US|MULTISECTION WHOLE BODY:FINDING:POINT IN TIME:^PATIENT:DOCUMENT:RADNUC.PET
C1715409|T060||SNOMEDCT_US|MULTISECTION WHOLE BODY:FIND:PT:^PATIENT:DOC:RADNUC.PET
C3263050|T060||SNOMEDCT_US|SPECT FOR TUMOR WB W RNC IV
C3263050|T060||SNOMEDCT_US|SPECT FOR TUMOR WHOLE BODY
C3263050|T060||SNOMEDCT_US|MULTISECTION FOR TUMOR WHOLE BODY^W RADIONUCLIDE IV:FIND:PT:^PATIENT:DOC:RADNUC.SPECT
C3263050|T060||SNOMEDCT_US|MULTISECTION FOR TUMOR WHOLE BODY^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:^PATIENT:DOCUMENT:RADNUC.SPECT
C1648951|T060||SNOMEDCT_US|SPECT WB W TC99MCEA IV
C1648951|T060||SNOMEDCT_US|SPECT WHOLE BODY W TC-99M ARCITUMOMAB IV
C1648951|T060||SNOMEDCT_US|MULTISECTION WHOLE BODY^W TC-99M ARCITUMOMAB INTRAVENOUS:FINDING:POINT IN TIME:^PATIENT:DOCUMENT:RADNUC.SPECT
C1648951|T060||SNOMEDCT_US|MULTISECTION WHOLE BODY^W TC-99M ARCITUMOMAB IV:FIND:PT:^PATIENT:DOC:RADNUC.SPECT
C1830259|T060||SNOMEDCT_US|MULTISECTION WHOLE BODY:FINDING:POINT IN TIME:^PATIENT:NARRATIVE:MRI
C1830259|T060||SNOMEDCT_US|MRI WHOLE BODY
C1830259|T060||SNOMEDCT_US|MRI WB
C1830259|T060||SNOMEDCT_US|MULTISECTION WHOLE BODY:FINDING:POINT IN TIME:^PATIENT:DOCUMENT:MRI
C1830259|T060||SNOMEDCT_US|MULTISECTION WHOLE BODY:FIND:PT:^PATIENT:DOC:MRI
C1714784|T060||SNOMEDCT_US|MULTISECTION FOR TUMOR WHOLE BODY:FIND:PT:^PATIENT:DOC:CT
C1714784|T060||SNOMEDCT_US|DEPRECATED CT FOR TUMOR WHOLE BODY
C1714784|T060||SNOMEDCT_US|MULTISECTION FOR TUMOR WHOLE BODY:FINDING:POINT IN TIME:^PATIENT:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1714784|T060||SNOMEDCT_US|DEPRECATED CT FOR TUMOR WB
C1542855|T060||SNOMEDCT_US|RI FOR TUMOR MUL AREAS W GA-67 IV
C1542855|T060||SNOMEDCT_US|VIEWS FOR TUMOR MULTIPLE AREAS^W GA-67 INTRAVENOUS:FINDING:POINT IN TIME:^PATIENT:DOCUMENT:RADNUC
C1542855|T060||SNOMEDCT_US|VIEWS FOR TUMOR MULTIPLE AREAS^W GA-67 IV:FIND:PT:^PATIENT:DOC:RADNUC
C1542855|T060||SNOMEDCT_US|SCAN FOR TUMOR MULTIPLE AREAS W GA-67 IV
C1626178|T060||SNOMEDCT_US|SCAN WHOLE BODY
C1626178|T060||SNOMEDCT_US|RI WB W RNC IV
C1626178|T060||SNOMEDCT_US|VIEWS WHOLE BODY^W RADIONUCLIDE IV:FIND:PT:^PATIENT:DOC:RADNUC
C1626178|T060||SNOMEDCT_US|VIEWS WHOLE BODY^W RADIONUCLIDE INTRAVENOUS:FINDING:POINT IN TIME:^PATIENT:DOCUMENT:RADNUC
C1543801|T060||SNOMEDCT_US|RI FOR TUMOR WB W TC99MMIBI IV
C1543801|T060||SNOMEDCT_US|SCAN FOR TUMOR WHOLE BODY W TC-99M SESTAMIBI IV
C1543801|T060||SNOMEDCT_US|VIEWS FOR TUMOR WHOLE BODY^W TC-99M SESTAMIBI INTRAVENOUS:FINDING:POINT IN TIME:^PATIENT:DOCUMENT:RADNUC
C1543801|T060||SNOMEDCT_US|VIEWS FOR TUMOR WHOLE BODY^W TC-99M SESTAMIBI IV:FIND:PT:^PATIENT:DOC:RADNUC
C1830206|T060||SNOMEDCT_US|WHOLE BODY CT
C1830206|T060||SNOMEDCT_US|MULTISECTION:FINDING:POINT IN TIME:WHOLE BODY:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1830206|T060||SNOMEDCT_US|MULTISECTION:FIND:PT:WHOLE BODY:DOC:CT
C0032743|T060|363678002|SNOMEDCT_US|POSITRON-EMISSION TOMOGRAPHY|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHY|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|PETT|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISS TOMOGR|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|TOMOGR POSITRON EMISS|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHIC IMAGING|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|PET SCAN|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|PET|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHY |POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISSION TOMOGRAM|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|IMAGING, PET|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|PET IMAGING|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|PET SCANS|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|PROTON MAGNETIC RESONANCE SPECTROSCOPIC IMAGING|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHY SCAN|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|TOMOGRAPHY, POSITRON-EMISSION|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|PET - POSITRON EMISSION TOMOGRAPHY|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION (QUALIFIER VALUE)|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHY, NOS|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|PET SCAN, NOS|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|SCAN, PET|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|SCANS, PET|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|TOMOGRAPHY, POSITRON EMISSION|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|MEDICAL IMAGING, POSITRON EMISSION TOMOGRAPHY|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C0032743|T060|363678002|SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHY (PET)|POSITRON EMISSION TOMOGRAPHIC IMAGING - ACTION
C2729424|T060||SNOMEDCT_US|PET TUMOR INIT TX STRAT
C2729424|T060||SNOMEDCT_US|POSITRON EMISSION TOMOGRAPHY (PET) OR PET/COMPUTED TOMOGRAPHY (CT) TO INFORM THE INITIAL TREATMENT STRATEGY OF TUMORS THAT ARE BIOPSY PROVEN OR STRONGLY SUSPECTED OF BEING CANCEROUS BASED ON OTHER DIAGNOSTIC TESTING
C0203669|T060|367385006|SNOMEDCT_US|WHOLE BODY SCANNING|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|TOTAL BODY SCAN|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|WHOLE BODY SCAN|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|WHOLE BODY IMAGING|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|TOTAL BODY SCAN |TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|SCAN NOS WHOLE BODY|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|RADIOISOTOPE SCAN OF TOTAL BODY|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|RADIOISOTOPE SCAN OF TOTAL BODY |TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|TOTAL BODY SCAN  [AMBIGUOUS]|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|IMAGING, WHOLE BODY|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|IMAGINGS, WHOLE BODY|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|SCAN, WHOLE BODY|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|SCANS, WHOLE BODY|TOTAL BODY SCAN (PROCEDURE)
C0203669|T060|367385006|SNOMEDCT_US|WHOLE BODY IMAGINGS|TOTAL BODY SCAN (PROCEDURE)
C1715435|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE OF ABSCESS:FINDING:POINT IN TIME:PERITONEAL SPACE:DOCUMENT:ULTRASOUND
C1715435|T060||SNOMEDCT_US|PERITONEAL SPACE US ABSCESS DRAIN GUID
C1715435|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE OF ABSCESS:FIND:PT:PERITONEAL SPACE:DOC:US
C1715435|T060||SNOMEDCT_US|US GUIDANCE FOR DRAINAGE OF ABSCESS OF PERITONEAL SPACE
C1645316|T060||SNOMEDCT_US|GUIDANCE FOR REMOVAL OF FLUID:FIND:PT:ABDOMEN:DOC:CT
C1645316|T060||SNOMEDCT_US|DEPRECATED CT GUIDANCE FOR REMOVAL OF FLUID FROM ABDOMEN
C1645316|T060||SNOMEDCT_US|GUIDANCE FOR REMOVAL OF FLUID:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1645316|T060||SNOMEDCT_US|DEPRECATED ABD CT FLD REM GUID
C1525261|T060||SNOMEDCT_US|ABD CT ASP+DRAIN TUBE PLAC GUID
C1525261|T060||SNOMEDCT_US|CT GUIDANCE FOR ASPIRATION AND PLACEMENT OF DRAINAGE TUBE OF ABDOMEN
C1525261|T060||SNOMEDCT_US|GUIDANCE FOR ASPIRATION & PLACEMENT OF DRAINAGE TUBE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1525261|T060||SNOMEDCT_US|GUIDANCE FOR ASPIRATION & PLACEMENT OF DRAINAGE TUBE:FIND:PT:ABDOMEN:DOC:CT
C3263037|T060||SNOMEDCT_US|ABD FLR BX NEEDLE GUID
C3263037|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR NEEDLE BIOPSY OF ABDOMEN
C3263037|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.NEEDLE:FIND:PT:ABDOMEN:DOC:XR.FLUOR
C3263037|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY.NEEDLE:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR.FLUOR
C1524289|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR BIOPSY OF ABDOMEN
C1524289|T060||SNOMEDCT_US|ABD FLR BX GUID
C1524289|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR.FLUOR
C1524289|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FIND:PT:ABDOMEN:DOC:XR.FLUOR
C1526193|T060||SNOMEDCT_US|ABD US BX GUID
C1526193|T060||SNOMEDCT_US|US GUIDANCE FOR BIOPSY OF ABDOMEN
C1526193|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FIND:PT:ABDOMEN:DOC:US
C1526193|T060||SNOMEDCT_US|GUIDANCE FOR BIOPSY:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:ULTRASOUND
C1639941|T060||SNOMEDCT_US|ABD FLR REPLAC OF PCS GUID
C1639941|T060||SNOMEDCT_US|FLUOROSCOPY GUIDANCE FOR REPLACEMENT OF PERCUTANEOUS CHOLECYSTOSTOMY IN ABDOMEN
C1639941|T060||SNOMEDCT_US|GUIDANCE FOR REPLACEMENT OF PERCUTANEOUS CHOLECYSTOSTOMY:FIND:PT:ABDOMEN:DOC:XR.FLUOR
C1639941|T060||SNOMEDCT_US|GUIDANCE FOR REPLACEMENT OF PERCUTANEOUS CHOLECYSTOSTOMY:FINDING:POINT IN TIME:ABDOMEN:DOCUMENT:XR.FLUOR
C1524316|T060||SNOMEDCT_US|ABD GB CT DRAIN GUID
C1524316|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE:FIND:PT:ABDOMEN>GALLBLADDER:DOC:CT
C1524316|T060||SNOMEDCT_US|GUIDANCE FOR DRAINAGE:FINDING:POINT IN TIME:ABDOMEN>GALLBLADDER:DOCUMENT:COMPUTERIZED TOMOGRAPHY
C1114635|T060||SNOMEDCT_US|VISCERAL ARTERY FLUOROSCOPIC ANGIOGRAM ANGIOPLASTY W CONTRAST IA
C1114635|T060||SNOMEDCT_US|VISCERAL A XRA ANGPSTY W CONTR IA
C1114635|T060||SNOMEDCT_US|ANGIOPLASTY^W CONTRAST IA:FIND:PT:VISCERAL ARTERY:DOC:XR.FLUOR.ANGIO
C1114635|T060||SNOMEDCT_US|ANGIOPLASTY^W CONTRAST INTRA-ARTERIAL:FINDING:POINT IN TIME:VISCERAL ARTERY:DOCUMENT:XR.FLUOR.ANGIO
