C0019682|T047|19030005|SNOMEDCT_US|HIV|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019693|T047|123321001|SNOMEDCT_US|HIV INFECTIONS|HTLV-III/LAV INFECTION (DISORDER)
C0019704|T047|243598007|SNOMEDCT_US|HIV-1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS 1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|AIDS VIRUS|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFIC VIRUS 1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS 001|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFIC VIRUS TYPE 1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HIV 01|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|IMMUNODEFIC VIRUS TYPE 1 HUMAN|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HIV 1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN T CELL LEUKEMIA VIRUS III|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE I -RETIRED-|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS 1 HIV-1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS HIV-1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 HIV 1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 HIV-1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 HIV1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1, HIV-1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE I HIV-1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE-1 HIV-1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-1 HIV-1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE I|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HIV1 - HUMAN IMMUNODEFICIENCY VIRUS TYPE 1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE I |HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 |HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|OLD NAME, BUT AT LEAST STILL REFERS TO THE RIGHT VIRUS|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN T-CELL LEUKAEMIA VIRUS III|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN T-CELL LEUKEMIA VIRUS III|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|IMMUNODEFICIENCY VIRUS TYPE 1, HUMAN|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HIV-I|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HIV1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 [AMBIGUOUS]|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019704|T047|243598007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS, TYPE 1|HUMAN IMMUNODEFICIENCY VIRUS TYPE 1 (ORGANISM)
C0019707|T047|123188003|SNOMEDCT_US|HIV-2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS 2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|IMMUNODEFIC VIRUS TYPE 2 HUMAN|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|LAV AA 02|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFIC VIRUS 2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFIC VIRUS TYPE 2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HIV 02|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HTLV WIV|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN LYMPHOTROPIC VIRUS TYPE IV A T|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS 002|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HIV 2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS 2 (HIV-2)|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 HIV-2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2, HIV-2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 |HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|LAV-2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|IMMUNODEFICIENCY VIRUS TYPE 2, HUMAN|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HIV-II|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HIV TYPE 2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HIV2 - HUMAN IMMUNODEFICIENCY VIRUS TYPE 2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HIV2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019707|T047|123188003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS, TYPE 2|HUMAN IMMUNODEFICIENCY VIRUS TYPE 2 -RETIRED-
C0019682|T047|19030005|SNOMEDCT_US|HIV|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|LYMPHADENOPATHY ASSOCIATED VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|LYMPHADENOPATHY-ASSOCIATED VIRUSES|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUS, LYMPHADENOPATHY-ASSOCIATED|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUSES, LYMPHADENOPATHY-ASSOCIATED|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HUMAN IMMUNODEFIC VIRUSES|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|IMMUNODEFIC VIRUSES HUMAN|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUS HUMAN IMMUNODEFIC|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HUMAN IMMUNODEFIC VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUSES HUMAN IMMUNODEFIC|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|IMMUNODEFIC VIRUS HUMAN|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|LAV|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS, NOS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HUMAN T CELL LEUKEMIA VIRUS TYPE III|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUS (HIV), HUMAN IMMUNODEFICIENCY|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV)|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HIV, HUMAN IMMUNODEFICIENCY VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|IMMUNODEFICIENCY VIRUSES, HUMAN|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|LAV-HTLV-III|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HUMAN T-CELL LEUKEMIA VIRUS TYPE III|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|IMMUNODEFICIENCY VIRUS, HUMAN|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|AIDS VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUSES|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|LYMPHADENOPATHY-ASSOCIATED VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUS, HUMAN IMMUNODEFICIENCY|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUSES, HUMAN IMMUNODEFICIENCY|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS |HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|LYMPHADENOPATHY-ASSOCIATED VIRUS (LAV)|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|LYMPHADENOPATHY-ASSOCIATED VIRUS, TYPE I (LAV-I)|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|AIDS VIRUSES|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUS, AIDS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUSES, AIDS|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0019682|T047|19030005|SNOMEDCT_US|VIRUS-HIV|HUMAN IMMUNODEFICIENCY VIRUS (ORGANISM)
C0497169|T047||SNOMEDCT_US|HIV/AIDS
C1989665|T047||SNOMEDCT_US|HIV PHENOTYPE &#X7C; ISOLATE
C1954120|T047||SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS GENOTYPE:SUSCEPTIBILITY:POINT IN TIME:ISOLATE:NOMINAL:GENOTYPING
C1954120|T047||SNOMEDCT_US|HIV GENTYP ISLT
C1954120|T047||SNOMEDCT_US|HIV GENOTYPE:SUSC:PT:ISOLATE:NOM:GENOTYPING
C1954120|T047||SNOMEDCT_US|HIV GENOTYPE [SUSCEPTIBILITY]
C0369501|T047||SNOMEDCT_US|HIV IDENTIFIED
C0369501|T047||SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS IDENTIFIED
C3534218|T047||SNOMEDCT_US|HIV 1 INTEGRASE GENE &#X7C; ISOLATE
C1440749|T047||SNOMEDCT_US|HIV REVERSE TRANSCRIPTASE+PROTEASE GENE
C1440733|T047||SNOMEDCT_US|HIV 1+2
C1440733|T047||SNOMEDCT_US|HIV 1 & 2
C1977331|T047||SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS GENOTYPE:SUSCEPTIBILITY:POINT IN TIME:ISOLATE:NARRATIVE:GENOTYPING
C1977331|T047||SNOMEDCT_US|HIV GENOTYPE:SUSC:PT:ISOLATE:NAR:GENOTYPING
C1977331|T047||SNOMEDCT_US|HIV GENOTYPE [SUSCEPTIBILITY] IN ISOLATE BY GENOTYPE METHOD NARRATIVE
C1977331|T047||SNOMEDCT_US|HIV GENTYP ISLT NAR
C3656356|T047||SNOMEDCT_US|HIV REVERSE TRANSCRIPTASE+PROTEASE+INTEGRASE GENE
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNO DEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNO-DEFICIENCY SYNDROMES|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROMES|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|AIDS|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|IMMUNO-DEFICIENCY SYNDROME, ACQUIRED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|IMMUNO-DEFICIENCY SYNDROMES, ACQUIRED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|IMMUNODEFICIENCY SYNDROMES, ACQUIRED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|SYNDROME, ACQUIRED IMMUNO-DEFICIENCY|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|SYNDROME, ACQUIRED IMMUNODEFICIENCY|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|SYNDROMES, ACQUIRED IMMUNO-DEFICIENCY|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|SYNDROMES, ACQUIRED IMMUNODEFICIENCY|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|AIDS |ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME (AIDS)|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|IMMUNODEFIC SYNDROME ACQUIRED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNO DEFIC SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFIC SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|IMMUNOL DEFIC SYNDROME ACQUIRED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFIC SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (HIV-1 STAGE 6)|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) |ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS)|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDR|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME [AIDS]|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME [DISEASE/FINDING]|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|IMMUNODEFICIENCY SYNDROME, ACQUIRED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNO-DEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|IMMUNOLOGIC DEFICIENCY SYNDROME, ACQUIRED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME |ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFIC. SYND.|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED HUMAN IMMUNODEFICIENCY VIRUS INFECTION SYNDROME NOS|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED HUMAN IMMUNODEFICIENCY VIRUS INFECTION SYNDROME NOS |ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFIC. SYNDR.|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME (AIDS) |ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY DISEASE|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|AIDS, ACQUIRED IMMUNODEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME, AIDS|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME NOS|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME, UNSPECIFIED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|AUTOIMMUNE DEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|AIDS - ACQUIRED IMMUNODEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|IMMUNODEFICIENCY DUE TO HUMAN IMMUNODEFICIENCY VIRUS INFECTION|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED; IMMUNODEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|AIDS, NOS|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME, NOS|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME, NOS|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0001175|T047|62479008|SNOMEDCT_US|ACQUIRED IMMUN-DEFICIENCY SYND|ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0596049|T047||SNOMEDCT_US|AIDS/HIV NEUROPATHY
C0019693|T047|123321001|SNOMEDCT_US|HIV INFECTION|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HIV INFECTIONS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV III LAV INFECTIONS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|INFECTION, HIV|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|INFECTION, HTLV-III-LAV|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|INFECTIONS, HIV|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|INFECTIONS, HTLV-III-LAV|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|UNSPECIFIED HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV III INFECT|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV WIII LAV INFECTIONS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV WIII INFECTIONS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HIV INFECT|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV III LAV INFECT|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV-III/LAV INFECTION, NOS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION |HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV-III/LAV INFECTION -RETIRED-|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|LYMPHADENOPATHY-ASSOCIATED VIRUS |HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|LYMPHADENOPATHY-ASSOCIATED VIRUS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION, UNSPECIFIED|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNO VIRUS DIS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HIV INFECTIONS [DISEASE/FINDING]|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV-III-LAV INFECTIONS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|INFECTION;HIV|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE (B20)|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV-III-LAV INFECTION|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|[X]HUMAN IMMUNODEFICIENCY VIRUS DISEASE |HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV-III/LAV INFECTION|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|[X]UNSPECIFIED HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|[X]UNSPECIFIED HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE |HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|[X]HUMAN IMMUNODEFICIENCY VIRUS DISEASE|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HTLV-III/LAV INFECTION |HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HIV|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS SYNDROME|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HIV DISEASE|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HIV INFECTION NOS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS INFECTION|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION |HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HIV DISEASE; DISEASE (I.E. CAUSED BY HIV DISEASE)|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HIV DISEASE; INFECTION|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|DISEASE (OR DISORDER); HIV DISEASE (RESULTING FROM HIV DISEASE)|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|DISEASE (OR DISORDER); RESULTING FROM HIV DISEASE|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS; DISEASE|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|IMMUNODEFICIENCY VIRUS DISEASE; HUMAN|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|INFECTION; HIV DISEASE AS CAUSE|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION, NOS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE|HTLV-III/LAV INFECTION (DISORDER)
C0019693|T047|123321001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS [HIV] INFECTION|HTLV-III/LAV INFECTION (DISORDER)
C0348209|T047|187445009|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER INFECTIOUS AND PARASITIC DISEASES|[X]HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS AND PARASITIC DISEASE (DISORDER)
C0348209|T047|187445009|SNOMEDCT_US|HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS OR PARASITIC DISEASE|[X]HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS AND PARASITIC DISEASE (DISORDER)
C0348209|T047|187445009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE RESULTING IN INFECTIOUS AND PARASITIC DISEASES|[X]HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS AND PARASITIC DISEASE (DISORDER)
C0348209|T047|187445009|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS AND PARASITIC DISEASE|[X]HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS AND PARASITIC DISEASE (DISORDER)
C0348209|T047|187445009|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS AND PARASITIC DISEASE |[X]HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS AND PARASITIC DISEASE (DISORDER)
C0348209|T047|187445009|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER INFECTIOUS AND PARASITIC DISEASES|[X]HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS AND PARASITIC DISEASE (DISORDER)
C0348209|T047|187445009|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER INFECTIOUS AND PARASITIC DISEASES |[X]HIV DISEASE RESULTING IN UNSPECIFIED INFECTIOUS AND PARASITIC DISEASE (DISORDER)
C0348213|T047|187449003|SNOMEDCT_US|HIV DISEASE RESULTING IN UNSPECIFIED MALIGNANT NEOPLASM|[X]HIV DISEASE RESULTING IN UNSPECIFIED MALIGNANT NEOPLASM (DISORDER)
C0348213|T047|187449003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE RESULTING IN MALIGNANT NEOPLASMS|[X]HIV DISEASE RESULTING IN UNSPECIFIED MALIGNANT NEOPLASM (DISORDER)
C0348213|T047|187449003|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN UNSPECIFIED MALIGNANT NEOPLASM|[X]HIV DISEASE RESULTING IN UNSPECIFIED MALIGNANT NEOPLASM (DISORDER)
C0348213|T047|187449003|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN UNSPECIFIED MALIGNANT NEOPLASM |[X]HIV DISEASE RESULTING IN UNSPECIFIED MALIGNANT NEOPLASM (DISORDER)
C0348213|T047|187449003|SNOMEDCT_US|HIV DISEASE; NEOPLASM, MALIGNANT|[X]HIV DISEASE RESULTING IN UNSPECIFIED MALIGNANT NEOPLASM (DISORDER)
C0494097|T047||SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE RESULTING IN OTHER CONDITIONS
C0494096|T047||SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE RESULTING IN OTHER SPECIFIED DISEASES
C0152983|T047||SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION CAUSING OTHER SPECIFIED CONDITIONS
C0152987|T047||SNOMEDCT_US|OTHER HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C1142553|T047||SNOMEDCT_US|PRIMARY HIV INFECTION
C0152979|T047||SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH SPECIFIED CONDITIONS
C0152988|T047||SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION CAUSING SPECIFIED ACUTE INFECTIONS
C0343752|T047|111880001|SNOMEDCT_US|ACUTE HIV INFECTION|ACUTE HIV INFECTION (DISORDER)
C0343752|T047|111880001|SNOMEDCT_US|ACUTE HIV INFECTION SYNDROME|ACUTE HIV INFECTION (DISORDER)
C0343752|T047|111880001|SNOMEDCT_US|ACUTE HUMAN IMMUNODEFICIENCY VIRUS INFECTION |ACUTE HIV INFECTION (DISORDER)
C0343752|T047|111880001|SNOMEDCT_US|ACUTE HIV INFECTION |ACUTE HIV INFECTION (DISORDER)
C0343752|T047|111880001|SNOMEDCT_US|HIV INFECTION ACUTE|ACUTE HIV INFECTION (DISORDER)
C0343752|T047|111880001|SNOMEDCT_US|ACUTE HIV INFECTION |ACUTE HIV INFECTION (DISORDER)
C0343752|T047|111880001|SNOMEDCT_US|ACUTE INFECTION WITH HIV|ACUTE HIV INFECTION (DISORDER)
C0343752|T047|111880001|SNOMEDCT_US|HIV SEROCONVERSION ILLNESS|ACUTE HIV INFECTION (DISORDER)
C0343752|T047|111880001|SNOMEDCT_US|ACUTE HUMAN IMMUNODEFICIENCY VIRUS INFECTION|ACUTE HIV INFECTION (DISORDER)
C0343752|T047|111880001|SNOMEDCT_US|ACUTE HUMAN IMMUNODEFICIENCY VIRUS SEROCONVERSION ILLNESS|ACUTE HIV INFECTION (DISORDER)
C0343751|T047|91947003|SNOMEDCT_US|ASYMPTOMATIC HIV INFECTION|ASYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0343751|T047|91947003|SNOMEDCT_US|HIV INFECTION ASYMPTOMATIC|ASYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0343751|T047|91947003|SNOMEDCT_US|ASYMPTOMATIC HIV INFECTION |ASYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0343751|T047|91947003|SNOMEDCT_US|ASYMPTOMATIC INFECTION WITH HIV|ASYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0343751|T047|91947003|SNOMEDCT_US|ASYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION|ASYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0343751|T047|91947003|SNOMEDCT_US|ASYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION |ASYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0864665|T047||SNOMEDCT_US|HIV INFECTION, SYMPTOMATIC
C0864665|T047||SNOMEDCT_US|SYMPTOMATIC HIV INFECTION
C0864665|T047||SNOMEDCT_US|HIV INFECTION SYMPTOMATIC
C0864665|T047||SNOMEDCT_US|SYMPTOMATIC HIV INFECTION 
C0001857|T047|266201009|SNOMEDCT_US|AIDS RELATED COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|AIDS-RELATED COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|COMPLEX, AIDS-RELATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|AIDS-LIKE SYNDROME |ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|AIDS RELAT COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|AIDS-RELATED COMPLEX [ARC]|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|AIDS-RELATED COMPLEX [DISEASE/FINDING]|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS)-LIKE SYNDROME |ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC])|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) |ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|AIDS-RELATED COMPLEX (ARC)|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME-LIKE SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME-LIKE SYNDROME |ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME-RELATED COMPLEX, UNSPECIFIED|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|AIDS-LIKE SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS)-LIKE SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED COMPLEX |ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME-LIKE SYNDROME |ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ARC - ACQUIRED IMMUNODEFICIENCY SYNDROME-RELATED COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0001857|T047|266201009|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME (& [ARC]) (DISORDER)
C0019699|T047|402916007|SNOMEDCT_US|AIDS SEROCONVERSIONS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|AIDS SEROPOSITIVITIES|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV SEROCONVERSIONS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV SEROPOSITIVITIES|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV SEROPOSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|SEROCONVERSION, AIDS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|SEROCONVERSION, HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|SEROCONVERSIONS, AIDS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|SEROCONVERSIONS, HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|SEROPOSITIVITIES, AIDS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|SEROPOSITIVITIES, HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|SEROPOSITIVITY, AIDS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|SEROPOSITIVITY, HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|ANTI HIV POSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|ANTI-HIV POSITIVITIES|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|ANTIBODY POSITIVITIES, HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|ANTIBODY POSITIVITY, HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV ANTIBODY POSITIVITIES|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|POSITIVITIES, ANTI-HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|POSITIVITIES, HIV ANTIBODY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|POSITIVITY, ANTI-HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|POSITIVITY, HIV ANTIBODY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV POSITIVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV POSITIVE |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV SEROPOSITIVITY |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) POSITIVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV ANTIBODY POS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HTLV III SEROPOS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|ANTIHIV POSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HTLV WIII SEROCONVERSION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV SEROPOS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|AIDS SEROPOS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HTLV WIII SEROPOSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|ANTI HIV POS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|SEROPOSITIVE (AIDS TEST)|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV TEST POSITIVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV POSITVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV TEST POSITVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV POSITIVE NOS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|AIDS SEROCONVERSION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HTLV-III SEROCONVERSION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV ANTIBODY POSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV SEROPOSITIVITY [DISEASE/FINDING]|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|ANTI-HIV POSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|AIDS SEROPOSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HTLV-III SEROPOSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV SEROCONVERSION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|ANTIBODY POSITIVE AIDS TEST|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|ANTIGEN POSITIVE AIDS TEST|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS POSITIVE |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) POSITIVE |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS POSITIVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV SEROPOSITIVITY |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS SEROPOSITIVITY |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS SEROPOSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|POSITIVE TEST FOR HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HTLV III TEST POSITIVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV SEROPOSITIVE NOS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV+|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV-TEST; POSITIVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV; POSITIVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV; TEST, POSITIVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|POSITIVE; HIV-TEST|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|POSITIVE; HIV|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|TEST; HIV, POSITIVE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0019699|T047|402916007|SNOMEDCT_US|HIV POSITIVITY|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROPOSITIVITY
C0001849|T047|192178000|SNOMEDCT_US|AIDS DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|COMPLEX, AIDS DEMENTIA|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA, HIV|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA IN HUMAN IMMUNODEFICIENCY VIRUS [HIV] DISEASE|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|ADC - ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS - ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED DEMENTIA|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA ASSOCIATED WITH AIDS|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA COMPLEX AIDS RELAT|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV ASSOC COGNITIVE MOTOR COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA COMPLEX ACQUIRED IMMUNE DEFIC SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|ACQUIRED IMMUNE DEFIC SYNDROME DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS RELAT DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) DEMENTIA|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) DEMENTIA |ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS DEMENTIA|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA COMPLEX, AIDS|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS RELATED DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|COMPLEX, AIDS-RELATED DEMENTIA|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA COMPLEX, AIDS RELATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIAS, HIV|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV DEMENTIAS|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA COMPLEX, AIDS-RELATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|ACQUIRED-IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS-RELATED DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA COMPLEX, ACQUIRED IMMUNE DEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS DEMENTIA COMPLEX [DISEASE/FINDING]|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV DEMENTIA|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV-ASSOCIATED COGNITIVE MOTOR COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV ASSOCIATED COGNITIVE MOTOR COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV ASSOCIATED COGNITIVE AND MOTOR COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS WITH DEMENTIA |ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX |ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS WITH DEMENTIA|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA ASSOCIATED WITH AIDS |ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME |ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV-RELATED DEMENTIA|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS-DEMENTIA COMPLEX|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS-RELATED DEMENTIA|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA DUE TO HIV DISEASE|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV DISEASE; DEMENTIA (ETIOLOGY)|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV DISEASE; DEMENTIA (MANIFESTATION)|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV DISEASE; RESULTING IN, DEMENTIA (ETIOLOGY)|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|HIV DISEASE; RESULTING IN, DEMENTIA (MANIFESTATION)|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA; HUMAN IMMUNODEFICIENCY VIRUS DISEASE (ETIOLOGY)|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|DEMENTIA; HUMAN IMMUNODEFICIENCY VIRUS DISEASE (MANIFESTATION)|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0001849|T047|192178000|SNOMEDCT_US|AIDS WITH DEMENTIA, NOS|ACQUIRED IMMUNE DEFICIENCY SYNDROME DEMENTIA COMPLEX (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS ASSOCIATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS-ASSOCIATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV ASSOCIATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV RELATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES, AIDS|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY, AIDS|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS ASSOCIATED NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV ASSOCIATED NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV RELATED NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES, AIDS ASSOCIATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES, HIV ASSOCIATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES, HIV RELATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY, AIDS ASSOCIATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY, HIV ASSOCIATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY, HIV RELATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV-ASSOCIATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS-RELATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV RELAT NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV RELAT NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY HIV RELAT|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY AIDS ASSOC|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY HIV ASSOC|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS ASSOC NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIVAN|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HUMAN IMMUNODEFIC VIRUS ASSOC NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES AIDS ASSOC|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES HIV RELAT|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS ASSOC NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV ASSOC NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES HIV ASSOC|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV-ASSOCIATED NEPHROPATHY |ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS-ASSOCIATED NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV-RELATED NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES, AIDS-ASSOCIATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV-ASSOCIATED NEPHROPATHIES|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES, HIV-ASSOCIATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV-RELATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHIES, HIV-RELATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY, AIDS-ASSOCIATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY, HIV-ASSOCIATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|NEPHROPATHY, HIV-RELATED|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS-ASSOCIATED NEPHROPATHY [DISEASE/FINDING]|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-ASSOCIATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS ASSOCIATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HIV NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-RELATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|AIDS - ACQUIRED IMMUNE DEFICIENCY SYND-RELATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0078911|T047|236406007|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY |ACQUIRED IMMUNE DEFICIENCY SYNDROME-RELATED NEPHROPATHY (DISORDER)
C0162526|T047||SNOMEDCT_US|AIDS-RELATED OPPORTUNISTIC INFECTIONS
C0162526|T047||SNOMEDCT_US|AIDS RELATED OPPORTUNISTIC INFECTIONS
C0162526|T047||SNOMEDCT_US|AIDS-RELATED OPPORTUNISTIC INFECTION
C0162526|T047||SNOMEDCT_US|OPPORTUNISTIC INFECTION, AIDS-RELATED
C0162526|T047||SNOMEDCT_US|OPPORTUNISTIC INFECTIONS, AIDS RELATED
C0162526|T047||SNOMEDCT_US|HIV RELATED OPPORTUNISTIC INFECTIONS
C0162526|T047||SNOMEDCT_US|HIV-RELATED OPPORTUNISTIC INFECTION
C0162526|T047||SNOMEDCT_US|INFECTION, HIV-RELATED OPPORTUNISTIC
C0162526|T047||SNOMEDCT_US|INFECTIONS, HIV-RELATED OPPORTUNISTIC
C0162526|T047||SNOMEDCT_US|OPPORTUNISTIC INFECTION, HIV-RELATED
C0162526|T047||SNOMEDCT_US|OPPORTUNISTIC INFECTIONS, HIV RELATED
C0162526|T047||SNOMEDCT_US|HIV RELAT OPPORTUNISTIC INFECT
C0162526|T047||SNOMEDCT_US|OPPORTUNISTIC INFECT AIDS RELAT
C0162526|T047||SNOMEDCT_US|AIDS RELAT OPPORTUNISTIC INFECT
C0162526|T047||SNOMEDCT_US|OPPORTUNISTIC INFECT HIV RELAT
C0162526|T047||SNOMEDCT_US|HIV-RELATED OPPORTUNISTIC INFECTIONS
C0162526|T047||SNOMEDCT_US|OPPORTUNISTIC INFECTIONS, HIV-RELATED
C0162526|T047||SNOMEDCT_US|AIDS-RELATED OPPORTUNISTIC INFECTIONS [DISEASE/FINDING]
C0162526|T047||SNOMEDCT_US|OPPORTUNISTIC INFECTIONS, AIDS-RELATED
C0162526|T047||SNOMEDCT_US|OPPORTUNISTIC INFECTIONS IN AIDS
C0162526|T047||SNOMEDCT_US|AIDS ASSOCIATED OPPORTUNISTIC INFECTION
C0162526|T047||SNOMEDCT_US|AIDS, OPPORTUNISTIC INFECTION
C0282616|T047|235726002|SNOMEDCT_US|AIDS ASSOCIATED ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|AIDS ENTEROPATHIES|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|AIDS-ASSOCIATED ENTEROPATHIES|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHIES, AIDS|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHIES, AIDS-ASSOCIATED|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHIES, HIV|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHIES, HIV-ASSOCIATED|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHY, AIDS|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHY, AIDS ASSOCIATED|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHY, HIV ASSOCIATED|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV ASSOCIATED ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV ENTEROPATHIES|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV-ASSOCIATED ENTEROPATHIES|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV ASSOC ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHY HIV ASSOC|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHY AIDS ASSOC|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|AIDS ASSOC ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|INFECTIOUS DIARRHEA OF HIV PATIENT|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|INFECTIOUS DIARRHEA OF HIV PATIENT |HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|AIDS ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|AIDS-ASSOCIATED ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHY, HIV|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHY, HIV-ASSOCIATED|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|IDIOPATHIC AIDS ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHY, AIDS-ASSOCIATED|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV ENTEROPATHY [DISEASE/FINDING]|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV-ASSOCIATED ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV ENTEROPATHY |HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|AIDS ENTEROPATHIES, IDIOPATHIC|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|AIDS ENTEROPATHY, IDIOPATHIC|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHIES, IDIOPATHIC AIDS|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|ENTEROPATHY, IDIOPATHIC AIDS|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|IDIOPATHIC AIDS ENTEROPATHIES|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS DIARRHEA|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS DIARRHOEA|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DIARRHEA|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DIARRHOEA|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS NON-PATHOGENIC DIARRHEA|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS NON-PATHOGENIC DIARRHOEA|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0282616|T047|235726002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY |HUMAN IMMUNODEFICIENCY VIRUS ENTEROPATHY (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HIV WASTING SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HIV DISEASE RESULTING IN WASTING SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|WASTING SYNDROME, AIDS|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|SLIM DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|CACHEXIA ASSOCIATED WITH AIDS|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HIV WASTING DIS|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|SLIM DIS|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|WASTING DIS HIV|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|AIDS WASTING SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HIV WASTING SYNDROME [DISEASE/FINDING]|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HIV WASTING DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|WASTING DISEASE, HIV|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|WASTING SYNDROME, HIV|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME |HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|AIDS WITH CACHEXIA|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|AIDS WITH CACHEXIA |HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|CACHEXIA ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|CACHEXIA ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME |HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|CACHEXIA ASSOCIATED WITH AIDS |HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HIV DISEASE; FAILURE TO THRIVE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HIV DISEASE; RESULTING IN, FAILURE TO THRIVE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|HIV DISEASE; RESULTING IN, WASTING SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|DISEASE (OR DISORDER); SLIM DISEASE (HIV)|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0343755|T047|186727001|SNOMEDCT_US|DISEASE; SLIM|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WASTING SYNDROME (DISORDER)
C0752330|T047||SNOMEDCT_US|AIDS ARTERITIS CNS
C0752330|T047||SNOMEDCT_US|CNS AIDS ARTERITIS
C0752330|T047||SNOMEDCT_US|AIDS ARTERITIS, CENTRAL NERVOUS SYSTEM
C0752330|T047||SNOMEDCT_US|CENTRAL NERVOUS SYSTEM AIDS ARTERITIS
C0752330|T047||SNOMEDCT_US|AIDS ARTERITIS, CENTRAL NERVOUS SYSTEM [DISEASE/FINDING]
C1136321|T047||SNOMEDCT_US|HIV ASSOC LIPODYSTROPHY SYNDROME
C1136321|T047||SNOMEDCT_US|HIV ASSOC LIPODYSTROPHY
C1136321|T047||SNOMEDCT_US|HIV LIPODYSTROPHY SYNDROME
C1136321|T047||SNOMEDCT_US|HIV-ASSOCIATED LIPODYSTROPHY SYNDROME
C1136321|T047||SNOMEDCT_US|HIV-ASSOCIATED LIPODYSTROPHY
C1136321|T047||SNOMEDCT_US|HIV-ASSOCIATED LIPODYSTROPHY SYNDROME [DISEASE/FINDING]
C1136321|T047||SNOMEDCT_US|LIPODYSTROPHY SYNDROME, HIV
C1136321|T047||SNOMEDCT_US|HIV ASSOCIATED LIPODYSTROPHY
C1136321|T047||SNOMEDCT_US|HIV ASSOCIATED LIPODYSTROPHY SYNDROME
C1136321|T047||SNOMEDCT_US|LIPODYSTROPHY SYNDROME, HIV-ASSOCIATED
C1136321|T047||SNOMEDCT_US|LIPODYSTROPHY, HIV-ASSOCIATED
C0520783|T047|52079000|SNOMEDCT_US|CONGENITAL HIV INFECTION|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0520783|T047|52079000|SNOMEDCT_US|HIV INFECTION CONGENITAL|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0520783|T047|52079000|SNOMEDCT_US|CONGENITAL HIV INFECTION |CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0520783|T047|52079000|SNOMEDCT_US|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS INFECTION|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0520783|T047|52079000|SNOMEDCT_US|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS INFECTION |CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C2319244|T047||SNOMEDCT_US|HIV INFECTION CDC CLASSIFICATION 
C2319244|T047||SNOMEDCT_US|HIV INFECTION CDC CLASSIFICATION
C2046425|T047||SNOMEDCT_US|HIV INFECTION, STAGE 0 
C2046425|T047||SNOMEDCT_US|HIV INFECTION, STAGE 0
C2046426|T047||SNOMEDCT_US|HIV INFECTION, STAGE 1 
C2046426|T047||SNOMEDCT_US|HIV INFECTION, STAGE 1
C2046427|T047||SNOMEDCT_US|HIV INFECTION, STAGE 2 (PGL) 
C2046427|T047||SNOMEDCT_US|PGL (PERSISTENT GENERALIZED LYMPHADENOPATHY) STAGE II OF HIV INFECTION
C2046427|T047||SNOMEDCT_US|HIV INFECTION, STAGE 2 (PGL)
C2240389|T047||SNOMEDCT_US|HIV INFECTION, STAGE 3 (PGL) 
C2240389|T047||SNOMEDCT_US|HIV INFECTION, STAGE 3 (PGL)
C2240389|T047||SNOMEDCT_US|PGL (PERSISTENT GENERALIZED LYMPHADENOPATHY) STAGE III OF HIV INFECTION
C2046428|T047||SNOMEDCT_US|HIV INFECTION, STAGE 4
C2046428|T047||SNOMEDCT_US|HIV INFECTION, STAGE 4 
C2046429|T047||SNOMEDCT_US|ARC (AIDS-RELATED COMPLEX) STAGE V OF HIV INFECTION
C2046429|T047||SNOMEDCT_US|HIV INFECTION, STAGE 5 (ARC)
C2046429|T047||SNOMEDCT_US|HIV INFECTION, STAGE 5 (ARC) 
C0276554|T047|421977001|SNOMEDCT_US|AIDS WITH LYMPHADENOPATHY|LYMPHADENOPATHY ASSOCIATED WITH AIDS
C0276554|T047|421977001|SNOMEDCT_US|AIDS WITH LYMPHADENOPATHY |LYMPHADENOPATHY ASSOCIATED WITH AIDS
C0276554|T047|421977001|SNOMEDCT_US|LYMPHADENOPATHY ASSOCIATED WITH AIDS |LYMPHADENOPATHY ASSOCIATED WITH AIDS
C0276554|T047|421977001|SNOMEDCT_US|LYMPHADENOPATHY ASSOCIATED WITH AIDS|LYMPHADENOPATHY ASSOCIATED WITH AIDS
C0276554|T047|421977001|SNOMEDCT_US|LYMPHADENOPATHY ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME |LYMPHADENOPATHY ASSOCIATED WITH AIDS
C0276554|T047|421977001|SNOMEDCT_US|LYMPHADENOPATHY ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME|LYMPHADENOPATHY ASSOCIATED WITH AIDS
C1834751|T047||SNOMEDCT_US|CORONARY ARTERY DISEASE, DEVELOPMENT OF, IN HIV
C1304455|T047|402901009|SNOMEDCT_US|ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HUMAN IMMUNODEFICIENCY VIRUS DISEASE |ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HIV DISEASE (DISORDER)
C1304455|T047|402901009|SNOMEDCT_US|ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HIV DISEASE |ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HIV DISEASE (DISORDER)
C1304455|T047|402901009|SNOMEDCT_US|ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HUMAN IMMUNODEFICIENCY VIRUS DISEASE|ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HIV DISEASE (DISORDER)
C1304455|T047|402901009|SNOMEDCT_US|ORAL HAIRY LEUCOPLAKIA ASSOCIATED WITH HUMAN IMMUNODEFICIENCY VIRUS DISEASE|ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HIV DISEASE (DISORDER)
C1304455|T047|402901009|SNOMEDCT_US|ORAL HAIRY LEUCOPLAKIA ASSOCIATED WITH HIV DISEASE|ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HIV DISEASE (DISORDER)
C1304455|T047|402901009|SNOMEDCT_US|ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HIV DISEASE|ORAL HAIRY LEUKOPLAKIA ASSOCIATED WITH HIV DISEASE (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|AIDS WITH KAPOSI'S SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|HIV DISEASE RESULTING IN KAPOSI'S SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|AIDS-RELATED KAPOSI SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|AIDS-RELATED KAPOSI'S SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI'S SARCOMA AIDS RELATED|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI SARCOMA ASSOCIATED WITH AIDS|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|HIV DISEASE RESULTING IN KAPOSI'S SARCOMA |KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|AIDS WITH KAPOSI'S SARCOMA |KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS |KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI'S SARCOMA ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME |KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI'S SARCOMA ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|MALIGNANT NEOPLASM SARCOMA KAPOSI'S ASSOCIATED WITH AIDS|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS |KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI'S SARCOMA EPIDEMIC TYPE|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|EPIDEMIC KAPOSI'S SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|AIDS RELATED KAPOSI'S SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|AIDS RELATED MULTIPLE HEMORRHAGIC SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|AIDS-ASSOCIATED KAPOSI'S SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI'S SARCOMA, AIDS RELATED|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI'S SARCOMA, EPIDEMIC|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|ACQUIRED IMMUNE DEFICIENCY SYNDROME RELATED KAPOSI'S SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|MULTIPLE HEMORRHAGIC SARCOMA, AIDS RELATED|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|SARCOMA, KAPOSI'S, AIDS RELATED|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|SARCOMA, MULTIPLE HEMORRHAGIC, AIDS RELATED|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|HIV DISEASE; KAPOSI'S SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|HIV DISEASE; SARCOMA, KAPOSI|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|KAPOSI; SARCOMA, RESULTING FROM HIV DISEASE|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|SARCOMA; KAPOSI, RESULTING FROM HIV DISEASE|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|AUTOIMMUNE DEFICIENCY SYNDROME-RELATED KAPOSI SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0276535|T047|420524008|SNOMEDCT_US|AIDS, KAPOSI'S SARCOMA|KAPOSI'S SARCOMA ASSOCIATED WITH AIDS (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA |HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|HIV DISEASE; PNEUMOCYSTOSIS|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|HIV DISEASE; RESULTING IN, PNEUMOCYSTIS CARINII PNEUMONIA|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|HIV DISEASE; RESULTING IN, INFECTION, PNEUMOCYSTIS CARINII (PNEUMONIA)|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|PNEUMOCYSTIS CARINII; INFECTION, RESULTING FROM HIV DISEASE|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|INFECTION; PNEUMOCYSTIS CARINII, RESULTING FROM HIV DISEASE|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|PNEUMOCYSTOSIS; PNEUMONIA, RESULTING FROM HIV DISEASE|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|PNEUMOCYSTOSIS; RESULTING FROM HIV DISEASE|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0348804|T047|186720004|SNOMEDCT_US|PNEUMONIA; PNEUMOCYSTOSIS, RESULTING FROM HIV DISEASE|HIV DISEASE RESULTING IN PNEUMOCYSTIS CARINII PNEUMONIA (DISORDER)
C0452192|T047|186724008|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER TYPES OF NON-HODGKIN'S LYMPHOMA|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN OTHER TYPES OF NON-HODGKIN'S LYMPHOMA
C0452192|T047|186724008|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER TYPES OF NON-HODGKIN'S LYMPHOMA |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN OTHER TYPES OF NON-HODGKIN'S LYMPHOMA
C0452192|T047|186724008|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN OTHER TYPES OF NON-HODGKIN'S LYMPHOMA |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN OTHER TYPES OF NON-HODGKIN'S LYMPHOMA
C0452192|T047|186724008|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN OTHER TYPES OF NON-HODGKIN'S LYMPHOMA|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN OTHER TYPES OF NON-HODGKIN'S LYMPHOMA
C0348983|T047|186716003|SNOMEDCT_US|HUMAN IMMUNODEF VIRUS RESULTING IN OTHER DISEASE |HUMAN IMMUNODEF VIRUS RESULTING IN OTHER DISEASE (DISORDER)
C0348983|T047|186716003|SNOMEDCT_US|HUMAN IMMUNODEF VIRUS RESULTING IN OTHER DISEASE|HUMAN IMMUNODEF VIRUS RESULTING IN OTHER DISEASE (DISORDER)
C0343749|T047|186714000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS WITH OTHER CLINICAL FINDINGS|HUMAN IMMUNODEFICIENCY VIRUS WITH OTHER CLINICAL FINDINGS (DISORDER)
C0343749|T047|186714000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS WITH OTHER CLINICAL FINDINGS |HUMAN IMMUNODEFICIENCY VIRUS WITH OTHER CLINICAL FINDINGS (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|HIV NEUROPATHY|HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY |HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY|HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY|HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|NEUROPATHY DUE TO HUMAN IMMUNODEFICIENCY VIRUS|HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|NEUROPATHY DUE TO HUMAN IMMUNODEFICIENCY VIRUS |HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|NEUROPATHY DUE TO HUMAN IMMUNODEFICIENCY VIRUS |HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|NEUROPATHY CAUSED BY HUMAN IMMUNODEFICIENCY VIRUS |HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|NEUROPATHY CAUSED BY HUMAN IMMUNODEFICIENCY VIRUS|HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|NEUROPATHY CAUSED BY HIV - HUMAN IMMUNODEFICIENCY VIRUS|HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C0343757|T047|240612001|SNOMEDCT_US|NEUROPATHY DUE TO HIV - HUMAN IMMUNODEFICIENCY VIRUS|HUMAN IMMUNODEFICIENCY VIRUS NEUROPATHY (DISORDER)
C3648901|T047||SNOMEDCT_US|HIV INFECTION COMPLICATING PREGNANCY, CHILDBIRTH, AND PUERPERIUM
C3648901|T047||SNOMEDCT_US|HIV INFECTION COMPLICATING PREGNANCY, CHILDBIRTH, AND PUERPERIUM 
C3648903|T047||SNOMEDCT_US|HIV INFECTION COMPLICATING CHILDBIRTH
C3648903|T047||SNOMEDCT_US|HIV INFECTION COMPLICATING CHILDBIRTH 
C3648900|T047||SNOMEDCT_US|HIV INFECTION COMPLICATING PUERPERIUM
C3648900|T047||SNOMEDCT_US|HIV INFECTION COMPLICATING PUERPERIUM 
C3661937|T047|81000119104|SNOMEDCT_US|SYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION |SYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C3661937|T047|81000119104|SNOMEDCT_US|SYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION|SYMPTOMATIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0343748|T047|186709004|SNOMEDCT_US|HIV INFECTION WITH SECONDARY CANCERS|HUMAN IMMUNODEFICIENCY VIRUS WITH SECONDARY CANCERS (DISORDER)
C0343748|T047|186709004|SNOMEDCT_US|HIV INFECTION WITH SECONDARY CANCERS |HUMAN IMMUNODEFICIENCY VIRUS WITH SECONDARY CANCERS (DISORDER)
C0343748|T047|186709004|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS WITH SECONDARY CANCERS|HUMAN IMMUNODEFICIENCY VIRUS WITH SECONDARY CANCERS (DISORDER)
C0343748|T047|186709004|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS WITH SECONDARY CANCERS |HUMAN IMMUNODEFICIENCY VIRUS WITH SECONDARY CANCERS (DISORDER)
C0343754|T047|186706006|SNOMEDCT_US|HIV INFECTION CONSTITUTIONAL DISEASE |HUMAN IMMUNODEFICIENCY VIRUS INFECTION CONSTITUTIONAL DISEASE (DISORDER)
C0343754|T047|186706006|SNOMEDCT_US|HIV INFECTION CONSTITUTIONAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION CONSTITUTIONAL DISEASE (DISORDER)
C0343754|T047|186706006|SNOMEDCT_US|HIV INFECTION WITH CONSTITUTIONAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION CONSTITUTIONAL DISEASE (DISORDER)
C0343754|T047|186706006|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS INFECTION CONSTITUTIONAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION CONSTITUTIONAL DISEASE (DISORDER)
C0343754|T047|186706006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION CONSTITUTIONAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION CONSTITUTIONAL DISEASE (DISORDER)
C0343754|T047|186706006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION CONSTITUTIONAL DISEASE |HUMAN IMMUNODEFICIENCY VIRUS INFECTION CONSTITUTIONAL DISEASE (DISORDER)
C1274337|T047|402915006|SNOMEDCT_US|HIV SEROCONVERSION EXANTHEM |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROCONVERSION EXANTHEM
C1274337|T047|402915006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROCONVERSION EXANTHEM |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROCONVERSION EXANTHEM
C1274337|T047|402915006|SNOMEDCT_US|HIV SEROCONVERSION EXANTHEM|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROCONVERSION EXANTHEM
C1274337|T047|402915006|SNOMEDCT_US|HIV SEROCONVERSION EXANTHEM |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROCONVERSION EXANTHEM
C1274337|T047|402915006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS SEROCONVERSION EXANTHEM|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROCONVERSION EXANTHEM
C1274337|T047|402915006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROCONVERSION EXANTHEM|HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROCONVERSION EXANTHEM
C1274337|T047|402915006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS SEROCONVERSION EXANTHEM |HUMAN IMMUNODEFICIENCY VIRUS (HIV) SEROCONVERSION EXANTHEM
C0276600|T047|315019000|SNOMEDCT_US|HIV INFECTION WITH ASEPTIC MENINGITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0276600|T047|315019000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0276600|T047|315019000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH ASEPTIC MENINGITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0276600|T047|315019000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH ASEPTIC MENINGITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0276600|T047|315019000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0276600|T047|315019000|SNOMEDCT_US|AIDS VIRUS WITH ASEPTIC MENINGITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0276600|T047|315019000|SNOMEDCT_US|AIDS VIRUS WITH ASEPTIC MENINGITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0276600|T047|315019000|SNOMEDCT_US|HIV INFECTION WITH ASEPTIC MENINGITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0276600|T047|315019000|SNOMEDCT_US|HIV INFECTION WITH ASEPTIC MENINGITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0276600|T047|315019000|SNOMEDCT_US|HIV INFECTION WITH ASEPTIC MENINGITIS  [AMBIGUOUS]|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ASEPTIC MENINGITIS
C0206019|T047|397763006|SNOMEDCT_US|HIV DISEASE RESULTING IN ENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|ENCEPH HIV|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|ENCEPH AIDS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HIV ENCEPH|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|AIDS ENCEPH|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HIV ENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) ENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) ENCEPHALOPATHY |HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|AIDS ENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|AIDS ENCEPHALOPATHIES|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|ENCEPHALOPATHIES, AIDS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|ENCEPHALOPATHIES, HIV|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HIV ENCEPHALOPATHIES|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|AIDS WITH ENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|AIDS WITH ENCEPHALOPATHY |HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HIV ENCEPHALOPATHY |HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS ENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS ENCEPHALOPATHY |HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY |HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|ENCEPHALOPATHY, HIV|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|ENCEPHALOPATHY, AIDS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HIV DISEASE; ENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|HIV DISEASE; RESULTING IN, ENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0206019|T047|397763006|SNOMEDCT_US|ENCEPHALOPATHY; RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALOPATHY (DISORDER)
C0399449|T047|235009000|SNOMEDCT_US|HIV ASSOCIATED PERIDONTITIS|HUMAN IMMUNODEFICIENCY VIRUS-ASSOCIATED PERIODONTITIS (DISORDER)
C0399449|T047|235009000|SNOMEDCT_US|HIV ASSOCIATED PERIDONTITIS |HUMAN IMMUNODEFICIENCY VIRUS-ASSOCIATED PERIODONTITIS (DISORDER)
C0399449|T047|235009000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-ASSOCIATED PERIODONTITIS|HUMAN IMMUNODEFICIENCY VIRUS-ASSOCIATED PERIODONTITIS (DISORDER)
C0399449|T047|235009000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-ASSOCIATED PERIODONTITIS |HUMAN IMMUNODEFICIENCY VIRUS-ASSOCIATED PERIODONTITIS (DISORDER)
C0348990|T047|186719005|SNOMEDCT_US|HIV DISEASE RESULTING IN CANDIDIASIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HIV DISEASE RESULTING IN CANDIDIASIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HIV INFECTION RESULTING IN CANDIDIASIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HIV INFECTION RESULTING IN CANDIDIASIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN CANDIDIASIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN CANDIDIASIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HIV DISEASE; CANDIDIASIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HIV DISEASE; RESULTING IN, CANDIDIASIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|HIV DISEASE; RESULTING IN, INFECTION, CANDIDA|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|CANDIDA; INFECTION, RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|CANDIDIASIS; RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0348990|T047|186719005|SNOMEDCT_US|INFECTION; CANDIDA, RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CANDIDIASIS
C0343747|T047|186707002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH NEUROLOGICAL DISEASE |HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH NEUROLOGICAL DISEASE (DISORDER)
C0343747|T047|186707002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS WITH NEUROLOGICAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH NEUROLOGICAL DISEASE (DISORDER)
C0343747|T047|186707002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH NEUROLOGICAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH NEUROLOGICAL DISEASE (DISORDER)
C0343747|T047|186707002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS WITH NEUROLOGICAL DISEASE |HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH NEUROLOGICAL DISEASE (DISORDER)
C0343747|T047|186707002|SNOMEDCT_US|HIV INFECTION WITH NEUROLOGICAL DISEASE |HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH NEUROLOGICAL DISEASE (DISORDER)
C0343747|T047|186707002|SNOMEDCT_US|HIV INFECTION WITH NEUROLOGICAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH NEUROLOGICAL DISEASE (DISORDER)
C0348969|T047|186717007|SNOMEDCT_US|HIV DISEASE RESULTING IN MYCOBACTERIAL INFECTION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HIV DISEASE RESULTING IN MYCOBACTERIAL INFECTION |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HIV INFECTION RESULTING IN MYCOBACTERIAL INFECTION |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HIV INFECTION RESULTING IN MYCOBACTERIAL INFECTION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN MYCOBACTERIAL INFECTION |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN MYCOBACTERIAL INFECTION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HIV DISEASE; MYCOBACTERIUM|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HIV DISEASE; RESULTING IN, INFECTION, MYCOBACTERIAL|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|HIV DISEASE; RESULTING IN, MYCOBACTERIAL INFECTION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|MYCOBACTERIUM; INFECTION, RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|MYCOBACTERIUM; RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|INFECTION; MYCOBACTERIUM, MYCOBACTERIAL, RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348969|T047|186717007|SNOMEDCT_US|INFECTION; TUBERCULOUS, RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MYCOBACTERIAL INFECTION
C0348982|T047|186718002|SNOMEDCT_US|HIV DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HIV DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HIV INFECTION RESULTING IN CYTOMEGALOVIRAL INFECTION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HIV INFECTION RESULTING IN CYTOMEGALOVIRAL INFECTION |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HIV DISEASE; CYTOMEGALOVIRAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HIV DISEASE; RESULTING IN, CYTOMEGALOVIRAL DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|HIV DISEASE; RESULTING IN, INFECTION, CYTOMEGALOVIRAL|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348982|T047|186718002|SNOMEDCT_US|CYTOMEGALOVIRAL DISEASE; RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN CYTOMEGALOVIRAL DISEASE
C0348821|T047|186726005|SNOMEDCT_US|HIV DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348821|T047|186726005|SNOMEDCT_US|HIV DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348821|T047|186726005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348821|T047|186726005|SNOMEDCT_US|HIV INFECTION RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348821|T047|186726005|SNOMEDCT_US|HIV INFECTION RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348821|T047|186726005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348821|T047|186726005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348821|T047|186726005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348821|T047|186726005|SNOMEDCT_US|HIV DISEASE; RESULTING IN, LYMPHOID INTERSTITIAL PNEUMONITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348821|T047|186726005|SNOMEDCT_US|HIV DISEASE; RESULTING IN, PNEUMONITIS, INTERSTITIAL, LYMPHATIC|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN LYMPHOID INTERSTITIAL PNEUMONITIS
C0348207|T047|186721000|SNOMEDCT_US|HIV DISEASE RESULTING IN MULTIPLE INFECTIONS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0348207|T047|186721000|SNOMEDCT_US|HIV DISEASE RESULTING IN MULTIPLE INFECTIONS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0348207|T047|186721000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0348207|T047|186721000|SNOMEDCT_US|HIV INFECTION RESULTING IN MULTIPLE INFECTIONS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0348207|T047|186721000|SNOMEDCT_US|HIV INFECTION RESULTING IN MULTIPLE INFECTIONS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0348207|T047|186721000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0348207|T047|186721000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN MULTIPLE INFECTIONS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0348207|T047|186721000|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN MULTIPLE INFECTIONS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0348207|T047|186721000|SNOMEDCT_US|HIV DISEASE; RESULTING IN MULTIPLE INFECTIONS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0348207|T047|186721000|SNOMEDCT_US|HIV DISEASE; RESULTING IN, INFECTION, MULTIPLE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE INFECTIONS
C0349036|T047|186725009|SNOMEDCT_US|HIV DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS
C0349036|T047|186725009|SNOMEDCT_US|HIV DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS
C0349036|T047|186725009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS
C0349036|T047|186725009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS
C0349036|T047|186725009|SNOMEDCT_US|HIV INFECTION RESULTING IN MULTIPLE MALIGNANT NEOPLASMS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS
C0349036|T047|186725009|SNOMEDCT_US|HIV INFECTION RESULTING IN MULTIPLE MALIGNANT NEOPLASMS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS
C0349036|T047|186725009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS
C0349036|T047|186725009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS
C0349036|T047|186725009|SNOMEDCT_US|HIV DISEASE; RESULTING IN, NEOPLASM, MALIGNANT, MULTIPLE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN MULTIPLE MALIGNANT NEOPLASMS
C0410223|T047|240103002|SNOMEDCT_US|HIV-ASSOCIATED MYOPATHY|HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY (DISORDER)
C0410223|T047|240103002|SNOMEDCT_US|HIV-ASSOCIATED MYOPATHY |HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY (DISORDER)
C0410223|T047|240103002|SNOMEDCT_US|HIV ASSOCIATED MYOPATHY|HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY (DISORDER)
C0410223|T047|240103002|SNOMEDCT_US|HIV ASSOCIATED MYOPATHY |HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY (DISORDER)
C0410223|T047|240103002|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY|HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY (DISORDER)
C0410223|T047|240103002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY|HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY (DISORDER)
C0410223|T047|240103002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY |HUMAN IMMUNODEFICIENCY VIRUS MYOPATHY (DISORDER)
C0276500|T047|40780007|SNOMEDCT_US|HIV I INFECTION|HUMAN IMMUNODEFICIENCY VIRUS I INFECTION (DISORDER)
C0276500|T047|40780007|SNOMEDCT_US|HIV I INFECTION |HUMAN IMMUNODEFICIENCY VIRUS I INFECTION (DISORDER)
C0276500|T047|40780007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS I INFECTION|HUMAN IMMUNODEFICIENCY VIRUS I INFECTION (DISORDER)
C0276500|T047|40780007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS I INFECTION |HUMAN IMMUNODEFICIENCY VIRUS I INFECTION (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HIV LEUKOENCEPHALOPATHY |HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HIV LEUKOENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS LEUCOENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS LEUKOENCEPHALOPATHY |HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HUMAN IMMUNODEFIENCY VIRUS LEUCOENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS LEUCOENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS LEUKOENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HIV - HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HIV - HUMAN IMMUNODEFIENCY VIRUS LEUCOENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY |HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0338422|T047|230180003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS LEUKOENCEPHALOPATHY|HUMAN IMMUNODEFIENCY VIRUS LEUKOENCEPHALOPATHY (DISORDER)
C0276501|T047|79019005|SNOMEDCT_US|HIV II INFECTION|HUMAN IMMUNODEFICIENCY VIRUS II INFECTION (DISORDER)
C0276501|T047|79019005|SNOMEDCT_US|HIV II INFECTION |HUMAN IMMUNODEFICIENCY VIRUS II INFECTION (DISORDER)
C0276501|T047|79019005|SNOMEDCT_US|HIV 2 INFECTION|HUMAN IMMUNODEFICIENCY VIRUS II INFECTION (DISORDER)
C0276501|T047|79019005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS II INFECTION|HUMAN IMMUNODEFICIENCY VIRUS II INFECTION (DISORDER)
C0276501|T047|79019005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS II INFECTION |HUMAN IMMUNODEFICIENCY VIRUS II INFECTION (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|HIV ENCEPHALITIS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|AIDS WITH ENCEPHALITIS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|AIDS WITH ENCEPHALITIS |HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|HIV - HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|HUMAN IMMUNODEFIENCY VIRUS SUBACUTE ENCEPHALITIS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|HIV ENCEPHALITIS |HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS ENCEPHALITIS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS |HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS ENCEPHALITIS|HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0276548|T047|398329009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS ENCEPHALITIS |HUMAN IMMUNODEFIENCY VIRUS ENCEPHALITIS (DISORDER)
C0452189|T047|186723002|SNOMEDCT_US|HIV DISEASE RESULTING IN BURKITT'S LYMPHOMA|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HIV DISEASE RESULTING IN BURKITT'S LYMPHOMA |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HIV INFECTION RESULTING IN BURKITT'S LYMPHOMA|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HIV INFECTION RESULTING IN BURKITT'S LYMPHOMA |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN BURKITT'S LYMPHOMA |HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS DISEASE RESULTING IN BURKITT'S LYMPHOMA|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT LYMPHOMA|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HIV DISEASE; BURKITT|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|HIV DISEASE; LYMPHOMA, BURKITT|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|BURKITT; LYMPHOMA, RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0452189|T047|186723002|SNOMEDCT_US|LYMPHOMA; BURKITT, RESULTING FROM HIV DISEASE|HUMAN IMMUNODEFICIENCY VIRUS (HIV) DISEASE RESULTING IN BURKITT'S LYMPHOMA
C0276601|T047|5810003|SNOMEDCT_US|HIV INFECTION WITH INFECTION BY ANOTHER VIRUS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HIV INFECTION WITH INFECTION BY ANOTHER VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HIV INFECTION WITH INFECTION BY ANOTHER VIRUS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH INFECTION CAUSED BY ANOTHER VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH INFECTION CAUSED BY ANOTHER VIRUS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION CAUSED BY ANOTHER VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH INFECTION BY ANOTHER VIRUS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH INFECTION BY ANOTHER VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|HIV INFECTION WITH INFECTION CAUSED BY ANOTHER VIRUS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0276601|T047|5810003|SNOMEDCT_US|AIDS VIRUS WITH VIRAL INFECTION|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTION BY ANOTHER VIRUS
C0343756|T047|230201009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRAL MYELITIS|HUMAN IMMUNODEFICIENCY VIRUS MYELITIS (DISORDER)
C0343756|T047|230201009|SNOMEDCT_US|HIV MYELITIS|HUMAN IMMUNODEFICIENCY VIRUS MYELITIS (DISORDER)
C0343756|T047|230201009|SNOMEDCT_US|HIV MYELITIS |HUMAN IMMUNODEFICIENCY VIRUS MYELITIS (DISORDER)
C0343756|T047|230201009|SNOMEDCT_US|HIV - HUMAN IMMUNODEFICIENCY VIRUS MYELITIS|HUMAN IMMUNODEFICIENCY VIRUS MYELITIS (DISORDER)
C0343756|T047|230201009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS MYELITIS|HUMAN IMMUNODEFICIENCY VIRUS MYELITIS (DISORDER)
C0343756|T047|230201009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS MYELITIS |HUMAN IMMUNODEFICIENCY VIRUS MYELITIS (DISORDER)
C0456101|T047|276666007|SNOMEDCT_US|HIV CONGENITAL POSITIVE STATUS SYNDROME|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS POSITIVE STATUS SYNDROME (DISORDER)
C0456101|T047|276666007|SNOMEDCT_US|CONGENITAL HIV POSITIVE STATUS SYNDROME |CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS POSITIVE STATUS SYNDROME (DISORDER)
C0456101|T047|276666007|SNOMEDCT_US|CONGENITAL HIV POSITIVE STATUS SYNDROME|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS POSITIVE STATUS SYNDROME (DISORDER)
C0456101|T047|276666007|SNOMEDCT_US|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS POSITIVE STATUS SYNDROME|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS POSITIVE STATUS SYNDROME (DISORDER)
C0456101|T047|276666007|SNOMEDCT_US|HIV - CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS POSITIVE STATUS SYNDROME|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS POSITIVE STATUS SYNDROME (DISORDER)
C0456101|T047|276666007|SNOMEDCT_US|CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS POSITIVE STATUS SYNDROME |CONGENITAL HUMAN IMMUNODEFICIENCY VIRUS POSITIVE STATUS SYNDROME (DISORDER)
C0276599|T047|87117006|SNOMEDCT_US|HIV INFECTION WITH ACUTE LYMPHADENITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS
C0276599|T047|87117006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS
C0276599|T047|87117006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH ACUTE LYMPHADENITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS
C0276599|T047|87117006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH ACUTE LYMPHADENITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS
C0276599|T047|87117006|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS
C0276599|T047|87117006|SNOMEDCT_US|AIDS VIRUS WITH ACUTE LYMPHADENITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS
C0276599|T047|87117006|SNOMEDCT_US|HIV INFECTION WITH ACUTE LYMPHADENITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS
C0276599|T047|87117006|SNOMEDCT_US|AIDS VIRUS WITH ACUTE LYMPHADENITIS|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS
C0276599|T047|87117006|SNOMEDCT_US|HIV INFECTION WITH ACUTE LYMPHADENITIS |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH ACUTE LYMPHADENITIS
C0276602|T047|48794007|SNOMEDCT_US|HIV INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME
C0276602|T047|48794007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME
C0276602|T047|48794007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME
C0276602|T047|48794007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME
C0276602|T047|48794007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME
C0276602|T047|48794007|SNOMEDCT_US|HIV INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME
C0276602|T047|48794007|SNOMEDCT_US|HIV INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME
C0276602|T047|48794007|SNOMEDCT_US|AIDS VIRUS WITH "INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME"|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION WITH INFECTIOUS MONONUCLEOSIS-LIKE SYNDROME
C0343746|T047|186708007|SNOMEDCT_US|HIV INFECTION WITH SECONDARY CLINICALLY INFECTIOUS DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH SECONDARY CLINICAL INFECTIOUS DISEASE (DISORDER)
C0343746|T047|186708007|SNOMEDCT_US|HIV INFECTION WITH SECONDARY CLINICALLY INFECTIOUS DISEASE |HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH SECONDARY CLINICAL INFECTIOUS DISEASE (DISORDER)
C0343746|T047|186708007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH SECONDARY CLINICAL INFECTIOUS DISEASE|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH SECONDARY CLINICAL INFECTIOUS DISEASE (DISORDER)
C0343746|T047|186708007|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH SECONDARY CLINICAL INFECTIOUS DISEASE |HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH SECONDARY CLINICAL INFECTIOUS DISEASE (DISORDER)
C1319296|T047|405631006|SNOMEDCT_US|PEDIATRIC HIV INFECTION|HIV INFECTION, PEDIATRIC
C1319296|T047|405631006|SNOMEDCT_US|HIV INFECTION PEDIATRIC|HIV INFECTION, PEDIATRIC
C1319296|T047|405631006|SNOMEDCT_US|PEDIATRIC HIV INFECTION |HIV INFECTION, PEDIATRIC
C1319296|T047|405631006|SNOMEDCT_US|HIV INFECTION, PAEDIATRIC|HIV INFECTION, PEDIATRIC
C1319296|T047|405631006|SNOMEDCT_US|HIV INFECTION, PEDIATRIC|HIV INFECTION, PEDIATRIC
C1319296|T047|405631006|SNOMEDCT_US|PAEDIATRIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION|HIV INFECTION, PEDIATRIC
C1319296|T047|405631006|SNOMEDCT_US|PEDIATRIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION |HIV INFECTION, PEDIATRIC
C1319296|T047|405631006|SNOMEDCT_US|PEDIATRIC HUMAN IMMUNODEFICIENCY VIRUS INFECTION|HIV INFECTION, PEDIATRIC
C3840061|T047|10755671000119100|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS IN MOTHER COMPLICATING CHILDBIRTH |HIV (HUMAN IMMUNODEFICIENCY VIRUS) IN CHILDBIRTH
C3840061|T047|10755671000119100|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS IN MOTHER COMPLICATING CHILDBIRTH|HIV (HUMAN IMMUNODEFICIENCY VIRUS) IN CHILDBIRTH
C3840061|T047|10755671000119100|SNOMEDCT_US|HIV (HUMAN IMMUNODEFICIENCY VIRUS) IN CHILDBIRTH|HIV (HUMAN IMMUNODEFICIENCY VIRUS) IN CHILDBIRTH
C3874345|T047|76991000119109|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION CATEGORY B2 |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION CATEGORY B2 (DISORDER)
C3874345|T047|76991000119109|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION CATEGORY B2|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION CATEGORY B2 (DISORDER)
C3874330|T047|76981000119106|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION CATEGORY B1 |HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION CATEGORY B1 (DISORDER)
C3874330|T047|76981000119106|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION CATEGORY B1|HUMAN IMMUNODEFICIENCY VIRUS (HIV) INFECTION CATEGORY B1 (DISORDER)
C3874341|T047|72631000119101|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) II INFECTION CATEGORY B2|HUMAN IMMUNODEFICIENCY VIRUS (HIV) II INFECTION CATEGORY B2 (DISORDER)
C3874341|T047|72631000119101|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS (HIV) II INFECTION CATEGORY B2 |HUMAN IMMUNODEFICIENCY VIRUS (HIV) II INFECTION CATEGORY B2 (DISORDER)
C4076110|T047|713484001|SNOMEDCT_US|DISORDER OF RESPIRATORY SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|DISORDER OF RESPIRATORY SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076110|T047|713484001|SNOMEDCT_US|DISORDER OF RESPIRATORY SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |DISORDER OF RESPIRATORY SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076215|T047|713342008|SNOMEDCT_US|INFECTION CAUSED BY SALMONELLA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |SALMONELLOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076215|T047|713342008|SNOMEDCT_US|SALMONELLOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|SALMONELLOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076215|T047|713342008|SNOMEDCT_US|INFECTION CAUSED BY SALMONELLA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|SALMONELLOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4075735|T047|713731001|SNOMEDCT_US|FEVER OF UNKNOWN ORIGIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|PYREXIA OF UNKNOWN ORIGIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075735|T047|713731001|SNOMEDCT_US|PYREXIA OF UNKNOWN ORIGIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|PYREXIA OF UNKNOWN ORIGIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075735|T047|713731001|SNOMEDCT_US|PYREXIA OF UNKNOWN ORIGIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |PYREXIA OF UNKNOWN ORIGIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075750|T047|713732008|SNOMEDCT_US|INFECTION CAUSED BY ASPERGILLUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY ASPERGILLUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075750|T047|713732008|SNOMEDCT_US|ASPERGILLOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY ASPERGILLUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075750|T047|713732008|SNOMEDCT_US|INFECTION CAUSED BY ASPERGILLUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |INFECTION CAUSED BY ASPERGILLUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076090|T047|713506004|SNOMEDCT_US|NEURITIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|NEURITIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076090|T047|713506004|SNOMEDCT_US|NEURITIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |NEURITIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075393|T047|714464009|SNOMEDCT_US|IMMUNE RECONSTITUTION INFLAMMATORY SYNDROME CAUSED BY HUMAN IMMUNODEFICIENCY VIRUS INFECTION|IMMUNE RECONSTITUTION INFLAMMATORY SYNDROME CAUSED BY HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075393|T047|714464009|SNOMEDCT_US|IMMUNE RECONSTITUTION INFLAMMATORY SYNDROME CAUSED BY HUMAN IMMUNODEFICIENCY VIRUS INFECTION |IMMUNE RECONSTITUTION INFLAMMATORY SYNDROME CAUSED BY HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075812|T047|713733003|SNOMEDCT_US|INFECTION CAUSED BY HERPES ZOSTER VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY HERPES ZOSTER VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075812|T047|713733003|SNOMEDCT_US|HERPES ZOSTER INFECTION CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY HERPES ZOSTER VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075812|T047|713733003|SNOMEDCT_US|INFECTION CAUSED BY HERPES ZOSTER VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |INFECTION CAUSED BY HERPES ZOSTER VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075921|T047|713571008|SNOMEDCT_US|DISORDER OF CENTRAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |DISORDER OF CENTRAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075921|T047|713571008|SNOMEDCT_US|DISORDER OF CENTRAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|DISORDER OF CENTRAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4074813|T047|713729005|SNOMEDCT_US|COCCIDIOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY COCCIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4074813|T047|713729005|SNOMEDCT_US|INFECTION CAUSED BY COCCIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |INFECTION CAUSED BY COCCIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4074813|T047|713729005|SNOMEDCT_US|INFECTION CAUSED BY COCCIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY COCCIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076083|T047|713510001|SNOMEDCT_US|HEPATOMEGALY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|LARGE LIVER CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076083|T047|713510001|SNOMEDCT_US|ENLARGEMENT OF LIVER CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|LARGE LIVER CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076083|T047|713510001|SNOMEDCT_US|ENLARGEMENT OF LIVER CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |LARGE LIVER CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076083|T047|713510001|SNOMEDCT_US|LARGE LIVER CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|LARGE LIVER CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076016|T047|713527009|SNOMEDCT_US|DISORDER OF PERIPHERAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |DISORDER OF PERIPHERAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076016|T047|713527009|SNOMEDCT_US|DISORDER OF PERIPHERAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|DISORDER OF PERIPHERAL NERVOUS SYSTEM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075583|T047|713967004|SNOMEDCT_US|DISSEMINATED ATYPICAL INFECTION CAUSED BY MYCOBACTERIUM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|DISSEMINATED ATYPICAL INFECTION CAUSED BY MYCOBACTERIUM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075583|T047|713967004|SNOMEDCT_US|DISSEMINATED ATYPICAL INFECTION CAUSED BY MYCOBACTERIUM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |DISSEMINATED ATYPICAL INFECTION CAUSED BY MYCOBACTERIUM CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076290|T047|713275003|SNOMEDCT_US|SPLENOMEGALY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |SPLENOMEGALY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076290|T047|713275003|SNOMEDCT_US|SPLENOMEGALY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|SPLENOMEGALY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076117|T047|713490002|SNOMEDCT_US|INFECTION CAUSED BY PNEUMOCYSTIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|PNEUMOCYSTOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076117|T047|713490002|SNOMEDCT_US|INFECTION CAUSED BY PNEUMOCYSTIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |PNEUMOCYSTOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076117|T047|713490002|SNOMEDCT_US|PNEUMOCYSTOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|PNEUMOCYSTOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076026|T047|713532005|SNOMEDCT_US|INFECTIVE ARTHRITIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |INFECTIVE ARTHRITIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076026|T047|713532005|SNOMEDCT_US|INFECTIVE ARTHRITIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTIVE ARTHRITIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075796|T047|713730000|SNOMEDCT_US|INFECTION CAUSED BY HERPES SIMPLEX VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |INFECTION CAUSED BY HERPES SIMPLEX VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075796|T047|713730000|SNOMEDCT_US|HERPES SIMPLEX VIRUS INFECTION CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY HERPES SIMPLEX VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075796|T047|713730000|SNOMEDCT_US|INFECTION CAUSED BY HERPES SIMPLEX VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY HERPES SIMPLEX VIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075629|T047|713881001|SNOMEDCT_US|MICROSPORIDIOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY MICROSPORIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075629|T047|713881001|SNOMEDCT_US|INFECTION CAUSED BY MICROSPORIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |INFECTION CAUSED BY MICROSPORIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075629|T047|713881001|SNOMEDCT_US|INFECTION CAUSED BY MICROSPORIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY MICROSPORIDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075653|T047|713880000|SNOMEDCT_US|OPPORTUNISTIC MYCOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|OPPORTUNISTIC MYCOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075653|T047|713880000|SNOMEDCT_US|OPPORTUNISTIC MYCOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |OPPORTUNISTIC MYCOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076086|T047|713497004|SNOMEDCT_US|CANDIDIASIS OF MOUTH CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |CANDIDIASIS OF MOUTH CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076086|T047|713497004|SNOMEDCT_US|CANDIDIASIS OF MOUTH CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|CANDIDIASIS OF MOUTH CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076155|T047|713444005|SNOMEDCT_US|HEMOPHAGOCYTIC SYNDROME CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|HEMOPHAGOCYTIC SYNDROME CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076155|T047|713444005|SNOMEDCT_US|HEMOPHAGOCYTIC SYNDROME CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |HEMOPHAGOCYTIC SYNDROME CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075982|T047|713545009|SNOMEDCT_US|NOCARDIOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY NOCARDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075982|T047|713545009|SNOMEDCT_US|INFECTION CAUSED BY NOCARDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |INFECTION CAUSED BY NOCARDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075982|T047|713545009|SNOMEDCT_US|INFECTION CAUSED BY NOCARDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY NOCARDIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076042|T047|713531003|SNOMEDCT_US|VISUAL IMPAIRMENT CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |VISUAL IMPAIRMENT CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076042|T047|713531003|SNOMEDCT_US|VISUAL IMPAIRMENT CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|VISUAL IMPAIRMENT CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075766|T047|713722001|SNOMEDCT_US|INFECTION CAUSED BY CYTOMEGALOVIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY CYTOMEGALOVIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075766|T047|713722001|SNOMEDCT_US|INFECTION CAUSED BY CYTOMEGALOVIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |INFECTION CAUSED BY CYTOMEGALOVIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075766|T047|713722001|SNOMEDCT_US|CYTOMEGALOVIRUS INFECTION CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY CYTOMEGALOVIRUS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075814|T047|713734009|SNOMEDCT_US|DERMATOPHYTOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY DERMATOPHYTE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075814|T047|713734009|SNOMEDCT_US|INFECTION CAUSED BY DERMATOPHYTE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|INFECTION CAUSED BY DERMATOPHYTE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075814|T047|713734009|SNOMEDCT_US|INFECTION CAUSED BY DERMATOPHYTE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |INFECTION CAUSED BY DERMATOPHYTE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076115|T047|713489006|SNOMEDCT_US|POLYNEUROPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|POLYNEUROPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076115|T047|713489006|SNOMEDCT_US|POLYNEUROPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |POLYNEUROPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076275|T047|713299003|SNOMEDCT_US|DISORDER OF EYE PROPER CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|DISORDER OF EYE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076275|T047|713299003|SNOMEDCT_US|DISORDER OF EYE PROPER CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |DISORDER OF EYE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076275|T047|713299003|SNOMEDCT_US|DISORDER OF EYE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|DISORDER OF EYE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076216|T047|713349004|SNOMEDCT_US|ANAEMIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|ANEMIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076216|T047|713349004|SNOMEDCT_US|ANEMIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |ANEMIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076216|T047|713349004|SNOMEDCT_US|ANEMIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|ANEMIA CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076274|T047|713298006|SNOMEDCT_US|HEART DISEASE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |HEART DISEASE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076274|T047|713298006|SNOMEDCT_US|HEART DISEASE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|HEART DISEASE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075781|T047|713339002|SNOMEDCT_US|INFECTION CAUSED BY STRONGYLOIDES CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |STRONGYLOIDIASIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4075781|T047|713339002|SNOMEDCT_US|INFECTION CAUSED BY STRONGYLOIDES CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|STRONGYLOIDIASIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4075781|T047|713339002|SNOMEDCT_US|STRONGYLOIDIASIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|STRONGYLOIDIASIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076265|T047|713300006|SNOMEDCT_US|DISORDER OF GASTROINTESTINAL TRACT CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|DISORDER OF GASTROINTESTINAL TRACT CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076265|T047|713300006|SNOMEDCT_US|DISORDER OF GASTROINTESTINAL TRACT CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |DISORDER OF GASTROINTESTINAL TRACT CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076101|T047|713507008|SNOMEDCT_US|LYMPHADENOPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|LYMPHADENOPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076101|T047|713507008|SNOMEDCT_US|LYMPHADENOPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |LYMPHADENOPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075933|T047|713572001|SNOMEDCT_US|MALIGNANT NEOPLASTIC DISEASE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |MALIGNANT NEOPLASTIC DISEASE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4075933|T047|713572001|SNOMEDCT_US|MALIGNANT NEOPLASTIC DISEASE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|MALIGNANT NEOPLASTIC DISEASE CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076103|T047|713504001|SNOMEDCT_US|NEPHROPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|NEPHROPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076103|T047|713504001|SNOMEDCT_US|DISORDER OF KIDNEY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|NEPHROPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076103|T047|713504001|SNOMEDCT_US|DISORDER OF KIDNEY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |NEPHROPATHY CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION
C4076222|T047|713340000|SNOMEDCT_US|DISORDER OF SKIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |DISORDER OF SKIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076222|T047|713340000|SNOMEDCT_US|DISORDER OF SKIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|DISORDER OF SKIN CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076020|T047|713530002|SNOMEDCT_US|AGRANULOCYTOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION |AGRANULOCYTOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C4076020|T047|713530002|SNOMEDCT_US|AGRANULOCYTOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION|AGRANULOCYTOSIS CO-OCCURRENT WITH HUMAN IMMUNODEFICIENCY VIRUS INFECTION (DISORDER)
C0856916|T047|95892003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH PERSISTENT GENERALISED LYMPHADENOPATHY|PERSISTENT GENERALIZED LYMPHADENOPATHY (DISORDER)
C0856916|T047|95892003|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS INFECTION WITH PERSISTENT GENERALIZED LYMPHADENOPATHY|PERSISTENT GENERALIZED LYMPHADENOPATHY (DISORDER)
C0686714|T047|91923005|SNOMEDCT_US|AIDS VIRUS INFECTION ASSOCIATED WITH PREGNANCY |ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) VIRUS INFECTION ASSOCIATED WITH PREGNANCY
C0686714|T047|91923005|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) VIRUS INFECTION ASSOCIATED WITH PREGNANCY|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) VIRUS INFECTION ASSOCIATED WITH PREGNANCY
C0686714|T047|91923005|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME VIRUS INFECTION ASSOCIATED WITH PREGNANCY |ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) VIRUS INFECTION ASSOCIATED WITH PREGNANCY
C0686714|T047|91923005|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) VIRUS INFECTION ASSOCIATED WITH PREGNANCY |ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) VIRUS INFECTION ASSOCIATED WITH PREGNANCY
C0686714|T047|91923005|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME VIRUS INFECTION ASSOCIATED WITH PREGNANCY|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) VIRUS INFECTION ASSOCIATED WITH PREGNANCY
C0686714|T047|91923005|SNOMEDCT_US|AIDS VIRUS INFECTION ASSOCIATED WITH PREGNANCY|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) VIRUS INFECTION ASSOCIATED WITH PREGNANCY
C0559284|T047|281390005|SNOMEDCT_US|HIV-RELATED GUT DISEASE - CAUSE UNKNOWN |HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED GUT DISEASE - CAUSE UNKNOWN
C0559284|T047|281390005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED GUT DISEASE - CAUSE UNKNOWN |HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED GUT DISEASE - CAUSE UNKNOWN
C0559284|T047|281390005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-RELATED GUT DISEASE - CAUSE UNKNOWN |HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED GUT DISEASE - CAUSE UNKNOWN
C0559284|T047|281390005|SNOMEDCT_US|HIV-RELATED GUT DISEASE - CAUSE UNKNOWN|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED GUT DISEASE - CAUSE UNKNOWN
C0559284|T047|281390005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED GUT DISEASE - CAUSE UNKNOWN|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED GUT DISEASE - CAUSE UNKNOWN
C0559284|T047|281390005|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-RELATED GUT DISEASE - CAUSE UNKNOWN|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED GUT DISEASE - CAUSE UNKNOWN
C0559283|T047|281388009|SNOMEDCT_US|HIV-RELATED SCLEROSING CHOLANGITIS |HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS
C0559283|T047|281388009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS
C0559283|T047|281388009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-RELATED SCLEROSING CHOLANGITIS |HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS
C0559283|T047|281388009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-RELATED SCLEROSING CHOLANGITIS|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS
C0559283|T047|281388009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS |HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS
C0559283|T047|281388009|SNOMEDCT_US|SCLEROSING CHOLANGITIS HUMAN IMMUNODEFICIENCY VIRUS-REALTED|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS
C0559283|T047|281388009|SNOMEDCT_US|HUMAN IMMUNODEFICIENCY VIRUS-RELATED SCLEROSING CHOLANGITIS |HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS
C0559283|T047|281388009|SNOMEDCT_US|HIV-RELATED SCLEROSING CHOLANGITIS|HUMAN IMMUNODEFICIENCY VIRUS HIV-RELATED SCLEROSING CHOLANGITIS
C0276605|T047|78466009|SNOMEDCT_US|POSITIVE SEROLOGICAL OR VIRAL CULTURE FINDINGS FOR HUMAN UMMUNODEFICIENCY VIRUS|POSITIVE SEROLOGICAL OR VIRAL CULTURE FINDINGS FOR HUMAN UMMUNODEFICIENCY VIRUS
C0276605|T047|78466009|SNOMEDCT_US|POSITIVE SEROLOGICAL AND/OR VIRAL CULTURE FINDINGS FOR HUMAN IMMUNODEFICIENCY VIRUS |POSITIVE SEROLOGICAL OR VIRAL CULTURE FINDINGS FOR HUMAN UMMUNODEFICIENCY VIRUS
C0276605|T047|78466009|SNOMEDCT_US|POSITIVE SEROLOGICAL AND/OR VIRAL CULTURE FINDINGS FOR HUMAN IMMUNODEFICIENCY VIRUS|POSITIVE SEROLOGICAL OR VIRAL CULTURE FINDINGS FOR HUMAN UMMUNODEFICIENCY VIRUS
C0276605|T047|78466009|SNOMEDCT_US|POSITIVE SEROLOGICAL OR VIRAL CULTURE FINDINGS FOR HUMAN IMMUNODEFICIENCY VIRUS|POSITIVE SEROLOGICAL OR VIRAL CULTURE FINDINGS FOR HUMAN UMMUNODEFICIENCY VIRUS
C0348204|T047|187439001|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER BACTERIAL INFECTIONS|[X]HIV DISEASE RESULTING IN OTHER BACTERIAL INFECTIONS (DISORDER)
C0348204|T047|187439001|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER BACTERIAL INFECTIONS|[X]HIV DISEASE RESULTING IN OTHER BACTERIAL INFECTIONS (DISORDER)
C0348204|T047|187439001|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER BACTERIAL INFECTIONS |[X]HIV DISEASE RESULTING IN OTHER BACTERIAL INFECTIONS (DISORDER)
C0348204|T047|187439001|SNOMEDCT_US|BACTERIAL; INFECTION, RESULTING FROM HIV DISEASE|[X]HIV DISEASE RESULTING IN OTHER BACTERIAL INFECTIONS (DISORDER)
C0348204|T047|187439001|SNOMEDCT_US|INFECTION; BACTERIAL, RESULTING FROM HIV DISEASE|[X]HIV DISEASE RESULTING IN OTHER BACTERIAL INFECTIONS (DISORDER)
C0348212|T047|187448006|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS (DISORDER)
C0348212|T047|187448006|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS (DISORDER)
C0348212|T047|187448006|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS |[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER MYCOSES|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER MYCOSES |[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER MYCOSES|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|HIV DISEASE; MYCOSIS|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|HIV DISEASE; RESULTING IN, INFECTION, FUNGUS|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|HIV DISEASE; RESULTING IN, INFECTION, MYCOTIC|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|HIV DISEASE; RESULTING IN, MYCOSIS|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|FUNGUS; INFECTION, RESULTING FROM HIV DISEASE|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|INFECTION; FUNGUS, RESULTING FROM HIV DISEASE|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|INFECTION; MYCOTIC, RESULTING FROM HIV DISEASE|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|MYCOSIS; RESULTING FROM HIV DISEASE|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348206|T047|187442007|SNOMEDCT_US|MYCOTIC; INFECTION, RESULTING FROM HIV DISEASE|[X]HIV DISEASE RESULTING IN OTHER MYCOSES (DISORDER)
C0348210|T047|187446005|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER NON-HODGKIN'S LYMPHOMA|[X]HIV DISEASE RESULTING IN OTHER NON-HODGKIN'S LYMPHOMA (DISORDER)
C0348210|T047|187446005|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER NON-HODGKIN'S LYMPHOMA |[X]HIV DISEASE RESULTING IN OTHER NON-HODGKIN'S LYMPHOMA (DISORDER)
C0276555|T047|111888008|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER SPECIFIED CONDITIONS|AIDS WITH OTHER SPECIFIED CONDITIONS (DISORDER)
C0276555|T047|111888008|SNOMEDCT_US|AIDS WITH OTHER SPECIFIED CONDITIONS -RETIRED-|AIDS WITH OTHER SPECIFIED CONDITIONS (DISORDER)
C0276555|T047|111888008|SNOMEDCT_US|AIDS WITH OTHER SPECIFIED CONDITIONS|AIDS WITH OTHER SPECIFIED CONDITIONS (DISORDER)
C0276555|T047|111888008|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER SPECIFIED CONDITIONS |AIDS WITH OTHER SPECIFIED CONDITIONS (DISORDER)
C0276555|T047|111888008|SNOMEDCT_US|AIDS WITH OTHER SPECIFIED CONDITIONS |AIDS WITH OTHER SPECIFIED CONDITIONS (DISORDER)
C0276555|T047|111888008|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER SPECIFIED CONDITIONS|AIDS WITH OTHER SPECIFIED CONDITIONS (DISORDER)
C0348205|T047|187441000|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER VIRAL INFECTIONS|[X]HIV DISEASE RESULTING IN OTHER VIRAL INFECTIONS (DISORDER)
C0348205|T047|187441000|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER VIRAL INFECTIONS|[X]HIV DISEASE RESULTING IN OTHER VIRAL INFECTIONS (DISORDER)
C0348205|T047|187441000|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER VIRAL INFECTIONS |[X]HIV DISEASE RESULTING IN OTHER VIRAL INFECTIONS (DISORDER)
C0348215|T047|186710009|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN HEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NOT ELSEWHERE CLASSIFIED|[X]HIV DISEASE RESULTING IN HAEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NOT ELSEWHERE CLASSIFIED (DISORDER)
C0348215|T047|186710009|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN HAEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NOT ELSEWHERE CLASSIFIED|[X]HIV DISEASE RESULTING IN HAEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NOT ELSEWHERE CLASSIFIED (DISORDER)
C0348215|T047|186710009|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN HAEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NOT ELSEWHERE CLASSIFIED |[X]HIV DISEASE RESULTING IN HAEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NOT ELSEWHERE CLASSIFIED (DISORDER)
C0348215|T047|186710009|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN HEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NOT ELSEWHERE CLASSIFIED |[X]HIV DISEASE RESULTING IN HAEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NOT ELSEWHERE CLASSIFIED (DISORDER)
C0348215|T047|186710009|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN HAEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NEC  IN SNOMEDCT_US_2016_03_01|[X]HIV DISEASE RESULTING IN HAEMATOLOGICAL AND IMMUNOLOGICAL ABNORMALITIES, NOT ELSEWHERE CLASSIFIED (DISORDER)
C0348211|T047|187447001|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE (DISORDER)
C0348211|T047|187447001|SNOMEDCT_US|HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE (DISORDER)
C0348211|T047|187447001|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE (DISORDER)
C0348211|T047|187447001|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE |[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE (DISORDER)
C0348211|T047|187447001|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE |[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE (DISORDER)
C0348211|T047|187447001|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HAEMATOPOIETIC AND RELATED TISSUE|[X]HIV DISEASE RESULTING IN OTHER MALIGNANT NEOPLASMS OF LYMPHOID, HEMATOPOIETIC AND RELATED TISSUE (DISORDER)
C0348214|T047|186711008|SNOMEDCT_US|HIV DISEASE RESULTING IN MULTIPLE DISEASES CLASSIFIED ELSEWHERE|[X]HIV DISEASE RESULTING IN MULTIPLE DISEASES CLASSIFIED ELSEWHERE (DISORDER)
C0348214|T047|186711008|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN MULTIPLE DISEASES CLASSIFIED ELSEWHERE |[X]HIV DISEASE RESULTING IN MULTIPLE DISEASES CLASSIFIED ELSEWHERE (DISORDER)
C0348214|T047|186711008|SNOMEDCT_US|[X]HIV DISEASE RESULTING IN MULTIPLE DISEASES CLASSIFIED ELSEWHERE|[X]HIV DISEASE RESULTING IN MULTIPLE DISEASES CLASSIFIED ELSEWHERE (DISORDER)
C0348214|T047|186711008|SNOMEDCT_US|HIV DISEASE; RESULTING IN, MULTIPLE, DISEASES CLASSIFIED ELSEWHERE|[X]HIV DISEASE RESULTING IN MULTIPLE DISEASES CLASSIFIED ELSEWHERE (DISORDER)
C0393489|T047|230202002|SNOMEDCT_US|CANNOT FIND ANY REFERENCES OF THIS BEING ASSOCIAED WITH ANY OTHER DIEASES BESIDES HIV SO WILL KEEP IT|VACUOLAR MYELOPATHY (DISORDER)
C0393489|T047|230202002|SNOMEDCT_US|VACUOLAR MYELOPATHY |VACUOLAR MYELOPATHY (DISORDER)
C0456100|T047|276665006|SNOMEDCT_US|AIDS - CONGENITAL ACQUIRED IMMUNE DEFICIENCY SYNDROME|CONGENITAL ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0456100|T047|276665006|SNOMEDCT_US|CONGENITAL ACQUIRED IMMUNE DEFICIENCY SYNDROME|CONGENITAL ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C0456100|T047|276665006|SNOMEDCT_US|CONGENITAL ACQUIRED IMMUNE DEFICIENCY SYNDROME |CONGENITAL ACQUIRED IMMUNE DEFICIENCY SYNDROME (DISORDER)
C1562915|T047|416491000|SNOMEDCT_US|UVEITIS IMMUNE RECOVERY|IMMUNE RECOVERY UVEITIS (DISORDER)
C1562915|T047|416491000|SNOMEDCT_US|IMMUNE RECOVERY UVEITIS|IMMUNE RECOVERY UVEITIS (DISORDER)
C1562915|T047|416491000|SNOMEDCT_US|IMMUNE RECOVERY UVEITIS |IMMUNE RECOVERY UVEITIS (DISORDER)
C1562915|T047|416491000|SNOMEDCT_US|IMMUNE RECOVERY UVEITIS |IMMUNE RECOVERY UVEITIS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|AIDS WITH VIRAL PNEUMONIA |VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|VIRAL PNEUMONIA ASSOCIATED WITH AIDS|VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) WITH VIRAL PNEUMONIA|VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|AIDS WITH VIRAL PNEUMONIA|VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME (AIDS) WITH VIRAL PNEUMONIA |VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|VIRAL PNEUMONIA ASSOCIATED WITH AIDS |VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|PNEUMONIA VIRAL ASSOCIATED WITH AIDS|VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|VIRAL PNEUMONIA ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME|VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|VIRAL PNEUMONIA ASSOCIATED WITH ACQUIRED IMMUNODEFICIENCY SYNDROME |VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|VIRAL PNEUMONIA ASSOCIATED WITH AIDS |VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C0276528|T047|421508002|SNOMEDCT_US|AIDS WITH VIRAL PNEUMONIA, NOS|VIRAL PNEUMONIA ASSOCIATED WITH AIDS (DISORDER)
C1720105|T047|420721002|SNOMEDCT_US|AIDS-ASSOCIATED DISORDER|AIDS COMPLICATION
C1720105|T047|420721002|SNOMEDCT_US|COMPLICATION OF AIDS|AIDS COMPLICATION
C1720105|T047|420721002|SNOMEDCT_US|AIDS COMPLICATION|AIDS COMPLICATION
C1720105|T047|420721002|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME-ASSOCIATED DISORDER |AIDS COMPLICATION
C1720105|T047|420721002|SNOMEDCT_US|AIDS-ASSOCIATED DISORDER |AIDS COMPLICATION
C1720105|T047|420721002|SNOMEDCT_US|ACQUIRED IMMUNODEFICIENCY SYNDROME-ASSOCIATED DISORDER|AIDS COMPLICATION
