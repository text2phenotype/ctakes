C0010403|T047|30911005|SNOMEDCT_US|CRYOGLOBULINEMIA|CRYOGLOBULINEMIA (DISORDER)
C0543697|T047||SNOMEDCT_US|MIXED CRYOGLOBULINEMIA
C0543697|T047||SNOMEDCT_US|MIXED CRYOGLOBULINAEMIA
C0010403|T047|30911005|SNOMEDCT_US|CRYOGLOBULINEMIA|CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOGLOBULINEMIAS|CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOGLOBULINAEMIA|CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOGLOBULINEMIA |CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOGLOBULINEMIA [DISEASE/FINDING]|CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOGLOBULINEMIA |CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOIMMUNOGLOBULINAEMIA|CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOIMMUNOGLOBULINEMIA|CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOGLOBULINEMIA, NOS|CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOIMMUNOGLOBULINEMIA, NOS|CRYOGLOBULINEMIA (DISORDER)
C0010403|T047|30911005|SNOMEDCT_US|CRYOGLOBULINAEMIA, NOS|CRYOGLOBULINEMIA (DISORDER)
C0340992|T047|190815001|SNOMEDCT_US|CRYOGLOBULINEMIC VASCULITIS |CRYOGLOBULINEMIC VASCULITIS (DISORDER)
C0340992|T047|190815001|SNOMEDCT_US|CRYOGLOBULINEMIC VASCULITIS|CRYOGLOBULINEMIC VASCULITIS (DISORDER)
C0340992|T047|190815001|SNOMEDCT_US|CRYOGLOBULINAEMIC VASCULITIS|CRYOGLOBULINEMIC VASCULITIS (DISORDER)
C0340992|T047|190815001|SNOMEDCT_US|CRYOGLOBULINEMIC VASCULITIS |CRYOGLOBULINEMIC VASCULITIS (DISORDER)
C0340992|T047|190815001|SNOMEDCT_US|CRYOGLOBULINEMIC; VASCULITIS|CRYOGLOBULINEMIC VASCULITIS (DISORDER)
C0340992|T047|190815001|SNOMEDCT_US|VASCULITIS; CRYOGLOBULINEMIC|CRYOGLOBULINEMIC VASCULITIS (DISORDER)
C0340979|T047|190814002|SNOMEDCT_US|CRYOGLOBULINEMIC PURPURA|CRYOGLOBULINEMIC PURPURA (DISORDER)
C0340979|T047|190814002|SNOMEDCT_US|CRYOGLOBULINEMIC PURPURA |CRYOGLOBULINEMIC PURPURA (DISORDER)
C0340979|T047|190814002|SNOMEDCT_US|CRYOGLOBULINAEMIC PURPURA|CRYOGLOBULINEMIC PURPURA (DISORDER)
C0340979|T047|190814002|SNOMEDCT_US|CRYOGLOBULINEMIC PURPURA |CRYOGLOBULINEMIC PURPURA (DISORDER)
C0340979|T047|190814002|SNOMEDCT_US|CRYOGLOBULINEMIC; PURPURA|CRYOGLOBULINEMIC PURPURA (DISORDER)
C0340979|T047|190814002|SNOMEDCT_US|PURPURA; CRYOGLOBULINEMIC|CRYOGLOBULINEMIC PURPURA (DISORDER)
C0343208|T047|239947001|SNOMEDCT_US|MIXED ESSENTIAL CRYOGLOBULINEMIA |ESSENTIAL MIXED CRYOGLOBULINEMIA (DISORDER)
C0343208|T047|239947001|SNOMEDCT_US|MIXED ESSENTIAL CRYOGLOBULINEMIA|ESSENTIAL MIXED CRYOGLOBULINEMIA (DISORDER)
C0343208|T047|239947001|SNOMEDCT_US|ESSENTIAL MIXED CRYOGLOBULINEMIA|ESSENTIAL MIXED CRYOGLOBULINEMIA (DISORDER)
C0343208|T047|239947001|SNOMEDCT_US|ESSENTIAL MIXED CRYOGLOBULINAEMIA|ESSENTIAL MIXED CRYOGLOBULINEMIA (DISORDER)
C0343208|T047|239947001|SNOMEDCT_US|ESSENTIAL CRYOGLOBULINAEMIC VASCULITIS|ESSENTIAL MIXED CRYOGLOBULINEMIA (DISORDER)
C0343208|T047|239947001|SNOMEDCT_US|ESSENTIAL CRYOGLOBULINEMIC VASCULITIS|ESSENTIAL MIXED CRYOGLOBULINEMIA (DISORDER)
C0343208|T047|239947001|SNOMEDCT_US|ESSENTIAL MIXED CRYOGLOBULINEMIA |ESSENTIAL MIXED CRYOGLOBULINEMIA (DISORDER)
C0272263|T047|10934005|SNOMEDCT_US|CRYOFIBRINOGENEMIA|CRYOFIBRINOGENEMIA (DISORDER)
C0272263|T047|10934005|SNOMEDCT_US|CRYOFIBRINOGENAEMIA|CRYOFIBRINOGENEMIA (DISORDER)
C0272263|T047|10934005|SNOMEDCT_US|CRYOFIBRINOGENEMIA |CRYOFIBRINOGENEMIA (DISORDER)
C0272263|T047|10934005|SNOMEDCT_US|CRYOFIBRINOGENEMIA, NOS|CRYOFIBRINOGENEMIA (DISORDER)
C1852456|T047||SNOMEDCT_US|CRYOGLOBULINEMIA, FAMILIAL MIXED
C1852456|T047||SNOMEDCT_US|MELTZER SYNDROME
C1852457|T047||SNOMEDCT_US|CRYOFIBRINOGENEMIA, FAMILIAL PRIMARY
C0272261|T047|57390009|SNOMEDCT_US|MIXED CRYOIMMUNOGLOBULINEMIA WITH MONOCLONAL COMPONENT|MIXED CRYOIMMUNOGLOBULINEMIA WITH MONOCLONAL COMPONENT (DISORDER)
C0272261|T047|57390009|SNOMEDCT_US|MIXED CRYOIMMUNOGLOBULINAEMIA WITH MONOCLONAL COMPONENT|MIXED CRYOIMMUNOGLOBULINEMIA WITH MONOCLONAL COMPONENT (DISORDER)
C0272261|T047|57390009|SNOMEDCT_US|MIXED CRYOIMMUNOGLOBULINEMIA WITH MONOCLONAL COMPONENT |MIXED CRYOIMMUNOGLOBULINEMIA WITH MONOCLONAL COMPONENT (DISORDER)
C0272262|T047|44371002|SNOMEDCT_US|MIXED POLYCLONAL CRYOIMMUNOGLOBULINEMIA|MIXED POLYCLONAL CRYOIMMUNOGLOBULINEMIA (DISORDER)
C0272262|T047|44371002|SNOMEDCT_US|MIXED POLYCLONAL CRYOIMMUNOGLOBULINAEMIA|MIXED POLYCLONAL CRYOIMMUNOGLOBULINEMIA (DISORDER)
C0272262|T047|44371002|SNOMEDCT_US|MIXED POLYCLONAL CRYOIMMUNOGLOBULINEMIA |MIXED POLYCLONAL CRYOIMMUNOGLOBULINEMIA (DISORDER)
C0272260|T047|38675009|SNOMEDCT_US|MONOCLONAL CRYOIMMUNOGLOBULINEMIA|MONOCLONAL CRYOIMMUNOGLOBULINEMIA (DISORDER)
C0272260|T047|38675009|SNOMEDCT_US|MONOCLONAL CRYOIMMUNOGLOBULINAEMIA|MONOCLONAL CRYOIMMUNOGLOBULINEMIA (DISORDER)
C0272260|T047|38675009|SNOMEDCT_US|MONOCLONAL CRYOIMMUNOGLOBULINEMIA |MONOCLONAL CRYOIMMUNOGLOBULINEMIA (DISORDER)
C0272258|T047|11352009|SNOMEDCT_US|PRIMARY CRYOGLOBULINEMIA|PRIMARY CRYOGLOBULINEMIA (DISORDER)
C0272258|T047|11352009|SNOMEDCT_US|PRIMARY CRYOGLOBULINAEMIA|PRIMARY CRYOGLOBULINEMIA (DISORDER)
C0272258|T047|11352009|SNOMEDCT_US|PRIMARY CRYOGLOBULINEMIA |PRIMARY CRYOGLOBULINEMIA (DISORDER)
C0272259|T047|28807005|SNOMEDCT_US|SECONDARY CRYOGLOBULINEMIA|SECONDARY CRYOGLOBULINEMIA (DISORDER)
C0272259|T047|28807005|SNOMEDCT_US|SECONDARY CRYOGLOBULINAEMIA|SECONDARY CRYOGLOBULINEMIA (DISORDER)
C0272259|T047|28807005|SNOMEDCT_US|SECONDARY CRYOGLOBULINEMIA |SECONDARY CRYOGLOBULINEMIA (DISORDER)
C1384927|T047||SNOMEDCT_US|DISEASE (OR DISORDER); GLOMERULAR, IN CRYOGLOBULINEMIA (ETIOLOGY)
C1384927|T047||SNOMEDCT_US|DISEASE (OR DISORDER); GLOMERULAR, IN CRYOGLOBULINEMIA (MANIFESTATION)
C1394252|T047||SNOMEDCT_US|CRYOGLOBULINEMIA; WITH LUNG INVOLVEMENT (ETIOLOGY)
C1394252|T047||SNOMEDCT_US|CRYOGLOBULINEMIA; WITH LUNG INVOLVEMENT (MANIFESTATION)
C1394252|T047||SNOMEDCT_US|DISEASE (OR DISORDER); LUNG, IN CRYOGLOBULINEMIA (ETIOLOGY)
C1394252|T047||SNOMEDCT_US|DISEASE (OR DISORDER); LUNG, IN CRYOGLOBULINEMIA (MANIFESTATION)
C1394252|T047||SNOMEDCT_US|LUNG; CRYOGLOBULINEMIA (ETIOLOGY)
C1394252|T047||SNOMEDCT_US|LUNG; CRYOGLOBULINEMIA (MANIFESTATION)
C1394252|T047||SNOMEDCT_US|LUNG; DISEASE, IN CRYOGLOBULINEMIA (MANIFESTATION)
C1385201|T047||SNOMEDCT_US|DISEASE (OR DISORDER); TUBULO-INTERSTITIAL, MIXED CRYOGLOBULINEMIA (ETIOLOGY)
C1385201|T047||SNOMEDCT_US|DISEASE (OR DISORDER); TUBULO-INTERSTITIAL, MIXED CRYOGLOBULINEMIA (MANIFESTATION)
C1394251|T047||SNOMEDCT_US|CRYOGLOBULINEMIA; GLOMERULONEPHRITIS (ETIOLOGY)
C1394251|T047||SNOMEDCT_US|CRYOGLOBULINEMIA; GLOMERULONEPHRITIS (MANIFESTATION)
C1394251|T047||SNOMEDCT_US|GLOMERULONEPHRITIS; CRYOGLOBULINEMIA (ETIOLOGY)
C1394251|T047||SNOMEDCT_US|GLOMERULONEPHRITIS; CRYOGLOBULINEMIA (MANIFESTATION)
C1394253|T047||SNOMEDCT_US|CRYOGLOBULINEMIA; PYELONEPHRITIS (ETIOLOGY)
C1394253|T047||SNOMEDCT_US|CRYOGLOBULINEMIA; PYELONEPHRITIS (MANIFESTATION)
C1394253|T047||SNOMEDCT_US|PYELONEPHRITIS; CRYOGLOBULINEMIA (ETIOLOGY)
C1394253|T047||SNOMEDCT_US|PYELONEPHRITIS; CRYOGLOBULINEMIA (MANIFESTATION)
C1398770|T047||SNOMEDCT_US|GLOMERULAR; DISEASE, IN CRYOGLOBULINEMIA (ETIOLOGY)
C1398770|T047||SNOMEDCT_US|GLOMERULAR; DISEASE, IN CRYOGLOBULINEMIA (MANIFESTATION)
C1407782|T047||SNOMEDCT_US|TUBULO-INTERSTITIAL; DISEASE, MIXED CRYOGLOBULINEMIA (ETIOLOGY)
C1407782|T047||SNOMEDCT_US|TUBULO-INTERSTITIAL; DISEASE, MIXED CRYOGLOBULINEMIA (MANIFESTATION)
