# CUI|TUI|CODE|SAB|TEXT|PREF_TEXT
# HBG - NOT FOUND
C0337443|T059|25197003|SNOMEDCT_US|SODIUM|SODIUM MEASUREMENT
C0202194|T059|59573005|SNOMEDCT_US|POTASSIUM|POTASSIUM MEASUREMENT
C0202059|T059|88645003|SNOMEDCT_US|BICARBONATE|BICARBONATE MEASUREMENT
C0201889|T059|25469001|SNOMEDCT_US|ANION GAP|ANION GAP MEASUREMENT
C0005845|T059|105011006|SNOMEDCT_US|UREA NITROGEN|BLOOD UREA NITROGEN MEASUREMENT
C0202239|T059|86228006|SNOMEDCT_US|URIC ACID|URIC ACID MEASUREMENT
C0202035|T059|69480007|SNOMEDCT_US|GAMMA GLUTAMYL TRANSFERASE|GAMMA GLUTAMYL TRANSFERASE MEASUREMENT
C0202113|T059|11274001|SNOMEDCT_US|LACTATE DEHYDROGENASE|LACTATE DEHYDROGENASE MEASUREMENT
C0523826|T059|104866001|SNOMEDCT_US|PHOSPHATE|PHOSPHATE MEASUREMENT
C0877347|T059|250707004|SNOMEDCT_US|GLOBULIN|GLOBULIN MEASUREMENT
# C0337439|T059|42950004|SNOMEDCT_US|IRON|IRON MEASUREMENT
C0201950|T059|77068002|SNOMEDCT_US|CHOLESTEROL|CHOLESTEROL MEASUREMENT
C0202236|T059|14740000|SNOMEDCT_US|TRIGLYCERIDES|TRIGLYCERIDES MEASUREMENT
C0523558|T059|313811003|SNOMEDCT_US|CHOLESTEROL/HDL RATIO SCREEN|CHOLESTEROL/HDL RATIO MEASUREMENT
C0202165|T059|81065003|SNOMEDCT_US|PH|PH MEASUREMENT
C0023516|T034|272170001|SNOMEDCT_US|WHITE COUNT|WHITE BLOOD CELL (CELL)
C1283004|T059|359846004|SNOMEDCT_US|PO2|PO2 MEASUREMENT
# C0337439|T059|42950004|SNOMEDCT_US|FE|IRON MEASUREMENT
C1277709|T059|165730006|SNOMEDCT_US|TRANSFERRIN SATURATION
C0201930|T059|38007001|SNOMEDCT_US|C02|CARBON DIOXIDE MEASUREMENT
C0030605|T059|42525009|SNOMEDCT_US|PTT|PARTIAL THROMBOPLASTIN TIME, ACTIVATED
C0036835|T034|LP32077-7|LNC|TOTAL IRON BINDING CAPACITY|IRON BINDING CAPACITY.TOTAL
C0002210|T034||LNC|ALPHA FETO PROTEIN LEVEL|ALPHA FETAL PROTEIN