C0237154|T053|160699002|SNOMEDCT_US|SHARING CONTAMINATED PERSONAL ITEMS|(HOUSING LACK) OR (HOMELESS) (FINDING)
