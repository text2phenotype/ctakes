C0015506|T037|89165002|SNOMEDCT_US|FOR HEMOPHILLIA|COAGULATION FACTOR VIII (SUBSTANCE)
C0086277|T037|44680008|SNOMEDCT_US|FACTOR VIII COAGULANT ANTIGEN|FACTOR VIII ANTIGEN (SUBSTANCE)
C0015491|T037|424562004|SNOMEDCT_US|FACTOR IX|FACTOR IX PRODUCTS
C1394921|T037||SNOMEDCT_US|COULD HAVE GOTTEN REPLACEMENT VIII
C4067217|T037||SNOMEDCT_US|ACQUIRED CLOTTING FACTOR INHIBITORS - FACTOR IX
C1394911|T037||SNOMEDCT_US|DEFICIENCY; CLOTTING FACTOR, IX (CONGENITAL) (FUNCTIONAL) (HEREDITARY) (WITH FUNCTIONAL DEFECT)
C0199967|T037|74287006|SNOMEDCT_US|TRANSFUSION OF COAGULATION FACTORS|TRANSFUSION OF COAGULATION FACTORS (PROCEDURE)
C0852255|T037||SNOMEDCT_US|BLOOD AND BLOOD PRODUCT TREATMENT
C0627512|T037||SNOMEDCT_US|CLOTTING FACTOR CONCENTRATE
C0633201|T037||SNOMEDCT_US|(DES-797-1562)-FACTOR VIII
C0633201|T037||SNOMEDCT_US|FACTOR VIII (DES-797-1562)
C0644521|T037||SNOMEDCT_US|FACTOR VIII DELTA II
C0644521|T037||SNOMEDCT_US|FACTOR VIII DELTAII
C0711027|T037||SNOMEDCT_US|KOATE-HP, HUMAN INTRAVENOUS POWDER FOR INJECTION
C0354641|T037|319871002|SNOMEDCT_US|FACTOR VIII FRACTION PRODUCTS|FACTOR VIII FRACTION PRODUCTS (SUBSTANCE)
C0354641|T037|319871002|SNOMEDCT_US|HUMAN ANTIHAEMOPHILIC FRACTION|FACTOR VIII FRACTION PRODUCTS (SUBSTANCE)
C0354641|T037|319871002|SNOMEDCT_US|HUMAN ANTIHEMOPHILIC FRACTION|FACTOR VIII FRACTION PRODUCTS (SUBSTANCE)
C0354641|T037|319871002|SNOMEDCT_US|HUMAN COAGULATION FACTOR VIII|FACTOR VIII FRACTION PRODUCTS (SUBSTANCE)
C0354641|T037|319871002|SNOMEDCT_US|FACTOR VIII FRACTION PRODUCTS |FACTOR VIII FRACTION PRODUCTS (SUBSTANCE)
C0354641|T037|319871002|SNOMEDCT_US|FACTOR VIII FRACTION PRODUCTS |FACTOR VIII FRACTION PRODUCTS (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|PORCINE FACTOR VIII|PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR, PORCINE|PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR,PORCINE|PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|PORCINE FACTOR VIII |PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|PORCINE FACTOR VIII |PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|PORCINE ANTIHAEMOPHILIC FACTOR AGENT|PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|PORCINE ANTIHAEMOPHILIC FACTOR|PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|PORCINE ANTIHEMOPHILIC FACTOR AGENT |PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|PORCINE ANTIHEMOPHILIC FACTOR AGENT|PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0724529|T037|412089003|SNOMEDCT_US|PORCINE ANTIHEMOPHILIC FACTOR|PORCINE ANTIHEMOPHILIC FACTOR AGENT (SUBSTANCE)
C0740130|T037||SNOMEDCT_US|HEMOFIL-M
C0740130|T037||SNOMEDCT_US|HEMOFIL
C0740130|T037||SNOMEDCT_US|HEMOPHIL
C0740130|T037||SNOMEDCT_US|HEMOFIL M
C0740130|T037||SNOMEDCT_US|HEMOFIL HM
C0795577|T037||SNOMEDCT_US|RECOMBINANT ANTIHEMOPHILIC FACTOR VIII
C0795577|T037||SNOMEDCT_US|FACTOR VIII RECOMBINANT
C0541364|T037||SNOMEDCT_US|FVIII ISE
C0541364|T037||SNOMEDCT_US|FACTOR VIII ISE
C0591821|T037||SNOMEDCT_US|MONOCLATE-P
C0591821|T037||SNOMEDCT_US|MONOCLATE-P (OBSOLETE)
C2342443|T037||SNOMEDCT_US|XYNTHA
C2342443|T037||SNOMEDCT_US|FACTOR VIII (XYNTHA)
C2342443|T037||SNOMEDCT_US|FACTOR VIII (XYNTHA) 
C0015514|T037|65738000|SNOMEDCT_US| I DON'T THINK ACTIVATED VIII IS GIVEN IN HEMOPHLIA, BUT I'M NOT CONFIDENT ENOUGH TO EXCLUDE AND WOULD BE SURPRISD IF YOU GOT FALSE POSITIVES|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|FACTOR VIII, THROMBIN ACTIVATED|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|FACTOR VIIIA|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|THROMBIN-ACTIVATED FACTOR VIII|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|BLOOD-COAGULATION FACTOR VIIIA, PROCOAGULANT|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|FACTOR VIIIA, COAGULATION|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|VIIIA, COAGULATION FACTOR|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|COAG FACTOR VIIIA|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|BLOOD COAG FACTOR VIII ACTIVATED|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|FACTOR VIIIA [CHEMICAL/INGREDIENT]|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|COAGULATION FACTOR VIIIA|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|FACTOR VIII, THROMBIN-ACTIVATED|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|FACTOR VIII, ACTIVATED|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|BLOOD COAGULATION FACTOR VIII, ACTIVATED|COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015514|T037|65738000|SNOMEDCT_US|COAGULATION FACTOR VIIIA |COAGULATION FACTOR VIIIA (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|FACTOR VIII|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|COAGULATION FACTOR VIII|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|BLOOD-COAGULATION FACTOR VIII, COMPLEX|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|COAG FACTOR VIII|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|BLOOD COAG FACTOR VIII|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR A|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|THROMBOPLASTINOGEN A|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|PLATELET COFACTOR I|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|HEMATOLOGICAL AGENTS ANTIHEMOPHILIC FACTORS|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|ANTIHEMOPHILIC FACTORS|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|ANTIHEMOPHILIC FACTORS |COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|THROMBOPLASTINOGEN|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|BLOOD COAGULATION FACTOR VIII|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|FACTOR VIII [CHEMICAL/INGREDIENT]|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|COAGULATION FACTOR VIII |COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|FACTOR VIII (ANTIHEMOPHILIC FACTOR, HUMAN) PER I.U.|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|AHF|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|AHG|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|ANTIHEMOPHILIC GLOBULIN|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|FACTOR VIII |COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR A|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|ANTIHAEMOPHILIC GLOBULIN|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|COAGULATION FACTOR VIII  [AMBIGUOUS]|COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|FACTOR VIII PRODUCT |COAGULATION FACTOR VIII (SUBSTANCE)
C0015506|T037|89165002|SNOMEDCT_US|FACTOR VIII PRODUCT|COAGULATION FACTOR VIII (SUBSTANCE)
C0020199|T037||SNOMEDCT_US|HYATE C
C0020199|T037||SNOMEDCT_US|HYATT C
C0020199|T037||SNOMEDCT_US|HYATE:C
C0020199|T037||SNOMEDCT_US|HYATE C (OBSOLETE)
C0020199|T037||SNOMEDCT_US|HYATEC
C0020199|T037||SNOMEDCT_US|HYATTC
C0020199|T037||SNOMEDCT_US|HYATE-C
C0020199|T037||SNOMEDCT_US|HYATT-C
C0020199|T037||SNOMEDCT_US|SPEYWOOD BRAND OF PORCINE FACTOR VIII PREPARATION
C2825466|T037||SNOMEDCT_US|MOROCTOCOG ALFA 
C2825466|T037||SNOMEDCT_US|MOROCTOCOG ALFA
C2825466|T037||SNOMEDCT_US|MOROCTOCOG ALFA 
C2825466|T037||SNOMEDCT_US|ANTIHEMOPHILIC FACTOR, HUMAN RECOMBINANT RESIDUES 743-1636 DELETED
C0971600|T037||SNOMEDCT_US|REFACTO
C0971600|T037||SNOMEDCT_US|REFACTO 
C0218184|T037||SNOMEDCT_US|KOGENATE
C0218184|T037||SNOMEDCT_US|KOGENATE BAYER
C0218184|T037||SNOMEDCT_US|KOGENATE (OBSOLETE)
C0218184|T037||SNOMEDCT_US|FACTOR VIII (KOGENATE)
C0218184|T037||SNOMEDCT_US|FACTOR VIII (KOGENATE) 
C0218184|T037||SNOMEDCT_US|RECOMBINANT ANTIHEMOPHILIC FACTOR VIII
C0700346|T037||SNOMEDCT_US|ANTIHEMOPHILIC FACTOR, HUMAN
C0700346|T037||SNOMEDCT_US|ANTIHEMOPHILIC FACTOR HUMAN
C0700346|T037||SNOMEDCT_US|ANTIHEMOPHILIC FACTOR,HUMAN
C2927721|T037||SNOMEDCT_US|FACTOR VIII/VON WILLEBRAND FACTOR COMPLEX HUMAN PLASMA
C2732002|T037|409259007|SNOMEDCT_US|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|RECOMBINANT ANTIHAEMOPHILIC FACTOR AGENT|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR, RECOMBINANT|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR, HUMAN RECOMBINANT|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|FVIII|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|FACTOR VIII|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR,RECOMBINANT|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|RECOMBINANT HUMAN FACTOR VIII - OCTOCOG ALPHA|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|DNA FACTOR VIII |RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|OCTOCOG ALPHA|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|RECOMBINANT ANTIHAEMOPHILIC FACTOR PREPARATION|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT |RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|RECOMBINANT ANTIHEMOPHILIC FACTOR PREPARATION|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|DNA FACTOR VIII |RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|RECOMBINANT ANTIHEMOPHILIC FACTOR PREPARATION |RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT |RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2732002|T037|409259007|SNOMEDCT_US|RECOMBINANT HUMAN FACTOR VIII|RECOMBINANT ANTIHEMOPHILIC FACTOR AGENT (PRODUCT)
C2601455|T037||SNOMEDCT_US|COAGULATION FACTOR VIII &#X7C; PLATELET POOR PLASMA
C2968287|T037||SNOMEDCT_US|FACTOR VIII &#X7C; PATIENT
C1985551|T037||SNOMEDCT_US|COAGULATION FACTOR VIII ACTIVITY.XA ACTIVATOR &#X7C; PLATELET POOR PLASMA
C1976512|T037||SNOMEDCT_US|TRANSFUSE FACTOR VIII &#X7C; PATIENT
C2968288|T037||SNOMEDCT_US|FACTOR VIII UNITS &#X7C; BLOOD PRODUCT UNIT
C1985549|T037||SNOMEDCT_US|COAGULATION FACTOR VIII AB &#X7C; PLATELET POOR PLASMA
C1985548|T037||SNOMEDCT_US|COAGULATION FACTOR VIII &#X7C; XXX
C2601456|T037||SNOMEDCT_US|COAGULATION FACTOR VIII ACTIVITY &#X7C; PLATELET POOR PLASMA
C1985550|T037||SNOMEDCT_US|COAGULATION FACTOR VIII ACTIVATED &#X7C; PLATELET POOR PLASMA
C2359705|T037||SNOMEDCT_US|TRANSFUSE FACTOR VIII &#X7C; BLOOD PRODUCT UNIT
C1307126|T037||SNOMEDCT_US|ANTIHEMOPHILIC FACTOR
C1307126|T037||SNOMEDCT_US|FACTOR VIII, HUMAN
C1307126|T037||SNOMEDCT_US|MOST ACCEPTED ABBREV IS FOR ANTIHEMOPHILIC FACTOR, PEOPLE MIGHT USE IN OTHER WAYS (ACUTE HEART FAILURE) BUT RARE
C1307126|T037||SNOMEDCT_US|F8 PROTEIN, HUMAN
C1307126|T037||SNOMEDCT_US|FVIII PROTEIN, HUMAN
C1307126|T037||SNOMEDCT_US|COAGULATION FACTOR VIII, PROCOAGULANT COMPONENT (HEMOPHILIA A) PROTEIN, HUMAN
C1307126|T037||SNOMEDCT_US|FACTOR VIII
C1307126|T037||SNOMEDCT_US|COAGULATION FACTOR VIII
C1307126|T037||SNOMEDCT_US|COAGULATION FACTOR VIIIC
C1307126|T037||SNOMEDCT_US|F8
C1307126|T037||SNOMEDCT_US|FACTOR VIII F8B
C1307126|T037||SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR
C1307126|T037||SNOMEDCT_US|PROCOAGULANT COMPONENT
C0086428|T037||SNOMEDCT_US|HUMATE-P
C0086428|T037||SNOMEDCT_US|HUMATE-P (OBSOLETE)
C2726511|T037||SNOMEDCT_US|FOR VWF DEFICENCY
C0594139|T037||SNOMEDCT_US|ALPHANATE
C0594139|T037||SNOMEDCT_US|ALPHANATE (OBSOLETE)
C3660038|T037||SNOMEDCT_US|N8-GP COMPOUND
C3529561|T037||SNOMEDCT_US|N8 RFVIII
C3529561|T037||SNOMEDCT_US|N8 RECOMBINANT FACTOR VIII
C3529561|T037||SNOMEDCT_US|RECOMBINANT FACTOR VIII N8
C1815380|T037||SNOMEDCT_US|OPTIVATE
C3849397|T037||SNOMEDCT_US|FACTOR VIII-FC FUSION PROTEIN
C3849397|T037||SNOMEDCT_US|RFVIIIFC PROTEIN
C3859470|T037||SNOMEDCT_US|OBIZUR
C3859426|T037|725746009|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR, PORCINE B-DOMAIN TRUNCATED RECOMBINANT|SUSOCTOCOG ALFA (SUBSTANCE)
C3859426|T037|725746009|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR PORCINE, B-DOMAIN TRUNCATED RECOMBINANT|SUSOCTOCOG ALFA (SUBSTANCE)
C4018188|T037||SNOMEDCT_US|NOVOEIGHT
C4031949|T037||SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (RECOMBINANT), PORCINE SEQUENCE 
C4031949|T037||SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (RECOMBINANT), PORCINE SEQUENCE
C3834170|T037|718943005|SNOMEDCT_US|FACTOR VIII (B-DOMAIN DELETED RECOMBINANT) FC FUSION PROTEIN|EFMOROCTOCOG ALFA (SUBSTANCE)
C3834170|T037|718943005|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR, RECOMBINANT FC FUSION PROTEIN|EFMOROCTOCOG ALFA (SUBSTANCE)
C3834170|T037|718943005|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (RECOMBINANT), FC FUSION PROTEIN |EFMOROCTOCOG ALFA (SUBSTANCE)
C3834170|T037|718943005|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (RECOMBINANT), FC FUSION PROTEIN|EFMOROCTOCOG ALFA (SUBSTANCE)
C3834170|T037|718943005|SNOMEDCT_US|EFMOROCTOCOG ALFA|EFMOROCTOCOG ALFA (SUBSTANCE)
C4038482|T037||SNOMEDCT_US|FACTOR VIII+VON WILLEBRAND FACTOR.RISTOCETIN COFACTOR
C4045418|T037||SNOMEDCT_US|BAY 94-9027
C4057564|T037||SNOMEDCT_US|KOATE
C0376176|T037||SNOMEDCT_US|MONOCLATE
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ 1000 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ 220-400 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ 250 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ 401-800 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ 500 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ KIT 250 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ KIT 500 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR HUMAN INTRAVENOUS POWDER FOR INJECTION|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (OBSOLETE) HUMAN INTRAVENOUS POWDER FOR INJECTION|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR AGENT 500 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT |ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR AGENT 1500 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT |ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR AGENT 500 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR AGENT 500 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR AGENT 1500 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT |ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR AGENT 1500 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII HUMAN 1 IU INTRAVENOUS POWDER FOR SOLUTION|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR,HUMAN INJ|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR,HUMAN INJ [VA PRODUCT]|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII HUMAN 1 IU INJECTION POWDER FOR SOLUTION|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII HUMAN INTRAVENOUS POWDER FOR SOLUTION|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII HUMAN 1 IU INJECTION POWDER FOR SOLUTION [FACTOR VIII:C]|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ 801-1500 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ 1501-2000 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII HUMAN/ANTIHEMOPHILIC FACTOR VIII:C HUMAN 1 IU-1 IU INTRAVENOUS POWDER FOR SOLUTION|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (HUMAN) FOR INJ 1700 UNIT|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|FACTOR VIII, HUMAN 1 UNT INJECTION|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR, HUMAN 1 UNT INJECTION|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR 500UNT/VIAL POWDER|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR 500UNT/VIAL POWDER |ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR 500UNT/VIAL POWDER|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C1300015|T037|427242002|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII:C HUMAN 1 IU INTRAVENOUS POWDER FOR SOLUTION|ANTIHEMOPHILIC FACTOR AGENT 1000 IU POWDER FOR INJECTION SOLUTION 5ML VIAL + DILUENT (PRODUCT)
C0543246|T037|347623003|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR (OBSOLETE) PORCINE INTRAVENOUS POWDER FOR INJECTION|PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR PORCINE INTRAVENOUS POWDER FOR INJECTION|PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|PORCINE FACTOR VIII 700IU INJECTION|PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII:C (PORCINE) 1 U INJECTION POWDER FOR SOLUTION|PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII (PORCINE) INJECTION POWDER FOR SOLUTION|PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII (PORCINE) 1 IU INJECTION POWDER FOR SOLUTION|PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR VIII (PORCINE) 1 U INTRAVENOUS POWDER FOR SOLUTION|PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|PORCINE FACTOR VIII 700IU POWDER FOR INJECTION SOLUTION VIAL |PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|PORCINE FACTOR VIII 700IU POWDER FOR INJECTION SOLUTION VIAL|PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|PORCINE FACTOR VIII 700IU INJECTION |PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C0543246|T037|347623003|SNOMEDCT_US|PORCINE FACTOR VIII 700IU INJECTION |PORCINE FACTOR VIII 700IU INJECTION (SUBSTANCE)
C4064080|T037|718853005|SNOMEDCT_US|SIMOCTOCOG ALFA|SIMOCTOCOG ALFA (SUBSTANCE)
C4064080|T037|718853005|SNOMEDCT_US|SIMOCTOCOG ALFA |SIMOCTOCOG ALFA (SUBSTANCE)
C4064080|T037|718853005|SNOMEDCT_US|ANTIHEMOPHILIC FACTORS SIMOCTOCOG ALFA|SIMOCTOCOG ALFA (SUBSTANCE)
C4064080|T037|718853005|SNOMEDCT_US|COAGULATION FACTOR VIII, B-DOMAIN DELETED RECOMBINANT|SIMOCTOCOG ALFA (SUBSTANCE)
C4074414|T037||SNOMEDCT_US|NUWIQ
C3529563|T037|735055007|SNOMEDCT_US|TUROCTOCOG ALFA|TUROCTOCOG ALFA (SUBSTANCE)
C3529563|T037|735055007|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR, HUMAN B-DOMAIN TRUNCATED RECOMBINANT|TUROCTOCOG ALFA (SUBSTANCE)
C0732093|T037|319925005|SNOMEDCT_US|FACTOR VIII + VON WILLEBRAND FACTOR|FACTOR VIII+VON WILLEBRAND FACTOR (SUBSTANCE)
C0732093|T037|319925005|SNOMEDCT_US|FACTOR VIII, VON WILLEBRAND FACTOR DRUG COMBINATION|FACTOR VIII+VON WILLEBRAND FACTOR (SUBSTANCE)
C0732093|T037|319925005|SNOMEDCT_US|FACTOR VIII - VON WILLEBRAND FACTOR|FACTOR VIII+VON WILLEBRAND FACTOR (SUBSTANCE)
C0732093|T037|319925005|SNOMEDCT_US|FACTOR VIII / VON WILLEBRAND FACTOR|FACTOR VIII+VON WILLEBRAND FACTOR (SUBSTANCE)
C0732093|T037|319925005|SNOMEDCT_US|FACTOR VIII+VON WILLEBRAND FACTOR|FACTOR VIII+VON WILLEBRAND FACTOR (SUBSTANCE)
C0732093|T037|319925005|SNOMEDCT_US|FACTOR VIII+VON WILLEBRAND FACTOR |FACTOR VIII+VON WILLEBRAND FACTOR (SUBSTANCE)
C0732093|T037|319925005|SNOMEDCT_US|FACTOR VIII+VON WILLEBRAND FACTOR |FACTOR VIII+VON WILLEBRAND FACTOR (SUBSTANCE)
C0358606|T037|346435001|SNOMEDCT_US|ACTIVATED PROTHROMBIN COMPLEX CONCENTRATE|FACTOR VIII BY-PASSING FRACTION PRODUCTS (SUBSTANCE)
C0358606|T037|346435001|SNOMEDCT_US|FACTOR VIII BY-PASSING FRACTION PRODUCTS|FACTOR VIII BY-PASSING FRACTION PRODUCTS (SUBSTANCE)
C0358606|T037|346435001|SNOMEDCT_US|FACTOR VIII BY-PASSING FRACTION PRODUCTS |FACTOR VIII BY-PASSING FRACTION PRODUCTS (SUBSTANCE)
C0358606|T037|346435001|SNOMEDCT_US|FACTOR VIII BY-PASSING FRACTION PRODUCTS |FACTOR VIII BY-PASSING FRACTION PRODUCTS (SUBSTANCE)
C0720828|T037||SNOMEDCT_US|HELIXATE
C0720828|T037||SNOMEDCT_US|HELIXATE (OBSOLETE)
C1815247|T037||SNOMEDCT_US|MONARC-M
C1815247|T037||SNOMEDCT_US|MONARC-M (OBSOLETE)
C0218182|T037||SNOMEDCT_US|RECOMBINATE
C0218182|T037||SNOMEDCT_US|RECOMBINATE (OBSOLETE)
C1691209|T037|422675008|SNOMEDCT_US|OCTOCOG ALFA|OCTOCOG ALFA (PRODUCT)
C1691209|T037|422675008|SNOMEDCT_US|OCTOCOG ALFA |OCTOCOG ALFA (PRODUCT)
C1691209|T037|422675008|SNOMEDCT_US|DNA FACTOR VIII|OCTOCOG ALFA (PRODUCT)
C1691209|T037|422675008|SNOMEDCT_US|DEOXYRIBONUCLEIC ACID FACTOR VIII|OCTOCOG ALFA (PRODUCT)
C1691209|T037|422675008|SNOMEDCT_US|DEOXYRIBONUCLEIC ACID FACTOR VIII |OCTOCOG ALFA (PRODUCT)
C1691209|T037|422675008|SNOMEDCT_US|OCTOCOG ALFA |OCTOCOG ALFA (PRODUCT)
C0056540|T037||SNOMEDCT_US|CRYOBULIN
C0056545|T037||SNOMEDCT_US|CRYOPRECIPITATE COAGULUM
C0961271|T037||SNOMEDCT_US|BAY 14-2222
C0961271|T037||SNOMEDCT_US|BAY-14-2222
C0961271|T037||SNOMEDCT_US|BAY14-2222
C0966326|T037||SNOMEDCT_US|MALMO PROTOCOL
C0966500|T037|441943001|SNOMEDCT_US|R-VIII SQ|MOROCTOCOG ALFA (PRODUCT)
C0966500|T037|441943001|SNOMEDCT_US|RECOMBINANT FACTOR VIII SQ|MOROCTOCOG ALFA (PRODUCT)
C1098523|T037||SNOMEDCT_US|RFVIII-FS
C1098523|T037||SNOMEDCT_US|RECOMBINANT FVIII, SUGAR FORMULATED
C1121470|T037||SNOMEDCT_US|B-DOMAIN-DELETED FACTOR VIII
C1121470|T037||SNOMEDCT_US|GC-RAHF
C1121470|T037||SNOMEDCT_US|RFVIII (B-DOMAIN-DELETED)
C1175691|T037||SNOMEDCT_US|8Y FACTOR VIII-VON WILLEBRAND FACTOR CONCENTRATE
C1175691|T037||SNOMEDCT_US|FACTOR VIII-VON WILLEBRAND FACTOR CONCENTRATE 8Y
C1175691|T037||SNOMEDCT_US|VWF-FVLLI 8Y
C0731320|T037||SNOMEDCT_US|HAEMATE P
C2002589|T037||SNOMEDCT_US|IMMUNATE SOLVENT DETERGENT, HUMAN
C1815260|T037||SNOMEDCT_US|ADVATE
C0015494|T037|63856005|SNOMEDCT_US|ACTIVATED FACTOR IX|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|FACTOR IXA|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|FACTOR IXA, COAGULATION|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|IXA, COAGULATION FACTOR|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|BLOOD COAG FACTOR IX ACTIVATED|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|COAG FACTOR IXA|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|FACTOR VIIIIA|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|FACTOR VIIII ACTIVATED|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|COAGULATION FACTOR VIIIIA|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|COAGULATION FACTOR IXA -RETIRED-|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|COAGULATION FACTOR IXA|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|FACTOR IX, ACTIVATED|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|BLOOD COAGULATION FACTOR IX, ACTIVATED|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|FACTOR IXA [CHEMICAL/INGREDIENT]|COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|COAGULATION FACTOR IXA |COAGULATION FACTOR IXA (SUBSTANCE)
C0015494|T037|63856005|SNOMEDCT_US|ACTIVATED CHRISTMAS FACTOR|COAGULATION FACTOR IXA (SUBSTANCE)
C0015491|T037|424562004|SNOMEDCT_US|FACTOR IX|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|CHRISTMAS FACTOR|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|COAGULATION FACTOR IX|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|BLOOD-COAGULATION FACTOR IX|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|COMPLEX, FACTOR IX|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|FRACTION, FACTOR IX|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|IX COMPLEX, FACTOR|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|IX FRACTION, FACTOR|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|FACTOR IX, COAGULATION|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|IX, COAGULATION FACTOR|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|COAGULATION FACTOR VIIII|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|COAG FACTOR IX|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|FACTOR VIIII|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|BLOOD COAG FACTOR IX|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR B|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|AUTOPROTHROMBIN II|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|THROMBOPLASTINOGEN B|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|FACTOR IX COMPLEX|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|PLASMA THROMBOPLASTIN COMPONENT|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|FACTOR IX FRACTION|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|BLOOD COAGULATION FACTOR IX|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|FACTOR IX [CHEMICAL/INGREDIENT]|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|PLATELET COFACTOR II|FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|COAGULATION FACTOR IX |FACTOR IX PRODUCTS
C0015491|T037|424562004|SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR B|FACTOR IX PRODUCTS
C1170091|T037||SNOMEDCT_US|BENEFIX
C1170091|T037||SNOMEDCT_US|BENEFIX (OBSOLETE)
C0060018|T037||SNOMEDCT_US|FACTOR IX LONG BEACH
C0060018|T037||SNOMEDCT_US|FIX-LB
C0082540|T037||SNOMEDCT_US|FACTOR IX-ANTITHROMBIN III COMPLEX
C0082540|T037||SNOMEDCT_US|FACTOR IX-ATIII COMPLEX
C0082536|T037||SNOMEDCT_US|FACTOR IX LEYDEN
C0082536|T037||SNOMEDCT_US|LEYDEN FACTOR IX
C0060011|T037||SNOMEDCT_US|BM LAKE ELSINORE FACTOR IX
C0060011|T037||SNOMEDCT_US|FACTOR IX BM LAKE ELSINORE
C0060011|T037||SNOMEDCT_US|FACTOR IX BMLE
C0060014|T037||SNOMEDCT_US|BLOOD-COAGULATION FACTOR IX CHAPEL HILL
C0060014|T037||SNOMEDCT_US|FACTOR IX CHAPEL HILL
C0297142|T037||SNOMEDCT_US|MONONINE
C0297142|T037||SNOMEDCT_US|MONONINE (OBSOLETE)
C0297142|T037||SNOMEDCT_US|MONONINE (OBSOLETE1)
C0289773|T037||SNOMEDCT_US|FACTOR IX (1-47)
C0251224|T037||SNOMEDCT_US|FACTOR IX STRASBOURG 2
C0117201|T037||SNOMEDCT_US|FACTOR IX MADRID
C0060013|T037||SNOMEDCT_US|FACTOR IX CARDIFF
C0117199|T037||SNOMEDCT_US|FACTOR IX CAMBRIDGE
C0117199|T037||SNOMEDCT_US|FACTOR IX PROPEPTIDE
C0718844|T037||SNOMEDCT_US|BEBULIN VH
C0718844|T037||SNOMEDCT_US|BEBULIN VH (OBSOLETE)
C0592047|T037||SNOMEDCT_US|REPLENINE
C2826076|T037|425189006|SNOMEDCT_US|FACTOR IX, RECOMBINANT|NONACOG ALFA (SUBSTANCE)
C2826076|T037|425189006|SNOMEDCT_US|COAGULATION FACTOR IX RECOMBINANT HUMAN|NONACOG ALFA (SUBSTANCE)
C2826076|T037|425189006|SNOMEDCT_US|FACTOR IX,RECOMBINANT|NONACOG ALFA (SUBSTANCE)
C2826076|T037|425189006|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMBINANT HUMAN)|NONACOG ALFA (SUBSTANCE)
C3666839|T037||SNOMEDCT_US|RIXUBIS
C3644708|T037||SNOMEDCT_US|KCENTRA
C0718417|T037||SNOMEDCT_US|ALPHANINE SD
C0718417|T037||SNOMEDCT_US|ALPHANINE SD (OBSOLETE)
C0718417|T037||SNOMEDCT_US|ALPHANINE SD (OBSOLETE1)
C2972532|T037||SNOMEDCT_US|TRANSFUSE FACTOR IX &#X7C; PATIENT
C1985535|T037||SNOMEDCT_US|COAGULATION FACTOR IX ACTIVATED &#X7C; PLATELET POOR PLASMA
C2601448|T037||SNOMEDCT_US|COAGULATION FACTOR IX &#X7C; PLATELET POOR PLASMA
C2972533|T037||SNOMEDCT_US|TRANSFUSE FACTOR IX UNITS &#X7C; BLOOD PRODUCT UNIT
C1985536|T037||SNOMEDCT_US|COAGULATION FACTOR IX AG &#X7C; PLATELET POOR PLASMA
C2601449|T037||SNOMEDCT_US|COAGULATION FACTOR IX ACTIVITY &#X7C; PLATELET POOR PLASMA
C2968286|T037||SNOMEDCT_US|FACTOR IX &#X7C; PATIENT
C2749016|T037||SNOMEDCT_US|THROMBOPHILIA, X-LINKED, DUE TO FACTOR IX DEFECT
C2749016|T037||SNOMEDCT_US|THPH8
C3657751|T037||SNOMEDCT_US|IB1001
C3657751|T037||SNOMEDCT_US|IB1001 TRENACOG ALFA
C4048712|T037|54144004|SNOMEDCT_US|FACTOR IX COMPLEX|FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|COAGULATION FACTOR IX|FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|FACTOR IX COMPLEX AGENT|FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|FACTOR IX COMPLEX, HUMAN|FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|FACTOR IX COMPLEX,HUMAN|FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|COAGULATION FACTOR IX COMPLEX HUMAN|FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|FACTOR IX COMPLEX PREPARATION|FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|FACTOR IX PREPARATION|FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|FACTOR IX COMPLEX AGENT |FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|FACTOR IX AGENT|FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C4048712|T037|54144004|SNOMEDCT_US|FACTOR IX COMPLEX PREPARATION |FACTOR IX COMPLEX PREPARATION (SUBSTANCE)
C3883805|T037|735232002|SNOMEDCT_US|N9-GP COMPOUND|NONACOG BETA PEGOL (SUBSTANCE)
C3883805|T037|735232002|SNOMEDCT_US|NONACOG BETA PEGOL|NONACOG BETA PEGOL (SUBSTANCE)
C3883952|T037||SNOMEDCT_US|FACTOR IX PADUA
C3883952|T037||SNOMEDCT_US|FACTOR IX-PADUA
C0722828|T037||SNOMEDCT_US|PROFILNINE SD
C4041753|T037||SNOMEDCT_US|RFIXFC PROTEIN
C4041753|T037||SNOMEDCT_US|FACTOR IX FC FUSION PROTEIN
C4051373|T037||SNOMEDCT_US|IXINITY
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMBINANT) FOR INJ 1000 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMBINANT) FOR INJ 250 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMBINANT) FOR INJ 500 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX RECOMBINANT INTRAVENOUS POWDER FOR INJECTION|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMBINANT) FOR INJ 2000 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT 1000 UNT/VIL INJ|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT 1000 UNT/VIL INJ [VA PRODUCT]|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX RECOMBINANT 1 IU INTRAVENOUS POWDER FOR SOLUTION|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX RECOMBINANT POWDER FOR SOLUTION FOR INJECTI WITH ALCOHOL PAD OR SWAB - IV ADMINISTRATION SET (UNSPECIFIED) - FILTER SPIKE - DOUBLE-ENDED NEEDLE - STERILE WATER FOR INJECTION -|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMBINANT) FOR INJ 3000 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT 3000 UNIT/VIL INJ|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT 2000 UNIT/VIL INJ|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT 2000 UNIT/VIL INJ [VA PRODUCT]|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT 3000 UNIT/VIL INJ [VA PRODUCT]|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMB) (RFIXFC) FOR INJ 500 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMB) (RFIXFC) FOR INJ 2000 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX RECOMBINANT LYOPHILISATE FOR SOLUTION FOR INJECTI WITH VIAL ADAPTER - DILUENT -|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMB) (RFIXFC) FOR INJ 1000 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMB) (RFIXFC) FOR INJ 3000 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMBINANT) FOR INJ 1500 UNIT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT (THR148) 1500 UNIT/VIL INJ [VA PRODUCT]|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT (THR148) 1000 UNIT/VIL INJ|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT (THR148) 500 UNIT/VIL INJ|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOM(THR148) 1000UNIT/VIL INJ|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOM(THR148) 1500UNIT/VIL INJ|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOM(THR148) 500UNIT/VIL INJ|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT (THR148) 1500 UNIT/VIL INJ|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT (THR148) 500 UNIT/VIL INJ [VA PRODUCT]|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|FACTOR IX,RECOMBINANT (THR148) 1000 UNIT/VIL INJ [VA PRODUCT]|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|COAGULATION FACTOR IX (RECOMBINANT HUMAN) 1 UNT INJECTION|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 1000IU INJECTION (PDR FOR RECON)+SOLVENT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 1000IU POWDER AND SOLVENT FOR INJECTION SOLUTION VIAL |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 1000IU POWDER AND SOLVENT FOR INJECTION SOLUTION VIAL|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 250IU INJECTION (PDR FOR RECON)+SOLVENT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 250IU POWDER AND SOLVENT FOR INJECTION SOLUTION VIAL |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 250IU POWDER AND SOLVENT FOR INJECTION SOLUTION VIAL|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 500IU INJECTION (PDR FOR RECON)+SOLVENT|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER AND SOLVENT FOR INJECTION SOLUTION VIAL |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER AND SOLVENT FOR INJECTION SOLUTION VIAL|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 1000IU INJECTION (PDR FOR RECON)+SOLVENT |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 1000IU INJECTION (PDR FOR RECON)+SOLVENT |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 250IU INJECTION (PDR FOR RECON)+SOLVENT |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 250IU INJECTION (PDR FOR RECON)+SOLVENT |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 500IU INJECTION (PDR FOR RECON)+SOLVENT |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 500IU INJECTION (PDR FOR RECON)+SOLVENT |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 1000IU POWDER FOR INJECTION SOLUTION VIAL |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 1000IU POWDER FOR INJECTION SOLUTION VIAL|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 250IU POWDER FOR INJECTION SOLUTION VIAL |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 250IU POWDER FOR INJECTION SOLUTION VIAL|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL |RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C1269927|T037|415244004|SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL|RECOMBINANT COAGULATION FACTOR IX 500IU POWDER FOR INJECTION SOLUTION VIAL
C0724584|T037||SNOMEDCT_US|FACTOR IX (HUMAN)
C0724584|T037||SNOMEDCT_US|COAGULATION FACTOR IX HUMAN
C0724584|T037||SNOMEDCT_US|FACTOR IX, HUMAN
C0724584|T037||SNOMEDCT_US|FACTOR 9
C0724584|T037||SNOMEDCT_US|PLASMA THROMBOPLASTIC COMPONENT
C0724584|T037||SNOMEDCT_US|PLASMA THROMBOPLASTIN COMPONENT
C0724584|T037||SNOMEDCT_US|COAGULATION FACTOR IX, HUMAN
C0724584|T037||SNOMEDCT_US|CHRISTMAS FACTOR
C0724584|T037||SNOMEDCT_US|FACTOR IX
C0724584|T037||SNOMEDCT_US|COAGULATION FACTOR IX
C0724584|T037||SNOMEDCT_US|EC 3.4.21.22
C0313501|T037|45807004|SNOMEDCT_US|COAGULATION FACTOR IX VARIANT |COAGULATION FACTOR IX VARIANT (SUBSTANCE)
C0313501|T037|45807004|SNOMEDCT_US|COAGULATION FACTOR IX VARIANT|COAGULATION FACTOR IX VARIANT (SUBSTANCE)
C0313501|T037|45807004|SNOMEDCT_US|COAGULATION FACTOR IX VARIANT, NOS|COAGULATION FACTOR IX VARIANT (SUBSTANCE)
C1273037|T037||SNOMEDCT_US|NONACOG ALFA
C1273037|T037||SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX
C1273037|T037||SNOMEDCT_US|COAGULATION FACTOR IX RECOMBINANT
C1273037|T037||SNOMEDCT_US|NONACOG ALFA 
C1273037|T037||SNOMEDCT_US|NONACOG ALFA 
C1273037|T037||SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX 
C1273037|T037||SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX PREPARATION 
C1273037|T037||SNOMEDCT_US|RECOMBINANT COAGULATION FACTOR IX PREPARATION
C1815181|T037||SNOMEDCT_US|KONYNE 80
C1815181|T037||SNOMEDCT_US|KONYNE 80 (OBSOLETE)
C0631906|T037||SNOMEDCT_US|FACTOR IX SEATTLE(2)
C0631906|T037||SNOMEDCT_US|FACTOR IX SEATTLE2
C0633767|T037||SNOMEDCT_US|FACTOR IX GLA-PEPTIDE
C0636372|T037||SNOMEDCT_US|FACTOR IX VANCOUVER
C0636589|T037||SNOMEDCT_US|FACTOR IX NIIGATA
C0636589|T037||SNOMEDCT_US|BLOOD COAGULATION FACTOR IX NIIGATA
C0636589|T037||SNOMEDCT_US|NIIGATA FACTOR IX
C0637620|T037||SNOMEDCT_US|FACTOR IX SAN DIMAS
C0637620|T037||SNOMEDCT_US|SAN DIMAS FACTOR IX
C0638162|T037||SNOMEDCT_US|FACTOR IX TROED-Y-RHIW
C0638164|T037||SNOMEDCT_US|FACTOR IX KAWACHINAGANO
C0638164|T037||SNOMEDCT_US|FACTOR IX KWC
C0639016|T037||SNOMEDCT_US|FACTOR IX BM NAGOYA
C0639016|T037||SNOMEDCT_US|IX NAGOYA
C0640832|T037||SNOMEDCT_US|FACTOR IX CHONGQING
C0641637|T037||SNOMEDCT_US|FACTOR IX ALABAMA
C0641676|T037||SNOMEDCT_US|FACTOR IX DEVENTER
C0641677|T037||SNOMEDCT_US|FACTOR IX BERGAMO
C0641681|T037||SNOMEDCT_US|FACTOR IX NOVARA
C0641682|T037||SNOMEDCT_US|FACTOR IX MILANO
C0643142|T037||SNOMEDCT_US|FACTOR IX HOLLYWOOD
C0643142|T037||SNOMEDCT_US|FACTOR IX (HW)
C0644057|T037||SNOMEDCT_US|FACTOR IX LINCOLN PARK
C0645143|T037||SNOMEDCT_US|FACTOR IX BASEL
C0645333|T037||SNOMEDCT_US|FACTOR IX NAGOYA 3
C0660527|T037||SNOMEDCT_US|FACTOR IX BM HILO
C0661606|T037||SNOMEDCT_US|PRECONATIV
C0383958|T037||SNOMEDCT_US|FACTOR IX ZUTPHEN
C1121564|T037||SNOMEDCT_US|FACTOR IX DENVER
C2743140|T037||SNOMEDCT_US|FACTOR IX, FACTOR VII, FACTOR X, PROTHROMBIN DRUG COMBINATION
C1394921|T037||SNOMEDCT_US|CLOTTING FACTOR; DEFICIENCY, VIII, WITH VASCULAR DEFECT
C1394921|T037||SNOMEDCT_US|DEFICIENCY; CLOTTING FACTOR, VIII, WITH VASCULAR DEFECT
C0200408|T037|165579001|SNOMEDCT_US|FACTOR IX ASSAY|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|FACTOR IX ASSAY |FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|FACTOR IX LEVEL|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|COAGULATION FACTOR IX LEVEL|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|CLOTTING; FACTOR IX (PTC OR CHRISTMAS)|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|COAGULATION FACTOR IX MEASUREMENT|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|CLOTTING FACTOR IX PTC/CHRISTMAS|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|FACTOR IX MEASUREMENT|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|CLOT FACTOR IX PTC/CHRSTMAS|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|ASSAY FOR CLOTTING FACTOR IX (PTC)|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|CLOTTING FACTOR IX (PTC OR CHRISTMAS) MEASUREMENT|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|FACTOR IX ASSAY |FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|CHRISTMAS FACTOR|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|FACTOR IX|FACTOR IX ASSAY (PROCEDURE)
C0200408|T037|165579001|SNOMEDCT_US|FACTIX|FACTOR IX ASSAY (PROCEDURE)
C1394911|T037||SNOMEDCT_US|CLOTTING FACTOR; DEFICIENCY, IX (CONGENITAL) (FUNCTIONAL) (HEREDITARY) (WITH FUNCTIONAL DEFECT)
C1394911|T037||SNOMEDCT_US|DEFICIENCY; CLOTTING FACTOR, IX (CONGENITAL) (FUNCTIONAL) (HEREDITARY) (WITH FUNCTIONAL DEFECT)
C0199967|T037|74287006|SNOMEDCT_US|CLOTTING FACTOR TRANSFUSION|TRANSFUSION OF COAGULATION FACTORS (PROCEDURE)
C0199967|T037|74287006|SNOMEDCT_US|COAG FACTOR TRANSFUSION|TRANSFUSION OF COAGULATION FACTORS (PROCEDURE)
C0199967|T037|74287006|SNOMEDCT_US|TRANSFUSION OF COAGULATION FACTORS|TRANSFUSION OF COAGULATION FACTORS (PROCEDURE)
C0199967|T037|74287006|SNOMEDCT_US|TRANSFUSION OF COAGULATION FACTOR|TRANSFUSION OF COAGULATION FACTORS (PROCEDURE)
C0199967|T037|74287006|SNOMEDCT_US|TRANSFUSION OF COAGULATION FACTORS |TRANSFUSION OF COAGULATION FACTORS (PROCEDURE)
C0199968|T037|274502001|SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR TRANSFUSION |ANTIHEMOPHILIC FACTOR TRANSFUSION (PROCEDURE)
C0199968|T037|274502001|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR TRANSFUSION|ANTIHEMOPHILIC FACTOR TRANSFUSION (PROCEDURE)
C0199968|T037|274502001|SNOMEDCT_US|TRANSFUSION OF ANTIHEMOPHILIC FACTOR|ANTIHEMOPHILIC FACTOR TRANSFUSION (PROCEDURE)
C0199968|T037|274502001|SNOMEDCT_US|TRANSFUSION OF ANTIHAEMOPHILIC FACTOR|ANTIHEMOPHILIC FACTOR TRANSFUSION (PROCEDURE)
C0199968|T037|274502001|SNOMEDCT_US|ANTIHAEMOPHILIC FACTOR TRANSFUSION|ANTIHEMOPHILIC FACTOR TRANSFUSION (PROCEDURE)
C0199968|T037|274502001|SNOMEDCT_US|TRANSFUSION OF ANTIHEMOPHILIC FACTOR |ANTIHEMOPHILIC FACTOR TRANSFUSION (PROCEDURE)
C0199968|T037|274502001|SNOMEDCT_US|ANTIHEMOPHILIC FACTOR TRANSFUSION |ANTIHEMOPHILIC FACTOR TRANSFUSION (PROCEDURE)
C2242940|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN 
C2242940|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN
C3161607|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN FACTOR XIII CONCENTRATE (HUMAN)
C3161607|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN FACTOR XIII CONCENTRATE (HUMAN) 
C2064859|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN FACTOR VIII (AHF, AHG)
C2064859|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN FACTOR VIII (AHF, AHG) 
C2064857|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN ALBUMIN, NORMAL SERUM 
C2064857|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN ALBUMIN, NORMAL SERUM
C2064858|T037||SNOMEDCT_US|PLASMA FRACTIONS, FACTOR IX COMPLEX (HUMAN)
C2064858|T037||SNOMEDCT_US|HUMAN FACTOR IX COMPLEX (HUMAN)
C2064858|T037||SNOMEDCT_US|HUMAN FACTOR IX COMPLEX (HUMAN) 
C2194217|T037||SNOMEDCT_US|FACTOR VIIA TRANSFUSION 
C2194217|T037||SNOMEDCT_US|FACTOR VIIA
C2194217|T037||SNOMEDCT_US|FACTOR VIIA 
C2069055|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN ALBUMIN + GLOBULIN 
C2069055|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN ALBUMIN + GLOBULIN
C2069056|T037||SNOMEDCT_US|PLASMA FRACTIONS, ANTITHROMBIN III (HUMAN) 
C2069056|T037||SNOMEDCT_US|PLASMA FRACTIONS, ANTITHROMBIN III (HUMAN)
C4064322|T037||SNOMEDCT_US|PLASMA FRACTIONS, COAGULATION FACTOR X (HUMAN) 
C4064322|T037||SNOMEDCT_US|PLASMA FRACTIONS, COAGULATION FACTOR X (HUMAN)
C4064322|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN FACTOR X
C1293889|T037|116797000|SNOMEDCT_US|COAGULATION FACTOR IX PRODUCT ADMINISTRATION BY INTRAVASCULAR INFUSION|TRANSFUSION OF FACTOR IX (PROCEDURE)
C1293889|T037|116797000|SNOMEDCT_US|TRANSFUSION OF FACTOR IX |TRANSFUSION OF FACTOR IX (PROCEDURE)
C1293889|T037|116797000|SNOMEDCT_US|TRANSFUSION OF FACTOR IX|TRANSFUSION OF FACTOR IX (PROCEDURE)
C1293888|T037|116798005|SNOMEDCT_US|COAGULATION FACTOR VII PRODUCT ADMINISTRATION BY INTRAVASCULAR INFUSION|TRANSFUSION OF FACTOR VII (PROCEDURE)
C1293888|T037|116798005|SNOMEDCT_US|TRANSFUSION OF FACTOR VII |TRANSFUSION OF FACTOR VII (PROCEDURE)
C1293888|T037|116798005|SNOMEDCT_US|TRANSFUSION OF FACTOR VII|TRANSFUSION OF FACTOR VII (PROCEDURE)
C1960763|T037|425524005|SNOMEDCT_US|TRANSFUSION ANTITHROMBIN III FACTOR |TRANSFUSION ANTITHROMBIN III FACTOR (PROCEDURE)
C1960763|T037|425524005|SNOMEDCT_US|TRANSFUSION ANTITHROMBIN III FACTOR|TRANSFUSION ANTITHROMBIN III FACTOR (PROCEDURE)
