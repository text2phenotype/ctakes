C0366777|T201|COMP|4544-3|LNCICU|Hematocrit|Hematocrit
C0362934|T201|COMP|804-5|LNCICU|White Blood Cells|Leukocytes
C0362923|T201|COMP|718-7|LNCICU|Hemoglobin|Hemoglobin
C0362994|T201|COMP|777-3|LNCICU|Platelet Count|Platelets
C0362906|T201|COMP|785-6|LNCICU|MCH|Erythrocyte mean corpuscular hemoglobin
C0362908|T201|COMP|787-2|LNCICU|MCV|Erythrocyte mean corpuscular volume
C0362910|T201|COMP|789-8|LNCICU|Red Blood Cells|Erythrocytes
C0362909|T201|COMP|788-0|LNCICU|RDW|Erythrocyte distribution width
C0364968|T201|COMP|2823-3|LNCICU|Potassium|Potassium
C0365095|T201|COMP|2951-2|LNCICU|Sodium|Sodium
C0364207|T201|COMP|2075-0|LNCICU|Chloride|Chloride
C0364096|T201|COMP|1963-8|LNCICU|Bicarbonate|Bicarbonate
C0363998|T201|COMP|1863-0|LNCICU|Anion Gap|Anion gap 4
C0365240|T201|COMP|3094-0|LNCICU|Urea Nitrogen|Urea nitrogen
C0364294|T201|COMP|2160-0|LNCICU|Creatinine|Creatinine
C0484731|T201|COMP|2345-7|LNCICU|Glucose|Glucose
C0364745|T201|COMP|2601-3|LNCICU|Magnesium|Magnesium
C0364133|T201|COMP|2000-8|LNCICU|Calcium, Total|Calcium
C1370010|T201|COMP|2777-1|LNCICU|Phosphate|Phosphate
C0486259|T201|COMP|5895-7|LNCICU|INR(PT)|Coagulation tissue factor induced.INR
C0482694|T201|COMP|5902-2|LNCICU|PT|Coagulation tissue factor induced
C0362947|T201|COMP|731-0|LNCICU|Lymphocytes|Lymphocytes
C0362958|T201|COMP|742-7|LNCICU|Monocytes|Monocytes
C0362978|T201|COMP|761-7|LNCICU|Neutrophils|Neutrophils
C0362892|T201|COMP|704-7|LNCICU|Basophils|Basophils
C0362900|T201|COMP|711-2|LNCICU|Eosinophils|Eosinophils
C0365392|T201|COMP|3173-2|LNCICU|PTT|Coagulation surface induced
C0364108|T201|COMP|1975-2|LNCICU|Bilirubin, Total|Bilirubin
C0368061|T201|COMP|5811-5|LNCICU|Specific Gravity|Specific gravity
C0550221|T201|COMP|11555-0|LNCICU|Base Excess|Base excess
C1369594|T201|COMP|34728-6|LNCICU|Calculated Total CO2|Carbon dioxide
C0550440|T201|COMP|11556-8|LNCICU|pO2|Oxygen
C0550246|T201|COMP|11557-6|LNCICU|pCO2|Carbon dioxide
C0363876|T201|COMP|1742-6|LNCICU|Alanine Aminotransferase (ALT)|Alanine aminotransferase
C0364055|T201|COMP|1920-8|LNCICU|Asparate Aminotransferase (AST)|Aspartate aminotransferase
C0484638|T201|COMP|6768-6|LNCICU|Alkaline Phosphatase|Alkaline phosphatase
C0368043|T201|COMP|5804-0|LNCICU|Protein|Protein
C0368032|T201|COMP|5797-6|LNCICU|Ketone|Ketones
C0368078|T201|COMP|5818-0|LNCICU|Urobilinogen|Urobilinogen
C0368018|T201|COMP|5792-7|LNCICU|Glucose|Glucose
C1315166|T201|COMP|32693-4|LNCICU|Lactate|Lactate
C0368002|T201|COMP|5778-6|LNCICU|Urine Color|Color
C0363885|T201|COMP|1751-7|LNCICU|Albumin|Albumin
C0367982|T201|COMP|5767-9|LNCICU|Urine Appearance|Appearance
C0368020|T201|COMP|5794-3|LNCICU|Blood|Hemoglobin
C0368040|T201|COMP|5802-4|LNCICU|Nitrite|Nitrite
C0367985|T201|COMP|5770-3|LNCICU|Bilirubin|Bilirubin
C0368080|T201|COMP|5822-2|LNCICU|Yeast|Yeast
C0368035|T201|COMP|5799-2|LNCICU|Leukocytes|Leukocyte esterase
C0368036|T201|COMP|5821-4|LNCICU|WBC|Leukocytes
C0368013|T201|COMP|5808-1|LNCICU|RBC|Erythrocytes
C0368011|T201|COMP|5787-7|LNCICU|Epithelial Cells|Epithelial cells
C0364961|T201|COMP|6298-4|LNCICU|Potassium, Whole Blood|Potassium
C0364127|T201|COMP|1994-3|LNCICU|Free Calcium|Calcium.ionized
C0364290|T201|COMP|2157-6|LNCICU|Creatine Kinase (CK)|Creatine kinase
C0364479|T201|COMP|2339-0|LNCICU|Glucose|Glucose
C0367984|T201|COMP|5769-5|LNCICU|Bacteria|Bacteria
C0362980|T201|COMP|763-3|LNCICU|Bands|Neutrophils.band form
C0484707|T201|COMP|6773-6|LNCICU|Creatine Kinase, MB Isoenzyme|Creatine kinase.MB
C0803379|T201|COMP|20570-8|LNCICU|Hematocrit, Calculated|Hematocrit
C0365091|T201|COMP|2947-0|LNCICU|Sodium, Whole Blood|Sodium
C0364674|T201|COMP|2532-0|LNCICU|Lactate Dehydrogenase (LD)|Lactate dehydrogenase
C0362933|T201|COMP|728-6|LNCICU|Hypochromia|Hypochromia
C0362954|T201|COMP|738-5|LNCICU|Macrocytes|Macrocytes
C0362890|T201|COMP|702-1|LNCICU|Anisocytosis|Anisocytosis
C0362957|T201|COMP|741-9|LNCICU|Microcytes|Microcytes
C0362949|T201|COMP|733-6|LNCICU|Atypical Lymphocytes|Lymphocytes.variant
C0944135|T201|COMP|28541-1|LNCICU|Metamyelocytes|Metamyelocytes/100 leukocytes
C0942460|T201|COMP|26498-6|LNCICU|Myelocytes|Myelocytes/100 leukocytes
C2363247|T201|COMP|779-9|LNCICU|Poikilocytosis|Poikilocytosis
C0365184|T201|COMP|3040-3|LNCICU|Lipase|Triacylglycerol lipase
C0364201|T201|COMP|2069-3|LNCICU|Chloride, Whole Blood|Chloride
C0484652|T201|COMP|1798-8|LNCICU|Amylase|Amylase
C0484851|T201|COMP|6598-7|LNCICU|Troponin T|Troponin T.cardiac
C0484448|T201|COMP|10378-8|LNCICU|Polychromasia|Polychromasia
C0802029|T201|COMP|13362-9|LNCICU|Length of Urine Collection|Collection duration
C0482705|T201|COMP|3255-7|LNCICU|Fibrinogen, Functional|Fibrinogen
C0362995|T201|COMP|778-1|LNCICU|Platelet Smear|Platelets
C0365160|T201|COMP|3016-3|LNCICU|Thyroid Stimulating Hormone|Thyrotropin
C1316377|T201|COMP|33914-3|LNCICU|Estimated GFR (MDRD equation)|Glomerular filtration rate/1.73 sq M.predicted
C0364101|T201|COMP|1968-7|LNCICU|Bilirubin, Direct|Bilirubin.glucuronidated+Bilirubin.albumin bound
C0364104|T201|COMP|1971-1|LNCICU|Bilirubin, Indirect|Bilirubin.non-glucuronidated
C0364295|T201|COMP|2161-8|LNCICU|Creatinine, Urine|Creatinine
C0363775|T201|COMP|1644-4|LNCICU|Triglycerides|Triglyceride^post 12H CFst
C0365099|T201|COMP|2955-3|LNCICU|Sodium, Urine|Sodium
C0364639|T201|COMP|2498-4|LNCICU|Iron|Iron
C0364708|T201|COMP|2093-3|LNCICU|Cholesterol, Total|Cholesterol
C0364411|T201|COMP|2276-4|LNCICU|Ferritin|Ferritin
C0364641|T201|COMP|2500-7|LNCICU|Iron Binding Capacity, Total|Iron binding capacity
C0803387|T201|COMP|20578-1|LNCICU|Vancomycin|Vancomycin
C0364221|T201|COMP|2085-9|LNCICU|Cholesterol, HDL|Cholesterol.in HDL
C0484684|T201|COMP|9322-9|LNCICU|Cholesterol Ratio (Total/HDL)|Cholesterol.total/Cholesterol.in HDL
C0366781|T201|COMP|4548-4|LNCICU|% Hemoglobin A1c|Hemoglobin A1c/Hemoglobin.total
C0364838|T201|COMP|2695-5|LNCICU|Osmolality, Urine|Osmolality
C2713147|T201|COMP|2090-9|LNCICU|Cholesterol, LDL, Calculated|Cholesterol.in LDL
C0368025|T201|COMP|5796-8|LNCICU|Hyaline Casts|Hyaline casts
C0362989|T201|COMP|772-4|LNCICU|Nucleated Red Cells|Erythrocytes.nucleated
C0486210|T201|COMP|8247-9|LNCICU|Urine Mucous|Mucus
C1642563|T201|COMP|42662-7|LNCICU|Benzodiazepine Screen|Benzodiazepines
C0365608|T201|COMP|3376-1|LNCICU|Barbiturate Screen|Barbiturates
C0366299|T201|COMP|4073-3|LNCICU|Tricyclic Antidepressant Screen|Tricyclic antidepressants
C0364304|T201|COMP|2170-9|LNCICU|Vitamin B12|Cyanocobalamin.true
C0365241|T201|COMP|3095-7|LNCICU|Urea Nitrogen, Urine|Urea nitrogen
C0364092|T201|COMP|1959-6|LNCICU|Calculated Bicarbonate, Whole Blood|Bicarbonate
C0362991|T201|COMP|774-0|LNCICU|Ovalocytes|Ovalocytes
C0803378|T201|COMP|20569-0|LNCICU|CK-MB Index|Creatine kinase.MB/Creatine kinase.total
C0365627|T201|COMP|3397-7|LNCICU|Cocaine, Urine|Cocaine
C0365620|T201|COMP|3390-2|LNCICU|Benzodiazepine Screen, Urine|Benzodiazepines
C0365583|T201|COMP|3349-8|LNCICU|Amphetamine Screen, Urine|Amphetamines
C0365609|T201|COMP|3377-9|LNCICU|Barbiturate Screen, Urine|Barbiturates
C0366106|T201|COMP|3879-4|LNCICU|Opiate Screen, Urine|Opiates
C0366000|T201|COMP|3773-9|LNCICU|Methadone, Urine|Methadone
C0365029|T201|COMP|2885-2|LNCICU|Protein, Total|Protein
C0364419|T201|COMP|2284-8|LNCICU|Folate|Folate
C0367799|T201|COMP|5642-4|LNCICU|Ethanol|Ethanol
C0800956|T201|COMP|17849-1|LNCICU|Reticulocyte Count, Automated|Reticulocytes/100 erythrocytes
C0365531|T201|COMP|3297-9|LNCICU|Acetaminophen|Acetaminophen
C0364971|T201|COMP|2828-2|LNCICU|Potassium, Urine|Potassium
C0366775|T201|COMP|4542-7|LNCICU|Haptoglobin|Haptoglobin
C0366250|T201|COMP|4023-8|LNCICU|Salicylate|Salicylates
C0484419|T201|COMP|7790-9|LNCICU|Burr Cells|Burr cells
C0364210|T201|COMP|2078-4|LNCICU|Chloride, Urine|Chloride
C0364275|T201|COMP|2143-6|LNCICU|Cortisol|Cortisol
C0363002|T201|COMP|800-3|LNCICU|Schistocytes|Schistocytes
C0364835|T201|COMP|2692-2|LNCICU|Osmolality, Measured|Osmolality
C0486200|T201|COMP|8246-1|LNCICU|Amorphous Crystals|Amorphous sediment
C0368021|T201|COMP|5793-5|LNCICU|Granular Casts|Granular casts
C0365168|T201|COMP|3024-7|LNCICU|Thyroxine (T4), Free|Thyroxine.free
C0364474|T201|COMP|2336-6|LNCICU|Globulin|Globulin
C0366770|T201|COMP|4537-7|LNCICU|Sedimentation Rate|Erythrocyte sedimentation rate
C0362997|T201|COMP|7791-7|LNCICU|Teardrop Cells|Dacryocytes
C1316226|T201|COMP|33762-6|LNCICU|NTproBNP|Natriuretic peptide.B prohormone N-Terminal
C0365228|T201|COMP|3084-1|LNCICU|Uric Acid|Urate
C1113987|T201|COMP|30089-7|LNCICU|Transitional Epithelial Cells|Transitional cells
C0366194|T201|COMP|3967-7|LNCICU|Phenytoin|Phenytoin
C0365031|T201|COMP|2887-8|LNCICU|Total Protein, Urine|Protein
C0364121|T201|COMP|1988-5|LNCICU|C-Reactive Protein|C reactive protein
C0484456|T201|COMP|10381-2|LNCICU|Target Cells|Target cells
C0365034|T201|COMP|2890-2|LNCICU|Protein/Creatinine Ratio|Protein/Creatinine
C0550543|T201|COMP|10839-9|LNCICU|Troponin I|Troponin I.cardiac
C0368404|T201|COMP|5196-1|LNCICU|Hepatitis B Surface Antigen|Hepatitis B virus surface Ag
C0799293|T201|COMP|16128-1|LNCICU|Hepatitis C Virus Antibody|Hepatitis C virus Ab
C0942430|T201|COMP|26465-5|LNCICU|WBC, CSF|Leukocytes
C0942441|T201|COMP|26479-6|LNCICU|Lymphs|Lymphocytes/100 leukocytes
C0942448|T201|COMP|26486-1|LNCICU|Monocytes|Monocytes/100 leukocytes
C0945364|T201|COMP|26517-3|LNCICU|Polys|Polymorphonuclear cells/100 leukocytes
C0368401|T201|COMP|5193-8|LNCICU|Hepatitis B Surface Antibody|Hepatitis B virus surface Ab
C0942423|T201|COMP|26454-9|LNCICU|RBC, CSF|Erythrocytes
C1953449|T201|COMP|48065-7|LNCICU|D-Dimer|Fibrin D-dimer FEU
C0365023|T201|COMP|2880-3|LNCICU|Total Protein, CSF|Protein
C0364482|T201|COMP|2342-4|LNCICU|Glucose, CSF|Glucose
C1114106|T201|COMP|30226-5|LNCICU|Fibrin Degradation Products|Fibrin+Fibrinogen fragments
C0484920|T201|COMP|10535-3|LNCICU|Digoxin|Digoxin
C0945182|T201|COMP|25156-1|LNCICU|Eosinophils|Eosinophils
C0368391|T201|COMP|5187-0|LNCICU|Hepatitis B Virus Core Antibody|Hepatitis B virus core Ab
C1114897|T201|COMP|30394-1|LNCICU|Granulocyte Count|Granulocytes
C0362891|T201|COMP|703-9|LNCICU|Basophilic Stippling|Basophilic stippling
C0365170|T201|COMP|3026-2|LNCICU|Thyroxine (T4)|Thyroxine
C0799525|T201|COMP|16362-6|LNCICU|Ammonia|Ammonia
C0364874|T201|COMP|2731-8|LNCICU|Parathyroid Hormone|Parathyrin.intact
C0881624|T201|COMP|24351-9|LNCICU|Protein Electrophoresis|Protein fractions panel
C0365000|T201|COMP|2857-1|LNCICU|Prostate Specific Antigen|Prostate specific Ag
C0364605|T201|COMP|2465-3|LNCICU|Immunoglobulin G|IgG
C0942079|T201|COMP|26052-1|LNCICU|Renal Epithelial Cells|Epithelial cells.renal
C0942432|T201|COMP|26467-1|LNCICU|WBC, Pleural|Leukocytes
C0942443|T201|COMP|26481-2|LNCICU|Lymphocytes|Lymphocytes/100 leukocytes
C0942477|T201|COMP|26519-9|LNCICU|Polys|Polymorphonuclear cells/100 leukocytes
C1315831|T201|COMP|33362-5|LNCICU|Monos|Monocytes/100 leukocytes
C0803372|T201|COMP|20563-3|LNCICU|Carboxyhemoglobin|Carboxyhemoglobin/Hemoglobin.total
C0484416|T201|COMP|7789-1|LNCICU|Acanthocytes|Acanthocytes
C0365026|T201|COMP|2882-9|LNCICU|Total Protein, Pleural|Protein
C0363004|T201|COMP|802-9|LNCICU|Spherocytes|Spherocytes
C0364672|T201|COMP|2530-4|LNCICU|Lactate Dehydrogenase, Pleural|Lactate dehydrogenase
C0942424|T201|COMP|26456-4|LNCICU|RBC, Pleural|Erythrocytes
C0364759|T201|COMP|2614-6|LNCICU|Methemoglobin|Methemoglobin/Hemoglobin.total
C1507819|T201|COMP|35668-3|LNCICU|Gentamicin|Gentamicin
C0367391|T201|COMP|5047-6|LNCICU|Anti-Nuclear Antibody|Nuclear Ab
C0364598|T201|COMP|2458-8|LNCICU|Immunoglobulin A|IgA
C0364459|T201|COMP|2324-2|LNCICU|Gamma Glutamyltransferase|Gamma glutamyl transferase
C1316630|T201|COMP|34167-7|LNCICU|Large Platelets|Platelets.large
C0364486|T201|COMP|2346-5|LNCICU|Glucose, Pleural|Glucose
C0364612|T201|COMP|2472-9|LNCICU|Immunoglobulin M|IgM
C2973277|T201|COMP|10330-9|LNCICU|Monos|Monocytes/100 leukocytes
C0549816|T201|COMP|11031-2|LNCICU|Lymphocytes|Lymphocytes/100 leukocytes
C0942476|T201|COMP|26518-1|LNCICU|Polys|Polymorphonuclear cells/100 leukocytes
C0365197|T201|COMP|3053-6|LNCICU|Triiodothyronine (T3)|Triiodothyronine
C0368455|T201|COMP|5220-9|LNCICU|HIV Antibody|HIV 1 Ab
C0363888|T201|COMP|1754-1|LNCICU|Albumin, Urine|Albumin
C1146797|T201|COMP|31112-6|LNCICU|Reticulocyte Count, Manual|Reticulocytes/100 erythrocytes
C0364171|T201|COMP|2039-6|LNCICU|Carcinoembyronic Antigen (CEA)|Carcinoembryonic Ag
C0368387|T201|COMP|5183-9|LNCICU|Hepatitis A Virus Antibody|Hepatitis A virus Ab
C0363968|T201|COMP|1834-1|LNCICU|Alpha-Fetoprotein|Alpha-1-Fetoprotein
C0801308|T201|COMP|18262-6|LNCICU|Cholesterol, LDL, Measured|Cholesterol.in LDL
C0550490|T201|COMP|13438-7|LNCICU|Prot. Electrophoresis, Urine|Protein pattern
C0798131|T201|COMP|14958-3|LNCICU|Albumin/Creatinine, Urine|Albumin/Creatinine
C0484426|T201|COMP|10373-9|LNCICU|Fragmented Cells|Fragments
C0945358|T201|COMP|26468-9|LNCICU|WBC, Ascites|Leukocytes
C0942444|T201|COMP|26482-0|LNCICU|Lymphocytes|Lymphocytes/100 leukocytes
C0942450|T201|COMP|26488-7|LNCICU|Monocytes|Monocytes/100 leukocytes
C0942478|T201|COMP|26520-7|LNCICU|Polys|Polymorphonuclear cells/100 leukocytes
C0362999|T201|COMP|781-5|LNCICU|Promyelocytes|Promyelocytes
C0942425|T201|COMP|26457-2|LNCICU|RBC, Ascites|Erythrocytes
C0942431|T201|COMP|26466-3|LNCICU|WBC, Other Fluid|Leukocytes
C1544494|T201|COMP|40520-9|LNCICU|Macrophages|Macrophages/100 leukocytes
C1114284|T201|COMP|30431-1|LNCICU|Mesothelial Cells|Mesothelial cells/100 leukocytes
C0367994|T201|COMP|5774-5|LNCICU|Calcium Oxalate Crystals|Calcium oxalate crystals
C0484417|T201|COMP|10371-3|LNCICU|Bite Cells|Bite cells
C0945355|T201|COMP|26455-6|LNCICU|RBC, Other Fluid|Erythrocytes
C0366727|T201|COMP|4498-2|LNCICU|C4|Complement C4
C0363882|T201|COMP|1748-3|LNCICU|Albumin, Pleural|Albumin
C0367699|T201|COMP|5567-3|LNCICU|Acetone|Acetone
C0802081|T201|COMP|19159-3|LNCICU|Urine Specimen Type|Urinalysis specimen collection method
C1544491|T201|COMP|40517-5|LNCICU|Macrophage|Macrophages/100 leukocytes
C0365027|T201|COMP|2883-7|LNCICU|Total Protein, Ascites|Protein
C0549819|T201|COMP|12230-9|LNCICU|Macrophage|Macrophages/100 leukocytes
C0366711|T201|COMP|4485-9|LNCICU|C3|Complement C3
C0368077|T201|COMP|5817-2|LNCICU|Uric Acid Crystals|Urate crystals
C1114285|T201|COMP|30432-9|LNCICU|Mesothelial Cell|Mesothelial cells/100 leukocytes
C0364923|T201|COMP|2778-9|LNCICU|Phosphate, Urine|Phosphate
C1114279|T201|COMP|30426-1|LNCICU|Macrophage|Macrophages/100 leukocytes
C0943674|T201|COMP|28009-9|LNCICU|Urine Volume|Specimen volume
C0363883|T201|COMP|1749-1|LNCICU|Albumin, Ascites|Albumin
C0364097|T201|COMP|1964-6|LNCICU|Bicarbonate, Urine|Bicarbonate
C0484553|T201|COMP|8127-3|LNCICU|CD4 Cells, Percent|Cells.CD4
C0484547|T201|COMP|8122-4|LNCICU|CD3 Cells, Percent|Cells.CD3
C0364673|T201|COMP|2531-2|LNCICU|Lactate Dehydrogenase, Ascites|Lactate dehydrogenase
C0364136|T201|COMP|2004-0|LNCICU|Calcium, Urine|Calcium
C0485879|T201|COMP|6928-6|LNCICU|Rheumatoid Factor|Rheumatoid factor
C0484444|T201|COMP|7795-8|LNCICU|Pappenheimer Bodies|Pappenheimer bodies
C0364487|T201|COMP|2347-3|LNCICU|Glucose, Ascites|Glucose
C1955034|T201|COMP|49275-1|LNCICU|Immunofixation|Interpretation
C0363931|T201|COMP|1797-0|LNCICU|Amylase, Ascites|Amylase
C0484567|T201|COMP|8137-2|LNCICU|CD8 Cells, Percent|Cells.CD8
C0942440|T201|COMP|26478-8|LNCICU|Lymphocytes, Percent|Lymphocytes/100 leukocytes
C0945357|T201|COMP|26464-8|LNCICU|WBC Count|Leukocytes
C0942437|T201|COMP|26474-7|LNCICU|Absolute Lymphocyte Count|Lymphocytes
C0484554|T201|COMP|8128-1|LNCICU|Absolute CD4 Count|Cells.CD4/100 cells
C0362945|T201|COMP|729-4|LNCICU|Other Cells|Leukocytes other
C0879885|T201|COMP|22314-9|LNCICU|Hepatitis A Virus IgM Antibody|Hepatitis A virus Ab.IgM
C0797153|T201|COMP|13965-9|LNCICU|Homocysteine|Homocysteine
C1370068|T201|COMP|35279-9|LNCICU|Anti-Neutrophil Cytoplasmic Antibody|Neutrophil cytoplasmic Ab
C1955035|T201|COMP|49276-9|LNCICU|Immunofixation, Urine|Interpretation
C0364239|T201|COMP|2119-6|LNCICU|Human Chorionic Gonadotropin|Choriogonadotropin
C1146889|T201|COMP|31204-1|LNCICU|Hepatitis B Core Antibody, IgM|Hepatitis B virus core Ab.IgM
C1114241|T201|COMP|30379-2|LNCICU|Eosinophils|Eosinophils/100 leukocytes
C0366312|T201|COMP|4086-5|LNCICU|Valproic Acid|Valproate
C0363930|T201|COMP|1796-2|LNCICU|Amylase, Pleural|Amylase
C0484550|T201|COMP|8124-0|LNCICU|Absolute CD3 Count|Cells.CD3/100 cells
C0484555|T201|COMP|8129-9|LNCICU|CD4/CD8 Ratio|Cells.CD4/Cells.CD8
C0484568|T201|COMP|8138-0|LNCICU|Absolute CD8 Count|Cells.CD8/100 cells
C0363929|T201|COMP|1795-4|LNCICU|Amylase, Body Fluid|Amylase
C0364236|T201|COMP|2106-3|LNCICU|HCG, Urine, Qualitative|Choriogonadotropin (pregnancy test)
C0942421|T201|COMP|26452-3|LNCICU|Eosinophils|Eosinophils/100 leukocytes
C0800930|T201|COMP|17823-6|LNCICU|CD45|Cells.CD45/100 cells
C0797600|T201|COMP|14422-0|LNCICU|Bilirubin, Total, Ascites|Bilirubin
C0942420|T201|COMP|26451-5|LNCICU|Eosinophils|Eosinophils/100 leukocytes
C0800936|T201|COMP|17829-3|LNCICU|CD19|Cells.CD19/100 cells
C0364296|T201|COMP|2162-6|LNCICU|24 hr Creatinine|Creatinine
C0485832|T201|COMP|8061-4|LNCICU|Anti-Nuclear Antibody, Titer|Nuclear Ab
C0364669|T201|COMP|2528-8|LNCICU|Lactate Dehydrogenase, CSF|Lactate dehydrogenase
C0800942|T201|COMP|17835-0|LNCICU|Monocytes|Monocytes/100 leukocytes
C0942433|T201|COMP|26469-7|LNCICU|WBC, Joint Fluid|Leukocytes
C0942445|T201|COMP|26483-8|LNCICU|Lymphocytes|Lymphocytes/100 leukocytes
C0945365|T201|COMP|26522-3|LNCICU|Polys|Polymorphonuclear cells/100 leukocytes
C0482696|T201|COMP|3243-3|LNCICU|Thrombin|Coagulation thrombin induced
C0365025|T201|COMP|2881-1|LNCICU|Total Protein, Body Fluid|Protein
C1544696|T201|COMP|40741-1|LNCICU|Platelet Clumps|Platelet clump
C0365230|T201|COMP|3086-6|LNCICU|Uric Acid, Urine|Urate
C0942426|T201|COMP|26458-0|LNCICU|RBC, Joint Fluid|Erythrocytes
C0364484|T201|COMP|2344-0|LNCICU|Glucose, Body Fluid|Glucose
C0365326|T201|COMP|3182-3|LNCICU|Anticardiolipin Antibody IgM|Cardiolipin Ab.IgM
C0485838|T201|COMP|8065-5|LNCICU|Anticardiolipin Antibody IgG|Cardiolipin Ab.IgG
C1114799|T201|COMP|31017-7|LNCICU|Tissue Transglutaminase Ab, IgA|Tissue transglutaminase Ab.IgA
C0484428|T201|COMP|7793-3|LNCICU|Howell-Jolly Bodies|Howell-Jolly bodies
C0945626|T201|COMP|28544-5|LNCICU|Mesothelial cells|Mesothelial cells/100 leukocytes
C1543046|T201|COMP|38924-7|LNCICU|H/O Smear|TBX5 gene targeted mutation analysis
C0362896|T201|COMP|708-8|LNCICU|Blasts|Blasts
C0364671|T201|COMP|2529-6|LNCICU|LD, Body Fluid|Lactate dehydrogenase
C0364742|T201|COMP|2598-1|LNCICU|Magnesium, Urine|Magnesium
C0363881|T201|COMP|1747-5|LNCICU|Albumin, Body Fluid|Albumin
C0366196|T201|COMP|3969-3|LNCICU|Phenytoin, Free|Phenytoin.free
C0484977|T201|COMP|10548-6|LNCICU|Phenytoin, Percent Free|Phenytoin.free/Phenytoin.total
C1114242|T201|COMP|30380-0|LNCICU|Eosinophils|Eosinophils/100 leukocytes
C0365171|T201|COMP|3027-0|LNCICU|Calculated TBG|Thyroxine/Thyroxine binding globulin
C0365194|T201|COMP|3050-2|LNCICU|Uptake Ratio|Triiodothyronine resin uptake (T3RU)
C1147899|T201|COMP|32215-6|LNCICU|Calculated Thyroxine (T4) Index|Thyroxine free index
C0797437|T201|COMP|14252-1|LNCICU|Anti-Smooth Muscle Antibody|Smooth muscle Ab
C0365137|T201|COMP|2986-8|LNCICU|Testosterone|Testosterone
C0797421|T201|COMP|14236-4|LNCICU|Anti-Mitochondrial Antibody|Mitochondria Ab
C0800933|T201|COMP|17826-9|LNCICU|CD3|Cells.CD3/100 cells
C0550284|T201|COMP|12191-3|LNCICU|Creatinine, Ascites|Creatinine
C0365750|T201|COMP|3521-2|LNCICU|Cyclosporin|cycloSPORINE
C0486211|T201|COMP|8248-7|LNCICU|Sperm|Spermatozoa
C1315158|T201|COMP|32684-3|LNCICU|Heparin, LMW|Heparin.low molecular weight
C0484675|T201|COMP|10334-1|LNCICU|CA-125|Cancer Ag 125
C2735785|T201|COMP|57418-6|LNCICU|CD20|Cells.CD20/100 cells
C1979282|T201|COMP|51217-8|LNCICU|CD10|Cells.CD10/100 cells
C2735790|T201|COMP|57423-6|LNCICU|CD5|Cells.CD5/100 cells
C0482602|T201|COMP|2842-3|LNCICU|Prolactin|Prolactin
C0943513|T201|COMP|27818-4|LNCICU|Protein C, Functional|Protein C actual/Normal
C0365135|T201|COMP|2991-8|LNCICU|Calculated Free Testosterone|Testosterone.free
C0367401|T201|COMP|5117-7|LNCICU|Cryoglobulin|Cryoglobulin
C0549840|T201|COMP|13047-6|LNCICU|Plasma Cells|Plasma cells/100 leukocytes
C0943506|T201|COMP|27811-9|LNCICU|Antithrombin|Antithrombin actual/Normal
C1979422|T201|COMP|51381-2|LNCICU|HLA-DR|Cells.HLA-DR+/100 cells
C0368065|T201|COMP|5814-9|LNCICU|Triple Phosphate Crystals|Triple phosphate crystals
C0881684|T201|COMP|24429-3|LNCICU|Blood Parasite Smear|Parasite identified
C1507821|T201|COMP|35670-9|LNCICU|Tobramycin|Tobramycin
C0366174|T201|COMP|3947-9|LNCICU|Phenobarbital|PHENobarbital
C0484790|T201|COMP|9618-0|LNCICU|Cholesterol, Pleural|Cholesterol
C1977710|T201|COMP|51269-9|LNCICU|CD23|Cells.CD23/100 cells
C0796707|T201|COMP|13513-7|LNCICU|Iron Stain|Iron.microscopic observation
C2735796|T201|COMP|57428-5|LNCICU|FMC-7|Cells.FMC7/100 cells
C0797578|T201|COMP|14399-0|LNCICU|Creatinine, Pleural|Creatinine
C1114269|T201|COMP|30416-2|LNCICU|Atypical Lymphocytes|Lymphocytes.variant/100 leukocytes
C1545207|T201|COMP|41284-1|LNCICU|Non-squamous Epithelial Cells|Epithelial cells.non-squamous
C0485103|T201|COMP|10346-5|LNCICU|Hemogloblin A|Hemoglobin A
C0366795|T201|COMP|4561-7|LNCICU|Hemoglobin C|Hemoglobin C/Hemoglobin.total
C0366857|T201|COMP|4622-7|LNCICU|Hemogloblin S|Hemoglobin S
C0797899|T201|COMP|14725-6|LNCICU|Fluid Type|Fluid
C0368034|T201|COMP|5820-6|LNCICU|WBC Casts|Leukocyte casts
C0365948|T201|COMP|3719-2|LNCICU|Lithium|Lithium
C1148230|T201|COMP|32546-4|LNCICU|Quantitative G6PD|Glucose-6-Phosphate dehydrogenase
C0364785|T201|COMP|2640-1|LNCICU|Myoglobin, Urine|Myoglobin
C0550836|T201|COMP|11153-4|LNCICU|Hematocrit, Other Fluid|Hematocrit
C0365661|T201|COMP|3432-2|LNCICU|Carbamazepine|carBAMazepine
C0482633|T201|COMP|3209-4|LNCICU|Factor VIII|Coagulation factor VIII activity actual/Normal
C0484445|T201|COMP|10377-0|LNCICU|Pencil Cells|Pencil cells
C0798239|T201|COMP|15067-2|LNCICU|Follicle Stimulating Hormone|Follitropin
C0942469|T201|COMP|26509-0|LNCICU|Bands|Neutrophils.band form/100 leukocytes
C1977718|T201|COMP|51340-8|LNCICU|CD45|Cells.CD45/100 cells
C2735792|T201|COMP|57425-1|LNCICU|CD7|Cells.CD7/100 cells
C0800934|T201|COMP|17827-7|LNCICU|CD2|Cells.CD2/100 cells
C1369982|T201|COMP|1974-5|LNCICU|Bilirubin, Total, Body Fluid|Bilirubin
C1148209|T201|COMP|32525-8|LNCICU|CD19|Cells.CD19/100 cells
C0362983|T201|COMP|766-6|LNCICU|Hypersegmented Neutrophils|Neutrophils.hypersegmented
C0484556|T201|COMP|8130-7|LNCICU|CD45|Cells.CD45/100 cells
C0484540|T201|COMP|8117-4|LNCICU|CD19|Cells.CD19/100 cells
C0944729|T201|COMP|29247-4|LNCICU|Rapamycin|Sirolimus
C0550281|T201|COMP|12190-5|LNCICU|Creatinine, Body Fluid|Creatinine
C0483101|T201|COMP|5380-1|LNCICU|Anti-Thyroglobulin Antibodies|Thyroglobulin Ab
C0367411|T201|COMP|5130-0|LNCICU|Double Stranded DNA|DNA double strand Ab
C1765334|T201|COMP|3427-2|LNCICU|Marijuana|Cannabinoids
C1979281|T201|COMP|51216-0|LNCICU|CD10|Cells.CD10/100 cells
C0942419|T201|COMP|26449-9|LNCICU|Eosinophil Count|Eosinophils
C1315845|T201|COMP|33376-5|LNCICU|Macrophage|Macrophages/100 leukocytes
C0484544|T201|COMP|8119-0|LNCICU|CD20|Cells.CD20/100 cells
C0484561|T201|COMP|8132-3|LNCICU|CD5|Cells.CD5/100 cells
C1979421|T201|COMP|51380-4|LNCICU|HLA-DR|Cells.HLA-DR+/100 cells
C0486204|T201|COMP|9842-6|LNCICU|Urine Casts, Other|Casts
C0364473|T201|COMP|2335-8|LNCICU|Blood, Occult|Hemoglobin.gastrointestinal
C1148213|T201|COMP|32529-0|LNCICU|CD3|Cells.CD3/100 cells
C1507792|T201|COMP|35640-2|LNCICU|CD5|Cells.CD5/100 cells
C0363731|T201|COMP|1599-0|LNCICU|Luteinizing Hormone|Lutropin^baseline
C0484528|T201|COMP|8107-5|LNCICU|CD10|Cells.CD10/100 cells
C0484792|T201|COMP|9619-8|LNCICU|Triglycerides, Pleural|Triglyceride
C1315202|T201|COMP|32731-2|LNCICU|Beta-2 Microglobulin|Beta 2 globulin
C1315095|T201|COMP|32621-5|LNCICU|HLA-DR|HLA-DR
C0881625|T201|COMP|24352-7|LNCICU|PEP, CSF|Protein fractions panel
C1146787|T201|COMP|31102-7|LNCICU|Protein S, Functional|Protein S actual/Normal
C0365033|T201|COMP|2889-4|LNCICU|24 hr Protein|Protein
C0368007|T201|COMP|5783-6|LNCICU|Urine Crystals, Other|Crystals.unidentified
C0551368|T201|COMP|8099-4|LNCICU|Thyroid Peroxidase Antibodies|Thyroperoxidase Ab
C1315839|T201|COMP|33370-8|LNCICU|Atypical Lymphocytes|Lymphocytes.variant/100 leukocytes
C1507793|T201|COMP|35641-0|LNCICU|CD7|Cells.CD7/100 cells
C0484565|T201|COMP|8135-6|LNCICU|CD7|Cells.CD7/100 cells
C0800949|T201|COMP|17842-6|LNCICU|Cancer Antigen 27.29|Cancer Ag 27-29
C1148211|T201|COMP|32527-4|LNCICU|CD2|Cells.CD2/100 cells
C0484542|T201|COMP|8118-2|LNCICU|CD2|Cells.CD2/100 cells
C0366878|T201|COMP|4644-1|LNCICU|Hemosiderin|Hemosiderin
C0800347|T201|COMP|17220-5|LNCICU|FMC-7|Cells.FMC7/100 cells
C1315838|T201|COMP|33369-0|LNCICU|Atypical Lymphocytes|Lymphocytes.variant/100 leukocytes
C0366275|T201|COMP|4049-3|LNCICU|Theophylline|Theophylline
C0797206|T201|COMP|14018-6|LNCICU|CD23|Cells.CD23/100 cells
C1977709|T201|COMP|51268-1|LNCICU|CD23|Cells.CD23/100 cells
C1369871|T201|COMP|35070-2|LNCICU|Basophils|Basophils/100 leukocytes
C1316027|T201|COMP|33558-8|LNCICU|Creatinine Clearance|Creatinine renal clearance
C1954411|T201|COMP|48778-5|LNCICU|NRBC|Erythrocytes.nucleated/100 cells
C2359896|T201|COMP|51633-6|LNCICU|Young Cells|Platelets.reticulated/100 platelets
C0942470|T201|COMP|26510-8|LNCICU|Bands|Neutrophils.band form/100 leukocytes
C0368079|T201|COMP|5819-8|LNCICU|Waxy Casts|Waxy casts
C2735535|T201|COMP|57400-4|LNCICU|CD34|Cells.CD34/100 cells
C1114236|T201|COMP|30374-3|LNCICU|Basophils|Basophils/100 leukocytes
C0482773|T201|COMP|6012-9|LNCICU|Von Willebrand Factor Antigen|von Willebrand factor Ag
C0365157|T201|COMP|3013-0|LNCICU|Thyroglobulin|Thyroglobulin
C1979107|T201|COMP|51237-6|LNCICU|CD13|Cells.CD13/100 cells
C0798373|T201|COMP|15202-5|LNCICU|Potassium, Stool|Potassium
C0798378|T201|COMP|15207-4|LNCICU|Sodium, Stool|Sodium
C0797624|T201|COMP|14447-7|LNCICU|Triglycerides, Ascites|Triglyceride
C1979344|T201|COMP|51301-0|LNCICU|CD4|Cells.CD4/100 cells
C1544496|T201|COMP|40522-5|LNCICU|Plasma Cells|Plasma cells/100 leukocytes
C1979336|T201|COMP|51293-9|LNCICU|CD33|Cells.CD33/100 cells
C0367986|T201|COMP|5771-1|LNCICU|Bilirubin Crystals|Bilirubin crystals
C0366785|T201|COMP|4552-6|LNCICU|Hemoglobin A2|Hemoglobin A2/Hemoglobin.total
C0364471|T201|COMP|2333-3|LNCICU|Gastrin|Gastrin
C1627309|T201|COMP|42866-4|LNCICU|CD117|Cells.CD117/100 cells
C1979413|T201|COMP|51372-1|LNCICU|CD8|Cells.CD8+HLA-DR+/100 cells
C0484562|T201|COMP|8133-1|LNCICU|CD56|Cells.CD56/100 cells
C0484438|T201|COMP|10376-2|LNCICU|MacroOvalocytes|Macrocytes.oval
C0800941|T201|COMP|17834-3|LNCICU|Eosinophils|Eosinophils/100 leukocytes
C0797599|T201|COMP|14421-2|LNCICU|Bilirubin, Total, Pleural|Bilirubin
C0944137|T201|COMP|28543-7|LNCICU|Basophils|Basophils/100 leukocytes
C1979303|T201|COMP|51251-7|LNCICU|CD15|Cells.CD15/100 cells
C0364836|T201|COMP|2693-0|LNCICU|Osmolality, Stool|Osmolality
C1148191|T201|COMP|32507-6|LNCICU|CD14|Cells.CD14/100 cells
C0485104|T201|COMP|9749-3|LNCICU|Hemoglobin F|Hemoglobin F
C0550841|T201|COMP|13055-9|LNCICU|Heparin|Heparin
C0365274|T201|COMP|3128-6|LNCICU|Serum Viscosity|Viscosity
C1369870|T201|COMP|35069-4|LNCICU|Basophils|Basophils/100 leukocytes
C0484673|T201|COMP|6874-2|LNCICU|24 hr Calcium|Calcium
C1114270|T201|COMP|30417-0|LNCICU|Atypical Lymphocytes|Lymphocytes.variant/100 leukocytes
C0484551|T201|COMP|8125-7|LNCICU|CD34|Cells.CD34/100 cells
C0943517|T201|COMP|27823-4|LNCICU|Protein S, Antigen|Protein S Ag actual/Normal
C0365094|T201|COMP|2950-4|LNCICU|Sodium, Body Fluid|Sodium
C0484522|T201|COMP|8102-6|LNCICU|CD33|Cells.CD33/100 cells
C0484534|T201|COMP|8110-9|LNCICU|CD13|Cells.CD13/100 cells
C1315673|T201|COMP|33202-3|LNCICU|CD11c|Cells.CD11c/100 cells
C0484535|T201|COMP|8111-7|LNCICU|CD14|Cells.CD14/100 cells
C1979405|T201|COMP|51365-5|LNCICU|CD64|Cells.CD64/100 cells
C0484533|T201|COMP|8109-1|LNCICU|CD11c|Cells.CD11c/100 cells
C0364964|T201|COMP|2821-7|LNCICU|Potassium|Potassium
C1979365|T201|COMP|51319-2|LNCICU|CD41|Cells.CD41/100 cells
C0800929|T201|COMP|17822-8|LNCICU|CD4|Cells.CD3+CD4+/100 cells
C0800931|T201|COMP|17824-4|LNCICU|CD8|Cells.CD3+CD8+/100 cells
C0364378|T201|COMP|2243-4|LNCICU|Estradiol|Estradiol
C1315679|T201|COMP|33208-0|LNCICU|Glyco A|Cells.CD235a/100 cells
C0482622|T201|COMP|3198-9|LNCICU|Factor VII|Coagulation factor VII activity actual/Normal
C1544492|T201|COMP|40518-3|LNCICU|Plasma|Plasma cells/100 leukocytes
C0366061|T201|COMP|3834-9|LNCICU|N-Acetylprocainamide (NAPA)|N-acetylprocainamide
C0366209|T201|COMP|3982-6|LNCICU|Procainamide|Procainamide
C0800245|T201|COMP|17117-3|LNCICU|CD15|Cells.CD15/100 cells
C0800275|T201|COMP|17148-8|LNCICU|CD41|Cells.CD41/100 cells
C0366892|T201|COMP|4659-9|LNCICU|Leukocyte Alkaline Phosphatase|Phosphatase.leukocyte
C0800235|T201|COMP|17107-4|LNCICU|CD117|Cells.CD117/100 cells
C0364490|T201|COMP|2350-7|LNCICU|Glucose, Urine|Glucose
C0484566|T201|COMP|8136-4|LNCICU|CD71|Cells.CD71/100 cells
C0800310|T201|COMP|17183-5|LNCICU|CD64|Cells.CD64/100 cells
C1146806|T201|COMP|17221-3|LNCICU|Glyco A|Cells.CD235a/100 cells
C0365239|T201|COMP|3093-2|LNCICU|Urea Nitrogen, Body Fluid|Urea nitrogen
C0482617|T201|COMP|3193-0|LNCICU|Factor V|Coagulation factor V activity actual/Normal
C0482641|T201|COMP|3218-5|LNCICU|Factor X|Coagulation factor X activity actual/Normal
C0550533|T201|COMP|12228-3|LNCICU|Triglycer|Triglyceride
C0798329|T201|COMP|15158-9|LNCICU|Chloride, Stool|Chloride
C0368012|T201|COMP|5807-3|LNCICU|RBC Casts|Erythrocyte casts
C0550585|T201|COMP|11067-6|LNCICU|Bleeding Time|Bleeding time
C0363933|T201|COMP|1799-6|LNCICU|Amylase, Urine|Amylase
C0364204|T201|COMP|2072-7|LNCICU|Chloride, Body Fluid|Chloride
C1316698|T201|COMP|34235-2|LNCICU|Amylase/Creatinine Ratio, Urine|Amylase/Creatinine
C0801313|T201|COMP|18267-5|LNCICU|CD16/56|Cells.CD16+CD56+/100 cells
C0364488|T201|COMP|2348-1|LNCICU|Glucose, Joint Fluid|Glucose
C0943515|T201|COMP|27820-0|LNCICU|Protein C, Antigen|Protein C Ag actual/Normal
C1114256|T201|COMP|30398-2|LNCICU|Hematocrit, CSF|Hematocrit
C1977102|T201|COMP|49790-9|LNCICU|Sodium, Ascites|Sodium
C0364325|T201|COMP|2191-5|LNCICU|DHEA-Sulfate|Dehydroepiandrosterone sulfate
C1315830|T201|COMP|33361-7|LNCICU|Bands|Neutrophils.band form/100 leukocytes
C0550247|T201|COMP|11211-0|LNCICU|Bicarbonate, Other Fluid|Carbon dioxide
C0797228|T201|COMP|14040-0|LNCICU|Bicarbonate, Stool|Carbon dioxide
C1114282|T201|COMP|30429-5|LNCICU|Mesothelial cells|Mesothelial cells/100 leukocytes
C0482612|T201|COMP|3188-0|LNCICU|Factor IX|Coagulation factor IX activity
C1977612|T201|COMP|49789-1|LNCICU|Potassium, Ascites|Potassium
C1953453|T201|COMP|48068-1|LNCICU|Heinz Body Prep|Heinz bodies
C1979108|T201|COMP|51238-4|LNCICU|CD13|Cells.CD13/100 cells
C0800302|T201|COMP|17175-1|LNCICU|CD55|Cells.CD55/100 cells
C0800304|T201|COMP|17177-7|LNCICU|CD59|Cells.CD59/100 cells
C0363880|T201|COMP|1746-7|LNCICU|<Albumin>|Albumin
C1315835|T201|COMP|33366-6|LNCICU|Chloride, Ascites|Chloride
C0799717|T201|COMP|16570-4|LNCICU|Centromere|Centromere Ab
C0801314|T201|COMP|18268-3|LNCICU|CD16/56|Cells.CD16+CD56+/100 cells
C2707103|T201|COMP|54360-3|LNCICU|Bicarbonate, Ascites|Bicarbonate
C2735791|T201|COMP|57424-4|LNCICU|CD56|Cells.CD56/100 cells
C1315195|T201|COMP|32724-7|LNCICU|Trichomonas|Trichomonas sp
C0364951|T201|COMP|2809-2|LNCICU|Porphobilinogen Screen|Porphobilinogen
C0482772|T201|COMP|3289-6|LNCICU|Factor II|Prothrombin.activity actual/Normal
C0365030|T201|COMP|2886-0|LNCICU|Total Protein, Joint Fluid|Protein
C1114228|T201|COMP|30366-9|LNCICU|Metamyelocytes|Metamyelocytes/100 leukocytes
C0801528|T201|COMP|18487-9|LNCICU|Broad Casts|Broad casts
C0485107|T201|COMP|6864-3|LNCICU|Sickle Cell Preparation|Hemoglobin S
C0363003|T201|COMP|801-1|LNCICU|Sickle Cells|Sickle cells
C1315834|T201|COMP|33365-8|LNCICU|Mesothelial Cells|Mesothelial cells/100 leukocytes
C1627310|T201|COMP|42867-2|LNCICU|CD117|Cells.CD117/100 cells
C0482649|T201|COMP|3226-8|LNCICU|Factor XI|Coagulation factor XI activity actual/Normal
C1979297|T201|COMP|51232-7|LNCICU|CD11c|Cells.CD11c/100 cells
C1979337|T201|COMP|51294-7|LNCICU|CD33|Cells.CD33/100 cells
C0364155|T201|COMP|2023-0|LNCICU|pCO2, Body Fluid|Carbon dioxide
C1628443|T201|COMP|42871-4|LNCICU|CD138|Cells.CD138/100 cells
C1831457|T201|COMP|47413-0|LNCICU|Plasma|Plasma cells/100 leukocytes
C1979304|T201|COMP|51252-5|LNCICU|CD15|Cells.CD15/100 cells
C0367999|T201|COMP|5775-2|LNCICU|Calcium Phosphate Crystals|Calcium phosphate crystals
C0484865|T201|COMP|6683-7|LNCICU|Reptilase Time|Coagulation reptilase induced
C1979406|T201|COMP|51366-3|LNCICU|CD64|Cells.CD64/100 cells
C0367802|T201|COMP|5644-0|LNCICU|Ethanol, Urine|Ethanol
C0484538|T201|COMP|8115-8|LNCICU|CD16|Cells.CD16/100 cells
C0551499|T201|COMP|12454-5|LNCICU|Ammonium Biurate|Urate crystals.amorphous
C1979300|T201|COMP|51248-3|LNCICU|CD14|Cells.CD14/100 cells
C0942849|T201|COMP|26969-6|LNCICU|Anti-Parietal Cell Antibody|Parietal cell Ab
C1315840|T201|COMP|33371-6|LNCICU|Atypical Lymphocytes|Lymphocytes.variant/100 leukocytes
C0797568|T201|COMP|14388-3|LNCICU|Amylase, Joint Fluid|Amylase
C0482663|T201|COMP|3240-9|LNCICU|Factor XIII|Coagulation factor XIII coagulum dissolution
C0485371|T201|COMP|7893-1|LNCICU|Anti-Gliadin Antibody, IgA|Gliadin Ab
C0482655|T201|COMP|3232-6|LNCICU|Factor XII|Coagulation factor XII activity actual/Normal
C0368062|T201|COMP|5812-3|LNCICU|Sulfonamides|Sulfonamide crystals
C0484552|T201|COMP|8126-5|LNCICU|CD38|Cells.CD38/100 cells
C0550555|T201|COMP|12265-5|LNCICU|Urea Nitrogen, Ascites|Urea nitrogen
C0800908|T201|COMP|17801-2|LNCICU|Metamyelocytes|Metamyelocytes/100 leukocytes
C1979307|T201|COMP|51255-8|LNCICU|CD16/56|Cells.CD16+CD56+/100 cells
C0550455|T201|COMP|12242-4|LNCICU|Phosphate, Body Fluid|Phosphate
C0363849|T201|COMP|1715-2|LNCICU|Acid Phosphatase|Acid phosphatase
C1953414|T201|COMP|48040-0|LNCICU|NRBC|Erythrocytes.nucleated/100 leukocytes
C1979342|T201|COMP|51299-6|LNCICU|CD38|Cells.CD38/100 cells
C1114298|T201|COMP|30447-7|LNCICU|Myelocytes|Myelocytes/100 leukocytes
C1979366|T201|COMP|51320-0|LNCICU|CD41|Cells.CD41/100 cells
C2735793|T201|COMP|57426-9|LNCICU|CD71|Cells.CD71/100 cells
C0797579|T201|COMP|14401-4|LNCICU|Creatinine, Joint Fluid|Creatinine
C0798383|T201|COMP|15212-4|LNCICU|Lipase, Body Fluid|Triacylglycerol lipase
C0800910|T201|COMP|17803-8|LNCICU|Plasma|Plasma cells/100 leukocytes
C0800940|T201|COMP|17833-5|LNCICU|Basophils|Basophils/100 leukocytes
C0364675|T201|COMP|2533-8|LNCICU|LD, Joint Fluid|Lactate dehydrogenase
C0942417|T201|COMP|26447-3|LNCICU|Blasts|Blasts/100 leukocytes
C0364849|T201|COMP|2706-0|LNCICU|pO2, Body Fluid|Oxygen
C0365086|T201|COMP|2942-1|LNCICU|Sex Hormone Binding Globulin|Sex hormone binding globulin
C1315193|T201|COMP|32722-1|LNCICU|Lipase, Ascites|Triacylglycerol lipase
C0366812|T201|COMP|4576-5|LNCICU|Fetal Hemoglobin|Hemoglobin F/Hemoglobin.total
C2735798|T201|COMP|57430-1|LNCICU|Glyco A|Cells.CD235a/100 cells
C0550266|T201|COMP|12183-0|LNCICU|Cholesterol, Body Fluid|Cholesterol
C0797205|T201|COMP|14017-8|LNCICU|CD22|Cells.CD22/100 cells
C0798371|T201|COMP|15200-9|LNCICU|Osmolality, Body Fluid|Osmolality
C0482628|T201|COMP|3204-5|LNCICU|Factor VIII Inhibitor|Coagulation factor VIII inhibitor
C0944827|T201|COMP|29365-4|LNCICU|Magnesium, Body Fluid|Magnesium
C1629585|T201|COMP|42875-5|LNCICU|CD22|Cells.CD22/100 cells
C0797618|T201|COMP|14441-0|LNCICU|Cholesterol, Ascites|Cholesterol
C0801312|T201|COMP|18266-7|LNCICU|CD4/CD8 Ratio|Cells.CD3+CD4+/Cells.CD3+CD8+
C2598765|T201|COMP|53627-6|LNCICU|Chloride, Pleural|Chloride
C0367990|T201|COMP|5773-7|LNCICU|Calcium Carbonate Crystals|Calcium carbonate crystals
C0798326|T201|COMP|15155-5|LNCICU|Calcium, Body Fluid|Calcium
C0800907|T201|COMP|17800-4|LNCICU|Myelocytes|Myelocytes/100 leukocytes
C0484987|T201|COMP|6694-4|LNCICU|Quinidine|quiNIDine
C0800916|T201|COMP|17809-5|LNCICU|Hematocrit|Hematocrit
C0368001|T201|COMP|5777-8|LNCICU|Cholesterol Crystals|Cholesterol crystals
C0797381|T201|COMP|14196-0|LNCICU|Reticulocyte Count, Absolute|Reticulocytes
C0942446|T201|COMP|26484-6|LNCICU|Monocyte Count|Monocytes
C1147726|T201|COMP|32042-4|LNCICU|ANTI-MC|Thyroperoxidase Ab
C1627311|T201|COMP|42869-8|LNCICU|CD138|Cells.CD138/100 cells
C1979286|T201|COMP|51221-0|LNCICU|CD103|Cells.CD103/100 cells
C2707104|T201|COMP|54361-1|LNCICU|Bicarbonate, Pleural|Bicarbonate
C0368006|T201|COMP|5782-8|LNCICU|Cysteine Crystals|Crystals
C0550517|T201|COMP|12260-6|LNCICU|Sugar Water Test|Sucrose hemolysis
C0800906|T201|COMP|17799-8|LNCICU|Promyelocytes|Promyelocytes/100 leukocytes
C0364106|T201|COMP|1973-7|LNCICU|Bilirubin, Total, CSF|Bilirubin
C1369827|T201|COMP|34964-7|LNCICU|Osmotic Fragility|Osmotic fragility
C0368075|T201|COMP|5815-6|LNCICU|Tyrosine Crystals|Tyrosine crystals
C0364834|T201|COMP|2691-4|LNCICU|Osmolality, Ascites|Osmolality
C1977722|T201|COMP|51344-0|LNCICU|CD55|Cells.CD55/100 cells
C1979398|T201|COMP|51358-0|LNCICU|CD59|Cells.CD59/100 cells
C0368033|T201|COMP|5798-4|LNCICU|Leucine Crystals|Leucine crystals
C0942467|T201|COMP|26506-6|LNCICU|Hypersegmented Neutrophils|Neutrophils.segmented/100 leukocytes
C1643606|T201|COMP|41865-7|LNCICU|Hyphenated Yeast|Yeast.hyphae
