C0551559|T102|strict|11488-4|LNC|Consult note|Consult note
C0551559|T102|strict|34099-2|LNC|Cardiology Consult note|Cardiology Consult note
C0551559|T102|strict|34756-7|LNC|Dentistry Consult note|Dentistry Consult note
C0551559|T102|strict|34758-3|LNC|Dermatology Consult note|Dermatology Consult note
C0551559|T102|strict|34760-9|LNC|Diabetology Consult note|Diabetology Consult note
C0551559|T102|strict|34879-7|LNC|Endocrinology Consult note|Endocrinology Consult note
C0551559|T102|strict|34761-7|LNC|Gastroenterology Consult note|Gastroenterology Consult note
C0551559|T102|strict|34764-1|LNC|General Medicine Consult note|General Medicine Consult note
C0551559|T102|strict|34776-5|LNC|Gerontology Consult note|Gerontology Consult note
C0551559|T102|strict|34779-9|LNC|Hematology + Medical Oncology Consult note|Hematology + Medical Oncology Consult note
C0551559|T102|strict|34781-5|LNC|Infectious Disease Consult note|Infectious Disease Consult note
C0551559|T102|strict|72555-6|LNC|Interventional Radiology Consult note|Interventional Radiology Consult note
C0551559|T102|strict|34783-1|LNC|Kinesiotherapy Consult note|Kinesiotherapy Consult note
C0551559|T102|strict|34785-6|LNC|Mental Health Consult note|Mental Health Consult note
C0551559|T102|strict|34795-5|LNC|Nephrology Consult note|Nephrology Consult note
C0551559|T102|strict|34798-9|LNC|Neurological Surgery Consult note|Neurological Surgery Consult note
C0551559|T102|strict|34797-1|LNC|Neurology Consult note|Neurology Consult note
C0551559|T102|strict|34800-3|LNC|Nutrition and Dietetics Consult note|Nutrition and Dietetics Consult note
C0551559|T102|strict|34777-3|LNC|Obstetrics and Gynecology Consult note|Obstetrics and Gynecology Consult note
C0551559|T102|strict|34803-7|LNC|Occupational Health Consult note|Occupational Health Consult note
C0551559|T102|strict|34855-7|LNC|Occupational Therapy Consult note|Occupational Therapy Consult note
C0551559|T102|strict|34805-2|LNC|Oncology Consult note|Oncology Consult note
C0551559|T102|strict|34807-8|LNC|Ophthalmology Consult note|Ophthalmology Consult note
C0551559|T102|strict|34810-2|LNC|Optometry Consult note|Optometry Consult note
C0551559|T102|strict|34812-8|LNC|Oromaxillofacial Surgery Consult note|Oromaxillofacial Surgery Consult note
C0551559|T102|strict|34814-4|LNC|Orthopedics Consult note|Orthopedics Consult note
C0551559|T102|strict|34816-9|LNC|Otorhinolaryngology Consult note|Otorhinolaryngology Consult note
C0551559|T102|strict|60570-9|LNC|Pathology Consult note|Pathology Consult note
C0551559|T102|strict|34820-1|LNC|Pharmacy Consult note|Pharmacy Consult note
C0551559|T102|strict|34822-7|LNC|Physical Medicine and Rehabilitation Consult note|Physical Medicine and Rehabilitation Consult note
C0551559|T102|strict|34824-3|LNC|Physical Therapy Consult note|Physical Therapy Consult note
C0551559|T102|strict|34826-8|LNC|Plastic Surgery Consult note|Plastic Surgery Consult note
C0551559|T102|strict|34828-4|LNC|Podiatry Consult note|Podiatry Consult note
C0551559|T102|strict|34788-0|LNC|Psychiatry Consult note|Psychiatry Consult note
C0551559|T102|strict|34791-4|LNC|Psychology Consult note|Psychology Consult note
C0551559|T102|strict|34103-2|LNC|Pulmonary Consult note|Pulmonary Consult note
C0551559|T102|strict|34831-8|LNC|Radiation Oncology Consult note|Radiation Oncology Consult note
C0551559|T102|strict|73575-3|LNC|Radiology Consult note|Radiology Consult note
C0551559|T102|strict|34833-4|LNC|Recreational Therapy Consult note|Recreational Therapy Consult note
C0551559|T102|strict|34835-9|LNC|Rehabilitation Consult note|Rehabilitation Consult note
C0551559|T102|strict|34837-5|LNC|Respiratory Therapy Consult note|Respiratory Therapy Consult note
C0551559|T102|strict|34839-1|LNC|Rheumatology Consult note|Rheumatology Consult note
C0551559|T102|strict|34841-7|LNC|Social Work Consult note|Social Work Consult note
C0551559|T102|strict|34845-8|LNC|Speech-language pathology+Audiology Consult note|Speech-language pathology+Audiology Consult note
C0551559|T102|strict|34847-4|LNC|Surgery Consult note|Surgery Consult note
C0551559|T102|strict|34849-0|LNC|Thoracic surgery Consult note|Thoracic surgery Consult note
C0551559|T102|strict|34851-6|LNC|Urology Consult note|Urology Consult note
C0551559|T102|strict|34853-2|LNC|Vascular surgery Consult note|Vascular surgery Consult note
C0551559|T102|strict|51846-4|LNC|Emergency department Consult note|Emergency department Consult note
C0551559|T102|strict|34104-0|LNC|Hospital Consult note|Hospital Consult note
C0551559|T102|strict|68619-6|LNC|Adolescent medicine Hospital Consult note|Adolescent medicine Hospital Consult note
C0551559|T102|strict|68633-7|LNC|Allergy and immunology Hospital Consult note|Allergy and immunology Hospital Consult note
C0551559|T102|strict|68639-4|LNC|Audiology Hospital Consult note|Audiology Hospital Consult note
C0551559|T102|strict|68486-0|LNC|Cardiovascular disease.medical student Hospital Consult note|Cardiovascular disease.medical student Hospital Consult note
C0551559|T102|strict|68648-5|LNC|Child and adolescent psychiatry Hospital Consult note|Child and adolescent psychiatry Hospital Consult note
C0551559|T102|strict|68651-9|LNC|Clinical biochemical genetics Hospital Consult note|Clinical biochemical genetics Hospital Consult note
C0551559|T102|strict|68661-8|LNC|Clinical genetics Hospital Consult note|Clinical genetics Hospital Consult note
C0551559|T102|strict|64072-2|LNC|Critical care medicine.medical student Hospital Consult note|Critical care medicine.medical student Hospital Consult note
C0551559|T102|strict|68551-1|LNC|Dermatology Hospital Consult note|Dermatology Hospital Consult note
C0551559|T102|strict|68670-9|LNC|Developmental-behavioral pediatrics Hospital Consult note|Developmental-behavioral pediatrics Hospital Consult note
C0551559|T102|strict|64056-5|LNC|General medicine.medical student Hospital Consult note|General medicine.medical student Hospital Consult note
C0551559|T102|strict|68681-6|LNC|Multi-specialty program Hospital Consult note|Multi-specialty program Hospital Consult note
C0551559|T102|strict|68685-7|LNC|Neonatal perinatal medicine Hospital Consult note|Neonatal perinatal medicine Hospital Consult note
C0551559|T102|strict|68694-9|LNC|Neurological surgery Hospital Consult note|Neurological surgery Hospital Consult note
C0551559|T102|strict|68705-3|LNC|Neurology with special qualifications in child neurology Hospital Consult note|Neurology with special qualifications in child neurology Hospital Consult note
C0551559|T102|strict|68566-9|LNC|Obstetrics and Gynecology Hospital Consult note|Obstetrics and Gynecology Hospital Consult note
C0551559|T102|strict|68570-1|LNC|Occupational therapy Hospital Consult note|Occupational therapy Hospital Consult note
C0551559|T102|strict|68575-0|LNC|Ophthalmology Hospital Consult note|Ophthalmology Hospital Consult note
C0551559|T102|strict|68584-2|LNC|Orthopedic surgery Hospital Consult note|Orthopedic surgery Hospital Consult note
C0551559|T102|strict|68716-0|LNC|Pain medicine Hospital Consult note|Pain medicine Hospital Consult note
C0551559|T102|strict|68469-6|LNC|Pastoral care Hospital Consult note|Pastoral care Hospital Consult note
C0551559|T102|strict|68727-7|LNC|Pediatric cardiology Hospital Consult note|Pediatric cardiology Hospital Consult note
C0551559|T102|strict|68892-9|LNC|Pediatric dermatology Hospital Consult note|Pediatric dermatology Hospital Consult note
C0551559|T102|strict|68897-8|LNC|Pediatric endocrinology Hospital Consult note|Pediatric endocrinology Hospital Consult note
C0551559|T102|strict|68746-7|LNC|Pediatric gastroenterology Hospital Consult note|Pediatric gastroenterology Hospital Consult note
C0551559|T102|strict|68757-4|LNC|Pediatric hematology-oncology Hospital Consult note|Pediatric hematology-oncology Hospital Consult note
C0551559|T102|strict|68765-7|LNC|Pediatric infectious diseases Hospital Consult note|Pediatric infectious diseases Hospital Consult note
C0551559|T102|strict|68869-7|LNC|Pediatric nephrology Hospital Consult note|Pediatric nephrology Hospital Consult note
C0551559|T102|strict|68874-7|LNC|Pediatric otolaryngology Hospital Consult note|Pediatric otolaryngology Hospital Consult note
C0551559|T102|strict|68787-1|LNC|Pediatric pulmonology Hospital Consult note|Pediatric pulmonology Hospital Consult note
C0551559|T102|strict|68879-6|LNC|Pediatric rheumatology Hospital Consult note|Pediatric rheumatology Hospital Consult note
C0551559|T102|strict|68802-8|LNC|Pediatric surgery Hospital Consult note|Pediatric surgery Hospital Consult note
C0551559|T102|strict|68864-8|LNC|Pediatric transplant hepatology Hospital Consult note|Pediatric transplant hepatology Hospital Consult note
C0551559|T102|strict|68812-7|LNC|Pediatric urology Hospital Consult note|Pediatric urology Hospital Consult note
C0551559|T102|strict|68821-8|LNC|Pediatrics Hospital Consult note|Pediatrics Hospital Consult note
C0551559|T102|strict|68586-7|LNC|Pharmacy Hospital Consult note|Pharmacy Hospital Consult note
C0551559|T102|strict|68590-9|LNC|Physical therapy Hospital Consult note|Physical therapy Hospital Consult note
C0551559|T102|strict|68597-4|LNC|Plastic surgery Hospital Consult note|Plastic surgery Hospital Consult note
C0551559|T102|strict|68837-4|LNC|Primary care Hospital Consult note|Primary care Hospital Consult note
C0551559|T102|strict|34102-4|LNC|Psychiatry Hospital Consult note|Psychiatry Hospital Consult note
C0551559|T102|strict|64080-5|LNC|Pulmonary disease.medical student Hospital Consult note|Pulmonary disease.medical student Hospital Consult note
C0551559|T102|strict|68846-5|LNC|Speech-language pathology Hospital Consult note|Speech-language pathology Hospital Consult note
C0551559|T102|strict|64068-0|LNC|Surgery medical student Hospital Consult note|Surgery medical student Hospital Consult note
C0551559|T102|strict|64076-3|LNC|Thoracic surgery.medical student Hospital Consult note|Thoracic surgery.medical student Hospital Consult note
C0551559|T102|strict|68852-3|LNC|Transplant surgery Hospital Consult note|Transplant surgery Hospital Consult note
C0551559|T102|strict|34100-8|LNC|Intensive care unit Consult note|Intensive care unit Consult note
C0551559|T102|strict|51854-8|LNC|Long term care facility Consult note|Long term care facility Consult note
C0551559|T102|strict|51845-6|LNC|Outpatient Consult note|Outpatient Consult note
C0551559|T102|strict|34749-2|LNC|Anesthesiology Outpatient Consult note|Anesthesiology Outpatient Consult note
C0551559|T102|strict|34101-6|LNC|General medicine Outpatient Consult note|General medicine Outpatient Consult note
C0551559|T102|relax|11488-4|LNC|Consult|Consult
C0551559|T102|relax|34099-2|LNC|Cardiology Consult|Cardiology Consult
C0551559|T102|relax|34756-7|LNC|Dentistry Consult|Dentistry Consult
C0551559|T102|relax|34758-3|LNC|Dermatology Consult|Dermatology Consult
C0551559|T102|relax|34760-9|LNC|Diabetes Consult|Diabetes Consult
C0551559|T102|relax|34879-7|LNC|Endocrinology Consult|Endocrinology Consult
C0551559|T102|relax|34761-7|LNC|Gastroenterology Consult|Gastroenterology Consult
C0551559|T102|relax|34764-1|LNC|General Medicine Consult|General Medicine Consult
C0551559|T102|relax|34776-5|LNC|Gerontology Consult|Gerontology Consult
C0551559|T102|relax|34779-9|LNC|Hematology Medical Oncology Consult|Hematology Medical Oncology Consult
C0551559|T102|relax|34781-5|LNC|Infectious Disease Consult|Infectious Disease Consult
C0551559|T102|relax|72555-6|LNC|Interventional Radiology Consult|Interventional Radiology Consult
C0551559|T102|relax|34783-1|LNC|Kinesiotherapy Consult|Kinesiotherapy Consult
C0551559|T102|relax|34785-6|LNC|Mental Health Consult|Mental Health Consult
C0551559|T102|relax|34795-5|LNC|Nephrology Consult|Nephrology Consult
C0551559|T102|relax|34798-9|LNC|Neurological Surgery Consult|Neurological Surgery Consult
C0551559|T102|relax|34797-1|LNC|Neurology Consult|Neurology Consult
C0551559|T102|relax|34800-3|LNC|Nutrition and Dietetics Consult|Nutrition and Dietetics Consult
C0551559|T102|relax|34777-3|LNC|Obstetrics and Gynecology Consult|Obstetrics and Gynecology Consult
C0551559|T102|relax|34803-7|LNC|Occupational Health Consult|Occupational Health Consult
C0551559|T102|relax|34855-7|LNC|Occupational Therapy Consult|Occupational Therapy Consult
C0551559|T102|relax|34805-2|LNC|Oncology Consult|Oncology Consult
C0551559|T102|relax|34807-8|LNC|Ophthalmology Consult|Ophthalmology Consult
C0551559|T102|relax|34810-2|LNC|Optometry Consult|Optometry Consult
C0551559|T102|relax|34812-8|LNC|Oromaxillofacial Surgery Consult|Oromaxillofacial Surgery Consult
C0551559|T102|relax|34814-4|LNC|Orthopedics Consult|Orthopedics Consult
C0551559|T102|relax|34816-9|LNC|Otorhinolaryngology Consult|Otorhinolaryngology Consult
C0551559|T102|relax|60570-9|LNC|Pathology Consult|Pathology Consult
C0551559|T102|relax|34820-1|LNC|Pharmacy Consult|Pharmacy Consult
C0551559|T102|relax|34822-7|LNC|Physical Medicine and Rehabilitation Consult|Physical Medicine and Rehabilitation Consult
C0551559|T102|relax|34824-3|LNC|Physical Therapy Consult|Physical Therapy Consult
C0551559|T102|relax|34826-8|LNC|Plastic Surgery Consult|Plastic Surgery Consult
C0551559|T102|relax|34828-4|LNC|Podiatry Consult|Podiatry Consult
C0551559|T102|relax|34788-0|LNC|Psychiatry Consult|Psychiatry Consult
C0551559|T102|relax|34791-4|LNC|Psychology Consult|Psychology Consult
C0551559|T102|relax|34103-2|LNC|Pulmonary Consult|Pulmonary Consult
C0551559|T102|relax|34831-8|LNC|Radiation Oncology Consult|Radiation Oncology Consult
C0551559|T102|relax|73575-3|LNC|Radiology Consult|Radiology Consult
C0551559|T102|relax|34833-4|LNC|Recreational Therapy Consult|Recreational Therapy Consult
C0551559|T102|relax|34835-9|LNC|Rehabilitation Consult|Rehabilitation Consult
C0551559|T102|relax|34837-5|LNC|Respiratory Therapy Consult|Respiratory Therapy Consult
C0551559|T102|relax|34839-1|LNC|Rheumatology Consult|Rheumatology Consult
C0551559|T102|relax|34841-7|LNC|Social Work Consult|Social Work Consult
C0551559|T102|relax|34845-8|LNC|Speech-language pathology+Audiology Consult|Speech-language pathology+Audiology Consult
C0551559|T102|relax|34847-4|LNC|Surgery Consult|Surgery Consult
C0551559|T102|relax|34849-0|LNC|Thoracic surgery Consult|Thoracic surgery Consult
C0551559|T102|relax|34851-6|LNC|Urology Consult|Urology Consult
C0551559|T102|relax|34853-2|LNC|Vascular surgery Consult|Vascular surgery Consult
C0551559|T102|relax|51846-4|LNC|Emergency department Consult|Emergency department Consult
C0551559|T102|relax|34104-0|LNC|Hospital Consult|Hospital Consult
C0551559|T102|relax|68619-6|LNC|Adolescent medicine Hospital Consult|Adolescent medicine Hospital Consult
C0551559|T102|relax|68633-7|LNC|Allergy and immunology Hospital Consult|Allergy and immunology Hospital Consult
C0551559|T102|relax|68639-4|LNC|Audiology Hospital Consult|Audiology Hospital Consult
C0551559|T102|relax|68486-0|LNC|Cardiovascular disease.medical student Hospital Consult|Cardiovascular disease.medical student Hospital Consult
C0551559|T102|relax|68648-5|LNC|Child and adolescent psychiatry Hospital Consult|Child and adolescent psychiatry Hospital Consult
C0551559|T102|relax|68651-9|LNC|Clinical biochemical genetics Hospital Consult|Clinical biochemical genetics Hospital Consult
C0551559|T102|relax|68661-8|LNC|Clinical genetics Hospital Consult|Clinical genetics Hospital Consult
C0551559|T102|relax|64072-2|LNC|Critical care medicine.medical student Hospital Consult|Critical care medicine.medical student Hospital Consult
C0551559|T102|relax|68551-1|LNC|Dermatology Hospital Consult|Dermatology Hospital Consult
C0551559|T102|relax|68670-9|LNC|Developmental-behavioral pediatrics Hospital Consult|Developmental-behavioral pediatrics Hospital Consult
C0551559|T102|relax|64056-5|LNC|General medicine.medical student Hospital Consult|General medicine.medical student Hospital Consult
C0551559|T102|relax|68681-6|LNC|Multi-specialty program Hospital Consult|Multi-specialty program Hospital Consult
C0551559|T102|relax|68685-7|LNC|Neonatal perinatal medicine Hospital Consult|Neonatal perinatal medicine Hospital Consult
C0551559|T102|relax|68694-9|LNC|Neurological surgery Hospital Consult|Neurological surgery Hospital Consult
C0551559|T102|relax|68705-3|LNC|Neurology with special qualifications in child neurology Hospital Consult|Neurology with special qualifications in child neurology Hospital Consult
C0551559|T102|relax|68566-9|LNC|Obstetrics and Gynecology Hospital Consult|Obstetrics and Gynecology Hospital Consult
C0551559|T102|relax|68570-1|LNC|Occupational therapy Hospital Consult|Occupational therapy Hospital Consult
C0551559|T102|relax|68575-0|LNC|Ophthalmology Hospital Consult|Ophthalmology Hospital Consult
C0551559|T102|relax|68584-2|LNC|Orthopedic surgery Hospital Consult|Orthopedic surgery Hospital Consult
C0551559|T102|relax|68716-0|LNC|Pain medicine Hospital Consult|Pain medicine Hospital Consult
C0551559|T102|relax|68469-6|LNC|Pastoral care Hospital Consult|Pastoral care Hospital Consult
C0551559|T102|relax|68727-7|LNC|Pediatric cardiology Hospital Consult|Pediatric cardiology Hospital Consult
C0551559|T102|relax|68892-9|LNC|Pediatric dermatology Hospital Consult|Pediatric dermatology Hospital Consult
C0551559|T102|relax|68897-8|LNC|Pediatric endocrinology Hospital Consult|Pediatric endocrinology Hospital Consult
C0551559|T102|relax|68746-7|LNC|Pediatric gastroenterology Hospital Consult|Pediatric gastroenterology Hospital Consult
C0551559|T102|relax|68757-4|LNC|Pediatric hematology-oncology Hospital Consult|Pediatric hematology-oncology Hospital Consult
C0551559|T102|relax|68765-7|LNC|Pediatric infectious diseases Hospital Consult|Pediatric infectious diseases Hospital Consult
C0551559|T102|relax|68869-7|LNC|Pediatric nephrology Hospital Consult|Pediatric nephrology Hospital Consult
C0551559|T102|relax|68874-7|LNC|Pediatric otolaryngology Hospital Consult|Pediatric otolaryngology Hospital Consult
C0551559|T102|relax|68787-1|LNC|Pediatric pulmonology Hospital Consult|Pediatric pulmonology Hospital Consult
C0551559|T102|relax|68879-6|LNC|Pediatric rheumatology Hospital Consult|Pediatric rheumatology Hospital Consult
C0551559|T102|relax|68802-8|LNC|Pediatric surgery Hospital Consult|Pediatric surgery Hospital Consult
C0551559|T102|relax|68864-8|LNC|Pediatric transplant hepatology Hospital Consult|Pediatric transplant hepatology Hospital Consult
C0551559|T102|relax|68812-7|LNC|Pediatric urology Hospital Consult|Pediatric urology Hospital Consult
C0551559|T102|relax|68821-8|LNC|Pediatrics Hospital Consult|Pediatrics Hospital Consult
C0551559|T102|relax|68586-7|LNC|Pharmacy Hospital Consult|Pharmacy Hospital Consult
C0551559|T102|relax|68590-9|LNC|Physical therapy Hospital Consult|Physical therapy Hospital Consult
C0551559|T102|relax|68597-4|LNC|Plastic surgery Hospital Consult|Plastic surgery Hospital Consult
C0551559|T102|relax|68837-4|LNC|Primary care Hospital Consult|Primary care Hospital Consult
C0551559|T102|relax|34102-4|LNC|Psychiatry Hospital Consult|Psychiatry Hospital Consult
C0551559|T102|relax|64080-5|LNC|Pulmonary disease.medical student Hospital Consult|Pulmonary disease.medical student Hospital Consult
C0551559|T102|relax|68846-5|LNC|Speech-language pathology Hospital Consult|Speech-language pathology Hospital Consult
C0551559|T102|relax|64068-0|LNC|Surgery medical student Hospital Consult|Surgery medical student Hospital Consult
C0551559|T102|relax|64076-3|LNC|Thoracic surgery.medical student Hospital Consult|Thoracic surgery.medical student Hospital Consult
C0551559|T102|relax|68852-3|LNC|Transplant surgery Hospital Consult|Transplant surgery Hospital Consult
C0551559|T102|relax|34100-8|LNC|Intensive care unit Consult|Intensive care unit Consult
C0551559|T102|relax|51854-8|LNC|Long term care facility Consult|Long term care facility Consult
C0551559|T102|relax|51845-6|LNC|Outpatient Consult|Outpatient Consult
C0551559|T102|relax|34749-2|LNC|Anesthesiology Outpatient Consult|Anesthesiology Outpatient Consult
C0551559|T102|relax|34101-6|LNC|General medicine Outpatient Consult|General medicine Outpatient Consult
C0801840|T102|strict|18842-5|LNC|Discharge summary|Discharge summary
C0801840|T102|strict|11490-0|LNC|Physician Discharge summary|Physician Discharge summary
C0801840|T102|strict|28655-9|LNC|Physician attending Discharge summary|Physician attending Discharge summary
C0801840|T102|strict|29761-4|LNC|Dentist Discharge summary|Dentist Discharge summary
C0801840|T102|strict|34745-0|LNC|Nurse Discharge summary|Nurse Discharge summary
C0801840|T102|strict|34105-7|LNC|Hospital Discharge summary|Hospital Discharge summary
C0801840|T102|strict|34106-5|LNC|Physician Hospital Discharge summary|Physician Hospital Discharge summary
C1316580|T102|strict|34117-2|LNC|History and physical note|History and physical note
C1316580|T102|strict|11492-6|LNC|Provider-unspecified, History and physical note|Provider-unspecified, History and physical note
C1316580|T102|strict|28626-0|LNC|Physician History and physical note|Physician History and physical note
C1316580|T102|strict|34774-0|LNC|Surgery History and physical note|Surgery History and physical note
C1316580|T102|strict|34115-6|LNC|Medical student Hospital History and physical note|Medical student Hospital History and physical note
C1316580|T102|strict|34116-4|LNC|Physician Nursing facility History and physical note|Physician Nursing facility History and physical note
C1316580|T102|strict|34095-0|LNC|Comprehensive history and physical note|Comprehensive history and physical note
C1316580|T102|strict|34096-8|LNC|Nursing facility Comprehensive history and physical note|Nursing facility Comprehensive history and physical note
C1316580|T102|strict|51849-8|LNC|Admission history and physical note|Admission history and physical note
C1316580|T102|strict|47039-3|LNC|Hospital Admission history and physical note|Hospital Admission history and physical note
C1316580|T102|strict|34763-3|LNC|General medicine Admission history and physical note|General medicine Admission history and physical note
C1316580|T102|strict|34094-3|LNC|Cardiology Hospital Admission history and physical note|Cardiology Hospital Admission history and physical note
C1316580|T102|strict|34138-8|LNC|Targeted history and physical note|Targeted history and physical note
C1316580|T102|relax|34117-2|LNC|History and physical|History and physical
C1316580|T102|relax|11492-6|LNC|Provider History and physical|Provider History and physical
C1316580|T102|relax|28626-0|LNC|Physician History and physical|Physician History and physical
C1316580|T102|relax|34774-0|LNC|Surgery History and physical|Surgery History and physical
C1316580|T102|relax|34115-6|LNC|Medical student Hospital History and physical|Medical student Hospital History and physical
C1316580|T102|relax|34116-4|LNC|Physician Nursing facility History and physical|Physician Nursing facility History and physical
C1316580|T102|relax|34095-0|LNC|Comprehensive history and physical|Comprehensive history and physical
C1316580|T102|relax|34096-8|LNC|Nursing facility Comprehensive history and physical|Nursing facility Comprehensive history and physical
C1316580|T102|relax|51849-8|LNC|Admission history and physical|Admission history and physical
C1316580|T102|relax|47039-3|LNC|Hospital Admission history and physical|Hospital Admission history and physical
C1316580|T102|relax|34763-3|LNC|General medicine Admission history and physical|General medicine Admission history and physical
C1316580|T102|relax|34094-3|LNC|Cardiology Hospital Admission history and physical|Cardiology Hospital Admission history and physical
C1316580|T102|relax|34138-8|LNC|Targeted history and physical|Targeted history and physical
C3483153|T102|strict|81192-7|LNC|Clinical pathology Consult note|Clinical pathology Consult note
C3483153|T102|strict|90010-0|LNC|Clinical pathology procedure note|Clinical pathology procedure note
C3483153|T102|strict|90011-8|LNC|Clinical pathology Progress note|Clinical pathology Progress note
C3483153|T102|strict|90013-4|LNC|Clinical pathology Initial evaluation note|Clinical pathology Initial evaluation note
C3483153|T102|strict|90015-9|LNC|Clinical pathology Telephone encounter Note|Clinical pathology Telephone encounter Note
C3483153|T102|strict|90371-6|LNC|Clinical pathology Note|Clinical pathology Note
C3483153|T102|relax|60570-9|LNC|Pathology Consult note|Pathology Consult note
C3483153|T102|relax|81192-7|LNC|pathology Consult note|pathology Consult note
C3483153|T102|relax|90010-0|LNC|pathology procedure note|pathology procedure note
C3483153|T102|relax|90011-8|LNC|pathology Progress note|pathology Progress note
C3483153|T102|relax|90013-4|LNC|pathology Initial evaluation note|pathology Initial evaluation note
C3483153|T102|relax|90015-9|LNC|pathology Telephone encounter|pathology Telephone encounter
C3483153|T102|relax|90371-6|LNC|pathology report|pathology report
C3853717|T102|strict|28570-0|LNC|Provider-unspecified Procedure note|Provider-unspecified Procedure note
C3853717|T102|strict|11505-5|LNC|Physician procedure note|Physician procedure note
C3853717|T102|strict|18744-3|LNC|Bronchoscopy study|Bronchoscopy study
C3853717|T102|strict|18745-0|LNC|Cardiac catheterization study|Cardiac catheterization study
C3853717|T102|strict|18746-8|LNC|Colonoscopy study|Colonoscopy study
C3853717|T102|strict|18751-8|LNC|Endoscopy study|Endoscopy study
C3853717|T102|strict|18753-4|LNC|Flexible sigmoidoscopy study|Flexible sigmoidoscopy study
C3853717|T102|strict|18836-7|LNC|Cardiac stress study Procedure|Cardiac stress study Procedure
C3853717|T102|strict|28577-5|LNC|Dentist procedure note|Dentist procedure note
C3853717|T102|strict|28625-2|LNC|Podiatry procedure note|Podiatry procedure note
C3853717|T102|strict|29757-2|LNC|Colposcopy study|Colposcopy study
C3853717|T102|strict|33721-2|LNC|Bone marrow Pathology biopsy report|Bone marrow Pathology biopsy report
C3853717|T102|strict|34121-4|LNC|Interventional procedure note|Interventional procedure note
C3853717|T102|strict|34896-1|LNC|Cardiovascular disease Interventional procedure note|Cardiovascular disease Interventional procedure note
C3853717|T102|strict|34899-5|LNC|Gastroenterology Interventional procedure note|Gastroenterology Interventional procedure note
C3853717|T102|strict|47048-4|LNC|Diagnostic interventional study report Interventional radiology|Diagnostic interventional study report Interventional radiology
C3853717|T102|strict|48807-2|LNC|Bone marrow aspiration report|Bone marrow aspiration report
C3853717|T102|relax|28570-0|LNC|Provider Procedure|Provider Procedure
C3853717|T102|relax|11505-5|LNC|Physician procedure|Physician procedure
C3853717|T102|relax|18745-0|LNC|Cardiac catheterization|Cardiac catheterization
C3853717|T102|relax|18746-8|LNC|Colonoscopy|Colonoscopy
C3853717|T102|relax|18751-8|LNC|Endoscopy|Endoscopy
C3853717|T102|relax|18753-4|LNC|Flexible sigmoidoscopy|Flexible sigmoidoscopy
C3853717|T102|relax|18836-7|LNC|Cardiac stress study|Cardiac stress study
C3853717|T102|relax|28577-5|LNC|Dentist procedure|Dentist procedure
C3853717|T102|relax|28625-2|LNC|Podiatry procedure|Podiatry procedure
C3853717|T102|relax|29757-2|LNC|Colposcopy|Colposcopy
C3853717|T102|relax|33721-2|LNC|Bone marrow biopsy|Bone marrow biopsy
C3853717|T102|relax|34121-4|LNC|Interventional procedure|Interventional procedure
C3853717|T102|relax|34896-1|LNC|Cardiovascular disease Interventional procedure|Cardiovascular disease Interventional procedure
C3853717|T102|relax|34899-5|LNC|Gastroenterology Interventional procedure|Gastroenterology Interventional procedure
C3853717|T102|relax|47048-4|LNC|Interventional radiology|Interventional radiology
C3853717|T102|relax|48807-2|LNC|Bone marrow aspiration|Bone marrow aspiration
C0551633|T102|strict|11506-3|LNC|Provider-unspecified Progress note|Provider-unspecified Progress note
C0551633|T102|strict|18733-6|LNC|Physician attending Progress note|Physician attending Progress note
C0551633|T102|strict|28569-2|LNC|Physician consulting Progress note|Physician consulting Progress note
C0551633|T102|strict|28617-9|LNC|Dentistry Progress note|Dentistry Progress note
C0551633|T102|strict|34900-1|LNC|General medicine Progress note|General medicine Progress note
C0551633|T102|strict|34904-3|LNC|Mental health Progress note|Mental health Progress note
C0551633|T102|strict|28623-7|LNC|Nurse Progress note|Nurse Progress note
C0551633|T102|strict|11507-1|LNC|Occupational therapy Progress note|Occupational therapy Progress note
C0551633|T102|strict|11508-9|LNC|Physical therapy Progress note|Physical therapy Progress note
C0551633|T102|strict|11509-7|LNC|Podiatry Progress note|Podiatry Progress note
C0551633|T102|strict|28627-8|LNC|Psychiatry Progress note|Psychiatry Progress note
C0551633|T102|strict|11510-5|LNC|Psychology Progress note|Psychology Progress note
C0551633|T102|strict|28656-7|LNC|Social work Progress note|Social work Progress note
C0551633|T102|strict|11512-1|LNC|Speech-language pathology Progress note|Speech-language pathology Progress note
C0551633|T102|strict|34126-3|LNC|Intensive care unit Progress note|Intensive care unit Progress note
C0551633|T102|strict|15507-7|LNC|Provider-unspecified ED Progress note|Provider-unspecified ED Progress note
C0551633|T102|strict|34129-7|LNC|Patient's home Progress note|Patient's home Progress note
C0551633|T102|strict|34125-5|LNC|Case manager Patient's home Progress note|Case manager Patient's home Progress note
C0551633|T102|strict|34130-5|LNC|Hospital Progress note|Hospital Progress note
C0551633|T102|strict|34131-3|LNC|Outpatient Progress note|Outpatient Progress note
C0551633|T102|strict|34124-8|LNC|Cardiology Outpatient Progress note|Cardiology Outpatient Progress note
C0551633|T102|strict|34127-1|LNC|Dentistry Hygienist Outpatient Progress note|Dentistry Hygienist Outpatient Progress note
C0551633|T102|strict|34128-9|LNC|Dentistry Outpatient Progress note|Dentistry Outpatient Progress note
C0551633|T102|strict|34901-9|LNC|General medicine Outpatient Progress note|General medicine Outpatient Progress note
C0551633|T102|strict|34132-1|LNC|Pharmacy Outpatient Progress note|Pharmacy Outpatient Progress note
C0551633|T102|strict|28580-9|LNC|Chiropractic medicine Progress note|Chiropractic medicine Progress note
C0551633|T102|strict|28575-9|LNC|Nurse practitioner Progress note|Nurse practitioner Progress note
C0551633|T102|relax|11506-3|LNC|Provider Progress|Provider Progress
C0551633|T102|relax|18733-6|LNC|Physician attending Progress|Physician attending Progress
C0551633|T102|relax|28569-2|LNC|Physician consulting Progress|Physician consulting Progress
C0551633|T102|relax|28617-9|LNC|Dentistry Progress|Dentistry Progress
C0551633|T102|relax|34900-1|LNC|General medicine Progress|General medicine Progress
C0551633|T102|relax|34904-3|LNC|Mental health progress|Mental health progress
C0551633|T102|relax|28623-7|LNC|Nurse progress|Nurse progress
C0551633|T102|relax|11507-1|LNC|Occupational therapy progress|Occupational therapy progress
C0551633|T102|relax|11508-9|LNC|Physical therapy progress|Physical therapy progress
C0551633|T102|relax|11509-7|LNC|Podiatry progress|Podiatry progress
C0551633|T102|relax|28627-8|LNC|Psychiatry progress|Psychiatry progress
C0551633|T102|relax|11510-5|LNC|Psychology progress|Psychology progress
C0551633|T102|relax|28656-7|LNC|Social work progress|Social work progress
C0551633|T102|relax|11512-1|LNC|Speech-language pathology progress|Speech-language pathology progress
C0551633|T102|relax|34126-3|LNC|Intensive care unit progress|Intensive care unit progress
C0551633|T102|relax|15507-7|LNC|Provider-unspecified ED progress|Provider-unspecified ED progress
C0551633|T102|relax|34129-7|LNC|Patient's home progress|Patient's home progress
C0551633|T102|relax|34125-5|LNC|Case manager Patient's home progress|Case manager Patient's home progress
C0551633|T102|relax|34130-5|LNC|Hospital progress|Hospital progress
C0551633|T102|relax|34131-3|LNC|Outpatient progress|Outpatient progress
C0551633|T102|relax|34124-8|LNC|Cardiology Outpatient progress|Cardiology Outpatient progress
C0551633|T102|relax|34127-1|LNC|Dentistry Hygienist Outpatient progress|Dentistry Hygienist Outpatient progress
C0551633|T102|relax|34128-9|LNC|Dentistry Outpatient progress|Dentistry Outpatient progress
C0551633|T102|relax|34901-9|LNC|General medicine Outpatient progress|General medicine Outpatient progress
C0551633|T102|relax|34132-1|LNC|Pharmacy Outpatient progress|Pharmacy Outpatient progress
C0551633|T102|relax|28580-9|LNC|Chiropractic medicine progress|Chiropractic medicine progress
C0551633|T102|relax|28575-9|LNC|Nurse practitioner progress|Nurse practitioner progress
C2735498|T102|strict|57133-1|LNC|Referral note|Referral note
C2735498|T102|strict|57170-3|LNC|Cardiovascular disease Referral note|Cardiovascular disease Referral note
C2735498|T102|strict|57178-6|LNC|Critical Care Medicine Referral note|Critical Care Medicine Referral note
C2735498|T102|strict|57134-9|LNC|Dentistry Referral note|Dentistry Referral note
C2735498|T102|strict|57135-6|LNC|Dermatology Referral note|Dermatology Referral note
C2735498|T102|strict|57136-4|LNC|Diabetology Referral note|Diabetology Referral note
C2735498|T102|strict|57137-2|LNC|Endocrinology Referral note|Endocrinology Referral note
C2735498|T102|strict|57138-0|LNC|Gastroenterology Referral note|Gastroenterology Referral note
C2735498|T102|strict|57139-8|LNC|General medicine Referral note|General medicine Referral note
C2735498|T102|strict|57171-1|LNC|Geriatric medicine Referral note|Geriatric medicine Referral note
C2735498|T102|strict|57141-4|LNC|Infectious disease Referral note|Infectious disease Referral note
C2735498|T102|strict|57142-2|LNC|Kinesiotherapy Referral note|Kinesiotherapy Referral note
C2735498|T102|strict|57143-0|LNC|Mental health Referral note|Mental health Referral note
C2735498|T102|strict|57144-8|LNC|Nephrology Referral note|Nephrology Referral note
C2735498|T102|strict|57146-3|LNC|Neurological surgery Referral note|Neurological surgery Referral note
C2735498|T102|strict|57145-5|LNC|Neurology Referral note|Neurology Referral note
C2735498|T102|strict|57173-7|LNC|Nutrition and dietetics Referral note|Nutrition and dietetics Referral note
C2735498|T102|strict|57179-4|LNC|Obstetrics and Gynecology Referral note|Obstetrics and Gynecology Referral note
C2735498|T102|strict|57147-1|LNC|Occupational health Referral note|Occupational health Referral note
C2735498|T102|strict|57148-9|LNC|Occupational therapy Referral note|Occupational therapy Referral note
C2735498|T102|strict|57149-7|LNC|Oncology Referral note|Oncology Referral note
C2735498|T102|strict|57150-5|LNC|Ophthalmology Referral note|Ophthalmology Referral note
C2735498|T102|strict|57151-3|LNC|Optometry Referral note|Optometry Referral note
C2735498|T102|strict|57174-5|LNC|Oral surgery Referral note|Oral surgery Referral note
C2735498|T102|strict|57175-2|LNC|Orthopedic surgery Referral note|Orthopedic surgery Referral note
C2735498|T102|strict|57176-0|LNC|Otolaryngology Referral note|Otolaryngology Referral note
C2735498|T102|strict|57152-1|LNC|Pharmacy Referral note|Pharmacy Referral note
C2735498|T102|strict|57153-9|LNC|Physical medicine and rehabilitation Referral note|Physical medicine and rehabilitation Referral note
C2735498|T102|strict|57154-7|LNC|Physical therapy Referral note|Physical therapy Referral note
C2735498|T102|strict|57155-4|LNC|Plastic surgery Referral note|Plastic surgery Referral note
C2735498|T102|strict|57156-2|LNC|Podiatry Referral note|Podiatry Referral note
C2735498|T102|strict|57157-0|LNC|Psychiatry Referral note|Psychiatry Referral note
C2735498|T102|strict|57158-8|LNC|Psychology Referral note|Psychology Referral note
C2735498|T102|strict|57177-8|LNC|Pulmonary disease Referral note|Pulmonary disease Referral note
C2735498|T102|strict|57159-6|LNC|Radiation oncology Referral note|Radiation oncology Referral note
C2735498|T102|strict|57160-4|LNC|Recreational therapy Referral note|Recreational therapy Referral note
C2735498|T102|strict|57161-2|LNC|Rehabilitation Referral note|Rehabilitation Referral note
C2735498|T102|strict|57162-0|LNC|Respiratory therapy Referral note|Respiratory therapy Referral note
C2735498|T102|strict|57163-8|LNC|Rheumatology Referral note|Rheumatology Referral note
C2735498|T102|strict|57164-6|LNC|Social work Referral note|Social work Referral note
C2735498|T102|strict|57166-1|LNC|Surgery Referral note|Surgery Referral note
C2735498|T102|strict|57167-9|LNC|Thoracic surgery Referral note|Thoracic surgery Referral note
C2735498|T102|strict|57168-7|LNC|Urology Referral note|Urology Referral note
C2735498|T102|strict|57169-5|LNC|Vascular surgery Referral note|Vascular surgery Referral note
C2735498|T102|strict|69438-0|LNC|Forensic medicine Referral note|Forensic medicine Referral note
C2735498|T102|relax|57133-1|LNC|Referral|Referral
C2735498|T102|relax|57170-3|LNC|Cardiovascular disease Referral|Cardiovascular disease Referral
C2735498|T102|relax|57178-6|LNC|Critical Care Medicine Referral|Critical Care Medicine Referral
C2735498|T102|relax|57134-9|LNC|Dentistry Referral|Dentistry Referral
C2735498|T102|relax|57135-6|LNC|Dermatology Referral|Dermatology Referral
C2735498|T102|relax|57136-4|LNC|Diabetology Referral|Diabetology Referral
C2735498|T102|relax|57137-2|LNC|Endocrinology Referral|Endocrinology Referral
C2735498|T102|relax|57138-0|LNC|Gastroenterology Referral|Gastroenterology Referral
C2735498|T102|relax|57139-8|LNC|General medicine Referral|General medicine Referral
C2735498|T102|relax|57171-1|LNC|Geriatric medicine Referral|Geriatric medicine Referral
C2735498|T102|relax|57141-4|LNC|Infectious disease Referral|Infectious disease Referral
C2735498|T102|relax|57142-2|LNC|Kinesiotherapy Referral|Kinesiotherapy Referral
C2735498|T102|relax|57143-0|LNC|Mental health Referral|Mental health Referral
C2735498|T102|relax|57144-8|LNC|Nephrology Referral|Nephrology Referral
C2735498|T102|relax|57146-3|LNC|Neurological surgery Referral|Neurological surgery Referral
C2735498|T102|relax|57145-5|LNC|Neurology Referral|Neurology Referral
C2735498|T102|relax|57173-7|LNC|Nutrition and dietetics Referral|Nutrition and dietetics Referral
C2735498|T102|relax|57179-4|LNC|Obstetrics and Gynecology Referral|Obstetrics and Gynecology Referral
C2735498|T102|relax|57147-1|LNC|Occupational health Referral|Occupational health Referral
C2735498|T102|relax|57148-9|LNC|Occupational therapy Referral|Occupational therapy Referral
C2735498|T102|relax|57149-7|LNC|Oncology Referral|Oncology Referral
C2735498|T102|relax|57150-5|LNC|Ophthalmology Referral|Ophthalmology Referral
C2735498|T102|relax|57151-3|LNC|Optometry Referral|Optometry Referral
C2735498|T102|relax|57174-5|LNC|Oral surgery Referral|Oral surgery Referral
C2735498|T102|relax|57175-2|LNC|Orthopedic surgery Referral|Orthopedic surgery Referral
C2735498|T102|relax|57176-0|LNC|Otolaryngology Referral|Otolaryngology Referral
C2735498|T102|relax|57152-1|LNC|Pharmacy Referral|Pharmacy Referral
C2735498|T102|relax|57153-9|LNC|Physical medicine and rehabilitation Referral|Physical medicine and rehabilitation Referral
C2735498|T102|relax|57154-7|LNC|Physical therapy Referral|Physical therapy Referral
C2735498|T102|relax|57155-4|LNC|Plastic surgery Referral|Plastic surgery Referral
C2735498|T102|relax|57156-2|LNC|Podiatry Referral|Podiatry Referral
C2735498|T102|relax|57157-0|LNC|Psychiatry Referral|Psychiatry Referral
C2735498|T102|relax|57158-8|LNC|Psychology Referral|Psychology Referral
C2735498|T102|relax|57177-8|LNC|Pulmonary disease Referral|Pulmonary disease Referral
C2735498|T102|relax|57159-6|LNC|Radiation oncology Referral|Radiation oncology Referral
C2735498|T102|relax|57160-4|LNC|Recreational therapy Referral|Recreational therapy Referral
C2735498|T102|relax|57161-2|LNC|Rehabilitation Referral|Rehabilitation Referral
C2735498|T102|relax|57162-0|LNC|Respiratory therapy Referral|Respiratory therapy Referral
C2735498|T102|relax|57163-8|LNC|Rheumatology Referral|Rheumatology Referral
C2735498|T102|relax|57164-6|LNC|Social work Referral|Social work Referral
C2735498|T102|relax|57166-1|LNC|Surgery Referral|Surgery Referral
C2735498|T102|relax|57167-9|LNC|Thoracic surgery Referral|Thoracic surgery Referral
C2735498|T102|relax|57168-7|LNC|Urology Referral|Urology Referral
C2735498|T102|relax|57169-5|LNC|Vascular surgery Referral|Vascular surgery Referral
C2735498|T102|relax|69438-0|LNC|Forensic medicine Referral|Forensic medicine Referral
C0551628|T102|strict|11504-8|LNC|Provider-unspecified Operation note|Provider-unspecified Operation note
C0551628|T102|strict|34137-0|LNC|Outpatient Surgical operation note|Outpatient Surgical operation note
C0551628|T102|strict|28583-3|LNC|Dentist Operation note|Dentist Operation note
C0551628|T102|strict|28624-5|LNC|Podiatry Operation note|Podiatry Operation note
C0551628|T102|strict|28573-4|LNC|Physician, Operation note|Physician, Operation note
C0551628|T102|strict|34877-1|LNC|Urology Surgical operation note|Urology Surgical operation note
C0551628|T102|strict|34874-8|LNC|Surgery Surgical operation note|Surgery Surgical operation note
C0551628|T102|strict|34870-6|LNC|Plastic surgery Surgical operation note|Plastic surgery Surgical operation note
C0551628|T102|strict|34868-0|LNC|Orthopaedic surgery Surgical operation note|Orthopaedic surgery Surgical operation note
C0551628|T102|strict|34818-5|LNC|Otolaryngology Surgical operation note|Otolaryngology Surgical operation note
C0551628|T102|relax|11504-8|LNC|Provider Operation|Provider Operation
C0551628|T102|relax|34137-0|LNC|Outpatient Surgical operation|Outpatient Surgical operation
C0551628|T102|relax|28583-3|LNC|Dentist Operation|Dentist Operation
C0551628|T102|relax|28624-5|LNC|Podiatry Operation|Podiatry Operation
C0551628|T102|relax|28573-4|LNC|Physician Operation|Physician Operation
C0551628|T102|relax|34877-1|LNC|Urology Surgical operation|Urology Surgical operation
C0551628|T102|relax|34874-8|LNC|Surgery Surgical operation|Surgery Surgical operation
C0551628|T102|relax|34870-6|LNC|Plastic surgery Surgical operation|Plastic surgery Surgical operation
C0551628|T102|relax|34868-0|LNC|Orthopaedic surgery Surgical operation|Orthopaedic surgery Surgical operation
C0551628|T102|relax|34818-5|LNC|Otolaryngology Surgical operation|Otolaryngology Surgical operation
C1316596|T102|strict|18761-7|LNC|Provider-unspecified Transfer summary|Provider-unspecified Transfer summary
C1316596|T102|strict|68618-8|LNC|Adolescent medicine Transfer summarization note|Adolescent medicine Transfer summarization note
C1316596|T102|strict|68632-9|LNC|Allergy and immunology Transfer summarization note|Allergy and immunology Transfer summarization note
C1316596|T102|strict|68647-7|LNC|Child and adolescent psychiatry Transfer summarization note|Child and adolescent psychiatry Transfer summarization note
C1316596|T102|strict|68660-0|LNC|Clinical genetics Transfer summarization note|Clinical genetics Transfer summarization note
C1316596|T102|strict|34755-9|LNC|Critical Care Medicine Transfer summarization note|Critical Care Medicine Transfer summarization note
C1316596|T102|strict|68669-1|LNC|Developmental-behavioral pediatrics Transfer summarization note|Developmental-behavioral pediatrics Transfer summarization note
C1316596|T102|strict|34770-8|LNC|General medicine Transfer summarization note|General medicine Transfer summarization note
C1316596|T102|strict|68680-8|LNC|Multi-specialty program Transfer summarization note|Multi-specialty program Transfer summarization note
C1316596|T102|strict|68704-6|LNC|Neurology with special qualifications in child neurology Transfer summary note|Neurology with special qualifications in child neurology Transfer summary note
C1316596|T102|strict|28651-8|LNC|Nurse Transfer note|Nurse Transfer note
C1316596|T102|strict|68565-1|LNC|Obstetrics and Gynecology Transfer summarization note|Obstetrics and Gynecology Transfer summarization note
C1316596|T102|strict|68569-3|LNC|Occupational therapy Transfer summarization note|Occupational therapy Transfer summarization note
C1316596|T102|strict|68887-9|LNC|Ophthalmology Transfer summarization note|Ophthalmology Transfer summarization note
C1316596|T102|strict|68583-4|LNC|Orthopedic surgery Transfer summarization note|Orthopedic surgery Transfer summarization note
C1316596|T102|strict|68715-2|LNC|Pain medicine Transfer summarization note|Pain medicine Transfer summarization note
C1316596|T102|strict|68726-9|LNC|Pediatric cardiology Transfer summarization note|Pediatric cardiology Transfer summarization note
C1316596|T102|strict|68737-6|LNC|Pediatric endocrinology Transfer summarization note|Pediatric endocrinology Transfer summarization note
C1316596|T102|strict|68745-9|LNC|Pediatric gastroenterology Transfer summarization note|Pediatric gastroenterology Transfer summarization note
C1316596|T102|strict|68756-6|LNC|Pediatric hematology-oncology Transfer summarization note|Pediatric hematology-oncology Transfer summarization note
C1316596|T102|strict|68764-0|LNC|Pediatric infectious diseases Transfer summarization note|Pediatric infectious diseases Transfer summarization note
C1316596|T102|strict|68772-3|LNC|Pediatric nephrology Transfer summarization note|Pediatric nephrology Transfer summarization note
C1316596|T102|strict|68777-2|LNC|Pediatric otolaryngology Transfer summarization note|Pediatric otolaryngology Transfer summarization note
C1316596|T102|strict|68786-3|LNC|Pediatric pulmonology Transfer summarization note|Pediatric pulmonology Transfer summarization note
C1316596|T102|strict|68793-9|LNC|Pediatric rheumatology Transfer summarization note|Pediatric rheumatology Transfer summarization note
C1316596|T102|strict|68801-0|LNC|Pediatric surgery Transfer summarization note|Pediatric surgery Transfer summarization note
C1316596|T102|strict|68863-0|LNC|Pediatric transplant hepatology Transfer summarization note|Pediatric transplant hepatology Transfer summarization note
C1316596|T102|strict|68811-9|LNC|Pediatric urology Transfer summarization note|Pediatric urology Transfer summarization note
C1316596|T102|strict|68883-8|LNC|Pediatrics Transfer summarization note|Pediatrics Transfer summarization note
C1316596|T102|strict|28616-1|LNC|Physician Transfer note|Physician Transfer note
C1316596|T102|strict|68596-6|LNC|Plastic surgery Transfer summarization note|Plastic surgery Transfer summarization note
C1316596|T102|strict|68482-9|LNC|Nurse Hospital Transfer summarization note|Nurse Hospital Transfer summarization note
C1316596|T102|strict|68884-6|LNC|Pediatrics Hospital Transfer summarization note|Pediatrics Hospital Transfer summarization note
C1316596|T102|relax|18761-7|LNC|Transfer summary|Transfer summary
C1316596|T102|relax|68618-8|LNC|Adolescent medicine Transfer|Adolescent medicine Transfer
C1316596|T102|relax|68632-9|LNC|Allergy and immunology Transfer|Allergy and immunology Transfer
C1316596|T102|relax|68647-7|LNC|Child and adolescent psychiatry Transfer|Child and adolescent psychiatry Transfer
C1316596|T102|relax|68660-0|LNC|Clinical genetics Transfer|Clinical genetics Transfer
C1316596|T102|relax|34755-9|LNC|Critical Care Medicine Transfer|Critical Care Medicine Transfer
C1316596|T102|relax|68669-1|LNC|Developmental-behavioral pediatrics Transfer|Developmental-behavioral pediatrics Transfer
C1316596|T102|relax|34770-8|LNC|General medicine Transfer|General medicine Transfer
C1316596|T102|relax|68680-8|LNC|Multi-specialty program Transfer|Multi-specialty program Transfer
C1316596|T102|relax|68704-6|LNC|Neurology Transfer summary|Neurology Transfer summary
C1316596|T102|relax|28651-8|LNC|Nurse Transfer note|Nurse Transfer note
C1316596|T102|relax|68565-1|LNC|Obstetrics and Gynecology Transfer|Obstetrics and Gynecology Transfer
C1316596|T102|relax|68569-3|LNC|Occupational therapy Transfer|Occupational therapy Transfer
C1316596|T102|relax|68887-9|LNC|Ophthalmology Transfer|Ophthalmology Transfer
C1316596|T102|relax|68583-4|LNC|Orthopedic surgery Transfer|Orthopedic surgery Transfer
C1316596|T102|relax|68715-2|LNC|Pain medicine Transfer|Pain medicine Transfer
C1316596|T102|relax|68726-9|LNC|Pediatric cardiology Transfer|Pediatric cardiology Transfer
C1316596|T102|relax|68737-6|LNC|Pediatric endocrinology Transfer|Pediatric endocrinology Transfer
C1316596|T102|relax|68745-9|LNC|Pediatric gastroenterology Transfer|Pediatric gastroenterology Transfer
C1316596|T102|relax|68756-6|LNC|Pediatric hematology oncology Transfer|Pediatric hematology oncology Transfer
C1316596|T102|relax|68764-0|LNC|Pediatric infectious diseases Transfer|Pediatric infectious diseases Transfer
C1316596|T102|relax|68772-3|LNC|Pediatric nephrology Transfer|Pediatric nephrology Transfer
C1316596|T102|relax|68777-2|LNC|Pediatric otolaryngology Transfer|Pediatric otolaryngology Transfer
C1316596|T102|relax|68786-3|LNC|Pediatric pulmonology Transfer|Pediatric pulmonology Transfer
C1316596|T102|relax|68793-9|LNC|Pediatric rheumatology Transfer|Pediatric rheumatology Transfer
C1316596|T102|relax|68801-0|LNC|Pediatric surgery Transfer|Pediatric surgery Transfer
C1316596|T102|relax|68863-0|LNC|Pediatric transplant hepatology Transfer|Pediatric transplant hepatology Transfer
C1316596|T102|relax|68811-9|LNC|Pediatric urology Transfer|Pediatric urology Transfer
C1316596|T102|relax|68883-8|LNC|Pediatrics Transfer|Pediatrics Transfer
C1316596|T102|relax|28616-1|LNC|Physician Transfer note|Physician Transfer note
C1316596|T102|relax|68596-6|LNC|Plastic surgery Transfer|Plastic surgery Transfer
C1316596|T102|relax|68482-9|LNC|Nurse Hospital Transfer|Nurse Hospital Transfer
C1316596|T102|relax|68884-6|LNC|Pediatrics Hospital Transfer|Pediatrics Hospital Transfer
C1547673|T102|strict|11369-6|LNC|History of Immunization|History of Immunization
C1547673|T102|strict|11485-0|LNC|Anesthesia records|Anesthesia records
C1547673|T102|strict|11486-8|LNC|Chemotherapy records|Chemotherapy records
C1547673|T102|strict|11488-4|LNC|Consult Note|Consult Note
C1547673|T102|strict|11506-3|LNC|Provider-unspecified progress note|Provider-unspecified progress note
C1547673|T102|strict|11543-6|LNC|Nursery records|Nursery records
C1547673|T102|strict|15508-5|LNC|Labor and delivery records|Labor and delivery records
C1547673|T102|strict|18726-0|LNC|Radiology studies (set)|Radiology studies (set)
C1547673|T102|strict|18761-7|LNC|Provider-unspecified transfer summary|Provider-unspecified transfer summary
C1547673|T102|strict|18842-5|LNC|Discharge summary|Discharge summary
C1547673|T102|strict|26436-6|LNC|Laboratory Studies (set)|Laboratory Studies (set)
C1547673|T102|strict|26441-6|LNC|Cardiology studies (set)|Cardiology studies (set)
C1547673|T102|strict|26442-4|LNC|Obstetrical studies (set)|Obstetrical studies (set)
C1547673|T102|strict|27895-2|LNC|Gastroenterology endoscopy studies (set)|Gastroenterology endoscopy studies (set)
C1547673|T102|strict|27896-0|LNC|Pulmonary studies (set)|Pulmonary studies (set)
C1547673|T102|strict|27897-8|LNC|Neuromuscular electrophysiology studies (set)|Neuromuscular electrophysiology studies (set)
C1547673|T102|strict|27898-6|LNC|Pathology studies (set)|Pathology studies (set)
C1547673|T102|strict|28570-0|LNC|Provider-unspecified procedure note|Provider-unspecified procedure note
C1547673|T102|strict|28619-5|LNC|Ophthalmology/optometry studies (set)|Ophthalmology/optometry studies (set)
C1547673|T102|strict|28634-4|LNC|Miscellaneous studies (set)|Miscellaneous studies (set)
C1547673|T102|strict|29749-9|LNC|Dialysis records|Dialysis records
C1547673|T102|strict|29750-7|LNC|Neonatal intensive care records|Neonatal intensive care records
C1547673|T102|strict|29751-5|LNC|Critical care records|Critical care records
C1547673|T102|strict|29752-3|LNC|Perioperative records|Perioperative records
C1547673|T102|strict|34109-9|LNC|Evaluation and management note|Evaluation and management note
C1547673|T102|strict|34117-2|LNC|Provider-unspecified, History and physical note|Provider-unspecified, History and physical note
C1547673|T102|strict|34121-4|LNC|Interventional procedure note|Interventional procedure note
C1547673|T102|strict|34122-2|LNC|Pathology procedure note|Pathology procedure note
C1547673|T102|strict|34133-9|LNC|Summarization of episode note|Summarization of episode note
C1547673|T102|strict|34140-4|LNC|Transfer of care referral note|Transfer of care referral note
C1547673|T102|strict|34748-4|LNC|Telephone encounter note|Telephone encounter note
C1547673|T102|strict|34775-7|LNC|General surgery Pre-operative evaluation and management note|General surgery Pre-operative evaluation and management note
C1547673|T102|strict|47039-3|LNC|Inpatient Admission history and physical note|Inpatient Admission history and physical note
C1547673|T102|strict|47042-7|LNC|Counseling note|Counseling note
C1547673|T102|strict|47045-0|LNC|Study report Document|Study report Document
C1547673|T102|strict|47046-8|LNC|Summary of death|Summary of death
C1547673|T102|strict|47049-2|LNC|Non-patient Communication|Non-patient Communication
C1547673|T102|strict|57017-6|LNC|Privacy Policy Organization Document|Privacy Policy Organization Document
C1547673|T102|strict|57016-8|LNC|Privacy Policy Acknowledgment Document|Privacy Policy Acknowledgment Document
C1547673|T102|strict|56445-0|LNC|Medication Summary Document|Medication Summary Document
C1547673|T102|strict|53576-5|LNC|Personal health monitoring report Document|Personal health monitoring report Document
C1547673|T102|strict|56447-6|LNC|Plan of care note|Plan of care note
C1547673|T102|strict|18748-4|LNC|Diagnostic imaging study|Diagnostic imaging study
C1547673|T102|strict|11504-8|LNC|Surgical operation note|Surgical operation note
C1547673|T102|strict|57133-1|LNC|Referral note|Referral note
C1547673|T102|relax|11488-4|LNC|Consult|Consult
C1547673|T102|relax|11506-3|LNC|Provider progress note|Provider progress note
C1547673|T102|relax|18726-0|LNC|Radiology studies|Radiology studies
C1547673|T102|relax|18761-7|LNC|Provider transfer summary|Provider transfer summary
C1547673|T102|relax|26436-6|LNC|Laboratory Studies|Laboratory Studies
C1547673|T102|relax|26441-6|LNC|Cardiology studies|Cardiology studies
C1547673|T102|relax|26442-4|LNC|Obstetrical studies|Obstetrical studies
C1547673|T102|relax|27895-2|LNC|Gastroenterology endoscopy studies|Gastroenterology endoscopy studies
C1547673|T102|relax|27896-0|LNC|Pulmonary studies|Pulmonary studies
C1547673|T102|relax|27897-8|LNC|Neuromuscular electrophysiology studies|Neuromuscular electrophysiology studies
C1547673|T102|relax|27898-6|LNC|Pathology studies|Pathology studies
C1547673|T102|relax|28570-0|LNC|Provider procedure note|Provider procedure note
C1547673|T102|relax|28619-5|LNC|Ophthalmology/optometry studies|Ophthalmology/optometry studies
C1547673|T102|relax|28634-4|LNC|Miscellaneous studies|Miscellaneous studies
C1547673|T102|relax|34109-9|LNC|Evaluation and management|Evaluation and management
C1547673|T102|relax|34117-2|LNC|Provider History and physical|Provider History and physical
C1547673|T102|relax|34121-4|LNC|Interventional procedure|Interventional procedure
C1547673|T102|relax|34122-2|LNC|Pathology procedure|Pathology procedure
C1547673|T102|relax|34133-9|LNC|Summarization of episode|Summarization of episode
C1547673|T102|relax|34140-4|LNC|Transfer of care referral|Transfer of care referral
C1547673|T102|relax|34748-4|LNC|Telephone encounter|Telephone encounter
C1547673|T102|relax|34775-7|LNC|Pre-operative evaluation and management|Pre-operative evaluation and management
C1547673|T102|relax|47039-3|LNC|Inpatient Admission history and physical|Inpatient Admission history and physical
C1547673|T102|relax|47045-0|LNC|Study report|Study report
C1547673|T102|relax|57017-6|LNC|Privacy Policy Document|Privacy Policy Document
C1547673|T102|relax|57016-8|LNC|Privacy Policy Acknowledgment|Privacy Policy Acknowledgment
C1547673|T102|relax|56445-0|LNC|Medication Summary|Medication Summary
C1547673|T102|relax|53576-5|LNC|Personal health monitoring report|Personal health monitoring report
C1547673|T102|relax|56447-6|LNC|Plan of care|Plan of care
C1547673|T102|relax|18748-4|LNC|Diagnostic imaging report|Diagnostic imaging report
C2826012|T102|strict|55107-7|LNC|Addendum Document|Addendum Document
C2826012|T102|strict|74155-3|LNC|ADHD action plan|ADHD action plan
C2826012|T102|strict|51851-4|LNC|Administrative note|Administrative note
C2826012|T102|strict|67851-6|LNC|Admission evaluation note|Admission evaluation note
C2826012|T102|strict|34744-3|LNC|Nurse Admission evaluation note|Nurse Admission evaluation note
C2826012|T102|strict|34873-0|LNC|Surgery Admission evaluation note|Surgery Admission evaluation note
C2826012|T102|strict|68552-9|LNC|Emergency medicine Emergency department Admission evaluation note|Emergency medicine Emergency department Admission evaluation note
C2826012|T102|strict|67852-4|LNC|Hospital Admission evaluation note|Hospital Admission evaluation note
C2826012|T102|strict|68471-2|LNC|Cardiology Hospital Admission evaluation note|Cardiology Hospital Admission evaluation note
C2826012|T102|strict|68483-7|LNC|Cardiology Medical student Hospital Admission evaluation note|Cardiology Medical student Hospital Admission evaluation note
C2826012|T102|strict|64058-1|LNC|Critical Care Medicine Hospital Admission evaluation note|Critical Care Medicine Hospital Admission evaluation note
C2826012|T102|strict|64070-6|LNC|Critical care medicine Medical student Hospital Admission evaluation note|Critical care medicine Medical student Hospital Admission evaluation note
C2826012|T102|strict|64053-2|LNC|General medicine Hospital Admission evaluation note|General medicine Hospital Admission evaluation note
C2826012|T102|strict|64054-0|LNC|General medicine Medical student Hospital Admission evaluation note|General medicine Medical student Hospital Admission evaluation note
C2826012|T102|strict|34862-3|LNC|General medicine Physician attending Hospital Admission evaluation note|General medicine Physician attending Hospital Admission evaluation note
C2826012|T102|strict|64062-3|LNC|Pulmonary Hospital Admission evaluation note|Pulmonary Hospital Admission evaluation note
C2826012|T102|strict|64078-9|LNC|Pulmonary Medical student Hospital Admission evaluation note|Pulmonary Medical student Hospital Admission evaluation note
C2826012|T102|strict|64066-4|LNC|Surgery Medical student Hospital Admission evaluation note|Surgery Medical student Hospital Admission evaluation note
C2826012|T102|strict|64060-7|LNC|Thoracic surgery Hospital Admission evaluation note|Thoracic surgery Hospital Admission evaluation note
C2826012|T102|strict|64074-8|LNC|Thoracic surgery Medical student Hospital Admission evaluation note|Thoracic surgery Medical student Hospital Admission evaluation note
C2826012|T102|strict|51849-8|LNC|Admission history and physical note|Admission history and physical note
C2826012|T102|strict|34763-3|LNC|General medicine Admission history and physical note|General medicine Admission history and physical note
C2826012|T102|strict|47039-3|LNC|Hospital Admission history and physical note|Hospital Admission history and physical note
C2826012|T102|strict|34094-3|LNC|Cardiology Hospital Admission history and physical note|Cardiology Hospital Admission history and physical note
C2826012|T102|strict|57830-2|LNC|Admission request Document|Admission request Document
C2826012|T102|strict|48765-2|LNC|Allergies and adverse reactions Document|Allergies and adverse reactions Document
C2826012|T102|strict|74152-0|LNC|Anaphylaxis action plan|Anaphylaxis action plan
C2826012|T102|strict|61359-6|LNC|Patient Anesthesia consent|Patient Anesthesia consent
C2826012|T102|strict|57055-6|LNC|Antepartum summary note|Antepartum summary note
C2826012|T102|strict|56446-8|LNC|Appointment summary Document|Appointment summary Document
C2826012|T102|strict|51848-0|LNC|Assessment note|Assessment note
C2826012|T102|strict|68814-3|LNC|Pediatrics Assessment note|Pediatrics Assessment note
C2826012|T102|strict|64064-9|LNC|Pastoral care Hospital Assessment note|Pastoral care Hospital Assessment note
C2826012|T102|strict|51847-2|LNC|Assessment + Plan note|Assessment + Plan note
C2826012|T102|strict|69981-9|LNC|Asthma action plan|Asthma action plan
C2826012|T102|strict|74154-6|LNC|Autism action plan|Autism action plan
C2826012|T102|strict|71230-7|LNC|Birth certificate Document|Birth certificate Document
C2826012|T102|strict|72134-0|LNC|Cancer event report|Cancer event report
C2826012|T102|strict|55108-5|LNC|Clinical presentation Document|Clinical presentation Document
C2826012|T102|strict|73568-8|LNC|Communication of critical results [Description] Document|Communication of critical results [Description] Document
C2826012|T102|strict|74144-7|LNC|Complex medical conditions action plan|Complex medical conditions action plan
C2826012|T102|strict|55109-3|LNC|Complications Document|Complications Document
C2826012|T102|strict|34095-0|LNC|Comprehensive history and physical note|Comprehensive history and physical note
C2826012|T102|strict|34096-8|LNC|Nursing facility Comprehensive history and physical note|Nursing facility Comprehensive history and physical note
C2826012|T102|strict|63485-7|LNC|Computer generated recommendation Document|Computer generated recommendation Document
C2826012|T102|strict|55110-1|LNC|Conclusions Document|Conclusions Document
C2826012|T102|strict|34098-4|LNC|Conference note|Conference note
C2826012|T102|strict|34097-6|LNC|Nursing facility Conference note|Nursing facility Conference note
C2826012|T102|strict|47040-1|LNC|Consultation 2nd opinion|Consultation 2nd opinion
C2826012|T102|strict|47041-9|LNC|Hospital Consultation 2nd opinion|Hospital Consultation 2nd opinion
C2826012|T102|strict|59284-0|LNC|Patient Consent|Patient Consent
C2826012|T102|strict|11488-4|LNC|Consult note|Consult note
C2826012|T102|strict|34099-2|LNC|Cardiology Consult note|Cardiology Consult note
C2826012|T102|strict|34756-7|LNC|Dentistry Consult note|Dentistry Consult note
C2826012|T102|strict|34758-3|LNC|Dermatology Consult note|Dermatology Consult note
C2826012|T102|strict|34760-9|LNC|Diabetology Consult note|Diabetology Consult note
C2826012|T102|strict|34879-7|LNC|Endocrinology Consult note|Endocrinology Consult note
C2826012|T102|strict|34761-7|LNC|Gastroenterology Consult note|Gastroenterology Consult note
C2826012|T102|strict|34764-1|LNC|General medicine Consult note|General medicine Consult note
C2826012|T102|strict|34776-5|LNC|Geriatric medicine Consult note|Geriatric medicine Consult note
C2826012|T102|strict|34779-9|LNC|Hematology+Medical Oncology Consult note|Hematology+Medical Oncology Consult note
C2826012|T102|strict|34781-5|LNC|Infectious disease Consult note|Infectious disease Consult note
C2826012|T102|strict|72555-6|LNC|Interventional radiology Consult note|Interventional radiology Consult note
C2826012|T102|strict|34783-1|LNC|Kinesiotherapy Consult note|Kinesiotherapy Consult note
C2826012|T102|strict|34785-6|LNC|Mental health Consult note|Mental health Consult note
C2826012|T102|strict|34795-5|LNC|Nephrology Consult note|Nephrology Consult note
C2826012|T102|strict|34798-9|LNC|Neurological surgery Consult note|Neurological surgery Consult note
C2826012|T102|strict|34797-1|LNC|Neurology Consult note|Neurology Consult note
C2826012|T102|strict|34800-3|LNC|Nutrition and dietetics Consult note|Nutrition and dietetics Consult note
C2826012|T102|strict|34777-3|LNC|Obstetrics and Gynecology Consult note|Obstetrics and Gynecology Consult note
C2826012|T102|strict|34803-7|LNC|Occupational medicine Consult note|Occupational medicine Consult note
C2826012|T102|strict|34855-7|LNC|Occupational therapy Consult note|Occupational therapy Consult note
C2826012|T102|strict|34805-2|LNC|Oncology Consult note|Oncology Consult note
C2826012|T102|strict|34807-8|LNC|Ophthalmology Consult note|Ophthalmology Consult note
C2826012|T102|strict|34810-2|LNC|Optometry Consult note|Optometry Consult note
C2826012|T102|strict|34812-8|LNC|Oral and Maxillofacial Surgery Consult note|Oral and Maxillofacial Surgery Consult note
C2826012|T102|strict|34814-4|LNC|Orthopaedic surgery Consult note|Orthopaedic surgery Consult note
C2826012|T102|strict|34816-9|LNC|Otolaryngology Consult note|Otolaryngology Consult note
C2826012|T102|strict|34820-1|LNC|Pharmacy Consult note|Pharmacy Consult note
C2826012|T102|strict|34822-7|LNC|Physical medicine and rehabilitation Consult note|Physical medicine and rehabilitation Consult note
C2826012|T102|strict|34824-3|LNC|Physical therapy Consult note|Physical therapy Consult note
C2826012|T102|strict|34826-8|LNC|Plastic surgery Consult note|Plastic surgery Consult note
C2826012|T102|strict|34828-4|LNC|Podiatry Consult note|Podiatry Consult note
C2826012|T102|strict|34788-0|LNC|Psychiatry Consult note|Psychiatry Consult note
C2826012|T102|strict|34791-4|LNC|Psychology Consult note|Psychology Consult note
C2826012|T102|strict|34103-2|LNC|Pulmonary Consult note|Pulmonary Consult note
C2826012|T102|strict|34831-8|LNC|Radiation oncology Consult note|Radiation oncology Consult note
C2826012|T102|strict|73575-3|LNC|Radiology Consult note|Radiology Consult note
C2826012|T102|strict|34833-4|LNC|Recreational therapy Consult note|Recreational therapy Consult note
C2826012|T102|strict|34837-5|LNC|Respiratory therapy Consult note|Respiratory therapy Consult note
C2826012|T102|strict|34839-1|LNC|Rheumatology Consult note|Rheumatology Consult note
C2826012|T102|strict|34841-7|LNC|Social work Consult note|Social work Consult note
C2826012|T102|strict|34845-8|LNC|Speech-language pathology+Audiology Consult note|Speech-language pathology+Audiology Consult note
C2826012|T102|strict|34847-4|LNC|Surgery Consult note|Surgery Consult note
C2826012|T102|strict|34849-0|LNC|Thoracic surgery Consult note|Thoracic surgery Consult note
C2826012|T102|strict|34851-6|LNC|Urology Consult note|Urology Consult note
C2826012|T102|strict|34853-2|LNC|Vascular surgery Consult note|Vascular surgery Consult note
C2826012|T102|strict|51846-4|LNC|Emergency department Consult note|Emergency department Consult note
C2826012|T102|strict|34104-0|LNC|Hospital Consult note|Hospital Consult note
C2826012|T102|strict|68619-6|LNC|Adolescent medicine Hospital Consult note|Adolescent medicine Hospital Consult note
C2826012|T102|strict|68633-7|LNC|Allergy and immunology Hospital Consult note|Allergy and immunology Hospital Consult note
C2826012|T102|strict|68639-4|LNC|Audiology Hospital Consult note|Audiology Hospital Consult note
C2826012|T102|strict|68486-0|LNC|Cardiology Medical student Hospital Consult note|Cardiology Medical student Hospital Consult note
C2826012|T102|strict|68648-5|LNC|Child and adolescent psychiatry Hospital Consult note|Child and adolescent psychiatry Hospital Consult note
C2826012|T102|strict|68651-9|LNC|Clinical biochemical genetics Hospital Consult note|Clinical biochemical genetics Hospital Consult note
C2826012|T102|strict|68661-8|LNC|Clinical genetics Hospital Consult note|Clinical genetics Hospital Consult note
C2826012|T102|strict|64072-2|LNC|Critical care medicine Medical student Hospital Consult note|Critical care medicine Medical student Hospital Consult note
C2826012|T102|strict|68551-1|LNC|Dermatology Hospital Consult note|Dermatology Hospital Consult note
C2826012|T102|strict|68670-9|LNC|Developmental-behavioral pediatrics Hospital Consult note|Developmental-behavioral pediatrics Hospital Consult note
C2826012|T102|strict|64056-5|LNC|General medicine Medical student Hospital Consult note|General medicine Medical student Hospital Consult note
C2826012|T102|strict|68681-6|LNC|Multi-specialty program Hospital Consult note|Multi-specialty program Hospital Consult note
C2826012|T102|strict|68685-7|LNC|Neonatal perinatal medicine Hospital Consult note|Neonatal perinatal medicine Hospital Consult note
C2826012|T102|strict|68694-9|LNC|Neurological surgery Hospital Consult note|Neurological surgery Hospital Consult note
C2826012|T102|strict|68705-3|LNC|Neurology with special qualifications in child neurology Hospital Consult note|Neurology with special qualifications in child neurology Hospital Consult note
C2826012|T102|strict|68566-9|LNC|Obstetrics and Gynecology Hospital Consult note|Obstetrics and Gynecology Hospital Consult note
C2826012|T102|strict|68570-1|LNC|Occupational therapy Hospital Consult note|Occupational therapy Hospital Consult note
C2826012|T102|strict|68575-0|LNC|Ophthalmology Hospital Consult note|Ophthalmology Hospital Consult note
C2826012|T102|strict|68716-0|LNC|Pain medicine Hospital Consult note|Pain medicine Hospital Consult note
C2826012|T102|strict|68469-6|LNC|Pastoral care Hospital Consult note|Pastoral care Hospital Consult note
C2826012|T102|strict|68727-7|LNC|Pediatric cardiology Hospital Consult note|Pediatric cardiology Hospital Consult note
C2826012|T102|strict|68892-9|LNC|Pediatric dermatology Hospital Consult note|Pediatric dermatology Hospital Consult note
C2826012|T102|strict|68897-8|LNC|Pediatric endocrinology Hospital Consult note|Pediatric endocrinology Hospital Consult note
C2826012|T102|strict|68746-7|LNC|Pediatric gastroenterology Hospital Consult note|Pediatric gastroenterology Hospital Consult note
C2826012|T102|strict|68757-4|LNC|Pediatric hematology-oncology Hospital Consult note|Pediatric hematology-oncology Hospital Consult note
C2826012|T102|strict|68765-7|LNC|Pediatric infectious diseases Hospital Consult note|Pediatric infectious diseases Hospital Consult note
C2826012|T102|strict|68869-7|LNC|Pediatric nephrology Hospital Consult note|Pediatric nephrology Hospital Consult note
C2826012|T102|strict|68874-7|LNC|Pediatric otolaryngology Hospital Consult note|Pediatric otolaryngology Hospital Consult note
C2826012|T102|strict|68787-1|LNC|Pediatric pulmonology Hospital Consult note|Pediatric pulmonology Hospital Consult note
C2826012|T102|strict|68879-6|LNC|Pediatric rheumatology Hospital Consult note|Pediatric rheumatology Hospital Consult note
C2826012|T102|strict|68802-8|LNC|Pediatric surgery Hospital Consult note|Pediatric surgery Hospital Consult note
C2826012|T102|strict|68864-8|LNC|Pediatric transplant hepatology Hospital Consult note|Pediatric transplant hepatology Hospital Consult note
C2826012|T102|strict|68812-7|LNC|Pediatric urology Hospital Consult note|Pediatric urology Hospital Consult note
C2826012|T102|strict|68821-8|LNC|Pediatrics Hospital Consult note|Pediatrics Hospital Consult note
C2826012|T102|strict|68586-7|LNC|Pharmacy Hospital Consult note|Pharmacy Hospital Consult note
C2826012|T102|strict|68590-9|LNC|Physical therapy Hospital Consult note|Physical therapy Hospital Consult note
C2826012|T102|strict|68597-4|LNC|Plastic surgery Hospital Consult note|Plastic surgery Hospital Consult note
C2826012|T102|strict|68837-4|LNC|Primary care Hospital Consult note|Primary care Hospital Consult note
C2826012|T102|strict|34102-4|LNC|Psychiatry Hospital Consult note|Psychiatry Hospital Consult note
C2826012|T102|strict|64080-5|LNC|Pulmonary Medical student Hospital Consult note|Pulmonary Medical student Hospital Consult note
C2826012|T102|strict|68846-5|LNC|Speech-language pathology Hospital Consult note|Speech-language pathology Hospital Consult note
C2826012|T102|strict|64068-0|LNC|Surgery Medical student Hospital Consult note|Surgery Medical student Hospital Consult note
C2826012|T102|strict|64076-3|LNC|Thoracic surgery Medical student Hospital Consult note|Thoracic surgery Medical student Hospital Consult note
C2826012|T102|strict|68852-3|LNC|Transplant surgery Hospital Consult note|Transplant surgery Hospital Consult note
C2826012|T102|strict|34100-8|LNC|Intensive care unit Consult note|Intensive care unit Consult note
C2826012|T102|strict|51854-8|LNC|Long term care facility Consult note|Long term care facility Consult note
C2826012|T102|strict|51845-6|LNC|Outpatient Consult note|Outpatient Consult note
C2826012|T102|strict|34749-2|LNC|Anesthesiology Outpatient Consult note|Anesthesiology Outpatient Consult note
C2826012|T102|strict|34101-6|LNC|General medicine Outpatient Consult note|General medicine Outpatient Consult note
C2826012|T102|strict|47042-7|LNC|Counseling note|Counseling note
C2826012|T102|strict|34864-9|LNC|Mental health Counseling note|Mental health Counseling note
C2826012|T102|strict|34869-8|LNC|Pharmacy Counseling note|Pharmacy Counseling note
C2826012|T102|strict|34865-6|LNC|Psychiatry Counseling note|Psychiatry Counseling note
C2826012|T102|strict|34866-4|LNC|Psychology Counseling note|Psychology Counseling note
C2826012|T102|strict|34872-2|LNC|Social work Counseling note|Social work Counseling note
C2826012|T102|strict|55111-9|LNC|Current imaging procedure descriptions Document|Current imaging procedure descriptions Document
C2826012|T102|strict|74148-8|LNC|Cystic fibrosis action plan|Cystic fibrosis action plan
C2826012|T102|strict|64297-5|LNC|Death certificate|Death certificate
C2826012|T102|strict|74208-0|LNC|Demographic information + History of occupation Document|Demographic information + History of occupation Document
C2826012|T102|strict|51899-3|LNC|Details Document|Details Document
C2826012|T102|strict|74150-4|LNC|Diabetes type I action plan|Diabetes type I action plan
C2826012|T102|strict|74151-2|LNC|Diabetes type II action plan|Diabetes type II action plan
C2826012|T102|strict|47048-4|LNC|Diagnostic interventional study report Interventional radiology|Diagnostic interventional study report Interventional radiology
C2826012|T102|strict|70004-7|LNC|Diagnostic study note|Diagnostic study note
C2826012|T102|strict|68611-3|LNC|Adolescent medicine Diagnostic study note|Adolescent medicine Diagnostic study note
C2826012|T102|strict|68625-3|LNC|Allergy and immunology Diagnostic study note|Allergy and immunology Diagnostic study note
C2826012|T102|strict|68635-2|LNC|Audiology Diagnostic study note|Audiology Diagnostic study note
C2826012|T102|strict|68641-0|LNC|Child and adolescent psychiatry Diagnostic study note|Child and adolescent psychiatry Diagnostic study note
C2826012|T102|strict|68652-7|LNC|Clinical genetics Diagnostic study note|Clinical genetics Diagnostic study note
C2826012|T102|strict|68673-3|LNC|Multi-specialty program Diagnostic study note|Multi-specialty program Diagnostic study note
C2826012|T102|strict|68687-3|LNC|Neurological surgery Diagnostic study note|Neurological surgery Diagnostic study note
C2826012|T102|strict|68556-0|LNC|Neurology Diagnostic study note|Neurology Diagnostic study note
C2826012|T102|strict|68696-4|LNC|Neurology with special qualifications in child neurology Diagnostic study note|Neurology with special qualifications in child neurology Diagnostic study note
C2826012|T102|strict|68557-8|LNC|Obstetrics and Gynecology Diagnostic study note|Obstetrics and Gynecology Diagnostic study note
C2826012|T102|strict|68577-6|LNC|Orthopaedic surgery Diagnostic study note|Orthopaedic surgery Diagnostic study note
C2826012|T102|strict|68708-7|LNC|Pain medicine Diagnostic study note|Pain medicine Diagnostic study note
C2826012|T102|strict|68718-6|LNC|Pediatric cardiology Diagnostic study note|Pediatric cardiology Diagnostic study note
C2826012|T102|strict|68748-3|LNC|Pediatric hematology-oncology Diagnostic study note|Pediatric hematology-oncology Diagnostic study note
C2826012|T102|strict|68767-3|LNC|Pediatric nephrology Diagnostic study note|Pediatric nephrology Diagnostic study note
C2826012|T102|strict|68778-0|LNC|Pediatric pulmonology Diagnostic study note|Pediatric pulmonology Diagnostic study note
C2826012|T102|strict|68794-7|LNC|Pediatric surgery Diagnostic study note|Pediatric surgery Diagnostic study note
C2826012|T102|strict|68855-6|LNC|Pediatric transplant hepatology Diagnostic study note|Pediatric transplant hepatology Diagnostic study note
C2826012|T102|strict|68804-4|LNC|Pediatric urology Diagnostic study note|Pediatric urology Diagnostic study note
C2826012|T102|strict|68604-8|LNC|Radiology Diagnostic study note|Radiology Diagnostic study note
C2826012|T102|strict|68640-2|LNC|Audiology Hospital Diagnostic study note|Audiology Hospital Diagnostic study note
C2826012|T102|strict|68706-1|LNC|Neurology with special qualifications in child neurology Hospital Diagnostic study note|Neurology with special qualifications in child neurology Hospital Diagnostic study note
C2826012|T102|strict|68788-9|LNC|Pediatric pulmonology Hospital Diagnostic study note|Pediatric pulmonology Hospital Diagnostic study note
C2826012|T102|strict|68822-6|LNC|Pediatrics Hospital Diagnostic study note|Pediatrics Hospital Diagnostic study note
C2826012|T102|strict|74213-0|LNC|Discharge instructions|Discharge instructions
C2826012|T102|strict|60280-5|LNC|Emergency department Discharge instructions|Emergency department Discharge instructions
C2826012|T102|strict|8653-8|LNC|Hospital Discharge instructions|Hospital Discharge instructions
C2826012|T102|strict|18842-5|LNC|Discharge summary|Discharge summary
C2826012|T102|strict|68612-1|LNC|Adolescent medicine Discharge summary|Adolescent medicine Discharge summary
C2826012|T102|strict|68626-1|LNC|Allergy and immunology Discharge summary|Allergy and immunology Discharge summary
C2826012|T102|strict|68642-8|LNC|Child and adolescent psychiatry Discharge summary|Child and adolescent psychiatry Discharge summary
C2826012|T102|strict|68653-5|LNC|Clinical genetics Discharge summary|Clinical genetics Discharge summary
C2826012|T102|strict|68663-4|LNC|Developmental-behavioral pediatrics Discharge summary|Developmental-behavioral pediatrics Discharge summary
C2826012|T102|strict|68674-1|LNC|Multi-specialty program Discharge summary|Multi-specialty program Discharge summary
C2826012|T102|strict|68688-1|LNC|Neurological surgery Discharge summary|Neurological surgery Discharge summary
C2826012|T102|strict|68697-2|LNC|Neurology with special qualifications in child neurology Discharge summary|Neurology with special qualifications in child neurology Discharge summary
C2826012|T102|strict|34745-0|LNC|Nurse Discharge summary|Nurse Discharge summary
C2826012|T102|strict|68558-6|LNC|Obstetrics and Gynecology Discharge summary|Obstetrics and Gynecology Discharge summary
C2826012|T102|strict|68572-7|LNC|Ophthalmology Discharge summary|Ophthalmology Discharge summary
C2826012|T102|strict|68578-4|LNC|Orthopaedic surgery Discharge summary|Orthopaedic surgery Discharge summary
C2826012|T102|strict|68709-5|LNC|Pain medicine Discharge summary|Pain medicine Discharge summary
C2826012|T102|strict|68719-4|LNC|Pediatric cardiology Discharge summary|Pediatric cardiology Discharge summary
C2826012|T102|strict|68733-5|LNC|Pediatric endocrinology Discharge summary|Pediatric endocrinology Discharge summary
C2826012|T102|strict|68738-4|LNC|Pediatric gastroenterology Discharge summary|Pediatric gastroenterology Discharge summary
C2826012|T102|strict|68749-1|LNC|Pediatric hematology-oncology Discharge summary|Pediatric hematology-oncology Discharge summary
C2826012|T102|strict|68768-1|LNC|Pediatric nephrology Discharge summary|Pediatric nephrology Discharge summary
C2826012|T102|strict|68773-1|LNC|Pediatric otolaryngology Discharge summary|Pediatric otolaryngology Discharge summary
C2826012|T102|strict|68779-8|LNC|Pediatric pulmonology Discharge summary|Pediatric pulmonology Discharge summary
C2826012|T102|strict|68795-4|LNC|Pediatric surgery Discharge summary|Pediatric surgery Discharge summary
C2826012|T102|strict|68856-4|LNC|Pediatric transplant hepatology Discharge summary|Pediatric transplant hepatology Discharge summary
C2826012|T102|strict|68805-1|LNC|Pediatric urology Discharge summary|Pediatric urology Discharge summary
C2826012|T102|strict|68815-0|LNC|Pediatrics Discharge summary|Pediatrics Discharge summary
C2826012|T102|strict|68591-7|LNC|Plastic surgery Discharge summary|Plastic surgery Discharge summary
C2826012|T102|strict|68831-7|LNC|Primary care Discharge summary|Primary care Discharge summary
C2826012|T102|strict|59259-2|LNC|Psychiatry Discharge summary|Psychiatry Discharge summary
C2826012|T102|strict|68841-6|LNC|Speech-language pathology Discharge summary|Speech-language pathology Discharge summary
C2826012|T102|strict|59258-4|LNC|Emergency department Discharge summary|Emergency department Discharge summary
C2826012|T102|strict|34105-7|LNC|Hospital Discharge summary|Hospital Discharge summary
C2826012|T102|strict|68823-4|LNC|Pediatrics Hospital Discharge summary|Pediatrics Hospital Discharge summary
C2826012|T102|strict|34106-5|LNC|Physician Hospital Discharge summary|Physician Hospital Discharge summary
C2826012|T102|strict|55112-7|LNC|Document summary|Document summary
C2826012|T102|strict|34895-3|LNC|Education note|Education note
C2826012|T102|strict|34897-9|LNC|Diabetology Education note|Diabetology Education note
C2826012|T102|strict|67854-0|LNC|Geriatric medicine Education note|Geriatric medicine Education note
C2826012|T102|strict|68477-9|LNC|Nurse Hospital Education note|Nurse Hospital Education note
C2826012|T102|strict|68605-5|LNC|Recreational therapy Hospital Education note|Recreational therapy Hospital Education note
C2826012|T102|strict|67855-7|LNC|Outpatient Education note|Outpatient Education note
C2826012|T102|strict|34902-7|LNC|Geriatric medicine Outpatient Education note|Geriatric medicine Outpatient Education note
C2826012|T102|strict|34107-3|LNC|Patient's home Education note|Patient's home Education note
C2826012|T102|strict|34856-5|LNC|Evaluation and management of anticoagulation note|Evaluation and management of anticoagulation note
C2826012|T102|strict|34859-9|LNC|Evaluation and management of hyperlipidemia|Evaluation and management of hyperlipidemia
C2826012|T102|strict|34860-7|LNC|Evaluation and management of hypertension|Evaluation and management of hypertension
C2826012|T102|strict|70005-4|LNC|Evaluation and management of smoking cessation|Evaluation and management of smoking cessation
C2826012|T102|strict|64142-3|LNC|Hospital Evaluation and management of smoking cessation|Hospital Evaluation and management of smoking cessation
C2826012|T102|strict|34857-3|LNC|Evaluation and management of substance abuse note|Evaluation and management of substance abuse note
C2826012|T102|strict|72267-8|LNC|Evaluation of mental and physical incapacity certificate Document|Evaluation of mental and physical incapacity certificate Document
C2826012|T102|strict|47420-5|LNC|Functional status assessment note|Functional status assessment note
C2826012|T102|strict|47043-5|LNC|Group counseling note|Group counseling note
C2826012|T102|strict|34787-2|LNC|Mental health Group counseling note|Mental health Group counseling note
C2826012|T102|strict|34790-6|LNC|Psychiatry Group counseling note|Psychiatry Group counseling note
C2826012|T102|strict|34793-0|LNC|Psychology Group counseling note|Psychology Group counseling note
C2826012|T102|strict|34843-3|LNC|Social work Group counseling note|Social work Group counseling note
C2826012|T102|strict|34114-9|LNC|Hospital Group counseling note|Hospital Group counseling note
C2826012|T102|strict|64290-0|LNC|Health insurance card|Health insurance card
C2826012|T102|strict|64291-8|LNC|Health insurance-related form|Health insurance-related form
C2826012|T102|strict|57024-2|LNC|Health Quality Measure document|Health Quality Measure document
C2826012|T102|strict|64289-2|LNC|Health record cover sheet|Health record cover sheet
C2826012|T102|strict|51897-7|LNC|Healthcare Associated Infection report Document|Healthcare Associated Infection report Document
C2826012|T102|strict|56444-3|LNC|Healthcare communication Document|Healthcare communication Document
C2826012|T102|strict|74146-2|LNC|Heart disease action plan|Heart disease action plan
C2826012|T102|strict|34117-2|LNC|History and physical note|History and physical note
C2826012|T102|strict|68614-7|LNC|Adolescent medicine History and physical note|Adolescent medicine History and physical note
C2826012|T102|strict|68622-0|LNC|Advanced heart failure and transplant cardiology History and physical note|Advanced heart failure and transplant cardiology History and physical note
C2826012|T102|strict|68628-7|LNC|Allergy and immunology History and physical note|Allergy and immunology History and physical note
C2826012|T102|strict|68637-8|LNC|Audiology History and physical note|Audiology History and physical note
C2826012|T102|strict|68644-4|LNC|Child and adolescent psychiatry History and physical note|Child and adolescent psychiatry History and physical note
C2826012|T102|strict|68655-0|LNC|Clinical genetics History and physical note|Clinical genetics History and physical note
C2826012|T102|strict|68665-9|LNC|Developmental-behavioral pediatrics History and physical note|Developmental-behavioral pediatrics History and physical note
C2826012|T102|strict|68676-6|LNC|Multi-specialty program History and physical note|Multi-specialty program History and physical note
C2826012|T102|strict|68683-2|LNC|Neonatal perinatal medicine History and physical note|Neonatal perinatal medicine History and physical note
C2826012|T102|strict|68690-7|LNC|Neurological surgery History and physical note|Neurological surgery History and physical note
C2826012|T102|strict|68699-8|LNC|Neurology with special qualifications in child neurology History and physical note|Neurology with special qualifications in child neurology History and physical note
C2826012|T102|strict|68560-2|LNC|Obstetrics and Gynecology History and physical note|Obstetrics and Gynecology History and physical note
C2826012|T102|strict|68573-5|LNC|Ophthalmology History and physical note|Ophthalmology History and physical note
C2826012|T102|strict|68580-0|LNC|Orthopaedic surgery History and physical note|Orthopaedic surgery History and physical note
C2826012|T102|strict|68711-1|LNC|Pain medicine History and physical note|Pain medicine History and physical note
C2826012|T102|strict|68721-0|LNC|Pediatric cardiology History and physical note|Pediatric cardiology History and physical note
C2826012|T102|strict|68731-9|LNC|Pediatric dermatology History and physical note|Pediatric dermatology History and physical note
C2826012|T102|strict|68735-0|LNC|Pediatric endocrinology History and physical note|Pediatric endocrinology History and physical note
C2826012|T102|strict|68740-0|LNC|Pediatric gastroenterology History and physical note|Pediatric gastroenterology History and physical note
C2826012|T102|strict|68751-7|LNC|Pediatric hematology-oncology History and physical note|Pediatric hematology-oncology History and physical note
C2826012|T102|strict|68760-8|LNC|Pediatric infectious diseases History and physical note|Pediatric infectious diseases History and physical note
C2826012|T102|strict|68770-7|LNC|Pediatric nephrology History and physical note|Pediatric nephrology History and physical note
C2826012|T102|strict|68775-6|LNC|Pediatric otolaryngology History and physical note|Pediatric otolaryngology History and physical note
C2826012|T102|strict|68781-4|LNC|Pediatric pulmonology History and physical note|Pediatric pulmonology History and physical note
C2826012|T102|strict|68791-3|LNC|Pediatric rheumatology History and physical note|Pediatric rheumatology History and physical note
C2826012|T102|strict|68797-0|LNC|Pediatric surgery History and physical note|Pediatric surgery History and physical note
C2826012|T102|strict|68858-0|LNC|Pediatric transplant hepatology History and physical note|Pediatric transplant hepatology History and physical note
C2826012|T102|strict|68807-7|LNC|Pediatric urology History and physical note|Pediatric urology History and physical note
C2826012|T102|strict|68817-6|LNC|Pediatrics History and physical note|Pediatrics History and physical note
C2826012|T102|strict|28626-0|LNC|Physician History and physical note|Physician History and physical note
C2826012|T102|strict|68592-5|LNC|Plastic surgery History and physical note|Plastic surgery History and physical note
C2826012|T102|strict|68833-3|LNC|Primary care History and physical note|Primary care History and physical note
C2826012|T102|strict|68599-0|LNC|Psychiatry History and physical note|Psychiatry History and physical note
C2826012|T102|strict|68843-2|LNC|Speech-language pathology History and physical note|Speech-language pathology History and physical note
C2826012|T102|strict|34774-0|LNC|Surgery History and physical note|Surgery History and physical note
C2826012|T102|strict|68849-9|LNC|Transplant surgery History and physical note|Transplant surgery History and physical note
C2826012|T102|strict|11492-6|LNC|Provider-unspecifed, History and physical note|Provider-unspecifed, History and physical note
C2826012|T102|strict|34115-6|LNC|Medical student Hospital History and physical note|Medical student Hospital History and physical note
C2826012|T102|strict|68825-9|LNC|Pediatrics Hospital History and physical note|Pediatrics Hospital History and physical note
C2826012|T102|strict|67856-5|LNC|Nursing facility History and physical note|Nursing facility History and physical note
C2826012|T102|strict|34116-4|LNC|Physician Nursing facility History and physical note|Physician Nursing facility History and physical note
C2826012|T102|strict|74264-3|LNC|HIV summary registry report Document|HIV summary registry report Document
C2826012|T102|strict|74149-6|LNC|Inflammatory bowel disease action plan|Inflammatory bowel disease action plan
C2826012|T102|strict|28636-9|LNC|Provider-unspecified Initial assessment|Provider-unspecified Initial assessment
C2826012|T102|strict|28581-7|LNC|Chiropractic medicine Initial assessment note|Chiropractic medicine Initial assessment note
C2826012|T102|strict|68553-7|LNC|Hematology+Medical Oncology Initial assessment note|Hematology+Medical Oncology Initial assessment note
C2826012|T102|strict|18740-1|LNC|Speech-language pathology Initial assessment note|Speech-language pathology Initial assessment note
C2826012|T102|strict|47044-3|LNC|Hospital Initial assessment note|Hospital Initial assessment note
C2826012|T102|strict|64065-6|LNC|Case manager Hospital Initial assessment note|Case manager Hospital Initial assessment note
C2826012|T102|strict|68470-4|LNC|Respiratory therapy Hospital Initial assessment note|Respiratory therapy Hospital Initial assessment note
C2826012|T102|strict|34119-8|LNC|Nursing facility Initial assessment note|Nursing facility Initial assessment note
C2826012|T102|strict|34120-6|LNC|Outpatient Initial assessment note|Outpatient Initial assessment note
C2826012|T102|strict|34118-0|LNC|Patient's home Initial assessment note|Patient's home Initial assessment note
C2826012|T102|strict|74209-8|LNC|Injury event summary Document|Injury event summary Document
C2826012|T102|strict|74188-4|LNC|InterRAI Acute Care (AC) Hospital Document|InterRAI Acute Care (AC) Hospital Document
C2826012|T102|strict|74194-2|LNC|InterRAI Community Health Assessment (CHA) Document|InterRAI Community Health Assessment (CHA) Document
C2826012|T102|strict|74191-8|LNC|InterRAI Community Health Assessment - Assisted Living Supplement (CHA-AL) Document|InterRAI Community Health Assessment - Assisted Living Supplement (CHA-AL) Document
C2826012|T102|strict|74190-0|LNC|InterRAI Community Health Assessment - Deafblind Supplement (CHA-Db) Document|InterRAI Community Health Assessment - Deafblind Supplement (CHA-Db) Document
C2826012|T102|strict|74193-4|LNC|InterRAI Community Health Assessment - Functional Supplement (CHA-FS) Document|InterRAI Community Health Assessment - Functional Supplement (CHA-FS) Document
C2826012|T102|strict|74192-6|LNC|InterRAI Community Health Assessment - Mental Health Supplement (CHA-MH) Document|InterRAI Community Health Assessment - Mental Health Supplement (CHA-MH) Document
C2826012|T102|strict|74197-5|LNC|InterRAI Contact Assessment (CA) Document|InterRAI Contact Assessment (CA) Document
C2826012|T102|strict|74187-6|LNC|InterRAI Emergency Screener for Psychiatry (ESP) Document|InterRAI Emergency Screener for Psychiatry (ESP) Document
C2826012|T102|strict|74196-7|LNC|InterRAI Home Care (HC) Document|InterRAI Home Care (HC) Document
C2826012|T102|strict|74195-9|LNC|InterRAI Long Term Care Facility (LTCF) Document|InterRAI Long Term Care Facility (LTCF) Document
C2826012|T102|strict|74189-2|LNC|InterRAI Palliative Care (PC) Document|InterRAI Palliative Care (PC) Document
C2826012|T102|strict|34121-4|LNC|Interventional procedure note|Interventional procedure note
C2826012|T102|strict|34896-1|LNC|Cardiology Interventional procedure note|Cardiology Interventional procedure note
C2826012|T102|strict|34899-5|LNC|Gastroenterology Interventional procedure note|Gastroenterology Interventional procedure note
C2826012|T102|strict|55113-5|LNC|Key images Document Radiology|Key images Document Radiology
C2826012|T102|strict|57056-4|LNC|Labor and delivery admission history and physical note|Labor and delivery admission history and physical note
C2826012|T102|strict|57057-2|LNC|Labor and delivery summary note|Labor and delivery summary note
C2826012|T102|strict|64299-1|LNC|Legal document|Legal document
C2826012|T102|strict|51852-2|LNC|Letter|Letter
C2826012|T102|strict|68684-0|LNC|Neonatal perinatal medicine Letter|Neonatal perinatal medicine Letter
C2826012|T102|strict|68866-3|LNC|Pediatric nephrology Letter|Pediatric nephrology Letter
C2826012|T102|strict|68593-3|LNC|Plastic surgery Letter|Plastic surgery Letter
C2826012|T102|strict|68609-7|LNC|Hospital Letter|Hospital Letter
C2826012|T102|strict|68620-4|LNC|Adolescent medicine Hospital Letter|Adolescent medicine Hospital Letter
C2826012|T102|strict|68624-6|LNC|Advanced heart failure and transplant cardiology Hospital Letter|Advanced heart failure and transplant cardiology Hospital Letter
C2826012|T102|strict|68634-5|LNC|Allergy and immunology Hospital Letter|Allergy and immunology Hospital Letter
C2826012|T102|strict|68649-3|LNC|Child and adolescent psychiatry Hospital Letter|Child and adolescent psychiatry Hospital Letter
C2826012|T102|strict|68662-6|LNC|Clinical genetics Hospital Letter|Clinical genetics Hospital Letter
C2826012|T102|strict|68671-7|LNC|Developmental-behavioral pediatrics Hospital Letter|Developmental-behavioral pediatrics Hospital Letter
C2826012|T102|strict|68555-2|LNC|Hematology+Medical Oncology Hospital Letter|Hematology+Medical Oncology Hospital Letter
C2826012|T102|strict|68682-4|LNC|Multi-specialty program Hospital Letter|Multi-specialty program Hospital Letter
C2826012|T102|strict|68686-5|LNC|Neonatal perinatal medicine Hospital Letter|Neonatal perinatal medicine Hospital Letter
C2826012|T102|strict|68695-6|LNC|Neurological surgery Hospital Letter|Neurological surgery Hospital Letter
C2826012|T102|strict|68707-9|LNC|Neurology with special qualifications in child neurology Hospital Letter|Neurology with special qualifications in child neurology Hospital Letter
C2826012|T102|strict|68567-7|LNC|Obstetrics and Gynecology Hospital Letter|Obstetrics and Gynecology Hospital Letter
C2826012|T102|strict|68571-9|LNC|Occupational therapy Hospital Letter|Occupational therapy Hospital Letter
C2826012|T102|strict|68576-8|LNC|Ophthalmology Hospital Letter|Ophthalmology Hospital Letter
C2826012|T102|strict|68585-9|LNC|Orthopaedic surgery Hospital Letter|Orthopaedic surgery Hospital Letter
C2826012|T102|strict|68717-8|LNC|Pain medicine Hospital Letter|Pain medicine Hospital Letter
C2826012|T102|strict|68728-5|LNC|Pediatric cardiology Hospital Letter|Pediatric cardiology Hospital Letter
C2826012|T102|strict|68893-7|LNC|Pediatric dermatology Hospital Letter|Pediatric dermatology Hospital Letter
C2826012|T102|strict|68898-6|LNC|Pediatric endocrinology Hospital Letter|Pediatric endocrinology Hospital Letter
C2826012|T102|strict|68747-5|LNC|Pediatric gastroenterology Hospital Letter|Pediatric gastroenterology Hospital Letter
C2826012|T102|strict|68758-2|LNC|Pediatric hematology-oncology Hospital Letter|Pediatric hematology-oncology Hospital Letter
C2826012|T102|strict|68766-5|LNC|Pediatric infectious diseases Hospital Letter|Pediatric infectious diseases Hospital Letter
C2826012|T102|strict|68870-5|LNC|Pediatric nephrology Hospital Letter|Pediatric nephrology Hospital Letter
C2826012|T102|strict|68875-4|LNC|Pediatric otolaryngology Hospital Letter|Pediatric otolaryngology Hospital Letter
C2826012|T102|strict|68789-7|LNC|Pediatric pulmonology Hospital Letter|Pediatric pulmonology Hospital Letter
C2826012|T102|strict|68880-4|LNC|Pediatric rheumatology Hospital Letter|Pediatric rheumatology Hospital Letter
C2826012|T102|strict|68803-6|LNC|Pediatric surgery Hospital Letter|Pediatric surgery Hospital Letter
C2826012|T102|strict|68865-5|LNC|Pediatric transplant hepatology Hospital Letter|Pediatric transplant hepatology Hospital Letter
C2826012|T102|strict|68813-5|LNC|Pediatric urology Hospital Letter|Pediatric urology Hospital Letter
C2826012|T102|strict|68826-7|LNC|Pediatrics Hospital Letter|Pediatrics Hospital Letter
C2826012|T102|strict|68598-2|LNC|Plastic surgery Hospital Letter|Plastic surgery Hospital Letter
C2826012|T102|strict|68838-2|LNC|Primary care Hospital Letter|Primary care Hospital Letter
C2826012|T102|strict|68847-3|LNC|Speech-language pathology Hospital Letter|Speech-language pathology Hospital Letter
C2826012|T102|strict|68853-1|LNC|Transplant surgery Hospital Letter|Transplant surgery Hospital Letter
C2826012|T102|strict|57058-0|LNC|Maternal discharge summary note|Maternal discharge summary note
C2826012|T102|strict|64285-0|LNC|Medical history screening form|Medical history screening form
C2826012|T102|strict|60590-7|LNC|Medication dispensed.brief Document|Medication dispensed.brief Document
C2826012|T102|strict|60593-1|LNC|Medication dispensed.extended Document|Medication dispensed.extended Document
C2826012|T102|strict|70006-2|LNC|Medication management note|Medication management note
C2826012|T102|strict|68587-5|LNC|Pharmacy Hospital Medication management note|Pharmacy Hospital Medication management note
C2826012|T102|strict|61357-0|LNC|Medication pharmaceutical advice.brief Document|Medication pharmaceutical advice.brief Document
C2826012|T102|strict|61356-2|LNC|Medication pharmaceutical advice.extended Document|Medication pharmaceutical advice.extended Document
C2826012|T102|strict|56445-0|LNC|Medication summary Document|Medication summary Document
C2826012|T102|strict|74145-4|LNC|Multiple sclerosis action plan|Multiple sclerosis action plan
C2826012|T102|strict|74147-0|LNC|Muscular dystrophy action plan|Muscular dystrophy action plan
C2826012|T102|strict|59268-3|LNC|Neonatal care report|Neonatal care report
C2826012|T102|strict|34109-9|LNC|Note|Note
C2826012|T102|strict|68615-4|LNC|Adolescent medicine Note|Adolescent medicine Note
C2826012|T102|strict|68621-2|LNC|Advanced heart failure and transplant cardiology Note|Advanced heart failure and transplant cardiology Note
C2826012|T102|strict|68629-5|LNC|Allergy and immunology Note|Allergy and immunology Note
C2826012|T102|strict|34750-0|LNC|Anesthesiology Note|Anesthesiology Note
C2826012|T102|strict|68636-0|LNC|Audiology Note|Audiology Note
C2826012|T102|strict|34752-6|LNC|Cardiology Note|Cardiology Note
C2826012|T102|strict|68645-1|LNC|Child and adolescent psychiatry Note|Child and adolescent psychiatry Note
C2826012|T102|strict|68650-1|LNC|Clinical biochemical genetics Note|Clinical biochemical genetics Note
C2826012|T102|strict|68656-8|LNC|Clinical genetics Note|Clinical genetics Note
C2826012|T102|strict|34754-2|LNC|Critical Care Medicine Note|Critical Care Medicine Note
C2826012|T102|strict|28618-7|LNC|Dentistry Note|Dentistry Note
C2826012|T102|strict|34759-1|LNC|Dermatology Note|Dermatology Note
C2826012|T102|strict|68666-7|LNC|Developmental-behavioral pediatrics Note|Developmental-behavioral pediatrics Note
C2826012|T102|strict|34861-5|LNC|Diabetology Note|Diabetology Note
C2826012|T102|strict|34878-9|LNC|Emergency medicine Note|Emergency medicine Note
C2826012|T102|strict|34898-7|LNC|Endocrinology Note|Endocrinology Note
C2826012|T102|strict|34762-5|LNC|Gastroenterology Note|Gastroenterology Note
C2826012|T102|strict|34765-8|LNC|General medicine Note|General medicine Note
C2826012|T102|strict|34767-4|LNC|General medicine Medical student Note|General medicine Medical student Note
C2826012|T102|strict|34768-2|LNC|General medicine Nurse Note|General medicine Nurse Note
C2826012|T102|strict|34769-0|LNC|General medicine Physician attending Note|General medicine Physician attending Note
C2826012|T102|strict|34780-7|LNC|Hematology+Medical Oncology Note|Hematology+Medical Oncology Note
C2826012|T102|strict|34782-3|LNC|Infectious disease Note|Infectious disease Note
C2826012|T102|strict|34794-8|LNC|Interdisciplinary Note|Interdisciplinary Note
C2826012|T102|strict|34784-9|LNC|Kinesiotherapy Note|Kinesiotherapy Note
C2826012|T102|strict|34786-4|LNC|Mental health Note|Mental health Note
C2826012|T102|strict|68677-4|LNC|Multi-specialty program Note|Multi-specialty program Note
C2826012|T102|strict|34796-3|LNC|Nephrology Note|Nephrology Note
C2826012|T102|strict|34799-7|LNC|Neurological surgery Note|Neurological surgery Note
C2826012|T102|strict|34905-0|LNC|Neurology Note|Neurology Note
C2826012|T102|strict|68700-4|LNC|Neurology with special qualifications in child neurology Note|Neurology with special qualifications in child neurology Note
C2826012|T102|strict|34746-8|LNC|Nurse Note|Nurse Note
C2826012|T102|strict|34801-1|LNC|Nutrition and dietetics Note|Nutrition and dietetics Note
C2826012|T102|strict|34778-1|LNC|Obstetrics and Gynecology Note|Obstetrics and Gynecology Note
C2826012|T102|strict|34802-9|LNC|Occupational medicine Note|Occupational medicine Note
C2826012|T102|strict|28578-3|LNC|Occupational therapy Note|Occupational therapy Note
C2826012|T102|strict|34806-0|LNC|Oncology Note|Oncology Note
C2826012|T102|strict|34808-6|LNC|Ophthalmology Note|Ophthalmology Note
C2826012|T102|strict|34811-0|LNC|Optometry Note|Optometry Note
C2826012|T102|strict|34813-6|LNC|Oral and Maxillofacial Surgery Note|Oral and Maxillofacial Surgery Note
C2826012|T102|strict|34815-1|LNC|Orthopaedic surgery Note|Orthopaedic surgery Note
C2826012|T102|strict|34817-7|LNC|Otolaryngology Note|Otolaryngology Note
C2826012|T102|strict|34858-1|LNC|Pain medicine Note|Pain medicine Note
C2826012|T102|strict|34906-8|LNC|Pastoral care Note|Pastoral care Note
C2826012|T102|strict|51855-5|LNC|Patient Note|Patient Note
C2826012|T102|strict|68722-8|LNC|Pediatric cardiology Note|Pediatric cardiology Note
C2826012|T102|strict|68889-5|LNC|Pediatric dermatology Note|Pediatric dermatology Note
C2826012|T102|strict|68894-5|LNC|Pediatric endocrinology Note|Pediatric endocrinology Note
C2826012|T102|strict|68741-8|LNC|Pediatric gastroenterology Note|Pediatric gastroenterology Note
C2826012|T102|strict|68752-5|LNC|Pediatric hematology-oncology Note|Pediatric hematology-oncology Note
C2826012|T102|strict|68761-6|LNC|Pediatric infectious diseases Note|Pediatric infectious diseases Note
C2826012|T102|strict|68867-1|LNC|Pediatric nephrology Note|Pediatric nephrology Note
C2826012|T102|strict|68871-3|LNC|Pediatric otolaryngology Note|Pediatric otolaryngology Note
C2826012|T102|strict|68782-2|LNC|Pediatric pulmonology Note|Pediatric pulmonology Note
C2826012|T102|strict|68854-9|LNC|Pediatric rehabilitation medicine Note|Pediatric rehabilitation medicine Note
C2826012|T102|strict|68876-2|LNC|Pediatric rheumatology Note|Pediatric rheumatology Note
C2826012|T102|strict|68881-2|LNC|Pediatric surgery Note|Pediatric surgery Note
C2826012|T102|strict|68859-8|LNC|Pediatric transplant hepatology Note|Pediatric transplant hepatology Note
C2826012|T102|strict|68882-0|LNC|Pediatric urology Note|Pediatric urology Note
C2826012|T102|strict|68818-4|LNC|Pediatrics Note|Pediatrics Note
C2826012|T102|strict|34821-9|LNC|Pharmacy Note|Pharmacy Note
C2826012|T102|strict|34823-5|LNC|Physical medicine and rehabilitation Note|Physical medicine and rehabilitation Note
C2826012|T102|strict|28579-1|LNC|Physical therapy Note|Physical therapy Note
C2826012|T102|strict|34827-6|LNC|Plastic surgery Note|Plastic surgery Note
C2826012|T102|strict|34829-2|LNC|Podiatry Note|Podiatry Note
C2826012|T102|strict|68834-1|LNC|Primary care Note|Primary care Note
C2826012|T102|strict|28628-6|LNC|Psychiatry Note|Psychiatry Note
C2826012|T102|strict|34792-2|LNC|Psychology Note|Psychology Note
C2826012|T102|strict|34830-0|LNC|Pulmonary Note|Pulmonary Note
C2826012|T102|strict|34832-6|LNC|Radiation oncology Note|Radiation oncology Note
C2826012|T102|strict|34834-2|LNC|Recreational therapy Note|Recreational therapy Note
C2826012|T102|strict|68839-0|LNC|Research Note|Research Note
C2826012|T102|strict|34838-3|LNC|Respiratory therapy Note|Respiratory therapy Note
C2826012|T102|strict|34840-9|LNC|Rheumatology Note|Rheumatology Note
C2826012|T102|strict|28653-4|LNC|Social work Note|Social work Note
C2826012|T102|strict|28571-8|LNC|Speech-language pathology Note|Speech-language pathology Note
C2826012|T102|strict|34846-6|LNC|Speech-language pathology+Audiology Note|Speech-language pathology+Audiology Note
C2826012|T102|strict|34848-2|LNC|Surgery Note|Surgery Note
C2826012|T102|strict|34773-2|LNC|Surgery Physician attending Note|Surgery Physician attending Note
C2826012|T102|strict|68848-1|LNC|Transplant surgery Note|Transplant surgery Note
C2826012|T102|strict|34852-4|LNC|Urology Note|Urology Note
C2826012|T102|strict|34111-5|LNC|Emergency department Note|Emergency department Note
C2826012|T102|strict|57053-1|LNC|Nurse Emergency department Note|Nurse Emergency department Note
C2826012|T102|strict|34112-3|LNC|Hospital Note|Hospital Note
C2826012|T102|strict|64069-8|LNC|Critical care medicine Physician attending Hospital Note|Critical care medicine Physician attending Hospital Note
C2826012|T102|strict|68827-5|LNC|Pediatrics Hospital Note|Pediatrics Hospital Note
C2826012|T102|strict|64077-1|LNC|Pulmonary Physician attending Hospital Note|Pulmonary Physician attending Hospital Note
C2826012|T102|strict|64073-0|LNC|Thoracic surgery Physician attending Hospital Note|Thoracic surgery Physician attending Hospital Note
C2826012|T102|strict|34113-1|LNC|Nursing facility Note|Nursing facility Note
C2826012|T102|strict|34108-1|LNC|Outpatient Note|Outpatient Note
C2826012|T102|strict|34753-4|LNC|Cardiology Outpatient Note|Cardiology Outpatient Note
C2826012|T102|strict|34110-7|LNC|Diabetology Outpatient Note|Diabetology Outpatient Note
C2826012|T102|strict|34766-6|LNC|General medicine Outpatient Note|General medicine Outpatient Note
C2826012|T102|strict|68601-4|LNC|Psychiatry Outpatient Note|Psychiatry Outpatient Note
C2826012|T102|strict|34850-8|LNC|Thoracic surgery Outpatient Note|Thoracic surgery Outpatient Note
C2826012|T102|strict|34854-0|LNC|Vascular surgery Outpatient Note|Vascular surgery Outpatient Note
C2826012|T102|strict|68672-5|LNC|Geriatric medicine Skilled nursing facility Note|Geriatric medicine Skilled nursing facility Note
C2826012|T102|strict|34748-4|LNC|Telephone encounter Note|Telephone encounter Note
C2826012|T102|strict|34139-6|LNC|Nurse Telephone encounter Note|Nurse Telephone encounter Note
C2826012|T102|strict|34844-1|LNC|Social work Telephone encounter Note|Social work Telephone encounter Note
C2826012|T102|strict|74166-0|LNC|Occupational summary note|Occupational summary note
C2826012|T102|strict|74156-1|LNC|Oncology treatment plan and summary Document|Oncology treatment plan and summary Document
C2826012|T102|strict|64300-7|LNC|Organ donation consent|Organ donation consent
C2826012|T102|strict|60591-5|LNC|Patient summary Document|Patient summary Document
C2826012|T102|strict|60592-3|LNC|Patient summary.unexpected contact Document|Patient summary.unexpected contact Document
C2826012|T102|strict|57834-4|LNC|Patient transportation request Document|Patient transportation request Document
C2826012|T102|strict|48768-6|LNC|Payment sources Document|Payment sources Document
C2826012|T102|strict|53576-5|LNC|Personal health monitoring report Document|Personal health monitoring report Document
C2826012|T102|strict|64296-7|LNC|Personal health monitoring report Automated|Personal health monitoring report Automated
C2826012|T102|strict|72170-4|LNC|Photographic image Unspecified body region Document|Photographic image Unspecified body region Document
C2826012|T102|strict|56447-6|LNC|Plan of care note|Plan of care note
C2826012|T102|strict|64295-9|LNC|Nurse Plan of care note|Nurse Plan of care note
C2826012|T102|strict|51900-9|LNC|Population Summary note|Population Summary note
C2826012|T102|strict|67860-7|LNC|Postoperative evaluation and management note|Postoperative evaluation and management note
C2826012|T102|strict|67861-5|LNC|Ophthalmology Postoperative evaluation and management note|Ophthalmology Postoperative evaluation and management note
C2826012|T102|strict|34875-5|LNC|Surgery Postoperative evaluation and management note|Surgery Postoperative evaluation and management note
C2826012|T102|strict|34880-5|LNC|Surgery Nurse Postoperative evaluation and management note|Surgery Nurse Postoperative evaluation and management note
C2826012|T102|strict|68610-5|LNC|Hospital Postoperative evaluation and management note|Hospital Postoperative evaluation and management note
C2826012|T102|strict|68606-3|LNC|Surgery Hospital Postoperative evaluation and management note|Surgery Hospital Postoperative evaluation and management note
C2826012|T102|strict|34867-2|LNC|Ophthalmology Outpatient Postoperative evaluation and management note|Ophthalmology Outpatient Postoperative evaluation and management note
C2826012|T102|strict|64298-3|LNC|Power of attorney|Power of attorney
C2826012|T102|strict|74207-2|LNC|Prehospital summary Document|Prehospital summary Document
C2826012|T102|strict|67862-3|LNC|Preoperative evaluation and management note|Preoperative evaluation and management note
C2826012|T102|strict|68616-2|LNC|Adolescent medicine Preoperative evaluation and management note|Adolescent medicine Preoperative evaluation and management note
C2826012|T102|strict|68623-8|LNC|Advanced heart failure and transplant cardiology Preoperative evaluation and management note|Advanced heart failure and transplant cardiology Preoperative evaluation and management note
C2826012|T102|strict|34751-8|LNC|Anesthesiology Preoperative evaluation and management note|Anesthesiology Preoperative evaluation and management note
C2826012|T102|strict|68638-6|LNC|Audiology Preoperative evaluation and management note|Audiology Preoperative evaluation and management note
C2826012|T102|strict|68657-6|LNC|Clinical genetics Preoperative evaluation and management note|Clinical genetics Preoperative evaluation and management note
C2826012|T102|strict|68550-3|LNC|Dermatology Preoperative evaluation and management note|Dermatology Preoperative evaluation and management note
C2826012|T102|strict|68678-2|LNC|Multi-specialty program Preoperative evaluation and management note|Multi-specialty program Preoperative evaluation and management note
C2826012|T102|strict|68691-5|LNC|Neurological surgery Preoperative evaluation and management note|Neurological surgery Preoperative evaluation and management note
C2826012|T102|strict|68701-2|LNC|Neurology with special qualifications in child neurology Preoperative evaluation and management note|Neurology with special qualifications in child neurology Preoperative evaluation and management note
C2826012|T102|strict|34747-6|LNC|Nurse Preoperative evaluation and management note|Nurse Preoperative evaluation and management note
C2826012|T102|strict|68562-8|LNC|Obstetrics and Gynecology Preoperative evaluation and management note|Obstetrics and Gynecology Preoperative evaluation and management note
C2826012|T102|strict|34809-4|LNC|Ophthalmology Preoperative evaluation and management note|Ophthalmology Preoperative evaluation and management note
C2826012|T102|strict|68581-8|LNC|Orthopaedic surgery Preoperative evaluation and management note|Orthopaedic surgery Preoperative evaluation and management note
C2826012|T102|strict|68713-7|LNC|Pain medicine Preoperative evaluation and management note|Pain medicine Preoperative evaluation and management note
C2826012|T102|strict|68723-6|LNC|Pediatric cardiology Preoperative evaluation and management note|Pediatric cardiology Preoperative evaluation and management note
C2826012|T102|strict|68732-7|LNC|Pediatric dermatology Preoperative evaluation and management note|Pediatric dermatology Preoperative evaluation and management note
C2826012|T102|strict|68736-8|LNC|Pediatric endocrinology Preoperative evaluation and management note|Pediatric endocrinology Preoperative evaluation and management note
C2826012|T102|strict|68742-6|LNC|Pediatric gastroenterology Preoperative evaluation and management note|Pediatric gastroenterology Preoperative evaluation and management note
C2826012|T102|strict|68753-3|LNC|Pediatric hematology-oncology Preoperative evaluation and management note|Pediatric hematology-oncology Preoperative evaluation and management note
C2826012|T102|strict|68762-4|LNC|Pediatric infectious diseases Preoperative evaluation and management note|Pediatric infectious diseases Preoperative evaluation and management note
C2826012|T102|strict|68771-5|LNC|Pediatric nephrology Preoperative evaluation and management note|Pediatric nephrology Preoperative evaluation and management note
C2826012|T102|strict|68776-4|LNC|Pediatric otolaryngology Preoperative evaluation and management note|Pediatric otolaryngology Preoperative evaluation and management note
C2826012|T102|strict|68783-0|LNC|Pediatric pulmonology Preoperative evaluation and management note|Pediatric pulmonology Preoperative evaluation and management note
C2826012|T102|strict|68792-1|LNC|Pediatric rheumatology Preoperative evaluation and management note|Pediatric rheumatology Preoperative evaluation and management note
C2826012|T102|strict|68798-8|LNC|Pediatric surgery Preoperative evaluation and management note|Pediatric surgery Preoperative evaluation and management note
C2826012|T102|strict|68860-6|LNC|Pediatric transplant hepatology Preoperative evaluation and management note|Pediatric transplant hepatology Preoperative evaluation and management note
C2826012|T102|strict|68808-5|LNC|Pediatric urology Preoperative evaluation and management note|Pediatric urology Preoperative evaluation and management note
C2826012|T102|strict|68819-2|LNC|Pediatrics Preoperative evaluation and management note|Pediatrics Preoperative evaluation and management note
C2826012|T102|strict|68594-1|LNC|Plastic surgery Preoperative evaluation and management note|Plastic surgery Preoperative evaluation and management note
C2826012|T102|strict|68835-8|LNC|Primary care Preoperative evaluation and management note|Primary care Preoperative evaluation and management note
C2826012|T102|strict|68844-0|LNC|Speech-language pathology Preoperative evaluation and management note|Speech-language pathology Preoperative evaluation and management note
C2826012|T102|strict|34876-3|LNC|Surgery Preoperative evaluation and management note|Surgery Preoperative evaluation and management note
C2826012|T102|strict|34881-3|LNC|Surgery Nurse Preoperative evaluation and management note|Surgery Nurse Preoperative evaluation and management note
C2826012|T102|strict|68850-7|LNC|Transplant surgery Preoperative evaluation and management note|Transplant surgery Preoperative evaluation and management note
C2826012|T102|strict|34123-0|LNC|Anesthesiology Hospital Preoperative evaluation and management note|Anesthesiology Hospital Preoperative evaluation and management note
C2826012|T102|strict|68828-3|LNC|Pediatrics Hospital Preoperative evaluation and management note|Pediatrics Hospital Preoperative evaluation and management note
C2826012|T102|strict|57832-8|LNC|Prescription for diagnostic or specialist care Document|Prescription for diagnostic or specialist care Document
C2826012|T102|strict|64288-4|LNC|Prescription for eyewear|Prescription for eyewear
C2826012|T102|strict|57829-4|LNC|Prescription for medical equipment or product Document|Prescription for medical equipment or product Document
C2826012|T102|strict|57833-6|LNC|Prescription for medication Document|Prescription for medication Document
C2826012|T102|strict|57831-0|LNC|Prescription for rehabilitation Document|Prescription for rehabilitation Document
C2826012|T102|strict|57828-6|LNC|Prescription list Document|Prescription list Document
C2826012|T102|strict|73709-8|LNC|Prescription request Pharmacy Document from Pharmacist|Prescription request Pharmacy Document from Pharmacist
C2826012|T102|strict|55114-3|LNC|Prior imaging procedure descriptions Document|Prior imaging procedure descriptions Document
C2826012|T102|strict|57017-6|LNC|Privacy policy Organization Document|Privacy policy Organization Document
C2826012|T102|strict|57016-8|LNC|Privacy policy acknowledgment Document|Privacy policy acknowledgment Document
C2826012|T102|strict|64293-4|LNC|Procedure consent|Procedure consent
C2826012|T102|strict|68630-3|LNC|Allergy and immunology procedure note|Allergy and immunology procedure note
C2826012|T102|strict|68658-4|LNC|Clinical genetics procedure note|Clinical genetics procedure note
C2826012|T102|strict|68667-5|LNC|Developmental-behavioral pediatrics procedure note|Developmental-behavioral pediatrics procedure note
C2826012|T102|strict|68692-3|LNC|Neurological surgery procedure note|Neurological surgery procedure note
C2826012|T102|strict|68702-0|LNC|Neurology with special qualifications in child neurology procedure note|Neurology with special qualifications in child neurology procedure note
C2826012|T102|strict|68563-6|LNC|Obstetrics and Gynecology procedure note|Obstetrics and Gynecology procedure note
C2826012|T102|strict|68714-5|LNC|Pain medicine procedure note|Pain medicine procedure note
C2826012|T102|strict|68724-4|LNC|Pediatric cardiology procedure note|Pediatric cardiology procedure note
C2826012|T102|strict|68890-3|LNC|Pediatric dermatology procedure note|Pediatric dermatology procedure note
C2826012|T102|strict|68895-2|LNC|Pediatric endocrinology procedure note|Pediatric endocrinology procedure note
C2826012|T102|strict|68743-4|LNC|Pediatric gastroenterology procedure note|Pediatric gastroenterology procedure note
C2826012|T102|strict|68754-1|LNC|Pediatric hematology-oncology procedure note|Pediatric hematology-oncology procedure note
C2826012|T102|strict|68868-9|LNC|Pediatric nephrology procedure note|Pediatric nephrology procedure note
C2826012|T102|strict|68872-1|LNC|Pediatric otolaryngology procedure note|Pediatric otolaryngology procedure note
C2826012|T102|strict|68784-8|LNC|Pediatric pulmonology procedure note|Pediatric pulmonology procedure note
C2826012|T102|strict|68877-0|LNC|Pediatric rheumatology procedure note|Pediatric rheumatology procedure note
C2826012|T102|strict|68799-6|LNC|Pediatric surgery procedure note|Pediatric surgery procedure note
C2826012|T102|strict|68861-4|LNC|Pediatric transplant hepatology procedure note|Pediatric transplant hepatology procedure note
C2826012|T102|strict|68809-3|LNC|Pediatric urology procedure note|Pediatric urology procedure note
C2826012|T102|strict|68820-0|LNC|Pediatrics procedure note|Pediatrics procedure note
C2826012|T102|strict|68836-6|LNC|Primary care procedure note|Primary care procedure note
C2826012|T102|strict|68851-5|LNC|Transplant surgery procedure note|Transplant surgery procedure note
C2826012|T102|strict|68729-3|LNC|Pediatric critical care medicine Hospital procedure note|Pediatric critical care medicine Hospital procedure note
C2826012|T102|strict|68829-1|LNC|Pediatrics Hospital procedure note|Pediatrics Hospital procedure note
C2826012|T102|strict|68607-1|LNC|Progress letter|Progress letter
C2826012|T102|strict|11506-3|LNC|Provider-unspecified Progress note|Provider-unspecified Progress note
C2826012|T102|strict|68617-0|LNC|Adolescent medicine Progress note|Adolescent medicine Progress note
C2826012|T102|strict|68631-1|LNC|Allergy and immunology Progress note|Allergy and immunology Progress note
C2826012|T102|strict|68646-9|LNC|Child and adolescent psychiatry Progress note|Child and adolescent psychiatry Progress note
C2826012|T102|strict|28580-9|LNC|Chiropractic medicine Progress note|Chiropractic medicine Progress note
C2826012|T102|strict|68659-2|LNC|Clinical genetics Progress note|Clinical genetics Progress note
C2826012|T102|strict|28617-9|LNC|Dentistry Progress note|Dentistry Progress note
C2826012|T102|strict|68668-3|LNC|Developmental-behavioral pediatrics Progress note|Developmental-behavioral pediatrics Progress note
C2826012|T102|strict|34900-1|LNC|General medicine Progress note|General medicine Progress note
C2826012|T102|strict|68554-5|LNC|Hematology+Medical Oncology Progress note|Hematology+Medical Oncology Progress note
C2826012|T102|strict|72556-4|LNC|Interventional radiology Progress note|Interventional radiology Progress note
C2826012|T102|strict|34904-3|LNC|Mental health Progress note|Mental health Progress note
C2826012|T102|strict|68679-0|LNC|Multi-specialty program Progress note|Multi-specialty program Progress note
C2826012|T102|strict|68693-1|LNC|Neurological surgery Progress note|Neurological surgery Progress note
C2826012|T102|strict|68703-8|LNC|Neurology with special qualifications in child neurology Progress note|Neurology with special qualifications in child neurology Progress note
C2826012|T102|strict|28623-7|LNC|Nurse Progress note|Nurse Progress note
C2826012|T102|strict|28575-9|LNC|Nurse practitioner Progress note|Nurse practitioner Progress note
C2826012|T102|strict|68564-4|LNC|Obstetrics and Gynecology Progress note|Obstetrics and Gynecology Progress note
C2826012|T102|strict|11507-1|LNC|Occupational therapy Progress note|Occupational therapy Progress note
C2826012|T102|strict|68574-3|LNC|Ophthalmology Progress note|Ophthalmology Progress note
C2826012|T102|strict|68582-6|LNC|Orthopaedic surgery Progress note|Orthopaedic surgery Progress note
C2826012|T102|strict|68725-1|LNC|Pediatric cardiology Progress note|Pediatric cardiology Progress note
C2826012|T102|strict|68891-1|LNC|Pediatric dermatology Progress note|Pediatric dermatology Progress note
C2826012|T102|strict|68896-0|LNC|Pediatric endocrinology Progress note|Pediatric endocrinology Progress note
C2826012|T102|strict|68744-2|LNC|Pediatric gastroenterology Progress note|Pediatric gastroenterology Progress note
C2826012|T102|strict|68755-8|LNC|Pediatric hematology-oncology Progress note|Pediatric hematology-oncology Progress note
C2826012|T102|strict|68763-2|LNC|Pediatric infectious diseases Progress note|Pediatric infectious diseases Progress note
C2826012|T102|strict|68873-9|LNC|Pediatric otolaryngology Progress note|Pediatric otolaryngology Progress note
C2826012|T102|strict|68785-5|LNC|Pediatric pulmonology Progress note|Pediatric pulmonology Progress note
C2826012|T102|strict|68878-8|LNC|Pediatric rheumatology Progress note|Pediatric rheumatology Progress note
C2826012|T102|strict|68800-2|LNC|Pediatric surgery Progress note|Pediatric surgery Progress note
C2826012|T102|strict|68862-2|LNC|Pediatric transplant hepatology Progress note|Pediatric transplant hepatology Progress note
C2826012|T102|strict|68810-1|LNC|Pediatric urology Progress note|Pediatric urology Progress note
C2826012|T102|strict|11508-9|LNC|Physical therapy Progress note|Physical therapy Progress note
C2826012|T102|strict|18733-6|LNC|Physician attending Progress note|Physician attending Progress note
C2826012|T102|strict|28569-2|LNC|Physician consulting Progress note|Physician consulting Progress note
C2826012|T102|strict|68595-8|LNC|Plastic surgery Progress note|Plastic surgery Progress note
C2826012|T102|strict|11509-7|LNC|Podiatry Progress note|Podiatry Progress note
C2826012|T102|strict|28627-8|LNC|Psychiatry Progress note|Psychiatry Progress note
C2826012|T102|strict|11510-5|LNC|Psychology Progress note|Psychology Progress note
C2826012|T102|strict|68840-8|LNC|Research Progress note|Research Progress note
C2826012|T102|strict|28656-7|LNC|Social work Progress note|Social work Progress note
C2826012|T102|strict|11512-1|LNC|Speech-language pathology Progress note|Speech-language pathology Progress note
C2826012|T102|strict|15507-7|LNC|Provider-unspecified ED Progress note|Provider-unspecified ED Progress note
C2826012|T102|strict|34130-5|LNC|Hospital Progress note|Hospital Progress note
C2826012|T102|strict|68472-0|LNC|Cardiology Hospital Progress note|Cardiology Hospital Progress note
C2826012|T102|strict|68485-2|LNC|Cardiology Medical student Hospital Progress note|Cardiology Medical student Hospital Progress note
C2826012|T102|strict|68484-5|LNC|Cardiology Physician attending Hospital Progress note|Cardiology Physician attending Hospital Progress note
C2826012|T102|strict|64059-9|LNC|Critical Care Medicine Hospital Progress note|Critical Care Medicine Hospital Progress note
C2826012|T102|strict|64071-4|LNC|Critical care medicine Medical student Hospital Progress note|Critical care medicine Medical student Hospital Progress note
C2826012|T102|strict|68473-8|LNC|Critical care medicine Physician attending Hospital Progress note|Critical care medicine Physician attending Hospital Progress note
C2826012|T102|strict|64055-7|LNC|General medicine Medical student Hospital Progress note|General medicine Medical student Hospital Progress note
C2826012|T102|strict|68475-3|LNC|General medicine Physician attending Hospital Progress note|General medicine Physician attending Hospital Progress note
C2826012|T102|strict|68830-9|LNC|Pediatrics Hospital Progress note|Pediatrics Hospital Progress note
C2826012|T102|strict|64063-1|LNC|Pulmonary Hospital Progress note|Pulmonary Hospital Progress note
C2826012|T102|strict|64079-7|LNC|Pulmonary Medical student Hospital Progress note|Pulmonary Medical student Hospital Progress note
C2826012|T102|strict|68478-7|LNC|Pulmonary Physician attending Hospital Progress note|Pulmonary Physician attending Hospital Progress note
C2826012|T102|strict|68479-5|LNC|Respiratory therapy Hospital Progress note|Respiratory therapy Hospital Progress note
C2826012|T102|strict|64057-3|LNC|Surgery Hospital Progress note|Surgery Hospital Progress note
C2826012|T102|strict|64067-2|LNC|Surgery Medical student Hospital Progress note|Surgery Medical student Hospital Progress note
C2826012|T102|strict|68480-3|LNC|Surgery Physician attending Hospital Progress note|Surgery Physician attending Hospital Progress note
C2826012|T102|strict|64061-5|LNC|Thoracic surgery Hospital Progress note|Thoracic surgery Hospital Progress note
C2826012|T102|strict|64075-5|LNC|Thoracic surgery Medical student Hospital Progress note|Thoracic surgery Medical student Hospital Progress note
C2826012|T102|strict|68481-1|LNC|Thoracic surgery Physician attending Hospital Progress note|Thoracic surgery Physician attending Hospital Progress note
C2826012|T102|strict|70238-1|LNC|Transplant surgery Hospital Progress note|Transplant surgery Hospital Progress note
C2826012|T102|strict|34126-3|LNC|Intensive care unit Progress note|Intensive care unit Progress note
C2826012|T102|strict|34131-3|LNC|Outpatient Progress note|Outpatient Progress note
C2826012|T102|strict|34124-8|LNC|Cardiology Outpatient Progress note|Cardiology Outpatient Progress note
C2826012|T102|strict|34128-9|LNC|Dentistry Outpatient Progress note|Dentistry Outpatient Progress note
C2826012|T102|strict|34127-1|LNC|Dentistry Hygienist Outpatient Progress note|Dentistry Hygienist Outpatient Progress note
C2826012|T102|strict|34901-9|LNC|General medicine Outpatient Progress note|General medicine Outpatient Progress note
C2826012|T102|strict|34132-1|LNC|Pharmacy Outpatient Progress note|Pharmacy Outpatient Progress note
C2826012|T102|strict|34129-7|LNC|Patient's home Progress note|Patient's home Progress note
C2826012|T102|strict|34125-5|LNC|Case manager Patient's home Progress note|Case manager Patient's home Progress note
C2826012|T102|strict|74468-0|LNC|Questionnaire form definition section Document|Questionnaire form definition section Document
C2826012|T102|strict|74465-6|LNC|Questionnaire response section Document|Questionnaire response section Document
C2826012|T102|strict|73569-6|LNC|Radiation exposure and protection information [Description] Document Diagnostic imaging|Radiation exposure and protection information [Description] Document Diagnostic imaging
C2826012|T102|strict|64294-2|LNC|Readiness for duty letter|Readiness for duty letter
C2826012|T102|strict|64284-3|LNC|Readiness for duty assessment|Readiness for duty assessment
C2826012|T102|strict|57133-1|LNC|Referral note|Referral note
C2826012|T102|strict|57170-3|LNC|Cardiology Referral note|Cardiology Referral note
C2826012|T102|strict|57178-6|LNC|Critical Care Medicine Referral note|Critical Care Medicine Referral note
C2826012|T102|strict|57134-9|LNC|Dentistry Referral note|Dentistry Referral note
C2826012|T102|strict|57135-6|LNC|Dermatology Referral note|Dermatology Referral note
C2826012|T102|strict|57136-4|LNC|Diabetology Referral note|Diabetology Referral note
C2826012|T102|strict|57137-2|LNC|Endocrinology Referral note|Endocrinology Referral note
C2826012|T102|strict|69438-0|LNC|Referral note Forensic medicine|Referral note Forensic medicine
C2826012|T102|strict|57138-0|LNC|Gastroenterology Referral note|Gastroenterology Referral note
C2826012|T102|strict|57139-8|LNC|General medicine Referral note|General medicine Referral note
C2826012|T102|strict|57171-1|LNC|Geriatric medicine Referral note|Geriatric medicine Referral note
C2826012|T102|strict|57172-9|LNC|Hematology+Medical Oncology Referral note|Hematology+Medical Oncology Referral note
C2826012|T102|strict|57141-4|LNC|Infectious disease Referral note|Infectious disease Referral note
C2826012|T102|strict|57142-2|LNC|Kinesiotherapy Referral note|Kinesiotherapy Referral note
C2826012|T102|strict|57143-0|LNC|Mental health Referral note|Mental health Referral note
C2826012|T102|strict|57144-8|LNC|Nephrology Referral note|Nephrology Referral note
C2826012|T102|strict|57146-3|LNC|Neurological surgery Referral note|Neurological surgery Referral note
C2826012|T102|strict|57145-5|LNC|Neurology Referral note|Neurology Referral note
C2826012|T102|strict|57173-7|LNC|Nutrition and dietetics Referral note|Nutrition and dietetics Referral note
C2826012|T102|strict|57179-4|LNC|Obstetrics and Gynecology Referral note|Obstetrics and Gynecology Referral note
C2826012|T102|strict|57147-1|LNC|Occupational medicine Referral note|Occupational medicine Referral note
C2826012|T102|strict|57148-9|LNC|Occupational therapy Referral note|Occupational therapy Referral note
C2826012|T102|strict|57149-7|LNC|Oncology Referral note|Oncology Referral note
C2826012|T102|strict|57150-5|LNC|Ophthalmology Referral note|Ophthalmology Referral note
C2826012|T102|strict|57151-3|LNC|Optometry Referral note|Optometry Referral note
C2826012|T102|strict|57174-5|LNC|Oral and Maxillofacial Surgery Referral note|Oral and Maxillofacial Surgery Referral note
C2826012|T102|strict|57175-2|LNC|Orthopaedic surgery Referral note|Orthopaedic surgery Referral note
C2826012|T102|strict|57176-0|LNC|Otolaryngology Referral note|Otolaryngology Referral note
C2826012|T102|strict|57152-1|LNC|Pharmacy Referral note|Pharmacy Referral note
C2826012|T102|strict|57153-9|LNC|Physical medicine and rehabilitation Referral note|Physical medicine and rehabilitation Referral note
C2826012|T102|strict|57154-7|LNC|Physical therapy Referral note|Physical therapy Referral note
C2826012|T102|strict|57155-4|LNC|Plastic surgery Referral note|Plastic surgery Referral note
C2826012|T102|strict|57156-2|LNC|Podiatry Referral note|Podiatry Referral note
C2826012|T102|strict|57157-0|LNC|Psychiatry Referral note|Psychiatry Referral note
C2826012|T102|strict|57158-8|LNC|Psychology Referral note|Psychology Referral note
C2826012|T102|strict|57177-8|LNC|Pulmonary Referral note|Pulmonary Referral note
C2826012|T102|strict|57159-6|LNC|Radiation oncology Referral note|Radiation oncology Referral note
C2826012|T102|strict|57160-4|LNC|Recreational therapy Referral note|Recreational therapy Referral note
C2826012|T102|strict|57162-0|LNC|Respiratory therapy Referral note|Respiratory therapy Referral note
C2826012|T102|strict|57163-8|LNC|Rheumatology Referral note|Rheumatology Referral note
C2826012|T102|strict|57164-6|LNC|Social work Referral note|Social work Referral note
C2826012|T102|strict|57165-3|LNC|Speech-language pathology Referral note|Speech-language pathology Referral note
C2826012|T102|strict|57166-1|LNC|Surgery Referral note|Surgery Referral note
C2826012|T102|strict|57167-9|LNC|Thoracic surgery Referral note|Thoracic surgery Referral note
C2826012|T102|strict|57168-7|LNC|Urology Referral note|Urology Referral note
C2826012|T102|strict|57169-5|LNC|Vascular surgery Referral note|Vascular surgery Referral note
C2826012|T102|strict|64292-6|LNC|Release of information consent|Release of information consent
C2826012|T102|strict|55115-0|LNC|Requested imaging studies information Document|Requested imaging studies information Document
C2826012|T102|strict|70007-0|LNC|Restraint note|Restraint note
C2826012|T102|strict|68476-1|LNC|Nurse Hospital Restraint note|Nurse Hospital Restraint note
C2826012|T102|strict|68474-6|LNC|Physician Hospital Restraint note|Physician Hospital Restraint note
C2826012|T102|strict|71482-4|LNC|Risk assessment Document|Risk assessment Document
C2826012|T102|strict|51898-5|LNC|Risk factors Document|Risk factors Document
C2826012|T102|strict|74153-8|LNC|Seizure disorder action plan|Seizure disorder action plan
C2826012|T102|strict|59282-4|LNC|Stress cardiac echo study report US|Stress cardiac echo study report US
C2826012|T102|strict|47045-0|LNC|Study report|Study report
C2826012|T102|strict|68608-9|LNC|Summary note|Summary note
C2826012|T102|strict|61143-4|LNC|Nurse Summary note|Nurse Summary note
C2826012|T102|strict|68602-2|LNC|Radiation oncology Summary note|Radiation oncology Summary note
C2826012|T102|strict|68603-0|LNC|Radiation oncology Hospital Summary note|Radiation oncology Hospital Summary note
C2826012|T102|strict|47046-8|LNC|Summary of death note|Summary of death note
C2826012|T102|strict|34133-9|LNC|Summary of episode note|Summary of episode note
C2826012|T102|strict|74211-4|LNC|Summary of episode note Emergency department+Hospital|Summary of episode note Emergency department+Hospital
C2826012|T102|strict|48764-5|LNC|Summary purpose CCD Document|Summary purpose CCD Document
C2826012|T102|strict|47047-6|LNC|Supervisory note|Supervisory note
C2826012|T102|strict|67865-6|LNC|Outpatient Supervisory note|Outpatient Supervisory note
C2826012|T102|strict|34135-4|LNC|Cardiology Physician attending Outpatient Supervisory note|Cardiology Physician attending Outpatient Supervisory note
C2826012|T102|strict|34136-2|LNC|Gastroenterology Physician attending Outpatient Supervisory note|Gastroenterology Physician attending Outpatient Supervisory note
C2826012|T102|strict|34134-7|LNC|Physician attending Outpatient Supervisory note|Physician attending Outpatient Supervisory note
C2826012|T102|strict|61358-8|LNC|Patient Surgical operation consent|Patient Surgical operation consent
C2826012|T102|strict|11504-8|LNC|Provider-unspecified Operation note|Provider-unspecified Operation note
C2826012|T102|strict|34868-0|LNC|Orthopaedic surgery Surgical operation note|Orthopaedic surgery Surgical operation note
C2826012|T102|strict|34818-5|LNC|Otolaryngology Surgical operation note|Otolaryngology Surgical operation note
C2826012|T102|strict|34870-6|LNC|Plastic surgery Surgical operation note|Plastic surgery Surgical operation note
C2826012|T102|strict|28624-5|LNC|Podiatry Operation note|Podiatry Operation note
C2826012|T102|strict|34874-8|LNC|Surgery Surgical operation note|Surgery Surgical operation note
C2826012|T102|strict|34877-1|LNC|Urology Surgical operation note|Urology Surgical operation note
C2826012|T102|strict|34137-0|LNC|Outpatient Surgical operation note|Outpatient Surgical operation note
C2826012|T102|strict|34138-8|LNC|Targeted history and physical note|Targeted history and physical note
C2826012|T102|strict|18761-7|LNC|Provider-unspecified Transfer summary|Provider-unspecified Transfer summary
C2826012|T102|strict|68618-8|LNC|Adolescent medicine Transfer summary note|Adolescent medicine Transfer summary note
C2826012|T102|strict|68632-9|LNC|Allergy and immunology Transfer summary note|Allergy and immunology Transfer summary note
C2826012|T102|strict|68647-7|LNC|Child and adolescent psychiatry Transfer summary note|Child and adolescent psychiatry Transfer summary note
C2826012|T102|strict|68660-0|LNC|Clinical genetics Transfer summary note|Clinical genetics Transfer summary note
C2826012|T102|strict|34755-9|LNC|Critical care medicine Transfer summary note|Critical care medicine Transfer summary note
C2826012|T102|strict|68669-1|LNC|Developmental-behavioral pediatrics Transfer summary note|Developmental-behavioral pediatrics Transfer summary note
C2826012|T102|strict|34770-8|LNC|General medicine Transfer summary note|General medicine Transfer summary note
C2826012|T102|strict|68680-8|LNC|Multi-specialty program Transfer summary note|Multi-specialty program Transfer summary note
C2826012|T102|strict|68704-6|LNC|Neurology with special qualifications in child neurology Transfer summary note|Neurology with special qualifications in child neurology Transfer summary note
C2826012|T102|strict|68565-1|LNC|Obstetrics and Gynecology Transfer summary note|Obstetrics and Gynecology Transfer summary note
C2826012|T102|strict|68569-3|LNC|Occupational therapy Transfer summary note|Occupational therapy Transfer summary note
C2826012|T102|strict|68887-9|LNC|Ophthalmology Transfer summary note|Ophthalmology Transfer summary note
C2826012|T102|strict|68583-4|LNC|Orthopaedic surgery Transfer summary note|Orthopaedic surgery Transfer summary note
C2826012|T102|strict|68715-2|LNC|Pain medicine Transfer summary note|Pain medicine Transfer summary note
C2826012|T102|strict|68726-9|LNC|Pediatric cardiology Transfer summary note|Pediatric cardiology Transfer summary note
C2826012|T102|strict|68737-6|LNC|Pediatric endocrinology Transfer summary note|Pediatric endocrinology Transfer summary note
C2826012|T102|strict|68745-9|LNC|Pediatric gastroenterology Transfer summary note|Pediatric gastroenterology Transfer summary note
C2826012|T102|strict|68756-6|LNC|Pediatric hematology-oncology Transfer summary note|Pediatric hematology-oncology Transfer summary note
C2826012|T102|strict|68764-0|LNC|Pediatric infectious diseases Transfer summary note|Pediatric infectious diseases Transfer summary note
C2826012|T102|strict|68772-3|LNC|Pediatric nephrology Transfer summary note|Pediatric nephrology Transfer summary note
C2826012|T102|strict|68777-2|LNC|Pediatric otolaryngology Transfer summary note|Pediatric otolaryngology Transfer summary note
C2826012|T102|strict|68786-3|LNC|Pediatric pulmonology Transfer summary note|Pediatric pulmonology Transfer summary note
C2826012|T102|strict|68793-9|LNC|Pediatric rheumatology Transfer summary note|Pediatric rheumatology Transfer summary note
C2826012|T102|strict|68801-0|LNC|Pediatric surgery Transfer summary note|Pediatric surgery Transfer summary note
C2826012|T102|strict|68863-0|LNC|Pediatric transplant hepatology Transfer summary note|Pediatric transplant hepatology Transfer summary note
C2826012|T102|strict|68811-9|LNC|Pediatric urology Transfer summary note|Pediatric urology Transfer summary note
C2826012|T102|strict|68883-8|LNC|Pediatrics Transfer summary note|Pediatrics Transfer summary note
C2826012|T102|strict|68596-6|LNC|Plastic surgery Transfer summary note|Plastic surgery Transfer summary note
C2826012|T102|strict|68482-9|LNC|Nurse Hospital Transfer summary note|Nurse Hospital Transfer summary note
C2826012|T102|strict|68884-6|LNC|Pediatrics Hospital Transfer summary note|Pediatrics Hospital Transfer summary note
C2826012|T102|strict|59281-6|LNC|Transthoracic cardiac echo study report US|Transthoracic cardiac echo study report US
C2826012|T102|strict|74198-3|LNC|Trauma summary registry report Document|Trauma summary registry report Document
C2826012|T102|strict|54094-8|LNC|Emergency department Triage note|Emergency department Triage note
C2826012|T102|strict|57054-9|LNC|Nurse Emergency department Triage+care note|Nurse Emergency department Triage+care note
C2826012|T102|strict|38932-0|LNC|VA Compensation and Pension (C and P) examination acromegaly|VA Compensation and Pension (C and P) examination acromegaly
C2826012|T102|strict|38933-8|LNC|VA Compensation and Pension (C and P) examination aid and attendance/housebound|VA Compensation and Pension (C and P) examination aid and attendance/housebound
C2826012|T102|strict|38934-6|LNC|VA Compensation and Pension (C and P) examination arrhythmias|VA Compensation and Pension (C and P) examination arrhythmias
C2826012|T102|strict|38936-1|LNC|VA Compensation and Pension (C and P) examination audio|VA Compensation and Pension (C and P) examination audio
C2826012|T102|strict|38937-9|LNC|VA Compensation and Pension (C and P) examination bones fractures/bone disease|VA Compensation and Pension (C and P) examination bones fractures/bone disease
C2826012|T102|strict|38938-7|LNC|VA Compensation and Pension (C and P) examination brain/spinal cord|VA Compensation and Pension (C and P) examination brain/spinal cord
C2826012|T102|strict|38939-5|LNC|VA Compensation and Pension (C and P) examination chronic fatigue syndrome|VA Compensation and Pension (C and P) examination chronic fatigue syndrome
C2826012|T102|strict|38940-3|LNC|VA Compensation and Pension (C and P) examination cold injury protocol|VA Compensation and Pension (C and P) examination cold injury protocol
C2826012|T102|strict|38941-1|LNC|VA Compensation and Pension (C and P) examination cranial nerves|VA Compensation and Pension (C and P) examination cranial nerves
C2826012|T102|strict|38942-9|LNC|VA Compensation and Pension (C and P) examination Cushings syndrome|VA Compensation and Pension (C and P) examination Cushings syndrome
C2826012|T102|strict|38943-7|LNC|VA Compensation and Pension (C and P) examination dental/oral|VA Compensation and Pension (C and P) examination dental/oral
C2826012|T102|strict|38944-5|LNC|VA Compensation and Pension (C and P) examination diabetes mellitus|VA Compensation and Pension (C and P) examination diabetes mellitus
C2826012|T102|strict|38956-9|LNC|VA Compensation and Pension (C and P) examination disability in gulf war veterans|VA Compensation and Pension (C and P) examination disability in gulf war veterans
C2826012|T102|strict|38946-0|LNC|VA Compensation and Pension (C and P) examination ear disease|VA Compensation and Pension (C and P) examination ear disease
C2826012|T102|strict|38949-4|LNC|VA Compensation and Pension (C and P) examination epilepsy/narcolepsy|VA Compensation and Pension (C and P) examination epilepsy/narcolepsy
C2826012|T102|strict|38950-2|LNC|VA Compensation and Pension (C and P) examination esophagus/hiatal hernia|VA Compensation and Pension (C and P) examination esophagus/hiatal hernia
C2826012|T102|strict|38966-8|LNC|VA Compensation and Pension (C and P) examination extremity joints|VA Compensation and Pension (C and P) examination extremity joints
C2826012|T102|strict|38951-0|LNC|VA Compensation and Pension (C and P) examination eye|VA Compensation and Pension (C and P) examination eye
C2826012|T102|strict|38952-8|LNC|VA Compensation and Pension (C and P) examination feet|VA Compensation and Pension (C and P) examination feet
C2826012|T102|strict|38953-6|LNC|VA Compensation and Pension (C and P) examination fibromyalgia|VA Compensation and Pension (C and P) examination fibromyalgia
C2826012|T102|strict|38954-4|LNC|VA Compensation and Pension (C and P) examination general medical|VA Compensation and Pension (C and P) examination general medical
C2826012|T102|strict|38969-2|LNC|VA Compensation and Pension (C and P) examination general mental disorders|VA Compensation and Pension (C and P) examination general mental disorders
C2826012|T102|strict|38955-1|LNC|VA Compensation and Pension (C and P) examination genitourinary|VA Compensation and Pension (C and P) examination genitourinary
C2826012|T102|strict|38957-7|LNC|VA Compensation and Pension (C and P) examination gynecological conditions/disorders of the breast|VA Compensation and Pension (C and P) examination gynecological conditions/disorders of the breast
C2826012|T102|strict|38958-5|LNC|VA Compensation and Pension (C and P) examination hand/thumb/fingers|VA Compensation and Pension (C and P) examination hand/thumb/fingers
C2826012|T102|strict|38959-3|LNC|VA Compensation and Pension (C and P) examination heart|VA Compensation and Pension (C and P) examination heart
C2826012|T102|strict|38960-1|LNC|VA Compensation and Pension (C and P) examination hemic disorders|VA Compensation and Pension (C and P) examination hemic disorders
C2826012|T102|strict|38961-9|LNC|VA Compensation and Pension (C and P) examination HIV-related illness|VA Compensation and Pension (C and P) examination HIV-related illness
C2826012|T102|strict|38962-7|LNC|VA Compensation and Pension (C and P) examination hypertension|VA Compensation and Pension (C and P) examination hypertension
C2826012|T102|strict|38963-5|LNC|VA Compensation and Pension (C and P) examination infectious/immune/nutritional disabilities|VA Compensation and Pension (C and P) examination infectious/immune/nutritional disabilities
C2826012|T102|strict|38964-3|LNC|VA Compensation and Pension (C and P) examination initial evaluation post-traumatic stress disorder|VA Compensation and Pension (C and P) examination initial evaluation post-traumatic stress disorder
C2826012|T102|strict|38965-0|LNC|VA Compensation and Pension (C and P) examination large/small intestines|VA Compensation and Pension (C and P) examination large/small intestines
C2826012|T102|strict|38967-6|LNC|VA Compensation and Pension (C and P) examination liver/gall bladder/pancreas|VA Compensation and Pension (C and P) examination liver/gall bladder/pancreas
C2826012|T102|strict|38968-4|LNC|VA Compensation and Pension (C and P) examination lymphatic disorders|VA Compensation and Pension (C and P) examination lymphatic disorders
C2826012|T102|strict|38947-8|LNC|VA Compensation and Pension (C and P) examination mental health eating disorders|VA Compensation and Pension (C and P) examination mental health eating disorders
C2826012|T102|strict|38935-3|LNC|VA Compensation and Pension (C and P) examination miscellaneous arteries/veins|VA Compensation and Pension (C and P) examination miscellaneous arteries/veins
C2826012|T102|strict|38945-2|LNC|VA Compensation and Pension (C and P) examination miscellaneous digestive conditions|VA Compensation and Pension (C and P) examination miscellaneous digestive conditions
C2826012|T102|strict|38948-6|LNC|VA Compensation and Pension (C and P) examination miscellaneous endocrine diseases|VA Compensation and Pension (C and P) examination miscellaneous endocrine diseases
C2826012|T102|strict|38972-6|LNC|VA Compensation and Pension (C and P) examination miscellaneous neurological disorders|VA Compensation and Pension (C and P) examination miscellaneous neurological disorders
C2826012|T102|strict|38980-9|LNC|VA Compensation and Pension (C and P) examination miscellaneous respiratory diseases|VA Compensation and Pension (C and P) examination miscellaneous respiratory diseases
C2826012|T102|strict|38970-0|LNC|VA Compensation and Pension (C and P) examination mouth/lips/tongue|VA Compensation and Pension (C and P) examination mouth/lips/tongue
C2826012|T102|strict|38971-8|LNC|VA Compensation and Pension (C and P) examination muscles|VA Compensation and Pension (C and P) examination muscles
C2826012|T102|strict|38973-4|LNC|VA Compensation and Pension (C and P) examination nose/sinus/larynx/pharynx|VA Compensation and Pension (C and P) examination nose/sinus/larynx/pharynx
C2826012|T102|strict|38979-1|LNC|VA Compensation and Pension (C and P) examination obstructive/restrictive/interstitial respiratory diseases|VA Compensation and Pension (C and P) examination obstructive/restrictive/interstitial respiratory diseases
C2826012|T102|strict|38974-2|LNC|VA Compensation and Pension (C and P) examination peripheral nerves|VA Compensation and Pension (C and P) examination peripheral nerves
C2826012|T102|strict|38975-9|LNC|VA Compensation and Pension (C and P) examination prisoner of war protocol|VA Compensation and Pension (C and P) examination prisoner of war protocol
C2826012|T102|strict|38976-7|LNC|VA Compensation and Pension (C and P) examination pulmonary tuberculosis/mycobacterial diseases|VA Compensation and Pension (C and P) examination pulmonary tuberculosis/mycobacterial diseases
C2826012|T102|strict|38977-5|LNC|VA Compensation and Pension (C and P) examination rectum/anus|VA Compensation and Pension (C and P) examination rectum/anus
C2826012|T102|strict|38978-3|LNC|VA Compensation and Pension (C and P) examination residuals of amputations|VA Compensation and Pension (C and P) examination residuals of amputations
C2826012|T102|strict|38981-7|LNC|VA Compensation and Pension (C and P) examination review evaluation post-traumatic stress disorder|VA Compensation and Pension (C and P) examination review evaluation post-traumatic stress disorder
C2826012|T102|strict|38982-5|LNC|VA Compensation and Pension (C and P) examination scars|VA Compensation and Pension (C and P) examination scars
C2826012|T102|strict|38983-3|LNC|VA Compensation and Pension (C and P) examination sense of smell/taste|VA Compensation and Pension (C and P) examination sense of smell/taste
C2826012|T102|strict|38984-1|LNC|VA Compensation and Pension (C and P) examination skin diseases other than scars|VA Compensation and Pension (C and P) examination skin diseases other than scars
C2826012|T102|strict|38985-8|LNC|VA Compensation and Pension (C and P) examination social/industrial survey|VA Compensation and Pension (C and P) examination social/industrial survey
C2826012|T102|strict|38986-6|LNC|VA Compensation and Pension (C and P) examination spine|VA Compensation and Pension (C and P) examination spine
C2826012|T102|strict|38987-4|LNC|VA Compensation and Pension (C and P) examination stomach/duodenum/peritoneal adhesions|VA Compensation and Pension (C and P) examination stomach/duodenum/peritoneal adhesions
C2826012|T102|strict|38988-2|LNC|VA Compensation and Pension (C and P) examination thyroid/parathyroid diseases|VA Compensation and Pension (C and P) examination thyroid/parathyroid diseases
C2826012|T102|strict|59283-2|LNC|Well child visit note|Well child visit note
C2826012|T102|strict|52027-0|LNC|Abortion consent|Abortion consent
C2826012|T102|strict|24754-4|LNC|Administration of vasodilator into catheter of Vein|Administration of vasodilator into catheter of Vein
C2826012|T102|strict|26376-4|LNC|Administration of vasodilator into catheter of Vein - bilateral|Administration of vasodilator into catheter of Vein - bilateral
C2826012|T102|strict|26377-2|LNC|Administration of vasodilator into catheter of Vein - left|Administration of vasodilator into catheter of Vein - left
C2826012|T102|strict|26378-0|LNC|Administration of vasodilator into catheter of Vein - right|Administration of vasodilator into catheter of Vein - right
C2826012|T102|strict|53243-2|LNC|Advanced beneficiary notice|Advanced beneficiary notice
C2826012|T102|strict|11485-0|LNC|Anesthesia records|Anesthesia records
C2826012|T102|strict|30649-8|LNC|Peripheral artery Fluoroscopic angiogram Additional angioplasty W contrast IA|Peripheral artery Fluoroscopic angiogram Additional angioplasty W contrast IA
C2826012|T102|strict|30641-5|LNC|Vein Fluoroscopic angiogram Additional angioplasty W contrast IV|Vein Fluoroscopic angiogram Additional angioplasty W contrast IV
C2826012|T102|strict|36760-7|LNC|AV shunt Fluoroscopic angiogram Angioplasty W contrast|AV shunt Fluoroscopic angiogram Angioplasty W contrast
C2826012|T102|strict|36762-3|LNC|Extremity vessel Fluoroscopic angiogram Angioplasty W contrast|Extremity vessel Fluoroscopic angiogram Angioplasty W contrast
C2826012|T102|strict|69067-7|LNC|Unspecified body region Fluoroscopic angiogram Angioplasty W contrast|Unspecified body region Fluoroscopic angiogram Angioplasty W contrast
C2826012|T102|strict|24543-1|LNC|Aorta Fluoroscopic angiogram Angioplasty W contrast IA|Aorta Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|24580-3|LNC|Brachiocephalic artery Fluoroscopic angiogram Angioplasty W contrast IA|Brachiocephalic artery Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|26368-1|LNC|Brachiocephalic artery - left Fluoroscopic angiogram Angioplasty W contrast IA|Brachiocephalic artery - left Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|26369-9|LNC|Brachiocephalic artery - right Fluoroscopic angiogram Angioplasty W contrast IA|Brachiocephalic artery - right Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|24614-0|LNC|Carotid artery extracranial Fluoroscopic angiogram Angioplasty W contrast IA|Carotid artery extracranial Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|24615-7|LNC|Carotid artery intracranial Fluoroscopic angiogram Angioplasty W contrast IA|Carotid artery intracranial Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|35881-2|LNC|Extremity artery Fluoroscopic angiogram Angioplasty W contrast IA|Extremity artery Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|24698-3|LNC|Femoral artery Fluoroscopic angiogram Angioplasty W contrast IA|Femoral artery Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|36763-1|LNC|Femoral artery and Popliteal artery Fluoroscopic angiogram Angioplasty W contrast IA|Femoral artery and Popliteal artery Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|24766-8|LNC|Iliac artery Fluoroscopic angiogram Angioplasty W contrast IA|Iliac artery Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|26370-7|LNC|Iliac artery - bilateral Fluoroscopic angiogram Angioplasty W contrast IA|Iliac artery - bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|26371-5|LNC|Iliac artery - left Fluoroscopic angiogram Angioplasty W contrast IA|Iliac artery - left Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|26372-3|LNC|Iliac artery - right Fluoroscopic angiogram Angioplasty W contrast IA|Iliac artery - right Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|24832-8|LNC|Mesenteric artery Fluoroscopic angiogram Angioplasty W contrast IA|Mesenteric artery Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|30648-0|LNC|Peripheral artery Fluoroscopic angiogram Angioplasty W contrast IA|Peripheral artery Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|25081-1|LNC|Renal vessel Fluoroscopic angiogram Angioplasty W contrast IA|Renal vessel Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|25012-6|LNC|Tibial artery Fluoroscopic angiogram Angioplasty W contrast IA|Tibial artery Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|26373-1|LNC|Tibial artery - bilateral Fluoroscopic angiogram Angioplasty W contrast IA|Tibial artery - bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|26374-9|LNC|Tibial artery - left Fluoroscopic angiogram Angioplasty W contrast IA|Tibial artery - left Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|26375-6|LNC|Tibial artery - right Fluoroscopic angiogram Angioplasty W contrast IA|Tibial artery - right Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|43793-9|LNC|Tibioperoneal arteries Fluoroscopic angiogram Angioplasty W contrast IA|Tibioperoneal arteries Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|43794-7|LNC|Tibioperoneal arteries - bilateral Fluoroscopic angiogram Angioplasty W contrast IA|Tibioperoneal arteries - bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|43795-4|LNC|Tibioperoneal arteries - left Fluoroscopic angiogram Angioplasty W contrast IA|Tibioperoneal arteries - left Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|43792-1|LNC|Tibioperoneal arteries - right Fluoroscopic angiogram Angioplasty W contrast IA|Tibioperoneal arteries - right Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|25064-7|LNC|Vessel Fluoroscopic angiogram Angioplasty W contrast IA|Vessel Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|30836-1|LNC|Visceral artery Fluoroscopic angiogram Angioplasty W contrast IA|Visceral artery Fluoroscopic angiogram Angioplasty W contrast IA
C2826012|T102|strict|37426-4|LNC|Lower extremity vein Fluoroscopic angiogram Angioplasty W contrast IV|Lower extremity vein Fluoroscopic angiogram Angioplasty W contrast IV
C2826012|T102|strict|30640-7|LNC|Vein Fluoroscopic angiogram Angioplasty W contrast IV|Vein Fluoroscopic angiogram Angioplasty W contrast IV
C2826012|T102|strict|35882-0|LNC|Inferior vena cava Fluoroscopic angiogram Angioplasty W contrast IV|Inferior vena cava Fluoroscopic angiogram Angioplasty W contrast IV
C2826012|T102|strict|52032-0|LNC|Appeal denial letter|Appeal denial letter
C2826012|T102|strict|36764-9|LNC|Femoral vessel and Popliteal artery Fluoroscopic angiogram Atherectomy W contrast|Femoral vessel and Popliteal artery Fluoroscopic angiogram Atherectomy W contrast
C2826012|T102|strict|69135-2|LNC|Iliac artery Fluoroscopic angiogram Atherectomy W contrast|Iliac artery Fluoroscopic angiogram Atherectomy W contrast
C2826012|T102|strict|69253-3|LNC|Renal vessels Fluoroscopic angiogram Atherectomy W contrast|Renal vessels Fluoroscopic angiogram Atherectomy W contrast
C2826012|T102|strict|36765-6|LNC|Vessel Fluoroscopic angiogram Atherectomy W contrast|Vessel Fluoroscopic angiogram Atherectomy W contrast
C2826012|T102|strict|35883-8|LNC|Aorta Fluoroscopic angiogram Atherectomy W contrast IA|Aorta Fluoroscopic angiogram Atherectomy W contrast IA
C2826012|T102|strict|36766-4|LNC|Coronary arteries Fluoroscopic angiogram Atherectomy W contrast IA|Coronary arteries Fluoroscopic angiogram Atherectomy W contrast IA
C2826012|T102|strict|24568-8|LNC|AV fistula Fluoroscopic angiogram Atherectomy W contrast IV|AV fistula Fluoroscopic angiogram Atherectomy W contrast IV
C2826012|T102|strict|28615-3|LNC|Audiology study|Audiology study
C2826012|T102|strict|52065-0|LNC|Automobile liability|Automobile liability
C2826012|T102|strict|18743-5|LNC|Autopsy report|Autopsy report
C2826012|T102|strict|36761-5|LNC|Biliary ducts Fluoroscopy Balloon dilatation W contrast|Biliary ducts Fluoroscopy Balloon dilatation W contrast
C2826012|T102|strict|33720-4|LNC|Blood bank consult|Blood bank consult
C2826012|T102|strict|52041-1|LNC|Blood glucose monitors|Blood glucose monitors
C2826012|T102|strict|38268-9|LNC|Skeletal system DXA Bone density|Skeletal system DXA Bone density
C2826012|T102|strict|43562-8|LNC|Skeletal system.axial Scan Bone density|Skeletal system.axial Scan Bone density
C2826012|T102|strict|43563-6|LNC|Skeletal system.peripheral Scan Bone density|Skeletal system.peripheral Scan Bone density
C2826012|T102|strict|48807-2|LNC|Bone marrow aspiration report|Bone marrow aspiration report
C2826012|T102|strict|24631-4|LNC|Unspecified body region Fluoroscopy Central vein catheter placement check|Unspecified body region Fluoroscopy Central vein catheter placement check
C2826012|T102|strict|53242-4|LNC|Charge ticket or encounter form|Charge ticket or encounter form
C2826012|T102|strict|54095-5|LNC|Chemotherapy effectiveness panel [Identifier] - Blood or Tissue|Chemotherapy effectiveness panel [Identifier] - Blood or Tissue
C2826012|T102|strict|11486-8|LNC|Chemotherapy records|Chemotherapy records
C2826012|T102|strict|71428-7|LNC|CMS - history of present illness panel|CMS - history of present illness panel
C2826012|T102|strict|71421-2|LNC|CMS - past family - social history panel|CMS - past family - social history panel
C2826012|T102|strict|71388-3|LNC|CMS - physical exam panel|CMS - physical exam panel
C2826012|T102|strict|71406-3|LNC|CMS - review of systems panel|CMS - review of systems panel
C2826012|T102|strict|25062-1|LNC|Unspecified body region X-ray Comparison view|Unspecified body region X-ray Comparison view
C2826012|T102|strict|24611-6|LNC|Outpatient Consultation 2nd opinion|Outpatient Consultation 2nd opinion
C2826012|T102|strict|60570-9|LNC|Pathology Consult note|Pathology Consult note
C2826012|T102|strict|60571-7|LNC|Pathology Consult note.synoptic|Pathology Consult note.synoptic
C2826012|T102|strict|52042-9|LNC|Continuous positive airway pressure (CPAP)|Continuous positive airway pressure (CPAP)
C2826012|T102|strict|25038-1|LNC|Unspecified body region Courtesy consultation|Unspecified body region Courtesy consultation
C2826012|T102|strict|29751-5|LNC|Critical care records|Critical care records
C2826012|T102|strict|50007-4|LNC|Cytology report of Bronchoalveolar lavage Cyto stain|Cytology report of Bronchoalveolar lavage Cyto stain
C2826012|T102|strict|47523-6|LNC|Cytology report of Body fluid Cyto stain|Cytology report of Body fluid Cyto stain
C2826012|T102|strict|47530-1|LNC|Cytology report of Breast ductal lavage Cyto stain|Cytology report of Breast ductal lavage Cyto stain
C2826012|T102|strict|47521-0|LNC|Cytology report of Breast fine needle aspirate Cyto stain|Cytology report of Breast fine needle aspirate Cyto stain
C2826012|T102|strict|50971-1|LNC|Cytology report of Bronchial brush Cyto stain|Cytology report of Bronchial brush Cyto stain
C2826012|T102|strict|47528-5|LNC|Cytology report of Cervical or vaginal smear or scraping Cyto stain|Cytology report of Cervical or vaginal smear or scraping Cyto stain
C2826012|T102|strict|47527-7|LNC|Cytology report of Cervical or vaginal smear or scraping Cyto stain.thin prep|Cytology report of Cervical or vaginal smear or scraping Cyto stain.thin prep
C2826012|T102|strict|47522-8|LNC|Cytology report of Nipple discharge Cyto stain|Cytology report of Nipple discharge Cyto stain
C2826012|T102|strict|47520-2|LNC|Cytology report of Sputum Cyto stain|Cytology report of Sputum Cyto stain
C2826012|T102|strict|47524-4|LNC|Cytology report of Thyroid fine needle aspirate Cyto stain|Cytology report of Thyroid fine needle aspirate Cyto stain
C2826012|T102|strict|47529-3|LNC|Cytology report of Tissue Other stain|Cytology report of Tissue Other stain
C2826012|T102|strict|33718-8|LNC|Cytology report of Tissue fine needle aspirate Cyto stain|Cytology report of Tissue fine needle aspirate Cyto stain
C2826012|T102|strict|47525-1|LNC|Cytology report of Urine Cyto stain|Cytology report of Urine Cyto stain
C2826012|T102|strict|47526-9|LNC|Cytology report of Unspecified specimen Cyto stain|Cytology report of Unspecified specimen Cyto stain
C2826012|T102|strict|52040-3|LNC|Dental X-rays and other images (not DICOM)|Dental X-rays and other images (not DICOM)
C2826012|T102|strict|29749-9|LNC|Dialysis records|Dialysis records
C2826012|T102|strict|28622-9|LNC|Nurse Discharge assessment|Nurse Discharge assessment
C2826012|T102|strict|28574-2|LNC|Discharge note|Discharge note
C2826012|T102|strict|29761-4|LNC|Dentist Discharge summary|Dentist Discharge summary
C2826012|T102|strict|11490-0|LNC|Physician Discharge summary|Physician Discharge summary
C2826012|T102|strict|28655-9|LNC|Physician attending Discharge summary|Physician attending Discharge summary
C2826012|T102|strict|53245-7|LNC|Driver license image|Driver license image
C2826012|T102|strict|53247-3|LNC|Eligibility acknowledgement|Eligibility acknowledgement
C2826012|T102|strict|24684-3|LNC|Extracranial vessels Fluoroscopic angiogram Embolectomy W contrast IA|Extracranial vessels Fluoroscopic angiogram Embolectomy W contrast IA
C2826012|T102|strict|24887-2|LNC|Pulmonary artery Fluoroscopic angiogram Embolectomy W contrast IA|Pulmonary artery Fluoroscopic angiogram Embolectomy W contrast IA
C2826012|T102|strict|24553-0|LNC|Vessel intracranial Fluoroscopic angiogram Embolectomy W contrast IV|Vessel intracranial Fluoroscopic angiogram Embolectomy W contrast IV
C2826012|T102|strict|24554-8|LNC|Artery Fluoroscopic angiogram Embolization W contrast IA|Artery Fluoroscopic angiogram Embolization W contrast IA
C2826012|T102|strict|52071-8|LNC|Employee assistance program|Employee assistance program
C2826012|T102|strict|67796-3|LNC|EMS patient care report - version 3.1 Document NEMSIS|EMS patient care report - version 3.1 Document NEMSIS
C2826012|T102|strict|52043-7|LNC|Enteral nutrition|Enteral nutrition
C2826012|T102|strict|30600-1|LNC|Small bowel CT Views Enteroclysis W contrast PO via duodenal intubation|Small bowel CT Views Enteroclysis W contrast PO via duodenal intubation
C2826012|T102|strict|24923-5|LNC|Small bowel Fluoroscopy Views Enteroclysis W contrast PO via duodenal intubation|Small bowel Fluoroscopy Views Enteroclysis W contrast PO via duodenal intubation
C2826012|T102|strict|52030-4|LNC|Explanation of benefits|Explanation of benefits
C2826012|T102|strict|52031-2|LNC|Explanation of benefits to subscriber|Explanation of benefits to subscriber
C2826012|T102|strict|52044-5|LNC|External infusion pump|External infusion pump
C2826012|T102|strict|29272-2|LNC|Eye ultrasound study|Eye ultrasound study
C2826012|T102|strict|52064-3|LNC|First report of injury|First report of injury
C2826012|T102|strict|57129-9|LNC|Full newborn screening summary report for display or printing|Full newborn screening summary report for display or printing
C2826012|T102|strict|52045-2|LNC|Gait trainers|Gait trainers
C2826012|T102|strict|52033-8|LNC|General correspondence|General correspondence
C2826012|T102|strict|51969-4|LNC|Genetic analysis summary report in Blood or Tissue Document by Molecular genetics method|Genetic analysis summary report in Blood or Tissue Document by Molecular genetics method
C2826012|T102|strict|46365-3|LNC|CT Guidance for ablation of tissue of Celiac plexus|CT Guidance for ablation of tissue of Celiac plexus
C2826012|T102|strict|44228-5|LNC|CT Guidance for ablation of tissue of Kidney|CT Guidance for ablation of tissue of Kidney
C2826012|T102|strict|44156-8|LNC|US Guidance for ablation of tissue of Kidney|US Guidance for ablation of tissue of Kidney
C2826012|T102|strict|44101-4|LNC|CT Guidance for ablation of tissue of Liver|CT Guidance for ablation of tissue of Liver
C2826012|T102|strict|44155-0|LNC|US Guidance for ablation of tissue of Liver|US Guidance for ablation of tissue of Liver
C2826012|T102|strict|58747-7|LNC|CT Guidance for ablation of tissue of Unspecified body region|CT Guidance for ablation of tissue of Unspecified body region
C2826012|T102|strict|58743-6|LNC|US Guidance for ablation of tissue of Unspecified body region|US Guidance for ablation of tissue of Unspecified body region
C2826012|T102|strict|35884-6|LNC|CT Guidance for abscess drainage of Abdomen|CT Guidance for abscess drainage of Abdomen
C2826012|T102|strict|42280-8|LNC|CT Guidance for abscess drainage of Appendix|CT Guidance for abscess drainage of Appendix
C2826012|T102|strict|42705-4|LNC|US Guidance for abscess drainage of Appendix|US Guidance for abscess drainage of Appendix
C2826012|T102|strict|42281-6|LNC|CT Guidance for abscess drainage of Chest|CT Guidance for abscess drainage of Chest
C2826012|T102|strict|42285-7|LNC|CT Guidance for abscess drainage of Kidney|CT Guidance for abscess drainage of Kidney
C2826012|T102|strict|44167-5|LNC|US Guidance for abscess drainage of Kidney|US Guidance for abscess drainage of Kidney
C2826012|T102|strict|42282-4|LNC|CT Guidance for abscess drainage of Liver|CT Guidance for abscess drainage of Liver
C2826012|T102|strict|42133-9|LNC|US Guidance for abscess drainage of Liver|US Guidance for abscess drainage of Liver
C2826012|T102|strict|39361-1|LNC|Fluoroscopy Guidance for abscess drainage of Liver|Fluoroscopy Guidance for abscess drainage of Liver
C2826012|T102|strict|69120-4|LNC|Fluoroscopy Guidance for abscess drainage of Neck|Fluoroscopy Guidance for abscess drainage of Neck
C2826012|T102|strict|69122-0|LNC|Fluoroscopy Guidance for abscess drainage of Pancreas|Fluoroscopy Guidance for abscess drainage of Pancreas
C2826012|T102|strict|42286-5|LNC|CT Guidance for abscess drainage of Pelvis|CT Guidance for abscess drainage of Pelvis
C2826012|T102|strict|44168-3|LNC|US Guidance for abscess drainage of Pelvis|US Guidance for abscess drainage of Pelvis
C2826012|T102|strict|44169-1|LNC|US Guidance for abscess drainage of Peritoneal space|US Guidance for abscess drainage of Peritoneal space
C2826012|T102|strict|42284-0|LNC|CT Guidance for abscess drainage of Pleural space|CT Guidance for abscess drainage of Pleural space
C2826012|T102|strict|69123-8|LNC|Fluoroscopy Guidance for abscess drainage of Pleural space|Fluoroscopy Guidance for abscess drainage of Pleural space
C2826012|T102|strict|43502-4|LNC|CT Guidance for abscess drainage of Subphrenic space|CT Guidance for abscess drainage of Subphrenic space
C2826012|T102|strict|44166-7|LNC|US Guidance for abscess drainage of Subphrenic space|US Guidance for abscess drainage of Subphrenic space
C2826012|T102|strict|30578-9|LNC|CT Guidance for abscess drainage of Unspecified body region|CT Guidance for abscess drainage of Unspecified body region
C2826012|T102|strict|39451-0|LNC|US Guidance for abscess drainage of Unspecified body region|US Guidance for abscess drainage of Unspecified body region
C2826012|T102|strict|35885-3|LNC|Fluoroscopy Guidance for abscess drainage of Unspecified body region|Fluoroscopy Guidance for abscess drainage of Unspecified body region
C2826012|T102|strict|39620-0|LNC|Scan Guidance for abscess localization limited|Scan Guidance for abscess localization limited
C2826012|T102|strict|39623-4|LNC|Scan Guidance for abscess localization whole body|Scan Guidance for abscess localization whole body
C2826012|T102|strict|39622-6|LNC|SPECT Guidance for abscess localization whole body|SPECT Guidance for abscess localization whole body
C2826012|T102|strict|39621-8|LNC|SPECT Guidance for abscess localization|SPECT Guidance for abscess localization
C2826012|T102|strict|72533-3|LNC|US Guidance for ambulatory phlebectomy of Extremity vein - left|US Guidance for ambulatory phlebectomy of Extremity vein - left
C2826012|T102|strict|72532-5|LNC|US Guidance for ambulatory phlebectomy of Extremity vein - right|US Guidance for ambulatory phlebectomy of Extremity vein - right
C2826012|T102|strict|24623-1|LNC|CT Guidance for anesthetic block injection of Celiac plexus|CT Guidance for anesthetic block injection of Celiac plexus
C2826012|T102|strict|42688-2|LNC|CT Guidance for anesthetic block injection of Spine|CT Guidance for anesthetic block injection of Spine
C2826012|T102|strict|35886-1|LNC|CT Guidance for aspiration of Breast|CT Guidance for aspiration of Breast
C2826012|T102|strict|24598-5|LNC|Mammogram Guidance for aspiration of Breast|Mammogram Guidance for aspiration of Breast
C2826012|T102|strict|43756-6|LNC|US Guidance for aspiration of Breast|US Guidance for aspiration of Breast
C2826012|T102|strict|69278-0|LNC|US Guidance for aspiration of Breast - bilateral|US Guidance for aspiration of Breast - bilateral
C2826012|T102|strict|69292-1|LNC|US Guidance for aspiration of Breast - left|US Guidance for aspiration of Breast - left
C2826012|T102|strict|69296-2|LNC|US Guidance for aspiration of Breast - right|US Guidance for aspiration of Breast - right
C2826012|T102|strict|35888-7|LNC|Fluoroscopy Guidance for aspiration of Hip|Fluoroscopy Guidance for aspiration of Hip
C2826012|T102|strict|24771-8|LNC|Fluoroscopy Guidance for aspiration of Joint space|Fluoroscopy Guidance for aspiration of Joint space
C2826012|T102|strict|48434-5|LNC|US Guidance for aspiration of Kidney|US Guidance for aspiration of Kidney
C2826012|T102|strict|24811-2|LNC|CT Guidance for aspiration of Liver|CT Guidance for aspiration of Liver
C2826012|T102|strict|24822-9|LNC|CT Guidance for aspiration of Lung|CT Guidance for aspiration of Lung
C2826012|T102|strict|69287-1|LNC|US Guidance for aspiration of Lymph node|US Guidance for aspiration of Lymph node
C2826012|T102|strict|24837-7|LNC|CT Guidance for aspiration of Neck|CT Guidance for aspiration of Neck
C2826012|T102|strict|39452-8|LNC|US Guidance for aspiration of Ovary|US Guidance for aspiration of Ovary
C2826012|T102|strict|24856-7|LNC|CT Guidance for aspiration of Pancreas|CT Guidance for aspiration of Pancreas
C2826012|T102|strict|24863-3|LNC|CT Guidance for aspiration of Pelvis|CT Guidance for aspiration of Pelvis
C2826012|T102|strict|30703-3|LNC|US Guidance for aspiration of Pericardial space|US Guidance for aspiration of Pericardial space
C2826012|T102|strict|37491-8|LNC|CT Guidance for aspiration of Pleural space|CT Guidance for aspiration of Pleural space
C2826012|T102|strict|24662-9|LNC|US Guidance for aspiration of Pleural space|US Guidance for aspiration of Pleural space
C2826012|T102|strict|37887-7|LNC|Fluoroscopy Guidance for aspiration of Pleural space|Fluoroscopy Guidance for aspiration of Pleural space
C2826012|T102|strict|24973-0|LNC|Fluoroscopy Guidance for aspiration of Spine Lumbar Space|Fluoroscopy Guidance for aspiration of Spine Lumbar Space
C2826012|T102|strict|42134-7|LNC|US Guidance for aspiration of Thyroid|US Guidance for aspiration of Thyroid
C2826012|T102|strict|25043-1|LNC|CT Guidance for aspiration of Unspecified body region|CT Guidance for aspiration of Unspecified body region
C2826012|T102|strict|30878-3|LNC|US Guidance for aspiration of Unspecified body region|US Guidance for aspiration of Unspecified body region
C2826012|T102|strict|36926-4|LNC|CT Guidance for aspiration and placement of drainage tube of Abdomen|CT Guidance for aspiration and placement of drainage tube of Abdomen
C2826012|T102|strict|37210-2|LNC|CT Guidance for aspiration of cyst of Abdomen|CT Guidance for aspiration of cyst of Abdomen
C2826012|T102|strict|69306-9|LNC|Fluoroscopy Guidance for aspiration of cyst of Bone|Fluoroscopy Guidance for aspiration of cyst of Bone
C2826012|T102|strict|24594-4|LNC|Mammogram Guidance for aspiration of cyst of Breast|Mammogram Guidance for aspiration of cyst of Breast
C2826012|T102|strict|69192-3|LNC|MRI Guidance for aspiration of cyst of Breast|MRI Guidance for aspiration of cyst of Breast
C2826012|T102|strict|30653-0|LNC|US Guidance for aspiration of cyst of Breast|US Guidance for aspiration of cyst of Breast
C2826012|T102|strict|26343-4|LNC|Mammogram Guidance for aspiration of cyst of Breast - bilateral|Mammogram Guidance for aspiration of cyst of Breast - bilateral
C2826012|T102|strict|38012-1|LNC|US Guidance for aspiration of cyst of Breast - bilateral|US Guidance for aspiration of cyst of Breast - bilateral
C2826012|T102|strict|26344-2|LNC|Mammogram Guidance for aspiration of cyst of Breast - left|Mammogram Guidance for aspiration of cyst of Breast - left
C2826012|T102|strict|42450-7|LNC|US Guidance for aspiration of cyst of Breast - left|US Guidance for aspiration of cyst of Breast - left
C2826012|T102|strict|26345-9|LNC|Mammogram Guidance for aspiration of cyst of Breast - right|Mammogram Guidance for aspiration of cyst of Breast - right
C2826012|T102|strict|42458-0|LNC|US Guidance for aspiration of cyst of Breast - right|US Guidance for aspiration of cyst of Breast - right
C2826012|T102|strict|38126-9|LNC|US Guidance for aspiration of cyst of Kidney|US Guidance for aspiration of cyst of Kidney
C2826012|T102|strict|69121-2|LNC|Fluoroscopy Guidance for aspiration of cyst of Ovary|Fluoroscopy Guidance for aspiration of cyst of Ovary
C2826012|T102|strict|38133-5|LNC|US Guidance for aspiration of cyst of Pancreas|US Guidance for aspiration of cyst of Pancreas
C2826012|T102|strict|42447-3|LNC|US Guidance for aspiration of cyst of Thyroid|US Guidance for aspiration of cyst of Thyroid
C2826012|T102|strict|35887-9|LNC|CT Guidance for aspiration of cyst of Unspecified body region|CT Guidance for aspiration of cyst of Unspecified body region
C2826012|T102|strict|30698-5|LNC|US Guidance for aspiration of cyst of Unspecified body region|US Guidance for aspiration of cyst of Unspecified body region
C2826012|T102|strict|24671-0|LNC|Fluoroscopy Guidance for aspiration of cyst of Unspecified body region|Fluoroscopy Guidance for aspiration of cyst of Unspecified body region
C2826012|T102|strict|25042-3|LNC|CT Guidance for aspiration or biopsy of Unspecified body region|CT Guidance for aspiration or biopsy of Unspecified body region
C2826012|T102|strict|25041-5|LNC|CT Guidance for aspiration or biopsy of Unspecified body region-- W contrast IV|CT Guidance for aspiration or biopsy of Unspecified body region-- W contrast IV
C2826012|T102|strict|46281-2|LNC|CT Guidance for aspiration or injection of cyst of Unspecified body region|CT Guidance for aspiration or injection of cyst of Unspecified body region
C2826012|T102|strict|46282-0|LNC|US Guidance for aspiration or injection of cyst of Unspecified body region|US Guidance for aspiration or injection of cyst of Unspecified body region
C2826012|T102|strict|30602-7|LNC|CT Guidance for fine needle aspiration of Abdomen|CT Guidance for fine needle aspiration of Abdomen
C2826012|T102|strict|44107-1|LNC|CT Guidance for fine needle aspiration of Abdomen retroperitoneum|CT Guidance for fine needle aspiration of Abdomen retroperitoneum
C2826012|T102|strict|44108-9|LNC|CT Guidance for fine needle aspiration of Adrenal gland|CT Guidance for fine needle aspiration of Adrenal gland
C2826012|T102|strict|46387-7|LNC|Mammogram Guidance for fine needle aspiration of Breast|Mammogram Guidance for fine needle aspiration of Breast
C2826012|T102|strict|44160-0|LNC|US Guidance for fine needle aspiration of Breast|US Guidance for fine needle aspiration of Breast
C2826012|T102|strict|46284-6|LNC|Mammogram Guidance for fine needle aspiration of Breast - left|Mammogram Guidance for fine needle aspiration of Breast - left
C2826012|T102|strict|38026-1|LNC|US Guidance for fine needle aspiration of Breast - left|US Guidance for fine needle aspiration of Breast - left
C2826012|T102|strict|46283-8|LNC|Mammogram Guidance for fine needle aspiration of Breast - right|Mammogram Guidance for fine needle aspiration of Breast - right
C2826012|T102|strict|38033-7|LNC|US Guidance for fine needle aspiration of Breast - right|US Guidance for fine needle aspiration of Breast - right
C2826012|T102|strict|38135-0|LNC|US Guidance for fine needle aspiration of Deep tissue|US Guidance for fine needle aspiration of Deep tissue
C2826012|T102|strict|44221-0|LNC|Fluoroscopy Guidance for fine needle aspiration of Deep tissue|Fluoroscopy Guidance for fine needle aspiration of Deep tissue
C2826012|T102|strict|43757-4|LNC|CT Guidance for fine needle aspiration of Kidney|CT Guidance for fine needle aspiration of Kidney
C2826012|T102|strict|44159-2|LNC|US Guidance for fine needle aspiration of Kidney|US Guidance for fine needle aspiration of Kidney
C2826012|T102|strict|44217-8|LNC|Fluoroscopy Guidance for fine needle aspiration of Kidney|Fluoroscopy Guidance for fine needle aspiration of Kidney
C2826012|T102|strict|30608-4|LNC|CT Guidance for fine needle aspiration of Kidney - bilateral|CT Guidance for fine needle aspiration of Kidney - bilateral
C2826012|T102|strict|30603-5|LNC|CT Guidance for fine needle aspiration of Liver|CT Guidance for fine needle aspiration of Liver
C2826012|T102|strict|44158-4|LNC|US Guidance for fine needle aspiration of Liver|US Guidance for fine needle aspiration of Liver
C2826012|T102|strict|44220-2|LNC|Fluoroscopy Guidance for fine needle aspiration of Liver|Fluoroscopy Guidance for fine needle aspiration of Liver
C2826012|T102|strict|30595-3|LNC|CT Guidance for fine needle aspiration of Lung|CT Guidance for fine needle aspiration of Lung
C2826012|T102|strict|44103-0|LNC|CT Guidance for fine needle aspiration of Lymph node|CT Guidance for fine needle aspiration of Lymph node
C2826012|T102|strict|44219-4|LNC|Fluoroscopy Guidance for fine needle aspiration of Lymph node|Fluoroscopy Guidance for fine needle aspiration of Lymph node
C2826012|T102|strict|44104-8|LNC|CT Guidance for fine needle aspiration of Mediastinum|CT Guidance for fine needle aspiration of Mediastinum
C2826012|T102|strict|44105-5|LNC|CT Guidance for fine needle aspiration of Muscle|CT Guidance for fine needle aspiration of Muscle
C2826012|T102|strict|30605-0|LNC|CT Guidance for fine needle aspiration of Pancreas|CT Guidance for fine needle aspiration of Pancreas
C2826012|T102|strict|44157-6|LNC|US Guidance for fine needle aspiration of Pancreas|US Guidance for fine needle aspiration of Pancreas
C2826012|T102|strict|44218-6|LNC|Fluoroscopy Guidance for fine needle aspiration of Pancreas|Fluoroscopy Guidance for fine needle aspiration of Pancreas
C2826012|T102|strict|30606-8|LNC|CT Guidance for fine needle aspiration of Pelvis|CT Guidance for fine needle aspiration of Pelvis
C2826012|T102|strict|44106-3|LNC|CT Guidance for fine needle aspiration of Prostate|CT Guidance for fine needle aspiration of Prostate
C2826012|T102|strict|38017-0|LNC|US Guidance for fine needle aspiration of Prostate|US Guidance for fine needle aspiration of Prostate
C2826012|T102|strict|30610-0|LNC|CT Guidance for fine needle aspiration of Spleen|CT Guidance for fine needle aspiration of Spleen
C2826012|T102|strict|38136-8|LNC|US Guidance for fine needle aspiration of Superficial tissue|US Guidance for fine needle aspiration of Superficial tissue
C2826012|T102|strict|69124-6|LNC|Fluoroscopy Guidance for fine needle aspiration of Superficial tissue|Fluoroscopy Guidance for fine needle aspiration of Superficial tissue
C2826012|T102|strict|38019-6|LNC|US Guidance for fine needle aspiration of Thyroid|US Guidance for fine needle aspiration of Thyroid
C2826012|T102|strict|44216-0|LNC|Fluoroscopy Guidance for fine needle aspiration of Thyroid|Fluoroscopy Guidance for fine needle aspiration of Thyroid
C2826012|T102|strict|30580-5|LNC|CT Guidance for fine needle aspiration of Unspecified body region|CT Guidance for fine needle aspiration of Unspecified body region
C2826012|T102|strict|38018-8|LNC|US Guidance for fine needle aspiration of Unspecified body region|US Guidance for fine needle aspiration of Unspecified body region
C2826012|T102|strict|44215-2|LNC|Fluoroscopy Guidance for fine needle aspiration of Unspecified body region|Fluoroscopy Guidance for fine needle aspiration of Unspecified body region
C2826012|T102|strict|24755-1|LNC|Fluoroscopic angiogram Guidance for atherectomy of Vein-- W contrast IV|Fluoroscopic angiogram Guidance for atherectomy of Vein-- W contrast IV
C2826012|T102|strict|26298-0|LNC|Fluoroscopic angiogram Guidance for atherectomy of Vein - bilateral-- W contrast IV|Fluoroscopic angiogram Guidance for atherectomy of Vein - bilateral-- W contrast IV
C2826012|T102|strict|26299-8|LNC|Fluoroscopic angiogram Guidance for atherectomy of Vein - left-- W contrast IV|Fluoroscopic angiogram Guidance for atherectomy of Vein - left-- W contrast IV
C2826012|T102|strict|26300-4|LNC|Fluoroscopic angiogram Guidance for atherectomy of Vein - right-- W contrast IV|Fluoroscopic angiogram Guidance for atherectomy of Vein - right-- W contrast IV
C2826012|T102|strict|30601-9|LNC|CT Guidance for biopsy of Abdomen|CT Guidance for biopsy of Abdomen
C2826012|T102|strict|37913-1|LNC|US Guidance for biopsy of Abdomen|US Guidance for biopsy of Abdomen
C2826012|T102|strict|35890-3|LNC|Fluoroscopy Guidance for biopsy of Abdomen|Fluoroscopy Guidance for biopsy of Abdomen
C2826012|T102|strict|44117-0|LNC|CT Guidance for biopsy of Abdomen retroperitoneum|CT Guidance for biopsy of Abdomen retroperitoneum
C2826012|T102|strict|44162-6|LNC|US Guidance for biopsy of Abdomen retroperitoneum|US Guidance for biopsy of Abdomen retroperitoneum
C2826012|T102|strict|36767-2|LNC|CT Guidance for biopsy of Adrenal gland|CT Guidance for biopsy of Adrenal gland
C2826012|T102|strict|35891-1|LNC|CT Guidance for biopsy of Bone|CT Guidance for biopsy of Bone
C2826012|T102|strict|69076-8|LNC|Fluoroscopy Guidance for biopsy of Bone|Fluoroscopy Guidance for biopsy of Bone
C2826012|T102|strict|37211-0|LNC|CT Guidance for biopsy of Bone marrow|CT Guidance for biopsy of Bone marrow
C2826012|T102|strict|35893-7|LNC|CT Guidance for biopsy of Breast|CT Guidance for biopsy of Breast
C2826012|T102|strict|24602-5|LNC|Mammogram Guidance for biopsy of Breast|Mammogram Guidance for biopsy of Breast
C2826012|T102|strict|37914-9|LNC|US Guidance for biopsy of Breast|US Guidance for biopsy of Breast
C2826012|T102|strict|26337-6|LNC|Mammogram Guidance for biopsy of Breast - bilateral|Mammogram Guidance for biopsy of Breast - bilateral
C2826012|T102|strict|69169-1|LNC|MRI Guidance for biopsy of Breast - bilateral|MRI Guidance for biopsy of Breast - bilateral
C2826012|T102|strict|37912-3|LNC|US Guidance for biopsy of Breast - bilateral|US Guidance for biopsy of Breast - bilateral
C2826012|T102|strict|26338-4|LNC|Mammogram Guidance for biopsy of Breast - left|Mammogram Guidance for biopsy of Breast - left
C2826012|T102|strict|69203-8|LNC|MRI Guidance for biopsy of Breast - left|MRI Guidance for biopsy of Breast - left
C2826012|T102|strict|42449-9|LNC|US Guidance for biopsy of Breast - left|US Guidance for biopsy of Breast - left
C2826012|T102|strict|26339-2|LNC|Mammogram Guidance for biopsy of Breast - right|Mammogram Guidance for biopsy of Breast - right
C2826012|T102|strict|69213-7|LNC|MRI Guidance for biopsy of Breast - right|MRI Guidance for biopsy of Breast - right
C2826012|T102|strict|42457-2|LNC|US Guidance for biopsy of Breast - right|US Guidance for biopsy of Breast - right
C2826012|T102|strict|35895-2|LNC|CT Guidance for biopsy of Chest|CT Guidance for biopsy of Chest
C2826012|T102|strict|37915-6|LNC|US Guidance for biopsy of Chest|US Guidance for biopsy of Chest
C2826012|T102|strict|35894-5|LNC|Fluoroscopy Guidance for biopsy of Chest|Fluoroscopy Guidance for biopsy of Chest
C2826012|T102|strict|37492-6|LNC|CT Guidance for biopsy of Chest.pleura|CT Guidance for biopsy of Chest.pleura
C2826012|T102|strict|42333-5|LNC|US Guidance for biopsy of Chest.pleura|US Guidance for biopsy of Chest.pleura
C2826012|T102|strict|43567-7|LNC|CT Guidance for biopsy of Deep bone|CT Guidance for biopsy of Deep bone
C2826012|T102|strict|43565-1|LNC|US Guidance for biopsy of Deep bone|US Guidance for biopsy of Deep bone
C2826012|T102|strict|44109-7|LNC|CT Guidance for biopsy of Deep muscle|CT Guidance for biopsy of Deep muscle
C2826012|T102|strict|42463-0|LNC|US Guidance for biopsy of Endomyocardium|US Guidance for biopsy of Endomyocardium
C2826012|T102|strict|37212-8|LNC|CT Guidance for biopsy of Epididymis|CT Guidance for biopsy of Epididymis
C2826012|T102|strict|69387-9|LNC|US Guidance for biopsy of Epididymis|US Guidance for biopsy of Epididymis
C2826012|T102|strict|36927-2|LNC|CT Guidance for biopsy of Facial bones and Maxilla|CT Guidance for biopsy of Facial bones and Maxilla
C2826012|T102|strict|35892-9|LNC|CT Guidance for biopsy of Head|CT Guidance for biopsy of Head
C2826012|T102|strict|42136-2|LNC|CT Guidance for biopsy of Heart|CT Guidance for biopsy of Heart
C2826012|T102|strict|42279-0|LNC|CT Guidance for biopsy of Kidney|CT Guidance for biopsy of Kidney
C2826012|T102|strict|24772-6|LNC|US Guidance for biopsy of Kidney|US Guidance for biopsy of Kidney
C2826012|T102|strict|35899-4|LNC|Fluoroscopy Guidance for biopsy of Kidney|Fluoroscopy Guidance for biopsy of Kidney
C2826012|T102|strict|38766-2|LNC|US Guidance for biopsy of Kidney transplant|US Guidance for biopsy of Kidney transplant
C2826012|T102|strict|30607-6|LNC|CT Guidance for biopsy of Kidney - bilateral|CT Guidance for biopsy of Kidney - bilateral
C2826012|T102|strict|26340-0|LNC|US Guidance for biopsy of Kidney - bilateral|US Guidance for biopsy of Kidney - bilateral
C2826012|T102|strict|26341-8|LNC|US Guidance for biopsy of Kidney - left|US Guidance for biopsy of Kidney - left
C2826012|T102|strict|26342-6|LNC|US Guidance for biopsy of Kidney - right|US Guidance for biopsy of Kidney - right
C2826012|T102|strict|24812-0|LNC|CT Guidance for biopsy of Liver|CT Guidance for biopsy of Liver
C2826012|T102|strict|24816-1|LNC|US Guidance for biopsy of Liver|US Guidance for biopsy of Liver
C2826012|T102|strict|35900-0|LNC|Fluoroscopy Guidance for biopsy of Liver|Fluoroscopy Guidance for biopsy of Liver
C2826012|T102|strict|38765-4|LNC|US Guidance for biopsy of Liver transplant|US Guidance for biopsy of Liver transplant
C2826012|T102|strict|35896-0|LNC|CT Guidance for biopsy of Lower extremity|CT Guidance for biopsy of Lower extremity
C2826012|T102|strict|24823-7|LNC|CT Guidance for biopsy of Lung|CT Guidance for biopsy of Lung
C2826012|T102|strict|44161-8|LNC|US Guidance for biopsy of Lung|US Guidance for biopsy of Lung
C2826012|T102|strict|30634-0|LNC|Fluoroscopy Guidance for biopsy of Lung|Fluoroscopy Guidance for biopsy of Lung
C2826012|T102|strict|35901-8|LNC|CT Guidance for biopsy of Lymph node|CT Guidance for biopsy of Lymph node
C2826012|T102|strict|39522-8|LNC|US Guidance for biopsy of Lymph node|US Guidance for biopsy of Lymph node
C2826012|T102|strict|37213-6|LNC|CT Guidance for biopsy of Mediastinum|CT Guidance for biopsy of Mediastinum
C2826012|T102|strict|42137-0|LNC|US Guidance for biopsy of Mediastinum|US Guidance for biopsy of Mediastinum
C2826012|T102|strict|36768-0|LNC|CT Guidance for biopsy of Muscle|CT Guidance for biopsy of Muscle
C2826012|T102|strict|37917-2|LNC|US Guidance for biopsy of Muscle|US Guidance for biopsy of Muscle
C2826012|T102|strict|24838-5|LNC|CT Guidance for biopsy of Neck|CT Guidance for biopsy of Neck
C2826012|T102|strict|37918-0|LNC|US Guidance for biopsy of Neck|US Guidance for biopsy of Neck
C2826012|T102|strict|30604-3|LNC|CT Guidance for biopsy of Pancreas|CT Guidance for biopsy of Pancreas
C2826012|T102|strict|37919-8|LNC|US Guidance for biopsy of Pancreas|US Guidance for biopsy of Pancreas
C2826012|T102|strict|35902-6|LNC|Fluoroscopy Guidance for biopsy of Pancreas|Fluoroscopy Guidance for biopsy of Pancreas
C2826012|T102|strict|24864-1|LNC|CT Guidance for biopsy of Pelvis|CT Guidance for biopsy of Pelvis
C2826012|T102|strict|69074-3|LNC|Fluoroscopy Guidance for biopsy of Pelvis|Fluoroscopy Guidance for biopsy of Pelvis
C2826012|T102|strict|35903-4|LNC|CT Guidance for biopsy of Prostate|CT Guidance for biopsy of Prostate
C2826012|T102|strict|24883-1|LNC|US Guidance for biopsy of Prostate|US Guidance for biopsy of Prostate
C2826012|T102|strict|41802-0|LNC|Fluoroscopy Guidance for biopsy of Prostate|Fluoroscopy Guidance for biopsy of Prostate
C2826012|T102|strict|35898-6|LNC|CT Guidance for biopsy of Salivary gland|CT Guidance for biopsy of Salivary gland
C2826012|T102|strict|37920-6|LNC|US Guidance for biopsy of Salivary gland|US Guidance for biopsy of Salivary gland
C2826012|T102|strict|69075-0|LNC|Fluoroscopy Guidance for biopsy of Salivary gland|Fluoroscopy Guidance for biopsy of Salivary gland
C2826012|T102|strict|38132-7|LNC|US Guidance for biopsy of Scrotum and Testicle|US Guidance for biopsy of Scrotum and Testicle
C2826012|T102|strict|69396-0|LNC|US Guidance for biopsy of Spinal cord|US Guidance for biopsy of Spinal cord
C2826012|T102|strict|24986-2|LNC|CT Guidance for biopsy of Spine|CT Guidance for biopsy of Spine
C2826012|T102|strict|35904-2|LNC|CT Guidance for biopsy of Spine Cervical|CT Guidance for biopsy of Spine Cervical
C2826012|T102|strict|35905-9|LNC|CT Guidance for biopsy of Spine Lumbar|CT Guidance for biopsy of Spine Lumbar
C2826012|T102|strict|35906-7|LNC|CT Guidance for biopsy of Spine Thoracic|CT Guidance for biopsy of Spine Thoracic
C2826012|T102|strict|30609-2|LNC|CT Guidance for biopsy of Spleen|CT Guidance for biopsy of Spleen
C2826012|T102|strict|35907-5|LNC|Fluoroscopy Guidance for biopsy of Spleen|Fluoroscopy Guidance for biopsy of Spleen
C2826012|T102|strict|42265-9|LNC|CT Guidance for biopsy of Superficial bone|CT Guidance for biopsy of Superficial bone
C2826012|T102|strict|42135-4|LNC|US Guidance for biopsy of Superficial bone|US Guidance for biopsy of Superficial bone
C2826012|T102|strict|38154-1|LNC|Fluoroscopy Guidance for biopsy of Superficial bone|Fluoroscopy Guidance for biopsy of Superficial bone
C2826012|T102|strict|43797-0|LNC|US Guidance for biopsy of Superficial lymph node|US Guidance for biopsy of Superficial lymph node
C2826012|T102|strict|43564-4|LNC|US Guidance for biopsy of Superficial muscle|US Guidance for biopsy of Superficial muscle
C2826012|T102|strict|37214-4|LNC|CT Guidance for biopsy of Superficial tissue|CT Guidance for biopsy of Superficial tissue
C2826012|T102|strict|35908-3|LNC|CT Guidance for biopsy of Thyroid|CT Guidance for biopsy of Thyroid
C2826012|T102|strict|25009-2|LNC|US Guidance for biopsy of Thyroid|US Guidance for biopsy of Thyroid
C2826012|T102|strict|35897-8|LNC|CT Guidance for biopsy of Upper extremity|CT Guidance for biopsy of Upper extremity
C2826012|T102|strict|25044-9|LNC|CT Guidance for biopsy of Unspecified body region|CT Guidance for biopsy of Unspecified body region
C2826012|T102|strict|25059-7|LNC|US Guidance for biopsy of Unspecified body region|US Guidance for biopsy of Unspecified body region
C2826012|T102|strict|25069-6|LNC|Fluoroscopy Guidance for biopsy of Unspecified body region|Fluoroscopy Guidance for biopsy of Unspecified body region
C2826012|T102|strict|24670-2|LNC|US Guidance for biopsy of cyst of Unspecified body region|US Guidance for biopsy of cyst of Unspecified body region
C2826012|T102|strict|30651-4|LNC|US Guidance for core needle biopsy of Breast|US Guidance for core needle biopsy of Breast
C2826012|T102|strict|24813-8|LNC|CT Guidance for core needle biopsy of Liver|CT Guidance for core needle biopsy of Liver
C2826012|T102|strict|69279-8|LNC|US Guidance for core needle biopsy of Lymph node|US Guidance for core needle biopsy of Lymph node
C2826012|T102|strict|46285-3|LNC|US Guidance for core needle biopsy of Thyroid|US Guidance for core needle biopsy of Thyroid
C2826012|T102|strict|38024-6|LNC|US Guidance for core needle biopsy of Unspecified body region|US Guidance for core needle biopsy of Unspecified body region
C2826012|T102|strict|69073-5|LNC|Fluoroscopy Guidance for core needle biopsy of Unspecified body region|Fluoroscopy Guidance for core needle biopsy of Unspecified body region
C2826012|T102|strict|42448-1|LNC|US Guidance for excisional biopsy of Breast|US Guidance for excisional biopsy of Breast
C2826012|T102|strict|30652-2|LNC|US Guidance for fine needle biopsy of Breast|US Guidance for fine needle biopsy of Breast
C2826012|T102|strict|42288-1|LNC|CT Guidance for needle biopsy of Abdomen|CT Guidance for needle biopsy of Abdomen
C2826012|T102|strict|69224-4|LNC|Fluoroscopy Guidance for needle biopsy of Abdomen|Fluoroscopy Guidance for needle biopsy of Abdomen
C2826012|T102|strict|46367-9|LNC|CT Guidance for needle biopsy of Adrenal gland|CT Guidance for needle biopsy of Adrenal gland
C2826012|T102|strict|46368-7|LNC|CT Guidance for needle biopsy of Breast|CT Guidance for needle biopsy of Breast
C2826012|T102|strict|46286-1|LNC|Mammogram Guidance for needle biopsy of Breast|Mammogram Guidance for needle biopsy of Breast
C2826012|T102|strict|38028-7|LNC|US Guidance for needle biopsy of Breast|US Guidance for needle biopsy of Breast
C2826012|T102|strict|41803-8|LNC|Fluoroscopy Guidance for needle biopsy of Breast|Fluoroscopy Guidance for needle biopsy of Breast
C2826012|T102|strict|43462-1|LNC|US Guidance for needle biopsy of Breast - left|US Guidance for needle biopsy of Breast - left
C2826012|T102|strict|43447-2|LNC|Mammogram Guidance for needle biopsy of Breast - right|Mammogram Guidance for needle biopsy of Breast - right
C2826012|T102|strict|69290-5|LNC|US Guidance for needle biopsy of Breast - right|US Guidance for needle biopsy of Breast - right
C2826012|T102|strict|38029-5|LNC|US Guidance for needle biopsy of Chest|US Guidance for needle biopsy of Chest
C2826012|T102|strict|69225-1|LNC|Fluoroscopy Guidance for needle biopsy of Chest|Fluoroscopy Guidance for needle biopsy of Chest
C2826012|T102|strict|69099-0|LNC|CT Guidance for needle biopsy of Chest.pleura|CT Guidance for needle biopsy of Chest.pleura
C2826012|T102|strict|44171-7|LNC|US Guidance for needle biopsy of Chest.pleura|US Guidance for needle biopsy of Chest.pleura
C2826012|T102|strict|69127-9|LNC|Fluoroscopy Guidance for needle biopsy of Chest.pleura|Fluoroscopy Guidance for needle biopsy of Chest.pleura
C2826012|T102|strict|43568-5|LNC|CT Guidance for needle biopsy of Deep bone|CT Guidance for needle biopsy of Deep bone
C2826012|T102|strict|42289-9|LNC|CT Guidance for needle biopsy of Kidney|CT Guidance for needle biopsy of Kidney
C2826012|T102|strict|38027-9|LNC|US Guidance for needle biopsy of Kidney - bilateral|US Guidance for needle biopsy of Kidney - bilateral
C2826012|T102|strict|69097-4|LNC|CT Guidance for needle biopsy of Liver|CT Guidance for needle biopsy of Liver
C2826012|T102|strict|69197-2|LNC|MRI Guidance for needle biopsy of Liver|MRI Guidance for needle biopsy of Liver
C2826012|T102|strict|44170-9|LNC|US Guidance for needle biopsy of Liver|US Guidance for needle biopsy of Liver
C2826012|T102|strict|69125-3|LNC|Fluoroscopy Guidance for needle biopsy of Liver|Fluoroscopy Guidance for needle biopsy of Liver
C2826012|T102|strict|42267-5|LNC|CT Guidance for needle biopsy of Lymph node|CT Guidance for needle biopsy of Lymph node
C2826012|T102|strict|37916-4|LNC|US Guidance for needle biopsy of Lymph node|US Guidance for needle biopsy of Lymph node
C2826012|T102|strict|69098-2|LNC|CT Guidance for needle biopsy of Muscle|CT Guidance for needle biopsy of Muscle
C2826012|T102|strict|69198-0|LNC|MRI Guidance for needle biopsy of Muscle|MRI Guidance for needle biopsy of Muscle
C2826012|T102|strict|69288-9|LNC|US Guidance for needle biopsy of Muscle|US Guidance for needle biopsy of Muscle
C2826012|T102|strict|69226-9|LNC|Fluoroscopy Guidance for needle biopsy of Muscle|Fluoroscopy Guidance for needle biopsy of Muscle
C2826012|T102|strict|46369-5|LNC|US Guidance for needle biopsy of Ovary|US Guidance for needle biopsy of Ovary
C2826012|T102|strict|42290-7|LNC|CT Guidance for needle biopsy of Pancreas|CT Guidance for needle biopsy of Pancreas
C2826012|T102|strict|69199-8|LNC|MRI Guidance for needle biopsy of Pancreas|MRI Guidance for needle biopsy of Pancreas
C2826012|T102|strict|69289-7|LNC|US Guidance for needle biopsy of Pancreas|US Guidance for needle biopsy of Pancreas
C2826012|T102|strict|69126-1|LNC|Fluoroscopy Guidance for needle biopsy of Pancreas|Fluoroscopy Guidance for needle biopsy of Pancreas
C2826012|T102|strict|46370-3|LNC|US Guidance for needle biopsy of Pelvis|US Guidance for needle biopsy of Pelvis
C2826012|T102|strict|69200-4|LNC|MRI Guidance for needle biopsy of Pleura|MRI Guidance for needle biopsy of Pleura
C2826012|T102|strict|69227-7|LNC|Fluoroscopy Guidance for needle biopsy of Pleura|Fluoroscopy Guidance for needle biopsy of Pleura
C2826012|T102|strict|46288-7|LNC|US Guidance for needle biopsy of Prostate|US Guidance for needle biopsy of Prostate
C2826012|T102|strict|69228-5|LNC|Fluoroscopy Guidance for needle biopsy of Prostate|Fluoroscopy Guidance for needle biopsy of Prostate
C2826012|T102|strict|69100-6|LNC|CT Guidance for needle biopsy of Salivary gland|CT Guidance for needle biopsy of Salivary gland
C2826012|T102|strict|69201-2|LNC|MRI Guidance for needle biopsy of Salivary gland|MRI Guidance for needle biopsy of Salivary gland
C2826012|T102|strict|69291-3|LNC|US Guidance for needle biopsy of Salivary gland|US Guidance for needle biopsy of Salivary gland
C2826012|T102|strict|69128-7|LNC|Fluoroscopy Guidance for needle biopsy of Salivary gland|Fluoroscopy Guidance for needle biopsy of Salivary gland
C2826012|T102|strict|43571-9|LNC|CT Guidance for needle biopsy of Soft bone|CT Guidance for needle biopsy of Soft bone
C2826012|T102|strict|69401-8|LNC|US Guidance for needle biopsy of Spinal cord|US Guidance for needle biopsy of Spinal cord
C2826012|T102|strict|38030-3|LNC|US Guidance for needle biopsy of Spleen|US Guidance for needle biopsy of Spleen
C2826012|T102|strict|42266-7|LNC|CT Guidance for needle biopsy of Superficial bone|CT Guidance for needle biopsy of Superficial bone
C2826012|T102|strict|69101-4|LNC|CT Guidance for needle biopsy of Thyroid|CT Guidance for needle biopsy of Thyroid
C2826012|T102|strict|69202-0|LNC|MRI Guidance for needle biopsy of Thyroid|MRI Guidance for needle biopsy of Thyroid
C2826012|T102|strict|38031-1|LNC|US Guidance for needle biopsy of Thyroid|US Guidance for needle biopsy of Thyroid
C2826012|T102|strict|69129-5|LNC|Fluoroscopy Guidance for needle biopsy of Thyroid|Fluoroscopy Guidance for needle biopsy of Thyroid
C2826012|T102|strict|46287-9|LNC|CT Guidance for needle biopsy of Unspecified body region|CT Guidance for needle biopsy of Unspecified body region
C2826012|T102|strict|30700-9|LNC|US Guidance for needle biopsy of Unspecified body region|US Guidance for needle biopsy of Unspecified body region
C2826012|T102|strict|44225-1|LNC|Fluoroscopy Guidance for needle biopsy of Liver-- W contrast IV|Fluoroscopy Guidance for needle biopsy of Liver-- W contrast IV
C2826012|T102|strict|24718-9|LNC|Fluoroscopy Guidance for transjugular biopsy of Liver-- W contrast IV|Fluoroscopy Guidance for transjugular biopsy of Liver-- W contrast IV
C2826012|T102|strict|35910-9|LNC|CT Guidance for biopsy of Chest-- W and WO contrast IV|CT Guidance for biopsy of Chest-- W and WO contrast IV
C2826012|T102|strict|46289-5|LNC|CT Guidance for biopsy of Unspecified body region-- W and WO contrast IV|CT Guidance for biopsy of Unspecified body region-- W and WO contrast IV
C2826012|T102|strict|35909-1|LNC|CT Guidance for biopsy of Chest-- W contrast IV|CT Guidance for biopsy of Chest-- W contrast IV
C2826012|T102|strict|69093-3|LNC|CT Guidance for biopsy of Pelvis-- W contrast IV|CT Guidance for biopsy of Pelvis-- W contrast IV
C2826012|T102|strict|42260-0|LNC|CT Guidance for biopsy of Unspecified body region-- W contrast IV|CT Guidance for biopsy of Unspecified body region-- W contrast IV
C2826012|T102|strict|46366-1|LNC|SPECT Guidance for biopsy of Bone|SPECT Guidance for biopsy of Bone
C2826012|T102|strict|46384-4|LNC|SPECT Guidance for biopsy of Superficial bone|SPECT Guidance for biopsy of Superficial bone
C2826012|T102|strict|69083-4|LNC|CT Guidance for biopsy of Abdomen-- WO contrast|CT Guidance for biopsy of Abdomen-- WO contrast
C2826012|T102|strict|35911-7|LNC|CT Guidance for biopsy of Chest-- WO contrast|CT Guidance for biopsy of Chest-- WO contrast
C2826012|T102|strict|69092-5|LNC|CT Guidance for biopsy of Liver-- WO contrast|CT Guidance for biopsy of Liver-- WO contrast
C2826012|T102|strict|69094-1|LNC|CT Guidance for biopsy of Pelvis-- WO contrast|CT Guidance for biopsy of Pelvis-- WO contrast
C2826012|T102|strict|46290-3|LNC|CT Guidance for biopsy of Unspecified body region-- WO contrast|CT Guidance for biopsy of Unspecified body region-- WO contrast
C2826012|T102|strict|35889-5|LNC|Fluoroscopy Guidance for bronchoscopy of Chest|Fluoroscopy Guidance for bronchoscopy of Chest
C2826012|T102|strict|64998-8|LNC|Fluoroscopy Guidance for catheterization of Fallopian tube - left-- transcervical|Fluoroscopy Guidance for catheterization of Fallopian tube - left-- transcervical
C2826012|T102|strict|64999-6|LNC|Fluoroscopy Guidance for catheterization of Fallopian tube -right-- transcervical|Fluoroscopy Guidance for catheterization of Fallopian tube -right-- transcervical
C2826012|T102|strict|30818-9|LNC|Fluoroscopy Guidance for catheterization of Fallopian tubes-- transcervical|Fluoroscopy Guidance for catheterization of Fallopian tubes-- transcervical
C2826012|T102|strict|30892-4|LNC|Fluoroscopy Guidance for catheterization of Biliary ducts and Pancreatic duct-- W contrast retrograde|Fluoroscopy Guidance for catheterization of Biliary ducts and Pancreatic duct-- W contrast retrograde
C2826012|T102|strict|24624-9|LNC|Fluoroscopic angiogram Guidance for change of central catheter in Central vein-- W contrast IV|Fluoroscopic angiogram Guidance for change of central catheter in Central vein-- W contrast IV
C2826012|T102|strict|26331-9|LNC|Fluoroscopic angiogram Guidance for change of central catheter in Central vein - bilateral-- W contrast IV|Fluoroscopic angiogram Guidance for change of central catheter in Central vein - bilateral-- W contrast IV
C2826012|T102|strict|26332-7|LNC|Fluoroscopic angiogram Guidance for change of central catheter in Central vein - left-- W contrast IV|Fluoroscopic angiogram Guidance for change of central catheter in Central vein - left-- W contrast IV
C2826012|T102|strict|26333-5|LNC|Fluoroscopic angiogram Guidance for change of central catheter in Central vein - right-- W contrast IV|Fluoroscopic angiogram Guidance for change of central catheter in Central vein - right-- W contrast IV
C2826012|T102|strict|43558-6|LNC|Fluoroscopy Guidance for change of dialysis catheter in Unspecified body region-- W contrast IV|Fluoroscopy Guidance for change of dialysis catheter in Unspecified body region-- W contrast IV
C2826012|T102|strict|36769-8|LNC|CT Guidance for change of nephrostomy tube in Kidney|CT Guidance for change of nephrostomy tube in Kidney
C2826012|T102|strict|24781-7|LNC|Fluoroscopy Guidance for change of percutaneous nephrostomy tube in Kidney - bilateral-- W contrast|Fluoroscopy Guidance for change of percutaneous nephrostomy tube in Kidney - bilateral-- W contrast
C2826012|T102|strict|46371-1|LNC|X-ray Guidance for change of percutaneous tube in Unspecified body region-- W contrast|X-ray Guidance for change of percutaneous tube in Unspecified body region-- W contrast
C2826012|T102|strict|30646-4|LNC|Fluoroscopy Guidance for change of tube in Sinus tract-- W contrast|Fluoroscopy Guidance for change of tube in Sinus tract-- W contrast
C2826012|T102|strict|69400-0|LNC|US Guidance for chorionic villus sampling|US Guidance for chorionic villus sampling
C2826012|T102|strict|69391-1|LNC|US Guidance for cordocentesis|US Guidance for cordocentesis
C2826012|T102|strict|38127-7|LNC|US Guidance for CSF aspiration of Spine|US Guidance for CSF aspiration of Spine
C2826012|T102|strict|70915-4|LNC|US Guidance for CSF aspiration of Spine Cervical|US Guidance for CSF aspiration of Spine Cervical
C2826012|T102|strict|70916-2|LNC|US Guidance for CSF aspiration of Spine Lumbar|US Guidance for CSF aspiration of Spine Lumbar
C2826012|T102|strict|70917-0|LNC|US Guidance for CSF aspiration of Spine Thoracic|US Guidance for CSF aspiration of Spine Thoracic
C2826012|T102|strict|24680-1|LNC|Fluoroscopy Guidance for dilation of Esophagus|Fluoroscopy Guidance for dilation of Esophagus
C2826012|T102|strict|35913-3|LNC|CT Guidance for drainage of Abdomen|CT Guidance for drainage of Abdomen
C2826012|T102|strict|42287-3|LNC|CT Guidance for drainage of Abdomen retroperitoneum|CT Guidance for drainage of Abdomen retroperitoneum
C2826012|T102|strict|41809-5|LNC|US Guidance for drainage of Abdomen retroperitoneum|US Guidance for drainage of Abdomen retroperitoneum
C2826012|T102|strict|35914-1|LNC|CT Guidance for drainage of Anus|CT Guidance for drainage of Anus
C2826012|T102|strict|35915-8|LNC|CT Guidance for drainage of Appendix|CT Guidance for drainage of Appendix
C2826012|T102|strict|36770-6|LNC|CT Guidance for drainage of Biliary ducts and Gallbladder|CT Guidance for drainage of Biliary ducts and Gallbladder
C2826012|T102|strict|35916-6|LNC|CT Guidance for drainage of Chest|CT Guidance for drainage of Chest
C2826012|T102|strict|69078-4|LNC|Fluoroscopy Guidance for drainage of Chest|Fluoroscopy Guidance for drainage of Chest
C2826012|T102|strict|24692-6|LNC|US Guidance for drainage of Extremity|US Guidance for drainage of Extremity
C2826012|T102|strict|26325-1|LNC|US Guidance for drainage of Extremity - bilateral|US Guidance for drainage of Extremity - bilateral
C2826012|T102|strict|26326-9|LNC|US Guidance for drainage of Extremity - left|US Guidance for drainage of Extremity - left
C2826012|T102|strict|26327-7|LNC|US Guidance for drainage of Extremity - right|US Guidance for drainage of Extremity - right
C2826012|T102|strict|35917-4|LNC|CT Guidance for drainage of Gallbladder|CT Guidance for drainage of Gallbladder
C2826012|T102|strict|69133-7|LNC|Fluoroscopy Guidance for drainage of Hip|Fluoroscopy Guidance for drainage of Hip
C2826012|T102|strict|35918-2|LNC|CT Guidance for drainage of Kidney|CT Guidance for drainage of Kidney
C2826012|T102|strict|24896-3|LNC|US Guidance for drainage of Kidney|US Guidance for drainage of Kidney
C2826012|T102|strict|26328-5|LNC|US Guidance for drainage of Kidney - bilateral|US Guidance for drainage of Kidney - bilateral
C2826012|T102|strict|26329-3|LNC|US Guidance for drainage of Kidney - left|US Guidance for drainage of Kidney - left
C2826012|T102|strict|26330-1|LNC|US Guidance for drainage of Kidney - right|US Guidance for drainage of Kidney - right
C2826012|T102|strict|35919-0|LNC|CT Guidance for drainage of Liver|CT Guidance for drainage of Liver
C2826012|T102|strict|35920-8|LNC|CT Guidance for drainage of Lymph node|CT Guidance for drainage of Lymph node
C2826012|T102|strict|42283-2|LNC|CT Guidance for drainage of Pancreas|CT Guidance for drainage of Pancreas
C2826012|T102|strict|44172-5|LNC|US Guidance for drainage of Pancreas|US Guidance for drainage of Pancreas
C2826012|T102|strict|35921-6|LNC|CT Guidance for drainage of Pelvis|CT Guidance for drainage of Pelvis
C2826012|T102|strict|24868-2|LNC|US Guidance for drainage of Pelvis|US Guidance for drainage of Pelvis
C2826012|T102|strict|41800-4|LNC|Fluoroscopy Guidance for drainage of Pharynx|Fluoroscopy Guidance for drainage of Pharynx
C2826012|T102|strict|41798-0|LNC|US Guidance for drainage of Prostate|US Guidance for drainage of Prostate
C2826012|T102|strict|35922-4|LNC|CT Guidance for drainage of Unspecified body region|CT Guidance for drainage of Unspecified body region
C2826012|T102|strict|30699-3|LNC|US Guidance for drainage of Unspecified body region|US Guidance for drainage of Unspecified body region
C2826012|T102|strict|43537-0|LNC|Fluoroscopy Guidance for drainage of Unspecified body region|Fluoroscopy Guidance for drainage of Unspecified body region
C2826012|T102|strict|42478-8|LNC|US Guidance for drainage of cyst of Kidney|US Guidance for drainage of cyst of Kidney
C2826012|T102|strict|46291-1|LNC|CT Guidance for drainage of Unspecified body region-- W and WO contrast IV|CT Guidance for drainage of Unspecified body region-- W and WO contrast IV
C2826012|T102|strict|35923-2|LNC|CT Guidance for drainage of Chest-- W contrast IV|CT Guidance for drainage of Chest-- W contrast IV
C2826012|T102|strict|46292-9|LNC|CT Guidance for drainage of Unspecified body region-- W contrast IV|CT Guidance for drainage of Unspecified body region-- W contrast IV
C2826012|T102|strict|35924-0|LNC|CT Guidance for drainage of Chest-- WO contrast|CT Guidance for drainage of Chest-- WO contrast
C2826012|T102|strict|46293-7|LNC|CT Guidance for drainage of Unspecified body region-- WO contrast|CT Guidance for drainage of Unspecified body region-- WO contrast
C2826012|T102|strict|35925-7|LNC|Fluoroscopy Guidance for endoscopy of Stomach|Fluoroscopy Guidance for endoscopy of Stomach
C2826012|T102|strict|43478-7|LNC|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 1.5 hours post contrast retrograde|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 1.5 hours post contrast retrograde
C2826012|T102|strict|43474-6|LNC|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 15 minutes post contrast retrograde|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 15 minutes post contrast retrograde
C2826012|T102|strict|43477-9|LNC|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 1 hour post contrast retrograde|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 1 hour post contrast retrograde
C2826012|T102|strict|43473-8|LNC|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 2 hours post contrast retrograde|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 2 hours post contrast retrograde
C2826012|T102|strict|43475-3|LNC|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 30 minutes post contrast retrograde|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 30 minutes post contrast retrograde
C2826012|T102|strict|43476-1|LNC|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 45 minutes post contrast retrograde|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 45 minutes post contrast retrograde
C2826012|T102|strict|72248-8|LNC|Abdomen MRCP with and without contrast IV|Abdomen MRCP with and without contrast IV
C2826012|T102|strict|44214-5|LNC|Fluoroscopy Guidance for endoscopy of Biliary ducts-- W contrast retrograde|Fluoroscopy Guidance for endoscopy of Biliary ducts-- W contrast retrograde
C2826012|T102|strict|30815-5|LNC|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- W contrast retrograde|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- W contrast retrograde
C2826012|T102|strict|44213-7|LNC|Fluoroscopy Guidance for endoscopy of Pancreatic duct-- W contrast retrograde|Fluoroscopy Guidance for endoscopy of Pancreatic duct-- W contrast retrograde
C2826012|T102|strict|58740-2|LNC|Abdomen MRCP WO contrast|Abdomen MRCP WO contrast
C2826012|T102|strict|72541-6|LNC|Fluoroscopy Guidance for facet joint denervation of Spine Cervical|Fluoroscopy Guidance for facet joint denervation of Spine Cervical
C2826012|T102|strict|72542-4|LNC|Fluoroscopy Guidance for facet joint denervation of Spine Lumbar|Fluoroscopy Guidance for facet joint denervation of Spine Lumbar
C2826012|T102|strict|72540-8|LNC|Fluoroscopy Guidance for facet joint denervation of Spine|Fluoroscopy Guidance for facet joint denervation of Spine
C2826012|T102|strict|35926-5|LNC|Fluoroscopy Guidance for gastrostomy of Stomach|Fluoroscopy Guidance for gastrostomy of Stomach
C2826012|T102|strict|30638-1|LNC|Fluoroscopy Guidance for injection of Hip|Fluoroscopy Guidance for injection of Hip
C2826012|T102|strict|24769-2|LNC|CT Guidance for injection of Joint space|CT Guidance for injection of Joint space
C2826012|T102|strict|42334-3|LNC|Fluoroscopy Guidance for injection of Mammary artery.internal - left|Fluoroscopy Guidance for injection of Mammary artery.internal - left
C2826012|T102|strict|42706-2|LNC|US Guidance for injection of Pleural space|US Guidance for injection of Pleural space
C2826012|T102|strict|24901-1|LNC|CT Guidance for injection of Sacroiliac Joint|CT Guidance for injection of Sacroiliac Joint
C2826012|T102|strict|35927-3|LNC|Fluoroscopy Guidance for injection of Sacroiliac Joint|Fluoroscopy Guidance for injection of Sacroiliac Joint
C2826012|T102|strict|26319-4|LNC|CT Guidance for injection of Sacroiliac joint - bilateral|CT Guidance for injection of Sacroiliac joint - bilateral
C2826012|T102|strict|26320-2|LNC|CT Guidance for injection of Sacroiliac joint - left|CT Guidance for injection of Sacroiliac joint - left
C2826012|T102|strict|26321-0|LNC|CT Guidance for injection of Sacroiliac joint - right|CT Guidance for injection of Sacroiliac joint - right
C2826012|T102|strict|48435-2|LNC|Fluoroscopy Guidance for injection of Salivary gland - bilateral|Fluoroscopy Guidance for injection of Salivary gland - bilateral
C2826012|T102|strict|46392-7|LNC|Fluoroscopy Guidance for injection of Sinuses|Fluoroscopy Guidance for injection of Sinuses
C2826012|T102|strict|37427-2|LNC|Fluoroscopy Guidance for injection of Spine|Fluoroscopy Guidance for injection of Spine
C2826012|T102|strict|30579-7|LNC|CT Guidance for injection of Spine facet joint|CT Guidance for injection of Spine facet joint
C2826012|T102|strict|24931-8|LNC|Fluoroscopy Guidance for injection of Spine facet joint|Fluoroscopy Guidance for injection of Spine facet joint
C2826012|T102|strict|26322-8|LNC|Fluoroscopy Guidance for injection of Spine facet joint - bilateral|Fluoroscopy Guidance for injection of Spine facet joint - bilateral
C2826012|T102|strict|26323-6|LNC|Fluoroscopy Guidance for injection of Spine facet joint - left|Fluoroscopy Guidance for injection of Spine facet joint - left
C2826012|T102|strict|26324-4|LNC|Fluoroscopy Guidance for injection of Spine facet joint - right|Fluoroscopy Guidance for injection of Spine facet joint - right
C2826012|T102|strict|70918-8|LNC|Fluoroscopy Guidance for injection of Spine Cervical|Fluoroscopy Guidance for injection of Spine Cervical
C2826012|T102|strict|30812-2|LNC|Fluoroscopy Guidance for injection of Spine Cervical Facet Joint|Fluoroscopy Guidance for injection of Spine Cervical Facet Joint
C2826012|T102|strict|37493-4|LNC|CT Guidance for injection of Spine.disc.cervical|CT Guidance for injection of Spine.disc.cervical
C2826012|T102|strict|70919-6|LNC|Fluoroscopy Guidance for injection of Spine Lumbar|Fluoroscopy Guidance for injection of Spine Lumbar
C2826012|T102|strict|30817-1|LNC|Fluoroscopy Guidance for injection of Spine Lumbar Facet Joint|Fluoroscopy Guidance for injection of Spine Lumbar Facet Joint
C2826012|T102|strict|70920-4|LNC|Fluoroscopy Guidance for injection of Spine Thoracic|Fluoroscopy Guidance for injection of Spine Thoracic
C2826012|T102|strict|30814-8|LNC|Fluoroscopy Guidance for injection of Spine Thoracic Facet Joint|Fluoroscopy Guidance for injection of Spine Thoracic Facet Joint
C2826012|T102|strict|30702-5|LNC|US Guidance for injection of Thyroid|US Guidance for injection of Thyroid
C2826012|T102|strict|72530-9|LNC|US Guidance for injection of Joint|US Guidance for injection of Joint
C2826012|T102|strict|36771-4|LNC|Fluoroscopy Guidance for injection of Joint|Fluoroscopy Guidance for injection of Joint
C2826012|T102|strict|37494-2|LNC|Fluoroscopy Guidance for injection of Tendon|Fluoroscopy Guidance for injection of Tendon
C2826012|T102|strict|72537-4|LNC|US Guidance for injection of sclerosing agent of Extremity vein - bilateral|US Guidance for injection of sclerosing agent of Extremity vein - bilateral
C2826012|T102|strict|72645-5|LNC|US Guidance for injection of sclerosing agent of Extremity vein - left|US Guidance for injection of sclerosing agent of Extremity vein - left
C2826012|T102|strict|72644-8|LNC|US Guidance for injection of sclerosing agent of Extremity vein - right|US Guidance for injection of sclerosing agent of Extremity vein - right
C2826012|T102|strict|72536-6|LNC|US Guidance for injection of sclerosing agent of Extremity veins - bilateral|US Guidance for injection of sclerosing agent of Extremity veins - bilateral
C2826012|T102|strict|72643-0|LNC|US Guidance for injection of sclerosing agent of Extremity veins - left|US Guidance for injection of sclerosing agent of Extremity veins - left
C2826012|T102|strict|72642-2|LNC|US Guidance for injection of sclerosing agent of Extremity veins - right|US Guidance for injection of sclerosing agent of Extremity veins - right
C2826012|T102|strict|72543-2|LNC|Fluoroscopy Guidance for intercostal nerve devervation of Spine Thoracic|Fluoroscopy Guidance for intercostal nerve devervation of Spine Thoracic
C2826012|T102|strict|72552-3|LNC|Fluoroscopy Guidance for kyphoplasty of Spine Lumbar|Fluoroscopy Guidance for kyphoplasty of Spine Lumbar
C2826012|T102|strict|72553-1|LNC|Fluoroscopy Guidance for kyphoplasty of Spine Thoracic|Fluoroscopy Guidance for kyphoplasty of Spine Thoracic
C2826012|T102|strict|72535-8|LNC|US Guidance for laser ablation of vein(s) of Extremity vein - left|US Guidance for laser ablation of vein(s) of Extremity vein - left
C2826012|T102|strict|72534-1|LNC|US Guidance for laser ablation of vein(s) of Extremity vein - right|US Guidance for laser ablation of vein(s) of Extremity vein - right
C2826012|T102|strict|48735-5|LNC|Mammogram Guidance for localization of Breast|Mammogram Guidance for localization of Breast
C2826012|T102|strict|43759-0|LNC|US Guidance for localization of Breast - bilateral|US Guidance for localization of Breast - bilateral
C2826012|T102|strict|35928-1|LNC|CT Guidance for localization of Breast - left|CT Guidance for localization of Breast - left
C2826012|T102|strict|42296-4|LNC|Mammogram Guidance for localization of Breast - left|Mammogram Guidance for localization of Breast - left
C2826012|T102|strict|43758-2|LNC|US Guidance for localization of Breast - left|US Guidance for localization of Breast - left
C2826012|T102|strict|35929-9|LNC|CT Guidance for localization of Breast - right|CT Guidance for localization of Breast - right
C2826012|T102|strict|42297-2|LNC|Mammogram Guidance for localization of Breast - right|Mammogram Guidance for localization of Breast - right
C2826012|T102|strict|43760-8|LNC|US Guidance for localization of Breast - right|US Guidance for localization of Breast - right
C2826012|T102|strict|37608-7|LNC|US Guidance for localization of foreign body of Eye|US Guidance for localization of foreign body of Eye
C2826012|T102|strict|42701-3|LNC|CT Guidance for localization of placenta of Uterus|CT Guidance for localization of placenta of Uterus
C2826012|T102|strict|39760-4|LNC|Scan Guidance for localization of tumor limited|Scan Guidance for localization of tumor limited
C2826012|T102|strict|39759-6|LNC|SPECT Guidance for localization of tumor limited|SPECT Guidance for localization of tumor limited
C2826012|T102|strict|39761-2|LNC|Scan Guidance for localization of tumor limited-- W Tc-99m Sestamibi IV|Scan Guidance for localization of tumor limited-- W Tc-99m Sestamibi IV
C2826012|T102|strict|39953-5|LNC|Scan Guidance for localization of tumor multiple areas|Scan Guidance for localization of tumor multiple areas
C2826012|T102|strict|39763-8|LNC|Scan Guidance for localization of tumor|Scan Guidance for localization of tumor
C2826012|T102|strict|39762-0|LNC|SPECT Guidance for localization of tumor|SPECT Guidance for localization of tumor
C2826012|T102|strict|39758-8|LNC|Scan Guidance for localization of tumor of Breast|Scan Guidance for localization of tumor of Breast
C2826012|T102|strict|44110-5|LNC|CT Guidance for needle localization of Breast|CT Guidance for needle localization of Breast
C2826012|T102|strict|24600-9|LNC|US Guidance for needle localization of Breast|US Guidance for needle localization of Breast
C2826012|T102|strict|69068-5|LNC|Mammogram Guidance for needle localization of Breast - bilateral|Mammogram Guidance for needle localization of Breast - bilateral
C2826012|T102|strict|26313-7|LNC|US Guidance for needle localization of Breast - bilateral|US Guidance for needle localization of Breast - bilateral
C2826012|T102|strict|26314-5|LNC|US Guidance for needle localization of Breast - left|US Guidance for needle localization of Breast - left
C2826012|T102|strict|26318-6|LNC|US Guidance for needle localization of Breast - right|US Guidance for needle localization of Breast - right
C2826012|T102|strict|37921-4|LNC|US Guidance for needle localization of Chest|US Guidance for needle localization of Chest
C2826012|T102|strict|42021-6|LNC|CT Guidance for needle localization of Spine Cervical|CT Guidance for needle localization of Spine Cervical
C2826012|T102|strict|42020-8|LNC|CT Guidance for needle localization of Spine Lumbar|CT Guidance for needle localization of Spine Lumbar
C2826012|T102|strict|39026-0|LNC|CT Guidance for needle localization of Unspecified body region|CT Guidance for needle localization of Unspecified body region
C2826012|T102|strict|39028-6|LNC|MRI Guidance for needle localization of Unspecified body region|MRI Guidance for needle localization of Unspecified body region
C2826012|T102|strict|38032-9|LNC|US Guidance for needle localization of Unspecified body region|US Guidance for needle localization of Unspecified body region
C2826012|T102|strict|39027-8|LNC|Fluoroscopy Guidance for needle localization of Unspecified body region|Fluoroscopy Guidance for needle localization of Unspecified body region
C2826012|T102|strict|24595-1|LNC|Mammogram Guidance for needle localization of mass of Breast|Mammogram Guidance for needle localization of mass of Breast
C2826012|T102|strict|26315-2|LNC|Mammogram Guidance for needle localization of mass of Breast - bilateral|Mammogram Guidance for needle localization of mass of Breast - bilateral
C2826012|T102|strict|26316-0|LNC|Mammogram Guidance for needle localization of mass of Breast - left|Mammogram Guidance for needle localization of mass of Breast - left
C2826012|T102|strict|26317-8|LNC|Mammogram Guidance for needle localization of mass of Breast - right|Mammogram Guidance for needle localization of mass of Breast - right
C2826012|T102|strict|44118-8|LNC|CT Guidance for needle localization of Breast-- W and WO contrast IV|CT Guidance for needle localization of Breast-- W and WO contrast IV
C2826012|T102|strict|35930-7|LNC|CT Guidance for nerve block of Abdomen|CT Guidance for nerve block of Abdomen
C2826012|T102|strict|35931-5|LNC|CT Guidance for nerve block of Pelvis|CT Guidance for nerve block of Pelvis
C2826012|T102|strict|70921-2|LNC|CT Guidance for nerve block of Spine Cervical|CT Guidance for nerve block of Spine Cervical
C2826012|T102|strict|35932-3|LNC|CT Guidance for nerve block of Spine Lumbar|CT Guidance for nerve block of Spine Lumbar
C2826012|T102|strict|70922-0|LNC|CT Guidance for nerve block of Spine Thoracic|CT Guidance for nerve block of Spine Thoracic
C2826012|T102|strict|69240-0|LNC|Fluoroscopy Guidance for percutaneous biopsy of Abdomen|Fluoroscopy Guidance for percutaneous biopsy of Abdomen
C2826012|T102|strict|42139-6|LNC|US Guidance for percutaneous biopsy of Muscle|US Guidance for percutaneous biopsy of Muscle
C2826012|T102|strict|24609-0|LNC|Mammogram Guidance for core needle percutaneous biopsy of Breast|Mammogram Guidance for core needle percutaneous biopsy of Breast
C2826012|T102|strict|26334-3|LNC|Mammogram Guidance for core needle percutaneous biopsy of Breast - bilateral|Mammogram Guidance for core needle percutaneous biopsy of Breast - bilateral
C2826012|T102|strict|26335-0|LNC|Mammogram Guidance for core needle percutaneous biopsy of Breast - left|Mammogram Guidance for core needle percutaneous biopsy of Breast - left
C2826012|T102|strict|38023-8|LNC|US Guidance for core needle percutaneous biopsy of Breast - left|US Guidance for core needle percutaneous biopsy of Breast - left
C2826012|T102|strict|26336-8|LNC|Mammogram Guidance for core needle percutaneous biopsy of Breast - right|Mammogram Guidance for core needle percutaneous biopsy of Breast - right
C2826012|T102|strict|38025-3|LNC|US Guidance for core needle percutaneous biopsy of Breast - right|US Guidance for core needle percutaneous biopsy of Breast - right
C2826012|T102|strict|44121-2|LNC|Mammogram Guidance for percutaneous needle biopsy of Breast|Mammogram Guidance for percutaneous needle biopsy of Breast
C2826012|T102|strict|69245-9|LNC|Fluoroscopy Guidance for percutaneous needle biopsy of Kidney|Fluoroscopy Guidance for percutaneous needle biopsy of Kidney
C2826012|T102|strict|69246-7|LNC|Fluoroscopy Guidance for percutaneous needle biopsy of Liver|Fluoroscopy Guidance for percutaneous needle biopsy of Liver
C2826012|T102|strict|44204-6|LNC|Fluoroscopy Guidance for percutaneous needle biopsy of Lung|Fluoroscopy Guidance for percutaneous needle biopsy of Lung
C2826012|T102|strict|69247-5|LNC|Fluoroscopy Guidance for percutaneous needle biopsy of Salivary gland|Fluoroscopy Guidance for percutaneous needle biopsy of Salivary gland
C2826012|T102|strict|46372-9|LNC|Fluoroscopy Guidance for percutaneous drainage of Biliary ducts|Fluoroscopy Guidance for percutaneous drainage of Biliary ducts
C2826012|T102|strict|62494-0|LNC|US Guidance for percutaneous drainage of Cavity|US Guidance for percutaneous drainage of Cavity
C2826012|T102|strict|24621-5|LNC|Fluoroscopy Guidance for percutaneous drainage of Cavity|Fluoroscopy Guidance for percutaneous drainage of Cavity
C2826012|T102|strict|69241-8|LNC|Fluoroscopy Guidance for percutaneous drainage of abscess of Abdomen|Fluoroscopy Guidance for percutaneous drainage of abscess of Abdomen
C2826012|T102|strict|69242-6|LNC|Fluoroscopy Guidance for percutaneous drainage of abscess of Appendix|Fluoroscopy Guidance for percutaneous drainage of abscess of Appendix
C2826012|T102|strict|42422-6|LNC|Fluoroscopy Guidance for percutaneous drainage of abscess of Breast|Fluoroscopy Guidance for percutaneous drainage of abscess of Breast
C2826012|T102|strict|43444-9|LNC|CT Guidance for percutaneous drainage of abscess of Cavity|CT Guidance for percutaneous drainage of abscess of Cavity
C2826012|T102|strict|42423-4|LNC|Fluoroscopy Guidance for percutaneous drainage of abscess of Chest|Fluoroscopy Guidance for percutaneous drainage of abscess of Chest
C2826012|T102|strict|69243-4|LNC|Fluoroscopy Guidance for percutaneous drainage of abscess of Lung|Fluoroscopy Guidance for percutaneous drainage of abscess of Lung
C2826012|T102|strict|44223-6|LNC|Fluoroscopy Guidance for percutaneous drainage of abscess of Ovary|Fluoroscopy Guidance for percutaneous drainage of abscess of Ovary
C2826012|T102|strict|69244-2|LNC|Fluoroscopy Guidance for percutaneous drainage of abscess of Pelvis|Fluoroscopy Guidance for percutaneous drainage of abscess of Pelvis
C2826012|T102|strict|42421-8|LNC|Fluoroscopy Guidance for percutaneous drainage of abscess of Unspecified body region|Fluoroscopy Guidance for percutaneous drainage of abscess of Unspecified body region
C2826012|T102|strict|35933-1|LNC|CT Guidance for percutaneous vertebroplasty of Spine|CT Guidance for percutaneous vertebroplasty of Spine
C2826012|T102|strict|35936-4|LNC|Fluoroscopy Guidance for percutaneous vertebroplasty of Spine|Fluoroscopy Guidance for percutaneous vertebroplasty of Spine
C2826012|T102|strict|70923-8|LNC|Fluoroscopy Guidance for percutaneous vertebroplasty of Spine Cervical|Fluoroscopy Guidance for percutaneous vertebroplasty of Spine Cervical
C2826012|T102|strict|35934-9|LNC|CT Guidance for percutaneous vertebroplasty of Spine Lumbar|CT Guidance for percutaneous vertebroplasty of Spine Lumbar
C2826012|T102|strict|70924-6|LNC|Fluoroscopy Guidance for percutaneous vertebroplasty of Spine Lumbar|Fluoroscopy Guidance for percutaneous vertebroplasty of Spine Lumbar
C2826012|T102|strict|35935-6|LNC|CT Guidance for percutaneous vertebroplasty of Spine Thoracic|CT Guidance for percutaneous vertebroplasty of Spine Thoracic
C2826012|T102|strict|70925-3|LNC|Fluoroscopy Guidance for percutaneous vertebroplasty of Spine Thoracic|Fluoroscopy Guidance for percutaneous vertebroplasty of Spine Thoracic
C2826012|T102|strict|72539-0|LNC|Fluoroscopy Guidance for peripheral nerve denervation of Unspecified body region|Fluoroscopy Guidance for peripheral nerve denervation of Unspecified body region
C2826012|T102|strict|30643-1|LNC|US Guidance for placement of catheter in Central vein|US Guidance for placement of catheter in Central vein
C2826012|T102|strict|35912-5|LNC|Fluoroscopy Guidance for placement of catheter in Unspecified body region|Fluoroscopy Guidance for placement of catheter in Unspecified body region
C2826012|T102|strict|25028-2|LNC|Fluoroscopic angiogram Guidance for placement of catheter for adminstration of thrombolytic in Vessel|Fluoroscopic angiogram Guidance for placement of catheter for adminstration of thrombolytic in Vessel
C2826012|T102|strict|25029-0|LNC|Fluoroscopic angiogram Guidance for placement of catheter for vasoconstrictor infusion in Vessels|Fluoroscopic angiogram Guidance for placement of catheter for vasoconstrictor infusion in Vessels
C2826012|T102|strict|24613-2|LNC|Fluoroscopic angiogram Guidance for placement of catheter in artery in Central cardiovascular artery|Fluoroscopic angiogram Guidance for placement of catheter in artery in Central cardiovascular artery
C2826012|T102|strict|30644-9|LNC|US Guidance for placement of catheter in Central vein-- Tunneled|US Guidance for placement of catheter in Central vein-- Tunneled
C2826012|T102|strict|25077-9|LNC|Fluoroscopic angiogram Guidance for placement of catheter in Hepatic artery-- W contrast IA|Fluoroscopic angiogram Guidance for placement of catheter in Hepatic artery-- W contrast IA
C2826012|T102|strict|24625-6|LNC|Fluoroscopic angiogram Guidance for placement of catheter in Central vein-- W contrast IV|Fluoroscopic angiogram Guidance for placement of catheter in Central vein-- W contrast IV
C2826012|T102|strict|26310-3|LNC|Fluoroscopic angiogram Guidance for placement of catheter in Central vein - bilateral-- W contrast IV|Fluoroscopic angiogram Guidance for placement of catheter in Central vein - bilateral-- W contrast IV
C2826012|T102|strict|26311-1|LNC|Fluoroscopic angiogram Guidance for placement of catheter in Central vein - left-- W contrast IV|Fluoroscopic angiogram Guidance for placement of catheter in Central vein - left-- W contrast IV
C2826012|T102|strict|26312-9|LNC|Fluoroscopic angiogram Guidance for placement of catheter in Central vein - right-- W contrast IV|Fluoroscopic angiogram Guidance for placement of catheter in Central vein - right-- W contrast IV
C2826012|T102|strict|41801-2|LNC|Fluoroscopic angiogram Guidance for placement of catheter in Portal vein-- W contrast IV|Fluoroscopic angiogram Guidance for placement of catheter in Portal vein-- W contrast IV
C2826012|T102|strict|24716-3|LNC|Fluoroscopy Guidance for placement of decompression tube in Gastrointestine|Fluoroscopy Guidance for placement of decompression tube in Gastrointestine
C2826012|T102|strict|62491-6|LNC|Fluoroscopic angiogram Guidance for placement of ilio-iliac tube endoprosthesis in Iliac artery - left-- W contrast IA|Fluoroscopic angiogram Guidance for placement of ilio-iliac tube endoprosthesis in Iliac artery - left-- W contrast IA
C2826012|T102|strict|62492-4|LNC|Fluoroscopic angiogram Guidance for placement of ilio-iliac tube endoprosthesis in Iliac artery - right-- W contrast IA|Fluoroscopic angiogram Guidance for placement of ilio-iliac tube endoprosthesis in Iliac artery - right-- W contrast IA
C2826012|T102|strict|25072-0|LNC|Guidance for placement of infusion port in Unspecified body region|Guidance for placement of infusion port in Unspecified body region
C2826012|T102|strict|62450-2|LNC|Fluoroscopic angiogram Guidance for placement of intraperitoneal catheter in Abdomen|Fluoroscopic angiogram Guidance for placement of intraperitoneal catheter in Abdomen
C2826012|T102|strict|25026-6|LNC|Fluoroscopic angiogram Guidance for placement of IVC filter in Inferior vena cava-- W contrast IV|Fluoroscopic angiogram Guidance for placement of IVC filter in Inferior vena cava-- W contrast IV
C2826012|T102|strict|25027-4|LNC|Guidance for placement of large bore catheter into vessel in Central vein|Guidance for placement of large bore catheter into vessel in Central vein
C2826012|T102|strict|26307-9|LNC|Guidance for placement of large bore catheter into vessel in Central vein - bilateral|Guidance for placement of large bore catheter into vessel in Central vein - bilateral
C2826012|T102|strict|26308-7|LNC|Guidance for placement of large bore catheter into vessel in Central vein - left|Guidance for placement of large bore catheter into vessel in Central vein - left
C2826012|T102|strict|26309-5|LNC|Guidance for placement of large bore catheter into vessel in Central vein - right|Guidance for placement of large bore catheter into vessel in Central vein - right
C2826012|T102|strict|25024-1|LNC|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein
C2826012|T102|strict|26304-6|LNC|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein - bilateral|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein - bilateral
C2826012|T102|strict|26305-3|LNC|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein - left|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein - left
C2826012|T102|strict|26306-1|LNC|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein - right|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein - right
C2826012|T102|strict|64993-9|LNC|US Guidance for placement of needle in Unspecified body region|US Guidance for placement of needle in Unspecified body region
C2826012|T102|strict|42456-4|LNC|US Guidance for placement of needle wire in Breast|US Guidance for placement of needle wire in Breast
C2826012|T102|strict|36772-2|LNC|CT Guidance for placement of nephrostomy tube in Kidney|CT Guidance for placement of nephrostomy tube in Kidney
C2826012|T102|strict|24779-1|LNC|Fluoroscopy Guidance for placement of percutaneous nephrostomy in Kidney - bilateral-- W contrast via tube|Fluoroscopy Guidance for placement of percutaneous nephrostomy in Kidney - bilateral-- W contrast via tube
C2826012|T102|strict|24782-5|LNC|Fluoroscopy Guidance for placement of percutaneous nephroureteral stent in Kidney - bilateral|Fluoroscopy Guidance for placement of percutaneous nephroureteral stent in Kidney - bilateral
C2826012|T102|strict|35937-2|LNC|CT Guidance for placement of radiation therapy fields in Unspecified body region|CT Guidance for placement of radiation therapy fields in Unspecified body region
C2826012|T102|strict|43487-8|LNC|US Guidance for placement of radiation therapy fields in Unspecified body region|US Guidance for placement of radiation therapy fields in Unspecified body region
C2826012|T102|strict|65797-3|LNC|Fluoroscopic angiogram Guidance for placement of stent in Artery - left|Fluoroscopic angiogram Guidance for placement of stent in Artery - left
C2826012|T102|strict|65798-1|LNC|Fluoroscopic angiogram Guidance for placement of stent in Artery - right|Fluoroscopic angiogram Guidance for placement of stent in Artery - right
C2826012|T102|strict|69134-5|LNC|Fluoroscopic angiogram Guidance for placement of stent in Iliac artery|Fluoroscopic angiogram Guidance for placement of stent in Iliac artery
C2826012|T102|strict|25078-7|LNC|Fluoroscopy Guidance for placement of stent in Intrahepatic portal system|Fluoroscopy Guidance for placement of stent in Intrahepatic portal system
C2826012|T102|strict|24756-9|LNC|Fluoroscopic angiogram Guidance for placement of stent in Vein|Fluoroscopic angiogram Guidance for placement of stent in Vein
C2826012|T102|strict|26301-2|LNC|Fluoroscopic angiogram Guidance for placement of stent in Vein - bilateral|Fluoroscopic angiogram Guidance for placement of stent in Vein - bilateral
C2826012|T102|strict|26302-0|LNC|Fluoroscopic angiogram Guidance for placement of stent in Vein - left|Fluoroscopic angiogram Guidance for placement of stent in Vein - left
C2826012|T102|strict|26303-8|LNC|Fluoroscopic angiogram Guidance for placement of stent in Vein - right|Fluoroscopic angiogram Guidance for placement of stent in Vein - right
C2826012|T102|strict|24555-5|LNC|Fluoroscopic angiogram Guidance for placement of stent in Artery|Fluoroscopic angiogram Guidance for placement of stent in Artery
C2826012|T102|strict|51391-1|LNC|Fluoroscopic angiogram Guidance for placement of transjugular intrahepatic portosystemic shunt in Portal vein and Hepatic vein|Fluoroscopic angiogram Guidance for placement of transjugular intrahepatic portosystemic shunt in Portal vein and Hepatic vein
C2826012|T102|strict|35938-0|LNC|CT Guidance for placement of tube in Chest|CT Guidance for placement of tube in Chest
C2826012|T102|strict|42140-4|LNC|US Guidance for placement of tube in Chest|US Guidance for placement of tube in Chest
C2826012|T102|strict|39362-9|LNC|Fluoroscopy Guidance for placement of tube in Chest|Fluoroscopy Guidance for placement of tube in Chest
C2826012|T102|strict|30637-3|LNC|Fluoroscopy Guidance for placement of tube in Gastrointestine|Fluoroscopy Guidance for placement of tube in Gastrointestine
C2826012|T102|strict|41799-8|LNC|Fluoroscopy Guidance for placement of tube in Liver|Fluoroscopy Guidance for placement of tube in Liver
C2826012|T102|strict|24995-3|LNC|Fluoroscopy Guidance for placement of tube in Stomach|Fluoroscopy Guidance for placement of tube in Stomach
C2826012|T102|strict|44224-4|LNC|Fluoroscopy Guidance for placement of tube in Unspecified body region|Fluoroscopy Guidance for placement of tube in Unspecified body region
C2826012|T102|strict|46373-7|LNC|SPECT Guidance for placement of tube in Chest|SPECT Guidance for placement of tube in Chest
C2826012|T102|strict|44102-2|LNC|CT Guidance for procedure of Joint space|CT Guidance for procedure of Joint space
C2826012|T102|strict|44222-8|LNC|Fluoroscopy Guidance for procedure of Joint space|Fluoroscopy Guidance for procedure of Joint space
C2826012|T102|strict|30629-0|LNC|Fluoroscopy Guidance for procedure of Unspecified body region|Fluoroscopy Guidance for procedure of Unspecified body region
C2826012|T102|strict|30581-3|LNC|CT Guidance for radiation treatment of Unspecified body region-- W contrast IV|CT Guidance for radiation treatment of Unspecified body region-- W contrast IV
C2826012|T102|strict|30664-7|LNC|MRI Guidance for radiation treatment of Unspecified body region-- W contrast IV|MRI Guidance for radiation treatment of Unspecified body region-- W contrast IV
C2826012|T102|strict|30582-1|LNC|CT Guidance for radiation treatment of Unspecified body region-- WO contrast|CT Guidance for radiation treatment of Unspecified body region-- WO contrast
C2826012|T102|strict|30665-4|LNC|MRI Guidance for radiation treatment of Unspecified body region-- WO contrast|MRI Guidance for radiation treatment of Unspecified body region-- WO contrast
C2826012|T102|strict|25053-0|LNC|CT Guidance for radiosurgery of Unspecified body region|CT Guidance for radiosurgery of Unspecified body region
C2826012|T102|strict|25054-8|LNC|CT Guidance for radiosurgery of Unspecified body region-- W contrast IV|CT Guidance for radiosurgery of Unspecified body region-- W contrast IV
C2826012|T102|strict|24537-3|LNC|US Guidance for removal of amniotic fluid from Uterus|US Guidance for removal of amniotic fluid from Uterus
C2826012|T102|strict|42141-2|LNC|US Guidance for removal of catheter from Central vein-- Tunneled|US Guidance for removal of catheter from Central vein-- Tunneled
C2826012|T102|strict|72549-9|LNC|Fluoroscopy Guidance for removal of catheter from Central vein-- Tunneled|Fluoroscopy Guidance for removal of catheter from Central vein-- Tunneled
C2826012|T102|strict|72548-1|LNC|Fluoroscopic angiogram Guidance for removal of catheter from Central vein-- W contrast IV|Fluoroscopic angiogram Guidance for removal of catheter from Central vein-- W contrast IV
C2826012|T102|strict|72547-3|LNC|Fluoroscopy Guidance for removal of CVA device obstruction from Central vein|Fluoroscopy Guidance for removal of CVA device obstruction from Central vein
C2826012|T102|strict|72546-5|LNC|Fluoroscopy Guidance for removal of CVA lumen obstruction from Central vein|Fluoroscopy Guidance for removal of CVA lumen obstruction from Central vein
C2826012|T102|strict|41810-3|LNC|CT Guidance for removal of fluid from Abdomen|CT Guidance for removal of fluid from Abdomen
C2826012|T102|strict|24559-7|LNC|US Guidance for removal of fluid from Abdomen|US Guidance for removal of fluid from Abdomen
C2826012|T102|strict|38142-6|LNC|US Guidance for removal of fluid from Chest|US Guidance for removal of fluid from Chest
C2826012|T102|strict|30628-2|LNC|Fluoroscopy Guidance for removal of foreign body from Unspecified body region|Fluoroscopy Guidance for removal of foreign body from Unspecified body region
C2826012|T102|strict|72538-2|LNC|Fluoroscopic angiogram Guidance for removal of longterm peripheral catheter from Central vein|Fluoroscopic angiogram Guidance for removal of longterm peripheral catheter from Central vein
C2826012|T102|strict|72544-0|LNC|Fluoroscopy Guidance for removal of percutaneous nephrostomy tube from Kidney - bilateral-- W contrast|Fluoroscopy Guidance for removal of percutaneous nephrostomy tube from Kidney - bilateral-- W contrast
C2826012|T102|strict|24885-6|LNC|US Guidance for repair of Pseudoaneurysm/AV fistula|US Guidance for repair of Pseudoaneurysm/AV fistula
C2826012|T102|strict|72550-7|LNC|Fluoroscopy Guidance for repair of CVA catheter with port or pump of Central vein|Fluoroscopy Guidance for repair of CVA catheter with port or pump of Central vein
C2826012|T102|strict|72551-5|LNC|Fluoroscopy Guidance for repair of CVA catheter without port or pump of Central vein|Fluoroscopy Guidance for repair of CVA catheter without port or pump of Central vein
C2826012|T102|strict|42017-4|LNC|Fluoroscopy Guidance for replacement of percutaneous cholecystostomy in Abdomen|Fluoroscopy Guidance for replacement of percutaneous cholecystostomy in Abdomen
C2826012|T102|strict|52790-3|LNC|CT Guidance for replacement of percutaneous drainage tube in Abdomen|CT Guidance for replacement of percutaneous drainage tube in Abdomen
C2826012|T102|strict|72545-7|LNC|Fluoroscopy Guidance for replacement of percutaneous drainage tube in Biliary ducts and Gallbladder|Fluoroscopy Guidance for replacement of percutaneous drainage tube in Biliary ducts and Gallbladder
C2826012|T102|strict|52791-1|LNC|CT Guidance for replacement of percutaneous drainage tube in Pelvis|CT Guidance for replacement of percutaneous drainage tube in Pelvis
C2826012|T102|strict|46294-5|LNC|Fluoroscopy Guidance for replacement of percutaneous drainage tube in Stomach|Fluoroscopy Guidance for replacement of percutaneous drainage tube in Stomach
C2826012|T102|strict|24996-1|LNC|Fluoroscopy Guidance for replacement of percutaneous gastrostomy in Stomach|Fluoroscopy Guidance for replacement of percutaneous gastrostomy in Stomach
C2826012|T102|strict|24626-4|LNC|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein-- W contrast IV|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein-- W contrast IV
C2826012|T102|strict|26295-6|LNC|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein - bilateral-- W contrast IV|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein - bilateral-- W contrast IV
C2826012|T102|strict|26296-4|LNC|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein - left-- W contrast IV|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein - left-- W contrast IV
C2826012|T102|strict|26297-2|LNC|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein - right-- W contrast IV|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein - right-- W contrast IV
C2826012|T102|strict|48740-5|LNC|Mammogram Guidance for sentinel lymph node injection of Breast|Mammogram Guidance for sentinel lymph node injection of Breast
C2826012|T102|strict|48736-3|LNC|Mammogram Guidance for sentinel lymph node injection of Breast - left|Mammogram Guidance for sentinel lymph node injection of Breast - left
C2826012|T102|strict|48739-7|LNC|Mammogram Guidance for sentinel lymph node injection of Breast - right|Mammogram Guidance for sentinel lymph node injection of Breast - right
C2826012|T102|strict|24570-4|LNC|Fluoroscopy Guidance for stone removal of Biliary duct common-- W contrast intra biliary duct|Fluoroscopy Guidance for stone removal of Biliary duct common-- W contrast intra biliary duct
C2826012|T102|strict|43763-2|LNC|Fluoroscopic angiogram Guidance for thrombectomy of Vein-- W contrast IV|Fluoroscopic angiogram Guidance for thrombectomy of Vein-- W contrast IV
C2826012|T102|strict|43761-6|LNC|Fluoroscopic angiogram Guidance for thrombectomy of Vein - bilateral-- W contrast IV|Fluoroscopic angiogram Guidance for thrombectomy of Vein - bilateral-- W contrast IV
C2826012|T102|strict|43762-4|LNC|Fluoroscopic angiogram Guidance for thrombectomy of Vein - left-- W contrast IV|Fluoroscopic angiogram Guidance for thrombectomy of Vein - left-- W contrast IV
C2826012|T102|strict|43764-0|LNC|Fluoroscopic angiogram Guidance for thrombectomy of Vein - right-- W contrast IV|Fluoroscopic angiogram Guidance for thrombectomy of Vein - right-- W contrast IV
C2826012|T102|strict|72554-9|LNC|Fluoroscopy Guidance for trigger point injection of Muscle|Fluoroscopy Guidance for trigger point injection of Muscle
C2826012|T102|strict|39138-3|LNC|Fluoroscopic angiogram Guidance for vascular access of Vessel|Fluoroscopic angiogram Guidance for vascular access of Vessel
C2826012|T102|strict|39139-1|LNC|US Guidance for vascular access of Unspecified body region|US Guidance for vascular access of Unspecified body region
C2826012|T102|strict|36936-3|LNC|MRI Guidance.stereotactic for biopsy of Brain|MRI Guidance.stereotactic for biopsy of Brain
C2826012|T102|strict|24603-3|LNC|Mammogram Guidance.stereotactic for biopsy of Breast|Mammogram Guidance.stereotactic for biopsy of Breast
C2826012|T102|strict|26292-3|LNC|Mammogram Guidance.stereotactic for biopsy of Breast - bilateral|Mammogram Guidance.stereotactic for biopsy of Breast - bilateral
C2826012|T102|strict|26293-1|LNC|Mammogram Guidance.stereotactic for biopsy of Breast - left|Mammogram Guidance.stereotactic for biopsy of Breast - left
C2826012|T102|strict|26294-9|LNC|Mammogram Guidance.stereotactic for biopsy of Breast - right|Mammogram Guidance.stereotactic for biopsy of Breast - right
C2826012|T102|strict|36928-0|LNC|CT Guidance.stereotactic for biopsy of Head|CT Guidance.stereotactic for biopsy of Head
C2826012|T102|strict|46296-0|LNC|Mammogram Guidance.stereotactic for core needle biopsy of Breast|Mammogram Guidance.stereotactic for core needle biopsy of Breast
C2826012|T102|strict|46295-2|LNC|Mammogram Guidance.stereotactic for core needle biopsy of Breast - left|Mammogram Guidance.stereotactic for core needle biopsy of Breast - left
C2826012|T102|strict|42433-3|LNC|Mammogram Guidance.stereotactic for core needle biopsy of Breast - right|Mammogram Guidance.stereotactic for core needle biopsy of Breast - right
C2826012|T102|strict|69160-0|LNC|Mammogram Guidance.stereotactic for needle biopsy of Breast|Mammogram Guidance.stereotactic for needle biopsy of Breast
C2826012|T102|strict|24585-2|LNC|CT Guidance.stereotactic for biopsy of Head-- W contrast IV|CT Guidance.stereotactic for biopsy of Head-- W contrast IV
C2826012|T102|strict|36929-8|LNC|CT Guidance.stereotactic for biopsy of Head-- WO contrast|CT Guidance.stereotactic for biopsy of Head-- WO contrast
C2826012|T102|strict|44122-0|LNC|MRI Guidance.stereotactic for localization in Brain-- W and WO contrast IV|MRI Guidance.stereotactic for localization in Brain-- W and WO contrast IV
C2826012|T102|strict|30656-3|LNC|MRI Guidance.stereotactic for localization in Brain-- W contrast IV|MRI Guidance.stereotactic for localization in Brain-- W contrast IV
C2826012|T102|strict|30800-7|LNC|MRI Guidance.stereotactic for localization in Brain-- WO contrast|MRI Guidance.stereotactic for localization in Brain-- WO contrast
C2826012|T102|strict|28632-8|LNC|Heterophoria study|Heterophoria study
C2826012|T102|strict|46264-8|LNC|History of medical device use|History of medical device use
C2826012|T102|strict|47519-4|LNC|History of Procedures Document|History of Procedures Document
C2826012|T102|strict|47245-6|LNC|HIV treatment form Document|HIV treatment form Document
C2826012|T102|strict|52035-3|LNC|Home health claims|Home health claims
C2826012|T102|strict|52036-1|LNC|Home health prior authorization|Home health prior authorization
C2826012|T102|strict|52046-0|LNC|Hospital beds|Hospital beds
C2826012|T102|strict|18841-7|LNC|Hospital consultations Document|Hospital consultations Document
C2826012|T102|strict|52028-8|LNC|Hysterectomy consent|Hysterectomy consent
C2826012|T102|strict|24655-3|LNC|Chest Fluoroscopy Image intensifier during surgery|Chest Fluoroscopy Image intensifier during surgery
C2826012|T102|strict|52047-8|LNC|Immunosuppressive drugs|Immunosuppressive drugs
C2826012|T102|strict|65806-2|LNC|Inhalation challenge test report Document --W methacholine inhaled|Inhalation challenge test report Document --W methacholine inhaled
C2826012|T102|strict|11500-6|LNC|Occupational therapy Initial assessment note at First encounter|Occupational therapy Initial assessment note at First encounter
C2826012|T102|strict|11495-9|LNC|Physical therapy Initial assessment note at First encounter|Physical therapy Initial assessment note at First encounter
C2826012|T102|strict|11494-2|LNC|Physician Initial assessment note at First encounter|Physician Initial assessment note at First encounter
C2826012|T102|strict|11496-7|LNC|Podiatry Initial assessment note at First encounter|Podiatry Initial assessment note at First encounter
C2826012|T102|strict|11497-5|LNC|Psychology Initial assessment note at First encounter|Psychology Initial assessment note at First encounter
C2826012|T102|strict|11498-3|LNC|Social work Initial assessment note at First encounter|Social work Initial assessment note at First encounter
C2826012|T102|strict|28572-6|LNC|Dentist Initial assessment note|Dentist Initial assessment note
C2826012|T102|strict|28621-1|LNC|Nurse practitioner Initial assessment note|Nurse practitioner Initial assessment note
C2826012|T102|strict|29753-1|LNC|Nurse Initial assessment note|Nurse Initial assessment note
C2826012|T102|strict|18734-4|LNC|Occupational therapy Initial assessment note|Occupational therapy Initial assessment note
C2826012|T102|strict|18735-1|LNC|Physical therapy Initial assessment note|Physical therapy Initial assessment note
C2826012|T102|strict|18736-9|LNC|Physician Initial assessment note|Physician Initial assessment note
C2826012|T102|strict|28654-2|LNC|Physician attending Initial assessment note|Physician attending Initial assessment note
C2826012|T102|strict|18763-3|LNC|Physician consulting Initial assessment note|Physician consulting Initial assessment note
C2826012|T102|strict|18737-7|LNC|Podiatry Initial assessment note|Podiatry Initial assessment note
C2826012|T102|strict|28635-1|LNC|Psychiatry Initial assessment note|Psychiatry Initial assessment note
C2826012|T102|strict|18738-5|LNC|Psychology Initial assessment note|Psychology Initial assessment note
C2826012|T102|strict|18739-3|LNC|Social work Initial assessment note|Social work Initial assessment note
C2826012|T102|strict|46214-3|LNC|Intracardiac ablation study|Intracardiac ablation study
C2826012|T102|strict|15508-5|LNC|Labor and delivery records|Labor and delivery records
C2826012|T102|strict|11502-2|LNC|Laboratory report|Laboratory report
C2826012|T102|strict|24717-1|LNC|Ileal conduit X-ray Loopogram|Ileal conduit X-ray Loopogram
C2826012|T102|strict|52048-6|LNC|Lymphedema pumps|Lymphedema pumps
C2826012|T102|strict|52049-4|LNC|Manual wheelchair|Manual wheelchair
C2826012|T102|strict|55186-1|LNC|Measure Document|Measure Document
C2826012|T102|strict|55185-3|LNC|Measure set Document|Measure set Document
C2826012|T102|strict|11503-0|LNC|Medical records|Medical records
C2826012|T102|strict|52037-9|LNC|Member ID card copy|Member ID card copy
C2826012|T102|strict|24672-8|LNC|Diaphragm US Motion|Diaphragm US Motion
C2826012|T102|strict|30632-4|LNC|Diaphragm Fluoroscopy Motion|Diaphragm Fluoroscopy Motion
C2826012|T102|strict|52050-2|LNC|Motorized wheelchair|Motorized wheelchair
C2826012|T102|strict|35990-1|LNC|Fetal MRI|Fetal MRI
C2826012|T102|strict|41806-1|LNC|Abdomen CT|Abdomen CT
C2826012|T102|strict|24556-3|LNC|Abdomen MRI|Abdomen MRI
C2826012|T102|strict|24558-9|LNC|Abdomen US|Abdomen US
C2826012|T102|strict|30762-9|LNC|Abdomen X-ray tomograph|Abdomen X-ray tomograph
C2826012|T102|strict|24566-2|LNC|Abdomen retroperitoneum CT|Abdomen retroperitoneum CT
C2826012|T102|strict|24531-6|LNC|Abdomen retroperitoneum US|Abdomen retroperitoneum US
C2826012|T102|strict|24532-4|LNC|Abdomen RUQ US|Abdomen RUQ US
C2826012|T102|strict|44115-4|LNC|Abdomen and Pelvis CT|Abdomen and Pelvis CT
C2826012|T102|strict|36781-3|LNC|Abdominal veins MRI angiogram|Abdominal veins MRI angiogram
C2826012|T102|strict|30864-3|LNC|Abdominal veins and IVC MRI angiogram|Abdominal veins and IVC MRI angiogram
C2826012|T102|strict|36791-2|LNC|Abdominal vessels MRI angiogram|Abdominal vessels MRI angiogram
C2826012|T102|strict|24534-0|LNC|Abdominal vessels US.doppler|Abdominal vessels US.doppler
C2826012|T102|strict|39494-0|LNC|Abdominal wall US|Abdominal wall US
C2826012|T102|strict|36930-6|LNC|Adrenal gland CT|Adrenal gland CT
C2826012|T102|strict|36931-4|LNC|Adrenal gland MRI|Adrenal gland MRI
C2826012|T102|strict|69277-2|LNC|Adrenal gland US|Adrenal gland US
C2826012|T102|strict|36792-0|LNC|Adrenal vessels MRI angiogram|Adrenal vessels MRI angiogram
C2826012|T102|strict|35940-6|LNC|Ankle CT|Ankle CT
C2826012|T102|strict|24538-1|LNC|Ankle MRI|Ankle MRI
C2826012|T102|strict|35939-8|LNC|Ankle X-ray tomograph|Ankle X-ray tomograph
C2826012|T102|strict|35941-4|LNC|Ankle - bilateral CT|Ankle - bilateral CT
C2826012|T102|strict|26208-9|LNC|Ankle - bilateral MRI|Ankle - bilateral MRI
C2826012|T102|strict|35942-2|LNC|Ankle - left CT|Ankle - left CT
C2826012|T102|strict|26209-7|LNC|Ankle - left MRI|Ankle - left MRI
C2826012|T102|strict|35943-0|LNC|Ankle - left X-ray tomograph|Ankle - left X-ray tomograph
C2826012|T102|strict|35944-8|LNC|Ankle - right CT|Ankle - right CT
C2826012|T102|strict|26210-5|LNC|Ankle - right MRI|Ankle - right MRI
C2826012|T102|strict|37674-9|LNC|Ankle - right X-ray tomograph|Ankle - right X-ray tomograph
C2826012|T102|strict|37222-7|LNC|Ankle and Foot MRI|Ankle and Foot MRI
C2826012|T102|strict|24542-3|LNC|Anus US|Anus US
C2826012|T102|strict|35945-5|LNC|Aorta CT|Aorta CT
C2826012|T102|strict|35947-1|LNC|Aorta MRI|Aorta MRI
C2826012|T102|strict|35946-3|LNC|Aorta MRI angiogram|Aorta MRI angiogram
C2826012|T102|strict|24547-2|LNC|Aorta US|Aorta US
C2826012|T102|strict|46388-5|LNC|Aorta US.doppler|Aorta US.doppler
C2826012|T102|strict|35948-9|LNC|Aorta abdominal CT|Aorta abdominal CT
C2826012|T102|strict|35949-7|LNC|Aorta abdominal MRI|Aorta abdominal MRI
C2826012|T102|strict|69276-4|LNC|Aorta abdominal US|Aorta abdominal US
C2826012|T102|strict|37216-9|LNC|Aorta.endograft CT|Aorta.endograft CT
C2826012|T102|strict|24544-9|LNC|Aorta thoracic CT|Aorta thoracic CT
C2826012|T102|strict|35950-5|LNC|Aorta thoracic MRI|Aorta thoracic MRI
C2826012|T102|strict|24660-3|LNC|Aorta thoracic MRI angiogram|Aorta thoracic MRI angiogram
C2826012|T102|strict|30863-5|LNC|Abdominal Aorta and Arteries MRI angiogram|Abdominal Aorta and Arteries MRI angiogram
C2826012|T102|strict|35951-3|LNC|Aortic arch MRI angiogram|Aortic arch MRI angiogram
C2826012|T102|strict|30861-9|LNC|Aortic arch and Neck vessels MRI angiogram|Aortic arch and Neck vessels MRI angiogram
C2826012|T102|strict|35952-1|LNC|Appendix CT|Appendix CT
C2826012|T102|strict|24548-0|LNC|Appendix US|Appendix US
C2826012|T102|strict|39040-1|LNC|AV fistula US|AV fistula US
C2826012|T102|strict|43508-1|LNC|Axilla - left MRI|Axilla - left MRI
C2826012|T102|strict|72529-1|LNC|Axilla - left US|Axilla - left US
C2826012|T102|strict|43510-7|LNC|Axilla - right MRI|Axilla - right MRI
C2826012|T102|strict|72528-3|LNC|Axilla - right US|Axilla - right US
C2826012|T102|strict|37219-3|LNC|Biliary ducts MRI|Biliary ducts MRI
C2826012|T102|strict|38021-2|LNC|Biliary ducts and Gallbladder US|Biliary ducts and Gallbladder US
C2826012|T102|strict|37220-1|LNC|Biliary ducts and Pancreatic duct MRI|Biliary ducts and Pancreatic duct MRI
C2826012|T102|strict|39039-3|LNC|Brachiocephalic artery US.doppler|Brachiocephalic artery US.doppler
C2826012|T102|strict|24590-2|LNC|Brain MRI|Brain MRI
C2826012|T102|strict|58748-5|LNC|Brain Functional MRI|Brain Functional MRI
C2826012|T102|strict|44138-6|LNC|Brain PET|Brain PET
C2826012|T102|strict|37217-7|LNC|Brain Stem and Nerves.cranial MRI|Brain Stem and Nerves.cranial MRI
C2826012|T102|strict|37218-5|LNC|Brain.temporal MRI|Brain.temporal MRI
C2826012|T102|strict|43772-3|LNC|Brain and Internal auditory canal MRI|Brain and Internal auditory canal MRI
C2826012|T102|strict|42385-5|LNC|Brain and Pituitary and Sella turcica MRI|Brain and Pituitary and Sella turcica MRI
C2826012|T102|strict|30794-2|LNC|Breast MRI|Breast MRI
C2826012|T102|strict|24601-7|LNC|Breast US|Breast US
C2826012|T102|strict|69165-9|LNC|Breast implant - bilateral MRI|Breast implant - bilateral MRI
C2826012|T102|strict|38057-6|LNC|Breast implant - left MRI|Breast implant - left MRI
C2826012|T102|strict|38058-4|LNC|Breast implant - right MRI|Breast implant - right MRI
C2826012|T102|strict|24596-9|LNC|Breast specimen US|Breast specimen US
C2826012|T102|strict|69397-8|LNC|Breast vessels US.doppler|Breast vessels US.doppler
C2826012|T102|strict|30795-9|LNC|Breast - bilateral MRI|Breast - bilateral MRI
C2826012|T102|strict|26214-7|LNC|Breast - bilateral US|Breast - bilateral US
C2826012|T102|strict|35954-7|LNC|Breast - left MRI|Breast - left MRI
C2826012|T102|strict|26215-4|LNC|Breast - left US|Breast - left US
C2826012|T102|strict|35955-4|LNC|Breast - right MRI|Breast - right MRI
C2826012|T102|strict|26216-2|LNC|Breast - right US|Breast - right US
C2826012|T102|strict|46299-4|LNC|Breast - unilateral MRI|Breast - unilateral MRI
C2826012|T102|strict|36010-7|LNC|Calcaneus CT|Calcaneus CT
C2826012|T102|strict|36011-5|LNC|Calcaneus X-ray tomograph|Calcaneus X-ray tomograph
C2826012|T102|strict|24616-5|LNC|Carotid artery US|Carotid artery US
C2826012|T102|strict|42146-1|LNC|Carotid artery US.doppler|Carotid artery US.doppler
C2826012|T102|strict|26217-0|LNC|Carotid artery - bilateral US|Carotid artery - bilateral US
C2826012|T102|strict|43765-7|LNC|Carotid artery - bilateral US.doppler|Carotid artery - bilateral US.doppler
C2826012|T102|strict|26218-8|LNC|Carotid artery - left US|Carotid artery - left US
C2826012|T102|strict|39427-0|LNC|Carotid artery - left US.doppler|Carotid artery - left US.doppler
C2826012|T102|strict|26219-6|LNC|Carotid artery - right US|Carotid artery - right US
C2826012|T102|strict|39437-9|LNC|Carotid artery - right US.doppler|Carotid artery - right US.doppler
C2826012|T102|strict|43552-9|LNC|Carotid artery - unilateral US|Carotid artery - unilateral US
C2826012|T102|strict|36793-8|LNC|Carotid vessel MRI angiogram|Carotid vessel MRI angiogram
C2826012|T102|strict|30859-3|LNC|Carotid vessels and Neck Vessels MRI angiogram|Carotid vessels and Neck Vessels MRI angiogram
C2826012|T102|strict|30865-0|LNC|Celiac vessels and Superior mesenteric Vessels MRI angiogram|Celiac vessels and Superior mesenteric Vessels MRI angiogram
C2826012|T102|strict|46374-5|LNC|Cerebral artery US|Cerebral artery US
C2826012|T102|strict|24627-2|LNC|Chest CT|Chest CT
C2826012|T102|strict|24629-8|LNC|Chest MRI|Chest MRI
C2826012|T102|strict|24630-6|LNC|Chest US|Chest US
C2826012|T102|strict|24657-9|LNC|Chest X-ray tomograph|Chest X-ray tomograph
C2826012|T102|strict|30862-7|LNC|Chest vessels MRI angiogram|Chest vessels MRI angiogram
C2826012|T102|strict|38016-2|LNC|Chest wall US|Chest wall US
C2826012|T102|strict|37235-9|LNC|Circle of Willis MRI angiogram|Circle of Willis MRI angiogram
C2826012|T102|strict|35960-4|LNC|Clavicle CT|Clavicle CT
C2826012|T102|strict|35961-2|LNC|Clavicle MRI|Clavicle MRI
C2826012|T102|strict|35959-6|LNC|Clavicle X-ray tomograph|Clavicle X-ray tomograph
C2826012|T102|strict|44120-4|LNC|Colon CT|Colon CT
C2826012|T102|strict|24757-7|LNC|Coronary arteries CT fast|Coronary arteries CT fast
C2826012|T102|strict|35962-0|LNC|Elbow CT|Elbow CT
C2826012|T102|strict|24674-4|LNC|Elbow MRI|Elbow MRI
C2826012|T102|strict|35963-8|LNC|Elbow X-ray tomograph|Elbow X-ray tomograph
C2826012|T102|strict|35965-3|LNC|Elbow - bilateral CT|Elbow - bilateral CT
C2826012|T102|strict|26220-4|LNC|Elbow - bilateral MRI|Elbow - bilateral MRI
C2826012|T102|strict|35964-6|LNC|Elbow - bilateral X-ray tomograph|Elbow - bilateral X-ray tomograph
C2826012|T102|strict|35966-1|LNC|Elbow - left CT|Elbow - left CT
C2826012|T102|strict|26221-2|LNC|Elbow - left MRI|Elbow - left MRI
C2826012|T102|strict|35967-9|LNC|Elbow - left X-ray tomograph|Elbow - left X-ray tomograph
C2826012|T102|strict|35968-7|LNC|Elbow - right CT|Elbow - right CT
C2826012|T102|strict|26222-0|LNC|Elbow - right MRI|Elbow - right MRI
C2826012|T102|strict|37688-9|LNC|Elbow - right X-ray tomograph|Elbow - right X-ray tomograph
C2826012|T102|strict|35969-5|LNC|Esophagus CT|Esophagus CT
C2826012|T102|strict|57823-7|LNC|Esophagus PET|Esophagus PET
C2826012|T102|strict|24690-0|LNC|Extremity CT|Extremity CT
C2826012|T102|strict|69193-1|LNC|Extremity MRI|Extremity MRI
C2826012|T102|strict|24693-4|LNC|Extremity US|Extremity US
C2826012|T102|strict|35970-3|LNC|Extremity X-ray tomograph|Extremity X-ray tomograph
C2826012|T102|strict|39042-7|LNC|Extremity artery US.doppler|Extremity artery US.doppler
C2826012|T102|strict|39031-0|LNC|Extremity artery - bilateral US.doppler|Extremity artery - bilateral US.doppler
C2826012|T102|strict|69293-9|LNC|Extremity artery - left US|Extremity artery - left US
C2826012|T102|strict|39428-8|LNC|Extremity artery - left US.doppler|Extremity artery - left US.doppler
C2826012|T102|strict|69297-0|LNC|Extremity artery - right US|Extremity artery - right US
C2826012|T102|strict|39439-5|LNC|Extremity artery - right US.doppler|Extremity artery - right US.doppler
C2826012|T102|strict|39449-4|LNC|Extremity vein US.doppler|Extremity vein US.doppler
C2826012|T102|strict|39418-9|LNC|Extremity vein - bilateral US.doppler|Extremity vein - bilateral US.doppler
C2826012|T102|strict|42145-3|LNC|Extremity vein - left US|Extremity vein - left US
C2826012|T102|strict|39429-6|LNC|Extremity vein - left US.doppler|Extremity vein - left US.doppler
C2826012|T102|strict|42144-6|LNC|Extremity vein - right US|Extremity vein - right US
C2826012|T102|strict|39440-3|LNC|Extremity vein - right US.doppler|Extremity vein - right US.doppler
C2826012|T102|strict|30876-7|LNC|Extremity veins MRI angiogram|Extremity veins MRI angiogram
C2826012|T102|strict|69283-0|LNC|Extremity veins - bilateral US.doppler|Extremity veins - bilateral US.doppler
C2826012|T102|strict|41835-0|LNC|Extremity veins - left US|Extremity veins - left US
C2826012|T102|strict|41816-0|LNC|Extremity veins - right US|Extremity veins - right US
C2826012|T102|strict|36794-6|LNC|Extremity vessels MRI angiogram|Extremity vessels MRI angiogram
C2826012|T102|strict|43771-5|LNC|Extremity vessels US.doppler|Extremity vessels US.doppler
C2826012|T102|strict|39495-7|LNC|Extremity vessels - bilateral US.doppler|Extremity vessels - bilateral US.doppler
C2826012|T102|strict|69398-6|LNC|Extremity vessels Left US.doppler|Extremity vessels Left US.doppler
C2826012|T102|strict|39503-8|LNC|Extremity vessels - right US.doppler|Extremity vessels - right US.doppler
C2826012|T102|strict|26224-6|LNC|Extremity - bilateral CT|Extremity - bilateral CT
C2826012|T102|strict|26223-8|LNC|Extremity - bilateral US|Extremity - bilateral US
C2826012|T102|strict|26226-1|LNC|Extremity - left CT|Extremity - left CT
C2826012|T102|strict|26225-3|LNC|Extremity - left US|Extremity - left US
C2826012|T102|strict|26231-1|LNC|Extremity - right CT|Extremity - right CT
C2826012|T102|strict|26230-3|LNC|Extremity - right US|Extremity - right US
C2826012|T102|strict|24853-4|LNC|Eye+Orbit - bilateral US|Eye+Orbit - bilateral US
C2826012|T102|strict|35953-9|LNC|Face MRI|Face MRI
C2826012|T102|strict|41808-7|LNC|Facial bones and Maxilla CT|Facial bones and Maxilla CT
C2826012|T102|strict|24696-7|LNC|Facial bones and Sinuses CT|Facial bones and Sinuses CT
C2826012|T102|strict|69389-5|LNC|Femoral artery and Popliteal artery US|Femoral artery and Popliteal artery US
C2826012|T102|strict|69399-4|LNC|Femoral vein and Popliteal vein US|Femoral vein and Popliteal vein US
C2826012|T102|strict|30871-8|LNC|Femoral vessels MRI angiogram|Femoral vessels MRI angiogram
C2826012|T102|strict|38134-3|LNC|Femoral vessels US|Femoral vessels US
C2826012|T102|strict|38128-5|LNC|Femoral vessels - bilateral US|Femoral vessels - bilateral US
C2826012|T102|strict|39498-1|LNC|Femoral vessels - left US.doppler|Femoral vessels - left US.doppler
C2826012|T102|strict|39504-6|LNC|Femoral vessels - right US.doppler|Femoral vessels - right US.doppler
C2826012|T102|strict|35984-4|LNC|Femur CT|Femur CT
C2826012|T102|strict|35985-1|LNC|Femur X-ray tomograph|Femur X-ray tomograph
C2826012|T102|strict|35986-9|LNC|Femur - bilateral X-ray tomograph|Femur - bilateral X-ray tomograph
C2826012|T102|strict|35987-7|LNC|Femur - left CT|Femur - left CT
C2826012|T102|strict|38037-8|LNC|Femur - left US|Femur - left US
C2826012|T102|strict|35988-5|LNC|Femur - left X-ray tomograph|Femur - left X-ray tomograph
C2826012|T102|strict|35989-3|LNC|Femur - right CT|Femur - right CT
C2826012|T102|strict|38048-5|LNC|Femur - right US|Femur - right US
C2826012|T102|strict|38768-8|LNC|Femur - right X-ray tomograph|Femur - right X-ray tomograph
C2826012|T102|strict|24705-6|LNC|Finger MRI|Finger MRI
C2826012|T102|strict|26238-6|LNC|Finger - bilateral MRI|Finger - bilateral MRI
C2826012|T102|strict|26239-4|LNC|Finger - left MRI|Finger - left MRI
C2826012|T102|strict|26240-2|LNC|Finger - right MRI|Finger - right MRI
C2826012|T102|strict|37221-9|LNC|Fistula CT|Fistula CT
C2826012|T102|strict|35991-9|LNC|Foot CT|Foot CT
C2826012|T102|strict|24707-2|LNC|Foot MRI|Foot MRI
C2826012|T102|strict|35992-7|LNC|Foot X-ray tomograph|Foot X-ray tomograph
C2826012|T102|strict|30872-6|LNC|Foot vessels MRI angiogram|Foot vessels MRI angiogram
C2826012|T102|strict|46362-0|LNC|Foot vessels US.doppler|Foot vessels US.doppler
C2826012|T102|strict|35993-5|LNC|Foot - bilateral CT|Foot - bilateral CT
C2826012|T102|strict|26241-0|LNC|Foot - bilateral MRI|Foot - bilateral MRI
C2826012|T102|strict|35994-3|LNC|Foot - left CT|Foot - left CT
C2826012|T102|strict|26242-8|LNC|Foot - left MRI|Foot - left MRI
C2826012|T102|strict|35995-0|LNC|Foot - left X-ray tomograph|Foot - left X-ray tomograph
C2826012|T102|strict|35996-8|LNC|Foot - right CT|Foot - right CT
C2826012|T102|strict|26243-6|LNC|Foot - right MRI|Foot - right MRI
C2826012|T102|strict|37706-9|LNC|Foot - right X-ray tomograph|Foot - right X-ray tomograph
C2826012|T102|strict|35997-6|LNC|Forearm CT|Forearm CT
C2826012|T102|strict|24710-6|LNC|Forearm MRI|Forearm MRI
C2826012|T102|strict|30873-4|LNC|Forearm vessels MRI angiogram|Forearm vessels MRI angiogram
C2826012|T102|strict|35998-4|LNC|Forearm - bilateral CT|Forearm - bilateral CT
C2826012|T102|strict|26244-4|LNC|Forearm - bilateral MRI|Forearm - bilateral MRI
C2826012|T102|strict|35999-2|LNC|Forearm - left CT|Forearm - left CT
C2826012|T102|strict|26245-1|LNC|Forearm - left MRI|Forearm - left MRI
C2826012|T102|strict|36000-8|LNC|Forearm - right CT|Forearm - right CT
C2826012|T102|strict|26246-9|LNC|Forearm - right MRI|Forearm - right MRI
C2826012|T102|strict|24711-4|LNC|Gallbladder US|Gallbladder US
C2826012|T102|strict|36001-6|LNC|Gallbladder X-ray tomograph|Gallbladder X-ray tomograph
C2826012|T102|strict|39415-5|LNC|Gastrointestine US|Gastrointestine US
C2826012|T102|strict|39416-3|LNC|Genitourinary system US|Genitourinary system US
C2826012|T102|strict|37236-7|LNC|Great vessel MRI|Great vessel MRI
C2826012|T102|strict|24719-7|LNC|Groin US|Groin US
C2826012|T102|strict|36002-4|LNC|Hand CT|Hand CT
C2826012|T102|strict|24720-5|LNC|Hand MRI|Hand MRI
C2826012|T102|strict|36003-2|LNC|Hand X-ray tomograph|Hand X-ray tomograph
C2826012|T102|strict|46382-8|LNC|Hand vessels US.doppler|Hand vessels US.doppler
C2826012|T102|strict|36004-0|LNC|Hand - bilateral CT|Hand - bilateral CT
C2826012|T102|strict|26247-7|LNC|Hand - bilateral MRI|Hand - bilateral MRI
C2826012|T102|strict|36005-7|LNC|Hand - left CT|Hand - left CT
C2826012|T102|strict|26248-5|LNC|Hand - left MRI|Hand - left MRI
C2826012|T102|strict|36006-5|LNC|Hand - left X-ray tomograph|Hand - left X-ray tomograph
C2826012|T102|strict|36007-3|LNC|Hand - right CT|Hand - right CT
C2826012|T102|strict|26249-3|LNC|Hand - right MRI|Hand - right MRI
C2826012|T102|strict|37717-6|LNC|Hand - right X-ray tomograph|Hand - right X-ray tomograph
C2826012|T102|strict|24725-4|LNC|Head CT|Head CT
C2826012|T102|strict|24728-8|LNC|Head CT cine|Head CT cine
C2826012|T102|strict|24731-2|LNC|Head US|Head US
C2826012|T102|strict|58741-0|LNC|Head to thigh PET|Head to thigh PET
C2826012|T102|strict|30858-5|LNC|Head veins MRI angiogram|Head veins MRI angiogram
C2826012|T102|strict|30856-9|LNC|Head vessels MRI angiogram|Head vessels MRI angiogram
C2826012|T102|strict|24733-8|LNC|Head vessels US.doppler|Head vessels US.doppler
C2826012|T102|strict|42304-6|LNC|Head vessels and Neck vessels MRI angiogram|Head vessels and Neck vessels MRI angiogram
C2826012|T102|strict|30880-9|LNC|Head vessels and Neck vessels US.doppler|Head vessels and Neck vessels US.doppler
C2826012|T102|strict|30655-5|LNC|Head Cistern MRI|Head Cistern MRI
C2826012|T102|strict|24746-0|LNC|Head Sagittal Sinus MRI|Head Sagittal Sinus MRI
C2826012|T102|strict|58742-8|LNC|Head and Neck PET|Head and Neck PET
C2826012|T102|strict|44164-2|LNC|Head and Neck US|Head and Neck US
C2826012|T102|strict|58744-4|LNC|Heart CT|Heart CT
C2826012|T102|strict|24748-6|LNC|Heart MRI|Heart MRI
C2826012|T102|strict|36009-9|LNC|Heart MRI angiogram|Heart MRI angiogram
C2826012|T102|strict|44137-8|LNC|Heart PET|Heart PET
C2826012|T102|strict|42148-7|LNC|Heart US|Heart US
C2826012|T102|strict|36014-9|LNC|Hip CT|Hip CT
C2826012|T102|strict|36013-1|LNC|Hip MRI|Hip MRI
C2826012|T102|strict|24760-1|LNC|Hip US|Hip US
C2826012|T102|strict|36012-3|LNC|Hip X-ray tomograph|Hip X-ray tomograph
C2826012|T102|strict|36016-4|LNC|Hip - bilateral CT|Hip - bilateral CT
C2826012|T102|strict|36017-2|LNC|Hip - bilateral MRI|Hip - bilateral MRI
C2826012|T102|strict|26250-1|LNC|Hip - bilateral US|Hip - bilateral US
C2826012|T102|strict|36015-6|LNC|Hip - bilateral X-ray tomograph|Hip - bilateral X-ray tomograph
C2826012|T102|strict|36018-0|LNC|Hip - left CT|Hip - left CT
C2826012|T102|strict|36020-6|LNC|Hip - left MRI|Hip - left MRI
C2826012|T102|strict|26251-9|LNC|Hip - left US|Hip - left US
C2826012|T102|strict|36019-8|LNC|Hip - left X-ray tomograph|Hip - left X-ray tomograph
C2826012|T102|strict|36021-4|LNC|Hip - right CT|Hip - right CT
C2826012|T102|strict|36022-2|LNC|Hip - right MRI|Hip - right MRI
C2826012|T102|strict|26252-7|LNC|Hip - right US|Hip - right US
C2826012|T102|strict|37735-8|LNC|Hip - right X-ray tomograph|Hip - right X-ray tomograph
C2826012|T102|strict|43566-9|LNC|Hip and Thigh US|Hip and Thigh US
C2826012|T102|strict|36024-8|LNC|Humerus X-ray tomograph|Humerus X-ray tomograph
C2826012|T102|strict|39425-4|LNC|Iliac artery US.doppler|Iliac artery US.doppler
C2826012|T102|strict|42147-9|LNC|Iliac graft US.doppler|Iliac graft US.doppler
C2826012|T102|strict|39497-3|LNC|Iliac vessels US.doppler|Iliac vessels US.doppler
C2826012|T102|strict|38129-3|LNC|Iliac vessels - bilateral US|Iliac vessels - bilateral US
C2826012|T102|strict|38137-6|LNC|Iliac vessels - left US|Iliac vessels - left US
C2826012|T102|strict|38141-8|LNC|Iliac vessels - right US|Iliac vessels - right US
C2826012|T102|strict|35958-8|LNC|Internal auditory canal CT|Internal auditory canal CT
C2826012|T102|strict|35956-2|LNC|Internal auditory canal MRI|Internal auditory canal MRI
C2826012|T102|strict|24767-6|LNC|Internal auditory canal X-ray tomograph|Internal auditory canal X-ray tomograph
C2826012|T102|strict|26253-5|LNC|Internal auditory canal - bilateral X-ray tomograph|Internal auditory canal - bilateral X-ray tomograph
C2826012|T102|strict|35957-0|LNC|Internal auditory canal - left CT|Internal auditory canal - left CT
C2826012|T102|strict|26254-3|LNC|Internal auditory canal - left X-ray tomograph|Internal auditory canal - left X-ray tomograph
C2826012|T102|strict|38767-0|LNC|Internal auditory canal - right CT|Internal auditory canal - right CT
C2826012|T102|strict|26255-0|LNC|Internal auditory canal - right X-ray tomograph|Internal auditory canal - right X-ray tomograph
C2826012|T102|strict|24735-3|LNC|Internal auditory canal and Posterior fossa MRI|Internal auditory canal and Posterior fossa MRI
C2826012|T102|strict|36033-9|LNC|Kidney MRI|Kidney MRI
C2826012|T102|strict|38036-0|LNC|Kidney US|Kidney US
C2826012|T102|strict|36032-1|LNC|Kidney X-ray tomograph|Kidney X-ray tomograph
C2826012|T102|strict|39032-8|LNC|Kidney transplant US|Kidney transplant US
C2826012|T102|strict|42477-0|LNC|Kidney vessels transplant US.doppler|Kidney vessels transplant US.doppler
C2826012|T102|strict|43767-3|LNC|Kidney - bilateral CT|Kidney - bilateral CT
C2826012|T102|strict|36034-7|LNC|Kidney - bilateral MRI|Kidney - bilateral MRI
C2826012|T102|strict|43774-9|LNC|Kidney - bilateral US|Kidney - bilateral US
C2826012|T102|strict|24789-0|LNC|Kidney - bilateral X-ray tomograph|Kidney - bilateral X-ray tomograph
C2826012|T102|strict|69402-6|LNC|Kidney Bilateral and Bladder US|Kidney Bilateral and Bladder US
C2826012|T102|strict|36035-4|LNC|Kidney - left MRI|Kidney - left MRI
C2826012|T102|strict|38038-6|LNC|Kidney - left US|Kidney - left US
C2826012|T102|strict|69113-9|LNC|Kidney - right CT|Kidney - right CT
C2826012|T102|strict|36036-2|LNC|Kidney - right MRI|Kidney - right MRI
C2826012|T102|strict|38049-3|LNC|Kidney - right US|Kidney - right US
C2826012|T102|strict|36037-0|LNC|Knee CT|Knee CT
C2826012|T102|strict|24802-1|LNC|Knee MRI|Knee MRI
C2826012|T102|strict|36038-8|LNC|Knee X-ray tomograph|Knee X-ray tomograph
C2826012|T102|strict|36799-5|LNC|Knee vessels MRI angiogram|Knee vessels MRI angiogram
C2826012|T102|strict|36800-1|LNC|Knee vessels - left MRI angiogram|Knee vessels - left MRI angiogram
C2826012|T102|strict|36801-9|LNC|Knee vessels - right MRI angiogram|Knee vessels - right MRI angiogram
C2826012|T102|strict|36040-4|LNC|Knee - bilateral CT|Knee - bilateral CT
C2826012|T102|strict|26256-8|LNC|Knee - bilateral MRI|Knee - bilateral MRI
C2826012|T102|strict|36039-6|LNC|Knee - bilateral X-ray tomograph|Knee - bilateral X-ray tomograph
C2826012|T102|strict|36041-2|LNC|Knee - left CT|Knee - left CT
C2826012|T102|strict|26257-6|LNC|Knee - left MRI|Knee - left MRI
C2826012|T102|strict|36042-0|LNC|Knee - left X-ray tomograph|Knee - left X-ray tomograph
C2826012|T102|strict|36043-8|LNC|Knee - right CT|Knee - right CT
C2826012|T102|strict|26258-4|LNC|Knee - right MRI|Knee - right MRI
C2826012|T102|strict|37760-6|LNC|Knee - right X-ray tomograph|Knee - right X-ray tomograph
C2826012|T102|strict|36045-3|LNC|Larynx MRI|Larynx MRI
C2826012|T102|strict|36044-6|LNC|Larynx X-ray tomograph|Larynx X-ray tomograph
C2826012|T102|strict|24814-6|LNC|Liver CT|Liver CT
C2826012|T102|strict|36046-1|LNC|Liver MRI|Liver MRI
C2826012|T102|strict|28614-6|LNC|Liver US|Liver US
C2826012|T102|strict|39454-4|LNC|Liver transplant US|Liver transplant US
C2826012|T102|strict|24818-7|LNC|Liver and Diaphragm US|Liver and Diaphragm US
C2826012|T102|strict|35971-1|LNC|Lower extremity CT|Lower extremity CT
C2826012|T102|strict|30692-8|LNC|Lower extremity MRI|Lower extremity MRI
C2826012|T102|strict|30709-0|LNC|Lower extremity US|Lower extremity US
C2826012|T102|strict|35972-9|LNC|Lower extremity X-ray tomograph|Lower extremity X-ray tomograph
C2826012|T102|strict|48693-6|LNC|Lower extremity artery US|Lower extremity artery US
C2826012|T102|strict|39434-6|LNC|Lower extremity artery US.doppler|Lower extremity artery US.doppler
C2826012|T102|strict|38130-1|LNC|Lower extremity artery - bilateral US|Lower extremity artery - bilateral US
C2826012|T102|strict|39421-3|LNC|Lower extremity artery - bilateral US.doppler|Lower extremity artery - bilateral US.doppler
C2826012|T102|strict|41834-3|LNC|Lower extremity artery - left US|Lower extremity artery - left US
C2826012|T102|strict|39499-9|LNC|Lower extremity artery - left US.doppler|Lower extremity artery - left US.doppler
C2826012|T102|strict|41815-2|LNC|Lower extremity artery - right US|Lower extremity artery - right US
C2826012|T102|strict|39505-3|LNC|Lower extremity artery - right US.doppler|Lower extremity artery - right US.doppler
C2826012|T102|strict|46363-8|LNC|Lower extremity vein US|Lower extremity vein US
C2826012|T102|strict|30881-7|LNC|Lower extremity vein US.doppler|Lower extremity vein US.doppler
C2826012|T102|strict|46364-6|LNC|Lower extremity vein - bilateral US|Lower extremity vein - bilateral US
C2826012|T102|strict|39420-5|LNC|Lower extremity vein - bilateral US.doppler|Lower extremity vein - bilateral US.doppler
C2826012|T102|strict|48692-8|LNC|Lower extremity vein - left US|Lower extremity vein - left US
C2826012|T102|strict|39432-0|LNC|Lower extremity vein - left US.doppler|Lower extremity vein - left US.doppler
C2826012|T102|strict|48691-0|LNC|Lower extremity vein - right US|Lower extremity vein - right US
C2826012|T102|strict|39443-7|LNC|Lower extremity vein - right US.doppler|Lower extremity vein - right US.doppler
C2826012|T102|strict|36079-2|LNC|Lower extremity veins MRI angiogram|Lower extremity veins MRI angiogram
C2826012|T102|strict|69385-3|LNC|Lower extremity veins - bilateral US|Lower extremity veins - bilateral US
C2826012|T102|strict|36784-7|LNC|Lower extremity veins - left MRI angiogram|Lower extremity veins - left MRI angiogram
C2826012|T102|strict|69392-9|LNC|Lower extremity veins - left US|Lower extremity veins - left US
C2826012|T102|strict|36785-4|LNC|Lower extremity veins - right MRI angiogram|Lower extremity veins - right MRI angiogram
C2826012|T102|strict|42461-4|LNC|Lower extremity vessel graft - left US.doppler|Lower extremity vessel graft - left US.doppler
C2826012|T102|strict|42462-2|LNC|Lower extremity vessel graft - right US.doppler|Lower extremity vessel graft - right US.doppler
C2826012|T102|strict|30874-2|LNC|Lower extremity vessels MRI angiogram|Lower extremity vessels MRI angiogram
C2826012|T102|strict|44174-1|LNC|Lower extremity vessels US.doppler|Lower extremity vessels US.doppler
C2826012|T102|strict|35974-5|LNC|Lower extremity vessels - bilateral MRI angiogram|Lower extremity vessels - bilateral MRI angiogram
C2826012|T102|strict|39422-1|LNC|Lower extremity vessels - bilateral US.doppler|Lower extremity vessels - bilateral US.doppler
C2826012|T102|strict|36795-3|LNC|Lower extremity vessels - left MRI angiogram|Lower extremity vessels - left MRI angiogram
C2826012|T102|strict|39431-2|LNC|Lower extremity vessels - left US.doppler|Lower extremity vessels - left US.doppler
C2826012|T102|strict|36796-1|LNC|Lower extremity vessels - right MRI angiogram|Lower extremity vessels - right MRI angiogram
C2826012|T102|strict|39442-9|LNC|Lower extremity vessels - right US.doppler|Lower extremity vessels - right US.doppler
C2826012|T102|strict|35973-7|LNC|Lower extremity - bilateral CT|Lower extremity - bilateral CT
C2826012|T102|strict|35975-2|LNC|Lower extremity - bilateral MRI|Lower extremity - bilateral MRI
C2826012|T102|strict|38013-9|LNC|Lower extremity - bilateral US|Lower extremity - bilateral US
C2826012|T102|strict|24687-6|LNC|Lower Extremity Joint MRI|Lower Extremity Joint MRI
C2826012|T102|strict|26227-9|LNC|Lower extremity joint - bilateral MRI|Lower extremity joint - bilateral MRI
C2826012|T102|strict|26228-7|LNC|Lower extremity joint - left MRI|Lower extremity joint - left MRI
C2826012|T102|strict|26229-5|LNC|Lower extremity joint - right MRI|Lower extremity joint - right MRI
C2826012|T102|strict|35976-0|LNC|Lower extremity - left CT|Lower extremity - left CT
C2826012|T102|strict|35978-6|LNC|Lower extremity - left MRI|Lower extremity - left MRI
C2826012|T102|strict|38040-2|LNC|Lower extremity - left US|Lower extremity - left US
C2826012|T102|strict|35977-8|LNC|Lower extremity - left X-ray tomograph|Lower extremity - left X-ray tomograph
C2826012|T102|strict|35979-4|LNC|Lower extremity - right CT|Lower extremity - right CT
C2826012|T102|strict|35980-2|LNC|Lower extremity - right MRI|Lower extremity - right MRI
C2826012|T102|strict|38051-9|LNC|Lower extremity - right US|Lower extremity - right US
C2826012|T102|strict|37766-3|LNC|Lower extremity - right X-ray tomograph|Lower extremity - right X-ray tomograph
C2826012|T102|strict|36074-3|LNC|Lower leg CT|Lower leg CT
C2826012|T102|strict|24821-1|LNC|Lower leg MRI|Lower leg MRI
C2826012|T102|strict|43513-1|LNC|Lower leg vessels - left MRI angiogram|Lower leg vessels - left MRI angiogram
C2826012|T102|strict|43556-0|LNC|Lower leg vessels - right MRI angiogram|Lower leg vessels - right MRI angiogram
C2826012|T102|strict|42696-5|LNC|Lower leg - bilateral MRI|Lower leg - bilateral MRI
C2826012|T102|strict|36075-0|LNC|Lower leg - left MRI|Lower leg - left MRI
C2826012|T102|strict|36076-8|LNC|Lower leg - right MRI|Lower leg - right MRI
C2826012|T102|strict|30866-8|LNC|Lumbar plexus MRI|Lumbar plexus MRI
C2826012|T102|strict|57822-9|LNC|Lung PET|Lung PET
C2826012|T102|strict|36047-9|LNC|Mandible CT|Mandible CT
C2826012|T102|strict|36048-7|LNC|Mandible X-ray tomograph|Mandible X-ray tomograph
C2826012|T102|strict|38043-6|LNC|Mastoid US|Mastoid US
C2826012|T102|strict|36776-3|LNC|Mastoid X-ray tomograph|Mastoid X-ray tomograph
C2826012|T102|strict|46298-6|LNC|Mastoid - bilateral CT|Mastoid - bilateral CT
C2826012|T102|strict|36050-3|LNC|Maxilla CT|Maxilla CT
C2826012|T102|strict|36049-5|LNC|Maxilla and Mandible CT|Maxilla and Mandible CT
C2826012|T102|strict|37234-2|LNC|Mediastinum MRI|Mediastinum MRI
C2826012|T102|strict|38044-4|LNC|Mediastinum US|Mediastinum US
C2826012|T102|strict|37233-4|LNC|Mediastinum X-ray tomograph|Mediastinum X-ray tomograph
C2826012|T102|strict|69394-5|LNC|Mesenteric artery US|Mesenteric artery US
C2826012|T102|strict|69211-1|LNC|Nasal bones MRI|Nasal bones MRI
C2826012|T102|strict|37606-1|LNC|Nasal bones X-ray tomograph|Nasal bones X-ray tomograph
C2826012|T102|strict|30860-1|LNC|Nasopharynx MRI|Nasopharynx MRI
C2826012|T102|strict|24835-1|LNC|Nasopharynx and Neck CT|Nasopharynx and Neck CT
C2826012|T102|strict|36051-1|LNC|Neck CT|Neck CT
C2826012|T102|strict|24839-3|LNC|Neck MRI|Neck MRI
C2826012|T102|strict|24842-7|LNC|Neck US|Neck US
C2826012|T102|strict|36788-8|LNC|Neck veins MRI angiogram|Neck veins MRI angiogram
C2826012|T102|strict|36085-9|LNC|Neck vessels MRI angiogram|Neck vessels MRI angiogram
C2826012|T102|strict|44175-8|LNC|Neck vessels US.doppler|Neck vessels US.doppler
C2826012|T102|strict|30857-7|LNC|Nerves cranial MRI|Nerves cranial MRI
C2826012|T102|strict|41807-9|LNC|Orbit CT|Orbit CT
C2826012|T102|strict|36777-1|LNC|Orbit MRI|Orbit MRI
C2826012|T102|strict|36802-7|LNC|Orbit vessels MRI angiogram|Orbit vessels MRI angiogram
C2826012|T102|strict|24848-4|LNC|Orbit - bilateral CT|Orbit - bilateral CT
C2826012|T102|strict|37611-1|LNC|Orbit - bilateral X-ray tomograph|Orbit - bilateral X-ray tomograph
C2826012|T102|strict|38836-3|LNC|Orbit - left MRI|Orbit - left MRI
C2826012|T102|strict|36778-9|LNC|Orbit - right MRI|Orbit - right MRI
C2826012|T102|strict|42303-8|LNC|Orbit and Face MRI|Orbit and Face MRI
C2826012|T102|strict|43530-5|LNC|Orbit and Face and Neck MRI|Orbit and Face and Neck MRI
C2826012|T102|strict|43455-5|LNC|Oropharynx MRI|Oropharynx MRI
C2826012|T102|strict|39502-0|LNC|Ovarian vessels US.doppler|Ovarian vessels US.doppler
C2826012|T102|strict|36779-7|LNC|Ovary MRI|Ovary MRI
C2826012|T102|strict|69390-3|LNC|Ovary US|Ovary US
C2826012|T102|strict|43506-5|LNC|Ovary - bilateral MRI|Ovary - bilateral MRI
C2826012|T102|strict|24857-5|LNC|Pancreas CT|Pancreas CT
C2826012|T102|strict|36052-9|LNC|Pancreas MRI|Pancreas MRI
C2826012|T102|strict|24859-1|LNC|Pancreas US|Pancreas US
C2826012|T102|strict|39509-5|LNC|Pancreas transplant US|Pancreas transplant US
C2826012|T102|strict|36053-7|LNC|Parathyroid MRI|Parathyroid MRI
C2826012|T102|strict|38045-1|LNC|Parathyroid US|Parathyroid US
C2826012|T102|strict|37223-5|LNC|Parotid gland CT|Parotid gland CT
C2826012|T102|strict|37224-3|LNC|Parotid gland MRI|Parotid gland MRI
C2826012|T102|strict|38138-4|LNC|Parotid gland US|Parotid gland US
C2826012|T102|strict|24865-8|LNC|Pelvis CT|Pelvis CT
C2826012|T102|strict|24867-4|LNC|Pelvis MRI|Pelvis MRI
C2826012|T102|strict|24869-0|LNC|Pelvis US|Pelvis US
C2826012|T102|strict|37632-7|LNC|Pelvis X-ray tomograph|Pelvis X-ray tomograph
C2826012|T102|strict|36789-6|LNC|Pelvis veins MRI angiogram|Pelvis veins MRI angiogram
C2826012|T102|strict|30867-6|LNC|Pelvis vessels MRI angiogram|Pelvis vessels MRI angiogram
C2826012|T102|strict|24870-8|LNC|Pelvis vessels US.doppler|Pelvis vessels US.doppler
C2826012|T102|strict|24872-4|LNC|Pelvis and Hip MRI|Pelvis and Hip MRI
C2826012|T102|strict|26259-2|LNC|Pelvis and Hip - bilateral MRI|Pelvis and Hip - bilateral MRI
C2826012|T102|strict|26260-0|LNC|Pelvis and Hip - left MRI|Pelvis and Hip - left MRI
C2826012|T102|strict|26261-8|LNC|Pelvis and Hip - right MRI|Pelvis and Hip - right MRI
C2826012|T102|strict|38140-0|LNC|Penis US|Penis US
C2826012|T102|strict|38139-2|LNC|Penis vessels US|Penis vessels US
C2826012|T102|strict|24877-3|LNC|Petrous bone CT|Petrous bone CT
C2826012|T102|strict|36932-2|LNC|Pituitary and Sella turcica CT|Pituitary and Sella turcica CT
C2826012|T102|strict|24880-7|LNC|Pituitary and Sella turcica MRI|Pituitary and Sella turcica MRI
C2826012|T102|strict|24881-5|LNC|Popliteal space US|Popliteal space US
C2826012|T102|strict|26262-6|LNC|Popliteal space - bilateral US|Popliteal space - bilateral US
C2826012|T102|strict|26263-4|LNC|Popliteal space - left US|Popliteal space - left US
C2826012|T102|strict|26264-2|LNC|Popliteal space - right US|Popliteal space - right US
C2826012|T102|strict|36077-6|LNC|Portal vein MRI angiogram|Portal vein MRI angiogram
C2826012|T102|strict|69284-8|LNC|Portal vein and Hepatic vein US.doppler|Portal vein and Hepatic vein US.doppler
C2826012|T102|strict|36055-2|LNC|Posterior fossa CT|Posterior fossa CT
C2826012|T102|strict|36056-0|LNC|Posterior fossa MRI|Posterior fossa MRI
C2826012|T102|strict|36057-8|LNC|Prostate CT|Prostate CT
C2826012|T102|strict|30675-3|LNC|Prostate MRI|Prostate MRI
C2826012|T102|strict|24884-9|LNC|Prostate US|Prostate US
C2826012|T102|strict|43445-6|LNC|Pulmonary system CT|Pulmonary system CT
C2826012|T102|strict|43454-8|LNC|Pulmonary system MRI|Pulmonary system MRI
C2826012|T102|strict|36803-5|LNC|Pulmonary vessels MRI angiogram|Pulmonary vessels MRI angiogram
C2826012|T102|strict|24892-2|LNC|Rectum US|Rectum US
C2826012|T102|strict|69294-7|LNC|Renal artery US|Renal artery US
C2826012|T102|strict|39435-3|LNC|Renal artery US.doppler|Renal artery US.doppler
C2826012|T102|strict|36078-4|LNC|Renal vein MRI angiogram|Renal vein MRI angiogram
C2826012|T102|strict|30868-4|LNC|Renal vessels MRI angiogram|Renal vessels MRI angiogram
C2826012|T102|strict|69295-4|LNC|Renal vessels US|Renal vessels US
C2826012|T102|strict|39426-2|LNC|Renal vessels US.doppler|Renal vessels US.doppler
C2826012|T102|strict|36804-3|LNC|Renal vessels - bilateral MRI angiogram|Renal vessels - bilateral MRI angiogram
C2826012|T102|strict|39419-7|LNC|Renal vessels - bilateral US.doppler|Renal vessels - bilateral US.doppler
C2826012|T102|strict|30619-1|LNC|Sacroiliac Joint CT|Sacroiliac Joint CT
C2826012|T102|strict|36031-3|LNC|Sacroiliac Joint MRI|Sacroiliac Joint MRI
C2826012|T102|strict|36058-6|LNC|Sacrum CT|Sacrum CT
C2826012|T102|strict|36059-4|LNC|Sacrum MRI|Sacrum MRI
C2826012|T102|strict|38053-5|LNC|Sacrum US|Sacrum US
C2826012|T102|strict|37653-3|LNC|Sacrum X-ray tomograph|Sacrum X-ray tomograph
C2826012|T102|strict|69116-2|LNC|Sacrum and Coccyx CT|Sacrum and Coccyx CT
C2826012|T102|strict|36060-2|LNC|Sacrum and Coccyx MRI|Sacrum and Coccyx MRI
C2826012|T102|strict|36933-0|LNC|Salivary gland MRI|Salivary gland MRI
C2826012|T102|strict|69298-8|LNC|Salivary gland US|Salivary gland US
C2826012|T102|strict|69117-0|LNC|Scapula CT|Scapula CT
C2826012|T102|strict|36061-0|LNC|Scapula MRI|Scapula MRI
C2826012|T102|strict|36073-5|LNC|Scrotum and Testicle MRI|Scrotum and Testicle MRI
C2826012|T102|strict|25002-7|LNC|Scrotum and Testicle US|Scrotum and Testicle US
C2826012|T102|strict|48742-1|LNC|Scrotum and Testicle US.doppler|Scrotum and Testicle US.doppler
C2826012|T102|strict|26271-7|LNC|Scrotum and Testicle - bilateral US|Scrotum and Testicle - bilateral US
C2826012|T102|strict|26272-5|LNC|Scrotum and Testicle - left US|Scrotum and Testicle - left US
C2826012|T102|strict|26273-3|LNC|Scrotum and Testicle - right US|Scrotum and Testicle - right US
C2826012|T102|strict|42437-4|LNC|Sella turcica X-ray tomograph|Sella turcica X-ray tomograph
C2826012|T102|strict|36062-8|LNC|Shoulder CT|Shoulder CT
C2826012|T102|strict|24905-2|LNC|Shoulder MRI|Shoulder MRI
C2826012|T102|strict|24907-8|LNC|Shoulder US|Shoulder US
C2826012|T102|strict|37850-5|LNC|Shoulder X-ray tomograph|Shoulder X-ray tomograph
C2826012|T102|strict|36805-0|LNC|Shoulder vessels MRI angiogram|Shoulder vessels MRI angiogram
C2826012|T102|strict|36806-8|LNC|Shoulder vessels - left MRI angiogram|Shoulder vessels - left MRI angiogram
C2826012|T102|strict|36807-6|LNC|Shoulder vessels - right MRI angiogram|Shoulder vessels - right MRI angiogram
C2826012|T102|strict|36063-6|LNC|Shoulder - bilateral CT|Shoulder - bilateral CT
C2826012|T102|strict|26266-7|LNC|Shoulder - bilateral MRI|Shoulder - bilateral MRI
C2826012|T102|strict|26265-9|LNC|Shoulder - bilateral US|Shoulder - bilateral US
C2826012|T102|strict|36064-4|LNC|Shoulder - left CT|Shoulder - left CT
C2826012|T102|strict|26268-3|LNC|Shoulder - left MRI|Shoulder - left MRI
C2826012|T102|strict|26267-5|LNC|Shoulder - left US|Shoulder - left US
C2826012|T102|strict|36065-1|LNC|Shoulder - left X-ray tomograph|Shoulder - left X-ray tomograph
C2826012|T102|strict|36066-9|LNC|Shoulder - right CT|Shoulder - right CT
C2826012|T102|strict|26270-9|LNC|Shoulder - right MRI|Shoulder - right MRI
C2826012|T102|strict|26269-1|LNC|Shoulder - right US|Shoulder - right US
C2826012|T102|strict|37811-7|LNC|Shoulder - right X-ray tomograph|Shoulder - right X-ray tomograph
C2826012|T102|strict|30588-8|LNC|Sinuses CT|Sinuses CT
C2826012|T102|strict|24914-4|LNC|Sinuses MRI|Sinuses MRI
C2826012|T102|strict|37866-1|LNC|Sinuses X-ray tomograph|Sinuses X-ray tomograph
C2826012|T102|strict|37874-5|LNC|Skull X-ray tomograph|Skull X-ray tomograph
C2826012|T102|strict|37495-9|LNC|Skull.base CT|Skull.base CT
C2826012|T102|strict|28566-8|LNC|Spine CT|Spine CT
C2826012|T102|strict|36067-7|LNC|Spine MRI|Spine MRI
C2826012|T102|strict|24926-8|LNC|Spine US|Spine US
C2826012|T102|strict|37497-5|LNC|Spine vessels MRI angiogram|Spine vessels MRI angiogram
C2826012|T102|strict|24932-6|LNC|Spine Cervical CT|Spine Cervical CT
C2826012|T102|strict|24935-9|LNC|Spine Cervical MRI|Spine Cervical MRI
C2826012|T102|strict|70926-1|LNC|Spine Cervical US|Spine Cervical US
C2826012|T102|strict|36068-5|LNC|Spine Cervical X-ray tomograph|Spine Cervical X-ray tomograph
C2826012|T102|strict|43457-1|LNC|Spine Cervical and Spine Thoracic MRI|Spine Cervical and Spine Thoracic MRI
C2826012|T102|strict|42698-1|LNC|Spine Cervical and Thoracic and Lumbar MRI|Spine Cervical and Thoracic and Lumbar MRI
C2826012|T102|strict|24963-1|LNC|Spine Lumbar CT|Spine Lumbar CT
C2826012|T102|strict|24968-0|LNC|Spine Lumbar MRI|Spine Lumbar MRI
C2826012|T102|strict|69393-7|LNC|Spine Lumbar US|Spine Lumbar US
C2826012|T102|strict|36069-3|LNC|Spine Lumbar X-ray tomograph|Spine Lumbar X-ray tomograph
C2826012|T102|strict|37232-6|LNC|Spine Lumbosacral Junction CT|Spine Lumbosacral Junction CT
C2826012|T102|strict|24978-9|LNC|Spine Thoracic CT|Spine Thoracic CT
C2826012|T102|strict|24980-5|LNC|Spine Thoracic MRI|Spine Thoracic MRI
C2826012|T102|strict|70927-9|LNC|Spine Thoracic US|Spine Thoracic US
C2826012|T102|strict|37911-5|LNC|Spine Thoracic X-ray tomograph|Spine Thoracic X-ray tomograph
C2826012|T102|strict|49565-5|LNC|Thoracic Spine vessels MRI angiogram|Thoracic Spine vessels MRI angiogram
C2826012|T102|strict|24988-8|LNC|Spleen CT|Spleen CT
C2826012|T102|strict|36070-1|LNC|Spleen MRI|Spleen MRI
C2826012|T102|strict|24990-4|LNC|Spleen US|Spleen US
C2826012|T102|strict|37225-0|LNC|Sternoclavicular Joint CT|Sternoclavicular Joint CT
C2826012|T102|strict|36071-9|LNC|Sternum CT|Sternum CT
C2826012|T102|strict|36072-7|LNC|Sternum MRI|Sternum MRI
C2826012|T102|strict|37885-1|LNC|Sternum X-ray tomograph|Sternum X-ray tomograph
C2826012|T102|strict|36782-1|LNC|Subclavian artery MRI angiogram|Subclavian artery MRI angiogram
C2826012|T102|strict|38131-9|LNC|Subclavian vessels - bilateral US|Subclavian vessels - bilateral US
C2826012|T102|strict|46359-6|LNC|Superior mesenteric vessels MRI angiogram|Superior mesenteric vessels MRI angiogram
C2826012|T102|strict|44235-0|LNC|Superior mesenteric vessels US.doppler|Superior mesenteric vessels US.doppler
C2826012|T102|strict|42468-9|LNC|Surgical specimen US|Surgical specimen US
C2826012|T102|strict|38059-2|LNC|Talus CT|Talus CT
C2826012|T102|strict|36773-0|LNC|Temporal bone CT|Temporal bone CT
C2826012|T102|strict|37226-8|LNC|Temporomandibular joint CT|Temporomandibular joint CT
C2826012|T102|strict|24999-5|LNC|Temporomandibular joint MRI|Temporomandibular joint MRI
C2826012|T102|strict|30719-9|LNC|Temporomandibular joint X-ray tomograph|Temporomandibular joint X-ray tomograph
C2826012|T102|strict|37228-4|LNC|Temporomandibular joint - bilateral MRI|Temporomandibular joint - bilateral MRI
C2826012|T102|strict|37227-6|LNC|Temporomandibular joint - bilateral X-ray tomograph|Temporomandibular joint - bilateral X-ray tomograph
C2826012|T102|strict|37230-0|LNC|Temporomandibular joint - left MRI|Temporomandibular joint - left MRI
C2826012|T102|strict|37229-2|LNC|Temporomandibular joint - left X-ray tomograph|Temporomandibular joint - left X-ray tomograph
C2826012|T102|strict|37231-8|LNC|Temporomandibular joint - right MRI|Temporomandibular joint - right MRI
C2826012|T102|strict|37819-0|LNC|Temporomandibular joint - right X-ray tomograph|Temporomandibular joint - right X-ray tomograph
C2826012|T102|strict|39446-0|LNC|Testicle vessels US.doppler|Testicle vessels US.doppler
C2826012|T102|strict|24702-3|LNC|Thigh MRI|Thigh MRI
C2826012|T102|strict|26235-2|LNC|Thigh - bilateral MRI|Thigh - bilateral MRI
C2826012|T102|strict|26236-0|LNC|Thigh - left MRI|Thigh - left MRI
C2826012|T102|strict|26237-8|LNC|Thigh - right MRI|Thigh - right MRI
C2826012|T102|strict|36054-5|LNC|Thoracic outlet CT|Thoracic outlet CT
C2826012|T102|strict|24582-9|LNC|Thoracic outlet MRI|Thoracic outlet MRI
C2826012|T102|strict|44163-4|LNC|Thoracic outlet US|Thoracic outlet US
C2826012|T102|strict|26211-3|LNC|Thoracic outlet - bilateral MRI|Thoracic outlet - bilateral MRI
C2826012|T102|strict|26212-1|LNC|Thoracic outlet - left MRI|Thoracic outlet - left MRI
C2826012|T102|strict|26213-9|LNC|Thoracic outlet - right MRI|Thoracic outlet - right MRI
C2826012|T102|strict|43507-3|LNC|Thymus gland MRI|Thymus gland MRI
C2826012|T102|strict|42300-4|LNC|Thyroid MRI|Thyroid MRI
C2826012|T102|strict|25010-0|LNC|Thyroid US|Thyroid US
C2826012|T102|strict|37898-4|LNC|Tibia and Fibula X-ray tomograph|Tibia and Fibula X-ray tomograph
C2826012|T102|strict|30888-2|LNC|Tibioperoneal vessels MRI angiogram|Tibioperoneal vessels MRI angiogram
C2826012|T102|strict|36780-5|LNC|Toe MRI|Toe MRI
C2826012|T102|strict|69285-5|LNC|Umbilical artery US.doppler|Umbilical artery US.doppler
C2826012|T102|strict|39508-7|LNC|Umbilical vessels US.doppler|Umbilical vessels US.doppler
C2826012|T102|strict|36023-0|LNC|Upper arm CT|Upper arm CT
C2826012|T102|strict|36025-5|LNC|Upper arm MRI|Upper arm MRI
C2826012|T102|strict|36026-3|LNC|Upper arm - bilateral CT|Upper arm - bilateral CT
C2826012|T102|strict|69180-8|LNC|Upper arm - bilateral MRI|Upper arm - bilateral MRI
C2826012|T102|strict|36027-1|LNC|Upper arm - left CT|Upper arm - left CT
C2826012|T102|strict|36028-9|LNC|Upper arm - left MRI|Upper arm - left MRI
C2826012|T102|strict|36029-7|LNC|Upper arm - right CT|Upper arm - right CT
C2826012|T102|strict|36030-5|LNC|Upper arm - right MRI|Upper arm - right MRI
C2826012|T102|strict|35981-0|LNC|Upper extremity CT|Upper extremity CT
C2826012|T102|strict|24688-4|LNC|Upper extremity MRI|Upper extremity MRI
C2826012|T102|strict|30710-8|LNC|Upper extremity US|Upper extremity US
C2826012|T102|strict|37923-0|LNC|Upper extremity X-ray tomograph|Upper extremity X-ray tomograph
C2826012|T102|strict|48448-5|LNC|Upper extremity artery US|Upper extremity artery US
C2826012|T102|strict|39447-8|LNC|Upper extremity artery US.doppler|Upper extremity artery US.doppler
C2826012|T102|strict|38014-7|LNC|Upper extremity artery - bilateral US|Upper extremity artery - bilateral US
C2826012|T102|strict|39423-9|LNC|Upper extremity artery - bilateral US.doppler|Upper extremity artery - bilateral US.doppler
C2826012|T102|strict|41833-5|LNC|Upper extremity artery - left US|Upper extremity artery - left US
C2826012|T102|strict|39500-4|LNC|Upper extremity artery - left US.doppler|Upper extremity artery - left US.doppler
C2826012|T102|strict|41814-5|LNC|Upper extremity artery - right US|Upper extremity artery - right US
C2826012|T102|strict|39506-1|LNC|Upper extremity artery - right US.doppler|Upper extremity artery - right US.doppler
C2826012|T102|strict|30882-5|LNC|Upper extremity vein US.doppler|Upper extremity vein US.doppler
C2826012|T102|strict|48690-2|LNC|Upper extremity vein - bilateral US|Upper extremity vein - bilateral US
C2826012|T102|strict|39496-5|LNC|Upper extremity vein - bilateral US.doppler|Upper extremity vein - bilateral US.doppler
C2826012|T102|strict|48689-4|LNC|Upper extremity vein - left US|Upper extremity vein - left US
C2826012|T102|strict|39501-2|LNC|Upper extremity vein - left US.doppler|Upper extremity vein - left US.doppler
C2826012|T102|strict|48688-6|LNC|Upper extremity vein - right US|Upper extremity vein - right US
C2826012|T102|strict|39507-9|LNC|Upper extremity vein - right US.doppler|Upper extremity vein - right US.doppler
C2826012|T102|strict|36080-0|LNC|Upper extremity veins MRI angiogram|Upper extremity veins MRI angiogram
C2826012|T102|strict|69395-2|LNC|Upper extremity veins US|Upper extremity veins US
C2826012|T102|strict|36786-2|LNC|Upper extremity veins - left MRI angiogram|Upper extremity veins - left MRI angiogram
C2826012|T102|strict|36787-0|LNC|Upper extremity veins - right MRI angiogram|Upper extremity veins - right MRI angiogram
C2826012|T102|strict|46385-1|LNC|Upper extremity vessel graft US.doppler|Upper extremity vessel graft US.doppler
C2826012|T102|strict|44236-8|LNC|Upper extremity vessel graft - bilateral US.doppler|Upper extremity vessel graft - bilateral US.doppler
C2826012|T102|strict|42475-4|LNC|Upper extremity vessel graft - left US.doppler|Upper extremity vessel graft - left US.doppler
C2826012|T102|strict|42476-2|LNC|Upper extremity vessel graft - right US.doppler|Upper extremity vessel graft - right US.doppler
C2826012|T102|strict|36084-2|LNC|Upper extremity vessels MRI angiogram|Upper extremity vessels MRI angiogram
C2826012|T102|strict|39448-6|LNC|Upper extremity vessels US.doppler|Upper extremity vessels US.doppler
C2826012|T102|strict|46379-4|LNC|Upper extremity vessels - bilateral US.doppler|Upper extremity vessels - bilateral US.doppler
C2826012|T102|strict|36797-9|LNC|Upper extremity vessels - left MRI angiogram|Upper extremity vessels - left MRI angiogram
C2826012|T102|strict|39433-8|LNC|Upper extremity vessels - left US.doppler|Upper extremity vessels - left US.doppler
C2826012|T102|strict|36798-7|LNC|Upper extremity vessels - right MRI angiogram|Upper extremity vessels - right MRI angiogram
C2826012|T102|strict|39444-5|LNC|Upper extremity vessels - right US.doppler|Upper extremity vessels - right US.doppler
C2826012|T102|strict|26232-9|LNC|Upper extremity - bilateral MRI|Upper extremity - bilateral MRI
C2826012|T102|strict|30875-9|LNC|Upper extremity .joint MRI|Upper extremity .joint MRI
C2826012|T102|strict|36774-8|LNC|Upper extremity joint - left MRI|Upper extremity joint - left MRI
C2826012|T102|strict|36775-5|LNC|Upper extremity joint - right MRI|Upper extremity joint - right MRI
C2826012|T102|strict|35982-8|LNC|Upper extremity - left CT|Upper extremity - left CT
C2826012|T102|strict|26233-7|LNC|Upper extremity - left MRI|Upper extremity - left MRI
C2826012|T102|strict|38041-0|LNC|Upper extremity - left US|Upper extremity - left US
C2826012|T102|strict|35983-6|LNC|Upper extremity - right CT|Upper extremity - right CT
C2826012|T102|strict|26234-5|LNC|Upper extremity - right MRI|Upper extremity - right MRI
C2826012|T102|strict|38052-7|LNC|Upper extremity - right US|Upper extremity - right US
C2826012|T102|strict|25019-1|LNC|Urinary bladder US|Urinary bladder US
C2826012|T102|strict|42301-2|LNC|Uterus MRI|Uterus MRI
C2826012|T102|strict|30705-8|LNC|Uterus and Fallopian tubes US|Uterus and Fallopian tubes US
C2826012|T102|strict|39036-9|LNC|Vein US|Vein US
C2826012|T102|strict|39525-1|LNC|Vein US.doppler|Vein US.doppler
C2826012|T102|strict|39030-2|LNC|Vein - bilateral US|Vein - bilateral US
C2826012|T102|strict|36783-9|LNC|Veins MRI angiogram|Veins MRI angiogram
C2826012|T102|strict|69222-8|LNC|Vena cava MRI|Vena cava MRI
C2826012|T102|strict|36081-8|LNC|Vena cava MRI angiogram|Vena cava MRI angiogram
C2826012|T102|strict|36083-4|LNC|Inferior vena cava MRI|Inferior vena cava MRI
C2826012|T102|strict|36082-6|LNC|Inferior vena cava MRI angiogram|Inferior vena cava MRI angiogram
C2826012|T102|strict|36790-4|LNC|Vena cava.inferior and Lower extremity veins MRI angiogram|Vena cava.inferior and Lower extremity veins MRI angiogram
C2826012|T102|strict|39445-2|LNC|Vessels US.doppler|Vessels US.doppler
C2826012|T102|strict|38054-3|LNC|Visceral artery US|Visceral artery US
C2826012|T102|strict|37428-0|LNC|Wrist CT|Wrist CT
C2826012|T102|strict|25033-2|LNC|Wrist MRI|Wrist MRI
C2826012|T102|strict|25036-5|LNC|Wrist US|Wrist US
C2826012|T102|strict|37932-1|LNC|Wrist X-ray tomograph|Wrist X-ray tomograph
C2826012|T102|strict|37430-6|LNC|Wrist - bilateral CT|Wrist - bilateral CT
C2826012|T102|strict|26277-4|LNC|Wrist - bilateral MRI|Wrist - bilateral MRI
C2826012|T102|strict|26278-2|LNC|Wrist - bilateral US|Wrist - bilateral US
C2826012|T102|strict|37429-8|LNC|Wrist - bilateral X-ray tomograph|Wrist - bilateral X-ray tomograph
C2826012|T102|strict|37431-4|LNC|Wrist - left CT|Wrist - left CT
C2826012|T102|strict|26279-0|LNC|Wrist - left MRI|Wrist - left MRI
C2826012|T102|strict|26280-8|LNC|Wrist - left US|Wrist - left US
C2826012|T102|strict|37432-2|LNC|Wrist - left X-ray tomograph|Wrist - left X-ray tomograph
C2826012|T102|strict|69209-5|LNC|Wrist - left and Hand - left MRI|Wrist - left and Hand - left MRI
C2826012|T102|strict|37433-0|LNC|Wrist - right CT|Wrist - right CT
C2826012|T102|strict|26281-6|LNC|Wrist - right MRI|Wrist - right MRI
C2826012|T102|strict|26282-4|LNC|Wrist - right US|Wrist - right US
C2826012|T102|strict|37644-2|LNC|Wrist - right X-ray tomograph|Wrist - right X-ray tomograph
C2826012|T102|strict|69219-4|LNC|Wrist - right and Hand - right MRI|Wrist - right and Hand - right MRI
C2826012|T102|strict|36008-1|LNC|Wrist and Hand MRI|Wrist and Hand MRI
C2826012|T102|strict|25045-6|LNC|Unspecified body region CT|Unspecified body region CT
C2826012|T102|strict|25040-7|LNC|Unspecified body region CT 3D|Unspecified body region CT 3D
C2826012|T102|strict|25056-3|LNC|Unspecified body region MRI|Unspecified body region MRI
C2826012|T102|strict|44136-0|LNC|Unspecified body region PET|Unspecified body region PET
C2826012|T102|strict|25061-3|LNC|Unspecified body region US|Unspecified body region US
C2826012|T102|strict|25071-2|LNC|Unspecified body region X-ray tomograph|Unspecified body region X-ray tomograph
C2826012|T102|strict|46375-2|LNC|Artery US|Artery US
C2826012|T102|strict|39523-6|LNC|Artery US.doppler|Artery US.doppler
C2826012|T102|strict|44229-3|LNC|Bones CT|Bones CT
C2826012|T102|strict|28576-7|LNC|Joint MRI|Joint MRI
C2826012|T102|strict|39453-6|LNC|Tendon US|Tendon US
C2826012|T102|strict|36957-9|LNC|Facial bones and Maxilla CT and 3D reconstruction|Facial bones and Maxilla CT and 3D reconstruction
C2826012|T102|strict|37294-6|LNC|Head CT and 3D reconstruction|Head CT and 3D reconstruction
C2826012|T102|strict|41804-6|LNC|Unspecified body region CT and 3D reconstruction|Unspecified body region CT and 3D reconstruction
C2826012|T102|strict|39043-5|LNC|Unspecified body region MRI and 3D reconstruction|Unspecified body region MRI and 3D reconstruction
C2826012|T102|strict|44165-9|LNC|Unspecified body region US and 3D reconstruction|Unspecified body region US and 3D reconstruction
C2826012|T102|strict|58745-1|LNC|Coronary arteries CT angiogram and 3D reconstruction W contrast IV|Coronary arteries CT angiogram and 3D reconstruction W contrast IV
C2826012|T102|strict|59255-0|LNC|Left atrium and Pulmonary veins CT angiogram and 3D reconstruction W contrast IV|Left atrium and Pulmonary veins CT angiogram and 3D reconstruction W contrast IV
C2826012|T102|strict|69082-6|LNC|Head CT and 3D reconstruction WO contrast|Head CT and 3D reconstruction WO contrast
C2826012|T102|strict|37295-3|LNC|Femur and Hip CT and anteversion measurement|Femur and Hip CT and anteversion measurement
C2826012|T102|strict|72830-3|LNC|Extremity arteries - bilateral US.doppler Multisection and physiologic artery study|Extremity arteries - bilateral US.doppler Multisection and physiologic artery study
C2826012|T102|strict|72832-9|LNC|Extremity arteries - bilateral US.doppler Multisection and physiologic artery study at rest and with exercise|Extremity arteries - bilateral US.doppler Multisection and physiologic artery study at rest and with exercise
C2826012|T102|strict|39879-2|LNC|Bone SPECT 1 phase|Bone SPECT 1 phase
C2826012|T102|strict|39881-8|LNC|Bone SPECT 3 phase whole body|Bone SPECT 3 phase whole body
C2826012|T102|strict|30760-3|LNC|Kidney - bilateral X-ray tomograph 3 views W contrast IV|Kidney - bilateral X-ray tomograph 3 views W contrast IV
C2826012|T102|strict|25055-5|LNC|Unspecified body region MRI additional sequence|Unspecified body region MRI additional sequence
C2826012|T102|strict|39408-0|LNC|Spine Thoracic X-ray tomograph AP|Spine Thoracic X-ray tomograph AP
C2826012|T102|strict|39862-8|LNC|Heart SPECT blood pool at rest and W radionuclide IV|Heart SPECT blood pool at rest and W radionuclide IV
C2826012|T102|strict|47378-5|LNC|Liver SPECT blood pool|Liver SPECT blood pool
C2826012|T102|strict|37435-5|LNC|Temporomandibular joint MRI cine|Temporomandibular joint MRI cine
C2826012|T102|strict|42693-2|LNC|Urinary Bladder and Urethra MRI cine|Urinary Bladder and Urethra MRI cine
C2826012|T102|strict|39140-9|LNC|Heart MRI cine for blood flow velocity mapping|Heart MRI cine for blood flow velocity mapping
C2826012|T102|strict|44126-1|LNC|Heart MRI cine for blood flow velocity mapping W contrast IV|Heart MRI cine for blood flow velocity mapping W contrast IV
C2826012|T102|strict|42386-3|LNC|Brain MRI cine for CSF flow|Brain MRI cine for CSF flow
C2826012|T102|strict|42387-1|LNC|Unspecified body region MRI cine for CSF flow|Unspecified body region MRI cine for CSF flow
C2826012|T102|strict|37434-8|LNC|Heart MRI cine for function|Heart MRI cine for function
C2826012|T102|strict|46300-0|LNC|Sinuses CT coronal|Sinuses CT coronal
C2826012|T102|strict|72139-9|LNC|Breast - bilateral FFD mammogram-tomosynthesis diagnostic|Breast - bilateral FFD mammogram-tomosynthesis diagnostic
C2826012|T102|strict|72138-1|LNC|Breast - left FFD mammogram-tomosynthesis diagnostic|Breast - left FFD mammogram-tomosynthesis diagnostic
C2826012|T102|strict|72137-3|LNC|Breast - right FFD mammogram-tomosynthesis diagnostic|Breast - right FFD mammogram-tomosynthesis diagnostic
C2826012|T102|strict|37436-3|LNC|Brain MRI diffusion weighted|Brain MRI diffusion weighted
C2826012|T102|strict|43555-2|LNC|Ankle - left MRI dynamic W contrast IV|Ankle - left MRI dynamic W contrast IV
C2826012|T102|strict|43449-8|LNC|Ankle - right MRI dynamic W contrast IV|Ankle - right MRI dynamic W contrast IV
C2826012|T102|strict|37437-1|LNC|Breast MRI dynamic W contrast IV|Breast MRI dynamic W contrast IV
C2826012|T102|strict|36114-7|LNC|Breast - bilateral MRI dynamic W contrast IV|Breast - bilateral MRI dynamic W contrast IV
C2826012|T102|strict|43450-6|LNC|Elbow - left MRI dynamic W contrast IV|Elbow - left MRI dynamic W contrast IV
C2826012|T102|strict|43451-4|LNC|Elbow - right MRI dynamic W contrast IV|Elbow - right MRI dynamic W contrast IV
C2826012|T102|strict|46394-3|LNC|Head CT dynamic W contrast IV|Head CT dynamic W contrast IV
C2826012|T102|strict|43452-2|LNC|Knee - left MRI dynamic W contrast IV|Knee - left MRI dynamic W contrast IV
C2826012|T102|strict|43453-0|LNC|Knee - right MRI dynamic W contrast IV|Knee - right MRI dynamic W contrast IV
C2826012|T102|strict|37438-9|LNC|Pituitary and Sella turcica CT dynamic W contrast IV|Pituitary and Sella turcica CT dynamic W contrast IV
C2826012|T102|strict|43527-1|LNC|Unspecified body region CT dynamic W contrast IV|Unspecified body region CT dynamic W contrast IV
C2826012|T102|strict|39637-4|LNC|Brain SPECT flow|Brain SPECT flow
C2826012|T102|strict|43655-0|LNC|Liver SPECT flow|Liver SPECT flow
C2826012|T102|strict|43652-7|LNC|Liver and Spleen SPECT flow|Liver and Spleen SPECT flow
C2826012|T102|strict|69235-0|LNC|Scrotum and Testicle SPECT flow|Scrotum and Testicle SPECT flow
C2826012|T102|strict|43670-9|LNC|Spleen SPECT flow|Spleen SPECT flow
C2826012|T102|strict|43673-3|LNC|Thyroid SPECT flow|Thyroid SPECT flow
C2826012|T102|strict|43662-6|LNC|Renal vessels SPECT flow W Tc-99m glucoheptonate IV|Renal vessels SPECT flow W Tc-99m glucoheptonate IV
C2826012|T102|strict|39684-6|LNC|SPECT for abscess W GA-67 IV|SPECT for abscess W GA-67 IV
C2826012|T102|strict|39811-5|LNC|SPECT for abscess|SPECT for abscess
C2826012|T102|strict|39141-7|LNC|Bone marrow MRI for blood flow|Bone marrow MRI for blood flow
C2826012|T102|strict|39656-4|LNC|Heart SPECT for infarct|Heart SPECT for infarct
C2826012|T102|strict|39654-9|LNC|Heart SPECT for infarct W Tc-99m PYP IV|Heart SPECT for infarct W Tc-99m PYP IV
C2826012|T102|strict|39655-6|LNC|Heart SPECT for infarct W Tc-99m Sestamibi IV|Heart SPECT for infarct W Tc-99m Sestamibi IV
C2826012|T102|strict|39675-4|LNC|SPECT for infection W GA-67 IV|SPECT for infection W GA-67 IV
C2826012|T102|strict|11525-3|LNC|US Pelvis and Fetus for pregnancy|US Pelvis and Fetus for pregnancy
C2826012|T102|strict|72251-2|LNC|Chest vessels CT Multisection for pulmonary embolus|Chest vessels CT Multisection for pulmonary embolus
C2826012|T102|strict|24889-8|LNC|Pylorus US for pyloric stenosis|Pylorus US for pyloric stenosis
C2826012|T102|strict|36934-8|LNC|Heart CT for scoring|Heart CT for scoring
C2826012|T102|strict|36935-5|LNC|Heart CT for scoring W contrast IV|Heart CT for scoring W contrast IV
C2826012|T102|strict|43446-4|LNC|CT for tumor whole body|CT for tumor whole body
C2826012|T102|strict|69237-6|LNC|SPECT for tumor whole body|SPECT for tumor whole body
C2826012|T102|strict|39678-8|LNC|SPECT for tumor W GA-67 IV|SPECT for tumor W GA-67 IV
C2826012|T102|strict|39748-9|LNC|SPECT for tumor W Tc-99m Sestamibi IV|SPECT for tumor W Tc-99m Sestamibi IV
C2826012|T102|strict|42292-3|LNC|SPECT for tumor W Tl-201 IV|SPECT for tumor W Tl-201 IV
C2826012|T102|strict|46395-0|LNC|Heart SPECT gated and ejection fraction at rest and W stress and W radionuclide IV|Heart SPECT gated and ejection fraction at rest and W stress and W radionuclide IV
C2826012|T102|strict|39913-9|LNC|Heart SPECT gated and ejection fraction|Heart SPECT gated and ejection fraction
C2826012|T102|strict|39918-8|LNC|Heart SPECT gated and wall motion|Heart SPECT gated and wall motion
C2826012|T102|strict|46396-8|LNC|Heart SPECT gated at rest and W Tc-99m Sestamibi IV|Heart SPECT gated at rest and W Tc-99m Sestamibi IV
C2826012|T102|strict|39916-2|LNC|Heart SPECT gated|Heart SPECT gated
C2826012|T102|strict|39930-3|LNC|Heart SPECT gated W stress and W radionuclide IV|Heart SPECT gated W stress and W radionuclide IV
C2826012|T102|strict|37439-7|LNC|Chest CT high resolution|Chest CT high resolution
C2826012|T102|strict|37440-5|LNC|Chest CT high resolution W contrast IV|Chest CT high resolution W contrast IV
C2826012|T102|strict|37441-3|LNC|Chest CT high resolution WO contrast|Chest CT high resolution WO contrast
C2826012|T102|strict|39409-8|LNC|Spine Thoracic X-ray tomograph lateral|Spine Thoracic X-ray tomograph lateral
C2826012|T102|strict|36086-7|LNC|Abdomen CT limited|Abdomen CT limited
C2826012|T102|strict|30704-1|LNC|Abdomen US limited|Abdomen US limited
C2826012|T102|strict|38047-7|LNC|Abdomen retroperitoneum US limited|Abdomen retroperitoneum US limited
C2826012|T102|strict|43572-7|LNC|Abdominal vessels US.doppler limited|Abdominal vessels US.doppler limited
C2826012|T102|strict|38011-3|LNC|Aorta US limited|Aorta US limited
C2826012|T102|strict|69280-6|LNC|Bladder US limited|Bladder US limited
C2826012|T102|strict|24599-3|LNC|Breast US limited|Breast US limited
C2826012|T102|strict|26286-5|LNC|Breast - bilateral US limited|Breast - bilateral US limited
C2826012|T102|strict|26288-1|LNC|Breast - left US limited|Breast - left US limited
C2826012|T102|strict|26290-7|LNC|Breast - right US limited|Breast - right US limited
C2826012|T102|strict|38015-4|LNC|Carotid artery US limited|Carotid artery US limited
C2826012|T102|strict|42149-5|LNC|Carotid artery - left US limited|Carotid artery - left US limited
C2826012|T102|strict|42151-1|LNC|Carotid artery - right US limited|Carotid artery - right US limited
C2826012|T102|strict|36089-1|LNC|Chest CT limited|Chest CT limited
C2826012|T102|strict|69281-4|LNC|Chest US limited|Chest US limited
C2826012|T102|strict|36090-9|LNC|Extremity CT limited|Extremity CT limited
C2826012|T102|strict|39526-9|LNC|Extremity US limited|Extremity US limited
C2826012|T102|strict|46301-8|LNC|Extremity vein - bilateral US.doppler limited|Extremity vein - bilateral US.doppler limited
C2826012|T102|strict|39424-7|LNC|Extremity vessels US.doppler limited|Extremity vessels US.doppler limited
C2826012|T102|strict|62451-0|LNC|Extremity - left US limited|Extremity - left US limited
C2826012|T102|strict|62452-8|LNC|Extremity - right US limited|Extremity - right US limited
C2826012|T102|strict|69286-3|LNC|Eye US limited|Eye US limited
C2826012|T102|strict|36937-1|LNC|Facial bones and Maxilla CT limited|Facial bones and Maxilla CT limited
C2826012|T102|strict|38020-4|LNC|Gallbladder US limited|Gallbladder US limited
C2826012|T102|strict|36087-5|LNC|Head CT limited|Head CT limited
C2826012|T102|strict|38034-5|LNC|Head US limited|Head US limited
C2826012|T102|strict|36808-4|LNC|Head vessels MRI angiogram limited|Head vessels MRI angiogram limited
C2826012|T102|strict|39044-3|LNC|Head vessels US.doppler limited|Head vessels US.doppler limited
C2826012|T102|strict|36091-7|LNC|Heart MRI limited|Heart MRI limited
C2826012|T102|strict|42707-0|LNC|Heart US limited|Heart US limited
C2826012|T102|strict|36092-5|LNC|Hip CT limited|Hip CT limited
C2826012|T102|strict|43776-4|LNC|Iliac artery US.doppler limited|Iliac artery US.doppler limited
C2826012|T102|strict|42150-3|LNC|Iliac graft US.doppler limited|Iliac graft US.doppler limited
C2826012|T102|strict|36088-3|LNC|Internal auditory canal MRI limited|Internal auditory canal MRI limited
C2826012|T102|strict|38035-2|LNC|Kidney US limited|Kidney US limited
C2826012|T102|strict|69300-2|LNC|Kidney transplant US limited|Kidney transplant US limited
C2826012|T102|strict|41812-9|LNC|Lower extremity artery US limited|Lower extremity artery US limited
C2826012|T102|strict|38042-8|LNC|Lower extremity artery US.doppler limited|Lower extremity artery US.doppler limited
C2826012|T102|strict|39430-4|LNC|Lower extremity vessels - left US.doppler limited|Lower extremity vessels - left US.doppler limited
C2826012|T102|strict|39441-1|LNC|Lower extremity vessels - right US.doppler limited|Lower extremity vessels - right US.doppler limited
C2826012|T102|strict|36093-3|LNC|Lower Extremity Joint MRI limited|Lower Extremity Joint MRI limited
C2826012|T102|strict|38039-4|LNC|Lower extremity - left US limited|Lower extremity - left US limited
C2826012|T102|strict|38050-1|LNC|Lower extremity - right US limited|Lower extremity - right US limited
C2826012|T102|strict|44116-2|LNC|Mandible CT limited|Mandible CT limited
C2826012|T102|strict|48461-8|LNC|Neck MRI limited|Neck MRI limited
C2826012|T102|strict|69212-9|LNC|Pelvis MRI limited|Pelvis MRI limited
C2826012|T102|strict|38046-9|LNC|Pelvis US limited|Pelvis US limited
C2826012|T102|strict|42152-9|LNC|Pelvis vessels US.doppler limited|Pelvis vessels US.doppler limited
C2826012|T102|strict|44173-3|LNC|Peripheral artery US limited|Peripheral artery US limited
C2826012|T102|strict|39436-1|LNC|Renal vessels US.doppler limited|Renal vessels US.doppler limited
C2826012|T102|strict|69299-6|LNC|Scrotum and Testicle US limited|Scrotum and Testicle US limited
C2826012|T102|strict|24913-6|LNC|Sinuses CT limited|Sinuses CT limited
C2826012|T102|strict|41813-7|LNC|Upper extremity artery US limited|Upper extremity artery US limited
C2826012|T102|strict|38143-4|LNC|Upper extremity artery US.doppler limited|Upper extremity artery US.doppler limited
C2826012|T102|strict|46302-6|LNC|Upper extremity artery - bilateral US.doppler limited|Upper extremity artery - bilateral US.doppler limited
C2826012|T102|strict|44237-6|LNC|Upper extremity vessel graft - bilateral US.doppler limited|Upper extremity vessel graft - bilateral US.doppler limited
C2826012|T102|strict|46303-4|LNC|Upper extremity vessels US.doppler limited|Upper extremity vessels US.doppler limited
C2826012|T102|strict|36094-1|LNC|Upper extremity .joint MRI limited|Upper extremity .joint MRI limited
C2826012|T102|strict|39045-0|LNC|Vein US limited|Vein US limited
C2826012|T102|strict|39524-4|LNC|Vein US.doppler limited|Vein US.doppler limited
C2826012|T102|strict|25039-9|LNC|Unspecified body region CT limited|Unspecified body region CT limited
C2826012|T102|strict|48460-0|LNC|Unspecified body region MRI limited|Unspecified body region MRI limited
C2826012|T102|strict|69282-2|LNC|Unspecified body region US.doppler limited|Unspecified body region US.doppler limited
C2826012|T102|strict|72831-1|LNC|Extremity arteries - bilateral US.doppler Multisection limited and physiologic artery study|Extremity arteries - bilateral US.doppler Multisection limited and physiologic artery study
C2826012|T102|strict|44127-9|LNC|Heart MRI limited cine for function|Heart MRI limited cine for function
C2826012|T102|strict|39046-8|LNC|Pelvis CT limited pelvimetry WO contrast|Pelvis CT limited pelvimetry WO contrast
C2826012|T102|strict|36102-2|LNC|Abdomen CT limited W and WO contrast IV|Abdomen CT limited W and WO contrast IV
C2826012|T102|strict|36095-8|LNC|Abdomen CT limited W contrast IV|Abdomen CT limited W contrast IV
C2826012|T102|strict|36096-6|LNC|Brain MRI limited W contrast IV|Brain MRI limited W contrast IV
C2826012|T102|strict|69096-6|LNC|Chest CT limited W contrast IV|Chest CT limited W contrast IV
C2826012|T102|strict|36098-2|LNC|Pelvis CT limited W contrast IV|Pelvis CT limited W contrast IV
C2826012|T102|strict|36099-0|LNC|Spine Cervical CT limited W contrast IV|Spine Cervical CT limited W contrast IV
C2826012|T102|strict|36100-6|LNC|Spine Lumbar MRI limited W contrast IV|Spine Lumbar MRI limited W contrast IV
C2826012|T102|strict|36101-4|LNC|Spine Thoracic MRI limited W contrast IV|Spine Thoracic MRI limited W contrast IV
C2826012|T102|strict|36097-4|LNC|Upper extremity CT limited W contrast IV|Upper extremity CT limited W contrast IV
C2826012|T102|strict|39681-2|LNC|SPECT limited W GA-67 IV|SPECT limited W GA-67 IV
C2826012|T102|strict|39813-1|LNC|Bone SPECT limited|Bone SPECT limited
C2826012|T102|strict|39821-4|LNC|Bone marrow SPECT limited|Bone marrow SPECT limited
C2826012|T102|strict|36103-0|LNC|Abdomen CT limited WO contrast|Abdomen CT limited WO contrast
C2826012|T102|strict|36105-5|LNC|Brain MRI limited WO contrast|Brain MRI limited WO contrast
C2826012|T102|strict|47366-0|LNC|Chest CT limited WO contrast|Chest CT limited WO contrast
C2826012|T102|strict|36938-9|LNC|Facial bones and Maxilla CT limited WO contrast|Facial bones and Maxilla CT limited WO contrast
C2826012|T102|strict|36104-8|LNC|Head CT limited WO contrast|Head CT limited WO contrast
C2826012|T102|strict|36106-3|LNC|Lower extremity CT limited WO contrast|Lower extremity CT limited WO contrast
C2826012|T102|strict|36107-1|LNC|Lower extremity joint - left MRI limited WO contrast|Lower extremity joint - left MRI limited WO contrast
C2826012|T102|strict|38769-6|LNC|Lower extremity joint - right MRI limited WO contrast|Lower extremity joint - right MRI limited WO contrast
C2826012|T102|strict|36108-9|LNC|Pelvis CT limited WO contrast|Pelvis CT limited WO contrast
C2826012|T102|strict|46304-2|LNC|Sinuses CT limited WO contrast|Sinuses CT limited WO contrast
C2826012|T102|strict|36109-7|LNC|Spine Cervical CT limited WO contrast|Spine Cervical CT limited WO contrast
C2826012|T102|strict|36110-5|LNC|Spine Lumbar CT limited WO contrast|Spine Lumbar CT limited WO contrast
C2826012|T102|strict|36111-3|LNC|Spine Lumbar MRI limited WO contrast|Spine Lumbar MRI limited WO contrast
C2826012|T102|strict|36112-1|LNC|Spine Thoracic MRI limited WO contrast|Spine Thoracic MRI limited WO contrast
C2826012|T102|strict|39905-5|LNC|Bone SPECT multiple areas|Bone SPECT multiple areas
C2826012|T102|strict|39906-3|LNC|Bone marrow SPECT multiple areas|Bone marrow SPECT multiple areas
C2826012|T102|strict|39527-7|LNC|Unspecified body region US of foreign body|Unspecified body region US of foreign body
C2826012|T102|strict|49569-7|LNC|Heart SPECT perfusion and wall motion at rest and W stress and W Tl-201 IV and W Tc-99m Sestamibi IV|Heart SPECT perfusion and wall motion at rest and W stress and W Tl-201 IV and W Tc-99m Sestamibi IV
C2826012|T102|strict|43659-2|LNC|Heart SPECT perfusion qualitative at rest and W radionuclide IV|Heart SPECT perfusion qualitative at rest and W radionuclide IV
C2826012|T102|strict|39725-7|LNC|Heart SPECT perfusion at rest and W adenosine and W Tl-201 IV|Heart SPECT perfusion at rest and W adenosine and W Tl-201 IV
C2826012|T102|strict|39718-2|LNC|Heart SPECT perfusion at rest and W radionuclide IV|Heart SPECT perfusion at rest and W radionuclide IV
C2826012|T102|strict|39724-0|LNC|Heart SPECT perfusion at rest and W stress and W radionuclide IV|Heart SPECT perfusion at rest and W stress and W radionuclide IV
C2826012|T102|strict|39723-2|LNC|Heart SPECT perfusion at rest and W stress and W Tl-201 IV|Heart SPECT perfusion at rest and W stress and W Tl-201 IV
C2826012|T102|strict|49568-9|LNC|Heart SPECT perfusion at rest and W stress and W Tl-201 IV and W Tc-99m Sestamibi IV|Heart SPECT perfusion at rest and W stress and W Tl-201 IV and W Tc-99m Sestamibi IV
C2826012|T102|strict|39729-9|LNC|Heart SPECT perfusion at rest and W Tl-201 IV|Heart SPECT perfusion at rest and W Tl-201 IV
C2826012|T102|strict|39700-0|LNC|Heart SPECT perfusion W adenosine and W radionuclide IV|Heart SPECT perfusion W adenosine and W radionuclide IV
C2826012|T102|strict|49567-1|LNC|Heart SPECT perfusion W adenosine and W Tc-99m Sestamibi IV|Heart SPECT perfusion W adenosine and W Tc-99m Sestamibi IV
C2826012|T102|strict|39142-5|LNC|Head CT perfusion W contrast IV|Head CT perfusion W contrast IV
C2826012|T102|strict|39712-5|LNC|Heart SPECT perfusion|Heart SPECT perfusion
C2826012|T102|strict|39734-9|LNC|Heart SPECT perfusion W stress and W radionuclide IV|Heart SPECT perfusion W stress and W radionuclide IV
C2826012|T102|strict|39736-4|LNC|Heart SPECT perfusion W stress and W Tc-99m Sestamibi IV|Heart SPECT perfusion W stress and W Tc-99m Sestamibi IV
C2826012|T102|strict|39710-9|LNC|Heart SPECT perfusion W Tc-99m Sestamibi IV|Heart SPECT perfusion W Tc-99m Sestamibi IV
C2826012|T102|strict|39711-7|LNC|Heart SPECT perfusion W Tl-201 IV|Heart SPECT perfusion W Tl-201 IV
C2826012|T102|strict|38060-0|LNC|Spine.lumbosacral+Cervical+Thoracic MRI sagittal|Spine.lumbosacral+Cervical+Thoracic MRI sagittal
C2826012|T102|strict|25052-2|LNC|Unspecified body region CT sagittal and coronal|Unspecified body region CT sagittal and coronal
C2826012|T102|strict|25050-6|LNC|Unspecified body region CT 3D sagittal and coronal disarticulation|Unspecified body region CT 3D sagittal and coronal disarticulation
C2826012|T102|strict|42132-1|LNC|Breast US screening|Breast US screening
C2826012|T102|strict|72142-3|LNC|Breast - bilateral FFD mammogram-tomosynthesis screening|Breast - bilateral FFD mammogram-tomosynthesis screening
C2826012|T102|strict|72141-5|LNC|Breast - left FFD mammogram-tomosynthesis screening|Breast - left FFD mammogram-tomosynthesis screening
C2826012|T102|strict|72140-7|LNC|Breast - right FFD mammogram-tomosynthesis screening|Breast - right FFD mammogram-tomosynthesis screening
C2826012|T102|strict|37442-1|LNC|Brain MRI spectroscopy|Brain MRI spectroscopy
C2826012|T102|strict|37443-9|LNC|Unspecified body region MRI spectroscopy|Unspecified body region MRI spectroscopy
C2826012|T102|strict|36939-7|LNC|Spine CT stereotactic|Spine CT stereotactic
C2826012|T102|strict|70929-5|LNC|Spine Cervical CT stereotactic|Spine Cervical CT stereotactic
C2826012|T102|strict|70928-7|LNC|Spine Lumbar CT stereotactic|Spine Lumbar CT stereotactic
C2826012|T102|strict|70930-3|LNC|Spine Thoracic CT stereotactic|Spine Thoracic CT stereotactic
C2826012|T102|strict|36940-5|LNC|Unspecified body region CT stereotactic|Unspecified body region CT stereotactic
C2826012|T102|strict|42455-6|LNC|Pelvis US transabdominal and transvaginal|Pelvis US transabdominal and transvaginal
C2826012|T102|strict|24677-7|LNC|Pelvis US transvaginal|Pelvis US transvaginal
C2826012|T102|strict|42390-5|LNC|Transvaginal MRI|Transvaginal MRI
C2826012|T102|strict|39838-8|LNC|Lung SPECT ventilation and perfusion W radionuclide inhaled and W radionuclide IV|Lung SPECT ventilation and perfusion W radionuclide inhaled and W radionuclide IV
C2826012|T102|strict|39898-2|LNC|Lung SPECT ventilation W radionuclide aerosol inhaled|Lung SPECT ventilation W radionuclide aerosol inhaled
C2826012|T102|strict|39872-7|LNC|Heart SPECT wall motion|Heart SPECT wall motion
C2826012|T102|strict|46305-9|LNC|CT whole body|CT whole body
C2826012|T102|strict|46358-8|LNC|MRI whole body|MRI whole body
C2826012|T102|strict|44139-4|LNC|PET whole body|PET whole body
C2826012|T102|strict|46306-7|LNC|CT whole body W contrast IV|CT whole body W contrast IV
C2826012|T102|strict|39680-4|LNC|SPECT whole body W GA-67 IV|SPECT whole body W GA-67 IV
C2826012|T102|strict|39816-4|LNC|Bone SPECT whole body|Bone SPECT whole body
C2826012|T102|strict|39825-5|LNC|Bone marrow SPECT whole body|Bone marrow SPECT whole body
C2826012|T102|strict|41837-6|LNC|SPECT whole body W Tc-99m Arcitumomab IV|SPECT whole body W Tc-99m Arcitumomab IV
C2826012|T102|strict|39658-0|LNC|Heart SPECT at rest and W radionuclide IV|Heart SPECT at rest and W radionuclide IV
C2826012|T102|strict|39662-2|LNC|Heart SPECT at rest and W stress and W Tc-99m Sestamibi IV|Heart SPECT at rest and W stress and W Tc-99m Sestamibi IV
C2826012|T102|strict|49566-3|LNC|Heart SPECT at rest and W Tc-99m Sestamibi IV|Heart SPECT at rest and W Tc-99m Sestamibi IV
C2826012|T102|strict|30711-6|LNC|Hip US developmental joint assessment|Hip US developmental joint assessment
C2826012|T102|strict|24732-0|LNC|Head US during surgery|Head US during surgery
C2826012|T102|strict|30706-6|LNC|Liver US during surgery|Liver US during surgery
C2826012|T102|strict|30701-7|LNC|Unspecified body region US during surgery|Unspecified body region US during surgery
C2826012|T102|strict|69388-7|LNC|Urinary bladder US post void|Urinary bladder US post void
C2826012|T102|strict|69086-7|LNC|Aorta CT W and WO contrast|Aorta CT W and WO contrast
C2826012|T102|strict|69108-9|LNC|Pulmonary vessels CT angiogram W and WO contrast|Pulmonary vessels CT angiogram W and WO contrast
C2826012|T102|strict|69085-9|LNC|Renal vessels CT angiogram W and WO contrast|Renal vessels CT angiogram W and WO contrast
C2826012|T102|strict|69207-9|LNC|Hip - left MRI W and WO contrast intraarticular|Hip - left MRI W and WO contrast intraarticular
C2826012|T102|strict|69217-8|LNC|Hip - right MRI W and WO contrast intraarticular|Hip - right MRI W and WO contrast intraarticular
C2826012|T102|strict|69208-7|LNC|Shoulder - left MRI W and WO contrast intraarticular|Shoulder - left MRI W and WO contrast intraarticular
C2826012|T102|strict|69218-6|LNC|Shoulder - right MRI W and WO contrast intraarticular|Shoulder - right MRI W and WO contrast intraarticular
C2826012|T102|strict|48442-8|LNC|Spine CT W and WO contrast IT|Spine CT W and WO contrast IT
C2826012|T102|strict|48450-1|LNC|Spine Cervical MRI W and WO contrast IT|Spine Cervical MRI W and WO contrast IT
C2826012|T102|strict|44114-7|LNC|Spine Lumbar CT W and WO contrast IT|Spine Lumbar CT W and WO contrast IT
C2826012|T102|strict|48452-7|LNC|Spine Lumbar MRI W and WO contrast IT|Spine Lumbar MRI W and WO contrast IT
C2826012|T102|strict|44113-9|LNC|Spine Thoracic CT W and WO contrast IT|Spine Thoracic CT W and WO contrast IT
C2826012|T102|strict|48441-0|LNC|Spine Thoracic MRI W and WO contrast IT|Spine Thoracic MRI W and WO contrast IT
C2826012|T102|strict|36267-3|LNC|Abdomen CT W and WO contrast IV|Abdomen CT W and WO contrast IV
C2826012|T102|strict|24557-1|LNC|Abdomen MRI W and WO contrast IV|Abdomen MRI W and WO contrast IV
C2826012|T102|strict|48743-9|LNC|Abdomen retroperitoneum CT W and WO contrast IV|Abdomen retroperitoneum CT W and WO contrast IV
C2826012|T102|strict|42274-1|LNC|Abdomen and Pelvis CT W and WO contrast IV|Abdomen and Pelvis CT W and WO contrast IV
C2826012|T102|strict|36846-4|LNC|Abdominal veins MRI angiogram W and WO contrast IV|Abdominal veins MRI angiogram W and WO contrast IV
C2826012|T102|strict|30805-6|LNC|Abdominal vessels CT angiogram W and WO contrast IV|Abdominal vessels CT angiogram W and WO contrast IV
C2826012|T102|strict|36855-5|LNC|Abdominal vessels MRI angiogram W and WO contrast IV|Abdominal vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|36950-4|LNC|Adrenal gland CT W and WO contrast IV|Adrenal gland CT W and WO contrast IV
C2826012|T102|strict|36951-2|LNC|Adrenal gland MRI W and WO contrast IV|Adrenal gland MRI W and WO contrast IV
C2826012|T102|strict|36268-1|LNC|Ankle CT W and WO contrast IV|Ankle CT W and WO contrast IV
C2826012|T102|strict|24539-9|LNC|Ankle MRI W and WO contrast IV|Ankle MRI W and WO contrast IV
C2826012|T102|strict|26187-5|LNC|Ankle - bilateral MRI W and WO contrast IV|Ankle - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36269-9|LNC|Ankle - left CT W and WO contrast IV|Ankle - left CT W and WO contrast IV
C2826012|T102|strict|26188-3|LNC|Ankle - left MRI W and WO contrast IV|Ankle - left MRI W and WO contrast IV
C2826012|T102|strict|36270-7|LNC|Ankle - right CT W and WO contrast IV|Ankle - right CT W and WO contrast IV
C2826012|T102|strict|26189-1|LNC|Ankle - right MRI W and WO contrast IV|Ankle - right MRI W and WO contrast IV
C2826012|T102|strict|44131-1|LNC|Aorta MRI angiogram W and WO contrast IV|Aorta MRI angiogram W and WO contrast IV
C2826012|T102|strict|36271-5|LNC|Aorta abdominal CT W and WO contrast IV|Aorta abdominal CT W and WO contrast IV
C2826012|T102|strict|36273-1|LNC|Aorta abdominal MRI W and WO contrast IV|Aorta abdominal MRI W and WO contrast IV
C2826012|T102|strict|36272-3|LNC|Aorta abdominal MRI angiogram W and WO contrast IV|Aorta abdominal MRI angiogram W and WO contrast IV
C2826012|T102|strict|36274-9|LNC|Aorta thoracic MRI angiogram W and WO contrast IV|Aorta thoracic MRI angiogram W and WO contrast IV
C2826012|T102|strict|30806-4|LNC|Aorta and Femoral artery - bilateral CT angiogram W and WO contrast IV|Aorta and Femoral artery - bilateral CT angiogram W and WO contrast IV
C2826012|T102|strict|46360-4|LNC|Aortic arch MRI angiogram W and WO contrast IV|Aortic arch MRI angiogram W and WO contrast IV
C2826012|T102|strict|43509-9|LNC|Axilla - left MRI W and WO contrast IV|Axilla - left MRI W and WO contrast IV
C2826012|T102|strict|43511-5|LNC|Axilla - right MRI W and WO contrast IV|Axilla - right MRI W and WO contrast IV
C2826012|T102|strict|36944-7|LNC|Biliary ducts and Pancreatic duct MRI W and WO contrast IV|Biliary ducts and Pancreatic duct MRI W and WO contrast IV
C2826012|T102|strict|24587-8|LNC|Brain MRI W and WO contrast IV|Brain MRI W and WO contrast IV
C2826012|T102|strict|48694-4|LNC|Brain.temporal MRI W and WO contrast IV|Brain.temporal MRI W and WO contrast IV
C2826012|T102|strict|43769-9|LNC|Brain and Internal auditory canal MRI W and WO contrast IV|Brain and Internal auditory canal MRI W and WO contrast IV
C2826012|T102|strict|42392-1|LNC|Brain and Pituitary and Sella turcica MRI W and WO contrast IV|Brain and Pituitary and Sella turcica MRI W and WO contrast IV
C2826012|T102|strict|36276-4|LNC|Breast MRI W and WO contrast IV|Breast MRI W and WO contrast IV
C2826012|T102|strict|69189-9|LNC|Breast implant MRI W and WO contrast IV|Breast implant MRI W and WO contrast IV
C2826012|T102|strict|69166-7|LNC|Breast implant - bilateral MRI W and WO contrast IV|Breast implant - bilateral MRI W and WO contrast IV
C2826012|T102|strict|38870-2|LNC|Breast implant - left MRI W and WO contrast IV|Breast implant - left MRI W and WO contrast IV
C2826012|T102|strict|38062-6|LNC|Breast implant - right MRI W and WO contrast IV|Breast implant - right MRI W and WO contrast IV
C2826012|T102|strict|36277-2|LNC|Breast - bilateral MRI W and WO contrast IV|Breast - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36278-0|LNC|Breast - left MRI W and WO contrast IV|Breast - left MRI W and WO contrast IV
C2826012|T102|strict|36279-8|LNC|Breast - right MRI W and WO contrast IV|Breast - right MRI W and WO contrast IV
C2826012|T102|strict|43528-9|LNC|Breast - unilateral MRI W and WO contrast IV|Breast - unilateral MRI W and WO contrast IV
C2826012|T102|strict|36358-0|LNC|Calcaneus CT W and WO contrast IV|Calcaneus CT W and WO contrast IV
C2826012|T102|strict|36280-6|LNC|Calcaneus - left CT W and WO contrast IV|Calcaneus - left CT W and WO contrast IV
C2826012|T102|strict|36281-4|LNC|Calcaneus - right CT W and WO contrast IV|Calcaneus - right CT W and WO contrast IV
C2826012|T102|strict|36856-3|LNC|Carotid vessel MRI angiogram W and WO contrast IV|Carotid vessel MRI angiogram W and WO contrast IV
C2826012|T102|strict|30598-7|LNC|Chest CT W and WO contrast IV|Chest CT W and WO contrast IV
C2826012|T102|strict|36283-0|LNC|Chest MRI W and WO contrast IV|Chest MRI W and WO contrast IV
C2826012|T102|strict|36848-0|LNC|Chest veins MRI angiogram W and WO contrast IV|Chest veins MRI angiogram W and WO contrast IV
C2826012|T102|strict|30804-9|LNC|Chest vessels CT angiogram W and WO contrast IV|Chest vessels CT angiogram W and WO contrast IV
C2826012|T102|strict|36420-8|LNC|Chest vessels MRI angiogram W and WO contrast IV|Chest vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|42277-4|LNC|Chest and Abdomen CT W and WO contrast IV|Chest and Abdomen CT W and WO contrast IV
C2826012|T102|strict|36284-8|LNC|Chest and Abdomen MRI W and WO contrast IV|Chest and Abdomen MRI W and WO contrast IV
C2826012|T102|strict|72252-0|LNC|Chest and Abdomen and Pelvis CT W and WO contrast IV|Chest and Abdomen and Pelvis CT W and WO contrast IV
C2826012|T102|strict|69161-8|LNC|Circle of Willis MRI angiogram W and WO contrast IV|Circle of Willis MRI angiogram W and WO contrast IV
C2826012|T102|strict|42299-8|LNC|Clavicle MRI W and WO contrast IV|Clavicle MRI W and WO contrast IV
C2826012|T102|strict|48455-0|LNC|Clavicle - left MRI W and WO contrast IV|Clavicle - left MRI W and WO contrast IV
C2826012|T102|strict|48454-3|LNC|Clavicle - right MRI W and WO contrast IV|Clavicle - right MRI W and WO contrast IV
C2826012|T102|strict|36285-5|LNC|Elbow CT W and WO contrast IV|Elbow CT W and WO contrast IV
C2826012|T102|strict|24675-1|LNC|Elbow MRI W and WO contrast IV|Elbow MRI W and WO contrast IV
C2826012|T102|strict|26193-3|LNC|Elbow - bilateral MRI W and WO contrast IV|Elbow - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36286-3|LNC|Elbow - left CT W and WO contrast IV|Elbow - left CT W and WO contrast IV
C2826012|T102|strict|26194-1|LNC|Elbow - left MRI W and WO contrast IV|Elbow - left MRI W and WO contrast IV
C2826012|T102|strict|36287-1|LNC|Elbow - right CT W and WO contrast IV|Elbow - right CT W and WO contrast IV
C2826012|T102|strict|26195-8|LNC|Elbow - right MRI W and WO contrast IV|Elbow - right MRI W and WO contrast IV
C2826012|T102|strict|42268-3|LNC|Extremity CT W and WO contrast IV|Extremity CT W and WO contrast IV
C2826012|T102|strict|24694-2|LNC|Face MRI W and WO contrast IV|Face MRI W and WO contrast IV
C2826012|T102|strict|30803-1|LNC|Facial bones and Maxilla CT W and WO contrast IV|Facial bones and Maxilla CT W and WO contrast IV
C2826012|T102|strict|36338-2|LNC|Femur CT W and WO contrast IV|Femur CT W and WO contrast IV
C2826012|T102|strict|36339-0|LNC|Femur - left CT W and WO contrast IV|Femur - left CT W and WO contrast IV
C2826012|T102|strict|36340-8|LNC|Femur - right CT W and WO contrast IV|Femur - right CT W and WO contrast IV
C2826012|T102|strict|69194-9|LNC|Finger MRI W and WO contrast IV|Finger MRI W and WO contrast IV
C2826012|T102|strict|69204-6|LNC|Finger - left MRI W and WO contrast IV|Finger - left MRI W and WO contrast IV
C2826012|T102|strict|69214-5|LNC|Finger - right MRI W and WO contrast IV|Finger - right MRI W and WO contrast IV
C2826012|T102|strict|36341-6|LNC|Foot CT W and WO contrast IV|Foot CT W and WO contrast IV
C2826012|T102|strict|30682-9|LNC|Foot MRI W and WO contrast IV|Foot MRI W and WO contrast IV
C2826012|T102|strict|36342-4|LNC|Foot - bilateral MRI W and WO contrast IV|Foot - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36343-2|LNC|Foot - left CT W and WO contrast IV|Foot - left CT W and WO contrast IV
C2826012|T102|strict|36344-0|LNC|Foot - left MRI W and WO contrast IV|Foot - left MRI W and WO contrast IV
C2826012|T102|strict|36345-7|LNC|Foot - right CT W and WO contrast IV|Foot - right CT W and WO contrast IV
C2826012|T102|strict|36346-5|LNC|Foot - right MRI W and WO contrast IV|Foot - right MRI W and WO contrast IV
C2826012|T102|strict|36347-3|LNC|Forearm CT W and WO contrast IV|Forearm CT W and WO contrast IV
C2826012|T102|strict|30684-5|LNC|Forearm MRI W and WO contrast IV|Forearm MRI W and WO contrast IV
C2826012|T102|strict|69174-1|LNC|Forearm - bilateral MRI W and WO contrast IV|Forearm - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36348-1|LNC|Forearm - left CT W and WO contrast IV|Forearm - left CT W and WO contrast IV
C2826012|T102|strict|36349-9|LNC|Forearm - left MRI W and WO contrast IV|Forearm - left MRI W and WO contrast IV
C2826012|T102|strict|36350-7|LNC|Forearm - right CT W and WO contrast IV|Forearm - right CT W and WO contrast IV
C2826012|T102|strict|36351-5|LNC|Forearm - right MRI W and WO contrast IV|Forearm - right MRI W and WO contrast IV
C2826012|T102|strict|36352-3|LNC|Hand CT W and WO contrast IV|Hand CT W and WO contrast IV
C2826012|T102|strict|30686-0|LNC|Hand MRI W and WO contrast IV|Hand MRI W and WO contrast IV
C2826012|T102|strict|69177-4|LNC|Hand - bilateral MRI W and WO contrast IV|Hand - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36353-1|LNC|Hand - left CT W and WO contrast IV|Hand - left CT W and WO contrast IV
C2826012|T102|strict|36354-9|LNC|Hand - left MRI W and WO contrast IV|Hand - left MRI W and WO contrast IV
C2826012|T102|strict|36355-6|LNC|Hand - right CT W and WO contrast IV|Hand - right CT W and WO contrast IV
C2826012|T102|strict|36356-4|LNC|Hand - right MRI W and WO contrast IV|Hand - right MRI W and WO contrast IV
C2826012|T102|strict|24726-2|LNC|Head CT W and WO contrast IV|Head CT W and WO contrast IV
C2826012|T102|strict|24729-6|LNC|Head CT cine W and WO contrast IV|Head CT cine W and WO contrast IV
C2826012|T102|strict|36847-2|LNC|Head veins MRI angiogram W and WO contrast IV|Head veins MRI angiogram W and WO contrast IV
C2826012|T102|strict|30593-8|LNC|Head vessels CT angiogram W and WO contrast IV|Head vessels CT angiogram W and WO contrast IV
C2826012|T102|strict|36857-1|LNC|Head vessels MRI angiogram W and WO contrast IV|Head vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|36357-2|LNC|Heart MRI W and WO contrast IV|Heart MRI W and WO contrast IV
C2826012|T102|strict|36359-8|LNC|Hip CT W and WO contrast IV|Hip CT W and WO contrast IV
C2826012|T102|strict|30688-6|LNC|Hip MRI W and WO contrast IV|Hip MRI W and WO contrast IV
C2826012|T102|strict|36360-6|LNC|Hip - bilateral CT W and WO contrast IV|Hip - bilateral CT W and WO contrast IV
C2826012|T102|strict|36361-4|LNC|Hip - bilateral MRI W and WO contrast IV|Hip - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36362-2|LNC|Hip - left CT W and WO contrast IV|Hip - left CT W and WO contrast IV
C2826012|T102|strict|36363-0|LNC|Hip - left MRI W and WO contrast IV|Hip - left MRI W and WO contrast IV
C2826012|T102|strict|36364-8|LNC|Hip - right CT W and WO contrast IV|Hip - right CT W and WO contrast IV
C2826012|T102|strict|36365-5|LNC|Hip - right MRI W and WO contrast IV|Hip - right MRI W and WO contrast IV
C2826012|T102|strict|36282-2|LNC|Internal auditory canal CT W and WO contrast IV|Internal auditory canal CT W and WO contrast IV
C2826012|T102|strict|30659-7|LNC|Internal auditory canal MRI W and WO contrast IV|Internal auditory canal MRI W and WO contrast IV
C2826012|T102|strict|24740-3|LNC|Internal auditory canal and Posterior fossa MRI W and WO contrast IV|Internal auditory canal and Posterior fossa MRI W and WO contrast IV
C2826012|T102|strict|43768-1|LNC|Kidney CT W and WO contrast IV|Kidney CT W and WO contrast IV
C2826012|T102|strict|43775-6|LNC|Kidney MRI W and WO contrast IV|Kidney MRI W and WO contrast IV
C2826012|T102|strict|36377-0|LNC|Kidney - bilateral CT W and WO contrast IV|Kidney - bilateral CT W and WO contrast IV
C2826012|T102|strict|36378-8|LNC|Kidney - bilateral MRI W and WO contrast IV|Kidney - bilateral MRI W and WO contrast IV
C2826012|T102|strict|24784-1|LNC|Kidney - bilateral X-ray tomograph W and WO contrast IV|Kidney - bilateral X-ray tomograph W and WO contrast IV
C2826012|T102|strict|36379-6|LNC|Knee CT W and WO contrast IV|Knee CT W and WO contrast IV
C2826012|T102|strict|24803-9|LNC|Knee MRI W and WO contrast IV|Knee MRI W and WO contrast IV
C2826012|T102|strict|38837-1|LNC|Knee vessels - left MRI angiogram W and WO contrast IV|Knee vessels - left MRI angiogram W and WO contrast IV
C2826012|T102|strict|36862-1|LNC|Knee vessels - right MRI angiogram W and WO contrast IV|Knee vessels - right MRI angiogram W and WO contrast IV
C2826012|T102|strict|26199-0|LNC|Knee - bilateral MRI W and WO contrast IV|Knee - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36380-4|LNC|Knee - left CT W and WO contrast IV|Knee - left CT W and WO contrast IV
C2826012|T102|strict|26200-6|LNC|Knee - left MRI W and WO contrast IV|Knee - left MRI W and WO contrast IV
C2826012|T102|strict|36381-2|LNC|Knee - right CT W and WO contrast IV|Knee - right CT W and WO contrast IV
C2826012|T102|strict|26201-4|LNC|Knee - right MRI W and WO contrast IV|Knee - right MRI W and WO contrast IV
C2826012|T102|strict|36382-0|LNC|Larynx MRI W and WO contrast IV|Larynx MRI W and WO contrast IV
C2826012|T102|strict|30612-6|LNC|Liver CT W and WO contrast IV|Liver CT W and WO contrast IV
C2826012|T102|strict|30670-4|LNC|Liver MRI W and WO contrast IV|Liver MRI W and WO contrast IV
C2826012|T102|strict|36288-9|LNC|Lower extremity CT W and WO contrast IV|Lower extremity CT W and WO contrast IV
C2826012|T102|strict|39291-0|LNC|Lower extremity MRI W and WO contrast IV|Lower extremity MRI W and WO contrast IV
C2826012|T102|strict|36416-6|LNC|Lower extremity veins MRI angiogram W and WO contrast IV|Lower extremity veins MRI angiogram W and WO contrast IV
C2826012|T102|strict|36849-8|LNC|Lower extremity veins - left MRI angiogram W and WO contrast IV|Lower extremity veins - left MRI angiogram W and WO contrast IV
C2826012|T102|strict|36850-6|LNC|Lower extremity veins - right MRI angiogram W and WO contrast IV|Lower extremity veins - right MRI angiogram W and WO contrast IV
C2826012|T102|strict|30807-2|LNC|Lower extremity vessels CT angiogram W and WO contrast IV|Lower extremity vessels CT angiogram W and WO contrast IV
C2826012|T102|strict|44128-7|LNC|Lower extremity vessels MRI angiogram W and WO contrast IV|Lower extremity vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|46308-3|LNC|Lower extremity vessels - left CT angiogram W and WO contrast IV|Lower extremity vessels - left CT angiogram W and WO contrast IV
C2826012|T102|strict|36858-9|LNC|Lower extremity vessels - left MRI angiogram W and WO contrast IV|Lower extremity vessels - left MRI angiogram W and WO contrast IV
C2826012|T102|strict|46307-5|LNC|Lower extremity vessels - right CT angiogram W and WO contrast IV|Lower extremity vessels - right CT angiogram W and WO contrast IV
C2826012|T102|strict|36859-7|LNC|Lower extremity vessels - right MRI angiogram W and WO contrast IV|Lower extremity vessels - right MRI angiogram W and WO contrast IV
C2826012|T102|strict|36289-7|LNC|Lower extremity - bilateral MRI W and WO contrast IV|Lower extremity - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36371-3|LNC|Lower Extremity Joint MRI W and WO contrast IV|Lower Extremity Joint MRI W and WO contrast IV
C2826012|T102|strict|36372-1|LNC|Lower extremity joint - left MRI W and WO contrast IV|Lower extremity joint - left MRI W and WO contrast IV
C2826012|T102|strict|36373-9|LNC|Lower extremity joint - right MRI W and WO contrast IV|Lower extremity joint - right MRI W and WO contrast IV
C2826012|T102|strict|36290-5|LNC|Lower extremity - left CT W and WO contrast IV|Lower extremity - left CT W and WO contrast IV
C2826012|T102|strict|36291-3|LNC|Lower extremity - left MRI W and WO contrast IV|Lower extremity - left MRI W and WO contrast IV
C2826012|T102|strict|36292-1|LNC|Lower extremity - right CT W and WO contrast IV|Lower extremity - right CT W and WO contrast IV
C2826012|T102|strict|36333-3|LNC|Lower extremity - right MRI W and WO contrast IV|Lower extremity - right MRI W and WO contrast IV
C2826012|T102|strict|36408-3|LNC|Lower leg CT W and WO contrast IV|Lower leg CT W and WO contrast IV
C2826012|T102|strict|30870-0|LNC|Lower leg MRI W and WO contrast IV|Lower leg MRI W and WO contrast IV
C2826012|T102|strict|42697-3|LNC|Lower leg - bilateral MRI W and WO contrast IV|Lower leg - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36409-1|LNC|Lower leg - left CT W and WO contrast IV|Lower leg - left CT W and WO contrast IV
C2826012|T102|strict|36410-9|LNC|Lower leg - left MRI W and WO contrast IV|Lower leg - left MRI W and WO contrast IV
C2826012|T102|strict|36411-7|LNC|Lower leg - right CT W and WO contrast IV|Lower leg - right CT W and WO contrast IV
C2826012|T102|strict|36412-5|LNC|Lower leg - right MRI W and WO contrast IV|Lower leg - right MRI W and WO contrast IV
C2826012|T102|strict|36383-8|LNC|Mandible CT W and WO contrast IV|Mandible CT W and WO contrast IV
C2826012|T102|strict|37272-2|LNC|Mediastinum MRI W and WO contrast IV|Mediastinum MRI W and WO contrast IV
C2826012|T102|strict|48443-6|LNC|Nasopharynx CT W and WO contrast IV|Nasopharynx CT W and WO contrast IV
C2826012|T102|strict|36384-6|LNC|Nasopharynx MRI W and WO contrast IV|Nasopharynx MRI W and WO contrast IV
C2826012|T102|strict|30586-2|LNC|Neck CT W and WO contrast IV|Neck CT W and WO contrast IV
C2826012|T102|strict|24840-1|LNC|Neck MRI W and WO contrast IV|Neck MRI W and WO contrast IV
C2826012|T102|strict|36853-0|LNC|Neck veins MRI angiogram W and WO contrast IV|Neck veins MRI angiogram W and WO contrast IV
C2826012|T102|strict|30594-6|LNC|Neck vessels CT angiogram W and WO contrast IV|Neck vessels CT angiogram W and WO contrast IV
C2826012|T102|strict|36423-2|LNC|Neck vessels MRI angiogram W and WO contrast IV|Neck vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|48451-9|LNC|Orbit CT W and WO contrast IV|Orbit CT W and WO contrast IV
C2826012|T102|strict|36842-3|LNC|Orbit MRI W and WO contrast IV|Orbit MRI W and WO contrast IV
C2826012|T102|strict|43458-9|LNC|Orbit vessels MRI angiogram W and WO contrast IV|Orbit vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|24849-2|LNC|Orbit - bilateral CT W and WO contrast IV|Orbit - bilateral CT W and WO contrast IV
C2826012|T102|strict|24851-8|LNC|Orbit - bilateral MRI W and WO contrast IV|Orbit - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36843-1|LNC|Orbit - left MRI W and WO contrast IV|Orbit - left MRI W and WO contrast IV
C2826012|T102|strict|36844-9|LNC|Orbit - right MRI W and WO contrast IV|Orbit - right MRI W and WO contrast IV
C2826012|T102|strict|39029-4|LNC|Orbit and Face MRI W and WO contrast IV|Orbit and Face MRI W and WO contrast IV
C2826012|T102|strict|46310-9|LNC|Orbit and Face and Neck MRI W and WO contrast IV|Orbit and Face and Neck MRI W and WO contrast IV
C2826012|T102|strict|36845-6|LNC|Ovary MRI W and WO contrast IV|Ovary MRI W and WO contrast IV
C2826012|T102|strict|30614-2|LNC|Pancreas CT W and WO contrast IV|Pancreas CT W and WO contrast IV
C2826012|T102|strict|36385-3|LNC|Pancreas MRI W and WO contrast IV|Pancreas MRI W and WO contrast IV
C2826012|T102|strict|46311-7|LNC|Parotid gland CT W and WO contrast IV|Parotid gland CT W and WO contrast IV
C2826012|T102|strict|37265-6|LNC|Parotid gland MRI W and WO contrast IV|Parotid gland MRI W and WO contrast IV
C2826012|T102|strict|30616-7|LNC|Pelvis CT W and WO contrast IV|Pelvis CT W and WO contrast IV
C2826012|T102|strict|30674-6|LNC|Pelvis MRI W and WO contrast IV|Pelvis MRI W and WO contrast IV
C2826012|T102|strict|36854-8|LNC|Pelvis veins MRI angiogram W and WO contrast IV|Pelvis veins MRI angiogram W and WO contrast IV
C2826012|T102|strict|30623-3|LNC|Pelvis vessels CT angiogram W and WO contrast IV|Pelvis vessels CT angiogram W and WO contrast IV
C2826012|T102|strict|36863-9|LNC|Pelvis vessels MRI angiogram W and WO contrast IV|Pelvis vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|30672-0|LNC|Pelvis and Hip MRI W and WO contrast IV|Pelvis and Hip MRI W and WO contrast IV
C2826012|T102|strict|36835-7|LNC|Petrous bone CT W and WO contrast IV|Petrous bone CT W and WO contrast IV
C2826012|T102|strict|24904-5|LNC|Pituitary and Sella turcica CT W and WO contrast IV|Pituitary and Sella turcica CT W and WO contrast IV
C2826012|T102|strict|24879-9|LNC|Pituitary and Sella turcica MRI W and WO contrast IV|Pituitary and Sella turcica MRI W and WO contrast IV
C2826012|T102|strict|36414-1|LNC|Portal vein MRI angiogram W and WO contrast IV|Portal vein MRI angiogram W and WO contrast IV
C2826012|T102|strict|36387-9|LNC|Posterior fossa CT W and WO contrast IV|Posterior fossa CT W and WO contrast IV
C2826012|T102|strict|36388-7|LNC|Posterior fossa MRI W and WO contrast IV|Posterior fossa MRI W and WO contrast IV
C2826012|T102|strict|36389-5|LNC|Prostate MRI W and WO contrast IV|Prostate MRI W and WO contrast IV
C2826012|T102|strict|36275-6|LNC|Renal artery MRI angiogram W and WO contrast IV|Renal artery MRI angiogram W and WO contrast IV
C2826012|T102|strict|36415-8|LNC|Renal vein MRI angiogram W and WO contrast IV|Renal vein MRI angiogram W and WO contrast IV
C2826012|T102|strict|44134-5|LNC|Renal vessels MRI angiogram W and WO contrast IV|Renal vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|36375-4|LNC|Sacroiliac Joint CT W and WO contrast IV|Sacroiliac Joint CT W and WO contrast IV
C2826012|T102|strict|36376-2|LNC|Sacroiliac Joint MRI W and WO contrast IV|Sacroiliac Joint MRI W and WO contrast IV
C2826012|T102|strict|36390-3|LNC|Sacrum CT W and WO contrast IV|Sacrum CT W and WO contrast IV
C2826012|T102|strict|36391-1|LNC|Sacrum MRI W and WO contrast IV|Sacrum MRI W and WO contrast IV
C2826012|T102|strict|36392-9|LNC|Sacrum and Coccyx MRI W and WO contrast IV|Sacrum and Coccyx MRI W and WO contrast IV
C2826012|T102|strict|36393-7|LNC|Scapula - left MRI W and WO contrast IV|Scapula - left MRI W and WO contrast IV
C2826012|T102|strict|36394-5|LNC|Scapula - right MRI W and WO contrast IV|Scapula - right MRI W and WO contrast IV
C2826012|T102|strict|36406-7|LNC|Scrotum and Testicle MRI W and WO contrast IV|Scrotum and Testicle MRI W and WO contrast IV
C2826012|T102|strict|36395-2|LNC|Shoulder CT W and WO contrast IV|Shoulder CT W and WO contrast IV
C2826012|T102|strict|24906-0|LNC|Shoulder MRI W and WO contrast IV|Shoulder MRI W and WO contrast IV
C2826012|T102|strict|36864-7|LNC|Shoulder vessels - left MRI angiogram W and WO contrast IV|Shoulder vessels - left MRI angiogram W and WO contrast IV
C2826012|T102|strict|36865-4|LNC|Shoulder vessels - right MRI angiogram W and WO contrast IV|Shoulder vessels - right MRI angiogram W and WO contrast IV
C2826012|T102|strict|26202-2|LNC|Shoulder - bilateral MRI W and WO contrast IV|Shoulder - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36396-0|LNC|Shoulder - left CT W and WO contrast IV|Shoulder - left CT W and WO contrast IV
C2826012|T102|strict|26203-0|LNC|Shoulder - left MRI W and WO contrast IV|Shoulder - left MRI W and WO contrast IV
C2826012|T102|strict|36397-8|LNC|Shoulder - right CT W and WO contrast IV|Shoulder - right CT W and WO contrast IV
C2826012|T102|strict|26204-8|LNC|Shoulder - right MRI W and WO contrast IV|Shoulder - right MRI W and WO contrast IV
C2826012|T102|strict|36398-6|LNC|Sinuses CT W and WO contrast IV|Sinuses CT W and WO contrast IV
C2826012|T102|strict|30663-9|LNC|Sinuses MRI W and WO contrast IV|Sinuses MRI W and WO contrast IV
C2826012|T102|strict|44111-3|LNC|Skull.base CT W and WO contrast IV|Skull.base CT W and WO contrast IV
C2826012|T102|strict|69220-2|LNC|Skull.base MRI W and WO contrast IV|Skull.base MRI W and WO contrast IV
C2826012|T102|strict|37277-1|LNC|Spinal vein MRI angiogram W and WO contrast IV|Spinal vein MRI angiogram W and WO contrast IV
C2826012|T102|strict|36399-4|LNC|Spine CT W and WO contrast IV|Spine CT W and WO contrast IV
C2826012|T102|strict|36400-0|LNC|Spine MRI W and WO contrast IV|Spine MRI W and WO contrast IV
C2826012|T102|strict|37505-5|LNC|Spine vessels MRI angiogram W and WO contrast IV|Spine vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|36401-8|LNC|Spine Cervical CT W and WO contrast IV|Spine Cervical CT W and WO contrast IV
C2826012|T102|strict|24937-5|LNC|Spine Cervical MRI W and WO contrast IV|Spine Cervical MRI W and WO contrast IV
C2826012|T102|strict|37506-3|LNC|Cervical Spine vessels MRI angiogram W and WO contrast IV|Cervical Spine vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|43456-3|LNC|Spine Cervical and Spine Thoracic MRI W and WO contrast IV|Spine Cervical and Spine Thoracic MRI W and WO contrast IV
C2826012|T102|strict|30855-1|LNC|Spine Cervical and Thoracic and Lumbar MRI W and WO contrast IV|Spine Cervical and Thoracic and Lumbar MRI W and WO contrast IV
C2826012|T102|strict|36402-6|LNC|Spine Lumbar CT W and WO contrast IV|Spine Lumbar CT W and WO contrast IV
C2826012|T102|strict|24967-2|LNC|Spine Lumbar MRI W and WO contrast IV|Spine Lumbar MRI W and WO contrast IV
C2826012|T102|strict|37507-1|LNC|Lumbar Spine vessels MRI angiogram W and WO contrast IV|Lumbar Spine vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|36403-4|LNC|Spine Thoracic CT W and WO contrast IV|Spine Thoracic CT W and WO contrast IV
C2826012|T102|strict|24981-3|LNC|Spine Thoracic MRI W and WO contrast IV|Spine Thoracic MRI W and WO contrast IV
C2826012|T102|strict|37508-9|LNC|Thoracic Spine vessels MRI angiogram W and WO contrast IV|Thoracic Spine vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|24989-6|LNC|Spleen CT W and WO contrast IV|Spleen CT W and WO contrast IV
C2826012|T102|strict|36404-2|LNC|Spleen MRI W and WO contrast IV|Spleen MRI W and WO contrast IV
C2826012|T102|strict|37266-4|LNC|Sternoclavicular Joint CT W and WO contrast IV|Sternoclavicular Joint CT W and WO contrast IV
C2826012|T102|strict|36405-9|LNC|Sternum CT W and WO contrast IV|Sternum CT W and WO contrast IV
C2826012|T102|strict|44231-9|LNC|Superior mesenteric vessels MRI angiogram W and WO contrast IV|Superior mesenteric vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|36837-3|LNC|Temporal bone CT W and WO contrast IV|Temporal bone CT W and WO contrast IV
C2826012|T102|strict|37267-2|LNC|Temporomandibular joint CT W and WO contrast IV|Temporomandibular joint CT W and WO contrast IV
C2826012|T102|strict|37268-0|LNC|Temporomandibular joint MRI W and WO contrast IV|Temporomandibular joint MRI W and WO contrast IV
C2826012|T102|strict|37269-8|LNC|Temporomandibular joint - bilateral MRI W and WO contrast IV|Temporomandibular joint - bilateral MRI W and WO contrast IV
C2826012|T102|strict|37270-6|LNC|Temporomandibular joint - left MRI W and WO contrast IV|Temporomandibular joint - left MRI W and WO contrast IV
C2826012|T102|strict|37271-4|LNC|Temporomandibular joint - right MRI W and WO contrast IV|Temporomandibular joint - right MRI W and WO contrast IV
C2826012|T102|strict|24703-1|LNC|Thigh MRI W and WO contrast IV|Thigh MRI W and WO contrast IV
C2826012|T102|strict|26196-6|LNC|Thigh - bilateral MRI W and WO contrast IV|Thigh - bilateral MRI W and WO contrast IV
C2826012|T102|strict|26197-4|LNC|Thigh - left MRI W and WO contrast IV|Thigh - left MRI W and WO contrast IV
C2826012|T102|strict|26198-2|LNC|Thigh - right MRI W and WO contrast IV|Thigh - right MRI W and WO contrast IV
C2826012|T102|strict|24583-7|LNC|Thoracic outlet MRI W and WO contrast IV|Thoracic outlet MRI W and WO contrast IV
C2826012|T102|strict|26190-9|LNC|Thoracic outlet - bilateral MRI W and WO contrast IV|Thoracic outlet - bilateral MRI W and WO contrast IV
C2826012|T102|strict|26191-7|LNC|Thoracic outlet - left MRI W and WO contrast IV|Thoracic outlet - left MRI W and WO contrast IV
C2826012|T102|strict|26192-5|LNC|Thoracic outlet - right MRI W and WO contrast IV|Thoracic outlet - right MRI W and WO contrast IV
C2826012|T102|strict|36407-5|LNC|Thyroid MRI W and WO contrast IV|Thyroid MRI W and WO contrast IV
C2826012|T102|strict|72241-3|LNC|Toes - left MRI W and WO contrast IV|Toes - left MRI W and WO contrast IV
C2826012|T102|strict|72238-9|LNC|Toes - right MRI W and WO contrast IV|Toes - right MRI W and WO contrast IV
C2826012|T102|strict|36366-3|LNC|Upper arm CT W and WO contrast IV|Upper arm CT W and WO contrast IV
C2826012|T102|strict|30690-2|LNC|Upper arm MRI W and WO contrast IV|Upper arm MRI W and WO contrast IV
C2826012|T102|strict|69181-6|LNC|Upper arm - bilateral MRI W and WO contrast IV|Upper arm - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36367-1|LNC|Upper arm - left CT W and WO contrast IV|Upper arm - left CT W and WO contrast IV
C2826012|T102|strict|36368-9|LNC|Upper arm - left MRI W and WO contrast IV|Upper arm - left MRI W and WO contrast IV
C2826012|T102|strict|36369-7|LNC|Upper arm - right CT W and WO contrast IV|Upper arm - right CT W and WO contrast IV
C2826012|T102|strict|36370-5|LNC|Upper arm - right MRI W and WO contrast IV|Upper arm - right MRI W and WO contrast IV
C2826012|T102|strict|36334-1|LNC|Upper extremity CT W and WO contrast IV|Upper extremity CT W and WO contrast IV
C2826012|T102|strict|39034-4|LNC|Upper extremity MRI W and WO contrast IV|Upper extremity MRI W and WO contrast IV
C2826012|T102|strict|36417-4|LNC|Upper extremity veins MRI angiogram W and WO contrast IV|Upper extremity veins MRI angiogram W and WO contrast IV
C2826012|T102|strict|36851-4|LNC|Upper extremity veins - left MRI angiogram W and WO contrast IV|Upper extremity veins - left MRI angiogram W and WO contrast IV
C2826012|T102|strict|36852-2|LNC|Upper extremity veins - right MRI angiogram W and WO contrast IV|Upper extremity veins - right MRI angiogram W and WO contrast IV
C2826012|T102|strict|36421-6|LNC|Upper extremity vessels CT angiogram W and WO contrast IV|Upper extremity vessels CT angiogram W and WO contrast IV
C2826012|T102|strict|36422-4|LNC|Upper extremity vessels MRI angiogram W and WO contrast IV|Upper extremity vessels MRI angiogram W and WO contrast IV
C2826012|T102|strict|46312-5|LNC|Upper extremity vessels - left CT angiogram W and WO contrast IV|Upper extremity vessels - left CT angiogram W and WO contrast IV
C2826012|T102|strict|36860-5|LNC|Upper extremity vessels - left MRI angiogram W and WO contrast IV|Upper extremity vessels - left MRI angiogram W and WO contrast IV
C2826012|T102|strict|46309-1|LNC|Upper extremity vessels - right CT angiogram W and WO contrast IV|Upper extremity vessels - right CT angiogram W and WO contrast IV
C2826012|T102|strict|36861-3|LNC|Upper extremity vessels - right MRI angiogram W and WO contrast IV|Upper extremity vessels - right MRI angiogram W and WO contrast IV
C2826012|T102|strict|69186-5|LNC|Upper extremity - bilateral MRI W and WO contrast IV|Upper extremity - bilateral MRI W and WO contrast IV
C2826012|T102|strict|36374-7|LNC|Upper extremity .joint MRI W and WO contrast IV|Upper extremity .joint MRI W and WO contrast IV
C2826012|T102|strict|36840-7|LNC|Upper extremity joint - left MRI W and WO contrast IV|Upper extremity joint - left MRI W and WO contrast IV
C2826012|T102|strict|36841-5|LNC|Upper extremity joint - right MRI W and WO contrast IV|Upper extremity joint - right MRI W and WO contrast IV
C2826012|T102|strict|36335-8|LNC|Upper extremity - left CT W and WO contrast IV|Upper extremity - left CT W and WO contrast IV
C2826012|T102|strict|38831-4|LNC|Upper extremity - left MRI W and WO contrast IV|Upper extremity - left MRI W and WO contrast IV
C2826012|T102|strict|36336-6|LNC|Upper extremity - right CT W and WO contrast IV|Upper extremity - right CT W and WO contrast IV
C2826012|T102|strict|36337-4|LNC|Upper extremity - right MRI W and WO contrast IV|Upper extremity - right MRI W and WO contrast IV
C2826012|T102|strict|36413-3|LNC|Uterus MRI W and WO contrast IV|Uterus MRI W and WO contrast IV
C2826012|T102|strict|36418-2|LNC|Inferior vena cava MRI W and WO contrast IV|Inferior vena cava MRI W and WO contrast IV
C2826012|T102|strict|36419-0|LNC|Superior vena cava MRI W and WO contrast IV|Superior vena cava MRI W and WO contrast IV
C2826012|T102|strict|37457-9|LNC|Wrist CT W and WO contrast IV|Wrist CT W and WO contrast IV
C2826012|T102|strict|25035-7|LNC|Wrist MRI W and WO contrast IV|Wrist MRI W and WO contrast IV
C2826012|T102|strict|26205-5|LNC|Wrist - bilateral MRI W and WO contrast IV|Wrist - bilateral MRI W and WO contrast IV
C2826012|T102|strict|37458-7|LNC|Wrist - left CT W and WO contrast IV|Wrist - left CT W and WO contrast IV
C2826012|T102|strict|26206-3|LNC|Wrist - left MRI W and WO contrast IV|Wrist - left MRI W and WO contrast IV
C2826012|T102|strict|38802-5|LNC|Wrist - right CT W and WO contrast IV|Wrist - right CT W and WO contrast IV
C2826012|T102|strict|26207-1|LNC|Wrist - right MRI W and WO contrast IV|Wrist - right MRI W and WO contrast IV
C2826012|T102|strict|42298-0|LNC|Unspecified body region MRI W and WO contrast IV|Unspecified body region MRI W and WO contrast IV
C2826012|T102|strict|24588-6|LNC|Brain MRI W and WO contrast IV and W anesthesia|Brain MRI W and WO contrast IV and W anesthesia
C2826012|T102|strict|72244-7|LNC|Pelvis MRI W and WO contrast IV and W endorectal coil|Pelvis MRI W and WO contrast IV and W endorectal coil
C2826012|T102|strict|43448-0|LNC|Liver MRI W and WO ferumoxides IV|Liver MRI W and WO ferumoxides IV
C2826012|T102|strict|46318-2|LNC|Abdomen CT W and WO reduced contrast volume IV|Abdomen CT W and WO reduced contrast volume IV
C2826012|T102|strict|46317-4|LNC|Chest CT W and WO reduced contrast volume IV|Chest CT W and WO reduced contrast volume IV
C2826012|T102|strict|46315-8|LNC|Facial bones and Maxilla CT W and WO reduced contrast volume IV|Facial bones and Maxilla CT W and WO reduced contrast volume IV
C2826012|T102|strict|46316-6|LNC|Head CT W and WO reduced contrast volume IV|Head CT W and WO reduced contrast volume IV
C2826012|T102|strict|46314-1|LNC|Internal auditory canal CT W and WO reduced contrast volume IV|Internal auditory canal CT W and WO reduced contrast volume IV
C2826012|T102|strict|46313-3|LNC|Pelvis CT W and WO reduced contrast volume IV|Pelvis CT W and WO reduced contrast volume IV
C2826012|T102|strict|60515-4|LNC|Rectum and Colon CT 3D W air contrast PR|Rectum and Colon CT 3D W air contrast PR
C2826012|T102|strict|24586-0|LNC|Brain MRI W anesthesia|Brain MRI W anesthesia
C2826012|T102|strict|24936-7|LNC|Spine Cervical MRI W anesthesia|Spine Cervical MRI W anesthesia
C2826012|T102|strict|24977-1|LNC|Spine Lumbar MRI W anesthesia|Spine Lumbar MRI W anesthesia
C2826012|T102|strict|25046-4|LNC|Unspecified body region CT W anesthesia|Unspecified body region CT W anesthesia
C2826012|T102|strict|38022-0|LNC|Gallbladder US W cholecystokinin|Gallbladder US W cholecystokinin
C2826012|T102|strict|25047-2|LNC|Unspecified body region CT W conscious sedation|Unspecified body region CT W conscious sedation
C2826012|T102|strict|25057-1|LNC|Unspecified body region MRI W conscious sedation|Unspecified body region MRI W conscious sedation
C2826012|T102|strict|30599-5|LNC|Abdomen CT W contrast|Abdomen CT W contrast
C2826012|T102|strict|24567-0|LNC|Abdomen retroperitoneum CT W contrast|Abdomen retroperitoneum CT W contrast
C2826012|T102|strict|38055-0|LNC|Unspecified body region US W contrast|Unspecified body region US W contrast
C2826012|T102|strict|36809-2|LNC|Hepatic artery CT angiogram W contrast IA|Hepatic artery CT angiogram W contrast IA
C2826012|T102|strict|69162-6|LNC|Pulmonary artery - bilateral MRI angiogram W contrast IA|Pulmonary artery - bilateral MRI angiogram W contrast IA
C2826012|T102|strict|69238-4|LNC|Urinary Bladder and Urethra SPECT W contrast intra bladder during voiding|Urinary Bladder and Urethra SPECT W contrast intra bladder during voiding
C2826012|T102|strict|30853-6|LNC|Breast duct US W contrast intra duct|Breast duct US W contrast intra duct
C2826012|T102|strict|36941-3|LNC|Salivary gland CT W contrast intra salivary duct|Salivary gland CT W contrast intra salivary duct
C2826012|T102|strict|37237-5|LNC|Sinus tract CT W contrast intra sinus tract|Sinus tract CT W contrast intra sinus tract
C2826012|T102|strict|36115-4|LNC|Ankle MRI W contrast intraarticular|Ankle MRI W contrast intraarticular
C2826012|T102|strict|69102-2|LNC|Ankle - left CT W contrast intraarticular|Ankle - left CT W contrast intraarticular
C2826012|T102|strict|36116-2|LNC|Ankle - left MRI W contrast intraarticular|Ankle - left MRI W contrast intraarticular
C2826012|T102|strict|69109-7|LNC|Ankle - right CT W contrast intraarticular|Ankle - right CT W contrast intraarticular
C2826012|T102|strict|36117-0|LNC|Ankle - right MRI W contrast intraarticular|Ankle - right MRI W contrast intraarticular
C2826012|T102|strict|46319-0|LNC|Elbow MRI W contrast intraarticular|Elbow MRI W contrast intraarticular
C2826012|T102|strict|69103-0|LNC|Elbow - left CT W contrast intraarticular|Elbow - left CT W contrast intraarticular
C2826012|T102|strict|36118-8|LNC|Elbow - left MRI W contrast intraarticular|Elbow - left MRI W contrast intraarticular
C2826012|T102|strict|69110-5|LNC|Elbow - right CT W contrast intraarticular|Elbow - right CT W contrast intraarticular
C2826012|T102|strict|36119-6|LNC|Elbow - right MRI W contrast intraarticular|Elbow - right MRI W contrast intraarticular
C2826012|T102|strict|36120-4|LNC|Hip MRI W contrast intraarticular|Hip MRI W contrast intraarticular
C2826012|T102|strict|69105-5|LNC|Hip - left CT W contrast intraarticular|Hip - left CT W contrast intraarticular
C2826012|T102|strict|36121-2|LNC|Hip - left MRI W contrast intraarticular|Hip - left MRI W contrast intraarticular
C2826012|T102|strict|69112-1|LNC|Hip - right CT W contrast intraarticular|Hip - right CT W contrast intraarticular
C2826012|T102|strict|36122-0|LNC|Hip - right MRI W contrast intraarticular|Hip - right MRI W contrast intraarticular
C2826012|T102|strict|36124-6|LNC|Knee CT W contrast intraarticular|Knee CT W contrast intraarticular
C2826012|T102|strict|36125-3|LNC|Knee MRI W contrast intraarticular|Knee MRI W contrast intraarticular
C2826012|T102|strict|69106-3|LNC|Knee - left CT W contrast intraarticular|Knee - left CT W contrast intraarticular
C2826012|T102|strict|36126-1|LNC|Knee - left MRI W contrast intraarticular|Knee - left MRI W contrast intraarticular
C2826012|T102|strict|69114-7|LNC|Knee - right CT W contrast intraarticular|Knee - right CT W contrast intraarticular
C2826012|T102|strict|36127-9|LNC|Knee - right MRI W contrast intraarticular|Knee - right MRI W contrast intraarticular
C2826012|T102|strict|37238-3|LNC|Lower Extremity Joint CT W contrast intraarticular|Lower Extremity Joint CT W contrast intraarticular
C2826012|T102|strict|69210-3|LNC|Lower Extremity Joint MRI W contrast intraarticular|Lower Extremity Joint MRI W contrast intraarticular
C2826012|T102|strict|36123-8|LNC|Sacroiliac Joint CT W contrast intraarticular|Sacroiliac Joint CT W contrast intraarticular
C2826012|T102|strict|36128-7|LNC|Shoulder CT W contrast intraarticular|Shoulder CT W contrast intraarticular
C2826012|T102|strict|36129-5|LNC|Shoulder MRI W contrast intraarticular|Shoulder MRI W contrast intraarticular
C2826012|T102|strict|38828-0|LNC|Shoulder - left CT W contrast intraarticular|Shoulder - left CT W contrast intraarticular
C2826012|T102|strict|36130-3|LNC|Shoulder - left MRI W contrast intraarticular|Shoulder - left MRI W contrast intraarticular
C2826012|T102|strict|36131-1|LNC|Shoulder - right CT W contrast intraarticular|Shoulder - right CT W contrast intraarticular
C2826012|T102|strict|36132-9|LNC|Shoulder - right MRI W contrast intraarticular|Shoulder - right MRI W contrast intraarticular
C2826012|T102|strict|36810-0|LNC|Upper Joint CT W contrast intraarticular|Upper Joint CT W contrast intraarticular
C2826012|T102|strict|37444-7|LNC|Wrist MRI W contrast intraarticular|Wrist MRI W contrast intraarticular
C2826012|T102|strict|69107-1|LNC|Wrist - left CT W contrast intraarticular|Wrist - left CT W contrast intraarticular
C2826012|T102|strict|37445-4|LNC|Wrist - left MRI W contrast intraarticular|Wrist - left MRI W contrast intraarticular
C2826012|T102|strict|69115-4|LNC|Wrist - right CT W contrast intraarticular|Wrist - right CT W contrast intraarticular
C2826012|T102|strict|37446-2|LNC|Wrist - right MRI W contrast intraarticular|Wrist - right MRI W contrast intraarticular
C2826012|T102|strict|36811-8|LNC|Joint CT W contrast intraarticular|Joint CT W contrast intraarticular
C2826012|T102|strict|36812-6|LNC|Joint MRI W contrast intraarticular|Joint MRI W contrast intraarticular
C2826012|T102|strict|39322-3|LNC|Spine CT W contrast intradisc|Spine CT W contrast intradisc
C2826012|T102|strict|37496-7|LNC|Spine Cervical CT W contrast intradisc|Spine Cervical CT W contrast intradisc
C2826012|T102|strict|37509-7|LNC|Spine Lumbar CT W contrast intradisc|Spine Lumbar CT W contrast intradisc
C2826012|T102|strict|70931-1|LNC|Spine Thoracic CT W contrast intradisc|Spine Thoracic CT W contrast intradisc
C2826012|T102|strict|24734-6|LNC|Head Cistern CT W contrast IT|Head Cistern CT W contrast IT
C2826012|T102|strict|47985-7|LNC|Spine CT W contrast IT|Spine CT W contrast IT
C2826012|T102|strict|24934-2|LNC|Spine Cervical CT W contrast IT|Spine Cervical CT W contrast IT
C2826012|T102|strict|48447-7|LNC|Spine Cervical MRI W contrast IT|Spine Cervical MRI W contrast IT
C2826012|T102|strict|24965-6|LNC|Spine Lumbar CT W contrast IT|Spine Lumbar CT W contrast IT
C2826012|T102|strict|48436-0|LNC|Spine Lumbar MRI W contrast IT|Spine Lumbar MRI W contrast IT
C2826012|T102|strict|30596-1|LNC|Spine Thoracic CT W contrast IT|Spine Thoracic CT W contrast IT
C2826012|T102|strict|48439-4|LNC|Spine Thoracic MRI W contrast IT|Spine Thoracic MRI W contrast IT
C2826012|T102|strict|36134-5|LNC|Abdomen MRI W contrast IV|Abdomen MRI W contrast IV
C2826012|T102|strict|36813-4|LNC|Abdomen and Pelvis CT W contrast IV|Abdomen and Pelvis CT W contrast IV
C2826012|T102|strict|36828-2|LNC|Abdominal vessels CT angiogram W contrast IV|Abdominal vessels CT angiogram W contrast IV
C2826012|T102|strict|24533-2|LNC|Abdominal vessels MRI angiogram W contrast IV|Abdominal vessels MRI angiogram W contrast IV
C2826012|T102|strict|69908-2|LNC|Abdominal vessels and Pelvis vessels CT angiogram W contrast IV|Abdominal vessels and Pelvis vessels CT angiogram W contrast IV
C2826012|T102|strict|36943-9|LNC|Adrenal gland CT W contrast IV|Adrenal gland CT W contrast IV
C2826012|T102|strict|44124-6|LNC|Adrenal gland MRI W contrast IV|Adrenal gland MRI W contrast IV
C2826012|T102|strict|36135-2|LNC|Ankle CT W contrast IV|Ankle CT W contrast IV
C2826012|T102|strict|36136-0|LNC|Ankle MRI W contrast IV|Ankle MRI W contrast IV
C2826012|T102|strict|69163-4|LNC|Ankle - bilateral MRI W contrast IV|Ankle - bilateral MRI W contrast IV
C2826012|T102|strict|36137-8|LNC|Ankle - left CT W contrast IV|Ankle - left CT W contrast IV
C2826012|T102|strict|36138-6|LNC|Ankle - left MRI W contrast IV|Ankle - left MRI W contrast IV
C2826012|T102|strict|36139-4|LNC|Ankle - right CT W contrast IV|Ankle - right CT W contrast IV
C2826012|T102|strict|36140-2|LNC|Ankle - right MRI W contrast IV|Ankle - right MRI W contrast IV
C2826012|T102|strict|36142-8|LNC|Aorta CT W contrast IV|Aorta CT W contrast IV
C2826012|T102|strict|36141-0|LNC|Aorta CT angiogram W contrast IV|Aorta CT angiogram W contrast IV
C2826012|T102|strict|36143-6|LNC|Aorta abdominal CT W contrast IV|Aorta abdominal CT W contrast IV
C2826012|T102|strict|24545-6|LNC|Aorta thoracic CT W contrast IV|Aorta thoracic CT W contrast IV
C2826012|T102|strict|72255-3|LNC|Aorta and Femoral artery - bilateral CT angiogram W contrast IV|Aorta and Femoral artery - bilateral CT angiogram W contrast IV
C2826012|T102|strict|43503-2|LNC|Aorta and Lower extremity vessels CT angiogram W contrast IV|Aorta and Lower extremity vessels CT angiogram W contrast IV
C2826012|T102|strict|36144-4|LNC|Aortic arch CT angiogram W contrast IV|Aortic arch CT angiogram W contrast IV
C2826012|T102|strict|37499-1|LNC|Aortic stent CT angiogram W contrast IV|Aortic stent CT angiogram W contrast IV
C2826012|T102|strict|36145-1|LNC|Appendix CT W contrast IV|Appendix CT W contrast IV
C2826012|T102|strict|43504-0|LNC|Axilla - left MRI W contrast IV|Axilla - left MRI W contrast IV
C2826012|T102|strict|43505-7|LNC|Axilla - right MRI W contrast IV|Axilla - right MRI W contrast IV
C2826012|T102|strict|44125-3|LNC|Biliary ducts and Pancreatic duct MRI W contrast IV|Biliary ducts and Pancreatic duct MRI W contrast IV
C2826012|T102|strict|69095-8|LNC|Bladder CT W contrast IV|Bladder CT W contrast IV
C2826012|T102|strict|24589-4|LNC|Brain MRI W contrast IV|Brain MRI W contrast IV
C2826012|T102|strict|48444-4|LNC|Brain.temporal MRI W contrast IV|Brain.temporal MRI W contrast IV
C2826012|T102|strict|37239-1|LNC|Brain and Internal auditory canal MRI W contrast IV|Brain and Internal auditory canal MRI W contrast IV
C2826012|T102|strict|37215-1|LNC|Brain and Larynx MRI W contrast IV|Brain and Larynx MRI W contrast IV
C2826012|T102|strict|42391-3|LNC|Brain and Pituitary and Sella turcica MRI W contrast IV|Brain and Pituitary and Sella turcica MRI W contrast IV
C2826012|T102|strict|36149-3|LNC|Breast MRI W contrast IV|Breast MRI W contrast IV
C2826012|T102|strict|69190-7|LNC|Breast implant MRI W contrast IV|Breast implant MRI W contrast IV
C2826012|T102|strict|69167-5|LNC|Breast implant - bilateral MRI W contrast IV|Breast implant - bilateral MRI W contrast IV
C2826012|T102|strict|36150-1|LNC|Breast - bilateral MRI W contrast IV|Breast - bilateral MRI W contrast IV
C2826012|T102|strict|36151-9|LNC|Breast - left MRI W contrast IV|Breast - left MRI W contrast IV
C2826012|T102|strict|36152-7|LNC|Breast - right MRI W contrast IV|Breast - right MRI W contrast IV
C2826012|T102|strict|46323-2|LNC|Breast - unilateral MRI W contrast IV|Breast - unilateral MRI W contrast IV
C2826012|T102|strict|36198-0|LNC|Calcaneus CT W contrast IV|Calcaneus CT W contrast IV
C2826012|T102|strict|36153-5|LNC|Calcaneus - left CT W contrast IV|Calcaneus - left CT W contrast IV
C2826012|T102|strict|36154-3|LNC|Calcaneus - right CT W contrast IV|Calcaneus - right CT W contrast IV
C2826012|T102|strict|36146-9|LNC|Carotid artery CT angiogram W contrast IV|Carotid artery CT angiogram W contrast IV
C2826012|T102|strict|36829-0|LNC|Carotid vessel MRI angiogram W contrast IV|Carotid vessel MRI angiogram W contrast IV
C2826012|T102|strict|24628-0|LNC|Chest CT W contrast IV|Chest CT W contrast IV
C2826012|T102|strict|36156-8|LNC|Chest MRI W contrast IV|Chest MRI W contrast IV
C2826012|T102|strict|36266-5|LNC|Chest vessels CT angiogram W contrast IV|Chest vessels CT angiogram W contrast IV
C2826012|T102|strict|24659-5|LNC|Chest vessels MRI angiogram W contrast IV|Chest vessels MRI angiogram W contrast IV
C2826012|T102|strict|42275-8|LNC|Chest and Abdomen CT W contrast IV|Chest and Abdomen CT W contrast IV
C2826012|T102|strict|36942-1|LNC|Chest and Abdomen MRI W contrast IV|Chest and Abdomen MRI W contrast IV
C2826012|T102|strict|72254-6|LNC|Chest and Abdomen and Pelvis CT W contrast IV|Chest and Abdomen and Pelvis CT W contrast IV
C2826012|T102|strict|37254-0|LNC|Circle of Willis MRI angiogram W contrast IV|Circle of Willis MRI angiogram W contrast IV
C2826012|T102|strict|42694-0|LNC|Clavicle MRI W contrast IV|Clavicle MRI W contrast IV
C2826012|T102|strict|48457-6|LNC|Clavicle - left MRI W contrast IV|Clavicle - left MRI W contrast IV
C2826012|T102|strict|48456-8|LNC|Clavicle - right MRI W contrast IV|Clavicle - right MRI W contrast IV
C2826012|T102|strict|36157-6|LNC|Elbow CT W contrast IV|Elbow CT W contrast IV
C2826012|T102|strict|36158-4|LNC|Elbow MRI W contrast IV|Elbow MRI W contrast IV
C2826012|T102|strict|69170-9|LNC|Elbow - bilateral MRI W contrast IV|Elbow - bilateral MRI W contrast IV
C2826012|T102|strict|36159-2|LNC|Elbow - left CT W contrast IV|Elbow - left CT W contrast IV
C2826012|T102|strict|36160-0|LNC|Elbow - left MRI W contrast IV|Elbow - left MRI W contrast IV
C2826012|T102|strict|36161-8|LNC|Elbow - right CT W contrast IV|Elbow - right CT W contrast IV
C2826012|T102|strict|36162-6|LNC|Elbow - right MRI W contrast IV|Elbow - right MRI W contrast IV
C2826012|T102|strict|24691-8|LNC|Extremity CT W contrast IV|Extremity CT W contrast IV
C2826012|T102|strict|26184-2|LNC|Extremity - bilateral CT W contrast IV|Extremity - bilateral CT W contrast IV
C2826012|T102|strict|26185-9|LNC|Extremity - left CT W contrast IV|Extremity - left CT W contrast IV
C2826012|T102|strict|26186-7|LNC|Extremity - right CT W contrast IV|Extremity - right CT W contrast IV
C2826012|T102|strict|36148-5|LNC|Face MRI W contrast IV|Face MRI W contrast IV
C2826012|T102|strict|30801-5|LNC|Facial bones and Maxilla CT W contrast IV|Facial bones and Maxilla CT W contrast IV
C2826012|T102|strict|24697-5|LNC|Facial bones and Sinuses CT W contrast IV|Facial bones and Sinuses CT W contrast IV
C2826012|T102|strict|36172-5|LNC|Femur CT W contrast IV|Femur CT W contrast IV
C2826012|T102|strict|69172-5|LNC|Femur - bilateral MRI W contrast IV|Femur - bilateral MRI W contrast IV
C2826012|T102|strict|36174-1|LNC|Femur - left CT W contrast IV|Femur - left CT W contrast IV
C2826012|T102|strict|36176-6|LNC|Femur - right CT W contrast IV|Femur - right CT W contrast IV
C2826012|T102|strict|69195-6|LNC|Finger MRI W contrast IV|Finger MRI W contrast IV
C2826012|T102|strict|69205-3|LNC|Finger - left MRI W contrast IV|Finger - left MRI W contrast IV
C2826012|T102|strict|69215-2|LNC|Finger - right MRI W contrast IV|Finger - right MRI W contrast IV
C2826012|T102|strict|36178-2|LNC|Foot CT W contrast IV|Foot CT W contrast IV
C2826012|T102|strict|36179-0|LNC|Foot MRI W contrast IV|Foot MRI W contrast IV
C2826012|T102|strict|36180-8|LNC|Foot - bilateral MRI W contrast IV|Foot - bilateral MRI W contrast IV
C2826012|T102|strict|36181-6|LNC|Foot - left CT W contrast IV|Foot - left CT W contrast IV
C2826012|T102|strict|36182-4|LNC|Foot - left MRI W contrast IV|Foot - left MRI W contrast IV
C2826012|T102|strict|36183-2|LNC|Foot - right CT W contrast IV|Foot - right CT W contrast IV
C2826012|T102|strict|36184-0|LNC|Foot - right MRI W contrast IV|Foot - right MRI W contrast IV
C2826012|T102|strict|36185-7|LNC|Forearm CT W contrast IV|Forearm CT W contrast IV
C2826012|T102|strict|36186-5|LNC|Forearm MRI W contrast IV|Forearm MRI W contrast IV
C2826012|T102|strict|69175-8|LNC|Forearm - bilateral MRI W contrast IV|Forearm - bilateral MRI W contrast IV
C2826012|T102|strict|36187-3|LNC|Forearm - left CT W contrast IV|Forearm - left CT W contrast IV
C2826012|T102|strict|36188-1|LNC|Forearm - left MRI W contrast IV|Forearm - left MRI W contrast IV
C2826012|T102|strict|36189-9|LNC|Forearm - right CT W contrast IV|Forearm - right CT W contrast IV
C2826012|T102|strict|36190-7|LNC|Forearm - right MRI W contrast IV|Forearm - right MRI W contrast IV
C2826012|T102|strict|36191-5|LNC|Hand CT W contrast IV|Hand CT W contrast IV
C2826012|T102|strict|36192-3|LNC|Hand MRI W contrast IV|Hand MRI W contrast IV
C2826012|T102|strict|69178-2|LNC|Hand - bilateral MRI W contrast IV|Hand - bilateral MRI W contrast IV
C2826012|T102|strict|36193-1|LNC|Hand - left CT W contrast IV|Hand - left CT W contrast IV
C2826012|T102|strict|36194-9|LNC|Hand - left MRI W contrast IV|Hand - left MRI W contrast IV
C2826012|T102|strict|36195-6|LNC|Hand - right CT W contrast IV|Hand - right CT W contrast IV
C2826012|T102|strict|36196-4|LNC|Hand - right MRI W contrast IV|Hand - right MRI W contrast IV
C2826012|T102|strict|24727-0|LNC|Head CT W contrast IV|Head CT W contrast IV
C2826012|T102|strict|36814-2|LNC|Head arteries CT angiogram W contrast IV|Head arteries CT angiogram W contrast IV
C2826012|T102|strict|36826-6|LNC|Head veins MRI angiogram W contrast IV|Head veins MRI angiogram W contrast IV
C2826012|T102|strict|36830-8|LNC|Head vessels CT angiogram W contrast IV|Head vessels CT angiogram W contrast IV
C2826012|T102|strict|24593-6|LNC|Head vessels MRI angiogram W contrast IV|Head vessels MRI angiogram W contrast IV
C2826012|T102|strict|37498-3|LNC|Head vessels and Neck vessels CT angiogram W contrast IV|Head vessels and Neck vessels CT angiogram W contrast IV
C2826012|T102|strict|24747-8|LNC|Head Sagittal Sinus MRI angiogram W contrast IV|Head Sagittal Sinus MRI angiogram W contrast IV
C2826012|T102|strict|36197-2|LNC|Heart MRI W contrast IV|Heart MRI W contrast IV
C2826012|T102|strict|36200-4|LNC|Hip CT W contrast IV|Hip CT W contrast IV
C2826012|T102|strict|36199-8|LNC|Hip MRI W contrast IV|Hip MRI W contrast IV
C2826012|T102|strict|36201-2|LNC|Hip - bilateral CT W contrast IV|Hip - bilateral CT W contrast IV
C2826012|T102|strict|36202-0|LNC|Hip - bilateral MRI W contrast IV|Hip - bilateral MRI W contrast IV
C2826012|T102|strict|36203-8|LNC|Hip - left CT W contrast IV|Hip - left CT W contrast IV
C2826012|T102|strict|36204-6|LNC|Hip - left MRI W contrast IV|Hip - left MRI W contrast IV
C2826012|T102|strict|36205-3|LNC|Hip - right CT W contrast IV|Hip - right CT W contrast IV
C2826012|T102|strict|36206-1|LNC|Hip - right MRI W contrast IV|Hip - right MRI W contrast IV
C2826012|T102|strict|30583-9|LNC|Internal auditory canal CT W contrast IV|Internal auditory canal CT W contrast IV
C2826012|T102|strict|36155-0|LNC|Internal auditory canal MRI W contrast IV|Internal auditory canal MRI W contrast IV
C2826012|T102|strict|46322-4|LNC|Kidney CT W contrast IV|Kidney CT W contrast IV
C2826012|T102|strict|36113-9|LNC|Kidney MRI W contrast IV|Kidney MRI W contrast IV
C2826012|T102|strict|43766-5|LNC|Kidney - bilateral CT W contrast IV|Kidney - bilateral CT W contrast IV
C2826012|T102|strict|36219-4|LNC|Kidney - bilateral MRI W contrast IV|Kidney - bilateral MRI W contrast IV
C2826012|T102|strict|24790-8|LNC|Kidney - bilateral X-ray tomograph W contrast IV|Kidney - bilateral X-ray tomograph W contrast IV
C2826012|T102|strict|36220-2|LNC|Kidney - left MRI W contrast IV|Kidney - left MRI W contrast IV
C2826012|T102|strict|36221-0|LNC|Kidney - right MRI W contrast IV|Kidney - right MRI W contrast IV
C2826012|T102|strict|36222-8|LNC|Knee CT W contrast IV|Knee CT W contrast IV
C2826012|T102|strict|36223-6|LNC|Knee MRI W contrast IV|Knee MRI W contrast IV
C2826012|T102|strict|69088-3|LNC|Knee - bilateral CT W contrast IV|Knee - bilateral CT W contrast IV
C2826012|T102|strict|36224-4|LNC|Knee - bilateral MRI W contrast IV|Knee - bilateral MRI W contrast IV
C2826012|T102|strict|36225-1|LNC|Knee - left CT W contrast IV|Knee - left CT W contrast IV
C2826012|T102|strict|36226-9|LNC|Knee - left MRI W contrast IV|Knee - left MRI W contrast IV
C2826012|T102|strict|36227-7|LNC|Knee - right CT W contrast IV|Knee - right CT W contrast IV
C2826012|T102|strict|36228-5|LNC|Knee - right MRI W contrast IV|Knee - right MRI W contrast IV
C2826012|T102|strict|36229-3|LNC|Larynx CT W contrast IV|Larynx CT W contrast IV
C2826012|T102|strict|36230-1|LNC|Larynx MRI W contrast IV|Larynx MRI W contrast IV
C2826012|T102|strict|24815-3|LNC|Liver CT W contrast IV|Liver CT W contrast IV
C2826012|T102|strict|36231-9|LNC|Liver MRI W contrast IV|Liver MRI W contrast IV
C2826012|T102|strict|30624-1|LNC|Lower extremity CT W contrast IV|Lower extremity CT W contrast IV
C2826012|T102|strict|39293-6|LNC|Lower extremity MRI W contrast IV|Lower extremity MRI W contrast IV
C2826012|T102|strict|36824-1|LNC|Lower extremity veins - left CT W contrast IV|Lower extremity veins - left CT W contrast IV
C2826012|T102|strict|36825-8|LNC|Lower extremity veins - right CT W contrast IV|Lower extremity veins - right CT W contrast IV
C2826012|T102|strict|36831-6|LNC|Lower extremity vessels CT angiogram W contrast IV|Lower extremity vessels CT angiogram W contrast IV
C2826012|T102|strict|46324-0|LNC|Lower extremity vessels MRI angiogram W contrast IV|Lower extremity vessels MRI angiogram W contrast IV
C2826012|T102|strict|44135-2|LNC|Lower extremity vessels - bilateral MRI angiogram W contrast IV|Lower extremity vessels - bilateral MRI angiogram W contrast IV
C2826012|T102|strict|50755-8|LNC|Lower extremity - bilateral CT W contrast IV|Lower extremity - bilateral CT W contrast IV
C2826012|T102|strict|36163-4|LNC|Lower extremity - bilateral MRI W contrast IV|Lower extremity - bilateral MRI W contrast IV
C2826012|T102|strict|36213-7|LNC|Lower Extremity Joint MRI W contrast IV|Lower Extremity Joint MRI W contrast IV
C2826012|T102|strict|36214-5|LNC|Lower extremity joint - left MRI W contrast IV|Lower extremity joint - left MRI W contrast IV
C2826012|T102|strict|36215-2|LNC|Lower extremity joint - right MRI W contrast IV|Lower extremity joint - right MRI W contrast IV
C2826012|T102|strict|36164-2|LNC|Lower extremity - left CT W contrast IV|Lower extremity - left CT W contrast IV
C2826012|T102|strict|36165-9|LNC|Lower extremity - left MRI W contrast IV|Lower extremity - left MRI W contrast IV
C2826012|T102|strict|36166-7|LNC|Lower extremity - right CT W contrast IV|Lower extremity - right CT W contrast IV
C2826012|T102|strict|36167-5|LNC|Lower extremity - right MRI W contrast IV|Lower extremity - right MRI W contrast IV
C2826012|T102|strict|36258-2|LNC|Lower leg CT W contrast IV|Lower leg CT W contrast IV
C2826012|T102|strict|36259-0|LNC|Lower leg MRI W contrast IV|Lower leg MRI W contrast IV
C2826012|T102|strict|24820-3|LNC|Lower leg vessels MRI angiogram W contrast IV|Lower leg vessels MRI angiogram W contrast IV
C2826012|T102|strict|43512-3|LNC|Lower leg vessels - bilateral MRI angiogram W contrast IV|Lower leg vessels - bilateral MRI angiogram W contrast IV
C2826012|T102|strict|42695-7|LNC|Lower leg - bilateral MRI W contrast IV|Lower leg - bilateral MRI W contrast IV
C2826012|T102|strict|36260-8|LNC|Lower leg - left CT W contrast IV|Lower leg - left CT W contrast IV
C2826012|T102|strict|36261-6|LNC|Lower leg - left MRI W contrast IV|Lower leg - left MRI W contrast IV
C2826012|T102|strict|36262-4|LNC|Lower leg - right CT W contrast IV|Lower leg - right CT W contrast IV
C2826012|T102|strict|36263-2|LNC|Lower leg - right MRI W contrast IV|Lower leg - right MRI W contrast IV
C2826012|T102|strict|36232-7|LNC|Mandible CT W contrast IV|Mandible CT W contrast IV
C2826012|T102|strict|48446-9|LNC|Nasopharynx CT W contrast IV|Nasopharynx CT W contrast IV
C2826012|T102|strict|36233-5|LNC|Nasopharynx MRI W contrast IV|Nasopharynx MRI W contrast IV
C2826012|T102|strict|24836-9|LNC|Nasopharynx and Neck CT W contrast IV|Nasopharynx and Neck CT W contrast IV
C2826012|T102|strict|36235-0|LNC|Neck CT W contrast IV|Neck CT W contrast IV
C2826012|T102|strict|24841-9|LNC|Neck MRI W contrast IV|Neck MRI W contrast IV
C2826012|T102|strict|36827-4|LNC|Neck veins MRI angiogram W contrast IV|Neck veins MRI angiogram W contrast IV
C2826012|T102|strict|36234-3|LNC|Neck vessels CT angiogram W contrast IV|Neck vessels CT angiogram W contrast IV
C2826012|T102|strict|24844-3|LNC|Neck vessels MRI angiogram W contrast IV|Neck vessels MRI angiogram W contrast IV
C2826012|T102|strict|48449-3|LNC|Orbit CT W contrast IV|Orbit CT W contrast IV
C2826012|T102|strict|36820-9|LNC|Orbit MRI W contrast IV|Orbit MRI W contrast IV
C2826012|T102|strict|36832-4|LNC|Orbit vessels MRI angiogram W contrast IV|Orbit vessels MRI angiogram W contrast IV
C2826012|T102|strict|24850-0|LNC|Orbit - bilateral CT W contrast IV|Orbit - bilateral CT W contrast IV
C2826012|T102|strict|24852-6|LNC|Orbit - bilateral MRI W contrast IV|Orbit - bilateral MRI W contrast IV
C2826012|T102|strict|36821-7|LNC|Orbit - left MRI W contrast IV|Orbit - left MRI W contrast IV
C2826012|T102|strict|36822-5|LNC|Orbit - right MRI W contrast IV|Orbit - right MRI W contrast IV
C2826012|T102|strict|46320-8|LNC|Orbit and Face CT W contrast IV|Orbit and Face CT W contrast IV
C2826012|T102|strict|39038-5|LNC|Orbit and Face MRI W contrast IV|Orbit and Face MRI W contrast IV
C2826012|T102|strict|46321-6|LNC|Orbit and Face and Neck MRI W contrast IV|Orbit and Face and Neck MRI W contrast IV
C2826012|T102|strict|36823-3|LNC|Ovary MRI W contrast IV|Ovary MRI W contrast IV
C2826012|T102|strict|24858-3|LNC|Pancreas CT W contrast IV|Pancreas CT W contrast IV
C2826012|T102|strict|36236-8|LNC|Pancreas MRI W contrast IV|Pancreas MRI W contrast IV
C2826012|T102|strict|37240-9|LNC|Parotid gland CT W contrast IV|Parotid gland CT W contrast IV
C2826012|T102|strict|37241-7|LNC|Parotid gland MRI W contrast IV|Parotid gland MRI W contrast IV
C2826012|T102|strict|24866-6|LNC|Pelvis CT W contrast IV|Pelvis CT W contrast IV
C2826012|T102|strict|36237-6|LNC|Pelvis MRI W contrast IV|Pelvis MRI W contrast IV
C2826012|T102|strict|42294-9|LNC|Pelvis vessels CT angiogram W contrast IV|Pelvis vessels CT angiogram W contrast IV
C2826012|T102|strict|24873-2|LNC|Pelvis vessels MRI angiogram W contrast IV|Pelvis vessels MRI angiogram W contrast IV
C2826012|T102|strict|24878-1|LNC|Petrous bone CT W contrast IV|Petrous bone CT W contrast IV
C2826012|T102|strict|30590-4|LNC|Pituitary and Sella turcica CT W contrast IV|Pituitary and Sella turcica CT W contrast IV
C2826012|T102|strict|36238-4|LNC|Pituitary and Sella turcica MRI W contrast IV|Pituitary and Sella turcica MRI W contrast IV
C2826012|T102|strict|36242-6|LNC|Posterior fossa CT W contrast IV|Posterior fossa CT W contrast IV
C2826012|T102|strict|36243-4|LNC|Posterior fossa MRI W contrast IV|Posterior fossa MRI W contrast IV
C2826012|T102|strict|36244-2|LNC|Prostate MRI W contrast IV|Prostate MRI W contrast IV
C2826012|T102|strict|36147-7|LNC|Pulmonary artery CT angiogram W contrast IV|Pulmonary artery CT angiogram W contrast IV
C2826012|T102|strict|36833-2|LNC|Renal vessels CT angiogram W contrast IV|Renal vessels CT angiogram W contrast IV
C2826012|T102|strict|30887-4|LNC|Renal vessels MRI angiogram W contrast IV|Renal vessels MRI angiogram W contrast IV
C2826012|T102|strict|36217-8|LNC|Sacroiliac Joint CT W contrast IV|Sacroiliac Joint CT W contrast IV
C2826012|T102|strict|36218-6|LNC|Sacroiliac Joint MRI W contrast IV|Sacroiliac Joint MRI W contrast IV
C2826012|T102|strict|36245-9|LNC|Sacrum CT W contrast IV|Sacrum CT W contrast IV
C2826012|T102|strict|36246-7|LNC|Sacrum MRI W contrast IV|Sacrum MRI W contrast IV
C2826012|T102|strict|36247-5|LNC|Sacrum and Coccyx MRI W contrast IV|Sacrum and Coccyx MRI W contrast IV
C2826012|T102|strict|36248-3|LNC|Scapula - left MRI W contrast IV|Scapula - left MRI W contrast IV
C2826012|T102|strict|36249-1|LNC|Scapula - right MRI W contrast IV|Scapula - right MRI W contrast IV
C2826012|T102|strict|69221-0|LNC|Scrotum and Testicle MRI W contrast IV|Scrotum and Testicle MRI W contrast IV
C2826012|T102|strict|36250-9|LNC|Shoulder CT W contrast IV|Shoulder CT W contrast IV
C2826012|T102|strict|36251-7|LNC|Shoulder MRI W contrast IV|Shoulder MRI W contrast IV
C2826012|T102|strict|69184-0|LNC|Shoulder - bilateral MRI W contrast IV|Shoulder - bilateral MRI W contrast IV
C2826012|T102|strict|36252-5|LNC|Shoulder - left CT W contrast IV|Shoulder - left CT W contrast IV
C2826012|T102|strict|38830-6|LNC|Shoulder - left MRI W contrast IV|Shoulder - left MRI W contrast IV
C2826012|T102|strict|36253-3|LNC|Shoulder - right CT W contrast IV|Shoulder - right CT W contrast IV
C2826012|T102|strict|36254-1|LNC|Shoulder - right MRI W contrast IV|Shoulder - right MRI W contrast IV
C2826012|T102|strict|36255-8|LNC|Sinuses CT W contrast IV|Sinuses CT W contrast IV
C2826012|T102|strict|24915-1|LNC|Sinuses MRI W contrast IV|Sinuses MRI W contrast IV
C2826012|T102|strict|48440-2|LNC|Skull.base MRI W contrast IV|Skull.base MRI W contrast IV
C2826012|T102|strict|37253-2|LNC|Soft tissue MRI W contrast IV|Soft tissue MRI W contrast IV
C2826012|T102|strict|24987-0|LNC|Spine CT W contrast IV|Spine CT W contrast IV
C2826012|T102|strict|36256-6|LNC|Spine MRI W contrast IV|Spine MRI W contrast IV
C2826012|T102|strict|37500-6|LNC|Spine vessels MRI angiogram W contrast IV|Spine vessels MRI angiogram W contrast IV
C2826012|T102|strict|24933-4|LNC|Spine Cervical CT W contrast IV|Spine Cervical CT W contrast IV
C2826012|T102|strict|24938-3|LNC|Spine Cervical MRI W contrast IV|Spine Cervical MRI W contrast IV
C2826012|T102|strict|37501-4|LNC|Cervical Spine vessels MRI angiogram W contrast IV|Cervical Spine vessels MRI angiogram W contrast IV
C2826012|T102|strict|38061-8|LNC|Spine Cervical and Spine Thoracic and Spine Lumbar and Sacrum MRI W contrast IV|Spine Cervical and Spine Thoracic and Spine Lumbar and Sacrum MRI W contrast IV
C2826012|T102|strict|24964-9|LNC|Spine Lumbar CT W contrast IV|Spine Lumbar CT W contrast IV
C2826012|T102|strict|30678-7|LNC|Spine Lumbar MRI W contrast IV|Spine Lumbar MRI W contrast IV
C2826012|T102|strict|37502-2|LNC|Lumbar Spine vessels MRI angiogram W contrast IV|Lumbar Spine vessels MRI angiogram W contrast IV
C2826012|T102|strict|24979-7|LNC|Spine Thoracic CT W contrast IV|Spine Thoracic CT W contrast IV
C2826012|T102|strict|24982-1|LNC|Spine Thoracic MRI W contrast IV|Spine Thoracic MRI W contrast IV
C2826012|T102|strict|37503-0|LNC|Thoracic Spine vessels MRI angiogram W contrast IV|Thoracic Spine vessels MRI angiogram W contrast IV
C2826012|T102|strict|30622-5|LNC|Spleen CT W contrast IV|Spleen CT W contrast IV
C2826012|T102|strict|37242-5|LNC|Sternoclavicular Joint CT W contrast IV|Sternoclavicular Joint CT W contrast IV
C2826012|T102|strict|36257-4|LNC|Sternum CT W contrast IV|Sternum CT W contrast IV
C2826012|T102|strict|36815-9|LNC|Temporal bone CT W contrast IV|Temporal bone CT W contrast IV
C2826012|T102|strict|38835-5|LNC|Temporal bone - left CT W contrast IV|Temporal bone - left CT W contrast IV
C2826012|T102|strict|36816-7|LNC|Temporal bone - right CT W contrast IV|Temporal bone - right CT W contrast IV
C2826012|T102|strict|37243-3|LNC|Temporomandibular joint CT W contrast IV|Temporomandibular joint CT W contrast IV
C2826012|T102|strict|37244-1|LNC|Temporomandibular joint MRI W contrast IV|Temporomandibular joint MRI W contrast IV
C2826012|T102|strict|37245-8|LNC|Temporomandibular joint - bilateral MRI W contrast IV|Temporomandibular joint - bilateral MRI W contrast IV
C2826012|T102|strict|37246-6|LNC|Temporomandibular joint - left CT W contrast IV|Temporomandibular joint - left CT W contrast IV
C2826012|T102|strict|37247-4|LNC|Temporomandibular joint - left MRI W contrast IV|Temporomandibular joint - left MRI W contrast IV
C2826012|T102|strict|37248-2|LNC|Temporomandibular joint - right CT W contrast IV|Temporomandibular joint - right CT W contrast IV
C2826012|T102|strict|37249-0|LNC|Temporomandibular joint - right MRI W contrast IV|Temporomandibular joint - right MRI W contrast IV
C2826012|T102|strict|36173-3|LNC|Thigh MRI W contrast IV|Thigh MRI W contrast IV
C2826012|T102|strict|25003-5|LNC|Thigh vessels MRI angiogram W contrast IV|Thigh vessels MRI angiogram W contrast IV
C2826012|T102|strict|36175-8|LNC|Thigh - left MRI W contrast IV|Thigh - left MRI W contrast IV
C2826012|T102|strict|36177-4|LNC|Thigh - right MRI W contrast IV|Thigh - right MRI W contrast IV
C2826012|T102|strict|36239-2|LNC|Thoracic outlet MRI W contrast IV|Thoracic outlet MRI W contrast IV
C2826012|T102|strict|24584-5|LNC|Thoracic outlet vessels MRI angiogram W contrast IV|Thoracic outlet vessels MRI angiogram W contrast IV
C2826012|T102|strict|26181-8|LNC|Thoracic outlet vessels - bilateral MRI angiogram W contrast IV|Thoracic outlet vessels - bilateral MRI angiogram W contrast IV
C2826012|T102|strict|26182-6|LNC|Thoracic outlet vessels - left MRI angiogram W contrast IV|Thoracic outlet vessels - left MRI angiogram W contrast IV
C2826012|T102|strict|26183-4|LNC|Thoracic outlet vessels - right MRI angiogram W contrast IV|Thoracic outlet vessels - right MRI angiogram W contrast IV
C2826012|T102|strict|36240-0|LNC|Thoracic outlet - left MRI W contrast IV|Thoracic outlet - left MRI W contrast IV
C2826012|T102|strict|36241-8|LNC|Thoracic outlet - right MRI W contrast IV|Thoracic outlet - right MRI W contrast IV
C2826012|T102|strict|72243-9|LNC|Toes - left MRI W contrast IV|Toes - left MRI W contrast IV
C2826012|T102|strict|72240-5|LNC|Toes - right MRI W contrast IV|Toes - right MRI W contrast IV
C2826012|T102|strict|36207-9|LNC|Upper arm CT W contrast IV|Upper arm CT W contrast IV
C2826012|T102|strict|36208-7|LNC|Upper arm MRI W contrast IV|Upper arm MRI W contrast IV
C2826012|T102|strict|69182-4|LNC|Upper arm - bilateral MRI W contrast IV|Upper arm - bilateral MRI W contrast IV
C2826012|T102|strict|36209-5|LNC|Upper arm - left CT W contrast IV|Upper arm - left CT W contrast IV
C2826012|T102|strict|36210-3|LNC|Upper arm - left MRI W contrast IV|Upper arm - left MRI W contrast IV
C2826012|T102|strict|36211-1|LNC|Upper arm - right CT W contrast IV|Upper arm - right CT W contrast IV
C2826012|T102|strict|36212-9|LNC|Upper arm - right MRI W contrast IV|Upper arm - right MRI W contrast IV
C2826012|T102|strict|30626-6|LNC|Upper extremity CT W contrast IV|Upper extremity CT W contrast IV
C2826012|T102|strict|39037-7|LNC|Upper extremity MRI W contrast IV|Upper extremity MRI W contrast IV
C2826012|T102|strict|42295-6|LNC|Upper extremity vessels CT angiogram W contrast IV|Upper extremity vessels CT angiogram W contrast IV
C2826012|T102|strict|24549-8|LNC|Upper extremity vessels MRI angiogram W contrast IV|Upper extremity vessels MRI angiogram W contrast IV
C2826012|T102|strict|36168-3|LNC|Upper extremity - bilateral CT W contrast IV|Upper extremity - bilateral CT W contrast IV
C2826012|T102|strict|69187-3|LNC|Upper extremity - bilateral MRI W contrast IV|Upper extremity - bilateral MRI W contrast IV
C2826012|T102|strict|36216-0|LNC|Upper extremity .joint MRI W contrast IV|Upper extremity .joint MRI W contrast IV
C2826012|T102|strict|36817-5|LNC|Upper extremity joint - bilateral MRI W contrast IV|Upper extremity joint - bilateral MRI W contrast IV
C2826012|T102|strict|36818-3|LNC|Upper extremity joint - left MRI W contrast IV|Upper extremity joint - left MRI W contrast IV
C2826012|T102|strict|36819-1|LNC|Upper extremity joint - right MRI W contrast IV|Upper extremity joint - right MRI W contrast IV
C2826012|T102|strict|36169-1|LNC|Upper extremity - left CT W contrast IV|Upper extremity - left CT W contrast IV
C2826012|T102|strict|38829-8|LNC|Upper extremity - left MRI W contrast IV|Upper extremity - left MRI W contrast IV
C2826012|T102|strict|36170-9|LNC|Upper extremity - right CT W contrast IV|Upper extremity - right CT W contrast IV
C2826012|T102|strict|36171-7|LNC|Upper extremity - right MRI W contrast IV|Upper extremity - right MRI W contrast IV
C2826012|T102|strict|36264-0|LNC|Uterus CT W contrast IV|Uterus CT W contrast IV
C2826012|T102|strict|36265-7|LNC|Uterus MRI W contrast IV|Uterus MRI W contrast IV
C2826012|T102|strict|36834-0|LNC|Vessel CT angiogram W contrast IV|Vessel CT angiogram W contrast IV
C2826012|T102|strict|37447-0|LNC|Wrist CT W contrast IV|Wrist CT W contrast IV
C2826012|T102|strict|37448-8|LNC|Wrist MRI W contrast IV|Wrist MRI W contrast IV
C2826012|T102|strict|69091-7|LNC|Wrist - bilateral CT W contrast IV|Wrist - bilateral CT W contrast IV
C2826012|T102|strict|37449-6|LNC|Wrist - bilateral MRI W contrast IV|Wrist - bilateral MRI W contrast IV
C2826012|T102|strict|37450-4|LNC|Wrist - left CT W contrast IV|Wrist - left CT W contrast IV
C2826012|T102|strict|37451-2|LNC|Wrist - left MRI W contrast IV|Wrist - left MRI W contrast IV
C2826012|T102|strict|37452-0|LNC|Wrist - right CT W contrast IV|Wrist - right CT W contrast IV
C2826012|T102|strict|37453-8|LNC|Wrist - right MRI W contrast IV|Wrist - right MRI W contrast IV
C2826012|T102|strict|24753-6|LNC|Unspecified body region CT W contrast IV|Unspecified body region CT W contrast IV
C2826012|T102|strict|49507-7|LNC|Unspecified body region MRI W contrast IV|Unspecified body region MRI W contrast IV
C2826012|T102|strict|25058-9|LNC|Unspecified body region MRI angiogram W contrast IV|Unspecified body region MRI angiogram W contrast IV
C2826012|T102|strict|72531-7|LNC|Rectum and Colon CT 3D W contrast IV and W air contrast PR|Rectum and Colon CT 3D W contrast IV and W air contrast PR
C2826012|T102|strict|39450-2|LNC|Gastrointestine US W contrast PO|Gastrointestine US W contrast PO
C2826012|T102|strict|72246-2|LNC|Abdomen and Pelvis MRI W contrast PO and W and WO contrast IV|Abdomen and Pelvis MRI W contrast PO and W and WO contrast IV
C2826012|T102|strict|72250-4|LNC|Abdomen and Pelvis CT W contrast PO and W contrast IV|Abdomen and Pelvis CT W contrast PO and W contrast IV
C2826012|T102|strict|72247-0|LNC|Abdomen and Pelvis MRI W contrast PO and WO contrast IV|Abdomen and Pelvis MRI W contrast PO and WO contrast IV
C2826012|T102|strict|72245-4|LNC|Pelvis MRI W contrast PR at rest and maxmal sphincter contraction during straining and defecation|Pelvis MRI W contrast PR at rest and maxmal sphincter contraction during straining and defecation
C2826012|T102|strict|39648-1|LNC|Heart SPECT W dipyridamole and W radionuclide IV|Heart SPECT W dipyridamole and W radionuclide IV
C2826012|T102|strict|44154-3|LNC|Heart SPECT W dipyridamole and W Tc-99m Sestamibi IV|Heart SPECT W dipyridamole and W Tc-99m Sestamibi IV
C2826012|T102|strict|42389-7|LNC|Pelvis MRI W endorectal coil|Pelvis MRI W endorectal coil
C2826012|T102|strict|42388-9|LNC|Prostate MRI W endorectal coil|Prostate MRI W endorectal coil
C2826012|T102|strict|42270-9|LNC|Spine Cervical MRI W flexion and W extension|Spine Cervical MRI W flexion and W extension
C2826012|T102|strict|39682-0|LNC|SPECT W GA-67 IV|SPECT W GA-67 IV
C2826012|T102|strict|39638-2|LNC|Brain SPECT W I-123 IV|Brain SPECT W I-123 IV
C2826012|T102|strict|39755-4|LNC|Thyroid SPECT W I-131 IV|Thyroid SPECT W I-131 IV
C2826012|T102|strict|39839-6|LNC|SPECT W I-131 MIBG IV|SPECT W I-131 MIBG IV
C2826012|T102|strict|39844-6|LNC|SPECT W In-111 Satumomab IV|SPECT W In-111 Satumomab IV
C2826012|T102|strict|41838-4|LNC|Prostate SPECT W In-111 Satumomab IV|Prostate SPECT W In-111 Satumomab IV
C2826012|T102|strict|41772-5|LNC|Bone SPECT W In-111 tagged WBC IV|Bone SPECT W In-111 tagged WBC IV
C2826012|T102|strict|46297-8|LNC|SPECT|SPECT
C2826012|T102|strict|39823-0|LNC|Bone marrow SPECT|Bone marrow SPECT
C2826012|T102|strict|24578-7|LNC|Bones SPECT|Bones SPECT
C2826012|T102|strict|39632-5|LNC|Brain SPECT|Brain SPECT
C2826012|T102|strict|39644-0|LNC|Breast SPECT|Breast SPECT
C2826012|T102|strict|39770-3|LNC|Gastrointestine SPECT|Gastrointestine SPECT
C2826012|T102|strict|39649-9|LNC|Heart SPECT|Heart SPECT
C2826012|T102|strict|42310-3|LNC|Kidney SPECT|Kidney SPECT
C2826012|T102|strict|39852-9|LNC|Kidney - bilateral SPECT|Kidney - bilateral SPECT
C2826012|T102|strict|39692-9|LNC|Liver SPECT|Liver SPECT
C2826012|T102|strict|39876-8|LNC|Liver and Spleen SPECT|Liver and Spleen SPECT
C2826012|T102|strict|39628-3|LNC|Meckels diverticulum SPECT|Meckels diverticulum SPECT
C2826012|T102|strict|39740-6|LNC|Parathyroid SPECT|Parathyroid SPECT
C2826012|T102|strict|43526-3|LNC|Unspecified body region SPECT|Unspecified body region SPECT
C2826012|T102|strict|39938-6|LNC|Joint SPECT|Joint SPECT
C2826012|T102|strict|46330-7|LNC|Abdomen CT W reduced contrast volume IV|Abdomen CT W reduced contrast volume IV
C2826012|T102|strict|46327-3|LNC|Chest CT W reduced contrast volume IV|Chest CT W reduced contrast volume IV
C2826012|T102|strict|46326-5|LNC|Facial bones and Maxilla CT W reduced contrast volume IV|Facial bones and Maxilla CT W reduced contrast volume IV
C2826012|T102|strict|46328-1|LNC|Head CT W reduced contrast volume IV|Head CT W reduced contrast volume IV
C2826012|T102|strict|46325-7|LNC|Internal auditory canal CT W reduced contrast volume IV|Internal auditory canal CT W reduced contrast volume IV
C2826012|T102|strict|46329-9|LNC|Pelvis CT W reduced contrast volume IV|Pelvis CT W reduced contrast volume IV
C2826012|T102|strict|42143-8|LNC|Uterus and Fallopian tubes US W saline intrauterine|Uterus and Fallopian tubes US W saline intrauterine
C2826012|T102|strict|58750-1|LNC|Heart MRI W stress|Heart MRI W stress
C2826012|T102|strict|58749-3|LNC|Heart MRI W stress and W and WO contrast IV|Heart MRI W stress and W and WO contrast IV
C2826012|T102|strict|39668-9|LNC|Heart SPECT W stress and W radionuclide IV|Heart SPECT W stress and W radionuclide IV
C2826012|T102|strict|44152-7|LNC|Brain SPECT W Tc-99m bicisate IV|Brain SPECT W Tc-99m bicisate IV
C2826012|T102|strict|39743-0|LNC|Prostate SPECT W Tc-99m capromab pendatide IV|Prostate SPECT W Tc-99m capromab pendatide IV
C2826012|T102|strict|39640-8|LNC|Brain SPECT W Tc-99m DTPA IV|Brain SPECT W Tc-99m DTPA IV
C2826012|T102|strict|39641-6|LNC|Brain SPECT W Tc-99m glucoheptonate IV|Brain SPECT W Tc-99m glucoheptonate IV
C2826012|T102|strict|44153-5|LNC|Kidney SPECT W Tc-99m glucoheptonate IV|Kidney SPECT W Tc-99m glucoheptonate IV
C2826012|T102|strict|39631-7|LNC|Brain SPECT W Tc-99m HMPAO IV|Brain SPECT W Tc-99m HMPAO IV
C2826012|T102|strict|24817-9|LNC|Liver SPECT W Tc-99m IV|Liver SPECT W Tc-99m IV
C2826012|T102|strict|39851-1|LNC|Kidney - bilateral SPECT W Tc-99m Mertiatide IV|Kidney - bilateral SPECT W Tc-99m Mertiatide IV
C2826012|T102|strict|69229-3|LNC|Liver SPECT W Tc-99m SC IV|Liver SPECT W Tc-99m SC IV
C2826012|T102|strict|44151-9|LNC|Heart SPECT W Tc-99m Sestamibi IV|Heart SPECT W Tc-99m Sestamibi IV
C2826012|T102|strict|39691-1|LNC|Liver SPECT W Tc-99m tagged RBC IV|Liver SPECT W Tc-99m tagged RBC IV
C2826012|T102|strict|69234-3|LNC|Spleen SPECT W Tc-99m tagged RBC IV|Spleen SPECT W Tc-99m tagged RBC IV
C2826012|T102|strict|39647-3|LNC|Heart SPECT W Tc-99m Tetrofosmin IV|Heart SPECT W Tc-99m Tetrofosmin IV
C2826012|T102|strict|39639-0|LNC|Brain SPECT W Tl-201 IV|Brain SPECT W Tl-201 IV
C2826012|T102|strict|42377-2|LNC|Brain CT W Xe-133 inhaled|Brain CT W Xe-133 inhaled
C2826012|T102|strict|46393-5|LNC|Liver CT W Xe-133 inhaled|Liver CT W Xe-133 inhaled
C2826012|T102|strict|42394-7|LNC|Pulmonary system CT W Xe-133 inhaled|Pulmonary system CT W Xe-133 inhaled
C2826012|T102|strict|36424-0|LNC|Abdomen CT WO contrast|Abdomen CT WO contrast
C2826012|T102|strict|30668-8|LNC|Abdomen MRI WO contrast|Abdomen MRI WO contrast
C2826012|T102|strict|42291-5|LNC|Abdomen retroperitoneum CT WO contrast|Abdomen retroperitoneum CT WO contrast
C2826012|T102|strict|36952-0|LNC|Abdomen and Pelvis CT WO contrast|Abdomen and Pelvis CT WO contrast
C2826012|T102|strict|36878-7|LNC|Abdominal vessels MRI angiogram WO contrast|Abdominal vessels MRI angiogram WO contrast
C2826012|T102|strict|36496-8|LNC|Acromioclavicular Joint MRI WO contrast|Acromioclavicular Joint MRI WO contrast
C2826012|T102|strict|36953-8|LNC|Adrenal gland CT WO contrast|Adrenal gland CT WO contrast
C2826012|T102|strict|36954-6|LNC|Adrenal gland MRI WO contrast|Adrenal gland MRI WO contrast
C2826012|T102|strict|36425-7|LNC|Ankle CT WO contrast|Ankle CT WO contrast
C2826012|T102|strict|30680-3|LNC|Ankle MRI WO contrast|Ankle MRI WO contrast
C2826012|T102|strict|36879-5|LNC|Ankle vessels MRI angiogram WO contrast|Ankle vessels MRI angiogram WO contrast
C2826012|T102|strict|69087-5|LNC|Ankle - bilateral CT WO contrast|Ankle - bilateral CT WO contrast
C2826012|T102|strict|69164-2|LNC|Ankle - bilateral MRI WO contrast|Ankle - bilateral MRI WO contrast
C2826012|T102|strict|36426-5|LNC|Ankle - left CT WO contrast|Ankle - left CT WO contrast
C2826012|T102|strict|36427-3|LNC|Ankle - left MRI WO contrast|Ankle - left MRI WO contrast
C2826012|T102|strict|36428-1|LNC|Ankle - right CT WO contrast|Ankle - right CT WO contrast
C2826012|T102|strict|36429-9|LNC|Ankle - right MRI WO contrast|Ankle - right MRI WO contrast
C2826012|T102|strict|36430-7|LNC|Aorta CT WO contrast|Aorta CT WO contrast
C2826012|T102|strict|44132-9|LNC|Aorta MRI angiogram WO contrast|Aorta MRI angiogram WO contrast
C2826012|T102|strict|36431-5|LNC|Aorta abdominal CT WO contrast|Aorta abdominal CT WO contrast
C2826012|T102|strict|36432-3|LNC|Aorta abdominal MRI angiogram WO contrast|Aorta abdominal MRI angiogram WO contrast
C2826012|T102|strict|69119-6|LNC|Aorta thoracic CT angiogram WO contrast|Aorta thoracic CT angiogram WO contrast
C2826012|T102|strict|36433-1|LNC|Aorta thoracic MRI angiogram WO contrast|Aorta thoracic MRI angiogram WO contrast
C2826012|T102|strict|44130-3|LNC|Aortic arch MRI angiogram WO contrast|Aortic arch MRI angiogram WO contrast
C2826012|T102|strict|36434-9|LNC|Appendix CT WO contrast|Appendix CT WO contrast
C2826012|T102|strict|44123-8|LNC|Biliary ducts and Pancreatic duct MRI WO contrast|Biliary ducts and Pancreatic duct MRI WO contrast
C2826012|T102|strict|30657-1|LNC|Brain MRI WO contrast|Brain MRI WO contrast
C2826012|T102|strict|48453-5|LNC|Brain.temporal MRI WO contrast|Brain.temporal MRI WO contrast
C2826012|T102|strict|37278-9|LNC|Brain and Internal auditory canal MRI WO contrast|Brain and Internal auditory canal MRI WO contrast
C2826012|T102|strict|37279-7|LNC|Brain and Larynx MRI WO contrast|Brain and Larynx MRI WO contrast
C2826012|T102|strict|42393-9|LNC|Brain and Pituitary and Sella turcica MRI WO contrast|Brain and Pituitary and Sella turcica MRI WO contrast
C2826012|T102|strict|36436-4|LNC|Breast MRI WO contrast|Breast MRI WO contrast
C2826012|T102|strict|69191-5|LNC|Breast implant MRI WO contrast|Breast implant MRI WO contrast
C2826012|T102|strict|69168-3|LNC|Breast implant - bilateral MRI WO contrast|Breast implant - bilateral MRI WO contrast
C2826012|T102|strict|38064-2|LNC|Breast implant - left MRI WO contrast|Breast implant - left MRI WO contrast
C2826012|T102|strict|38817-3|LNC|Breast implant - right MRI WO contrast|Breast implant - right MRI WO contrast
C2826012|T102|strict|44119-6|LNC|Breast - bilateral CT WO contrast|Breast - bilateral CT WO contrast
C2826012|T102|strict|36437-2|LNC|Breast - bilateral MRI WO contrast|Breast - bilateral MRI WO contrast
C2826012|T102|strict|36438-0|LNC|Breast - left MRI WO contrast|Breast - left MRI WO contrast
C2826012|T102|strict|36439-8|LNC|Breast - right MRI WO contrast|Breast - right MRI WO contrast
C2826012|T102|strict|46333-1|LNC|Breast - unilateral MRI WO contrast|Breast - unilateral MRI WO contrast
C2826012|T102|strict|36483-6|LNC|Calcaneus CT WO contrast|Calcaneus CT WO contrast
C2826012|T102|strict|36440-6|LNC|Calcaneus - left CT WO contrast|Calcaneus - left CT WO contrast
C2826012|T102|strict|36441-4|LNC|Calcaneus - right CT WO contrast|Calcaneus - right CT WO contrast
C2826012|T102|strict|36880-3|LNC|Carotid vessel MRI angiogram WO contrast|Carotid vessel MRI angiogram WO contrast
C2826012|T102|strict|29252-4|LNC|Chest CT WO contrast|Chest CT WO contrast
C2826012|T102|strict|36442-2|LNC|Chest MRI WO contrast|Chest MRI WO contrast
C2826012|T102|strict|69084-2|LNC|Chest vessels CT angiogram WO contrast|Chest vessels CT angiogram WO contrast
C2826012|T102|strict|36547-8|LNC|Chest vessels MRI angiogram WO contrast|Chest vessels MRI angiogram WO contrast
C2826012|T102|strict|42276-6|LNC|Chest and Abdomen CT WO contrast|Chest and Abdomen CT WO contrast
C2826012|T102|strict|72253-8|LNC|Chest and Abdomen and Pelvis CT WO contrast|Chest and Abdomen and Pelvis CT WO contrast
C2826012|T102|strict|42302-0|LNC|Clavicle MRI WO contrast|Clavicle MRI WO contrast
C2826012|T102|strict|48459-2|LNC|Clavicle - left MRI WO contrast|Clavicle - left MRI WO contrast
C2826012|T102|strict|48458-4|LNC|Clavicle - right MRI WO contrast|Clavicle - right MRI WO contrast
C2826012|T102|strict|36443-0|LNC|Elbow CT WO contrast|Elbow CT WO contrast
C2826012|T102|strict|30796-7|LNC|Elbow MRI WO contrast|Elbow MRI WO contrast
C2826012|T102|strict|36444-8|LNC|Elbow - bilateral CT WO contrast|Elbow - bilateral CT WO contrast
C2826012|T102|strict|69171-7|LNC|Elbow - bilateral MRI WO contrast|Elbow - bilateral MRI WO contrast
C2826012|T102|strict|36445-5|LNC|Elbow - left CT WO contrast|Elbow - left CT WO contrast
C2826012|T102|strict|36446-3|LNC|Elbow - left MRI WO contrast|Elbow - left MRI WO contrast
C2826012|T102|strict|36447-1|LNC|Elbow - right CT WO contrast|Elbow - right CT WO contrast
C2826012|T102|strict|36448-9|LNC|Elbow - right MRI WO contrast|Elbow - right MRI WO contrast
C2826012|T102|strict|42278-2|LNC|Extremity CT WO contrast|Extremity CT WO contrast
C2826012|T102|strict|69104-8|LNC|Extremity - left CT WO contrast|Extremity - left CT WO contrast
C2826012|T102|strict|69111-3|LNC|Extremity - right CT WO contrast|Extremity - right CT WO contrast
C2826012|T102|strict|36435-6|LNC|Face MRI WO contrast|Face MRI WO contrast
C2826012|T102|strict|30802-3|LNC|Facial bones and Maxilla CT WO contrast|Facial bones and Maxilla CT WO contrast
C2826012|T102|strict|72249-6|LNC|Facial bones and Sinuses CT WO contrast|Facial bones and Sinuses CT WO contrast
C2826012|T102|strict|36460-4|LNC|Femur CT WO contrast|Femur CT WO contrast
C2826012|T102|strict|69173-3|LNC|Femur - bilateral MRI WO contrast|Femur - bilateral MRI WO contrast
C2826012|T102|strict|36462-0|LNC|Femur - left CT WO contrast|Femur - left CT WO contrast
C2826012|T102|strict|36464-6|LNC|Femur - right CT WO contrast|Femur - right CT WO contrast
C2826012|T102|strict|69196-4|LNC|Finger MRI WO contrast|Finger MRI WO contrast
C2826012|T102|strict|69206-1|LNC|Finger - left MRI WO contrast|Finger - left MRI WO contrast
C2826012|T102|strict|69216-0|LNC|Finger - right MRI WO contrast|Finger - right MRI WO contrast
C2826012|T102|strict|36466-1|LNC|Foot CT WO contrast|Foot CT WO contrast
C2826012|T102|strict|30681-1|LNC|Foot MRI WO contrast|Foot MRI WO contrast
C2826012|T102|strict|36467-9|LNC|Foot - bilateral MRI WO contrast|Foot - bilateral MRI WO contrast
C2826012|T102|strict|36468-7|LNC|Foot - left CT WO contrast|Foot - left CT WO contrast
C2826012|T102|strict|36469-5|LNC|Foot - left MRI WO contrast|Foot - left MRI WO contrast
C2826012|T102|strict|36470-3|LNC|Foot - right CT WO contrast|Foot - right CT WO contrast
C2826012|T102|strict|36471-1|LNC|Foot - right MRI WO contrast|Foot - right MRI WO contrast
C2826012|T102|strict|36472-9|LNC|Forearm CT WO contrast|Forearm CT WO contrast
C2826012|T102|strict|30683-7|LNC|Forearm MRI WO contrast|Forearm MRI WO contrast
C2826012|T102|strict|69176-6|LNC|Forearm - bilateral MRI WO contrast|Forearm - bilateral MRI WO contrast
C2826012|T102|strict|36473-7|LNC|Forearm - left CT WO contrast|Forearm - left CT WO contrast
C2826012|T102|strict|36474-5|LNC|Forearm - left MRI WO contrast|Forearm - left MRI WO contrast
C2826012|T102|strict|36475-2|LNC|Forearm - right CT WO contrast|Forearm - right CT WO contrast
C2826012|T102|strict|36476-0|LNC|Forearm - right MRI WO contrast|Forearm - right MRI WO contrast
C2826012|T102|strict|36477-8|LNC|Hand CT WO contrast|Hand CT WO contrast
C2826012|T102|strict|30685-2|LNC|Hand MRI WO contrast|Hand MRI WO contrast
C2826012|T102|strict|69179-0|LNC|Hand - bilateral MRI WO contrast|Hand - bilateral MRI WO contrast
C2826012|T102|strict|36478-6|LNC|Hand - left CT WO contrast|Hand - left CT WO contrast
C2826012|T102|strict|36479-4|LNC|Hand - left MRI WO contrast|Hand - left MRI WO contrast
C2826012|T102|strict|36480-2|LNC|Hand - right CT WO contrast|Hand - right CT WO contrast
C2826012|T102|strict|36481-0|LNC|Hand - right MRI WO contrast|Hand - right MRI WO contrast
C2826012|T102|strict|30799-1|LNC|Head CT WO contrast|Head CT WO contrast
C2826012|T102|strict|36876-1|LNC|Head veins MRI angiogram WO contrast|Head veins MRI angiogram WO contrast
C2826012|T102|strict|42293-1|LNC|Head vessels CT angiogram WO contrast|Head vessels CT angiogram WO contrast
C2826012|T102|strict|36881-1|LNC|Head vessels MRI angiogram WO contrast|Head vessels MRI angiogram WO contrast
C2826012|T102|strict|36482-8|LNC|Heart MRI WO contrast|Heart MRI WO contrast
C2826012|T102|strict|36484-4|LNC|Hip CT WO contrast|Hip CT WO contrast
C2826012|T102|strict|30687-8|LNC|Hip MRI WO contrast|Hip MRI WO contrast
C2826012|T102|strict|36485-1|LNC|Hip - bilateral CT WO contrast|Hip - bilateral CT WO contrast
C2826012|T102|strict|36486-9|LNC|Hip - bilateral MRI WO contrast|Hip - bilateral MRI WO contrast
C2826012|T102|strict|36487-7|LNC|Hip - left CT WO contrast|Hip - left CT WO contrast
C2826012|T102|strict|36488-5|LNC|Hip - left MRI WO contrast|Hip - left MRI WO contrast
C2826012|T102|strict|36489-3|LNC|Hip - right CT WO contrast|Hip - right CT WO contrast
C2826012|T102|strict|36490-1|LNC|Hip - right MRI WO contrast|Hip - right MRI WO contrast
C2826012|T102|strict|30584-7|LNC|Internal auditory canal CT WO contrast|Internal auditory canal CT WO contrast
C2826012|T102|strict|30658-9|LNC|Internal auditory canal MRI WO contrast|Internal auditory canal MRI WO contrast
C2826012|T102|strict|43770-7|LNC|Kidney CT WO contrast|Kidney CT WO contrast
C2826012|T102|strict|43773-1|LNC|Kidney MRI WO contrast|Kidney MRI WO contrast
C2826012|T102|strict|36503-1|LNC|Kidney - bilateral CT WO contrast|Kidney - bilateral CT WO contrast
C2826012|T102|strict|36504-9|LNC|Kidney - bilateral MRI WO contrast|Kidney - bilateral MRI WO contrast
C2826012|T102|strict|39359-5|LNC|Kidney - bilateral X-ray tomograph WO contrast|Kidney - bilateral X-ray tomograph WO contrast
C2826012|T102|strict|36505-6|LNC|Knee CT WO contrast|Knee CT WO contrast
C2826012|T102|strict|30691-0|LNC|Knee MRI WO contrast|Knee MRI WO contrast
C2826012|T102|strict|69089-1|LNC|Knee - bilateral CT WO contrast|Knee - bilateral CT WO contrast
C2826012|T102|strict|36506-4|LNC|Knee - bilateral MRI WO contrast|Knee - bilateral MRI WO contrast
C2826012|T102|strict|36507-2|LNC|Knee - left CT WO contrast|Knee - left CT WO contrast
C2826012|T102|strict|36508-0|LNC|Knee - left MRI WO contrast|Knee - left MRI WO contrast
C2826012|T102|strict|36509-8|LNC|Knee - right CT WO contrast|Knee - right CT WO contrast
C2826012|T102|strict|36510-6|LNC|Knee - right MRI WO contrast|Knee - right MRI WO contrast
C2826012|T102|strict|36511-4|LNC|Larynx CT WO contrast|Larynx CT WO contrast
C2826012|T102|strict|48445-1|LNC|Larynx MRI WO contrast|Larynx MRI WO contrast
C2826012|T102|strict|30611-8|LNC|Liver CT WO contrast|Liver CT WO contrast
C2826012|T102|strict|30669-6|LNC|Liver MRI WO contrast|Liver MRI WO contrast
C2826012|T102|strict|30625-8|LNC|Lower extremity CT WO contrast|Lower extremity CT WO contrast
C2826012|T102|strict|39292-8|LNC|Lower extremity MRI WO contrast|Lower extremity MRI WO contrast
C2826012|T102|strict|44129-5|LNC|Lower extremity vessels MRI angiogram WO contrast|Lower extremity vessels MRI angiogram WO contrast
C2826012|T102|strict|36450-5|LNC|Lower extremity vessels - bilateral MRI angiogram WO contrast|Lower extremity vessels - bilateral MRI angiogram WO contrast
C2826012|T102|strict|36882-9|LNC|Lower extremity vessels - left MRI angiogram WO contrast|Lower extremity vessels - left MRI angiogram WO contrast
C2826012|T102|strict|38773-8|LNC|Lower extremity vessels - right MRI angiogram WO contrast|Lower extremity vessels - right MRI angiogram WO contrast
C2826012|T102|strict|36449-7|LNC|Lower extremity - bilateral CT WO contrast|Lower extremity - bilateral CT WO contrast
C2826012|T102|strict|36451-3|LNC|Lower extremity - bilateral MRI WO contrast|Lower extremity - bilateral MRI WO contrast
C2826012|T102|strict|36497-6|LNC|Lower Extremity Joint MRI WO contrast|Lower Extremity Joint MRI WO contrast
C2826012|T102|strict|36498-4|LNC|Lower extremity joint - left MRI WO contrast|Lower extremity joint - left MRI WO contrast
C2826012|T102|strict|36499-2|LNC|Lower extremity joint - right MRI WO contrast|Lower extremity joint - right MRI WO contrast
C2826012|T102|strict|36452-1|LNC|Lower extremity - left CT WO contrast|Lower extremity - left CT WO contrast
C2826012|T102|strict|36453-9|LNC|Lower extremity - left MRI WO contrast|Lower extremity - left MRI WO contrast
C2826012|T102|strict|36454-7|LNC|Lower extremity - right CT WO contrast|Lower extremity - right CT WO contrast
C2826012|T102|strict|36455-4|LNC|Lower extremity - right MRI WO contrast|Lower extremity - right MRI WO contrast
C2826012|T102|strict|36537-9|LNC|Lower leg CT WO contrast|Lower leg CT WO contrast
C2826012|T102|strict|30869-2|LNC|Lower leg MRI WO contrast|Lower leg MRI WO contrast
C2826012|T102|strict|69185-7|LNC|Lower leg - bilateral MRI WO contrast|Lower leg - bilateral MRI WO contrast
C2826012|T102|strict|36538-7|LNC|Lower leg - left CT WO contrast|Lower leg - left CT WO contrast
C2826012|T102|strict|36539-5|LNC|Lower leg - left MRI WO contrast|Lower leg - left MRI WO contrast
C2826012|T102|strict|36540-3|LNC|Lower leg - right CT WO contrast|Lower leg - right CT WO contrast
C2826012|T102|strict|36541-1|LNC|Lower leg - right MRI WO contrast|Lower leg - right MRI WO contrast
C2826012|T102|strict|36512-2|LNC|Mandible CT WO contrast|Mandible CT WO contrast
C2826012|T102|strict|36513-0|LNC|Nasopharynx MRI WO contrast|Nasopharynx MRI WO contrast
C2826012|T102|strict|30585-4|LNC|Nasopharynx and Neck CT WO contrast|Nasopharynx and Neck CT WO contrast
C2826012|T102|strict|36514-8|LNC|Neck CT WO contrast|Neck CT WO contrast
C2826012|T102|strict|30660-5|LNC|Neck MRI WO contrast|Neck MRI WO contrast
C2826012|T102|strict|36877-9|LNC|Neck veins MRI angiogram WO contrast|Neck veins MRI angiogram WO contrast
C2826012|T102|strict|36549-4|LNC|Neck vessels MRI angiogram WO contrast|Neck vessels MRI angiogram WO contrast
C2826012|T102|strict|46331-5|LNC|Orbit CT WO contrast|Orbit CT WO contrast
C2826012|T102|strict|36872-0|LNC|Orbit MRI WO contrast|Orbit MRI WO contrast
C2826012|T102|strict|30587-0|LNC|Orbit - bilateral CT WO contrast|Orbit - bilateral CT WO contrast
C2826012|T102|strict|30661-3|LNC|Orbit - bilateral MRI WO contrast|Orbit - bilateral MRI WO contrast
C2826012|T102|strict|36873-8|LNC|Orbit - left MRI WO contrast|Orbit - left MRI WO contrast
C2826012|T102|strict|36874-6|LNC|Orbit - right MRI WO contrast|Orbit - right MRI WO contrast
C2826012|T102|strict|36956-1|LNC|Orbit and Face MRI WO contrast|Orbit and Face MRI WO contrast
C2826012|T102|strict|46332-3|LNC|Orbit and Face and Neck MRI WO contrast|Orbit and Face and Neck MRI WO contrast
C2826012|T102|strict|36875-3|LNC|Ovary MRI WO contrast|Ovary MRI WO contrast
C2826012|T102|strict|30613-4|LNC|Pancreas CT WO contrast|Pancreas CT WO contrast
C2826012|T102|strict|36515-5|LNC|Pancreas MRI WO contrast|Pancreas MRI WO contrast
C2826012|T102|strict|37280-5|LNC|Parotid gland CT WO contrast|Parotid gland CT WO contrast
C2826012|T102|strict|37281-3|LNC|Parotid gland MRI WO contrast|Parotid gland MRI WO contrast
C2826012|T102|strict|30615-9|LNC|Pelvis CT WO contrast|Pelvis CT WO contrast
C2826012|T102|strict|30673-8|LNC|Pelvis MRI WO contrast|Pelvis MRI WO contrast
C2826012|T102|strict|36883-7|LNC|Pelvis vessels MRI angiogram WO contrast|Pelvis vessels MRI angiogram WO contrast
C2826012|T102|strict|30671-2|LNC|Pelvis and Hip MRI WO contrast|Pelvis and Hip MRI WO contrast
C2826012|T102|strict|30589-6|LNC|Petrous bone CT WO contrast|Petrous bone CT WO contrast
C2826012|T102|strict|30591-2|LNC|Pituitary and Sella turcica CT WO contrast|Pituitary and Sella turcica CT WO contrast
C2826012|T102|strict|30666-2|LNC|Pituitary and Sella turcica MRI WO contrast|Pituitary and Sella turcica MRI WO contrast
C2826012|T102|strict|36543-7|LNC|Portal vein MRI angiogram WO contrast|Portal vein MRI angiogram WO contrast
C2826012|T102|strict|36517-1|LNC|Posterior fossa CT WO contrast|Posterior fossa CT WO contrast
C2826012|T102|strict|36518-9|LNC|Posterior fossa MRI WO contrast|Posterior fossa MRI WO contrast
C2826012|T102|strict|36519-7|LNC|Prostate MRI WO contrast|Prostate MRI WO contrast
C2826012|T102|strict|36544-5|LNC|Renal vein MRI angiogram WO contrast|Renal vein MRI angiogram WO contrast
C2826012|T102|strict|44133-7|LNC|Renal vessels MRI angiogram WO contrast|Renal vessels MRI angiogram WO contrast
C2826012|T102|strict|36501-5|LNC|Sacroiliac Joint CT WO contrast|Sacroiliac Joint CT WO contrast
C2826012|T102|strict|36502-3|LNC|Sacroiliac Joint MRI WO contrast|Sacroiliac Joint MRI WO contrast
C2826012|T102|strict|36520-5|LNC|Sacrum CT WO contrast|Sacrum CT WO contrast
C2826012|T102|strict|36521-3|LNC|Sacrum MRI WO contrast|Sacrum MRI WO contrast
C2826012|T102|strict|36522-1|LNC|Sacrum and Coccyx MRI WO contrast|Sacrum and Coccyx MRI WO contrast
C2826012|T102|strict|69118-8|LNC|Scapula CT WO contrast|Scapula CT WO contrast
C2826012|T102|strict|36523-9|LNC|Scapula - left MRI WO contrast|Scapula - left MRI WO contrast
C2826012|T102|strict|38770-4|LNC|Scapula - right MRI WO contrast|Scapula - right MRI WO contrast
C2826012|T102|strict|36535-3|LNC|Scrotum and Testicle MRI WO contrast|Scrotum and Testicle MRI WO contrast
C2826012|T102|strict|36524-7|LNC|Shoulder CT WO contrast|Shoulder CT WO contrast
C2826012|T102|strict|30693-6|LNC|Shoulder MRI WO contrast|Shoulder MRI WO contrast
C2826012|T102|strict|69090-9|LNC|Shoulder - bilateral CT WO contrast|Shoulder - bilateral CT WO contrast
C2826012|T102|strict|36525-4|LNC|Shoulder - bilateral MRI WO contrast|Shoulder - bilateral MRI WO contrast
C2826012|T102|strict|36526-2|LNC|Shoulder - left CT WO contrast|Shoulder - left CT WO contrast
C2826012|T102|strict|38834-8|LNC|Shoulder - left MRI WO contrast|Shoulder - left MRI WO contrast
C2826012|T102|strict|36527-0|LNC|Shoulder - right CT WO contrast|Shoulder - right CT WO contrast
C2826012|T102|strict|36528-8|LNC|Shoulder - right MRI WO contrast|Shoulder - right MRI WO contrast
C2826012|T102|strict|36529-6|LNC|Sinuses CT WO contrast|Sinuses CT WO contrast
C2826012|T102|strict|30662-1|LNC|Sinuses MRI WO contrast|Sinuses MRI WO contrast
C2826012|T102|strict|44112-1|LNC|Skull.base CT WO contrast|Skull.base CT WO contrast
C2826012|T102|strict|48687-8|LNC|Skull.base MRI WO contrast|Skull.base MRI WO contrast
C2826012|T102|strict|37293-8|LNC|Soft tissue MRI WO contrast|Soft tissue MRI WO contrast
C2826012|T102|strict|36530-4|LNC|Spine CT WO contrast|Spine CT WO contrast
C2826012|T102|strict|36531-2|LNC|Spine MRI WO contrast|Spine MRI WO contrast
C2826012|T102|strict|37510-5|LNC|Spine vessels MRI angiogram WO contrast|Spine vessels MRI angiogram WO contrast
C2826012|T102|strict|30592-0|LNC|Spine Cervical CT WO contrast|Spine Cervical CT WO contrast
C2826012|T102|strict|30667-0|LNC|Spine Cervical MRI WO contrast|Spine Cervical MRI WO contrast
C2826012|T102|strict|37511-3|LNC|Cervical Spine vessels MRI angiogram WO contrast|Cervical Spine vessels MRI angiogram WO contrast
C2826012|T102|strict|30854-4|LNC|Spine Cervical and Thoracic and Lumbar MRI WO contrast|Spine Cervical and Thoracic and Lumbar MRI WO contrast
C2826012|T102|strict|30620-9|LNC|Spine Lumbar CT WO contrast|Spine Lumbar CT WO contrast
C2826012|T102|strict|30679-5|LNC|Spine Lumbar MRI WO contrast|Spine Lumbar MRI WO contrast
C2826012|T102|strict|37994-1|LNC|Lumbar Spine vessels MRI angiogram WO contrast|Lumbar Spine vessels MRI angiogram WO contrast
C2826012|T102|strict|37288-8|LNC|Spine Lumbosacral Junction CT WO contrast|Spine Lumbosacral Junction CT WO contrast
C2826012|T102|strict|30597-9|LNC|Spine Thoracic CT WO contrast|Spine Thoracic CT WO contrast
C2826012|T102|strict|36532-0|LNC|Spine Thoracic MRI WO contrast|Spine Thoracic MRI WO contrast
C2826012|T102|strict|37512-1|LNC|Thoracic Spine vessels MRI angiogram WO contrast|Thoracic Spine vessels MRI angiogram WO contrast
C2826012|T102|strict|30621-7|LNC|Spleen CT WO contrast|Spleen CT WO contrast
C2826012|T102|strict|36533-8|LNC|Spleen MRI WO contrast|Spleen MRI WO contrast
C2826012|T102|strict|37282-1|LNC|Sternoclavicular Joint CT WO contrast|Sternoclavicular Joint CT WO contrast
C2826012|T102|strict|36534-6|LNC|Sternum CT WO contrast|Sternum CT WO contrast
C2826012|T102|strict|44230-1|LNC|Superior mesenteric vessels MRI angiogram WO contrast|Superior mesenteric vessels MRI angiogram WO contrast
C2826012|T102|strict|36866-2|LNC|Temporal bone CT WO contrast|Temporal bone CT WO contrast
C2826012|T102|strict|36867-0|LNC|Temporal bone - left CT WO contrast|Temporal bone - left CT WO contrast
C2826012|T102|strict|36868-8|LNC|Temporal bone - right CT WO contrast|Temporal bone - right CT WO contrast
C2826012|T102|strict|37283-9|LNC|Temporomandibular joint CT WO contrast|Temporomandibular joint CT WO contrast
C2826012|T102|strict|37284-7|LNC|Temporomandibular joint MRI WO contrast|Temporomandibular joint MRI WO contrast
C2826012|T102|strict|37285-4|LNC|Temporomandibular joint - bilateral MRI WO contrast|Temporomandibular joint - bilateral MRI WO contrast
C2826012|T102|strict|37286-2|LNC|Temporomandibular joint - left MRI WO contrast|Temporomandibular joint - left MRI WO contrast
C2826012|T102|strict|37287-0|LNC|Temporomandibular joint - right MRI WO contrast|Temporomandibular joint - right MRI WO contrast
C2826012|T102|strict|36461-2|LNC|Thigh MRI WO contrast|Thigh MRI WO contrast
C2826012|T102|strict|43514-9|LNC|Thigh vessels - left MRI angiogram WO contrast|Thigh vessels - left MRI angiogram WO contrast
C2826012|T102|strict|43515-6|LNC|Thigh vessels - right MRI angiogram WO contrast|Thigh vessels - right MRI angiogram WO contrast
C2826012|T102|strict|36463-8|LNC|Thigh - left MRI WO contrast|Thigh - left MRI WO contrast
C2826012|T102|strict|36465-3|LNC|Thigh - right MRI WO contrast|Thigh - right MRI WO contrast
C2826012|T102|strict|30654-8|LNC|Thoracic outlet MRI WO contrast|Thoracic outlet MRI WO contrast
C2826012|T102|strict|38833-0|LNC|Thoracic outlet - left MRI WO contrast|Thoracic outlet - left MRI WO contrast
C2826012|T102|strict|36516-3|LNC|Thoracic outlet - right MRI WO contrast|Thoracic outlet - right MRI WO contrast
C2826012|T102|strict|36955-3|LNC|Thyroid CT WO contrast|Thyroid CT WO contrast
C2826012|T102|strict|36536-1|LNC|Thyroid MRI WO contrast|Thyroid MRI WO contrast
C2826012|T102|strict|72242-1|LNC|Toes - left MRI WO contrast|Toes - left MRI WO contrast
C2826012|T102|strict|72239-7|LNC|Toes - right MRI WO contrast|Toes - right MRI WO contrast
C2826012|T102|strict|36491-9|LNC|Upper arm CT WO contrast|Upper arm CT WO contrast
C2826012|T102|strict|30689-4|LNC|Upper arm MRI WO contrast|Upper arm MRI WO contrast
C2826012|T102|strict|69183-2|LNC|Upper arm - bilateral MRI WO contrast|Upper arm - bilateral MRI WO contrast
C2826012|T102|strict|36492-7|LNC|Upper arm - left CT WO contrast|Upper arm - left CT WO contrast
C2826012|T102|strict|36493-5|LNC|Upper arm - left MRI WO contrast|Upper arm - left MRI WO contrast
C2826012|T102|strict|36494-3|LNC|Upper arm - right CT WO contrast|Upper arm - right CT WO contrast
C2826012|T102|strict|36495-0|LNC|Upper arm - right MRI WO contrast|Upper arm - right MRI WO contrast
C2826012|T102|strict|30627-4|LNC|Upper extremity CT WO contrast|Upper extremity CT WO contrast
C2826012|T102|strict|39033-6|LNC|Upper extremity MRI WO contrast|Upper extremity MRI WO contrast
C2826012|T102|strict|36548-6|LNC|Upper extremity vessels MRI angiogram WO contrast|Upper extremity vessels MRI angiogram WO contrast
C2826012|T102|strict|36456-2|LNC|Upper extremity - bilateral CT WO contrast|Upper extremity - bilateral CT WO contrast
C2826012|T102|strict|69188-1|LNC|Upper extremity - bilateral MRI WO contrast|Upper extremity - bilateral MRI WO contrast
C2826012|T102|strict|36500-7|LNC|Upper extremity .joint MRI WO contrast|Upper extremity .joint MRI WO contrast
C2826012|T102|strict|36869-6|LNC|Upper extremity joint - left MRI WO contrast|Upper extremity joint - left MRI WO contrast
C2826012|T102|strict|36870-4|LNC|Upper extremity joint - right MRI WO contrast|Upper extremity joint - right MRI WO contrast
C2826012|T102|strict|36457-0|LNC|Upper extremity - left CT WO contrast|Upper extremity - left CT WO contrast
C2826012|T102|strict|38832-2|LNC|Upper extremity - left MRI WO contrast|Upper extremity - left MRI WO contrast
C2826012|T102|strict|36458-8|LNC|Upper extremity - right CT WO contrast|Upper extremity - right CT WO contrast
C2826012|T102|strict|36459-6|LNC|Upper extremity - right MRI WO contrast|Upper extremity - right MRI WO contrast
C2826012|T102|strict|36542-9|LNC|Uterus MRI WO contrast|Uterus MRI WO contrast
C2826012|T102|strict|36545-2|LNC|Inferior vena cava MRI WO contrast|Inferior vena cava MRI WO contrast
C2826012|T102|strict|36546-0|LNC|Superior vena cava MRI WO contrast|Superior vena cava MRI WO contrast
C2826012|T102|strict|37459-5|LNC|Wrist CT WO contrast|Wrist CT WO contrast
C2826012|T102|strict|37460-3|LNC|Wrist MRI WO contrast|Wrist MRI WO contrast
C2826012|T102|strict|43516-4|LNC|Wrist vessels - left MRI angiogram WO contrast|Wrist vessels - left MRI angiogram WO contrast
C2826012|T102|strict|43517-2|LNC|Wrist vessels - right MRI angiogram WO contrast|Wrist vessels - right MRI angiogram WO contrast
C2826012|T102|strict|37461-1|LNC|Wrist - bilateral CT WO contrast|Wrist - bilateral CT WO contrast
C2826012|T102|strict|37462-9|LNC|Wrist - bilateral MRI WO contrast|Wrist - bilateral MRI WO contrast
C2826012|T102|strict|37463-7|LNC|Wrist - left CT WO contrast|Wrist - left CT WO contrast
C2826012|T102|strict|37464-5|LNC|Wrist - left MRI WO contrast|Wrist - left MRI WO contrast
C2826012|T102|strict|37465-2|LNC|Wrist - right CT WO contrast|Wrist - right CT WO contrast
C2826012|T102|strict|37466-0|LNC|Wrist - right MRI WO contrast|Wrist - right MRI WO contrast
C2826012|T102|strict|43525-5|LNC|Unspecified body region CT WO contrast|Unspecified body region CT WO contrast
C2826012|T102|strict|69223-6|LNC|Unspecified body region MRI WO contrast|Unspecified body region MRI WO contrast
C2826012|T102|strict|36871-2|LNC|Joint MRI WO contrast|Joint MRI WO contrast
C2826012|T102|strict|24787-4|LNC|Kidney - bilateral X-ray tomograph WO contrast and 10M post contrast IV|Kidney - bilateral X-ray tomograph WO contrast and 10M post contrast IV
C2826012|T102|strict|30712-4|LNC|Hip US WO developmental joint assessment|Hip US WO developmental joint assessment
C2826012|T102|strict|25051-4|LNC|Unspecified body region CT Multisectional sagittal|Unspecified body region CT Multisectional sagittal
C2826012|T102|strict|29750-7|LNC|Neonatal intensive care records|Neonatal intensive care records
C2826012|T102|strict|25060-5|LNC|Unspecified body region US No charge|Unspecified body region US No charge
C2826012|T102|strict|52072-6|LNC|Non-emergency transportation|Non-emergency transportation
C2826012|T102|strict|53246-5|LNC|Non-medical services|Non-medical services
C2826012|T102|strict|46210-1|LNC|Case manager Note|Case manager Note
C2826012|T102|strict|34819-3|LNC|Pathology Evaluation and management note|Pathology Evaluation and management note
C2826012|T102|strict|46215-0|LNC|Wound care management Note|Wound care management Note
C2826012|T102|strict|28568-4|LNC|Physician Emergency department Note|Physician Emergency department Note
C2826012|T102|strict|11536-0|LNC|Nurse Notes|Nurse Notes
C2826012|T102|strict|52066-8|LNC|Notice of Discharge Medicare Appeal Rights (NODMAR) form|Notice of Discharge Medicare Appeal Rights (NODMAR) form
C2826012|T102|strict|53244-0|LNC|Notice of privacy practices receipt|Notice of privacy practices receipt
C2826012|T102|strict|11543-6|LNC|Nursery records|Nursery records
C2826012|T102|strict|46208-5|LNC|Nursing notes|Nursing notes
C2826012|T102|strict|52051-0|LNC|Orthotics/Prosthetics|Orthotics/Prosthetics
C2826012|T102|strict|52052-8|LNC|Osteogenesis stimulators|Osteogenesis stimulators
C2826012|T102|strict|52053-6|LNC|Oxygen|Oxygen
C2826012|T102|strict|52054-4|LNC|Parenteral|Parenteral
C2826012|T102|strict|52067-6|LNC|Past filing limit justification|Past filing limit justification
C2826012|T102|strict|24620-7|LNC|Catheter Fluoroscopy Patency check W contrast via catheter|Catheter Fluoroscopy Patency check W contrast via catheter
C2826012|T102|strict|33721-2|LNC|Bone marrow Pathology biopsy report|Bone marrow Pathology biopsy report
C2826012|T102|strict|34122-2|LNC|Pathology procedure note|Pathology procedure note
C2826012|T102|strict|55188-7|LNC|Patient data Document|Patient data Document
C2826012|T102|strict|55750-4|LNC|Patient safety report Event Document|Patient safety report Event Document
C2826012|T102|strict|52034-6|LNC|Payer letter|Payer letter
C2826012|T102|strict|24882-3|LNC|Popliteal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA|Popliteal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA
C2826012|T102|strict|69252-5|LNC|Pulmonary artery Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA|Pulmonary artery Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA
C2826012|T102|strict|69248-3|LNC|Renal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA|Renal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA
C2826012|T102|strict|42018-2|LNC|Vein Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA|Vein Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA
C2826012|T102|strict|69301-0|LNC|Upper extremity vein Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IV|Upper extremity vein Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IV
C2826012|T102|strict|28629-4|LNC|Perimetry study|Perimetry study
C2826012|T102|strict|74030-8|LNC|Periodontal service attachment|Periodontal service attachment
C2826012|T102|strict|29752-3|LNC|Perioperative records|Perioperative records
C2826012|T102|strict|24875-7|LNC|Peripheral vessel US.doppler Peripheral plane|Peripheral vessel US.doppler Peripheral plane
C2826012|T102|strict|51965-2|LNC|Pharmacogenetic analysis report in Blood or Tissue Document by Molecular genetics method|Pharmacogenetic analysis report in Blood or Tissue Document by Molecular genetics method
C2826012|T102|strict|51850-6|LNC|Physical findings of Head and Ears and Eyes and Nose and Throat|Physical findings of Head and Ears and Eyes and Nose and Throat
C2826012|T102|strict|24998-7|LNC|Placement check of gastrostomy tube W contrast via GI tube|Placement check of gastrostomy tube W contrast via GI tube
C2826012|T102|strict|52055-1|LNC|Power operated vehicles|Power operated vehicles
C2826012|T102|strict|52063-5|LNC|Prescription for durable medical equipment (DME)|Prescription for durable medical equipment (DME)
C2826012|T102|strict|18836-7|LNC|Cardiac stress study Procedure|Cardiac stress study Procedure
C2826012|T102|strict|28570-0|LNC|Provider-unspecified Procedure note|Provider-unspecified Procedure note
C2826012|T102|strict|28577-5|LNC|Dentist procedure note|Dentist procedure note
C2826012|T102|strict|11505-5|LNC|Physician procedure note|Physician procedure note
C2826012|T102|strict|28625-2|LNC|Podiatry procedure note|Podiatry procedure note
C2826012|T102|strict|52068-4|LNC|Property and casualty state mandated forms|Property and casualty state mandated forms
C2826012|T102|strict|46209-3|LNC|Provider orders|Provider orders
C2826012|T102|strict|55751-2|LNC|Public health case report Document|Public health case report Document
C2826012|T102|strict|52075-9|LNC|Purchase invoice|Purchase invoice
C2826012|T102|strict|55184-6|LNC|Quality Reporting Document Architecture calculated summary report population Document|Quality Reporting Document Architecture calculated summary report population Document
C2826012|T102|strict|55182-0|LNC|Quality Reporting Document Architecture incidence report Document|Quality Reporting Document Architecture incidence report Document
C2826012|T102|strict|55183-8|LNC|Quality Reporting Document Architecture patient list report population Document|Quality Reporting Document Architecture patient list report population Document
C2826012|T102|strict|62385-0|LNC|Recommendation [interpretation] Document|Recommendation [interpretation] Document
C2826012|T102|strict|11514-7|LNC|Chiropractic Records total Encounter|Chiropractic Records total Encounter
C2826012|T102|strict|11521-2|LNC|Occupational therapy Records total Encounter|Occupational therapy Records total Encounter
C2826012|T102|strict|11515-4|LNC|Physical therapy Records total Encounter|Physical therapy Records total Encounter
C2826012|T102|strict|11516-2|LNC|Physician Records total Encounter|Physician Records total Encounter
C2826012|T102|strict|11517-0|LNC|Podiatry Records total Encounter|Podiatry Records total Encounter
C2826012|T102|strict|11518-8|LNC|Psychology Records total Encounter|Psychology Records total Encounter
C2826012|T102|strict|11519-6|LNC|Social service Records total Encounter|Social service Records total Encounter
C2826012|T102|strict|11520-4|LNC|Speech therapy Records total Encounter|Speech therapy Records total Encounter
C2826012|T102|strict|44226-9|LNC|Colon Fluoroscopy Reduction W views W barium contrast PR|Colon Fluoroscopy Reduction W views W barium contrast PR
C2826012|T102|strict|30636-5|LNC|Colon Fluoroscopy Reduction W views W contrast PR|Colon Fluoroscopy Reduction W views W contrast PR
C2826012|T102|strict|18823-5|LNC|Alcohol and/or substance abuse service attachment|Alcohol and/or substance abuse service attachment
C2826012|T102|strict|18824-3|LNC|Cardiac service attachment|Cardiac service attachment
C2826012|T102|strict|18825-0|LNC|Medical social services attachment|Medical social services attachment
C2826012|T102|strict|18826-8|LNC|Occupational therapy service attachment|Occupational therapy service attachment
C2826012|T102|strict|19002-5|LNC|Physical therapy service attachment|Physical therapy service attachment
C2826012|T102|strict|18594-2|LNC|Psychiatric service attachment|Psychiatric service attachment
C2826012|T102|strict|52184-9|LNC|Pulmonary therapy service attachment|Pulmonary therapy service attachment
C2826012|T102|strict|19003-3|LNC|Respiratory therapy service attachment|Respiratory therapy service attachment
C2826012|T102|strict|19004-1|LNC|Skilled nursing service attachment|Skilled nursing service attachment
C2826012|T102|strict|29206-0|LNC|Speech therapy service attachment|Speech therapy service attachment
C2826012|T102|strict|25073-8|LNC|Vessel Fluoroscopic angiogram Removal of foreign body from vascular space|Vessel Fluoroscopic angiogram Removal of foreign body from vascular space
C2826012|T102|strict|52056-9|LNC|Repair of durable medical equipment|Repair of durable medical equipment
C2826012|T102|strict|25015-9|LNC|Upper GI tract Replacement of percutaneous gastrojejunostomy|Upper GI tract Replacement of percutaneous gastrojejunostomy
C2826012|T102|strict|60569-1|LNC|Report addendum.synoptic Document|Report addendum.synoptic Document
C2826012|T102|strict|55187-9|LNC|Reporting parameters Document|Reporting parameters Document
C2826012|T102|strict|52057-7|LNC|Seat lift mechanism|Seat lift mechanism
C2826012|T102|strict|52058-5|LNC|Seating systems|Seating systems
C2826012|T102|strict|52039-5|LNC|Skilled Nursing Facility (SNF) record|Skilled Nursing Facility (SNF) record
C2826012|T102|strict|52059-3|LNC|Speech generating device|Speech generating device
C2826012|T102|strict|52060-1|LNC|Standers/standing frames|Standers/standing frames
C2826012|T102|strict|52029-6|LNC|Sterilization consent|Sterilization consent
C2826012|T102|strict|55228-1|LNC|Cytogenetics study|Cytogenetics study
C2826012|T102|strict|18752-6|LNC|Exercise stress test study|Exercise stress test study
C2826012|T102|strict|29755-6|LNC|Nerve conduction study|Nerve conduction study
C2826012|T102|strict|11526-1|LNC|Pathology study|Pathology study
C2826012|T102|strict|28633-6|LNC|Polysomnography (sleep) study|Polysomnography (sleep) study
C2826012|T102|strict|11527-9|LNC|Psychiatry study|Psychiatry study
C2826012|T102|strict|58477-1|LNC|Pulmonary function report|Pulmonary function report
C2826012|T102|strict|11529-5|LNC|Surgical pathology study|Surgical pathology study
C2826012|T102|strict|55230-7|LNC|Immunophenotyping study|Immunophenotyping study
C2826012|T102|strict|11523-8|LNC|EEG study|EEG study
C2826012|T102|strict|11541-0|LNC|MRI Brain study|MRI Brain study
C2826012|T102|strict|29757-2|LNC|Colposcopy study|Colposcopy study
C2826012|T102|strict|33717-0|LNC|Cytology Cervical or vaginal smear or scraping study|Cytology Cervical or vaginal smear or scraping study
C2826012|T102|strict|18745-0|LNC|Cardiac catheterization study|Cardiac catheterization study
C2826012|T102|strict|11524-6|LNC|EKG study|EKG study
C2826012|T102|strict|18750-0|LNC|Electrophysiology study|Electrophysiology study
C2826012|T102|strict|18754-2|LNC|Holter monitor study|Holter monitor study
C2826012|T102|strict|18746-8|LNC|Colonoscopy study|Colonoscopy study
C2826012|T102|strict|18753-4|LNC|Flexible sigmoidoscopy study|Flexible sigmoidoscopy study
C2826012|T102|strict|29756-4|LNC|Peritoneoscopy study|Peritoneoscopy study
C2826012|T102|strict|18744-3|LNC|Bronchoscopy study|Bronchoscopy study
C2826012|T102|strict|18759-1|LNC|Spirometry study|Spirometry study
C2826012|T102|strict|38269-7|LNC|Study report Skeletal system DXA|Study report Skeletal system DXA
C2826012|T102|strict|18756-7|LNC|MRI Spine study|MRI Spine study
C2826012|T102|strict|17787-3|LNC|Thyroid Scan Study report|Thyroid Scan Study report
C2826012|T102|strict|55229-9|LNC|Immune stain study|Immune stain study
C2826012|T102|strict|18751-8|LNC|Endoscopy study|Endoscopy study
C2826012|T102|strict|18742-7|LNC|Arthroscopy study|Arthroscopy study
C2826012|T102|strict|33716-2|LNC|Non-gynecological cytology method study|Non-gynecological cytology method study
C2826012|T102|strict|18748-4|LNC|Diagnostic imaging study|Diagnostic imaging study
C2826012|T102|strict|18749-2|LNC|Electromyogram study|Electromyogram study
C2826012|T102|strict|33719-6|LNC|Flow cytometry study|Flow cytometry study
C2826012|T102|strict|29754-9|LNC|Nystagmogram study|Nystagmogram study
C2826012|T102|strict|52038-7|LNC|Subscriber Information including retroactive and presumptive eligibility|Subscriber Information including retroactive and presumptive eligibility
C2826012|T102|strict|52061-9|LNC|Support surfaces|Support surfaces
C2826012|T102|strict|28583-3|LNC|Dentist Operation note|Dentist Operation note
C2826012|T102|strict|28573-4|LNC|Physician, Operation note|Physician, Operation note
C2826012|T102|strict|60568-3|LNC|Synoptic report|Synoptic report
C2826012|T102|strict|52069-2|LNC|Tax ID number - IRS form W9|Tax ID number - IRS form W9
C2826012|T102|strict|11534-5|LNC|Temperature charts|Temperature charts
C2826012|T102|strict|46213-5|LNC|Tilt table study|Tilt table study
C2826012|T102|strict|28630-2|LNC|Tonometry study|Tonometry study
C2826012|T102|strict|52062-7|LNC|Transcutaneous electrical neural stimulation (TENS)|Transcutaneous electrical neural stimulation (TENS)
C2826012|T102|strict|28651-8|LNC|Nurse Transfer note|Nurse Transfer note
C2826012|T102|strict|28616-1|LNC|Physician Transfer note|Physician Transfer note
C2826012|T102|strict|69409-1|LNC|U.S. standard certificate of death - 2003 revision|U.S. standard certificate of death - 2003 revision
C2826012|T102|strict|24783-3|LNC|Kidney - bilateral Fluoroscopy Urodynamics|Kidney - bilateral Fluoroscopy Urodynamics
C2826012|T102|strict|25065-4|LNC|Unspecified body region Fluoroscopy 15 minutes|Unspecified body region Fluoroscopy 15 minutes
C2826012|T102|strict|25068-8|LNC|Unspecified body region Fluoroscopy 1 hour|Unspecified body region Fluoroscopy 1 hour
C2826012|T102|strict|43471-2|LNC|Unspecified body region Fluoroscopy 2 hour|Unspecified body region Fluoroscopy 2 hour
C2826012|T102|strict|25066-2|LNC|Unspecified body region Fluoroscopy 30 minutes|Unspecified body region Fluoroscopy 30 minutes
C2826012|T102|strict|25067-0|LNC|Unspecified body region Fluoroscopy 45 minutes|Unspecified body region Fluoroscopy 45 minutes
C2826012|T102|strict|43472-0|LNC|Unspecified body region Fluoroscopy 90 minutes|Unspecified body region Fluoroscopy 90 minutes
C2826012|T102|strict|42702-1|LNC|Unspecified body region Fluoroscopy Greater than 1 hour|Unspecified body region Fluoroscopy Greater than 1 hour
C2826012|T102|strict|42703-9|LNC|Unspecified body region Fluoroscopy Less than 1 hour|Unspecified body region Fluoroscopy Less than 1 hour
C2826012|T102|strict|36550-2|LNC|Abdomen X-ray Single view|Abdomen X-ray Single view
C2826012|T102|strict|36551-0|LNC|Ankle X-ray Single view|Ankle X-ray Single view
C2826012|T102|strict|69307-7|LNC|Ankle - left X-ray Single view|Ankle - left X-ray Single view
C2826012|T102|strict|69314-3|LNC|Ankle - right X-ray Single view|Ankle - right X-ray Single view
C2826012|T102|strict|46335-6|LNC|Breast - bilateral Mammogram Single view|Breast - bilateral Mammogram Single view
C2826012|T102|strict|46336-4|LNC|Breast - left Mammogram Single view|Breast - left Mammogram Single view
C2826012|T102|strict|46337-2|LNC|Breast - right Mammogram Single view|Breast - right Mammogram Single view
C2826012|T102|strict|46338-0|LNC|Breast - unilateral Mammogram Single view|Breast - unilateral Mammogram Single view
C2826012|T102|strict|36564-3|LNC|Calcaneus X-ray Single view|Calcaneus X-ray Single view
C2826012|T102|strict|69311-9|LNC|Calcaneus - left X-ray Single view|Calcaneus - left X-ray Single view
C2826012|T102|strict|69319-2|LNC|Calcaneus - right X-ray Single view|Calcaneus - right X-ray Single view
C2826012|T102|strict|36554-4|LNC|Chest X-ray Single view|Chest X-ray Single view
C2826012|T102|strict|42699-9|LNC|Chest and Abdomen X-ray Single view|Chest and Abdomen X-ray Single view
C2826012|T102|strict|36555-1|LNC|Clavicle X-ray Single view|Clavicle X-ray Single view
C2826012|T102|strict|36556-9|LNC|Elbow X-ray Single view|Elbow X-ray Single view
C2826012|T102|strict|69308-5|LNC|Elbow - left X-ray Single view|Elbow - left X-ray Single view
C2826012|T102|strict|69315-0|LNC|Elbow - right X-ray Single view|Elbow - right X-ray Single view
C2826012|T102|strict|42153-7|LNC|Extremity X-ray Single view|Extremity X-ray Single view
C2826012|T102|strict|36559-3|LNC|Femur X-ray Single view|Femur X-ray Single view
C2826012|T102|strict|36560-1|LNC|Femur - left X-ray Single view|Femur - left X-ray Single view
C2826012|T102|strict|37689-7|LNC|Femur - right X-ray Single view|Femur - right X-ray Single view
C2826012|T102|strict|36561-9|LNC|Foot X-ray Single view|Foot X-ray Single view
C2826012|T102|strict|69309-3|LNC|Foot - left X-ray Single view|Foot - left X-ray Single view
C2826012|T102|strict|69316-8|LNC|Foot - right X-ray Single view|Foot - right X-ray Single view
C2826012|T102|strict|36563-5|LNC|Hand X-ray Single view|Hand X-ray Single view
C2826012|T102|strict|69310-1|LNC|Hand - left X-ray Single view|Hand - left X-ray Single view
C2826012|T102|strict|69318-4|LNC|Hand - right X-ray Single view|Hand - right X-ray Single view
C2826012|T102|strict|24761-9|LNC|Hip X-ray Single view|Hip X-ray Single view
C2826012|T102|strict|26400-2|LNC|Hip - bilateral X-ray Single view|Hip - bilateral X-ray Single view
C2826012|T102|strict|26401-0|LNC|Hip - left X-ray Single view|Hip - left X-ray Single view
C2826012|T102|strict|26402-8|LNC|Hip - right X-ray Single view|Hip - right X-ray Single view
C2826012|T102|strict|36565-0|LNC|Humerus X-ray Single view|Humerus X-ray Single view
C2826012|T102|strict|69312-7|LNC|Humerus - left X-ray Single view|Humerus - left X-ray Single view
C2826012|T102|strict|69320-0|LNC|Humerus - right X-ray Single view|Humerus - right X-ray Single view
C2826012|T102|strict|36566-8|LNC|Knee - bilateral X-ray Single view|Knee - bilateral X-ray Single view
C2826012|T102|strict|36567-6|LNC|Knee - left X-ray Single view|Knee - left X-ray Single view
C2826012|T102|strict|37741-6|LNC|Knee - right X-ray Single view|Knee - right X-ray Single view
C2826012|T102|strict|36557-7|LNC|Lower extremity - bilateral X-ray Single view|Lower extremity - bilateral X-ray Single view
C2826012|T102|strict|36558-5|LNC|Lower extremity - left X-ray Single view|Lower extremity - left X-ray Single view
C2826012|T102|strict|37764-8|LNC|Lower extremity - right X-ray Single view|Lower extremity - right X-ray Single view
C2826012|T102|strict|37614-5|LNC|Patella X-ray Single view|Patella X-ray Single view
C2826012|T102|strict|69152-7|LNC|Patella - left X-ray Single view|Patella - left X-ray Single view
C2826012|T102|strict|69260-8|LNC|Patella - right X-ray Single view|Patella - right X-ray Single view
C2826012|T102|strict|37616-0|LNC|Pelvis X-ray Single view|Pelvis X-ray Single view
C2826012|T102|strict|69317-6|LNC|Radius - right and Ulna - right X-ray Single view|Radius - right and Ulna - right X-ray Single view
C2826012|T102|strict|42313-7|LNC|Ribs - left X-ray Single view|Ribs - left X-ray Single view
C2826012|T102|strict|42314-5|LNC|Ribs - right X-ray Single view|Ribs - right X-ray Single view
C2826012|T102|strict|37654-1|LNC|Scapula X-ray Single view|Scapula X-ray Single view
C2826012|T102|strict|30748-8|LNC|Shoulder X-ray Single view|Shoulder X-ray Single view
C2826012|T102|strict|36568-4|LNC|Shoulder - bilateral X-ray Single view|Shoulder - bilateral X-ray Single view
C2826012|T102|strict|36569-2|LNC|Shoulder - left X-ray Single view|Shoulder - left X-ray Single view
C2826012|T102|strict|37792-9|LNC|Shoulder - right X-ray Single view|Shoulder - right X-ray Single view
C2826012|T102|strict|37851-3|LNC|Sinuses X-ray Single view|Sinuses X-ray Single view
C2826012|T102|strict|24917-7|LNC|Skull X-ray Single view|Skull X-ray Single view
C2826012|T102|strict|48695-1|LNC|Skull.base X-ray Single view|Skull.base X-ray Single view
C2826012|T102|strict|37875-2|LNC|Spine X-ray Single view|Spine X-ray Single view
C2826012|T102|strict|24940-9|LNC|Spine Cervical X-ray Single view|Spine Cervical X-ray Single view
C2826012|T102|strict|30773-6|LNC|Spine Lumbar X-ray Single view|Spine Lumbar X-ray Single view
C2826012|T102|strict|37904-0|LNC|Spine Thoracic X-ray Single view|Spine Thoracic X-ray Single view
C2826012|T102|strict|38121-0|LNC|Spine Thoracic and Lumbar X-ray Single view|Spine Thoracic and Lumbar X-ray Single view
C2826012|T102|strict|69313-5|LNC|Tibia - left and Fibula - left X-ray Single view|Tibia - left and Fibula - left X-ray Single view
C2826012|T102|strict|69321-8|LNC|Tibia - right and Fibula - right X-ray Single view|Tibia - right and Fibula - right X-ray Single view
C2826012|T102|strict|37894-3|LNC|Tibia and Fibula X-ray Single view|Tibia and Fibula X-ray Single view
C2826012|T102|strict|37924-8|LNC|Wrist X-ray Single view|Wrist X-ray Single view
C2826012|T102|strict|42419-2|LNC|Wrist - bilateral X-ray Single view|Wrist - bilateral X-ray Single view
C2826012|T102|strict|36570-0|LNC|Wrist - left X-ray Single view|Wrist - left X-ray Single view
C2826012|T102|strict|37825-7|LNC|Wrist - right X-ray Single view|Wrist - right X-ray Single view
C2826012|T102|strict|30642-3|LNC|Unspecified body region Fluoroscopy Single view|Unspecified body region Fluoroscopy Single view
C2826012|T102|strict|30787-6|LNC|Joint X-ray Single view|Joint X-ray Single view
C2826012|T102|strict|44176-6|LNC|Hip X-ray Single view portable|Hip X-ray Single view portable
C2826012|T102|strict|41775-8|LNC|Pelvis X-ray Single view portable|Pelvis X-ray Single view portable
C2826012|T102|strict|30749-6|LNC|Shoulder X-ray Single view portable|Shoulder X-ray Single view portable
C2826012|T102|strict|30722-3|LNC|Skull X-ray Single view portable|Skull X-ray Single view portable
C2826012|T102|strict|30724-9|LNC|Spine Cervical X-ray Single view portable|Spine Cervical X-ray Single view portable
C2826012|T102|strict|30774-4|LNC|Spine Lumbar X-ray Single view portable|Spine Lumbar X-ray Single view portable
C2826012|T102|strict|70932-9|LNC|Spine Thoracic X-ray Single view portable|Spine Thoracic X-ray Single view portable
C2826012|T102|strict|25063-9|LNC|Vessel Fluoroscopic angiogram Single view W contrast IA|Vessel Fluoroscopic angiogram Single view W contrast IA
C2826012|T102|strict|69268-1|LNC|Breast duct Mammogram Single view W contrast intra duct|Breast duct Mammogram Single view W contrast intra duct
C2826012|T102|strict|49510-1|LNC|Breast duct - left Mammogram Single view W contrast intra duct|Breast duct - left Mammogram Single view W contrast intra duct
C2826012|T102|strict|49509-3|LNC|Breast duct - right Mammogram Single view W contrast intra duct|Breast duct - right Mammogram Single view W contrast intra duct
C2826012|T102|strict|24715-5|LNC|Gastrointestine upper Fluoroscopy Single view W contrast PO|Gastrointestine upper Fluoroscopy Single view W contrast PO
C2826012|T102|strict|37513-9|LNC|Tibia - bilateral X-ray 10 degree caudal angle|Tibia - bilateral X-ray 10 degree caudal angle
C2826012|T102|strict|37514-7|LNC|Tibia - left X-ray 10 degree caudal angle|Tibia - left X-ray 10 degree caudal angle
C2826012|T102|strict|38806-6|LNC|Tibia - right X-ray 10 degree caudal angle|Tibia - right X-ray 10 degree caudal angle
C2826012|T102|strict|37467-8|LNC|Acromioclavicular Joint X-ray 10 degree cephalic angle|Acromioclavicular Joint X-ray 10 degree cephalic angle
C2826012|T102|strict|37468-6|LNC|Shoulder - bilateral X-ray 30 degree caudal angle|Shoulder - bilateral X-ray 30 degree caudal angle
C2826012|T102|strict|42431-7|LNC|Knee - right X-ray 30 degree standing|Knee - right X-ray 30 degree standing
C2826012|T102|strict|69079-2|LNC|Clavicle X-ray 45 degree cephalic angle|Clavicle X-ray 45 degree cephalic angle
C2826012|T102|strict|37469-4|LNC|Clavicle - bilateral X-ray 45 degree cephalic angle|Clavicle - bilateral X-ray 45 degree cephalic angle
C2826012|T102|strict|37470-2|LNC|Clavicle - left X-ray 45 degree cephalic angle|Clavicle - left X-ray 45 degree cephalic angle
C2826012|T102|strict|38803-3|LNC|Clavicle - right X-ray 45 degree cephalic angle|Clavicle - right X-ray 45 degree cephalic angle
C2826012|T102|strict|24799-9|LNC|Abdomen X-ray AP single view|Abdomen X-ray AP single view
C2826012|T102|strict|36583-3|LNC|Acromioclavicular joint - left X-ray AP single view|Acromioclavicular joint - left X-ray AP single view
C2826012|T102|strict|37662-4|LNC|Acromioclavicular joint - right X-ray AP single view|Acromioclavicular joint - right X-ray AP single view
C2826012|T102|strict|36571-8|LNC|Ankle X-ray AP single view|Ankle X-ray AP single view
C2826012|T102|strict|36572-6|LNC|Chest X-ray AP single view|Chest X-ray AP single view
C2826012|T102|strict|36573-4|LNC|Clavicle X-ray AP single view|Clavicle X-ray AP single view
C2826012|T102|strict|36575-9|LNC|Femur X-ray AP single view|Femur X-ray AP single view
C2826012|T102|strict|36576-7|LNC|Finger fifth X-ray AP single view|Finger fifth X-ray AP single view
C2826012|T102|strict|36577-5|LNC|Finger fourth X-ray AP single view|Finger fourth X-ray AP single view
C2826012|T102|strict|36578-3|LNC|Finger third X-ray AP single view|Finger third X-ray AP single view
C2826012|T102|strict|36579-1|LNC|Foot X-ray AP single view|Foot X-ray AP single view
C2826012|T102|strict|36580-9|LNC|Foot - bilateral X-ray AP single view|Foot - bilateral X-ray AP single view
C2826012|T102|strict|36581-7|LNC|Hip X-ray AP single view|Hip X-ray AP single view
C2826012|T102|strict|36582-5|LNC|Hip - left X-ray AP single view|Hip - left X-ray AP single view
C2826012|T102|strict|37726-7|LNC|Hip - right X-ray AP single view|Hip - right X-ray AP single view
C2826012|T102|strict|36584-1|LNC|Knee X-ray AP single view|Knee X-ray AP single view
C2826012|T102|strict|36585-8|LNC|Knee - bilateral X-ray AP single view|Knee - bilateral X-ray AP single view
C2826012|T102|strict|48462-6|LNC|Knee - left X-ray AP single view|Knee - left X-ray AP single view
C2826012|T102|strict|48463-4|LNC|Knee - right X-ray AP single view|Knee - right X-ray AP single view
C2826012|T102|strict|36574-2|LNC|Lower extremity X-ray AP single view|Lower extremity X-ray AP single view
C2826012|T102|strict|42439-0|LNC|Neck X-ray AP single view|Neck X-ray AP single view
C2826012|T102|strict|37622-8|LNC|Pelvis X-ray AP single view|Pelvis X-ray AP single view
C2826012|T102|strict|39050-0|LNC|Ribs X-ray AP single view|Ribs X-ray AP single view
C2826012|T102|strict|36958-7|LNC|Ribs - bilateral X-ray AP single view|Ribs - bilateral X-ray AP single view
C2826012|T102|strict|36959-5|LNC|Ribs - left X-ray AP single view|Ribs - left X-ray AP single view
C2826012|T102|strict|37783-8|LNC|Ribs - right X-ray AP single view|Ribs - right X-ray AP single view
C2826012|T102|strict|39048-4|LNC|Scapula X-ray AP single view|Scapula X-ray AP single view
C2826012|T102|strict|37842-2|LNC|Shoulder X-ray AP single view|Shoulder X-ray AP single view
C2826012|T102|strict|36586-6|LNC|Shoulder - bilateral X-ray AP single view|Shoulder - bilateral X-ray AP single view
C2826012|T102|strict|36587-4|LNC|Shoulder - left X-ray AP single view|Shoulder - left X-ray AP single view
C2826012|T102|strict|37798-6|LNC|Shoulder - right X-ray AP single view|Shoulder - right X-ray AP single view
C2826012|T102|strict|69269-9|LNC|Skull X-ray AP single view|Skull X-ray AP single view
C2826012|T102|strict|37877-8|LNC|Spine X-ray AP single view|Spine X-ray AP single view
C2826012|T102|strict|30725-6|LNC|Spine Cervical X-ray AP single view|Spine Cervical X-ray AP single view
C2826012|T102|strict|24948-2|LNC|Spine Cervical Odontoid and Cervical axis X-ray AP single view|Spine Cervical Odontoid and Cervical axis X-ray AP single view
C2826012|T102|strict|30777-7|LNC|Spine Lumbar X-ray AP single view|Spine Lumbar X-ray AP single view
C2826012|T102|strict|30752-0|LNC|Spine Thoracic X-ray AP single view|Spine Thoracic X-ray AP single view
C2826012|T102|strict|39049-2|LNC|Spine Thoracic and Lumbar X-ray AP single view|Spine Thoracic and Lumbar X-ray AP single view
C2826012|T102|strict|37880-2|LNC|Sternoclavicular Joint X-ray AP single view|Sternoclavicular Joint X-ray AP single view
C2826012|T102|strict|37890-1|LNC|Thumb X-ray AP single view|Thumb X-ray AP single view
C2826012|T102|strict|37897-6|LNC|Tibia and Fibula X-ray AP single view|Tibia and Fibula X-ray AP single view
C2826012|T102|strict|39402-3|LNC|Shoulder X-ray AP (W internal rotation and W external rotation)|Shoulder X-ray AP (W internal rotation and W external rotation)
C2826012|T102|strict|37634-3|LNC|Pelvis X-ray AP 20 degree cephalic angle|Pelvis X-ray AP 20 degree cephalic angle
C2826012|T102|strict|30734-8|LNC|Chest X-ray AP lateral-decubitus|Chest X-ray AP lateral-decubitus
C2826012|T102|strict|30735-5|LNC|Chest X-ray AP lateral-decubitus portable|Chest X-ray AP lateral-decubitus portable
C2826012|T102|strict|24561-3|LNC|Abdomen X-ray AP left lateral-decubitus|Abdomen X-ray AP left lateral-decubitus
C2826012|T102|strict|24637-1|LNC|Chest X-ray AP left lateral-decubitus|Chest X-ray AP left lateral-decubitus
C2826012|T102|strict|24560-5|LNC|Abdomen X-ray AP left lateral-decubitus portable|Abdomen X-ray AP left lateral-decubitus portable
C2826012|T102|strict|24636-3|LNC|Chest X-ray AP left lateral-decubitus portable|Chest X-ray AP left lateral-decubitus portable
C2826012|T102|strict|36588-2|LNC|Abdomen X-ray AP portable single view|Abdomen X-ray AP portable single view
C2826012|T102|strict|36589-0|LNC|Chest X-ray AP portable single view|Chest X-ray AP portable single view
C2826012|T102|strict|30727-2|LNC|Spine Cervical X-ray AP portable single view|Spine Cervical X-ray AP portable single view
C2826012|T102|strict|30729-8|LNC|Spine Cervical Odontoid and Cervical axis X-ray AP portable single view|Spine Cervical Odontoid and Cervical axis X-ray AP portable single view
C2826012|T102|strict|30755-3|LNC|Spine Thoracic X-ray AP portable single view|Spine Thoracic X-ray AP portable single view
C2826012|T102|strict|24563-9|LNC|Abdomen X-ray AP right lateral-decubitus|Abdomen X-ray AP right lateral-decubitus
C2826012|T102|strict|43466-2|LNC|Chest X-ray AP right lateral-decubitus|Chest X-ray AP right lateral-decubitus
C2826012|T102|strict|24652-0|LNC|Chest X-ray AP right lateral-decubitus portable|Chest X-ray AP right lateral-decubitus portable
C2826012|T102|strict|43778-0|LNC|Chest X-ray AP supine portable|Chest X-ray AP supine portable
C2826012|T102|strict|24564-7|LNC|Abdomen X-ray AP upright portable|Abdomen X-ray AP upright portable
C2826012|T102|strict|36960-3|LNC|Chest X-ray AP upright portable|Chest X-ray AP upright portable
C2826012|T102|strict|24807-0|LNC|Knee X-ray AP single view standing|Knee X-ray AP single view standing
C2826012|T102|strict|26358-2|LNC|Knee - bilateral X-ray AP single view standing|Knee - bilateral X-ray AP single view standing
C2826012|T102|strict|26359-0|LNC|Knee - left X-ray AP single view standing|Knee - left X-ray AP single view standing
C2826012|T102|strict|26360-8|LNC|Knee - right X-ray AP single view standing|Knee - right X-ray AP single view standing
C2826012|T102|strict|44177-4|LNC|Lower extremity - bilateral X-ray AP single view standing|Lower extremity - bilateral X-ray AP single view standing
C2826012|T102|strict|38849-6|LNC|Lower extremity - left X-ray AP single view standing|Lower extremity - left X-ray AP single view standing
C2826012|T102|strict|37733-3|LNC|Lower extremity - right X-ray AP single view standing|Lower extremity - right X-ray AP single view standing
C2826012|T102|strict|42420-0|LNC|Pelvis X-ray AP single view standing|Pelvis X-ray AP single view standing
C2826012|T102|strict|42378-0|LNC|Spine Lumbar X-ray AP single view W left bending|Spine Lumbar X-ray AP single view W left bending
C2826012|T102|strict|39410-6|LNC|Spine Thoracic X-ray AP single view W left bending|Spine Thoracic X-ray AP single view W left bending
C2826012|T102|strict|42379-8|LNC|Spine Lumbar X-ray AP single view W right bending|Spine Lumbar X-ray AP single view W right bending
C2826012|T102|strict|39411-4|LNC|Spine Thoracic X-ray AP single view W right bending|Spine Thoracic X-ray AP single view W right bending
C2826012|T102|strict|24723-9|LNC|Hand X-ray arthritis|Hand X-ray arthritis
C2826012|T102|strict|26355-8|LNC|Hand - bilateral X-ray arthritis|Hand - bilateral X-ray arthritis
C2826012|T102|strict|26356-6|LNC|Hand - left X-ray arthritis|Hand - left X-ray arthritis
C2826012|T102|strict|26357-4|LNC|Hand - right X-ray arthritis|Hand - right X-ray arthritis
C2826012|T102|strict|42395-4|LNC|Foot sesamoid bones - bilateral X-ray axial|Foot sesamoid bones - bilateral X-ray axial
C2826012|T102|strict|42396-2|LNC|Foot sesamoid bones - left X-ray axial|Foot sesamoid bones - left X-ray axial
C2826012|T102|strict|36962-9|LNC|Breast Mammogram axillary|Breast Mammogram axillary
C2826012|T102|strict|37849-7|LNC|Shoulder X-ray axillary|Shoulder X-ray axillary
C2826012|T102|strict|36963-7|LNC|Shoulder - bilateral X-ray axillary|Shoulder - bilateral X-ray axillary
C2826012|T102|strict|36964-5|LNC|Shoulder - left X-ray axillary|Shoulder - left X-ray axillary
C2826012|T102|strict|37800-0|LNC|Shoulder - right X-ray axillary|Shoulder - right X-ray axillary
C2826012|T102|strict|36965-2|LNC|Hand X-ray Ball Catcher|Hand X-ray Ball Catcher
C2826012|T102|strict|37471-0|LNC|Hand - bilateral X-ray Bora|Hand - bilateral X-ray Bora
C2826012|T102|strict|37472-8|LNC|Hand - left X-ray Bora|Hand - left X-ray Bora
C2826012|T102|strict|38804-1|LNC|Hand - right X-ray Bora|Hand - right X-ray Bora
C2826012|T102|strict|36966-0|LNC|Hand - bilateral X-ray Brewerton|Hand - bilateral X-ray Brewerton
C2826012|T102|strict|36967-8|LNC|Hand - left X-ray Brewerton|Hand - left X-ray Brewerton
C2826012|T102|strict|38775-3|LNC|Hand - right X-ray Brewerton|Hand - right X-ray Brewerton
C2826012|T102|strict|37928-9|LNC|Wrist X-ray Brewerton|Wrist X-ray Brewerton
C2826012|T102|strict|37857-0|LNC|Sinuses X-ray Caldwell|Sinuses X-ray Caldwell
C2826012|T102|strict|69132-9|LNC|Hip X-ray Danelius Miller|Hip X-ray Danelius Miller
C2826012|T102|strict|69141-0|LNC|Hip - left X-ray Danelius Miller|Hip - left X-ray Danelius Miller
C2826012|T102|strict|39514-5|LNC|Hip - right X-ray Danelius Miller|Hip - right X-ray Danelius Miller
C2826012|T102|strict|37625-1|LNC|Pelvis X-ray Ferguson|Pelvis X-ray Ferguson
C2826012|T102|strict|37650-9|LNC|Sacroiliac Joint X-ray Ferguson|Sacroiliac Joint X-ray Ferguson
C2826012|T102|strict|65799-9|LNC|Kidney - bilateral Fluoroscopy View for cyst examination|Kidney - bilateral Fluoroscopy View for cyst examination
C2826012|T102|strict|65800-5|LNC|Kidney - left Fluoroscopy View for cyst examination|Kidney - left Fluoroscopy View for cyst examination
C2826012|T102|strict|65801-3|LNC|Kidney - right Fluoroscopy View for cyst examination|Kidney - right Fluoroscopy View for cyst examination
C2826012|T102|strict|37297-9|LNC|Abdomen and Fetus X-ray View for fetal age|Abdomen and Fetus X-ray View for fetal age
C2826012|T102|strict|39149-0|LNC|Gastrointestinal system and Respiratory system X-ray for foreign body|Gastrointestinal system and Respiratory system X-ray for foreign body
C2826012|T102|strict|36973-6|LNC|Hip X-ray Friedman|Hip X-ray Friedman
C2826012|T102|strict|37843-0|LNC|Shoulder X-ray Garth|Shoulder X-ray Garth
C2826012|T102|strict|36974-4|LNC|Shoulder - left X-ray Garth|Shoulder - left X-ray Garth
C2826012|T102|strict|37801-8|LNC|Shoulder - right X-ray Garth|Shoulder - right X-ray Garth
C2826012|T102|strict|37844-8|LNC|Shoulder X-ray Grashey|Shoulder X-ray Grashey
C2826012|T102|strict|37035-3|LNC|Shoulder - bilateral X-ray Grashey|Shoulder - bilateral X-ray Grashey
C2826012|T102|strict|37473-6|LNC|Shoulder - left X-ray Grashey|Shoulder - left X-ray Grashey
C2826012|T102|strict|38805-8|LNC|Shoulder - right X-ray Grashey|Shoulder - right X-ray Grashey
C2826012|T102|strict|36975-1|LNC|Calcaneus - bilateral X-ray Harris|Calcaneus - bilateral X-ray Harris
C2826012|T102|strict|36977-7|LNC|Calcaneus - left X-ray Harris|Calcaneus - left X-ray Harris
C2826012|T102|strict|38776-1|LNC|Calcaneus - right X-ray Harris|Calcaneus - right X-ray Harris
C2826012|T102|strict|36976-9|LNC|Foot X-ray Harris|Foot X-ray Harris
C2826012|T102|strict|36978-5|LNC|Knee X-ray Holmblad|Knee X-ray Holmblad
C2826012|T102|strict|37628-5|LNC|Pelvis X-ray inlet|Pelvis X-ray inlet
C2826012|T102|strict|36979-3|LNC|Elbow X-ray Jones|Elbow X-ray Jones
C2826012|T102|strict|36980-1|LNC|Elbow - left X-ray Jones|Elbow - left X-ray Jones
C2826012|T102|strict|38777-9|LNC|Elbow - right X-ray Jones|Elbow - right X-ray Jones
C2826012|T102|strict|36981-9|LNC|Hip X-ray Judet|Hip X-ray Judet
C2826012|T102|strict|36982-7|LNC|Hip - bilateral X-ray Judet|Hip - bilateral X-ray Judet
C2826012|T102|strict|36983-5|LNC|Hip - left X-ray Judet|Hip - left X-ray Judet
C2826012|T102|strict|37732-5|LNC|Hip - right X-ray Judet|Hip - right X-ray Judet
C2826012|T102|strict|36620-3|LNC|Chest X-ray left anterior oblique|Chest X-ray left anterior oblique
C2826012|T102|strict|36591-6|LNC|Abdomen X-ray lateral|Abdomen X-ray lateral
C2826012|T102|strict|36592-4|LNC|Ankle X-ray lateral|Ankle X-ray lateral
C2826012|T102|strict|39051-8|LNC|Chest X-ray lateral|Chest X-ray lateral
C2826012|T102|strict|36593-2|LNC|Femur X-ray lateral|Femur X-ray lateral
C2826012|T102|strict|36594-0|LNC|Finger fifth X-ray lateral|Finger fifth X-ray lateral
C2826012|T102|strict|36595-7|LNC|Finger fourth X-ray lateral|Finger fourth X-ray lateral
C2826012|T102|strict|36596-5|LNC|Finger second X-ray lateral|Finger second X-ray lateral
C2826012|T102|strict|36597-3|LNC|Finger third X-ray lateral|Finger third X-ray lateral
C2826012|T102|strict|36598-1|LNC|Foot - left X-ray lateral|Foot - left X-ray lateral
C2826012|T102|strict|37703-6|LNC|Foot - right X-ray lateral|Foot - right X-ray lateral
C2826012|T102|strict|36599-9|LNC|Hand X-ray lateral|Hand X-ray lateral
C2826012|T102|strict|36600-5|LNC|Hand - bilateral X-ray lateral|Hand - bilateral X-ray lateral
C2826012|T102|strict|36601-3|LNC|Hand - left X-ray lateral|Hand - left X-ray lateral
C2826012|T102|strict|37712-7|LNC|Hand - right X-ray lateral|Hand - right X-ray lateral
C2826012|T102|strict|36602-1|LNC|Hip X-ray lateral|Hip X-ray lateral
C2826012|T102|strict|36603-9|LNC|Hip - left X-ray lateral|Hip - left X-ray lateral
C2826012|T102|strict|37730-9|LNC|Hip - right X-ray lateral|Hip - right X-ray lateral
C2826012|T102|strict|36604-7|LNC|Knee X-ray lateral|Knee X-ray lateral
C2826012|T102|strict|36605-4|LNC|Knee - bilateral X-ray lateral|Knee - bilateral X-ray lateral
C2826012|T102|strict|36606-2|LNC|Knee - left X-ray lateral|Knee - left X-ray lateral
C2826012|T102|strict|37751-5|LNC|Knee - right X-ray lateral|Knee - right X-ray lateral
C2826012|T102|strict|24843-5|LNC|Neck X-ray lateral|Neck X-ray lateral
C2826012|T102|strict|37629-3|LNC|Pelvis X-ray lateral|Pelvis X-ray lateral
C2826012|T102|strict|39053-4|LNC|Ribs X-ray lateral|Ribs X-ray lateral
C2826012|T102|strict|38857-9|LNC|Ribs - left X-ray lateral|Ribs - left X-ray lateral
C2826012|T102|strict|37784-6|LNC|Ribs - right X-ray lateral|Ribs - right X-ray lateral
C2826012|T102|strict|37858-8|LNC|Sinuses X-ray lateral|Sinuses X-ray lateral
C2826012|T102|strict|24920-1|LNC|Skull X-ray lateral|Skull X-ray lateral
C2826012|T102|strict|39052-6|LNC|Spine X-ray lateral|Spine X-ray lateral
C2826012|T102|strict|24943-3|LNC|Spine Cervical X-ray lateral|Spine Cervical X-ray lateral
C2826012|T102|strict|24969-8|LNC|Spine Lumbar X-ray lateral|Spine Lumbar X-ray lateral
C2826012|T102|strict|30756-1|LNC|Spine Thoracic X-ray lateral|Spine Thoracic X-ray lateral
C2826012|T102|strict|37891-9|LNC|Thumb X-ray lateral|Thumb X-ray lateral
C2826012|T102|strict|37893-5|LNC|Tibia and Fibula X-ray lateral|Tibia and Fibula X-ray lateral
C2826012|T102|strict|37930-5|LNC|Wrist X-ray lateral|Wrist X-ray lateral
C2826012|T102|strict|36984-3|LNC|Abdomen X-ray lateral crosstable|Abdomen X-ray lateral crosstable
C2826012|T102|strict|36985-0|LNC|Hip X-ray lateral crosstable|Hip X-ray lateral crosstable
C2826012|T102|strict|36986-8|LNC|Hip - bilateral X-ray lateral crosstable|Hip - bilateral X-ray lateral crosstable
C2826012|T102|strict|36987-6|LNC|Hip - left X-ray lateral crosstable|Hip - left X-ray lateral crosstable
C2826012|T102|strict|37727-5|LNC|Hip - right X-ray lateral crosstable|Hip - right X-ray lateral crosstable
C2826012|T102|strict|36988-4|LNC|Knee X-ray lateral crosstable|Knee X-ray lateral crosstable
C2826012|T102|strict|37872-9|LNC|Skull X-ray lateral crosstable|Skull X-ray lateral crosstable
C2826012|T102|strict|37878-6|LNC|Spine X-ray lateral crosstable|Spine X-ray lateral crosstable
C2826012|T102|strict|36989-2|LNC|Spine Cervical X-ray lateral crosstable|Spine Cervical X-ray lateral crosstable
C2826012|T102|strict|36990-0|LNC|Spine Lumbar X-ray lateral crosstable|Spine Lumbar X-ray lateral crosstable
C2826012|T102|strict|37903-2|LNC|Spine Thoracic X-ray lateral crosstable|Spine Thoracic X-ray lateral crosstable
C2826012|T102|strict|36991-8|LNC|Spine Cervical X-ray lateral crosstable portable|Spine Cervical X-ray lateral crosstable portable
C2826012|T102|strict|36992-6|LNC|Spine Lumbar X-ray lateral crosstable portable|Spine Lumbar X-ray lateral crosstable portable
C2826012|T102|strict|30786-8|LNC|Hip X-ray lateral frog|Hip X-ray lateral frog
C2826012|T102|strict|36993-4|LNC|Hip - bilateral X-ray lateral frog|Hip - bilateral X-ray lateral frog
C2826012|T102|strict|36994-2|LNC|Hip - left X-ray lateral frog|Hip - left X-ray lateral frog
C2826012|T102|strict|37729-1|LNC|Hip - right X-ray lateral frog|Hip - right X-ray lateral frog
C2826012|T102|strict|37626-9|LNC|Pelvis X-ray lateral frog|Pelvis X-ray lateral frog
C2826012|T102|strict|36999-1|LNC|Knee - bilateral X-ray lateral hyperextension|Knee - bilateral X-ray lateral hyperextension
C2826012|T102|strict|37000-7|LNC|Knee - left X-ray lateral hyperextension|Knee - left X-ray lateral hyperextension
C2826012|T102|strict|37750-7|LNC|Knee - right X-ray lateral hyperextension|Knee - right X-ray lateral hyperextension
C2826012|T102|strict|37909-9|LNC|Spine Thoracic X-ray lateral hyperextension|Spine Thoracic X-ray lateral hyperextension
C2826012|T102|strict|41774-1|LNC|Neck X-ray lateral portable|Neck X-ray lateral portable
C2826012|T102|strict|30757-9|LNC|Spine Thoracic X-ray lateral portable|Spine Thoracic X-ray lateral portable
C2826012|T102|strict|37515-4|LNC|Spine Lumbosacral Junction X-ray lateral spot|Spine Lumbosacral Junction X-ray lateral spot
C2826012|T102|strict|37516-2|LNC|Spine Lumbosacral Junction X-ray lateral spot standing|Spine Lumbosacral Junction X-ray lateral spot standing
C2826012|T102|strict|38066-7|LNC|Hip - left X-ray lateral during surgery|Hip - left X-ray lateral during surgery
C2826012|T102|strict|38819-9|LNC|Hip - right X-ray lateral during surgery|Hip - right X-ray lateral during surgery
C2826012|T102|strict|37001-5|LNC|Foot X-ray lateral standing|Foot X-ray lateral standing
C2826012|T102|strict|37002-3|LNC|Knee - left X-ray lateral standing|Knee - left X-ray lateral standing
C2826012|T102|strict|37754-9|LNC|Knee - right X-ray lateral standing|Knee - right X-ray lateral standing
C2826012|T102|strict|42442-4|LNC|Spine X-ray lateral standing|Spine X-ray lateral standing
C2826012|T102|strict|37003-1|LNC|Spine Lumbar X-ray lateral standing|Spine Lumbar X-ray lateral standing
C2826012|T102|strict|37910-7|LNC|Spine Thoracic X-ray lateral standing|Spine Thoracic X-ray lateral standing
C2826012|T102|strict|36997-5|LNC|Spine Cervical X-ray lateral W extension|Spine Cervical X-ray lateral W extension
C2826012|T102|strict|36971-0|LNC|Wrist - left X-ray lateral W extension|Wrist - left X-ray lateral W extension
C2826012|T102|strict|37833-1|LNC|Wrist - right X-ray lateral W extension|Wrist - right X-ray lateral W extension
C2826012|T102|strict|36998-3|LNC|Spine Cervical X-ray lateral W flexion|Spine Cervical X-ray lateral W flexion
C2826012|T102|strict|36972-8|LNC|Wrist - left X-ray lateral W flexion|Wrist - left X-ray lateral W flexion
C2826012|T102|strict|37834-9|LNC|Wrist - right X-ray lateral W flexion|Wrist - right X-ray lateral W flexion
C2826012|T102|strict|37004-9|LNC|Knee X-ray Laurin|Knee X-ray Laurin
C2826012|T102|strict|36995-9|LNC|Abdomen X-ray left lateral|Abdomen X-ray left lateral
C2826012|T102|strict|30737-1|LNC|Chest X-ray left lateral|Chest X-ray left lateral
C2826012|T102|strict|30738-9|LNC|Chest X-ray left lateral portable|Chest X-ray left lateral portable
C2826012|T102|strict|24639-7|LNC|Chest X-ray left lateral upright|Chest X-ray left lateral upright
C2826012|T102|strict|24638-9|LNC|Chest X-ray left lateral upright portable|Chest X-ray left lateral upright portable
C2826012|T102|strict|37008-0|LNC|Chest X-ray left oblique|Chest X-ray left oblique
C2826012|T102|strict|37009-8|LNC|Spine Lumbar X-ray left oblique|Spine Lumbar X-ray left oblique
C2826012|T102|strict|24641-3|LNC|Chest X-ray left oblique portable|Chest X-ray left oblique portable
C2826012|T102|strict|24640-5|LNC|Chest X-ray lordotic|Chest X-ray lordotic
C2826012|T102|strict|38069-1|LNC|Abdomen X-ray left posterior oblique|Abdomen X-ray left posterior oblique
C2826012|T102|strict|37005-6|LNC|Breast - left Mammogram magnification|Breast - left Mammogram magnification
C2826012|T102|strict|37773-9|LNC|Breast - right Mammogram magnification|Breast - right Mammogram magnification
C2826012|T102|strict|42441-6|LNC|Neck X-ray magnification|Neck X-ray magnification
C2826012|T102|strict|24801-3|LNC|Knee X-ray Merchants|Knee X-ray Merchants
C2826012|T102|strict|26283-2|LNC|Knee - bilateral X-ray Merchants|Knee - bilateral X-ray Merchants
C2826012|T102|strict|26284-0|LNC|Knee - left X-ray Merchants|Knee - left X-ray Merchants
C2826012|T102|strict|26285-7|LNC|Knee - right X-ray Merchants|Knee - right X-ray Merchants
C2826012|T102|strict|37006-4|LNC|Breast - bilateral Mammogram MLO|Breast - bilateral Mammogram MLO
C2826012|T102|strict|37007-2|LNC|Ankle X-ray Mortise|Ankle X-ray Mortise
C2826012|T102|strict|37475-1|LNC|Ankle - left X-ray Mortise W manual stress|Ankle - left X-ray Mortise W manual stress
C2826012|T102|strict|37671-5|LNC|Ankle - right X-ray Mortise W manual stress|Ankle - right X-ray Mortise W manual stress
C2826012|T102|strict|38067-5|LNC|Breast - bilateral Mammogram nipple profile|Breast - bilateral Mammogram nipple profile
C2826012|T102|strict|36607-0|LNC|Abdomen X-ray oblique single view|Abdomen X-ray oblique single view
C2826012|T102|strict|36609-6|LNC|Femur X-ray oblique single view|Femur X-ray oblique single view
C2826012|T102|strict|36610-4|LNC|Finger fifth X-ray oblique single view|Finger fifth X-ray oblique single view
C2826012|T102|strict|36611-2|LNC|Finger fourth X-ray oblique single view|Finger fourth X-ray oblique single view
C2826012|T102|strict|36612-0|LNC|Finger second X-ray oblique single view|Finger second X-ray oblique single view
C2826012|T102|strict|36613-8|LNC|Finger third X-ray oblique single view|Finger third X-ray oblique single view
C2826012|T102|strict|36614-6|LNC|Foot X-ray oblique single view|Foot X-ray oblique single view
C2826012|T102|strict|36615-3|LNC|Foot - left X-ray oblique single view|Foot - left X-ray oblique single view
C2826012|T102|strict|37704-4|LNC|Foot - right X-ray oblique single view|Foot - right X-ray oblique single view
C2826012|T102|strict|36616-1|LNC|Hand X-ray oblique single view|Hand X-ray oblique single view
C2826012|T102|strict|36617-9|LNC|Hip X-ray oblique single view|Hip X-ray oblique single view
C2826012|T102|strict|36618-7|LNC|Hip - bilateral X-ray oblique single view|Hip - bilateral X-ray oblique single view
C2826012|T102|strict|42689-0|LNC|Spine X-ray oblique single view|Spine X-ray oblique single view
C2826012|T102|strict|30778-5|LNC|Spine Lumbar X-ray oblique single view|Spine Lumbar X-ray oblique single view
C2826012|T102|strict|30758-7|LNC|Spine Thoracic X-ray oblique single view|Spine Thoracic X-ray oblique single view
C2826012|T102|strict|37892-7|LNC|Thumb X-ray oblique single view|Thumb X-ray oblique single view
C2826012|T102|strict|44178-2|LNC|Spine Lumbar X-ray oblique view and (views W right bending and W left bending)|Spine Lumbar X-ray oblique view and (views W right bending and W left bending)
C2826012|T102|strict|37545-1|LNC|Hip - left X-ray oblique crosstable|Hip - left X-ray oblique crosstable
C2826012|T102|strict|37728-3|LNC|Hip - right X-ray oblique crosstable|Hip - right X-ray oblique crosstable
C2826012|T102|strict|30759-5|LNC|Spine Thoracic X-ray oblique portable|Spine Thoracic X-ray oblique portable
C2826012|T102|strict|37631-9|LNC|Pelvis X-ray outlet|Pelvis X-ray outlet
C2826012|T102|strict|37845-5|LNC|Shoulder X-ray outlet|Shoulder X-ray outlet
C2826012|T102|strict|37012-2|LNC|Shoulder - bilateral X-ray outlet|Shoulder - bilateral X-ray outlet
C2826012|T102|strict|37013-0|LNC|Shoulder - left X-ray outlet|Shoulder - left X-ray outlet
C2826012|T102|strict|37802-6|LNC|Shoulder - right X-ray outlet|Shoulder - right X-ray outlet
C2826012|T102|strict|36621-1|LNC|Hand X-ray PA|Hand X-ray PA
C2826012|T102|strict|36622-9|LNC|Hand - bilateral X-ray PA|Hand - bilateral X-ray PA
C2826012|T102|strict|36623-7|LNC|Hand - left X-ray PA|Hand - left X-ray PA
C2826012|T102|strict|37714-3|LNC|Hand - right X-ray PA|Hand - right X-ray PA
C2826012|T102|strict|69270-7|LNC|Skull X-ray PA|Skull X-ray PA
C2826012|T102|strict|37931-3|LNC|Wrist X-ray PA|Wrist X-ray PA
C2826012|T102|strict|36624-5|LNC|Wrist - bilateral X-ray PA|Wrist - bilateral X-ray PA
C2826012|T102|strict|37015-5|LNC|Abdomen X-ray PA prone|Abdomen X-ray PA prone
C2826012|T102|strict|24648-8|LNC|Chest X-ray PA upright|Chest X-ray PA upright
C2826012|T102|strict|37014-8|LNC|Knee - left X-ray PA standing|Knee - left X-ray PA standing
C2826012|T102|strict|37755-6|LNC|Knee - right X-ray PA standing|Knee - right X-ray PA standing
C2826012|T102|strict|37477-7|LNC|Knee X-ray PA standing and W 45 degree flexion|Knee X-ray PA standing and W 45 degree flexion
C2826012|T102|strict|37476-9|LNC|Knee X-ray PA W 45 degree flexion|Knee X-ray PA W 45 degree flexion
C2826012|T102|strict|39324-9|LNC|Wrist - left X-ray PA W clenched fist|Wrist - left X-ray PA W clenched fist
C2826012|T102|strict|69263-2|LNC|Wrist - right X-ray PA W clenched fist|Wrist - right X-ray PA W clenched fist
C2826012|T102|strict|24828-6|LNC|Mandible X-ray panorex|Mandible X-ray panorex
C2826012|T102|strict|24871-6|LNC|Pelvis X-ray pelvimetry|Pelvis X-ray pelvimetry
C2826012|T102|strict|37998-2|LNC|Elbow X-ray radial head capitellar|Elbow X-ray radial head capitellar
C2826012|T102|strict|37999-0|LNC|Elbow - bilateral X-ray radial head capitellar|Elbow - bilateral X-ray radial head capitellar
C2826012|T102|strict|38000-6|LNC|Elbow - left X-ray radial head capitellar|Elbow - left X-ray radial head capitellar
C2826012|T102|strict|38006-3|LNC|Elbow - right X-ray radial head capitellar|Elbow - right X-ray radial head capitellar
C2826012|T102|strict|38068-3|LNC|Chest X-ray right anterior oblique|Chest X-ray right anterior oblique
C2826012|T102|strict|36996-7|LNC|Abdomen X-ray right lateral|Abdomen X-ray right lateral
C2826012|T102|strict|37010-6|LNC|Chest X-ray right oblique|Chest X-ray right oblique
C2826012|T102|strict|37011-4|LNC|Spine Lumbar X-ray right oblique|Spine Lumbar X-ray right oblique
C2826012|T102|strict|37018-9|LNC|Knee X-ray Rosenberg standing|Knee X-ray Rosenberg standing
C2826012|T102|strict|37020-5|LNC|Knee - bilateral X-ray Rosenberg standing|Knee - bilateral X-ray Rosenberg standing
C2826012|T102|strict|37019-7|LNC|Knee - left X-ray Rosenberg standing|Knee - left X-ray Rosenberg standing
C2826012|T102|strict|37752-3|LNC|Knee - right X-ray Rosenberg standing|Knee - right X-ray Rosenberg standing
C2826012|T102|strict|39323-1|LNC|Abdomen X-ray right posterior oblique|Abdomen X-ray right posterior oblique
C2826012|T102|strict|49511-9|LNC|Femoral artery Fluoroscopic angiogram runoff W and WO contrast IA|Femoral artery Fluoroscopic angiogram runoff W and WO contrast IA
C2826012|T102|strict|24699-1|LNC|Femoral artery Fluoroscopic angiogram runoff W contrast IA|Femoral artery Fluoroscopic angiogram runoff W contrast IA
C2826012|T102|strict|26178-4|LNC|Femoral artery - bilateral Fluoroscopic angiogram runoff W contrast IA|Femoral artery - bilateral Fluoroscopic angiogram runoff W contrast IA
C2826012|T102|strict|26179-2|LNC|Femoral artery - left Fluoroscopic angiogram runoff W contrast IA|Femoral artery - left Fluoroscopic angiogram runoff W contrast IA
C2826012|T102|strict|26180-0|LNC|Femoral artery - right Fluoroscopic angiogram runoff W contrast IA|Femoral artery - right Fluoroscopic angiogram runoff W contrast IA
C2826012|T102|strict|42812-8|LNC|Wrist X-ray scaphoid single view|Wrist X-ray scaphoid single view
C2826012|T102|strict|42813-6|LNC|Wrist - bilateral X-ray scaphoid single view|Wrist - bilateral X-ray scaphoid single view
C2826012|T102|strict|42814-4|LNC|Wrist - left X-ray scaphoid single view|Wrist - left X-ray scaphoid single view
C2826012|T102|strict|42811-0|LNC|Wrist - right X-ray scaphoid single view|Wrist - right X-ray scaphoid single view
C2826012|T102|strict|44206-1|LNC|Spine Thoracic and Lumbar X-ray scoliosis single view|Spine Thoracic and Lumbar X-ray scoliosis single view
C2826012|T102|strict|30714-0|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP|Spine Thoracic and Lumbar X-ray scoliosis AP
C2826012|T102|strict|42426-7|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP sitting|Spine Thoracic and Lumbar X-ray scoliosis AP sitting
C2826012|T102|strict|37659-0|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP standing|Spine Thoracic and Lumbar X-ray scoliosis AP standing
C2826012|T102|strict|42428-3|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP standing and in brace|Spine Thoracic and Lumbar X-ray scoliosis AP standing and in brace
C2826012|T102|strict|42429-1|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP standing and W right bending|Spine Thoracic and Lumbar X-ray scoliosis AP standing and W right bending
C2826012|T102|strict|42427-5|LNC|Spine Thoracic and Lumbar X-ray scoliosis lateral sitting|Spine Thoracic and Lumbar X-ray scoliosis lateral sitting
C2826012|T102|strict|37660-8|LNC|Spine Thoracic and Lumbar X-ray scoliosis lateral standing|Spine Thoracic and Lumbar X-ray scoliosis lateral standing
C2826012|T102|strict|37846-3|LNC|Sternoclavicular Joint X-ray Serendipity|Sternoclavicular Joint X-ray Serendipity
C2826012|T102|strict|37298-7|LNC|Sternoclavicular joint - bilateral X-ray Serendipity|Sternoclavicular joint - bilateral X-ray Serendipity
C2826012|T102|strict|37299-5|LNC|Sternoclavicular joint - left X-ray Serendipity|Sternoclavicular joint - left X-ray Serendipity
C2826012|T102|strict|37808-3|LNC|Sternoclavicular joint - right X-ray Serendipity|Sternoclavicular joint - right X-ray Serendipity
C2826012|T102|strict|43671-7|LNC|Thyroid Scan spot|Thyroid Scan spot
C2826012|T102|strict|42471-3|LNC|Pelvis X-ray stereo|Pelvis X-ray stereo
C2826012|T102|strict|42474-7|LNC|Skull X-ray stereo|Skull X-ray stereo
C2826012|T102|strict|39516-0|LNC|Shoulder X-ray Stryker Notch|Shoulder X-ray Stryker Notch
C2826012|T102|strict|37024-7|LNC|Shoulder - bilateral X-ray Stryker Notch|Shoulder - bilateral X-ray Stryker Notch
C2826012|T102|strict|37025-4|LNC|Shoulder - left X-ray Stryker Notch|Shoulder - left X-ray Stryker Notch
C2826012|T102|strict|37791-1|LNC|Shoulder - right X-ray Stryker Notch|Shoulder - right X-ray Stryker Notch
C2826012|T102|strict|39517-8|LNC|Shoulder X-ray Stryker Notch and West Point|Shoulder X-ray Stryker Notch and West Point
C2826012|T102|strict|37861-2|LNC|Sinuses X-ray submentovertex|Sinuses X-ray submentovertex
C2826012|T102|strict|37026-2|LNC|Skull X-ray submentovertex|Skull X-ray submentovertex
C2826012|T102|strict|43780-6|LNC|Knee X-ray Sunrise|Knee X-ray Sunrise
C2826012|T102|strict|37027-0|LNC|Knee - bilateral X-ray Sunrise|Knee - bilateral X-ray Sunrise
C2826012|T102|strict|43779-8|LNC|Knee - left X-ray Sunrise|Knee - left X-ray Sunrise
C2826012|T102|strict|69256-6|LNC|Knee - right X-ray Sunrise|Knee - right X-ray Sunrise
C2826012|T102|strict|69239-2|LNC|Patella X-ray Sunrise|Patella X-ray Sunrise
C2826012|T102|strict|69069-3|LNC|Patella - bilateral X-ray Sunrise|Patella - bilateral X-ray Sunrise
C2826012|T102|strict|69064-4|LNC|Knee - bilateral X-ray Sunrise and (views standing)|Knee - bilateral X-ray Sunrise and (views standing)
C2826012|T102|strict|69149-3|LNC|Knee - left X-ray Sunrise and (views standing)|Knee - left X-ray Sunrise and (views standing)
C2826012|T102|strict|42432-5|LNC|Knee - right X-ray Sunrise and (views standing)|Knee - right X-ray Sunrise and (views standing)
C2826012|T102|strict|24944-1|LNC|Spine Cervical X-ray Swimmers|Spine Cervical X-ray Swimmers
C2826012|T102|strict|37028-8|LNC|Breast Mammogram tangential|Breast Mammogram tangential
C2826012|T102|strict|37029-6|LNC|Breast - bilateral Mammogram tangential|Breast - bilateral Mammogram tangential
C2826012|T102|strict|37030-4|LNC|Breast - left Mammogram tangential|Breast - left Mammogram tangential
C2826012|T102|strict|37770-5|LNC|Breast - right Mammogram tangential|Breast - right Mammogram tangential
C2826012|T102|strict|37870-3|LNC|Skull X-ray Towne|Skull X-ray Towne
C2826012|T102|strict|24668-6|LNC|Colon Fluoroscopy transit Post solid contrast|Colon Fluoroscopy transit Post solid contrast
C2826012|T102|strict|37031-2|LNC|Humerus X-ray transthoracic|Humerus X-ray transthoracic
C2826012|T102|strict|37032-0|LNC|Humerus - bilateral X-ray transthoracic|Humerus - bilateral X-ray transthoracic
C2826012|T102|strict|37033-8|LNC|Humerus - left X-ray transthoracic|Humerus - left X-ray transthoracic
C2826012|T102|strict|38007-1|LNC|Humerus - right X-ray transthoracic|Humerus - right X-ray transthoracic
C2826012|T102|strict|37034-6|LNC|Shoulder - left X-ray transthoracic|Shoulder - left X-ray transthoracic
C2826012|T102|strict|38779-5|LNC|Shoulder - right X-ray transthoracic|Shoulder - right X-ray transthoracic
C2826012|T102|strict|37300-1|LNC|Spine Lumbosacral Junction X-ray true AP|Spine Lumbosacral Junction X-ray true AP
C2826012|T102|strict|37037-9|LNC|Breast Mammogram true lateral|Breast Mammogram true lateral
C2826012|T102|strict|37038-7|LNC|Breast - bilateral Mammogram true lateral|Breast - bilateral Mammogram true lateral
C2826012|T102|strict|38855-3|LNC|Breast - left Mammogram true lateral|Breast - left Mammogram true lateral
C2826012|T102|strict|37771-3|LNC|Breast - right Mammogram true lateral|Breast - right Mammogram true lateral
C2826012|T102|strict|37039-5|LNC|Hip X-ray true lateral|Hip X-ray true lateral
C2826012|T102|strict|37040-3|LNC|Hip - left X-ray true lateral|Hip - left X-ray true lateral
C2826012|T102|strict|38772-0|LNC|Hip - right X-ray true lateral|Hip - right X-ray true lateral
C2826012|T102|strict|30790-0|LNC|Knee X-ray tunnel|Knee X-ray tunnel
C2826012|T102|strict|37041-1|LNC|Knee - bilateral X-ray tunnel|Knee - bilateral X-ray tunnel
C2826012|T102|strict|37042-9|LNC|Knee - left X-ray tunnel|Knee - left X-ray tunnel
C2826012|T102|strict|37761-4|LNC|Knee - right X-ray tunnel|Knee - right X-ray tunnel
C2826012|T102|strict|38842-1|LNC|Wrist - left X-ray tunnel.carpal|Wrist - left X-ray tunnel.carpal
C2826012|T102|strict|37677-2|LNC|Wrist - right X-ray tunnel.carpal|Wrist - right X-ray tunnel.carpal
C2826012|T102|strict|37043-7|LNC|Knee - left X-ray tunnel standing|Knee - left X-ray tunnel standing
C2826012|T102|strict|37756-4|LNC|Knee - right X-ray tunnel standing|Knee - right X-ray tunnel standing
C2826012|T102|strict|37044-5|LNC|Wrist - left X-ray ulnar deviation|Wrist - left X-ray ulnar deviation
C2826012|T102|strict|37645-9|LNC|Wrist - right X-ray ulnar deviation|Wrist - right X-ray ulnar deviation
C2826012|T102|strict|37045-2|LNC|Wrist - bilateral X-ray ulnar variance|Wrist - bilateral X-ray ulnar variance
C2826012|T102|strict|37046-0|LNC|Abdomen X-ray upright|Abdomen X-ray upright
C2826012|T102|strict|37047-8|LNC|Shoulder - bilateral X-ray Velpeau axillary|Shoulder - bilateral X-ray Velpeau axillary
C2826012|T102|strict|37048-6|LNC|Shoulder - left X-ray Velpeau axillary|Shoulder - left X-ray Velpeau axillary
C2826012|T102|strict|38780-3|LNC|Shoulder - right X-ray Velpeau axillary|Shoulder - right X-ray Velpeau axillary
C2826012|T102|strict|37049-4|LNC|Hip X-ray Von rossen|Hip X-ray Von rossen
C2826012|T102|strict|37613-7|LNC|Orbit - bilateral X-ray Waters|Orbit - bilateral X-ray Waters
C2826012|T102|strict|37863-8|LNC|Sinuses X-ray Waters|Sinuses X-ray Waters
C2826012|T102|strict|24921-9|LNC|Skull X-ray Waters|Skull X-ray Waters
C2826012|T102|strict|42473-9|LNC|Sinuses X-ray Waters stereo|Sinuses X-ray Waters stereo
C2826012|T102|strict|38117-8|LNC|Sinuses X-ray Waters upright|Sinuses X-ray Waters upright
C2826012|T102|strict|30751-2|LNC|Shoulder X-ray West Point|Shoulder X-ray West Point
C2826012|T102|strict|37050-2|LNC|Shoulder - bilateral X-ray West Point|Shoulder - bilateral X-ray West Point
C2826012|T102|strict|37051-0|LNC|Shoulder - left X-ray West Point|Shoulder - left X-ray West Point
C2826012|T102|strict|37809-1|LNC|Shoulder - right X-ray West Point|Shoulder - right X-ray West Point
C2826012|T102|strict|42680-9|LNC|Breast Mammogram XCCL|Breast Mammogram XCCL
C2826012|T102|strict|37052-8|LNC|Breast - bilateral Mammogram XCCL|Breast - bilateral Mammogram XCCL
C2826012|T102|strict|37053-6|LNC|Breast - left Mammogram XCCL|Breast - left Mammogram XCCL
C2826012|T102|strict|37772-1|LNC|Breast - right Mammogram XCCL|Breast - right Mammogram XCCL
C2826012|T102|strict|37656-6|LNC|Scapula X-ray Y|Scapula X-ray Y
C2826012|T102|strict|37055-1|LNC|Scapula - bilateral X-ray Y|Scapula - bilateral X-ray Y
C2826012|T102|strict|37054-4|LNC|Scapula - left X-ray Y|Scapula - left X-ray Y
C2826012|T102|strict|37790-3|LNC|Scapula - right X-ray Y|Scapula - right X-ray Y
C2826012|T102|strict|37847-1|LNC|Shoulder X-ray Y|Shoulder X-ray Y
C2826012|T102|strict|38858-7|LNC|Shoulder - left X-ray Y|Shoulder - left X-ray Y
C2826012|T102|strict|37805-9|LNC|Shoulder - right X-ray Y|Shoulder - right X-ray Y
C2826012|T102|strict|37848-9|LNC|Acromioclavicular Joint X-ray Zanca|Acromioclavicular Joint X-ray Zanca
C2826012|T102|strict|37056-9|LNC|Acromioclavicular joint - bilateral X-ray Zanca|Acromioclavicular joint - bilateral X-ray Zanca
C2826012|T102|strict|37057-7|LNC|Acromioclavicular joint - left X-ray Zanca|Acromioclavicular joint - left X-ray Zanca
C2826012|T102|strict|37810-9|LNC|Acromioclavicular joint - right X-ray Zanca|Acromioclavicular joint - right X-ray Zanca
C2826012|T102|strict|41793-1|LNC|Abdomen X-ray during surgery|Abdomen X-ray during surgery
C2826012|T102|strict|41790-7|LNC|Chest X-ray during surgery|Chest X-ray during surgery
C2826012|T102|strict|24656-1|LNC|Chest Fluoroscopy during surgery|Chest Fluoroscopy during surgery
C2826012|T102|strict|39047-6|LNC|Hip Fluoroscopy during surgery|Hip Fluoroscopy during surgery
C2826012|T102|strict|38065-9|LNC|Hip - left X-ray during surgery|Hip - left X-ray during surgery
C2826012|T102|strict|38818-1|LNC|Hip - right X-ray during surgery|Hip - right X-ray during surgery
C2826012|T102|strict|42008-3|LNC|Humerus X-ray during surgery|Humerus X-ray during surgery
C2826012|T102|strict|24893-0|LNC|Rectum Fluoroscopy post contrast PR during defecation|Rectum Fluoroscopy post contrast PR during defecation
C2826012|T102|strict|37058-5|LNC|Calcaneus - bilateral X-ray standing|Calcaneus - bilateral X-ray standing
C2826012|T102|strict|37059-3|LNC|Hip - bilateral X-ray standing|Hip - bilateral X-ray standing
C2826012|T102|strict|37207-8|LNC|Hip - left X-ray standing|Hip - left X-ray standing
C2826012|T102|strict|37731-7|LNC|Hip - right X-ray standing|Hip - right X-ray standing
C2826012|T102|strict|44205-3|LNC|Lower extremity - bilateral X-ray standing|Lower extremity - bilateral X-ray standing
C2826012|T102|strict|38850-4|LNC|Lower extremity - left X-ray standing|Lower extremity - left X-ray standing
C2826012|T102|strict|37734-1|LNC|Lower extremity - right X-ray standing|Lower extremity - right X-ray standing
C2826012|T102|strict|37633-5|LNC|Pelvis X-ray standing|Pelvis X-ray standing
C2826012|T102|strict|39144-1|LNC|Gastrointestine upper Fluoroscopy W air contrast PO|Gastrointestine upper Fluoroscopy W air contrast PO
C2826012|T102|strict|41795-6|LNC|Upper Gastrointestine and Small bowel Fluoroscopy W air contrast PO|Upper Gastrointestine and Small bowel Fluoroscopy W air contrast PO
C2826012|T102|strict|69302-8|LNC|Wrist X-ray W clenched fist|Wrist X-ray W clenched fist
C2826012|T102|strict|36968-6|LNC|Wrist - bilateral X-ray W clenched fist|Wrist - bilateral X-ray W clenched fist
C2826012|T102|strict|30639-9|LNC|Vessel Fluoroscopic angiogram W contrast|Vessel Fluoroscopic angiogram W contrast
C2826012|T102|strict|42470-5|LNC|Gastrointestine upper and Gallbladder Fluoroscopy W contrast PO|Gastrointestine upper and Gallbladder Fluoroscopy W contrast PO
C2826012|T102|strict|30809-8|LNC|Upper Gastrointestine and Small bowel Fluoroscopy W contrast PO|Upper Gastrointestine and Small bowel Fluoroscopy W contrast PO
C2826012|T102|strict|42469-7|LNC|Gastrointestine upper and Small bowel and Gallbladder Fluoroscopy W contrast PO|Gastrointestine upper and Small bowel and Gallbladder Fluoroscopy W contrast PO
C2826012|T102|strict|38001-4|LNC|Chest X-ray W expiration|Chest X-ray W expiration
C2826012|T102|strict|38002-2|LNC|Chest X-ray W inspiration|Chest X-ray W inspiration
C2826012|T102|strict|37060-1|LNC|Fetal X-ray|Fetal X-ray
C2826012|T102|strict|37636-8|LNC|Abdomen X-ray|Abdomen X-ray
C2826012|T102|strict|46341-4|LNC|Abdomen Fluoroscopy|Abdomen Fluoroscopy
C2826012|T102|strict|24535-7|LNC|Acetabulum X-ray|Acetabulum X-ray
C2826012|T102|strict|26133-9|LNC|Acetabulum - bilateral X-ray|Acetabulum - bilateral X-ray
C2826012|T102|strict|26134-7|LNC|Acetabulum - left X-ray|Acetabulum - left X-ray
C2826012|T102|strict|26135-4|LNC|Acetabulum - right X-ray|Acetabulum - right X-ray
C2826012|T102|strict|24536-5|LNC|Acromioclavicular Joint X-ray|Acromioclavicular Joint X-ray
C2826012|T102|strict|26136-2|LNC|Acromioclavicular joint - bilateral X-ray|Acromioclavicular joint - bilateral X-ray
C2826012|T102|strict|26137-0|LNC|Acromioclavicular joint - left X-ray|Acromioclavicular joint - left X-ray
C2826012|T102|strict|26138-8|LNC|Acromioclavicular joint - right X-ray|Acromioclavicular joint - right X-ray
C2826012|T102|strict|24541-5|LNC|Ankle X-ray|Ankle X-ray
C2826012|T102|strict|26097-6|LNC|Ankle - bilateral X-ray|Ankle - bilateral X-ray
C2826012|T102|strict|26098-4|LNC|Ankle - left X-ray|Ankle - left X-ray
C2826012|T102|strict|51395-2|LNC|Ankle - left and Foot.left X-ray|Ankle - left and Foot.left X-ray
C2826012|T102|strict|26099-2|LNC|Ankle - right X-ray|Ankle - right X-ray
C2826012|T102|strict|51394-5|LNC|Ankle - right and Foot - right X-ray|Ankle - right and Foot - right X-ray
C2826012|T102|strict|36625-2|LNC|Breast Mammogram|Breast Mammogram
C2826012|T102|strict|46342-2|LNC|Breast FFD mammogram|Breast FFD mammogram
C2826012|T102|strict|38070-9|LNC|Breast implant Mammogram|Breast implant Mammogram
C2826012|T102|strict|38071-7|LNC|Breast implant - bilateral Mammogram|Breast implant - bilateral Mammogram
C2826012|T102|strict|38072-5|LNC|Breast implant - left Mammogram|Breast implant - left Mammogram
C2826012|T102|strict|38820-7|LNC|Breast implant - right Mammogram|Breast implant - right Mammogram
C2826012|T102|strict|46380-2|LNC|Breast Implant - unilateral Mammogram|Breast Implant - unilateral Mammogram
C2826012|T102|strict|24597-7|LNC|Breast specimen Mammogram|Breast specimen Mammogram
C2826012|T102|strict|38079-0|LNC|Breast specimen - bilateral Mammogram|Breast specimen - bilateral Mammogram
C2826012|T102|strict|38080-8|LNC|Breast specimen - left Mammogram|Breast specimen - left Mammogram
C2826012|T102|strict|38821-5|LNC|Breast specimen - right Mammogram|Breast specimen - right Mammogram
C2826012|T102|strict|36626-0|LNC|Breast - bilateral Mammogram|Breast - bilateral Mammogram
C2826012|T102|strict|36627-8|LNC|Breast - left Mammogram|Breast - left Mammogram
C2826012|T102|strict|37774-7|LNC|Breast - right Mammogram|Breast - right Mammogram
C2826012|T102|strict|46339-8|LNC|Breast - unilateral Mammogram|Breast - unilateral Mammogram
C2826012|T102|strict|24612-4|LNC|Calcaneus X-ray|Calcaneus X-ray
C2826012|T102|strict|26100-8|LNC|Calcaneus - bilateral X-ray|Calcaneus - bilateral X-ray
C2826012|T102|strict|26101-6|LNC|Calcaneus - left X-ray|Calcaneus - left X-ray
C2826012|T102|strict|26102-4|LNC|Calcaneus - right X-ray|Calcaneus - right X-ray
C2826012|T102|strict|30745-4|LNC|Chest X-ray|Chest X-ray
C2826012|T102|strict|30631-6|LNC|Chest Fluoroscopy|Chest Fluoroscopy
C2826012|T102|strict|42269-1|LNC|Chest and Abdomen X-ray|Chest and Abdomen X-ray
C2826012|T102|strict|24664-5|LNC|Clavicle X-ray|Clavicle X-ray
C2826012|T102|strict|26106-5|LNC|Clavicle - bilateral X-ray|Clavicle - bilateral X-ray
C2826012|T102|strict|26107-3|LNC|Clavicle - left X-ray|Clavicle - left X-ray
C2826012|T102|strict|26108-1|LNC|Clavicle - right X-ray|Clavicle - right X-ray
C2826012|T102|strict|30883-3|LNC|Coccyx X-ray|Coccyx X-ray
C2826012|T102|strict|24676-9|LNC|Elbow X-ray|Elbow X-ray
C2826012|T102|strict|26109-9|LNC|Elbow - bilateral X-ray|Elbow - bilateral X-ray
C2826012|T102|strict|26110-7|LNC|Elbow - left X-ray|Elbow - left X-ray
C2826012|T102|strict|26111-5|LNC|Elbow - right X-ray|Elbow - right X-ray
C2826012|T102|strict|46381-0|LNC|Elbow+Radius+Ulna X-ray|Elbow+Radius+Ulna X-ray
C2826012|T102|strict|37637-6|LNC|Extremity X-ray|Extremity X-ray
C2826012|T102|strict|24695-9|LNC|Facial bones X-ray|Facial bones X-ray
C2826012|T102|strict|37303-5|LNC|Facial bones and Zygomatic arch X-ray|Facial bones and Zygomatic arch X-ray
C2826012|T102|strict|24704-9|LNC|Femur X-ray|Femur X-ray
C2826012|T102|strict|26118-0|LNC|Femur - bilateral X-ray|Femur - bilateral X-ray
C2826012|T102|strict|26120-6|LNC|Femur - left X-ray|Femur - left X-ray
C2826012|T102|strict|26122-2|LNC|Femur - right X-ray|Femur - right X-ray
C2826012|T102|strict|24706-4|LNC|Finger X-ray|Finger X-ray
C2826012|T102|strict|26124-8|LNC|Finger - bilateral X-ray|Finger - bilateral X-ray
C2826012|T102|strict|30783-5|LNC|Finger fifth X-ray|Finger fifth X-ray
C2826012|T102|strict|37517-0|LNC|Finger fifth - bilateral X-ray|Finger fifth - bilateral X-ray
C2826012|T102|strict|37518-8|LNC|Finger fifth - left X-ray|Finger fifth - left X-ray
C2826012|T102|strict|38147-5|LNC|Finger fifth - right X-ray|Finger fifth - right X-ray
C2826012|T102|strict|30782-7|LNC|Finger fourth X-ray|Finger fourth X-ray
C2826012|T102|strict|37519-6|LNC|Finger fourth - bilateral X-ray|Finger fourth - bilateral X-ray
C2826012|T102|strict|37520-4|LNC|Finger fourth - left X-ray|Finger fourth - left X-ray
C2826012|T102|strict|38146-7|LNC|Finger fourth - right X-ray|Finger fourth - right X-ray
C2826012|T102|strict|26125-5|LNC|Finger - left X-ray|Finger - left X-ray
C2826012|T102|strict|26126-3|LNC|Finger - right X-ray|Finger - right X-ray
C2826012|T102|strict|30780-1|LNC|Finger second X-ray|Finger second X-ray
C2826012|T102|strict|37521-2|LNC|Finger second - bilateral X-ray|Finger second - bilateral X-ray
C2826012|T102|strict|37522-0|LNC|Finger second - left X-ray|Finger second - left X-ray
C2826012|T102|strict|38144-2|LNC|Finger second - right X-ray|Finger second - right X-ray
C2826012|T102|strict|30781-9|LNC|Finger third X-ray|Finger third X-ray
C2826012|T102|strict|37523-8|LNC|Finger third - bilateral X-ray|Finger third - bilateral X-ray
C2826012|T102|strict|37524-6|LNC|Finger third - left X-ray|Finger third - left X-ray
C2826012|T102|strict|38145-9|LNC|Finger third - right X-ray|Finger third - right X-ray
C2826012|T102|strict|24709-8|LNC|Foot X-ray|Foot X-ray
C2826012|T102|strict|26127-1|LNC|Foot - bilateral X-ray|Foot - bilateral X-ray
C2826012|T102|strict|26128-9|LNC|Foot - left X-ray|Foot - left X-ray
C2826012|T102|strict|26129-7|LNC|Foot - right X-ray|Foot - right X-ray
C2826012|T102|strict|42399-6|LNC|Foot sesamoid bones X-ray|Foot sesamoid bones X-ray
C2826012|T102|strict|42400-2|LNC|Foot sesamoid bones - bilateral X-ray|Foot sesamoid bones - bilateral X-ray
C2826012|T102|strict|43641-0|LNC|Foot sesamoid bones - left X-ray|Foot sesamoid bones - left X-ray
C2826012|T102|strict|42434-1|LNC|Foot sesamoid bones - right X-ray|Foot sesamoid bones - right X-ray
C2826012|T102|strict|37532-9|LNC|Great toe - bilateral X-ray|Great toe - bilateral X-ray
C2826012|T102|strict|37533-7|LNC|Great toe - left X-ray|Great toe - left X-ray
C2826012|T102|strict|38152-5|LNC|Great toe - right X-ray|Great toe - right X-ray
C2826012|T102|strict|28582-5|LNC|Hand X-ray|Hand X-ray
C2826012|T102|strict|36629-4|LNC|Hand - bilateral X-ray|Hand - bilateral X-ray
C2826012|T102|strict|36630-2|LNC|Hand - left X-ray|Hand - left X-ray
C2826012|T102|strict|37716-8|LNC|Hand - right X-ray|Hand - right X-ray
C2826012|T102|strict|24752-8|LNC|Heart Fluoroscopy video|Heart Fluoroscopy video
C2826012|T102|strict|24762-7|LNC|Hip X-ray|Hip X-ray
C2826012|T102|strict|26130-5|LNC|Hip - bilateral X-ray|Hip - bilateral X-ray
C2826012|T102|strict|26131-3|LNC|Hip - left X-ray|Hip - left X-ray
C2826012|T102|strict|26132-1|LNC|Hip - right X-ray|Hip - right X-ray
C2826012|T102|strict|28567-6|LNC|Humerus X-ray|Humerus X-ray
C2826012|T102|strict|37319-1|LNC|Humerus bicipital groove X-ray|Humerus bicipital groove X-ray
C2826012|T102|strict|37321-7|LNC|Humerus bicipital groove - bilateral X-ray|Humerus bicipital groove - bilateral X-ray
C2826012|T102|strict|37320-9|LNC|Humerus bicipital groove - left X-ray|Humerus bicipital groove - left X-ray
C2826012|T102|strict|38797-7|LNC|Humerus bicipital groove - right X-ray|Humerus bicipital groove - right X-ray
C2826012|T102|strict|37062-7|LNC|Humerus - bilateral X-ray|Humerus - bilateral X-ray
C2826012|T102|strict|36632-8|LNC|Humerus - left X-ray|Humerus - left X-ray
C2826012|T102|strict|37738-2|LNC|Humerus - right X-ray|Humerus - right X-ray
C2826012|T102|strict|36628-6|LNC|Internal auditory canal X-ray|Internal auditory canal X-ray
C2826012|T102|strict|28565-0|LNC|Knee X-ray|Knee X-ray
C2826012|T102|strict|36635-1|LNC|Knee - bilateral X-ray|Knee - bilateral X-ray
C2826012|T102|strict|36636-9|LNC|Knee - left X-ray|Knee - left X-ray
C2826012|T102|strict|37758-0|LNC|Knee - right X-ray|Knee - right X-ray
C2826012|T102|strict|48465-9|LNC|Larynx Fluoroscopy|Larynx Fluoroscopy
C2826012|T102|strict|24686-8|LNC|Lower extremity X-ray|Lower extremity X-ray
C2826012|T102|strict|26112-3|LNC|Lower extremity - bilateral X-ray|Lower extremity - bilateral X-ray
C2826012|T102|strict|26113-1|LNC|Lower extremity - left X-ray|Lower extremity - left X-ray
C2826012|T102|strict|26114-9|LNC|Lower extremity - right X-ray|Lower extremity - right X-ray
C2826012|T102|strict|24829-4|LNC|Mandible X-ray|Mandible X-ray
C2826012|T102|strict|48745-4|LNC|Mandible - left X-ray|Mandible - left X-ray
C2826012|T102|strict|43533-9|LNC|Mandible - right X-ray|Mandible - right X-ray
C2826012|T102|strict|24830-2|LNC|Mastoid X-ray|Mastoid X-ray
C2826012|T102|strict|26139-6|LNC|Mastoid - bilateral X-ray|Mastoid - bilateral X-ray
C2826012|T102|strict|26140-4|LNC|Mastoid - left X-ray|Mastoid - left X-ray
C2826012|T102|strict|26141-2|LNC|Mastoid - right X-ray|Mastoid - right X-ray
C2826012|T102|strict|36637-7|LNC|Maxilla X-ray|Maxilla X-ray
C2826012|T102|strict|24834-4|LNC|Nasal bones X-ray|Nasal bones X-ray
C2826012|T102|strict|37639-2|LNC|Neck X-ray|Neck X-ray
C2826012|T102|strict|37332-4|LNC|Olecranon - left X-ray|Olecranon - left X-ray
C2826012|T102|strict|38798-5|LNC|Olecranon - right X-ray|Olecranon - right X-ray
C2826012|T102|strict|24846-8|LNC|Optic foramen X-ray|Optic foramen X-ray
C2826012|T102|strict|26142-0|LNC|Optic foramen - bilateral X-ray|Optic foramen - bilateral X-ray
C2826012|T102|strict|26143-8|LNC|Optic foramen - left X-ray|Optic foramen - left X-ray
C2826012|T102|strict|26144-6|LNC|Optic foramen - right X-ray|Optic foramen - right X-ray
C2826012|T102|strict|36886-0|LNC|Orbit X-ray|Orbit X-ray
C2826012|T102|strict|24854-2|LNC|Orbit - bilateral X-ray|Orbit - bilateral X-ray
C2826012|T102|strict|36887-8|LNC|Orbit - left X-ray|Orbit - left X-ray
C2826012|T102|strict|38774-6|LNC|Orbit - right X-ray|Orbit - right X-ray
C2826012|T102|strict|43529-7|LNC|Orbit + Facial bones X-ray|Orbit + Facial bones X-ray
C2826012|T102|strict|24855-9|LNC|Oropharynx Fluoroscopy video|Oropharynx Fluoroscopy video
C2826012|T102|strict|30791-8|LNC|Patella X-ray|Patella X-ray
C2826012|T102|strict|36638-5|LNC|Patella - bilateral X-ray|Patella - bilateral X-ray
C2826012|T102|strict|36639-3|LNC|Patella - left X-ray|Patella - left X-ray
C2826012|T102|strict|37777-0|LNC|Patella - right X-ray|Patella - right X-ray
C2826012|T102|strict|28561-9|LNC|Pelvis X-ray|Pelvis X-ray
C2826012|T102|strict|30885-8|LNC|Pelvis symphysis pubis X-ray|Pelvis symphysis pubis X-ray
C2826012|T102|strict|30767-8|LNC|Pelvis and Hip X-ray|Pelvis and Hip X-ray
C2826012|T102|strict|30768-6|LNC|Pelvis and Hip - bilateral X-ray|Pelvis and Hip - bilateral X-ray
C2826012|T102|strict|36631-0|LNC|Pelvis and Hip - left X-ray|Pelvis and Hip - left X-ray
C2826012|T102|strict|38771-2|LNC|Pelvis and Hip - right X-ray|Pelvis and Hip - right X-ray
C2826012|T102|strict|47984-0|LNC|Pelvis and Spine Lumbar X-ray|Pelvis and Spine Lumbar X-ray
C2826012|T102|strict|24745-2|LNC|Petrous bone X-ray|Petrous bone X-ray
C2826012|T102|strict|26146-1|LNC|Radius - bilateral and Ulna - bilateral X-ray|Radius - bilateral and Ulna - bilateral X-ray
C2826012|T102|strict|26148-7|LNC|Radius - left and Ulna.left X-ray|Radius - left and Ulna.left X-ray
C2826012|T102|strict|26150-3|LNC|Radius - right and Ulna - right X-ray|Radius - right and Ulna - right X-ray
C2826012|T102|strict|24891-4|LNC|Radius and Ulna X-ray|Radius and Ulna X-ray
C2826012|T102|strict|24899-7|LNC|Ribs X-ray|Ribs X-ray
C2826012|T102|strict|37937-0|LNC|Ribs anterior X-ray|Ribs anterior X-ray
C2826012|T102|strict|38073-3|LNC|Ribs anterior - bilateral X-ray|Ribs anterior - bilateral X-ray
C2826012|T102|strict|38074-1|LNC|Ribs anterior - left X-ray|Ribs anterior - left X-ray
C2826012|T102|strict|37963-6|LNC|Ribs anterior - right X-ray|Ribs anterior - right X-ray
C2826012|T102|strict|38868-6|LNC|Ribs anterior and posterior - left X-ray|Ribs anterior and posterior - left X-ray
C2826012|T102|strict|37962-8|LNC|Ribs anterior and posterior - right X-ray|Ribs anterior and posterior - right X-ray
C2826012|T102|strict|26151-1|LNC|Ribs - bilateral X-ray|Ribs - bilateral X-ray
C2826012|T102|strict|69071-9|LNC|Ribs - bilateral and Chest X-ray|Ribs - bilateral and Chest X-ray
C2826012|T102|strict|26152-9|LNC|Ribs - left X-ray|Ribs - left X-ray
C2826012|T102|strict|39326-4|LNC|Ribs - left and Chest X-ray|Ribs - left and Chest X-ray
C2826012|T102|strict|38866-0|LNC|Ribs lower - left X-ray|Ribs lower - left X-ray
C2826012|T102|strict|39489-0|LNC|Ribs lower posterior X-ray|Ribs lower posterior X-ray
C2826012|T102|strict|42381-4|LNC|Ribs lower posterior - left X-ray|Ribs lower posterior - left X-ray
C2826012|T102|strict|39493-2|LNC|Ribs lower posterior - right X-ray|Ribs lower posterior - right X-ray
C2826012|T102|strict|37960-2|LNC|Ribs lower - right X-ray|Ribs lower - right X-ray
C2826012|T102|strict|37938-8|LNC|Ribs posterior X-ray|Ribs posterior X-ray
C2826012|T102|strict|39352-0|LNC|Ribs posterior - bilateral X-ray|Ribs posterior - bilateral X-ray
C2826012|T102|strict|38869-4|LNC|Ribs posterior - left X-ray|Ribs posterior - left X-ray
C2826012|T102|strict|37964-4|LNC|Ribs posterior - right X-ray|Ribs posterior - right X-ray
C2826012|T102|strict|26153-7|LNC|Ribs - right X-ray|Ribs - right X-ray
C2826012|T102|strict|39351-2|LNC|Ribs upper anterior and posterior - left X-ray|Ribs upper anterior and posterior - left X-ray
C2826012|T102|strict|39491-6|LNC|Ribs upper anterior and posterior - right X-ray|Ribs upper anterior and posterior - right X-ray
C2826012|T102|strict|38867-8|LNC|Ribs upper - left X-ray|Ribs upper - left X-ray
C2826012|T102|strict|39353-8|LNC|Ribs upper posterior - left X-ray|Ribs upper posterior - left X-ray
C2826012|T102|strict|39492-4|LNC|Ribs upper posterior - right X-ray|Ribs upper posterior - right X-ray
C2826012|T102|strict|37961-0|LNC|Ribs upper - right X-ray|Ribs upper - right X-ray
C2826012|T102|strict|24900-3|LNC|Sacroiliac Joint X-ray|Sacroiliac Joint X-ray
C2826012|T102|strict|36633-6|LNC|Sacroiliac joint - bilateral X-ray|Sacroiliac joint - bilateral X-ray
C2826012|T102|strict|36634-4|LNC|Sacroiliac joint - left X-ray|Sacroiliac joint - left X-ray
C2826012|T102|strict|37786-1|LNC|Sacroiliac joint - right X-ray|Sacroiliac joint - right X-ray
C2826012|T102|strict|30884-1|LNC|Sacrum X-ray|Sacrum X-ray
C2826012|T102|strict|24665-2|LNC|Sacrum and Coccyx X-ray|Sacrum and Coccyx X-ray
C2826012|T102|strict|39058-3|LNC|Salivary gland X-ray|Salivary gland X-ray
C2826012|T102|strict|24903-7|LNC|Scapula X-ray|Scapula X-ray
C2826012|T102|strict|26154-5|LNC|Scapula - bilateral X-ray|Scapula - bilateral X-ray
C2826012|T102|strict|26155-2|LNC|Scapula - left X-ray|Scapula - left X-ray
C2826012|T102|strict|26156-0|LNC|Scapula - right X-ray|Scapula - right X-ray
C2826012|T102|strict|42159-4|LNC|Sella turcica X-ray|Sella turcica X-ray
C2826012|T102|strict|24909-4|LNC|Shoulder X-ray|Shoulder X-ray
C2826012|T102|strict|26157-8|LNC|Shoulder - bilateral X-ray|Shoulder - bilateral X-ray
C2826012|T102|strict|26158-6|LNC|Shoulder - left X-ray|Shoulder - left X-ray
C2826012|T102|strict|26159-4|LNC|Shoulder - right X-ray|Shoulder - right X-ray
C2826012|T102|strict|42160-2|LNC|Shunt X-ray|Shunt X-ray
C2826012|T102|strict|24911-0|LNC|Shunt Fluoroscopy|Shunt Fluoroscopy
C2826012|T102|strict|24916-9|LNC|Sinuses X-ray|Sinuses X-ray
C2826012|T102|strict|28564-3|LNC|Skull X-ray|Skull X-ray
C2826012|T102|strict|48697-7|LNC|Skull.base X-ray|Skull.base X-ray
C2826012|T102|strict|37338-1|LNC|Skull and Facial bones and Mandible X-ray|Skull and Facial bones and Mandible X-ray
C2826012|T102|strict|28613-8|LNC|Spine X-ray|Spine X-ray
C2826012|T102|strict|24946-6|LNC|Spine Cervical X-ray|Spine Cervical X-ray
C2826012|T102|strict|36640-1|LNC|Spine Cervical Fluoroscopy|Spine Cervical Fluoroscopy
C2826012|T102|strict|43538-8|LNC|Spine Cervical Fluoroscopy video|Spine Cervical Fluoroscopy video
C2826012|T102|strict|37481-9|LNC|Spine Cervical and Spine Thoracic X-ray|Spine Cervical and Spine Thoracic X-ray
C2826012|T102|strict|38008-9|LNC|Spine Cervical and Thoracic and Lumbar X-ray|Spine Cervical and Thoracic and Lumbar X-ray
C2826012|T102|strict|43781-4|LNC|Spine Cervicothoracic Junction X-ray|Spine Cervicothoracic Junction X-ray
C2826012|T102|strict|24972-2|LNC|Spine Lumbar X-ray|Spine Lumbar X-ray
C2826012|T102|strict|43536-2|LNC|Spine Lumbar Fluoroscopy video|Spine Lumbar Fluoroscopy video
C2826012|T102|strict|24975-5|LNC|Spine.lumbar and Sacroiliac joint - bilateral X-ray|Spine.lumbar and Sacroiliac joint - bilateral X-ray
C2826012|T102|strict|37340-7|LNC|Spine Lumbar and Sacrum X-ray|Spine Lumbar and Sacrum X-ray
C2826012|T102|strict|37341-5|LNC|Spine Lumbar and Sacrum and Coccyx X-ray|Spine Lumbar and Sacrum and Coccyx X-ray
C2826012|T102|strict|37342-3|LNC|Spine Lumbar and Sacrum and Sacroiliac Joint and Coccyx X-ray|Spine Lumbar and Sacrum and Sacroiliac Joint and Coccyx X-ray
C2826012|T102|strict|46340-6|LNC|Spine Lumbosacral Junction X-ray|Spine Lumbosacral Junction X-ray
C2826012|T102|strict|24983-9|LNC|Spine Thoracic X-ray|Spine Thoracic X-ray
C2826012|T102|strict|42692-4|LNC|Spine Thoracic and Lumbar X-ray|Spine Thoracic and Lumbar X-ray
C2826012|T102|strict|37975-0|LNC|Spine Thoracolumbar Junction X-ray|Spine Thoracolumbar Junction X-ray
C2826012|T102|strict|37323-3|LNC|Sternoclavicular joint - bilateral X-ray|Sternoclavicular joint - bilateral X-ray
C2826012|T102|strict|37324-1|LNC|Sternoclavicular joint - left X-ray|Sternoclavicular joint - left X-ray
C2826012|T102|strict|37965-1|LNC|Sternoclavicular joint - right X-ray|Sternoclavicular joint - right X-ray
C2826012|T102|strict|24993-8|LNC|Sternoclavicular Joints X-ray|Sternoclavicular Joints X-ray
C2826012|T102|strict|24994-6|LNC|Sternum X-ray|Sternum X-ray
C2826012|T102|strict|72876-6|LNC|Surgical specimen X-ray|Surgical specimen X-ray
C2826012|T102|strict|25000-1|LNC|Temporomandibular joint X-ray|Temporomandibular joint X-ray
C2826012|T102|strict|37325-8|LNC|Temporomandibular joint - bilateral X-ray|Temporomandibular joint - bilateral X-ray
C2826012|T102|strict|30889-0|LNC|Temporomandibular joint - left X-ray|Temporomandibular joint - left X-ray
C2826012|T102|strict|30890-8|LNC|Temporomandibular joint - right X-ray|Temporomandibular joint - right X-ray
C2826012|T102|strict|25006-8|LNC|Thumb X-ray|Thumb X-ray
C2826012|T102|strict|26160-2|LNC|Thumb - bilateral X-ray|Thumb - bilateral X-ray
C2826012|T102|strict|26161-0|LNC|Thumb - left X-ray|Thumb - left X-ray
C2826012|T102|strict|26162-8|LNC|Thumb - right X-ray|Thumb - right X-ray
C2826012|T102|strict|26163-6|LNC|Tibia - bilateral and Fibula - bilateral X-ray|Tibia - bilateral and Fibula - bilateral X-ray
C2826012|T102|strict|26164-4|LNC|Tibia - left and Fibula - left X-ray|Tibia - left and Fibula - left X-ray
C2826012|T102|strict|26165-1|LNC|Tibia - right and Fibula - right X-ray|Tibia - right and Fibula - right X-ray
C2826012|T102|strict|25011-8|LNC|Tibia and Fibula X-ray|Tibia and Fibula X-ray
C2826012|T102|strict|37530-3|LNC|Toe fifth - left X-ray|Toe fifth - left X-ray
C2826012|T102|strict|38151-7|LNC|Toe fifth - right X-ray|Toe fifth - right X-ray
C2826012|T102|strict|37531-1|LNC|Toe fourth - left X-ray|Toe fourth - left X-ray
C2826012|T102|strict|38150-9|LNC|Toe fourth - right X-ray|Toe fourth - right X-ray
C2826012|T102|strict|37534-5|LNC|Toe second - left X-ray|Toe second - left X-ray
C2826012|T102|strict|38148-3|LNC|Toe second - right X-ray|Toe second - right X-ray
C2826012|T102|strict|37535-2|LNC|Toe third - left X-ray|Toe third - left X-ray
C2826012|T102|strict|38149-1|LNC|Toe third - right X-ray|Toe third - right X-ray
C2826012|T102|strict|25013-4|LNC|Toes X-ray|Toes X-ray
C2826012|T102|strict|26166-9|LNC|Toes - bilateral X-ray|Toes - bilateral X-ray
C2826012|T102|strict|26167-7|LNC|Toes - left X-ray|Toes - left X-ray
C2826012|T102|strict|26168-5|LNC|Toes - right X-ray|Toes - right X-ray
C2826012|T102|strict|44238-4|LNC|Trachea X-ray|Trachea X-ray
C2826012|T102|strict|48464-2|LNC|Trachea Fluoroscopy|Trachea Fluoroscopy
C2826012|T102|strict|24689-2|LNC|Upper extremity X-ray|Upper extremity X-ray
C2826012|T102|strict|26115-6|LNC|Upper extremity - bilateral X-ray|Upper extremity - bilateral X-ray
C2826012|T102|strict|26116-4|LNC|Upper extremity - left X-ray|Upper extremity - left X-ray
C2826012|T102|strict|26117-2|LNC|Upper extremity - right X-ray|Upper extremity - right X-ray
C2826012|T102|strict|24619-9|LNC|Wrist X-ray|Wrist X-ray
C2826012|T102|strict|26169-3|LNC|Wrist - bilateral X-ray|Wrist - bilateral X-ray
C2826012|T102|strict|26170-1|LNC|Wrist - left X-ray|Wrist - left X-ray
C2826012|T102|strict|51392-9|LNC|Wrist - left and Hand - left X-ray|Wrist - left and Hand - left X-ray
C2826012|T102|strict|26171-9|LNC|Wrist - right X-ray|Wrist - right X-ray
C2826012|T102|strict|51388-7|LNC|Wrist - right and Hand - right X-ray|Wrist - right and Hand - right X-ray
C2826012|T102|strict|43468-8|LNC|Unspecified body region X-ray|Unspecified body region X-ray
C2826012|T102|strict|49512-7|LNC|Unspecified body region Fluoroscopy|Unspecified body region Fluoroscopy
C2826012|T102|strict|25074-6|LNC|Zygomatic arch X-ray|Zygomatic arch X-ray
C2826012|T102|strict|26172-7|LNC|Zygomatic arch - bilateral X-ray|Zygomatic arch - bilateral X-ray
C2826012|T102|strict|26173-5|LNC|Zygomatic arch - left X-ray|Zygomatic arch - left X-ray
C2826012|T102|strict|26174-3|LNC|Zygomatic arch - right X-ray|Zygomatic arch - right X-ray
C2826012|T102|strict|51387-9|LNC|Knee - bilateral X-ray and (AP view standing)|Knee - bilateral X-ray and (AP view standing)
C2826012|T102|strict|39370-2|LNC|Ankle - right X-ray and (view W manual stress)|Ankle - right X-ray and (view W manual stress)
C2826012|T102|strict|30635-7|LNC|Gastrointestine upper Fluoroscopy and AP W contrast PO|Gastrointestine upper Fluoroscopy and AP W contrast PO
C2826012|T102|strict|42162-8|LNC|Gastrointestine upper Fluoroscopy and AP W water soluble contrast PO|Gastrointestine upper Fluoroscopy and AP W water soluble contrast PO
C2826012|T102|strict|39400-7|LNC|Wrist - right X-ray and carpal tunnel|Wrist - right X-ray and carpal tunnel
C2826012|T102|strict|69131-1|LNC|Hip X-ray and Danelius Miller|Hip X-ray and Danelius Miller
C2826012|T102|strict|69140-2|LNC|Hip - left X-ray and Danelius Miller|Hip - left X-ray and Danelius Miller
C2826012|T102|strict|39513-7|LNC|Hip - right X-ray and Danelius Miller|Hip - right X-ray and Danelius Miller
C2826012|T102|strict|39360-3|LNC|Pelvis X-ray and inlet and outlet|Pelvis X-ray and inlet and outlet
C2826012|T102|strict|69059-4|LNC|Hip - bilateral X-ray and lateral crosstable|Hip - bilateral X-ray and lateral crosstable
C2826012|T102|strict|69139-4|LNC|Hip - left X-ray and lateral crosstable|Hip - left X-ray and lateral crosstable
C2826012|T102|strict|39377-7|LNC|Hip - right X-ray and lateral crosstable|Hip - right X-ray and lateral crosstable
C2826012|T102|strict|37583-2|LNC|Pelvis and Hip - bilateral X-ray and lateral frog|Pelvis and Hip - bilateral X-ray and lateral frog
C2826012|T102|strict|39372-8|LNC|Ankle - right X-ray and Mortise|Ankle - right X-ray and Mortise
C2826012|T102|strict|39373-6|LNC|Elbow - right X-ray and oblique|Elbow - right X-ray and oblique
C2826012|T102|strict|39390-0|LNC|Knee - right X-ray and oblique|Knee - right X-ray and oblique
C2826012|T102|strict|39511-1|LNC|Pelvis X-ray and oblique|Pelvis X-ray and oblique
C2826012|T102|strict|39376-9|LNC|Radius - right and Ulna - right X-ray and oblique|Radius - right and Ulna - right X-ray and oblique
C2826012|T102|strict|42164-4|LNC|Spine Cervical X-ray and oblique|Spine Cervical X-ray and oblique
C2826012|T102|strict|42163-6|LNC|Spine Lumbar X-ray and oblique|Spine Lumbar X-ray and oblique
C2826012|T102|strict|39414-8|LNC|Spine Thoracic X-ray and oblique|Spine Thoracic X-ray and oblique
C2826012|T102|strict|39398-3|LNC|Tibia - right and Fibula - right X-ray and oblique|Tibia - right and Fibula - right X-ray and oblique
C2826012|T102|strict|69056-0|LNC|Elbow - bilateral X-ray and obliques|Elbow - bilateral X-ray and obliques
C2826012|T102|strict|41811-1|LNC|Ribs - bilateral and Chest X-ray and PA chest|Ribs - bilateral and Chest X-ray and PA chest
C2826012|T102|strict|41832-7|LNC|Ribs - left and Chest X-ray and PA chest|Ribs - left and Chest X-ray and PA chest
C2826012|T102|strict|42010-9|LNC|Ribs - right and Chest X-ray and PA chest|Ribs - right and Chest X-ray and PA chest
C2826012|T102|strict|42165-1|LNC|Ribs and Chest X-ray and PA chest|Ribs and Chest X-ray and PA chest
C2826012|T102|strict|46389-3|LNC|Elbow - bilateral X-ray and radial head capitellar|Elbow - bilateral X-ray and radial head capitellar
C2826012|T102|strict|39391-8|LNC|Knee - right X-ray and Sunrise|Knee - right X-ray and Sunrise
C2826012|T102|strict|39412-2|LNC|Spine Thoracic X-ray and Swimmers|Spine Thoracic X-ray and Swimmers
C2826012|T102|strict|69148-5|LNC|Knee - left X-ray and tunnel|Knee - left X-ray and tunnel
C2826012|T102|strict|39389-2|LNC|Knee - right X-ray and tunnel|Knee - right X-ray and tunnel
C2826012|T102|strict|30694-4|LNC|Thyroid Scan and uptake.single|Thyroid Scan and uptake.single
C2826012|T102|strict|42271-7|LNC|Thyroid Scan and uptake W I-123 IV|Thyroid Scan and uptake W I-123 IV
C2826012|T102|strict|60527-9|LNC|Thyroid Scan and uptake W I-123 PO|Thyroid Scan and uptake W I-123 PO
C2826012|T102|strict|25008-4|LNC|Thyroid Scan and uptake W I-131 IV|Thyroid Scan and uptake W I-131 IV
C2826012|T102|strict|69236-8|LNC|Thyroid Scan and uptake W I-131 PO|Thyroid Scan and uptake W I-131 PO
C2826012|T102|strict|43672-5|LNC|Thyroid Scan and uptake|Thyroid Scan and uptake
C2826012|T102|strict|44147-7|LNC|Thyroid Scan and uptake W Tc-99m pertechnetate IV|Thyroid Scan and uptake W Tc-99m pertechnetate IV
C2826012|T102|strict|42405-1|LNC|Knee X-ray (AP^standing) and (lateral^W hyperextension)|Knee X-ray (AP^standing) and (lateral^W hyperextension)
C2826012|T102|strict|42401-0|LNC|Spine Lumbar X-ray (AP W R-bending and W L-bending and WO bending) and Lateral|Spine Lumbar X-ray (AP W R-bending and W L-bending and WO bending) and Lateral
C2826012|T102|strict|42411-9|LNC|Spine Lumbar X-ray (AP^W R-bending and W L-bending) and (lateral^W flexion and W extension)|Spine Lumbar X-ray (AP^W R-bending and W L-bending) and (lateral^W flexion and W extension)
C2826012|T102|strict|39392-6|LNC|Shoulder - right X-ray (W internal rotation and W external rotation) and axillary|Shoulder - right X-ray (W internal rotation and W external rotation) and axillary
C2826012|T102|strict|44199-8|LNC|Facial bones X-ray 1 or 2 views|Facial bones X-ray 1 or 2 views
C2826012|T102|strict|44198-0|LNC|Knee X-ray 1 or 2 views|Knee X-ray 1 or 2 views
C2826012|T102|strict|47373-6|LNC|Knee - left X-ray 1 or 2 views|Knee - left X-ray 1 or 2 views
C2826012|T102|strict|47375-1|LNC|Knee - right X-ray 1 or 2 views|Knee - right X-ray 1 or 2 views
C2826012|T102|strict|43521-4|LNC|Mandible X-ray 1 or 2 views|Mandible X-ray 1 or 2 views
C2826012|T102|strict|47983-2|LNC|Mastoid - bilateral X-ray 1 or 2 views|Mastoid - bilateral X-ray 1 or 2 views
C2826012|T102|strict|48489-9|LNC|Mastoid - left X-ray 1 or 2 views|Mastoid - left X-ray 1 or 2 views
C2826012|T102|strict|48488-1|LNC|Mastoid - right X-ray 1 or 2 views|Mastoid - right X-ray 1 or 2 views
C2826012|T102|strict|43522-2|LNC|Pelvis X-ray 1 or 2 views|Pelvis X-ray 1 or 2 views
C2826012|T102|strict|48467-5|LNC|Sacroiliac Joint X-ray 1 or 2 views|Sacroiliac Joint X-ray 1 or 2 views
C2826012|T102|strict|43523-0|LNC|Sinuses X-ray 1 or 2 views|Sinuses X-ray 1 or 2 views
C2826012|T102|strict|44202-0|LNC|Knee X-ray 1 or 2 views portable|Knee X-ray 1 or 2 views portable
C2826012|T102|strict|44201-2|LNC|Pelvis X-ray 1 or 2 views portable|Pelvis X-ray 1 or 2 views portable
C2826012|T102|strict|36641-9|LNC|Abdomen X-ray 2 views|Abdomen X-ray 2 views
C2826012|T102|strict|37064-3|LNC|Acetabulum - left X-ray 2 views|Acetabulum - left X-ray 2 views
C2826012|T102|strict|37664-0|LNC|Acetabulum - right X-ray 2 views|Acetabulum - right X-ray 2 views
C2826012|T102|strict|36665-8|LNC|Acromioclavicular joint - left X-ray 2 views|Acromioclavicular joint - left X-ray 2 views
C2826012|T102|strict|37661-6|LNC|Acromioclavicular joint - right X-ray 2 views|Acromioclavicular joint - right X-ray 2 views
C2826012|T102|strict|24540-7|LNC|Ankle X-ray 2 views|Ankle X-ray 2 views
C2826012|T102|strict|26385-5|LNC|Ankle - bilateral X-ray 2 views|Ankle - bilateral X-ray 2 views
C2826012|T102|strict|26386-3|LNC|Ankle - left X-ray 2 views|Ankle - left X-ray 2 views
C2826012|T102|strict|26387-1|LNC|Ankle - right X-ray 2 views|Ankle - right X-ray 2 views
C2826012|T102|strict|36642-7|LNC|Breast - left Mammogram 2 views|Breast - left Mammogram 2 views
C2826012|T102|strict|37768-9|LNC|Breast - right Mammogram 2 views|Breast - right Mammogram 2 views
C2826012|T102|strict|36661-7|LNC|Calcaneus X-ray 2 views|Calcaneus X-ray 2 views
C2826012|T102|strict|48433-7|LNC|Calcaneus - bilateral X-ray 2 views|Calcaneus - bilateral X-ray 2 views
C2826012|T102|strict|36662-5|LNC|Calcaneus - left X-ray 2 views|Calcaneus - left X-ray 2 views
C2826012|T102|strict|37718-4|LNC|Calcaneus - right X-ray 2 views|Calcaneus - right X-ray 2 views
C2826012|T102|strict|36643-5|LNC|Chest X-ray 2 views|Chest X-ray 2 views
C2826012|T102|strict|36644-3|LNC|Chest Fluoroscopy 2 views|Chest Fluoroscopy 2 views
C2826012|T102|strict|36645-0|LNC|Clavicle X-ray 2 views|Clavicle X-ray 2 views
C2826012|T102|strict|36646-8|LNC|Clavicle - left X-ray 2 views|Clavicle - left X-ray 2 views
C2826012|T102|strict|37679-8|LNC|Clavicle - right X-ray 2 views|Clavicle - right X-ray 2 views
C2826012|T102|strict|36647-6|LNC|Coccyx X-ray 2 views|Coccyx X-ray 2 views
C2826012|T102|strict|36648-4|LNC|Elbow X-ray 2 views|Elbow X-ray 2 views
C2826012|T102|strict|36649-2|LNC|Elbow - bilateral X-ray 2 views|Elbow - bilateral X-ray 2 views
C2826012|T102|strict|36650-0|LNC|Elbow - left X-ray 2 views|Elbow - left X-ray 2 views
C2826012|T102|strict|37681-4|LNC|Elbow - right X-ray 2 views|Elbow - right X-ray 2 views
C2826012|T102|strict|36652-6|LNC|Femur X-ray 2 views|Femur X-ray 2 views
C2826012|T102|strict|36653-4|LNC|Femur - bilateral X-ray 2 views|Femur - bilateral X-ray 2 views
C2826012|T102|strict|36654-2|LNC|Femur - left X-ray 2 views|Femur - left X-ray 2 views
C2826012|T102|strict|37690-5|LNC|Femur - right X-ray 2 views|Femur - right X-ray 2 views
C2826012|T102|strict|36655-9|LNC|Finger X-ray 2 views|Finger X-ray 2 views
C2826012|T102|strict|36656-7|LNC|Finger - left X-ray 2 views|Finger - left X-ray 2 views
C2826012|T102|strict|37694-7|LNC|Finger - right X-ray 2 views|Finger - right X-ray 2 views
C2826012|T102|strict|30784-3|LNC|Foot X-ray 2 views|Foot X-ray 2 views
C2826012|T102|strict|36657-5|LNC|Foot - bilateral X-ray 2 views|Foot - bilateral X-ray 2 views
C2826012|T102|strict|38846-2|LNC|Foot - left X-ray 2 views|Foot - left X-ray 2 views
C2826012|T102|strict|37697-0|LNC|Foot - right X-ray 2 views|Foot - right X-ray 2 views
C2826012|T102|strict|24721-3|LNC|Hand X-ray 2 views|Hand X-ray 2 views
C2826012|T102|strict|26388-9|LNC|Hand - bilateral X-ray 2 views|Hand - bilateral X-ray 2 views
C2826012|T102|strict|26389-7|LNC|Hand - left X-ray 2 views|Hand - left X-ray 2 views
C2826012|T102|strict|26390-5|LNC|Hand - right X-ray 2 views|Hand - right X-ray 2 views
C2826012|T102|strict|36663-3|LNC|Hip X-ray 2 views|Hip X-ray 2 views
C2826012|T102|strict|69058-6|LNC|Hip - bilateral X-ray 2 views|Hip - bilateral X-ray 2 views
C2826012|T102|strict|36664-1|LNC|Hip - left X-ray 2 views|Hip - left X-ray 2 views
C2826012|T102|strict|37721-8|LNC|Hip - right X-ray 2 views|Hip - right X-ray 2 views
C2826012|T102|strict|24765-0|LNC|Humerus X-ray 2 views|Humerus X-ray 2 views
C2826012|T102|strict|26391-3|LNC|Humerus - bilateral X-ray 2 views|Humerus - bilateral X-ray 2 views
C2826012|T102|strict|26392-1|LNC|Humerus - left X-ray 2 views|Humerus - left X-ray 2 views
C2826012|T102|strict|26393-9|LNC|Humerus - right X-ray 2 views|Humerus - right X-ray 2 views
C2826012|T102|strict|24806-2|LNC|Knee X-ray 2 views|Knee X-ray 2 views
C2826012|T102|strict|26394-7|LNC|Knee - bilateral X-ray 2 views|Knee - bilateral X-ray 2 views
C2826012|T102|strict|26395-4|LNC|Knee - left X-ray 2 views|Knee - left X-ray 2 views
C2826012|T102|strict|26396-2|LNC|Knee - right X-ray 2 views|Knee - right X-ray 2 views
C2826012|T102|strict|36651-8|LNC|Lower extremity X-ray 2 views|Lower extremity X-ray 2 views
C2826012|T102|strict|69257-4|LNC|Lower extremity - right X-ray 2 views|Lower extremity - right X-ray 2 views
C2826012|T102|strict|24861-7|LNC|Patella X-ray 2 views|Patella X-ray 2 views
C2826012|T102|strict|26397-0|LNC|Patella - bilateral X-ray 2 views|Patella - bilateral X-ray 2 views
C2826012|T102|strict|26398-8|LNC|Patella - left X-ray 2 views|Patella - left X-ray 2 views
C2826012|T102|strict|26399-6|LNC|Patella - right X-ray 2 views|Patella - right X-ray 2 views
C2826012|T102|strict|37617-8|LNC|Pelvis X-ray 2 views|Pelvis X-ray 2 views
C2826012|T102|strict|42685-8|LNC|Pelvis and Hip - left X-ray 2 views|Pelvis and Hip - left X-ray 2 views
C2826012|T102|strict|42686-6|LNC|Pelvis and Hip - right X-ray 2 views|Pelvis and Hip - right X-ray 2 views
C2826012|T102|strict|36659-1|LNC|Radius - bilateral and Ulna - bilateral X-ray 2 views|Radius - bilateral and Ulna - bilateral X-ray 2 views
C2826012|T102|strict|36660-9|LNC|Radius - left and Ulna.left X-ray 2 views|Radius - left and Ulna.left X-ray 2 views
C2826012|T102|strict|37707-7|LNC|Radius - right and Ulna - right X-ray 2 views|Radius - right and Ulna - right X-ray 2 views
C2826012|T102|strict|36658-3|LNC|Radius and Ulna X-ray 2 views|Radius and Ulna X-ray 2 views
C2826012|T102|strict|39060-9|LNC|Ribs X-ray 2 views|Ribs X-ray 2 views
C2826012|T102|strict|42687-4|LNC|Ribs - bilateral X-ray 2 views|Ribs - bilateral X-ray 2 views
C2826012|T102|strict|37066-8|LNC|Ribs - left X-ray 2 views|Ribs - left X-ray 2 views
C2826012|T102|strict|37780-4|LNC|Ribs - right X-ray 2 views|Ribs - right X-ray 2 views
C2826012|T102|strict|37651-7|LNC|Sacrum X-ray 2 views|Sacrum X-ray 2 views
C2826012|T102|strict|44179-0|LNC|Sacrum and Coccyx X-ray 2 views|Sacrum and Coccyx X-ray 2 views
C2826012|T102|strict|37655-8|LNC|Scapula X-ray 2 views|Scapula X-ray 2 views
C2826012|T102|strict|36666-6|LNC|Scapula - left X-ray 2 views|Scapula - left X-ray 2 views
C2826012|T102|strict|37787-9|LNC|Scapula - right X-ray 2 views|Scapula - right X-ray 2 views
C2826012|T102|strict|42435-8|LNC|Sella turcica X-ray 2 views|Sella turcica X-ray 2 views
C2826012|T102|strict|37840-6|LNC|Shoulder X-ray 2 views|Shoulder X-ray 2 views
C2826012|T102|strict|36667-4|LNC|Shoulder - bilateral X-ray 2 views|Shoulder - bilateral X-ray 2 views
C2826012|T102|strict|36668-2|LNC|Shoulder - left X-ray 2 views|Shoulder - left X-ray 2 views
C2826012|T102|strict|37793-7|LNC|Shoulder - right X-ray 2 views|Shoulder - right X-ray 2 views
C2826012|T102|strict|37853-9|LNC|Sinuses X-ray 2 views|Sinuses X-ray 2 views
C2826012|T102|strict|37867-9|LNC|Skull X-ray 2 views|Skull X-ray 2 views
C2826012|T102|strict|37879-4|LNC|Spine X-ray 2 views|Spine X-ray 2 views
C2826012|T102|strict|36669-0|LNC|Spine Cervical X-ray 2 views|Spine Cervical X-ray 2 views
C2826012|T102|strict|43784-8|LNC|Spine Cervical and Thoracic and Lumbar X-ray 2 views|Spine Cervical and Thoracic and Lumbar X-ray 2 views
C2826012|T102|strict|36670-8|LNC|Spine Lumbar X-ray 2 views|Spine Lumbar X-ray 2 views
C2826012|T102|strict|37905-7|LNC|Spine Thoracic X-ray 2 views|Spine Thoracic X-ray 2 views
C2826012|T102|strict|24984-7|LNC|Spine Thoracic and Lumbar X-ray 2 views|Spine Thoracic and Lumbar X-ray 2 views
C2826012|T102|strict|69273-1|LNC|Spine Thoracolumbar Junction X-ray 2 views|Spine Thoracolumbar Junction X-ray 2 views
C2826012|T102|strict|37883-6|LNC|Sternum X-ray 2 views|Sternum X-ray 2 views
C2826012|T102|strict|36671-6|LNC|Tibia - bilateral and Fibula - bilateral X-ray 2 views|Tibia - bilateral and Fibula - bilateral X-ray 2 views
C2826012|T102|strict|36672-4|LNC|Tibia - left and Fibula - left X-ray 2 views|Tibia - left and Fibula - left X-ray 2 views
C2826012|T102|strict|37815-8|LNC|Tibia - right and Fibula - right X-ray 2 views|Tibia - right and Fibula - right X-ray 2 views
C2826012|T102|strict|37895-0|LNC|Tibia and Fibula X-ray 2 views|Tibia and Fibula X-ray 2 views
C2826012|T102|strict|37902-4|LNC|Toes X-ray 2 views|Toes X-ray 2 views
C2826012|T102|strict|37348-0|LNC|Toes - bilateral X-ray 2 views|Toes - bilateral X-ray 2 views
C2826012|T102|strict|36673-2|LNC|Toes - left X-ray 2 views|Toes - left X-ray 2 views
C2826012|T102|strict|37821-6|LNC|Toes - right X-ray 2 views|Toes - right X-ray 2 views
C2826012|T102|strict|37922-2|LNC|Upper extremity X-ray 2 views|Upper extremity X-ray 2 views
C2826012|T102|strict|37925-5|LNC|Wrist X-ray 2 views|Wrist X-ray 2 views
C2826012|T102|strict|37482-7|LNC|Wrist - bilateral X-ray 2 views|Wrist - bilateral X-ray 2 views
C2826012|T102|strict|37483-5|LNC|Wrist - left X-ray 2 views|Wrist - left X-ray 2 views
C2826012|T102|strict|37826-5|LNC|Wrist - right X-ray 2 views|Wrist - right X-ray 2 views
C2826012|T102|strict|69305-1|LNC|Zygomatic arch X-ray 2 views|Zygomatic arch X-ray 2 views
C2826012|T102|strict|42430-9|LNC|Knee - right X-ray 2 views and (views standing)|Knee - right X-ray 2 views and (views standing)
C2826012|T102|strict|42009-1|LNC|Chest X-ray 2 views and apical|Chest X-ray 2 views and apical
C2826012|T102|strict|39378-5|LNC|Knee - right X-ray 2 views and oblique|Knee - right X-ray 2 views and oblique
C2826012|T102|strict|48468-3|LNC|Ribs - bilateral and Chest X-ray 2 views and PA chest|Ribs - bilateral and Chest X-ray 2 views and PA chest
C2826012|T102|strict|43467-0|LNC|Chest X-ray 2 views and right oblique and left oblique|Chest X-ray 2 views and right oblique and left oblique
C2826012|T102|strict|69060-2|LNC|Knee - bilateral X-ray 2 views and Sunrise|Knee - bilateral X-ray 2 views and Sunrise
C2826012|T102|strict|69142-8|LNC|Knee - left X-ray 2 views and Sunrise|Knee - left X-ray 2 views and Sunrise
C2826012|T102|strict|39379-3|LNC|Knee - right X-ray 2 views and Sunrise|Knee - right X-ray 2 views and Sunrise
C2826012|T102|strict|39380-1|LNC|Knee - right X-ray 2 views and Sunrise and tunnel|Knee - right X-ray 2 views and Sunrise and tunnel
C2826012|T102|strict|69061-0|LNC|Knee - bilateral X-ray 2 views and tunnel|Knee - bilateral X-ray 2 views and tunnel
C2826012|T102|strict|41819-4|LNC|Knee - left X-ray 2 views and tunnel|Knee - left X-ray 2 views and tunnel
C2826012|T102|strict|39381-9|LNC|Knee - right X-ray 2 views and tunnel|Knee - right X-ray 2 views and tunnel
C2826012|T102|strict|69143-6|LNC|Knee - left X-ray 2 views and tunnel standing|Knee - left X-ray 2 views and tunnel standing
C2826012|T102|strict|39382-7|LNC|Knee - right X-ray 2 views and tunnel standing|Knee - right X-ray 2 views and tunnel standing
C2826012|T102|strict|38118-6|LNC|Neck X-ray 2 views lateral|Neck X-ray 2 views lateral
C2826012|T102|strict|38844-7|LNC|Elbow - left X-ray 2 views Oblique|Elbow - left X-ray 2 views Oblique
C2826012|T102|strict|37686-3|LNC|Elbow - right X-ray 2 views Oblique|Elbow - right X-ray 2 views Oblique
C2826012|T102|strict|38871-0|LNC|Knee - left X-ray 2 views Oblique|Knee - left X-ray 2 views Oblique
C2826012|T102|strict|38108-7|LNC|Knee - right X-ray 2 views Oblique|Knee - right X-ray 2 views Oblique
C2826012|T102|strict|38874-4|LNC|Tibia - left and Fibula - left X-ray 2 views Oblique|Tibia - left and Fibula - left X-ray 2 views Oblique
C2826012|T102|strict|38114-5|LNC|Tibia - right and Fibula - right X-ray 2 views Oblique|Tibia - right and Fibula - right X-ray 2 views Oblique
C2826012|T102|strict|44181-6|LNC|Sacroiliac Joint X-ray 2 or 3 views|Sacroiliac Joint X-ray 2 or 3 views
C2826012|T102|strict|43539-6|LNC|Spine Cervical X-ray 2 or 3 views|Spine Cervical X-ray 2 or 3 views
C2826012|T102|strict|48469-1|LNC|Spine Lumbar X-ray 2 or 3 views|Spine Lumbar X-ray 2 or 3 views
C2826012|T102|strict|39880-0|LNC|Bone Scan 2 views phase|Bone Scan 2 views phase
C2826012|T102|strict|44184-0|LNC|Elbow X-ray 2 views portable|Elbow X-ray 2 views portable
C2826012|T102|strict|44182-4|LNC|Hand X-ray 2 views portable|Hand X-ray 2 views portable
C2826012|T102|strict|44183-2|LNC|Radius and Ulna X-ray 2 views portable|Radius and Ulna X-ray 2 views portable
C2826012|T102|strict|36674-0|LNC|Spine Lumbar X-ray 2 views portable|Spine Lumbar X-ray 2 views portable
C2826012|T102|strict|37658-2|LNC|Spine Thoracic and Lumbar X-ray 2 views scoliosis|Spine Thoracic and Lumbar X-ray 2 views scoliosis
C2826012|T102|strict|38843-9|LNC|Wrist - left X-ray 2 views tunnel.carpal|Wrist - left X-ray 2 views tunnel.carpal
C2826012|T102|strict|37678-0|LNC|Wrist - right X-ray 2 views tunnel.carpal|Wrist - right X-ray 2 views tunnel.carpal
C2826012|T102|strict|42166-9|LNC|Heart Scan 2 views at rest and W Tl-201 IV|Heart Scan 2 views at rest and W Tl-201 IV
C2826012|T102|strict|38841-3|LNC|Ankle - left X-ray 2 views standing|Ankle - left X-ray 2 views standing
C2826012|T102|strict|37675-6|LNC|Ankle - right X-ray 2 views standing|Ankle - right X-ray 2 views standing
C2826012|T102|strict|37068-4|LNC|Foot - bilateral X-ray 2 views standing|Foot - bilateral X-ray 2 views standing
C2826012|T102|strict|37069-2|LNC|Foot - left X-ray 2 views standing|Foot - left X-ray 2 views standing
C2826012|T102|strict|37698-8|LNC|Foot - right X-ray 2 views standing|Foot - right X-ray 2 views standing
C2826012|T102|strict|36945-4|LNC|Knee - bilateral X-ray 2 views standing|Knee - bilateral X-ray 2 views standing
C2826012|T102|strict|38851-2|LNC|Knee - left X-ray 2 views standing|Knee - left X-ray 2 views standing
C2826012|T102|strict|37762-2|LNC|Knee - right X-ray 2 views standing|Knee - right X-ray 2 views standing
C2826012|T102|strict|36946-2|LNC|Spine Lumbar X-ray 2 views standing|Spine Lumbar X-ray 2 views standing
C2826012|T102|strict|69274-9|LNC|Spine Thoracic X-ray 2 views standing|Spine Thoracic X-ray 2 views standing
C2826012|T102|strict|38840-5|LNC|Ankle - left X-ray 2 views W manual stress|Ankle - left X-ray 2 views W manual stress
C2826012|T102|strict|37672-3|LNC|Ankle - right X-ray 2 views W manual stress|Ankle - right X-ray 2 views W manual stress
C2826012|T102|strict|37067-6|LNC|Chest X-ray 2 views W nipple markers|Chest X-ray 2 views W nipple markers
C2826012|T102|strict|36293-9|LNC|Abdomen X-ray 3 views|Abdomen X-ray 3 views
C2826012|T102|strict|37635-0|LNC|Acetabulum X-ray 3 views|Acetabulum X-ray 3 views
C2826012|T102|strict|36294-7|LNC|Ankle X-ray 3 views|Ankle X-ray 3 views
C2826012|T102|strict|36295-4|LNC|Ankle - bilateral X-ray 3 views|Ankle - bilateral X-ray 3 views
C2826012|T102|strict|36296-2|LNC|Ankle - left X-ray 3 views|Ankle - left X-ray 3 views
C2826012|T102|strict|37665-7|LNC|Ankle - right X-ray 3 views|Ankle - right X-ray 3 views
C2826012|T102|strict|36298-8|LNC|Chest X-ray 3 views|Chest X-ray 3 views
C2826012|T102|strict|36299-6|LNC|Elbow X-ray 3 views|Elbow X-ray 3 views
C2826012|T102|strict|36300-2|LNC|Elbow - bilateral X-ray 3 views|Elbow - bilateral X-ray 3 views
C2826012|T102|strict|36301-0|LNC|Elbow - left X-ray 3 views|Elbow - left X-ray 3 views
C2826012|T102|strict|37682-2|LNC|Elbow - right X-ray 3 views|Elbow - right X-ray 3 views
C2826012|T102|strict|36297-0|LNC|Facial bones X-ray 3 views|Facial bones X-ray 3 views
C2826012|T102|strict|36302-8|LNC|Femur X-ray 3 views|Femur X-ray 3 views
C2826012|T102|strict|36303-6|LNC|Finger X-ray 3 views|Finger X-ray 3 views
C2826012|T102|strict|36304-4|LNC|Finger - left X-ray 3 views|Finger - left X-ray 3 views
C2826012|T102|strict|37695-4|LNC|Finger - right X-ray 3 views|Finger - right X-ray 3 views
C2826012|T102|strict|36305-1|LNC|Foot X-ray 3 views|Foot X-ray 3 views
C2826012|T102|strict|36306-9|LNC|Foot - bilateral X-ray 3 views|Foot - bilateral X-ray 3 views
C2826012|T102|strict|36307-7|LNC|Foot - left X-ray 3 views|Foot - left X-ray 3 views
C2826012|T102|strict|37699-6|LNC|Foot - right X-ray 3 views|Foot - right X-ray 3 views
C2826012|T102|strict|24722-1|LNC|Hand X-ray 3 views|Hand X-ray 3 views
C2826012|T102|strict|26379-8|LNC|Hand - bilateral X-ray 3 views|Hand - bilateral X-ray 3 views
C2826012|T102|strict|26380-6|LNC|Hand - left X-ray 3 views|Hand - left X-ray 3 views
C2826012|T102|strict|26381-4|LNC|Hand - right X-ray 3 views|Hand - right X-ray 3 views
C2826012|T102|strict|36308-5|LNC|Hip - bilateral X-ray 3 views|Hip - bilateral X-ray 3 views
C2826012|T102|strict|36309-3|LNC|Hip - left X-ray 3 views|Hip - left X-ray 3 views
C2826012|T102|strict|37722-6|LNC|Hip - right X-ray 3 views|Hip - right X-ray 3 views
C2826012|T102|strict|30788-4|LNC|Knee X-ray 3 views|Knee X-ray 3 views
C2826012|T102|strict|36310-1|LNC|Knee - bilateral X-ray 3 views|Knee - bilateral X-ray 3 views
C2826012|T102|strict|36311-9|LNC|Knee - left X-ray 3 views|Knee - left X-ray 3 views
C2826012|T102|strict|37742-4|LNC|Knee - right X-ray 3 views|Knee - right X-ray 3 views
C2826012|T102|strict|36312-7|LNC|Mandible X-ray 3 views|Mandible X-ray 3 views
C2826012|T102|strict|36838-1|LNC|Mastoid X-ray 3 views|Mastoid X-ray 3 views
C2826012|T102|strict|48470-9|LNC|Mastoid - left X-ray 3 views|Mastoid - left X-ray 3 views
C2826012|T102|strict|48471-7|LNC|Mastoid - right X-ray 3 views|Mastoid - right X-ray 3 views
C2826012|T102|strict|37604-6|LNC|Nasal bones X-ray 3 views|Nasal bones X-ray 3 views
C2826012|T102|strict|69261-6|LNC|Patella - right X-ray 3 views|Patella - right X-ray 3 views
C2826012|T102|strict|30766-0|LNC|Pelvis X-ray 3 views|Pelvis X-ray 3 views
C2826012|T102|strict|37256-5|LNC|Pelvis and Spine Lumbar X-ray 3 views|Pelvis and Spine Lumbar X-ray 3 views
C2826012|T102|strict|39062-5|LNC|Ribs X-ray 3 views|Ribs X-ray 3 views
C2826012|T102|strict|36313-5|LNC|Ribs - bilateral X-ray 3 views|Ribs - bilateral X-ray 3 views
C2826012|T102|strict|36314-3|LNC|Ribs - left X-ray 3 views|Ribs - left X-ray 3 views
C2826012|T102|strict|37781-2|LNC|Ribs - right X-ray 3 views|Ribs - right X-ray 3 views
C2826012|T102|strict|37648-3|LNC|Sacroiliac Joint X-ray 3 views|Sacroiliac Joint X-ray 3 views
C2826012|T102|strict|39061-7|LNC|Sacrum and Coccyx X-ray 3 views|Sacrum and Coccyx X-ray 3 views
C2826012|T102|strict|24908-6|LNC|Shoulder X-ray 3 views|Shoulder X-ray 3 views
C2826012|T102|strict|26382-2|LNC|Shoulder - bilateral X-ray 3 views|Shoulder - bilateral X-ray 3 views
C2826012|T102|strict|26383-0|LNC|Shoulder - left X-ray 3 views|Shoulder - left X-ray 3 views
C2826012|T102|strict|26384-8|LNC|Shoulder - right X-ray 3 views|Shoulder - right X-ray 3 views
C2826012|T102|strict|37854-7|LNC|Sinuses X-ray 3 views|Sinuses X-ray 3 views
C2826012|T102|strict|24918-5|LNC|Skull X-ray 3 views|Skull X-ray 3 views
C2826012|T102|strict|24941-7|LNC|Spine Cervical X-ray 3 views|Spine Cervical X-ray 3 views
C2826012|T102|strict|30775-1|LNC|Spine Lumbar X-ray 3 views|Spine Lumbar X-ray 3 views
C2826012|T102|strict|37257-3|LNC|Spine Lumbar and Sacroiliac Joint X-ray 3 views|Spine Lumbar and Sacroiliac Joint X-ray 3 views
C2826012|T102|strict|37259-9|LNC|Spine Lumbar and Sacrum X-ray 3 views|Spine Lumbar and Sacrum X-ray 3 views
C2826012|T102|strict|37260-7|LNC|Spine Lumbar and Sacrum and Coccyx X-ray 3 views|Spine Lumbar and Sacrum and Coccyx X-ray 3 views
C2826012|T102|strict|37261-5|LNC|Spine Lumbar and Sacrum and Sacroiliac Joint and Coccyx X-ray 3 views|Spine Lumbar and Sacrum and Sacroiliac Joint and Coccyx X-ray 3 views
C2826012|T102|strict|37906-5|LNC|Spine Thoracic X-ray 3 views|Spine Thoracic X-ray 3 views
C2826012|T102|strict|37881-0|LNC|Sternoclavicular Joint X-ray 3 views|Sternoclavicular Joint X-ray 3 views
C2826012|T102|strict|37888-5|LNC|Thumb X-ray 3 views|Thumb X-ray 3 views
C2826012|T102|strict|36315-0|LNC|Thumb - left X-ray 3 views|Thumb - left X-ray 3 views
C2826012|T102|strict|37812-5|LNC|Thumb - right X-ray 3 views|Thumb - right X-ray 3 views
C2826012|T102|strict|36316-8|LNC|Toes - left X-ray 3 views|Toes - left X-ray 3 views
C2826012|T102|strict|37820-8|LNC|Toes - right X-ray 3 views|Toes - right X-ray 3 views
C2826012|T102|strict|37926-3|LNC|Wrist X-ray 3 views|Wrist X-ray 3 views
C2826012|T102|strict|37454-6|LNC|Wrist - bilateral X-ray 3 views|Wrist - bilateral X-ray 3 views
C2826012|T102|strict|48738-9|LNC|Wrist - bilateral and Hand - bilateral X-ray 3 views|Wrist - bilateral and Hand - bilateral X-ray 3 views
C2826012|T102|strict|37455-3|LNC|Wrist - left X-ray 3 views|Wrist - left X-ray 3 views
C2826012|T102|strict|37827-3|LNC|Wrist - right X-ray 3 views|Wrist - right X-ray 3 views
C2826012|T102|strict|48737-1|LNC|Wrist and Hand X-ray 3 views|Wrist and Hand X-ray 3 views
C2826012|T102|strict|37933-9|LNC|Zygomatic arch X-ray 3 views|Zygomatic arch X-ray 3 views
C2826012|T102|strict|69154-3|LNC|Shoulder - left X-ray 3 views and axillary|Shoulder - left X-ray 3 views and axillary
C2826012|T102|strict|39393-4|LNC|Shoulder - right X-ray 3 views and axillary|Shoulder - right X-ray 3 views and axillary
C2826012|T102|strict|39399-1|LNC|Wrist - right X-ray 3 views and carpal tunnel|Wrist - right X-ray 3 views and carpal tunnel
C2826012|T102|strict|39364-5|LNC|Wrist - right X-ray 3 views and radial deviation|Wrist - right X-ray 3 views and radial deviation
C2826012|T102|strict|39404-9|LNC|Sinuses X-ray 3 views and submentovertex|Sinuses X-ray 3 views and submentovertex
C2826012|T102|strict|39383-5|LNC|Knee - right X-ray 3 views and Sunrise|Knee - right X-ray 3 views and Sunrise
C2826012|T102|strict|48472-5|LNC|Spine Thoracic X-ray 3 views and Swimmers|Spine Thoracic X-ray 3 views and Swimmers
C2826012|T102|strict|39365-2|LNC|Wrist - right X-ray 3 views and ulnar deviation|Wrist - right X-ray 3 views and ulnar deviation
C2826012|T102|strict|69155-0|LNC|Shoulder - left X-ray 3 views and Y|Shoulder - left X-ray 3 views and Y
C2826012|T102|strict|39394-2|LNC|Shoulder - right X-ray 3 views and Y|Shoulder - right X-ray 3 views and Y
C2826012|T102|strict|43499-3|LNC|Foot - left X-ray 3 or 4 views|Foot - left X-ray 3 or 4 views
C2826012|T102|strict|43483-7|LNC|Foot - right X-ray 3 or 4 views|Foot - right X-ray 3 or 4 views
C2826012|T102|strict|39901-4|LNC|Bone Scan 3 views phase multiple areas|Bone Scan 3 views phase multiple areas
C2826012|T102|strict|39902-2|LNC|Bone Scan 3 views phase single area|Bone Scan 3 views phase single area
C2826012|T102|strict|39882-6|LNC|Bone Scan 3 views phase whole body|Bone Scan 3 views phase whole body
C2826012|T102|strict|39883-4|LNC|Bone Scan 3 views phase|Bone Scan 3 views phase
C2826012|T102|strict|30776-9|LNC|Spine Lumbar X-ray 3 views portable|Spine Lumbar X-ray 3 views portable
C2826012|T102|strict|69151-9|LNC|Wrist - left X-ray 3 views scaphoid|Wrist - left X-ray 3 views scaphoid
C2826012|T102|strict|24778-3|LNC|Kidney - bilateral X-ray 3 views serial W and WO contrast IV|Kidney - bilateral X-ray 3 views serial W and WO contrast IV
C2826012|T102|strict|69138-6|LNC|Ankle - left X-ray 3 views standing|Ankle - left X-ray 3 views standing
C2826012|T102|strict|69254-1|LNC|Ankle - right X-ray 3 views standing|Ankle - right X-ray 3 views standing
C2826012|T102|strict|36947-0|LNC|Foot - bilateral X-ray 3 views standing|Foot - bilateral X-ray 3 views standing
C2826012|T102|strict|36948-8|LNC|Foot - left X-ray 3 views standing|Foot - left X-ray 3 views standing
C2826012|T102|strict|37700-2|LNC|Foot - right X-ray 3 views standing|Foot - right X-ray 3 views standing
C2826012|T102|strict|36949-6|LNC|Spine Lumbar X-ray 3 views standing|Spine Lumbar X-ray 3 views standing
C2826012|T102|strict|42443-2|LNC|Spine Thoracic X-ray 3 views standing|Spine Thoracic X-ray 3 views standing
C2826012|T102|strict|36317-6|LNC|Ankle X-ray 4 views|Ankle X-ray 4 views
C2826012|T102|strict|36319-2|LNC|Breast Mammogram 4 views|Breast Mammogram 4 views
C2826012|T102|strict|36320-0|LNC|Chest X-ray 4 views|Chest X-ray 4 views
C2826012|T102|strict|36321-8|LNC|Chest Fluoroscopy 4 views|Chest Fluoroscopy 4 views
C2826012|T102|strict|36322-6|LNC|Elbow - bilateral X-ray 4 views|Elbow - bilateral X-ray 4 views
C2826012|T102|strict|36323-4|LNC|Elbow - left X-ray 4 views|Elbow - left X-ray 4 views
C2826012|T102|strict|37683-0|LNC|Elbow - right X-ray 4 views|Elbow - right X-ray 4 views
C2826012|T102|strict|36318-4|LNC|Facial bones X-ray 4 views|Facial bones X-ray 4 views
C2826012|T102|strict|36324-2|LNC|Femur - left X-ray 4 views|Femur - left X-ray 4 views
C2826012|T102|strict|37691-3|LNC|Femur - right X-ray 4 views|Femur - right X-ray 4 views
C2826012|T102|strict|30789-2|LNC|Knee X-ray 4 views|Knee X-ray 4 views
C2826012|T102|strict|36325-9|LNC|Knee - bilateral X-ray 4 views|Knee - bilateral X-ray 4 views
C2826012|T102|strict|36326-7|LNC|Knee - left X-ray 4 views|Knee - left X-ray 4 views
C2826012|T102|strict|37743-2|LNC|Knee - right X-ray 4 views|Knee - right X-ray 4 views
C2826012|T102|strict|36327-5|LNC|Mandible X-ray 4 views|Mandible X-ray 4 views
C2826012|T102|strict|43534-7|LNC|Mandible - left X-ray 4 views|Mandible - left X-ray 4 views
C2826012|T102|strict|43535-4|LNC|Mandible - right X-ray 4 views|Mandible - right X-ray 4 views
C2826012|T102|strict|36839-9|LNC|Mastoid X-ray 4 views|Mastoid X-ray 4 views
C2826012|T102|strict|37609-5|LNC|Optic foramen X-ray 4 views|Optic foramen X-ray 4 views
C2826012|T102|strict|37612-9|LNC|Orbit - bilateral X-ray 4 views|Orbit - bilateral X-ray 4 views
C2826012|T102|strict|36328-3|LNC|Ribs - bilateral X-ray 4 views|Ribs - bilateral X-ray 4 views
C2826012|T102|strict|69265-7|LNC|Shoulder X-ray 4 views|Shoulder X-ray 4 views
C2826012|T102|strict|36329-1|LNC|Shoulder - bilateral X-ray 4 views|Shoulder - bilateral X-ray 4 views
C2826012|T102|strict|36330-9|LNC|Shoulder - left X-ray 4 views|Shoulder - left X-ray 4 views
C2826012|T102|strict|37794-5|LNC|Shoulder - right X-ray 4 views|Shoulder - right X-ray 4 views
C2826012|T102|strict|37855-4|LNC|Sinuses X-ray 4 views|Sinuses X-ray 4 views
C2826012|T102|strict|37868-7|LNC|Skull X-ray 4 views|Skull X-ray 4 views
C2826012|T102|strict|37876-0|LNC|Spine X-ray 4 views|Spine X-ray 4 views
C2826012|T102|strict|36331-7|LNC|Spine Cervical X-ray 4 views|Spine Cervical X-ray 4 views
C2826012|T102|strict|36332-5|LNC|Spine Lumbar X-ray 4 views|Spine Lumbar X-ray 4 views
C2826012|T102|strict|48473-3|LNC|Spine Lumbar and Sacrum X-ray 4 views|Spine Lumbar and Sacrum X-ray 4 views
C2826012|T102|strict|37907-3|LNC|Spine Thoracic X-ray 4 views|Spine Thoracic X-ray 4 views
C2826012|T102|strict|37882-8|LNC|Sternoclavicular Joint X-ray 4 views|Sternoclavicular Joint X-ray 4 views
C2826012|T102|strict|38155-8|LNC|Wrist X-ray 4 views|Wrist X-ray 4 views
C2826012|T102|strict|37070-0|LNC|Wrist - bilateral X-ray 4 views|Wrist - bilateral X-ray 4 views
C2826012|T102|strict|37071-8|LNC|Wrist - left X-ray 4 views|Wrist - left X-ray 4 views
C2826012|T102|strict|37828-1|LNC|Wrist - right X-ray 4 views|Wrist - right X-ray 4 views
C2826012|T102|strict|37934-7|LNC|Zygomatic arch X-ray 4 views|Zygomatic arch X-ray 4 views
C2826012|T102|strict|69144-4|LNC|Knee - left X-ray 4 views and AP standing|Knee - left X-ray 4 views and AP standing
C2826012|T102|strict|39384-3|LNC|Knee - right X-ray 4 views and AP standing|Knee - right X-ray 4 views and AP standing
C2826012|T102|strict|39385-0|LNC|Knee - right X-ray 4 views and oblique|Knee - right X-ray 4 views and oblique
C2826012|T102|strict|39413-0|LNC|Spine Thoracic X-ray 4 views and oblique|Spine Thoracic X-ray 4 views and oblique
C2826012|T102|strict|39099-7|LNC|Ribs - bilateral and Chest X-ray 4 views and PA chest|Ribs - bilateral and Chest X-ray 4 views and PA chest
C2826012|T102|strict|69063-6|LNC|Knee - bilateral X-ray 4 views and Sunrise and tunnel|Knee - bilateral X-ray 4 views and Sunrise and tunnel
C2826012|T102|strict|39387-6|LNC|Knee - right X-ray 4 views and Sunrise and tunnel|Knee - right X-ray 4 views and Sunrise and tunnel
C2826012|T102|strict|69145-1|LNC|Knee - left X-ray 4 views and tunnel|Knee - left X-ray 4 views and tunnel
C2826012|T102|strict|39386-8|LNC|Knee - right X-ray 4 views and tunnel|Knee - right X-ray 4 views and tunnel
C2826012|T102|strict|69062-8|LNC|Knee - bilateral X-ray 4 views standing|Knee - bilateral X-ray 4 views standing
C2826012|T102|strict|38852-0|LNC|Knee - left X-ray 4 views standing|Knee - left X-ray 4 views standing
C2826012|T102|strict|37763-0|LNC|Knee - right X-ray 4 views standing|Knee - right X-ray 4 views standing
C2826012|T102|strict|36675-7|LNC|Facial bones X-ray 5 views|Facial bones X-ray 5 views
C2826012|T102|strict|36676-5|LNC|Knee - left X-ray 5 views|Knee - left X-ray 5 views
C2826012|T102|strict|37744-0|LNC|Knee - right X-ray 5 views|Knee - right X-ray 5 views
C2826012|T102|strict|36890-2|LNC|Mastoid X-ray 5 views|Mastoid X-ray 5 views
C2826012|T102|strict|37351-4|LNC|Pelvis and Spine Lumbar X-ray 5 views|Pelvis and Spine Lumbar X-ray 5 views
C2826012|T102|strict|30750-4|LNC|Shoulder X-ray 5 views|Shoulder X-ray 5 views
C2826012|T102|strict|36677-3|LNC|Shoulder - left X-ray 5 views|Shoulder - left X-ray 5 views
C2826012|T102|strict|37795-2|LNC|Shoulder - right X-ray 5 views|Shoulder - right X-ray 5 views
C2826012|T102|strict|37856-2|LNC|Sinuses X-ray 5 views|Sinuses X-ray 5 views
C2826012|T102|strict|24922-7|LNC|Skull X-ray 5 views|Skull X-ray 5 views
C2826012|T102|strict|24939-1|LNC|Spine Cervical X-ray 5 views|Spine Cervical X-ray 5 views
C2826012|T102|strict|30797-5|LNC|Spine Lumbar X-ray 5 views|Spine Lumbar X-ray 5 views
C2826012|T102|strict|37353-0|LNC|Spine Lumbar and Sacroiliac Joint X-ray 5 views|Spine Lumbar and Sacroiliac Joint X-ray 5 views
C2826012|T102|strict|37355-5|LNC|Spine Lumbar and Sacrum X-ray 5 views|Spine Lumbar and Sacrum X-ray 5 views
C2826012|T102|strict|37356-3|LNC|Spine Lumbar and Sacrum and Coccyx X-ray 5 views|Spine Lumbar and Sacrum and Coccyx X-ray 5 views
C2826012|T102|strict|37357-1|LNC|Spine Lumbar and Sacrum and Sacroiliac Joint and Coccyx X-ray 5 views|Spine Lumbar and Sacrum and Sacroiliac Joint and Coccyx X-ray 5 views
C2826012|T102|strict|37350-6|LNC|Temporomandibular joint - bilateral X-ray 5 views|Temporomandibular joint - bilateral X-ray 5 views
C2826012|T102|strict|37072-6|LNC|Wrist - left X-ray 5 views|Wrist - left X-ray 5 views
C2826012|T102|strict|37829-9|LNC|Wrist - right X-ray 5 views|Wrist - right X-ray 5 views
C2826012|T102|strict|39407-2|LNC|Spine Thoracic X-ray 5 views and oblique|Spine Thoracic X-ray 5 views and oblique
C2826012|T102|strict|69081-8|LNC|Spine Cervical X-ray 5 views and Swimmers|Spine Cervical X-ray 5 views and Swimmers
C2826012|T102|strict|37073-4|LNC|Spine Lumbar X-ray 5 views standing|Spine Lumbar X-ray 5 views standing
C2826012|T102|strict|69080-0|LNC|Spine Cervical X-ray 5 views W flexion and W extension|Spine Cervical X-ray 5 views W flexion and W extension
C2826012|T102|strict|39063-3|LNC|Spine Lumbar X-ray 5 views W flexion and W extension|Spine Lumbar X-ray 5 views W flexion and W extension
C2826012|T102|strict|42273-3|LNC|Ankle - bilateral X-ray 6 views|Ankle - bilateral X-ray 6 views
C2826012|T102|strict|36678-1|LNC|Knee - bilateral X-ray 6 views|Knee - bilateral X-ray 6 views
C2826012|T102|strict|36679-9|LNC|Shoulder - left X-ray 6 views|Shoulder - left X-ray 6 views
C2826012|T102|strict|37796-0|LNC|Shoulder - right X-ray 6 views|Shoulder - right X-ray 6 views
C2826012|T102|strict|42691-6|LNC|Spine Cervical X-ray 6 views|Spine Cervical X-ray 6 views
C2826012|T102|strict|38156-6|LNC|Wrist X-ray 6 views|Wrist X-ray 6 views
C2826012|T102|strict|37074-2|LNC|Wrist - left X-ray 6 views|Wrist - left X-ray 6 views
C2826012|T102|strict|37830-7|LNC|Wrist - right X-ray 6 views|Wrist - right X-ray 6 views
C2826012|T102|strict|36680-7|LNC|Spine Cervical X-ray 7 views|Spine Cervical X-ray 7 views
C2826012|T102|strict|36681-5|LNC|Spine Lumbar X-ray 7 views|Spine Lumbar X-ray 7 views
C2826012|T102|strict|36682-3|LNC|Knee - bilateral X-ray 8 views|Knee - bilateral X-ray 8 views
C2826012|T102|strict|36683-1|LNC|Wrist - left X-ray 8 views|Wrist - left X-ray 8 views
C2826012|T102|strict|37831-5|LNC|Wrist - right X-ray 8 views|Wrist - right X-ray 8 views
C2826012|T102|strict|42412-7|LNC|Shoulder - left X-ray 90 degree abduction|Shoulder - left X-ray 90 degree abduction
C2826012|T102|strict|39064-1|LNC|Ribs X-ray anterior and lateral|Ribs X-ray anterior and lateral
C2826012|T102|strict|69070-1|LNC|Ribs - bilateral X-ray anterior and lateral|Ribs - bilateral X-ray anterior and lateral
C2826012|T102|strict|38856-1|LNC|Ribs - left X-ray anterior and lateral|Ribs - left X-ray anterior and lateral
C2826012|T102|strict|37782-0|LNC|Ribs - right X-ray anterior and lateral|Ribs - right X-ray anterior and lateral
C2826012|T102|strict|24796-5|LNC|Abdomen X-ray AP and AP left lateral-decubitus|Abdomen X-ray AP and AP left lateral-decubitus
C2826012|T102|strict|24792-4|LNC|Abdomen X-ray AP and AP left lateral-decubitus portable|Abdomen X-ray AP and AP left lateral-decubitus portable
C2826012|T102|strict|24653-8|LNC|Chest X-ray AP and AP right lateral-decubitus|Chest X-ray AP and AP right lateral-decubitus
C2826012|T102|strict|24654-6|LNC|Chest X-ray AP and AP right lateral-decubitus portable|Chest X-ray AP and AP right lateral-decubitus portable
C2826012|T102|strict|37080-9|LNC|Shoulder - bilateral X-ray AP and axillary|Shoulder - bilateral X-ray AP and axillary
C2826012|T102|strict|37081-7|LNC|Shoulder - bilateral X-ray AP and axillary and outlet|Shoulder - bilateral X-ray AP and axillary and outlet
C2826012|T102|strict|37082-5|LNC|Shoulder - left X-ray AP and axillary and outlet|Shoulder - left X-ray AP and axillary and outlet
C2826012|T102|strict|38781-1|LNC|Shoulder - right X-ray AP and axillary and outlet|Shoulder - right X-ray AP and axillary and outlet
C2826012|T102|strict|39339-7|LNC|Shoulder - bilateral X-ray AP and axillary and outlet and 30 degree caudal angle|Shoulder - bilateral X-ray AP and axillary and outlet and 30 degree caudal angle
C2826012|T102|strict|37083-3|LNC|Shoulder - left X-ray AP and axillary and outlet and Zanca|Shoulder - left X-ray AP and axillary and outlet and Zanca
C2826012|T102|strict|38782-9|LNC|Shoulder - right X-ray AP and axillary and outlet and Zanca|Shoulder - right X-ray AP and axillary and outlet and Zanca
C2826012|T102|strict|37126-0|LNC|Shoulder - bilateral X-ray AP and axillary and Y|Shoulder - bilateral X-ray AP and axillary and Y
C2826012|T102|strict|37084-1|LNC|Shoulder - left X-ray AP and axillary and Y|Shoulder - left X-ray AP and axillary and Y
C2826012|T102|strict|38783-7|LNC|Shoulder - right X-ray AP and axillary and Y|Shoulder - right X-ray AP and axillary and Y
C2826012|T102|strict|39512-9|LNC|Hip - right X-ray AP and Danelius Miller|Hip - right X-ray AP and Danelius Miller
C2826012|T102|strict|39401-5|LNC|Shoulder X-ray AP and Grashey and axillary|Shoulder X-ray AP and Grashey and axillary
C2826012|T102|strict|69153-5|LNC|Shoulder - left X-ray AP and Grashey and axillary|Shoulder - left X-ray AP and Grashey and axillary
C2826012|T102|strict|69262-4|LNC|Shoulder - right X-ray AP and Grashey and axillary|Shoulder - right X-ray AP and Grashey and axillary
C2826012|T102|strict|37618-6|LNC|Pelvis X-ray AP and inlet|Pelvis X-ray AP and inlet
C2826012|T102|strict|37623-6|LNC|Pelvis X-ray AP and inlet and outlet|Pelvis X-ray AP and inlet and outlet
C2826012|T102|strict|39065-8|LNC|Pelvis X-ray AP and inlet and outlet and oblique|Pelvis X-ray AP and inlet and outlet and oblique
C2826012|T102|strict|37619-4|LNC|Pelvis X-ray AP and Judet|Pelvis X-ray AP and Judet
C2826012|T102|strict|24794-0|LNC|Abdomen X-ray AP and lateral|Abdomen X-ray AP and lateral
C2826012|T102|strict|30779-3|LNC|Ankle X-ray AP and lateral|Ankle X-ray AP and lateral
C2826012|T102|strict|36684-9|LNC|Ankle - bilateral X-ray AP and lateral|Ankle - bilateral X-ray AP and lateral
C2826012|T102|strict|36685-6|LNC|Ankle - left X-ray AP and lateral|Ankle - left X-ray AP and lateral
C2826012|T102|strict|37667-3|LNC|Ankle - right X-ray AP and lateral|Ankle - right X-ray AP and lateral
C2826012|T102|strict|36686-4|LNC|Calcaneus - bilateral X-ray AP and lateral|Calcaneus - bilateral X-ray AP and lateral
C2826012|T102|strict|36701-1|LNC|Calcaneus - left X-ray AP and lateral|Calcaneus - left X-ray AP and lateral
C2826012|T102|strict|37719-2|LNC|Calcaneus - right X-ray AP and lateral|Calcaneus - right X-ray AP and lateral
C2826012|T102|strict|36687-2|LNC|Chest X-ray AP and lateral|Chest X-ray AP and lateral
C2826012|T102|strict|39066-6|LNC|Chest Fluoroscopy AP and lateral|Chest Fluoroscopy AP and lateral
C2826012|T102|strict|36688-0|LNC|Coccyx X-ray AP and lateral|Coccyx X-ray AP and lateral
C2826012|T102|strict|36689-8|LNC|Elbow X-ray AP and lateral|Elbow X-ray AP and lateral
C2826012|T102|strict|36690-6|LNC|Elbow - bilateral X-ray AP and lateral|Elbow - bilateral X-ray AP and lateral
C2826012|T102|strict|36691-4|LNC|Elbow - left X-ray AP and lateral|Elbow - left X-ray AP and lateral
C2826012|T102|strict|37684-8|LNC|Elbow - right X-ray AP and lateral|Elbow - right X-ray AP and lateral
C2826012|T102|strict|36693-0|LNC|Femur X-ray AP and lateral|Femur X-ray AP and lateral
C2826012|T102|strict|36694-8|LNC|Femur - bilateral X-ray AP and lateral|Femur - bilateral X-ray AP and lateral
C2826012|T102|strict|36695-5|LNC|Femur - left X-ray AP and lateral|Femur - left X-ray AP and lateral
C2826012|T102|strict|37692-1|LNC|Femur - right X-ray AP and lateral|Femur - right X-ray AP and lateral
C2826012|T102|strict|39069-0|LNC|Foot X-ray AP and lateral|Foot X-ray AP and lateral
C2826012|T102|strict|36696-3|LNC|Foot - bilateral X-ray AP and lateral|Foot - bilateral X-ray AP and lateral
C2826012|T102|strict|36697-1|LNC|Foot - left X-ray AP and lateral|Foot - left X-ray AP and lateral
C2826012|T102|strict|37701-0|LNC|Foot - right X-ray AP and lateral|Foot - right X-ray AP and lateral
C2826012|T102|strict|42409-3|LNC|Foot sesamoid bones X-ray AP and lateral|Foot sesamoid bones X-ray AP and lateral
C2826012|T102|strict|69130-3|LNC|Hand X-ray AP and lateral|Hand X-ray AP and lateral
C2826012|T102|strict|48474-1|LNC|Hand - bilateral X-ray AP and lateral|Hand - bilateral X-ray AP and lateral
C2826012|T102|strict|38847-0|LNC|Hand - left X-ray AP and lateral|Hand - left X-ray AP and lateral
C2826012|T102|strict|37710-1|LNC|Hand - right X-ray AP and lateral|Hand - right X-ray AP and lateral
C2826012|T102|strict|36702-9|LNC|Hip X-ray AP and lateral|Hip X-ray AP and lateral
C2826012|T102|strict|36703-7|LNC|Hip - bilateral X-ray AP and lateral|Hip - bilateral X-ray AP and lateral
C2826012|T102|strict|36704-5|LNC|Hip - left X-ray AP and lateral|Hip - left X-ray AP and lateral
C2826012|T102|strict|37725-9|LNC|Hip - right X-ray AP and lateral|Hip - right X-ray AP and lateral
C2826012|T102|strict|36706-0|LNC|Humerus X-ray AP and lateral|Humerus X-ray AP and lateral
C2826012|T102|strict|36707-8|LNC|Humerus - bilateral X-ray AP and lateral|Humerus - bilateral X-ray AP and lateral
C2826012|T102|strict|36708-6|LNC|Humerus - left X-ray AP and lateral|Humerus - left X-ray AP and lateral
C2826012|T102|strict|37736-6|LNC|Humerus - right X-ray AP and lateral|Humerus - right X-ray AP and lateral
C2826012|T102|strict|36709-4|LNC|Knee X-ray AP and lateral|Knee X-ray AP and lateral
C2826012|T102|strict|36590-8|LNC|Knee - bilateral X-ray AP and lateral|Knee - bilateral X-ray AP and lateral
C2826012|T102|strict|36710-2|LNC|Knee - left X-ray AP and lateral|Knee - left X-ray AP and lateral
C2826012|T102|strict|37745-7|LNC|Knee - right X-ray AP and lateral|Knee - right X-ray AP and lateral
C2826012|T102|strict|36692-2|LNC|Lower extremity X-ray AP and lateral|Lower extremity X-ray AP and lateral
C2826012|T102|strict|69258-2|LNC|Lower extremity - right X-ray AP and lateral|Lower extremity - right X-ray AP and lateral
C2826012|T102|strict|36711-0|LNC|Mandible X-ray AP and lateral|Mandible X-ray AP and lateral
C2826012|T102|strict|42438-2|LNC|Neck X-ray AP and lateral|Neck X-ray AP and lateral
C2826012|T102|strict|36712-8|LNC|Patella - bilateral X-ray AP and lateral|Patella - bilateral X-ray AP and lateral
C2826012|T102|strict|36713-6|LNC|Patella - left X-ray AP and lateral|Patella - left X-ray AP and lateral
C2826012|T102|strict|37776-2|LNC|Patella - right X-ray AP and lateral|Patella - right X-ray AP and lateral
C2826012|T102|strict|37620-2|LNC|Pelvis X-ray AP and lateral|Pelvis X-ray AP and lateral
C2826012|T102|strict|36705-2|LNC|Pelvis and Hip X-ray AP and lateral|Pelvis and Hip X-ray AP and lateral
C2826012|T102|strict|36699-7|LNC|Radius - bilateral and Ulna - bilateral X-ray AP and lateral|Radius - bilateral and Ulna - bilateral X-ray AP and lateral
C2826012|T102|strict|36700-3|LNC|Radius - left and Ulna.left X-ray AP and lateral|Radius - left and Ulna.left X-ray AP and lateral
C2826012|T102|strict|37708-5|LNC|Radius - right and Ulna - right X-ray AP and lateral|Radius - right and Ulna - right X-ray AP and lateral
C2826012|T102|strict|36698-9|LNC|Radius and Ulna X-ray AP and lateral|Radius and Ulna X-ray AP and lateral
C2826012|T102|strict|37652-5|LNC|Sacrum X-ray AP and lateral|Sacrum X-ray AP and lateral
C2826012|T102|strict|36714-4|LNC|Scapula - bilateral X-ray AP and lateral|Scapula - bilateral X-ray AP and lateral
C2826012|T102|strict|36715-1|LNC|Scapula - left X-ray AP and lateral|Scapula - left X-ray AP and lateral
C2826012|T102|strict|37788-7|LNC|Scapula - right X-ray AP and lateral|Scapula - right X-ray AP and lateral
C2826012|T102|strict|37841-4|LNC|Shoulder X-ray AP and lateral|Shoulder X-ray AP and lateral
C2826012|T102|strict|36716-9|LNC|Shoulder - bilateral X-ray AP and lateral|Shoulder - bilateral X-ray AP and lateral
C2826012|T102|strict|24919-3|LNC|Skull X-ray AP and lateral|Skull X-ray AP and lateral
C2826012|T102|strict|24928-4|LNC|Spine X-ray AP and lateral|Spine X-ray AP and lateral
C2826012|T102|strict|24942-5|LNC|Spine Cervical X-ray AP and lateral|Spine Cervical X-ray AP and lateral
C2826012|T102|strict|37361-3|LNC|Spine Cervical and Spine Thoracic X-ray AP and lateral|Spine Cervical and Spine Thoracic X-ray AP and lateral
C2826012|T102|strict|39067-4|LNC|Spine Cervical and Thoracic and Lumbar X-ray AP and lateral|Spine Cervical and Thoracic and Lumbar X-ray AP and lateral
C2826012|T102|strict|43785-5|LNC|Spine Cervicothoracic Junction X-ray AP and lateral|Spine Cervicothoracic Junction X-ray AP and lateral
C2826012|T102|strict|24970-6|LNC|Spine Lumbar X-ray AP and lateral|Spine Lumbar X-ray AP and lateral
C2826012|T102|strict|30753-8|LNC|Spine Thoracic X-ray AP and lateral|Spine Thoracic X-ray AP and lateral
C2826012|T102|strict|38123-6|LNC|Spine Thoracic and Lumbar X-ray AP and lateral|Spine Thoracic and Lumbar X-ray AP and lateral
C2826012|T102|strict|37974-3|LNC|Spine Thoracolumbar Junction X-ray AP and lateral|Spine Thoracolumbar Junction X-ray AP and lateral
C2826012|T102|strict|37889-3|LNC|Thumb X-ray AP and lateral|Thumb X-ray AP and lateral
C2826012|T102|strict|36717-7|LNC|Tibia - bilateral and Fibula - bilateral X-ray AP and lateral|Tibia - bilateral and Fibula - bilateral X-ray AP and lateral
C2826012|T102|strict|36718-5|LNC|Tibia - left and Fibula - left X-ray AP and lateral|Tibia - left and Fibula - left X-ray AP and lateral
C2826012|T102|strict|37816-6|LNC|Tibia - right and Fibula - right X-ray AP and lateral|Tibia - right and Fibula - right X-ray AP and lateral
C2826012|T102|strict|37896-8|LNC|Tibia and Fibula X-ray AP and lateral|Tibia and Fibula X-ray AP and lateral
C2826012|T102|strict|36719-3|LNC|Toes - left X-ray AP and lateral|Toes - left X-ray AP and lateral
C2826012|T102|strict|37822-4|LNC|Toes - right X-ray AP and lateral|Toes - right X-ray AP and lateral
C2826012|T102|strict|30793-4|LNC|Wrist X-ray AP and lateral|Wrist X-ray AP and lateral
C2826012|T102|strict|38860-3|LNC|Wrist - left X-ray AP and lateral|Wrist - left X-ray AP and lateral
C2826012|T102|strict|37832-3|LNC|Wrist - right X-ray AP and lateral|Wrist - right X-ray AP and lateral
C2826012|T102|strict|37839-8|LNC|Shoulder X-ray AP and lateral and axillary|Shoulder X-ray AP and lateral and axillary
C2826012|T102|strict|39070-8|LNC|Chest X-ray AP and lateral and lordotic|Chest X-ray AP and lateral and lordotic
C2826012|T102|strict|42404-4|LNC|Hip - left X-ray AP and lateral and measurement|Hip - left X-ray AP and lateral and measurement
C2826012|T102|strict|39071-6|LNC|Knee X-ray AP and lateral and Merchants|Knee X-ray AP and lateral and Merchants
C2826012|T102|strict|37095-7|LNC|Ankle X-ray AP and lateral and Mortise|Ankle X-ray AP and lateral and Mortise
C2826012|T102|strict|37096-5|LNC|Ankle - bilateral X-ray AP and lateral and Mortise|Ankle - bilateral X-ray AP and lateral and Mortise
C2826012|T102|strict|37097-3|LNC|Ankle - left X-ray AP and lateral and Mortise|Ankle - left X-ray AP and lateral and Mortise
C2826012|T102|strict|37666-5|LNC|Ankle - right X-ray AP and lateral and Mortise|Ankle - right X-ray AP and lateral and Mortise
C2826012|T102|strict|39072-4|LNC|Ankle X-ray AP and lateral and oblique|Ankle X-ray AP and lateral and oblique
C2826012|T102|strict|36720-1|LNC|Ankle - bilateral X-ray AP and lateral and oblique|Ankle - bilateral X-ray AP and lateral and oblique
C2826012|T102|strict|36721-9|LNC|Ankle - left X-ray AP and lateral and oblique|Ankle - left X-ray AP and lateral and oblique
C2826012|T102|strict|37668-1|LNC|Ankle - right X-ray AP and lateral and oblique|Ankle - right X-ray AP and lateral and oblique
C2826012|T102|strict|36731-8|LNC|Calcaneus X-ray AP and lateral and oblique|Calcaneus X-ray AP and lateral and oblique
C2826012|T102|strict|36722-7|LNC|Elbow X-ray AP and lateral and oblique|Elbow X-ray AP and lateral and oblique
C2826012|T102|strict|36723-5|LNC|Elbow - bilateral X-ray AP and lateral and oblique|Elbow - bilateral X-ray AP and lateral and oblique
C2826012|T102|strict|36724-3|LNC|Elbow - left X-ray AP and lateral and oblique|Elbow - left X-ray AP and lateral and oblique
C2826012|T102|strict|37685-5|LNC|Elbow - right X-ray AP and lateral and oblique|Elbow - right X-ray AP and lateral and oblique
C2826012|T102|strict|36725-0|LNC|Finger X-ray AP and lateral and oblique|Finger X-ray AP and lateral and oblique
C2826012|T102|strict|36726-8|LNC|Finger - bilateral X-ray AP and lateral and oblique|Finger - bilateral X-ray AP and lateral and oblique
C2826012|T102|strict|36727-6|LNC|Finger - left X-ray AP and lateral and oblique|Finger - left X-ray AP and lateral and oblique
C2826012|T102|strict|37696-2|LNC|Finger - right X-ray AP and lateral and oblique|Finger - right X-ray AP and lateral and oblique
C2826012|T102|strict|36728-4|LNC|Foot X-ray AP and lateral and oblique|Foot X-ray AP and lateral and oblique
C2826012|T102|strict|36729-2|LNC|Foot - bilateral X-ray AP and lateral and oblique|Foot - bilateral X-ray AP and lateral and oblique
C2826012|T102|strict|36730-0|LNC|Foot - left X-ray AP and lateral and oblique|Foot - left X-ray AP and lateral and oblique
C2826012|T102|strict|37702-8|LNC|Foot - right X-ray AP and lateral and oblique|Foot - right X-ray AP and lateral and oblique
C2826012|T102|strict|69057-8|LNC|Hand - bilateral X-ray AP and lateral and oblique|Hand - bilateral X-ray AP and lateral and oblique
C2826012|T102|strict|38848-8|LNC|Hand - left X-ray AP and lateral and oblique|Hand - left X-ray AP and lateral and oblique
C2826012|T102|strict|37711-9|LNC|Hand - right X-ray AP and lateral and oblique|Hand - right X-ray AP and lateral and oblique
C2826012|T102|strict|36732-6|LNC|Knee - bilateral X-ray AP and lateral and oblique|Knee - bilateral X-ray AP and lateral and oblique
C2826012|T102|strict|36733-4|LNC|Knee - left X-ray AP and lateral and oblique|Knee - left X-ray AP and lateral and oblique
C2826012|T102|strict|37748-1|LNC|Knee - right X-ray AP and lateral and oblique|Knee - right X-ray AP and lateral and oblique
C2826012|T102|strict|37624-4|LNC|Pelvis X-ray AP and lateral and oblique|Pelvis X-ray AP and lateral and oblique
C2826012|T102|strict|36734-2|LNC|Spine Cervical X-ray AP and lateral and oblique|Spine Cervical X-ray AP and lateral and oblique
C2826012|T102|strict|36735-9|LNC|Spine Lumbar X-ray AP and lateral and oblique|Spine Lumbar X-ray AP and lateral and oblique
C2826012|T102|strict|37908-1|LNC|Spine Thoracic X-ray AP and lateral and oblique|Spine Thoracic X-ray AP and lateral and oblique
C2826012|T102|strict|36736-7|LNC|Thumb - left X-ray AP and lateral and oblique|Thumb - left X-ray AP and lateral and oblique
C2826012|T102|strict|37813-3|LNC|Thumb - right X-ray AP and lateral and oblique|Thumb - right X-ray AP and lateral and oblique
C2826012|T102|strict|37927-1|LNC|Wrist X-ray AP and lateral and oblique|Wrist X-ray AP and lateral and oblique
C2826012|T102|strict|37099-9|LNC|Spine Cervical X-ray AP and lateral and oblique and odontoid|Spine Cervical X-ray AP and lateral and oblique and odontoid
C2826012|T102|strict|38083-2|LNC|Spine Cervical X-ray AP and lateral and oblique and odontoid and swimmer|Spine Cervical X-ray AP and lateral and oblique and odontoid and swimmer
C2826012|T102|strict|37101-3|LNC|Spine Lumbar X-ray AP and lateral and oblique and spot|Spine Lumbar X-ray AP and lateral and oblique and spot
C2826012|T102|strict|42410-1|LNC|Spine Lumbar X-ray AP and lateral and oblique and spot standing|Spine Lumbar X-ray AP and lateral and oblique and spot standing
C2826012|T102|strict|37102-1|LNC|Knee - bilateral X-ray AP and lateral and oblique and Sunrise|Knee - bilateral X-ray AP and lateral and oblique and Sunrise
C2826012|T102|strict|37118-7|LNC|Knee - bilateral X-ray AP and lateral and oblique and Sunrise and tunnel|Knee - bilateral X-ray AP and lateral and oblique and Sunrise and tunnel
C2826012|T102|strict|37115-3|LNC|Knee X-ray AP and lateral and oblique and tunnel|Knee X-ray AP and lateral and oblique and tunnel
C2826012|T102|strict|69137-8|LNC|Ankle - left X-ray AP and lateral and oblique standing|Ankle - left X-ray AP and lateral and oblique standing
C2826012|T102|strict|39371-0|LNC|Ankle - right X-ray AP and lateral and oblique standing|Ankle - right X-ray AP and lateral and oblique standing
C2826012|T102|strict|39334-8|LNC|Foot - left X-ray AP and lateral and oblique standing|Foot - left X-ray AP and lateral and oblique standing
C2826012|T102|strict|39375-1|LNC|Foot - right X-ray AP and lateral and oblique standing|Foot - right X-ray AP and lateral and oblique standing
C2826012|T102|strict|42417-6|LNC|Ankle - bilateral X-ray AP and lateral and oblique W manual stress|Ankle - bilateral X-ray AP and lateral and oblique W manual stress
C2826012|T102|strict|42418-4|LNC|Ankle - left X-ray AP and lateral and oblique W manual stress|Ankle - left X-ray AP and lateral and oblique W manual stress
C2826012|T102|strict|39369-4|LNC|Ankle - right X-ray AP and lateral and oblique W manual stress|Ankle - right X-ray AP and lateral and oblique W manual stress
C2826012|T102|strict|37103-9|LNC|Spine Cervical X-ray AP and lateral and odontoid|Spine Cervical X-ray AP and lateral and odontoid
C2826012|T102|strict|37079-1|LNC|Spine Cervical X-ray AP and lateral and odontoid portable|Spine Cervical X-ray AP and lateral and odontoid portable
C2826012|T102|strict|39074-0|LNC|Chest X-ray AP and lateral and right oblique and left oblique|Chest X-ray AP and lateral and right oblique and left oblique
C2826012|T102|strict|39073-2|LNC|Knee X-ray AP and lateral and right oblique and left oblique|Knee X-ray AP and lateral and right oblique and left oblique
C2826012|T102|strict|69147-7|LNC|Knee - left X-ray AP and lateral and right oblique and left oblique|Knee - left X-ray AP and lateral and right oblique and left oblique
C2826012|T102|strict|39388-4|LNC|Knee - right X-ray AP and lateral and right oblique and left oblique|Knee - right X-ray AP and lateral and right oblique and left oblique
C2826012|T102|strict|37105-4|LNC|Spine Lumbar X-ray AP and lateral and spot|Spine Lumbar X-ray AP and lateral and spot
C2826012|T102|strict|37106-2|LNC|Knee X-ray AP and lateral and Sunrise|Knee X-ray AP and lateral and Sunrise
C2826012|T102|strict|37107-0|LNC|Knee - bilateral X-ray AP and lateral and Sunrise|Knee - bilateral X-ray AP and lateral and Sunrise
C2826012|T102|strict|37108-8|LNC|Knee - left X-ray AP and lateral and Sunrise|Knee - left X-ray AP and lateral and Sunrise
C2826012|T102|strict|37749-9|LNC|Knee - right X-ray AP and lateral and Sunrise|Knee - right X-ray AP and lateral and Sunrise
C2826012|T102|strict|37109-6|LNC|Patella - bilateral X-ray AP and lateral and Sunrise|Patella - bilateral X-ray AP and lateral and Sunrise
C2826012|T102|strict|37110-4|LNC|Patella - left X-ray AP and lateral and Sunrise|Patella - left X-ray AP and lateral and Sunrise
C2826012|T102|strict|38786-0|LNC|Patella - right X-ray AP and lateral and Sunrise|Patella - right X-ray AP and lateral and Sunrise
C2826012|T102|strict|37111-2|LNC|Knee X-ray AP and lateral and Sunrise and tunnel|Knee X-ray AP and lateral and Sunrise and tunnel
C2826012|T102|strict|37116-1|LNC|Knee - bilateral X-ray AP and lateral and Sunrise and tunnel|Knee - bilateral X-ray AP and lateral and Sunrise and tunnel
C2826012|T102|strict|37117-9|LNC|Knee - left X-ray AP and lateral and Sunrise and tunnel|Knee - left X-ray AP and lateral and Sunrise and tunnel
C2826012|T102|strict|37740-8|LNC|Knee - right X-ray AP and lateral and Sunrise and tunnel|Knee - right X-ray AP and lateral and Sunrise and tunnel
C2826012|T102|strict|38009-7|LNC|Spine Thoracic X-ray AP and lateral and Swimmers|Spine Thoracic X-ray AP and lateral and Swimmers
C2826012|T102|strict|37112-0|LNC|Knee X-ray AP and lateral and tunnel|Knee X-ray AP and lateral and tunnel
C2826012|T102|strict|37113-8|LNC|Knee - bilateral X-ray AP and lateral and tunnel|Knee - bilateral X-ray AP and lateral and tunnel
C2826012|T102|strict|37114-6|LNC|Knee - left X-ray AP and lateral and tunnel|Knee - left X-ray AP and lateral and tunnel
C2826012|T102|strict|37747-3|LNC|Knee - right X-ray AP and lateral and tunnel|Knee - right X-ray AP and lateral and tunnel
C2826012|T102|strict|69065-1|LNC|Abdomen X-ray AP and lateral crosstable|Abdomen X-ray AP and lateral crosstable
C2826012|T102|strict|37086-6|LNC|Hip X-ray AP and lateral crosstable|Hip X-ray AP and lateral crosstable
C2826012|T102|strict|37087-4|LNC|Hip - left X-ray AP and lateral crosstable|Hip - left X-ray AP and lateral crosstable
C2826012|T102|strict|37723-4|LNC|Hip - right X-ray AP and lateral crosstable|Hip - right X-ray AP and lateral crosstable
C2826012|T102|strict|37090-8|LNC|Knee X-ray AP and lateral crosstable|Knee X-ray AP and lateral crosstable
C2826012|T102|strict|69146-9|LNC|Knee - left X-ray AP and lateral crosstable|Knee - left X-ray AP and lateral crosstable
C2826012|T102|strict|37089-0|LNC|Pelvis and Hip X-ray AP and lateral crosstable|Pelvis and Hip X-ray AP and lateral crosstable
C2826012|T102|strict|37088-2|LNC|Pelvis and Hip - left X-ray AP and lateral crosstable|Pelvis and Hip - left X-ray AP and lateral crosstable
C2826012|T102|strict|38784-5|LNC|Pelvis and Hip - right X-ray AP and lateral crosstable|Pelvis and Hip - right X-ray AP and lateral crosstable
C2826012|T102|strict|30763-7|LNC|Abdomen X-ray AP and lateral crosstable portable|Abdomen X-ray AP and lateral crosstable portable
C2826012|T102|strict|37077-5|LNC|Hip X-ray AP and lateral crosstable portable|Hip X-ray AP and lateral crosstable portable
C2826012|T102|strict|37091-6|LNC|Hip X-ray AP and lateral frog|Hip X-ray AP and lateral frog
C2826012|T102|strict|37092-4|LNC|Hip - bilateral X-ray AP and lateral frog|Hip - bilateral X-ray AP and lateral frog
C2826012|T102|strict|37093-2|LNC|Hip - left X-ray AP and lateral frog|Hip - left X-ray AP and lateral frog
C2826012|T102|strict|37724-2|LNC|Hip - right X-ray AP and lateral frog|Hip - right X-ray AP and lateral frog
C2826012|T102|strict|30770-2|LNC|Pelvis and Hip X-ray AP and lateral frog|Pelvis and Hip X-ray AP and lateral frog
C2826012|T102|strict|42167-7|LNC|Pelvis and Hip - bilateral X-ray AP and lateral frog|Pelvis and Hip - bilateral X-ray AP and lateral frog
C2826012|T102|strict|37094-0|LNC|Pelvis and Hip - left X-ray AP and lateral frog|Pelvis and Hip - left X-ray AP and lateral frog
C2826012|T102|strict|38785-2|LNC|Pelvis and Hip - right X-ray AP and lateral frog|Pelvis and Hip - right X-ray AP and lateral frog
C2826012|T102|strict|41776-6|LNC|Pelvis and Hip - right X-ray AP and lateral frog portable|Pelvis and Hip - right X-ray AP and lateral frog portable
C2826012|T102|strict|24793-2|LNC|Abdomen X-ray AP and lateral portable|Abdomen X-ray AP and lateral portable
C2826012|T102|strict|44185-7|LNC|Femur X-ray AP and lateral portable|Femur X-ray AP and lateral portable
C2826012|T102|strict|44186-5|LNC|Foot X-ray AP and lateral portable|Foot X-ray AP and lateral portable
C2826012|T102|strict|41817-8|LNC|Hip - left X-ray AP and lateral portable|Hip - left X-ray AP and lateral portable
C2826012|T102|strict|41777-4|LNC|Hip - right X-ray AP and lateral portable|Hip - right X-ray AP and lateral portable
C2826012|T102|strict|30726-4|LNC|Spine Cervical X-ray AP and lateral portable|Spine Cervical X-ray AP and lateral portable
C2826012|T102|strict|37078-3|LNC|Spine Lumbar X-ray AP and lateral portable|Spine Lumbar X-ray AP and lateral portable
C2826012|T102|strict|30754-6|LNC|Spine Thoracic X-ray AP and lateral portable|Spine Thoracic X-ray AP and lateral portable
C2826012|T102|strict|39330-6|LNC|Ankle - bilateral X-ray AP and lateral standing|Ankle - bilateral X-ray AP and lateral standing
C2826012|T102|strict|42380-6|LNC|Ankle - left X-ray AP and lateral standing|Ankle - left X-ray AP and lateral standing
C2826012|T102|strict|39368-6|LNC|Ankle - right X-ray AP and lateral standing|Ankle - right X-ray AP and lateral standing
C2826012|T102|strict|39068-2|LNC|Foot X-ray AP and lateral standing|Foot X-ray AP and lateral standing
C2826012|T102|strict|39331-4|LNC|Foot - bilateral X-ray AP and lateral standing|Foot - bilateral X-ray AP and lateral standing
C2826012|T102|strict|39332-2|LNC|Foot - left X-ray AP and lateral standing|Foot - left X-ray AP and lateral standing
C2826012|T102|strict|39374-4|LNC|Foot - right X-ray AP and lateral standing|Foot - right X-ray AP and lateral standing
C2826012|T102|strict|24805-4|LNC|Knee X-ray AP and lateral standing|Knee X-ray AP and lateral standing
C2826012|T102|strict|26364-0|LNC|Knee - bilateral X-ray AP and lateral standing|Knee - bilateral X-ray AP and lateral standing
C2826012|T102|strict|26365-7|LNC|Knee - left X-ray AP and lateral standing|Knee - left X-ray AP and lateral standing
C2826012|T102|strict|26366-5|LNC|Knee - right X-ray AP and lateral standing|Knee - right X-ray AP and lateral standing
C2826012|T102|strict|39333-0|LNC|Spine Lumbar X-ray AP and lateral standing|Spine Lumbar X-ray AP and lateral standing
C2826012|T102|strict|38084-0|LNC|Abdomen X-ray AP and left posterior oblique|Abdomen X-ray AP and left posterior oblique
C2826012|T102|strict|37119-5|LNC|Abdomen X-ray AP and oblique|Abdomen X-ray AP and oblique
C2826012|T102|strict|39076-5|LNC|Foot X-ray AP and oblique|Foot X-ray AP and oblique
C2826012|T102|strict|37621-0|LNC|Pelvis X-ray AP and oblique|Pelvis X-ray AP and oblique
C2826012|T102|strict|37649-1|LNC|Sacroiliac Joint X-ray AP and oblique|Sacroiliac Joint X-ray AP and oblique
C2826012|T102|strict|39075-7|LNC|Toes X-ray AP and oblique|Toes X-ray AP and oblique
C2826012|T102|strict|37098-1|LNC|Spine Cervical X-ray AP and oblique and lateral W flexion and W extension|Spine Cervical X-ray AP and oblique and lateral W flexion and W extension
C2826012|T102|strict|44187-3|LNC|Spine Cervical X-ray AP and oblique and odontoid and lateral portable W flexion and W extension|Spine Cervical X-ray AP and oblique and odontoid and lateral portable W flexion and W extension
C2826012|T102|strict|37100-5|LNC|Spine Cervical X-ray AP and oblique and odontoid and lateral W flexion and W extension|Spine Cervical X-ray AP and oblique and odontoid and lateral W flexion and W extension
C2826012|T102|strict|24797-3|LNC|Abdomen X-ray AP and oblique prone|Abdomen X-ray AP and oblique prone
C2826012|T102|strict|37120-3|LNC|Spine Cervical X-ray AP and odontoid and lateral crosstable|Spine Cervical X-ray AP and odontoid and lateral crosstable
C2826012|T102|strict|37104-7|LNC|Spine Cervical X-ray AP and odontoid and lateral W flexion and W extension|Spine Cervical X-ray AP and odontoid and lateral W flexion and W extension
C2826012|T102|strict|42011-7|LNC|Chest and Abdomen X-ray AP and PA chest|Chest and Abdomen X-ray AP and PA chest
C2826012|T102|strict|24642-1|LNC|Chest X-ray AP and PA upright|Chest X-ray AP and PA upright
C2826012|T102|strict|24808-8|LNC|Knee X-ray AP and PA standing|Knee X-ray AP and PA standing
C2826012|T102|strict|26361-6|LNC|Knee - bilateral X-ray AP and PA standing|Knee - bilateral X-ray AP and PA standing
C2826012|T102|strict|26362-4|LNC|Knee - left X-ray AP and PA standing|Knee - left X-ray AP and PA standing
C2826012|T102|strict|26363-2|LNC|Knee - right X-ray AP and PA standing|Knee - right X-ray AP and PA standing
C2826012|T102|strict|37121-1|LNC|Clavicle - left X-ray AP and Serendipity|Clavicle - left X-ray AP and Serendipity
C2826012|T102|strict|37680-6|LNC|Clavicle - right X-ray AP and Serendipity|Clavicle - right X-ray AP and Serendipity
C2826012|T102|strict|37122-9|LNC|Shoulder - left X-ray AP and Stryker Notch|Shoulder - left X-ray AP and Stryker Notch
C2826012|T102|strict|37797-8|LNC|Shoulder - right X-ray AP and Stryker Notch|Shoulder - right X-ray AP and Stryker Notch
C2826012|T102|strict|37485-0|LNC|Humerus X-ray AP and transthoracic|Humerus X-ray AP and transthoracic
C2826012|T102|strict|39077-3|LNC|Shoulder X-ray AP and transthoracic|Shoulder X-ray AP and transthoracic
C2826012|T102|strict|46349-7|LNC|Shoulder - bilateral X-ray AP and transthoracic|Shoulder - bilateral X-ray AP and transthoracic
C2826012|T102|strict|38082-4|LNC|Shoulder - left X-ray AP and transthoracic|Shoulder - left X-ray AP and transthoracic
C2826012|T102|strict|38822-3|LNC|Shoulder - right X-ray AP and transthoracic|Shoulder - right X-ray AP and transthoracic
C2826012|T102|strict|37123-7|LNC|Shoulder - left X-ray AP and West Point|Shoulder - left X-ray AP and West Point
C2826012|T102|strict|38787-8|LNC|Shoulder - right X-ray AP and West Point|Shoulder - right X-ray AP and West Point
C2826012|T102|strict|36961-1|LNC|Shoulder - left X-ray AP and West Point and outlet|Shoulder - left X-ray AP and West Point and outlet
C2826012|T102|strict|37799-4|LNC|Shoulder - right X-ray AP and West Point and outlet|Shoulder - right X-ray AP and West Point and outlet
C2826012|T102|strict|37124-5|LNC|Scapula - left X-ray AP and Y|Scapula - left X-ray AP and Y
C2826012|T102|strict|37789-5|LNC|Scapula - right X-ray AP and Y|Scapula - right X-ray AP and Y
C2826012|T102|strict|69266-5|LNC|Shoulder X-ray AP and Y|Shoulder X-ray AP and Y
C2826012|T102|strict|37125-2|LNC|Shoulder - left X-ray AP and Y|Shoulder - left X-ray AP and Y
C2826012|T102|strict|38788-6|LNC|Shoulder - right X-ray AP and Y|Shoulder - right X-ray AP and Y
C2826012|T102|strict|24562-1|LNC|Abdomen X-ray AP (left lateral-decubitus and right lateral-decubitus)|Abdomen X-ray AP (left lateral-decubitus and right lateral-decubitus)
C2826012|T102|strict|24650-4|LNC|Chest X-ray AP (right lateral-decubitus and left lateral-decubitus)|Chest X-ray AP (right lateral-decubitus and left lateral-decubitus)
C2826012|T102|strict|24649-6|LNC|Chest X-ray AP (right lateral-decubitus and left lateral-decubitus) portable|Chest X-ray AP (right lateral-decubitus and left lateral-decubitus) portable
C2826012|T102|strict|37085-8|LNC|Abdomen X-ray AP (supine and lateral-decubitus)|Abdomen X-ray AP (supine and lateral-decubitus)
C2826012|T102|strict|37076-7|LNC|Abdomen X-ray AP (supine and lateral-decubitus) portable|Abdomen X-ray AP (supine and lateral-decubitus) portable
C2826012|T102|strict|24798-1|LNC|Abdomen X-ray AP (supine and upright)|Abdomen X-ray AP (supine and upright)
C2826012|T102|strict|43463-9|LNC|Chest and Abdomen X-ray AP (supine and upright) and PA chest|Chest and Abdomen X-ray AP (supine and upright) and PA chest
C2826012|T102|strict|24795-7|LNC|Abdomen X-ray AP (supine and upright) portable|Abdomen X-ray AP (supine and upright) portable
C2826012|T102|strict|42019-0|LNC|Abdomen X-ray AP (upright and left lateral decubitus)|Abdomen X-ray AP (upright and left lateral decubitus)
C2826012|T102|strict|39329-8|LNC|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation)|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation)
C2826012|T102|strict|39328-0|LNC|Shoulder - left X-ray AP (W internal rotation and W external rotation)|Shoulder - left X-ray AP (W internal rotation and W external rotation)
C2826012|T102|strict|39395-9|LNC|Shoulder - right X-ray AP (W internal rotation and W external rotation)|Shoulder - right X-ray AP (W internal rotation and W external rotation)
C2826012|T102|strict|39321-5|LNC|Shoulder X-ray AP (W internal rotation and W external rotation) and axillary|Shoulder X-ray AP (W internal rotation and W external rotation) and axillary
C2826012|T102|strict|39336-3|LNC|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and axillary|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and axillary
C2826012|T102|strict|39335-5|LNC|Shoulder - left X-ray AP (W internal rotation and W external rotation) and axillary|Shoulder - left X-ray AP (W internal rotation and W external rotation) and axillary
C2826012|T102|strict|39337-1|LNC|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and axillary and outlet|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and axillary and outlet
C2826012|T102|strict|39344-7|LNC|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and axillary and Y|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and axillary and Y
C2826012|T102|strict|39338-9|LNC|Shoulder - left X-ray AP (W internal rotation and W external rotation) and axillary and Y|Shoulder - left X-ray AP (W internal rotation and W external rotation) and axillary and Y
C2826012|T102|strict|39397-5|LNC|Shoulder - right X-ray AP (W internal rotation and W external rotation) and West Point|Shoulder - right X-ray AP (W internal rotation and W external rotation) and West Point
C2826012|T102|strict|39343-9|LNC|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and Y|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and Y
C2826012|T102|strict|39348-8|LNC|Shoulder - left X-ray AP (W internal rotation and W external rotation) and Y|Shoulder - left X-ray AP (W internal rotation and W external rotation) and Y
C2826012|T102|strict|39325-6|LNC|Shoulder - left X-ray AP (W internal rotation) and Grashey and axillary and outlet|Shoulder - left X-ray AP (W internal rotation) and Grashey and axillary and outlet
C2826012|T102|strict|39346-2|LNC|Shoulder - bilateral X-ray AP (W internal rotation) and West Point|Shoulder - bilateral X-ray AP (W internal rotation) and West Point
C2826012|T102|strict|39347-0|LNC|Shoulder - left X-ray AP (W internal rotation) and West Point|Shoulder - left X-ray AP (W internal rotation) and West Point
C2826012|T102|strict|39396-7|LNC|Shoulder - right X-ray AP (W internal rotation) and West Point|Shoulder - right X-ray AP (W internal rotation) and West Point
C2826012|T102|strict|24632-2|LNC|Chest X-ray AP portable|Chest X-ray AP portable
C2826012|T102|strict|37075-9|LNC|Hip X-ray AP portable|Hip X-ray AP portable
C2826012|T102|strict|43561-0|LNC|Chest and Abdomen X-ray AP upright and AP chest|Chest and Abdomen X-ray AP upright and AP chest
C2826012|T102|strict|38003-0|LNC|Foot - left X-ray AP standing|Foot - left X-ray AP standing
C2826012|T102|strict|38815-7|LNC|Foot - right X-ray AP standing|Foot - right X-ray AP standing
C2826012|T102|strict|42406-9|LNC|Spine Lumbar X-ray AP W and WO left bending|Spine Lumbar X-ray AP W and WO left bending
C2826012|T102|strict|42407-7|LNC|Spine Lumbar X-ray AP W and WO right bending|Spine Lumbar X-ray AP W and WO right bending
C2826012|T102|strict|42445-7|LNC|Spine Thoracic X-ray AP W left bending and WO bending|Spine Thoracic X-ray AP W left bending and WO bending
C2826012|T102|strict|37484-3|LNC|Knee - left X-ray AP W manual stress|Knee - left X-ray AP W manual stress
C2826012|T102|strict|37746-5|LNC|Knee - right X-ray AP W manual stress|Knee - right X-ray AP W manual stress
C2826012|T102|strict|42403-6|LNC|Spine Lumbar X-ray AP W right bending and W left bending|Spine Lumbar X-ray AP W right bending and W left bending
C2826012|T102|strict|42408-5|LNC|Spine Lumbar X-ray AP W right bending and W left bending and WO bending|Spine Lumbar X-ray AP W right bending and W left bending and WO bending
C2826012|T102|strict|42444-0|LNC|Spine Thoracic X-ray AP W right bending and W left bending and WO bending|Spine Thoracic X-ray AP W right bending and W left bending and WO bending
C2826012|T102|strict|42446-5|LNC|Spine Thoracic X-ray AP W right bending and WO bending|Spine Thoracic X-ray AP W right bending and WO bending
C2826012|T102|strict|39403-1|LNC|Shoulder X-ray axillary and transcapular|Shoulder X-ray axillary and transcapular
C2826012|T102|strict|37127-8|LNC|Shoulder - bilateral X-ray axillary and Y|Shoulder - bilateral X-ray axillary and Y
C2826012|T102|strict|37128-6|LNC|Shoulder - left X-ray axillary and Y|Shoulder - left X-ray axillary and Y
C2826012|T102|strict|37807-5|LNC|Shoulder - right X-ray axillary and Y|Shoulder - right X-ray axillary and Y
C2826012|T102|strict|46386-9|LNC|Teeth X-ray bitewing|Teeth X-ray bitewing
C2826012|T102|strict|39884-2|LNC|Bone Scan blood pool|Bone Scan blood pool
C2826012|T102|strict|39861-0|LNC|Heart Scan blood pool|Heart Scan blood pool
C2826012|T102|strict|42709-6|LNC|Liver Scan blood pool|Liver Scan blood pool
C2826012|T102|strict|39860-2|LNC|Heart Scan blood pool W stress and W radionuclide IV|Heart Scan blood pool W stress and W radionuclide IV
C2826012|T102|strict|26352-5|LNC|Wrist - bilateral and Hand - bilateral X-ray bone age|Wrist - bilateral and Hand - bilateral X-ray bone age
C2826012|T102|strict|26353-3|LNC|Wrist - left and Hand - left X-ray bone age|Wrist - left and Hand - left X-ray bone age
C2826012|T102|strict|26354-1|LNC|Wrist - right and Hand - right X-ray bone age|Wrist - right and Hand - right X-ray bone age
C2826012|T102|strict|24724-7|LNC|Wrist and Hand X-ray bone age|Wrist and Hand X-ray bone age
C2826012|T102|strict|37362-1|LNC|Bones X-ray bone age|Bones X-ray bone age
C2826012|T102|strict|24591-0|LNC|Brain Scan brain death protocol W Tc-99m HMPAO IV|Brain Scan brain death protocol W Tc-99m HMPAO IV
C2826012|T102|strict|37996-6|LNC|Calcaneus X-ray Broden|Calcaneus X-ray Broden
C2826012|T102|strict|37995-8|LNC|Calcaneus - bilateral X-ray Broden|Calcaneus - bilateral X-ray Broden
C2826012|T102|strict|37997-4|LNC|Calcaneus - left X-ray Broden|Calcaneus - left X-ray Broden
C2826012|T102|strict|38814-0|LNC|Calcaneus - right X-ray Broden|Calcaneus - right X-ray Broden
C2826012|T102|strict|37486-8|LNC|Ankle X-ray Broden W manual stress|Ankle X-ray Broden W manual stress
C2826012|T102|strict|37852-1|LNC|Sinuses X-ray Caldwell and Waters|Sinuses X-ray Caldwell and Waters
C2826012|T102|strict|39859-4|LNC|Brain Scan delayed static|Brain Scan delayed static
C2826012|T102|strict|39875-0|LNC|Scan delayed W GA-67 IV|Scan delayed W GA-67 IV
C2826012|T102|strict|39840-4|LNC|Scan delayed W I-131 MIBG IV|Scan delayed W I-131 MIBG IV
C2826012|T102|strict|39842-0|LNC|Scan delayed W In-111 Satumomab IV|Scan delayed W In-111 Satumomab IV
C2826012|T102|strict|39874-3|LNC|Head Cistern Scan delayed W radionuclide IT|Head Cistern Scan delayed W radionuclide IT
C2826012|T102|strict|39819-8|LNC|Bone Scan delayed|Bone Scan delayed
C2826012|T102|strict|39741-4|LNC|Parathyroid Scan delayed|Parathyroid Scan delayed
C2826012|T102|strict|24605-8|LNC|Breast Mammogram diagnostic|Breast Mammogram diagnostic
C2826012|T102|strict|39152-4|LNC|Breast FFD mammogram diagnostic|Breast FFD mammogram diagnostic
C2826012|T102|strict|69158-4|LNC|Breast implant X-ray diagnostic|Breast implant X-ray diagnostic
C2826012|T102|strict|48475-8|LNC|Breast implant - bilateral Mammogram diagnostic|Breast implant - bilateral Mammogram diagnostic
C2826012|T102|strict|69150-1|LNC|Breast implant - left Mammogram diagnostic|Breast implant - left Mammogram diagnostic
C2826012|T102|strict|69259-0|LNC|Breast implant - right Mammogram diagnostic|Breast implant - right Mammogram diagnostic
C2826012|T102|strict|26346-7|LNC|Breast - bilateral Mammogram diagnostic|Breast - bilateral Mammogram diagnostic
C2826012|T102|strict|39154-0|LNC|Breast - bilateral FFD mammogram diagnostic|Breast - bilateral FFD mammogram diagnostic
C2826012|T102|strict|26347-5|LNC|Breast - left Mammogram diagnostic|Breast - left Mammogram diagnostic
C2826012|T102|strict|42169-3|LNC|Breast - left FFD mammogram diagnostic|Breast - left FFD mammogram diagnostic
C2826012|T102|strict|26348-3|LNC|Breast - right Mammogram diagnostic|Breast - right Mammogram diagnostic
C2826012|T102|strict|42168-5|LNC|Breast - right FFD mammogram diagnostic|Breast - right FFD mammogram diagnostic
C2826012|T102|strict|46350-5|LNC|Breast - unilateral Mammogram diagnostic|Breast - unilateral Mammogram diagnostic
C2826012|T102|strict|24604-1|LNC|Breast Mammogram diagnostic limited|Breast Mammogram diagnostic limited
C2826012|T102|strict|26349-1|LNC|Breast - bilateral Mammogram diagnostic limited|Breast - bilateral Mammogram diagnostic limited
C2826012|T102|strict|26350-9|LNC|Breast - left Mammogram diagnostic limited|Breast - left Mammogram diagnostic limited
C2826012|T102|strict|26351-7|LNC|Breast - right Mammogram diagnostic limited|Breast - right Mammogram diagnostic limited
C2826012|T102|strict|46351-3|LNC|Breast implant - bilateral Mammogram displacement|Breast implant - bilateral Mammogram displacement
C2826012|T102|strict|39895-8|LNC|Gallbladder Scan ejection fraction W Tc-99m DISIDA IV|Gallbladder Scan ejection fraction W Tc-99m DISIDA IV
C2826012|T102|strict|39887-5|LNC|Heart Scan first pass and ejection fraction at rest and W radionuclide IV|Heart Scan first pass and ejection fraction at rest and W radionuclide IV
C2826012|T102|strict|39889-1|LNC|Heart Scan first pass and ejection fraction|Heart Scan first pass and ejection fraction
C2826012|T102|strict|39885-9|LNC|Heart Scan first pass and ventricular volume|Heart Scan first pass and ventricular volume
C2826012|T102|strict|39910-5|LNC|Heart Scan first pass and wall motion and ejection fraction|Heart Scan first pass and wall motion and ejection fraction
C2826012|T102|strict|39912-1|LNC|Heart Scan first pass and wall motion and ventricular volume and ejection fraction|Heart Scan first pass and wall motion and ventricular volume and ejection fraction
C2826012|T102|strict|39909-7|LNC|Heart Scan first pass and wall motion and ventricular volume and ejection fraction W stress and W radionuclide IV|Heart Scan first pass and wall motion and ventricular volume and ejection fraction W stress and W radionuclide IV
C2826012|T102|strict|39908-9|LNC|Heart Scan first pass and wall motion and ventricular volume W stress and W radionuclide IV|Heart Scan first pass and wall motion and ventricular volume W stress and W radionuclide IV
C2826012|T102|strict|39886-7|LNC|Heart Scan first pass and wall motion at rest and W radionuclide IV|Heart Scan first pass and wall motion at rest and W radionuclide IV
C2826012|T102|strict|39890-9|LNC|Heart Scan first pass and wall motion|Heart Scan first pass and wall motion
C2826012|T102|strict|39888-3|LNC|Heart Scan first pass and wall motion W stress and W radionuclide IV|Heart Scan first pass and wall motion W stress and W radionuclide IV
C2826012|T102|strict|39867-7|LNC|Heart Scan first pass at rest and W radionuclide IV|Heart Scan first pass at rest and W radionuclide IV
C2826012|T102|strict|39863-6|LNC|Heart Scan first pass at rest and W stress and W radionuclide IV|Heart Scan first pass at rest and W stress and W radionuclide IV
C2826012|T102|strict|39866-9|LNC|Heart Scan first pass at rest and W Tc-99m Sestamibi IV|Heart Scan first pass at rest and W Tc-99m Sestamibi IV
C2826012|T102|strict|39864-4|LNC|Heart Scan first pass|Heart Scan first pass
C2826012|T102|strict|39865-1|LNC|Left ventricle Scan first pass|Left ventricle Scan first pass
C2826012|T102|strict|39869-3|LNC|Heart Scan first pass W stress and W radionuclide IV|Heart Scan first pass W stress and W radionuclide IV
C2826012|T102|strict|39868-5|LNC|Heart Scan first pass W stress and W Tc-99m Sestamibi IV|Heart Scan first pass W stress and W Tc-99m Sestamibi IV
C2826012|T102|strict|39893-3|LNC|Heart Scan flow for shunt detection|Heart Scan flow for shunt detection
C2826012|T102|strict|43644-4|LNC|Brain Scan flow limited|Brain Scan flow limited
C2826012|T102|strict|39858-6|LNC|Bone Scan flow|Bone Scan flow
C2826012|T102|strict|39636-6|LNC|Brain Scan flow|Brain Scan flow
C2826012|T102|strict|39871-9|LNC|Heart Scan flow|Heart Scan flow
C2826012|T102|strict|42261-8|LNC|Kidney - bilateral Scan flow|Kidney - bilateral Scan flow
C2826012|T102|strict|42262-6|LNC|Liver Scan flow|Liver Scan flow
C2826012|T102|strict|43653-5|LNC|Liver and Spleen Scan flow|Liver and Spleen Scan flow
C2826012|T102|strict|39847-9|LNC|Parotid gland Scan flow|Parotid gland Scan flow
C2826012|T102|strict|39899-0|LNC|Salivary gland Scan flow|Salivary gland Scan flow
C2826012|T102|strict|42308-7|LNC|Scrotum and Testicle Scan flow|Scrotum and Testicle Scan flow
C2826012|T102|strict|42263-4|LNC|Spleen Scan flow|Spleen Scan flow
C2826012|T102|strict|39856-0|LNC|Thyroid Scan flow|Thyroid Scan flow
C2826012|T102|strict|43500-8|LNC|Vessel Scan flow|Vessel Scan flow
C2826012|T102|strict|44148-5|LNC|Brain Scan flow W Tc-99m bicisate IV|Brain Scan flow W Tc-99m bicisate IV
C2826012|T102|strict|43642-8|LNC|Brain Scan flow W Tc-99m DTPA IV|Brain Scan flow W Tc-99m DTPA IV
C2826012|T102|strict|43664-2|LNC|Renal vessels Scan flow W Tc-99m DTPA IV|Renal vessels Scan flow W Tc-99m DTPA IV
C2826012|T102|strict|43643-6|LNC|Brain Scan flow W Tc-99m glucoheptonate IV|Brain Scan flow W Tc-99m glucoheptonate IV
C2826012|T102|strict|43666-7|LNC|Kidney - bilateral and Renal vessels Scan flow W Tc-99m glucoheptonate IV|Kidney - bilateral and Renal vessels Scan flow W Tc-99m glucoheptonate IV
C2826012|T102|strict|43663-4|LNC|Renal vessels Scan flow W Tc-99m glucoheptonate IV|Renal vessels Scan flow W Tc-99m glucoheptonate IV
C2826012|T102|strict|43665-9|LNC|Renal vessels Scan flow W Tc-99m Mertiatide IV|Renal vessels Scan flow W Tc-99m Mertiatide IV
C2826012|T102|strict|39870-1|LNC|Heart Scan flow W Tc-99m pertechnetate IV|Heart Scan flow W Tc-99m pertechnetate IV
C2826012|T102|strict|43654-3|LNC|Liver Scan flow W Tc-99m tagged RBC IV|Liver Scan flow W Tc-99m tagged RBC IV
C2826012|T102|strict|39685-3|LNC|Scan for abscess W GA-67 IV|Scan for abscess W GA-67 IV
C2826012|T102|strict|39940-2|LNC|Lung Scan Clearance W Tc-99m DTPA aerosol inhaled|Lung Scan Clearance W Tc-99m DTPA aerosol inhaled
C2826012|T102|strict|43787-1|LNC|Skull and Facial bones and Mandible X-ray for dental measurement|Skull and Facial bones and Mandible X-ray for dental measurement
C2826012|T102|strict|43648-5|LNC|Scan for endocrine tumor multiple areas W I-131 MIBG IV|Scan for endocrine tumor multiple areas W I-131 MIBG IV
C2826012|T102|strict|43649-3|LNC|Scan for endocrine tumor multiple areas W In-111 pentetreotide IV|Scan for endocrine tumor multiple areas W In-111 pentetreotide IV
C2826012|T102|strict|39827-1|LNC|Scan for endocrine tumor whole body W I-131 MIBG IV|Scan for endocrine tumor whole body W I-131 MIBG IV
C2826012|T102|strict|39828-9|LNC|Scan for endocrine tumor whole body W In-111 pentetreotide IV|Scan for endocrine tumor whole body W In-111 pentetreotide IV
C2826012|T102|strict|39327-2|LNC|Abdomen and Fetus X-ray for fetal age|Abdomen and Fetus X-ray for fetal age
C2826012|T102|strict|44208-7|LNC|Orbit X-ray for foreign body|Orbit X-ray for foreign body
C2826012|T102|strict|30720-7|LNC|Orbit - bilateral X-ray for foreign body|Orbit - bilateral X-ray for foreign body
C2826012|T102|strict|42311-1|LNC|Orbit - left X-ray for foreign body|Orbit - left X-ray for foreign body
C2826012|T102|strict|42312-9|LNC|Orbit - right X-ray for foreign body|Orbit - right X-ray for foreign body
C2826012|T102|strict|39768-7|LNC|Stomach Scan for gastric emptying W Tc-99m SC PO|Stomach Scan for gastric emptying W Tc-99m SC PO
C2826012|T102|strict|39767-9|LNC|Stomach Scan for gastric emptying liquid phase W radionuclide PO|Stomach Scan for gastric emptying liquid phase W radionuclide PO
C2826012|T102|strict|24997-9|LNC|Stomach Scan for gastric emptying solid phase W Tc-99m SC PO|Stomach Scan for gastric emptying solid phase W Tc-99m SC PO
C2826012|T102|strict|39769-5|LNC|Stomach Scan for gastric emptying W radionuclide PO|Stomach Scan for gastric emptying W radionuclide PO
C2826012|T102|strict|39892-5|LNC|Heart Scan for infarct and first pass|Heart Scan for infarct and first pass
C2826012|T102|strict|39891-7|LNC|Heart Scan for infarct and first pass W Tc-99m PYP IV|Heart Scan for infarct and first pass W Tc-99m PYP IV
C2826012|T102|strict|43646-9|LNC|Heart Scan for infarct qualitative and quantitative|Heart Scan for infarct qualitative and quantitative
C2826012|T102|strict|43645-1|LNC|Heart Scan for infarct qualitative|Heart Scan for infarct qualitative
C2826012|T102|strict|43647-7|LNC|Heart Scan for infarct quantitative|Heart Scan for infarct quantitative
C2826012|T102|strict|39653-1|LNC|Heart Scan for infarct|Heart Scan for infarct
C2826012|T102|strict|39657-2|LNC|Heart Scan for infarct W Tc-99m PYP IV|Heart Scan for infarct W Tc-99m PYP IV
C2826012|T102|strict|39933-7|LNC|Scan for infection multiple areas W GA-67 IV|Scan for infection multiple areas W GA-67 IV
C2826012|T102|strict|39830-5|LNC|Scan for infection whole body W GA-67 IV|Scan for infection whole body W GA-67 IV
C2826012|T102|strict|39677-0|LNC|Scan for infection W GA-67 IV|Scan for infection W GA-67 IV
C2826012|T102|strict|39490-8|LNC|Femur - right and Tibia - right X-ray for leg length|Femur - right and Tibia - right X-ray for leg length
C2826012|T102|strict|24700-7|LNC|Femur and Tibia X-ray for leg length|Femur and Tibia X-ray for leg length
C2826012|T102|strict|39686-1|LNC|Scan for lymphoma W GA-67 IV|Scan for lymphoma W GA-67 IV
C2826012|T102|strict|42170-1|LNC|Scan for lymphoma|Scan for lymphoma
C2826012|T102|strict|39672-1|LNC|Esophagus Scan for motility W radionuclide PO|Esophagus Scan for motility W radionuclide PO
C2826012|T102|strict|72256-1|LNC|Abdomen X-ray for motility with radioopaque markers|Abdomen X-ray for motility with radioopaque markers
C2826012|T102|strict|24571-2|LNC|Biliary ducts and Gallbladder Scan for patency of biliary structures and ejection fraction W sincalide and W radionuclide IV|Biliary ducts and Gallbladder Scan for patency of biliary structures and ejection fraction W sincalide and W radionuclide IV
C2826012|T102|strict|24572-0|LNC|Biliary ducts and Gallbladder Scan for patency of biliary structures W Tc-99m IV|Biliary ducts and Gallbladder Scan for patency of biliary structures W Tc-99m IV
C2826012|T102|strict|43788-9|LNC|Tube Fluoroscopy for patency W contrast via tube|Tube Fluoroscopy for patency W contrast via tube
C2826012|T102|strict|43789-7|LNC|Liver and Biliary ducts and Gallbladder Scan for patency W Tc-99m IV|Liver and Biliary ducts and Gallbladder Scan for patency W Tc-99m IV
C2826012|T102|strict|39673-9|LNC|Esophagus Scan for reflux W radionuclide PO|Esophagus Scan for reflux W radionuclide PO
C2826012|T102|strict|30650-6|LNC|Unspecified body region Fluoroscopy for shunt|Unspecified body region Fluoroscopy for shunt
C2826012|T102|strict|39665-5|LNC|Heart Scan for shunt detection|Heart Scan for shunt detection
C2826012|T102|strict|39664-8|LNC|Heart Scan for shunt detection W Tc-99m MAA IV|Heart Scan for shunt detection W Tc-99m MAA IV
C2826012|T102|strict|39848-7|LNC|Peritoneovenous shunt Scan for patency W In-111 IT|Peritoneovenous shunt Scan for patency W In-111 IT
C2826012|T102|strict|39849-5|LNC|Peritoneovenous shunt Scan for patency W radionuclide IT|Peritoneovenous shunt Scan for patency W radionuclide IT
C2826012|T102|strict|24876-5|LNC|Peritoneovenous shunt Scan for patency W Tc-99m DTPA IT|Peritoneovenous shunt Scan for patency W Tc-99m DTPA IT
C2826012|T102|strict|44149-3|LNC|Peritoneovenous shunt Scan for patency W Tc-99m MAA inj|Peritoneovenous shunt Scan for patency W Tc-99m MAA inj
C2826012|T102|strict|39954-3|LNC|Vein Scan for thrombosis|Vein Scan for thrombosis
C2826012|T102|strict|44140-2|LNC|Abdomen and Pelvis Scan for tumor|Abdomen and Pelvis Scan for tumor
C2826012|T102|strict|39831-3|LNC|Scan for tumor limited W GA-67 IV|Scan for tumor limited W GA-67 IV
C2826012|T102|strict|39951-9|LNC|Scan for tumor multiple area W Tc-99m Sestamibi IV|Scan for tumor multiple area W Tc-99m Sestamibi IV
C2826012|T102|strict|39934-5|LNC|Scan for tumor multiple areas W GA-67 IV|Scan for tumor multiple areas W GA-67 IV
C2826012|T102|strict|39829-7|LNC|Scan for tumor whole body W GA-67 IV|Scan for tumor whole body W GA-67 IV
C2826012|T102|strict|42171-9|LNC|Scan for tumor whole body|Scan for tumor whole body
C2826012|T102|strict|39749-7|LNC|Scan for tumor whole body W Tc-99m Sestamibi IV|Scan for tumor whole body W Tc-99m Sestamibi IV
C2826012|T102|strict|39679-6|LNC|Scan for tumor W GA-67 IV|Scan for tumor W GA-67 IV
C2826012|T102|strict|39750-5|LNC|Scan for tumor W Tc-99m Sestamibi IV|Scan for tumor W Tc-99m Sestamibi IV
C2826012|T102|strict|42305-3|LNC|Scan for tumor W Tl-201 IV|Scan for tumor W Tl-201 IV
C2826012|T102|strict|42397-0|LNC|Chest X-ray frontal stereo|Chest X-ray frontal stereo
C2826012|T102|strict|39923-8|LNC|Heart Scan gated and ejection fraction at rest and W radionuclide IV|Heart Scan gated and ejection fraction at rest and W radionuclide IV
C2826012|T102|strict|39917-0|LNC|Heart Scan gated and ejection fraction|Heart Scan gated and ejection fraction
C2826012|T102|strict|39919-6|LNC|Heart Scan gated and first pass|Heart Scan gated and first pass
C2826012|T102|strict|39925-3|LNC|Heart Scan gated and wall motion and ejection fraction at rest and W radionuclide IV|Heart Scan gated and wall motion and ejection fraction at rest and W radionuclide IV
C2826012|T102|strict|39931-1|LNC|Heart Scan gated and wall motion and ejection fraction|Heart Scan gated and wall motion and ejection fraction
C2826012|T102|strict|42306-1|LNC|Heart Scan gated and wall motion|Heart Scan gated and wall motion
C2826012|T102|strict|39929-5|LNC|Heart Scan gated and wall motion W stress and W radionuclide IV|Heart Scan gated and wall motion W stress and W radionuclide IV
C2826012|T102|strict|39921-2|LNC|Heart Scan gated at rest and W radionuclide IV|Heart Scan gated at rest and W radionuclide IV
C2826012|T102|strict|39924-6|LNC|Heart Scan gated at rest and W stress and W radionuclide IV|Heart Scan gated at rest and W stress and W radionuclide IV
C2826012|T102|strict|39922-0|LNC|Heart Scan gated at rest and W Tc-99m pertechnetate IV|Heart Scan gated at rest and W Tc-99m pertechnetate IV
C2826012|T102|strict|39920-4|LNC|Heart Scan gated at rest and W Tc-99m Sestamibi IV|Heart Scan gated at rest and W Tc-99m Sestamibi IV
C2826012|T102|strict|39915-4|LNC|Heart Scan gated|Heart Scan gated
C2826012|T102|strict|39928-7|LNC|Heart Scan gated W stress and W radionuclide IV|Heart Scan gated W stress and W radionuclide IV
C2826012|T102|strict|39927-9|LNC|Heart Scan gated W stress and W Tc-99m pertechnetate IV|Heart Scan gated W stress and W Tc-99m pertechnetate IV
C2826012|T102|strict|39914-7|LNC|Heart Scan gated W Tc-99m Sestamibi IV|Heart Scan gated W Tc-99m Sestamibi IV
C2826012|T102|strict|46348-9|LNC|Chest X-ray GE 2 and PA and Lateral views|Chest X-ray GE 2 and PA and Lateral views
C2826012|T102|strict|44210-3|LNC|Ankle X-ray GE 3 views|Ankle X-ray GE 3 views
C2826012|T102|strict|48480-8|LNC|Ankle - bilateral X-ray GE 3 views|Ankle - bilateral X-ray GE 3 views
C2826012|T102|strict|46390-1|LNC|Ankle - left X-ray GE 3 views|Ankle - left X-ray GE 3 views
C2826012|T102|strict|46347-1|LNC|Ankle - right X-ray GE 3 views|Ankle - right X-ray GE 3 views
C2826012|T102|strict|48481-6|LNC|Elbow - bilateral X-ray GE 3 views|Elbow - bilateral X-ray GE 3 views
C2826012|T102|strict|46344-8|LNC|Elbow - left X-ray GE 3 views|Elbow - left X-ray GE 3 views
C2826012|T102|strict|46345-5|LNC|Elbow - right X-ray GE 3 views|Elbow - right X-ray GE 3 views
C2826012|T102|strict|48479-0|LNC|Facial bones X-ray GE 3 views|Facial bones X-ray GE 3 views
C2826012|T102|strict|43492-8|LNC|Finger fifth - left X-ray GE 3 views|Finger fifth - left X-ray GE 3 views
C2826012|T102|strict|43497-7|LNC|Finger fifth - right X-ray GE 3 views|Finger fifth - right X-ray GE 3 views
C2826012|T102|strict|43491-0|LNC|Finger fourth - left X-ray GE 3 views|Finger fourth - left X-ray GE 3 views
C2826012|T102|strict|43496-9|LNC|Finger fourth - right X-ray GE 3 views|Finger fourth - right X-ray GE 3 views
C2826012|T102|strict|43489-4|LNC|Finger second - left X-ray GE 3 views|Finger second - left X-ray GE 3 views
C2826012|T102|strict|43494-4|LNC|Finger second - right X-ray GE 3 views|Finger second - right X-ray GE 3 views
C2826012|T102|strict|43490-2|LNC|Finger third - left X-ray GE 3 views|Finger third - left X-ray GE 3 views
C2826012|T102|strict|43495-1|LNC|Finger third - right X-ray GE 3 views|Finger third - right X-ray GE 3 views
C2826012|T102|strict|44188-1|LNC|Foot X-ray GE 3 views|Foot X-ray GE 3 views
C2826012|T102|strict|48478-2|LNC|Foot - bilateral X-ray GE 3 views|Foot - bilateral X-ray GE 3 views
C2826012|T102|strict|48477-4|LNC|Foot - left X-ray GE 3 views|Foot - left X-ray GE 3 views
C2826012|T102|strict|48476-6|LNC|Foot - right X-ray GE 3 views|Foot - right X-ray GE 3 views
C2826012|T102|strict|47370-2|LNC|Hand - left X-ray GE 3 views|Hand - left X-ray GE 3 views
C2826012|T102|strict|47371-0|LNC|Hand - right X-ray GE 3 views|Hand - right X-ray GE 3 views
C2826012|T102|strict|43498-5|LNC|Knee - left X-ray GE 3 views|Knee - left X-ray GE 3 views
C2826012|T102|strict|43482-9|LNC|Knee - right X-ray GE 3 views|Knee - right X-ray GE 3 views
C2826012|T102|strict|47381-9|LNC|Mastoid X-ray GE 3 views|Mastoid X-ray GE 3 views
C2826012|T102|strict|43543-8|LNC|Pelvis X-ray GE 3 views|Pelvis X-ray GE 3 views
C2826012|T102|strict|44189-9|LNC|Sacroiliac Joint X-ray GE 3 views|Sacroiliac Joint X-ray GE 3 views
C2826012|T102|strict|48746-2|LNC|Sacroiliac joint - bilateral X-ray GE 3 views|Sacroiliac joint - bilateral X-ray GE 3 views
C2826012|T102|strict|43486-0|LNC|Sinuses X-ray GE 3 views|Sinuses X-ray GE 3 views
C2826012|T102|strict|46377-8|LNC|Skull X-ray GE 3 views|Skull X-ray GE 3 views
C2826012|T102|strict|48482-4|LNC|Sternoclavicular Joints X-ray GE 3 views|Sternoclavicular Joints X-ray GE 3 views
C2826012|T102|strict|43488-6|LNC|Thumb - left X-ray GE 3 views|Thumb - left X-ray GE 3 views
C2826012|T102|strict|43493-6|LNC|Thumb - right X-ray GE 3 views|Thumb - right X-ray GE 3 views
C2826012|T102|strict|44190-7|LNC|Wrist X-ray GE 3 views|Wrist X-ray GE 3 views
C2826012|T102|strict|48483-2|LNC|Wrist - bilateral X-ray GE 3 views|Wrist - bilateral X-ray GE 3 views
C2826012|T102|strict|46346-3|LNC|Wrist - left X-ray GE 3 views|Wrist - left X-ray GE 3 views
C2826012|T102|strict|46343-0|LNC|Wrist - right X-ray GE 3 views|Wrist - right X-ray GE 3 views
C2826012|T102|strict|48485-7|LNC|Ribs - bilateral and Chest X-ray GE 3 and PA Chest views|Ribs - bilateral and Chest X-ray GE 3 and PA Chest views
C2826012|T102|strict|48486-5|LNC|Ribs - left and Chest X-ray GE 3 and PA Chest views|Ribs - left and Chest X-ray GE 3 and PA Chest views
C2826012|T102|strict|48484-0|LNC|Ribs - right and Chest X-ray GE 3 and PA Chest views|Ribs - right and Chest X-ray GE 3 and PA Chest views
C2826012|T102|strict|44191-5|LNC|Ribs and Chest X-ray GE 3 and PA Chest views|Ribs and Chest X-ray GE 3 and PA Chest views
C2826012|T102|strict|44239-2|LNC|Ribs - unilateral and Chest X-ray Ge 3 and PA Chest Portable views|Ribs - unilateral and Chest X-ray Ge 3 and PA Chest Portable views
C2826012|T102|strict|44193-1|LNC|Hand X-ray GE 3 Portable views|Hand X-ray GE 3 Portable views
C2826012|T102|strict|44192-3|LNC|Pelvis X-ray GE 3 Portable views|Pelvis X-ray GE 3 Portable views
C2826012|T102|strict|44211-1|LNC|Chest X-ray GE 4 views|Chest X-ray GE 4 views
C2826012|T102|strict|47367-8|LNC|Chest Fluoroscopy GE 4 views|Chest Fluoroscopy GE 4 views
C2826012|T102|strict|47374-4|LNC|Knee - left X-ray GE 4 views|Knee - left X-ray GE 4 views
C2826012|T102|strict|47376-9|LNC|Knee - right X-ray GE 4 views|Knee - right X-ray GE 4 views
C2826012|T102|strict|47379-3|LNC|Mandible X-ray GE 4 views|Mandible X-ray GE 4 views
C2826012|T102|strict|48747-0|LNC|Orbit - bilateral X-ray GE 4 views|Orbit - bilateral X-ray GE 4 views
C2826012|T102|strict|48487-3|LNC|Skull X-ray GE 4 views|Skull X-ray GE 4 views
C2826012|T102|strict|44212-9|LNC|Spine Cervical X-ray GE 4 views|Spine Cervical X-ray GE 4 views
C2826012|T102|strict|47382-7|LNC|Spine Lumbar X-ray GE 4 views|Spine Lumbar X-ray GE 4 views
C2826012|T102|strict|47368-6|LNC|Chest X-ray GE 4 and Pa and Lateral views|Chest X-ray GE 4 and Pa and Lateral views
C2826012|T102|strict|44194-9|LNC|Spine X-ray GE 4 views W right bending and W left bending|Spine X-ray GE 4 views W right bending and W left bending
C2826012|T102|strict|44195-6|LNC|Knee X-ray GE 5 views|Knee X-ray GE 5 views
C2826012|T102|strict|43524-8|LNC|Skull X-ray GE 5 views|Skull X-ray GE 5 views
C2826012|T102|strict|44197-2|LNC|Knee - bilateral X-ray GE 5 views standing|Knee - bilateral X-ray GE 5 views standing
C2826012|T102|strict|44196-4|LNC|Spine Lumbar X-ray GE 5 views W right bending and W left bending|Spine Lumbar X-ray GE 5 views W right bending and W left bending
C2826012|T102|strict|49570-5|LNC|Ankle - bilateral X-ray GE 6 views|Ankle - bilateral X-ray GE 6 views
C2826012|T102|strict|37160-9|LNC|Shoulder - left X-ray Grashey and axillary|Shoulder - left X-ray Grashey and axillary
C2826012|T102|strict|38793-6|LNC|Shoulder - right X-ray Grashey and axillary|Shoulder - right X-ray Grashey and axillary
C2826012|T102|strict|37158-3|LNC|Shoulder - left X-ray Grashey and axillary and outlet|Shoulder - left X-ray Grashey and axillary and outlet
C2826012|T102|strict|37806-7|LNC|Shoulder - right X-ray Grashey and axillary and outlet|Shoulder - right X-ray Grashey and axillary and outlet
C2826012|T102|strict|37161-7|LNC|Shoulder - bilateral X-ray Grashey and axillary and outlet and Zanca|Shoulder - bilateral X-ray Grashey and axillary and outlet and Zanca
C2826012|T102|strict|69267-3|LNC|Shoulder X-ray Grashey and axillary and Y|Shoulder X-ray Grashey and axillary and Y
C2826012|T102|strict|37538-6|LNC|Shoulder - left X-ray Grashey and axillary and Y|Shoulder - left X-ray Grashey and axillary and Y
C2826012|T102|strict|38789-4|LNC|Shoulder - right X-ray Grashey and axillary and Y|Shoulder - right X-ray Grashey and axillary and Y
C2826012|T102|strict|37157-5|LNC|Shoulder - left X-ray Grashey and outlet|Shoulder - left X-ray Grashey and outlet
C2826012|T102|strict|38791-0|LNC|Shoulder - right X-ray Grashey and outlet|Shoulder - right X-ray Grashey and outlet
C2826012|T102|strict|39350-4|LNC|Shoulder - bilateral X-ray Grashey and outlet and Serendipity|Shoulder - bilateral X-ray Grashey and outlet and Serendipity
C2826012|T102|strict|37162-5|LNC|Shoulder - left X-ray Grashey and outlet and Serendipity|Shoulder - left X-ray Grashey and outlet and Serendipity
C2826012|T102|strict|38794-4|LNC|Shoulder - right X-ray Grashey and outlet and Serendipity|Shoulder - right X-ray Grashey and outlet and Serendipity
C2826012|T102|strict|37167-4|LNC|Shoulder - left X-ray Grashey and West Point|Shoulder - left X-ray Grashey and West Point
C2826012|T102|strict|38795-1|LNC|Shoulder - right X-ray Grashey and West Point|Shoulder - right X-ray Grashey and West Point
C2826012|T102|strict|69156-8|LNC|Shoulder - left X-ray Grashey and Y|Shoulder - left X-ray Grashey and Y
C2826012|T102|strict|43790-5|LNC|Shoulder - right X-ray Grashey and Y|Shoulder - right X-ray Grashey and Y
C2826012|T102|strict|38004-8|LNC|Shoulder - left X-ray Grashey W and WO weight|Shoulder - left X-ray Grashey W and WO weight
C2826012|T102|strict|38816-5|LNC|Shoulder - right X-ray Grashey W and WO weight|Shoulder - right X-ray Grashey W and WO weight
C2826012|T102|strict|37539-4|LNC|Breast Mammogram grid|Breast Mammogram grid
C2826012|T102|strict|37540-2|LNC|Knee - bilateral X-ray Holmblad standing|Knee - bilateral X-ray Holmblad standing
C2826012|T102|strict|30771-0|LNC|Pelvis X-ray inlet and outlet|Pelvis X-ray inlet and outlet
C2826012|T102|strict|37627-7|LNC|Pelvis X-ray inlet and outlet and oblique|Pelvis X-ray inlet and outlet and oblique
C2826012|T102|strict|37164-1|LNC|Facial bones X-ray lateral and Caldwell and Waters|Facial bones X-ray lateral and Caldwell and Waters
C2826012|T102|strict|37864-6|LNC|Sinuses X-ray lateral and Caldwell and Waters|Sinuses X-ray lateral and Caldwell and Waters
C2826012|T102|strict|37165-8|LNC|Facial bones X-ray lateral and Caldwell and Waters and submentovertex|Facial bones X-ray lateral and Caldwell and Waters and submentovertex
C2826012|T102|strict|37166-6|LNC|Facial bones X-ray lateral and Caldwell and Waters and submentovertex and Towne|Facial bones X-ray lateral and Caldwell and Waters and submentovertex and Towne
C2826012|T102|strict|37871-1|LNC|Skull X-ray lateral and Caldwell and Waters and Towne|Skull X-ray lateral and Caldwell and Waters and Towne
C2826012|T102|strict|37134-4|LNC|Ankle - bilateral X-ray lateral and Mortise|Ankle - bilateral X-ray lateral and Mortise
C2826012|T102|strict|37135-1|LNC|Ankle - left X-ray lateral and Mortise|Ankle - left X-ray lateral and Mortise
C2826012|T102|strict|37670-7|LNC|Ankle - right X-ray lateral and Mortise|Ankle - right X-ray lateral and Mortise
C2826012|T102|strict|42382-2|LNC|Ankle - left X-ray lateral and Mortise and Broden W manual stress|Ankle - left X-ray lateral and Mortise and Broden W manual stress
C2826012|T102|strict|39366-0|LNC|Scapula X-ray lateral and outlet|Scapula X-ray lateral and outlet
C2826012|T102|strict|43464-7|LNC|Ribs - bilateral and Chest X-ray lateral and PA chest|Ribs - bilateral and Chest X-ray lateral and PA chest
C2826012|T102|strict|37603-8|LNC|Ribs - left and Chest X-ray lateral and PA chest|Ribs - left and Chest X-ray lateral and PA chest
C2826012|T102|strict|39100-3|LNC|Ribs - right and Chest X-ray lateral and PA chest|Ribs - right and Chest X-ray lateral and PA chest
C2826012|T102|strict|39101-1|LNC|Ribs and Chest X-ray lateral and PA chest|Ribs and Chest X-ray lateral and PA chest
C2826012|T102|strict|39341-3|LNC|Chest X-ray lateral and PA W inspiration and expiration|Chest X-ray lateral and PA W inspiration and expiration
C2826012|T102|strict|39406-4|LNC|Sternum X-ray lateral and right anterior oblique|Sternum X-ray lateral and right anterior oblique
C2826012|T102|strict|39405-6|LNC|Sternum X-ray lateral and right oblique and left oblique|Sternum X-ray lateral and right oblique and left oblique
C2826012|T102|strict|42436-6|LNC|Sella turcica X-ray lateral and Towne|Sella turcica X-ray lateral and Towne
C2826012|T102|strict|37869-5|LNC|Skull X-ray lateral and Towne|Skull X-ray lateral and Towne
C2826012|T102|strict|37605-3|LNC|Nasal bones X-ray lateral and Waters|Nasal bones X-ray lateral and Waters
C2826012|T102|strict|37862-0|LNC|Sinuses X-ray lateral and Waters|Sinuses X-ray lateral and Waters
C2826012|T102|strict|37136-9|LNC|Shoulder - left X-ray lateral and Y|Shoulder - left X-ray lateral and Y
C2826012|T102|strict|37803-4|LNC|Shoulder - right X-ray lateral and Y|Shoulder - right X-ray lateral and Y
C2826012|T102|strict|39340-5|LNC|Spine Lumbar X-ray lateral standing and W flexion and W extension|Spine Lumbar X-ray lateral standing and W flexion and W extension
C2826012|T102|strict|37133-6|LNC|Spine Cervical X-ray lateral W flexion and W extension|Spine Cervical X-ray lateral W flexion and W extension
C2826012|T102|strict|37132-8|LNC|Spine Lumbar X-ray lateral W flexion and W extension|Spine Lumbar X-ray lateral W flexion and W extension
C2826012|T102|strict|38010-5|LNC|Spine Thoracic X-ray lateral W flexion and W extension|Spine Thoracic X-ray lateral W flexion and W extension
C2826012|T102|strict|37929-7|LNC|Wrist X-ray lateral W flexion and W extension|Wrist X-ray lateral W flexion and W extension
C2826012|T102|strict|69157-6|LNC|Wrist - left X-ray lateral W flexion and W extension|Wrist - left X-ray lateral W flexion and W extension
C2826012|T102|strict|39515-2|LNC|Wrist - right X-ray lateral W flexion and W extension|Wrist - right X-ray lateral W flexion and W extension
C2826012|T102|strict|37474-4|LNC|Ankle - left X-ray lateral W manual stress|Ankle - left X-ray lateral W manual stress
C2826012|T102|strict|37669-9|LNC|Ankle - right X-ray lateral W manual stress|Ankle - right X-ray lateral W manual stress
C2826012|T102|strict|43480-3|LNC|Joint X-ray lateral W manual stress|Joint X-ray lateral W manual stress
C2826012|T102|strict|37541-0|LNC|Mastoid - bilateral X-ray law and Mayer and Stenver and Towne|Mastoid - bilateral X-ray law and Mayer and Stenver and Towne
C2826012|T102|strict|47380-1|LNC|Mandible X-ray LE 3 views|Mandible X-ray LE 3 views
C2826012|T102|strict|43470-4|LNC|Skull X-ray LE 3 views|Skull X-ray LE 3 views
C2826012|T102|strict|47377-7|LNC|Knee - right X-ray LE 4 views|Knee - right X-ray LE 4 views
C2826012|T102|strict|24610-8|LNC|Breast Mammogram limited|Breast Mammogram limited
C2826012|T102|strict|26287-3|LNC|Breast - bilateral Mammogram limited|Breast - bilateral Mammogram limited
C2826012|T102|strict|26289-9|LNC|Breast - left Mammogram limited|Breast - left Mammogram limited
C2826012|T102|strict|26291-5|LNC|Breast - right Mammogram limited|Breast - right Mammogram limited
C2826012|T102|strict|41826-9|LNC|Elbow - left X-ray limited|Elbow - left X-ray limited
C2826012|T102|strict|41785-7|LNC|Elbow - right X-ray limited|Elbow - right X-ray limited
C2826012|T102|strict|36737-5|LNC|Facial bones X-ray limited|Facial bones X-ray limited
C2826012|T102|strict|41830-1|LNC|Hand - left X-ray limited|Hand - left X-ray limited
C2826012|T102|strict|41789-9|LNC|Hand - right X-ray limited|Hand - right X-ray limited
C2826012|T102|strict|36738-3|LNC|Mandible X-ray limited|Mandible X-ray limited
C2826012|T102|strict|36893-6|LNC|Mastoid X-ray limited|Mastoid X-ray limited
C2826012|T102|strict|42007-5|LNC|Mastoid - bilateral X-ray limited|Mastoid - bilateral X-ray limited
C2826012|T102|strict|37646-7|LNC|Sacroiliac Joint X-ray limited|Sacroiliac Joint X-ray limited
C2826012|T102|strict|44209-5|LNC|Sinuses X-ray limited|Sinuses X-ray limited
C2826012|T102|strict|48466-7|LNC|Skull X-ray limited|Skull X-ray limited
C2826012|T102|strict|42710-4|LNC|Spine Cervical X-ray limited|Spine Cervical X-ray limited
C2826012|T102|strict|36739-1|LNC|Wrist - bilateral X-ray limited|Wrist - bilateral X-ray limited
C2826012|T102|strict|38838-9|LNC|Wrist - left X-ray limited|Wrist - left X-ray limited
C2826012|T102|strict|37642-6|LNC|Wrist - right X-ray limited|Wrist - right X-ray limited
C2826012|T102|strict|41797-2|LNC|Colon Fluoroscopy limited W air and barium contrast PR|Colon Fluoroscopy limited W air and barium contrast PR
C2826012|T102|strict|42335-0|LNC|Spine Cervical Fluoroscopy limited W contrast IT|Spine Cervical Fluoroscopy limited W contrast IT
C2826012|T102|strict|38125-1|LNC|Spine Cervical and Thoracic and Lumbar Fluoroscopy limited W contrast IT|Spine Cervical and Thoracic and Lumbar Fluoroscopy limited W contrast IT
C2826012|T102|strict|38120-2|LNC|Spine Thoracic Fluoroscopy limited W contrast IT|Spine Thoracic Fluoroscopy limited W contrast IT
C2826012|T102|strict|37137-7|LNC|Kidney X-ray limited W contrast IV|Kidney X-ray limited W contrast IV
C2826012|T102|strict|39687-9|LNC|Scan limited W GA-67 IV|Scan limited W GA-67 IV
C2826012|T102|strict|39754-7|LNC|Thyroid Scan limited W I-131 IV|Thyroid Scan limited W I-131 IV
C2826012|T102|strict|49571-3|LNC|Scan limited W I-131 MIBG IV|Scan limited W I-131 MIBG IV
C2826012|T102|strict|39843-8|LNC|Scan limited W In-111 Satumomab IV|Scan limited W In-111 Satumomab IV
C2826012|T102|strict|41836-8|LNC|Bone Scan limited W In-111 tagged WBC IV|Bone Scan limited W In-111 tagged WBC IV
C2826012|T102|strict|39627-5|LNC|Bone Scan limited|Bone Scan limited
C2826012|T102|strict|39822-2|LNC|Bone marrow Scan limited|Bone marrow Scan limited
C2826012|T102|strict|39645-7|LNC|Breast Scan limited|Breast Scan limited
C2826012|T102|strict|39695-2|LNC|Lung Scan limited|Lung Scan limited
C2826012|T102|strict|39936-0|LNC|Joint Scan limited|Joint Scan limited
C2826012|T102|strict|37542-8|LNC|Breast Mammogram magnification|Breast Mammogram magnification
C2826012|T102|strict|37543-6|LNC|Breast - bilateral Mammogram magnification|Breast - bilateral Mammogram magnification
C2826012|T102|strict|37554-3|LNC|Breast - bilateral Mammogram magnification and spot|Breast - bilateral Mammogram magnification and spot
C2826012|T102|strict|38854-6|LNC|Breast - left Mammogram magnification and spot|Breast - left Mammogram magnification and spot
C2826012|T102|strict|37769-7|LNC|Breast - right Mammogram magnification and spot|Breast - right Mammogram magnification and spot
C2826012|T102|strict|30769-4|LNC|Pelvis and Hip - bilateral X-ray max abduction|Pelvis and Hip - bilateral X-ray max abduction
C2826012|T102|strict|38086-5|LNC|Knee X-ray Merchants 30 and 45 and 60 degrees|Knee X-ray Merchants 30 and 45 and 60 degrees
C2826012|T102|strict|39935-2|LNC|Scan multiple areas W GA-67 IV|Scan multiple areas W GA-67 IV
C2826012|T102|strict|39949-3|LNC|Scan multiple areas W In-111 Satumomab IV|Scan multiple areas W In-111 Satumomab IV
C2826012|T102|strict|39904-8|LNC|Bone Scan multiple areas|Bone Scan multiple areas
C2826012|T102|strict|39907-1|LNC|Bone marrow Scan multiple areas|Bone marrow Scan multiple areas
C2826012|T102|strict|39937-8|LNC|Joint Scan multiple areas|Joint Scan multiple areas
C2826012|T102|strict|39950-1|LNC|Prostate Scan multiple areas W Tc-99m capromab pendatide IV|Prostate Scan multiple areas W Tc-99m capromab pendatide IV
C2826012|T102|strict|36608-8|LNC|Elbow X-ray oblique|Elbow X-ray oblique
C2826012|T102|strict|36740-9|LNC|Elbow - bilateral X-ray oblique|Elbow - bilateral X-ray oblique
C2826012|T102|strict|36741-7|LNC|Elbow - left X-ray oblique|Elbow - left X-ray oblique
C2826012|T102|strict|37687-1|LNC|Elbow - right X-ray oblique|Elbow - right X-ray oblique
C2826012|T102|strict|36744-1|LNC|Humerus - left X-ray oblique|Humerus - left X-ray oblique
C2826012|T102|strict|37737-4|LNC|Humerus - right X-ray oblique|Humerus - right X-ray oblique
C2826012|T102|strict|36619-5|LNC|Knee X-ray oblique|Knee X-ray oblique
C2826012|T102|strict|36745-8|LNC|Knee - bilateral X-ray oblique|Knee - bilateral X-ray oblique
C2826012|T102|strict|36746-6|LNC|Knee - left X-ray oblique|Knee - left X-ray oblique
C2826012|T102|strict|37757-2|LNC|Knee - right X-ray oblique|Knee - right X-ray oblique
C2826012|T102|strict|36747-4|LNC|Mandible X-ray oblique|Mandible X-ray oblique
C2826012|T102|strict|37630-1|LNC|Pelvis X-ray oblique|Pelvis X-ray oblique
C2826012|T102|strict|36742-5|LNC|Radius - bilateral and Ulna - bilateral X-ray oblique|Radius - bilateral and Ulna - bilateral X-ray oblique
C2826012|T102|strict|36743-3|LNC|Radius - left and Ulna.left X-ray oblique|Radius - left and Ulna.left X-ray oblique
C2826012|T102|strict|37709-3|LNC|Radius - right and Ulna - right X-ray oblique|Radius - right and Ulna - right X-ray oblique
C2826012|T102|strict|48748-8|LNC|Spine X-ray oblique|Spine X-ray oblique
C2826012|T102|strict|36748-2|LNC|Spine Cervical X-ray oblique|Spine Cervical X-ray oblique
C2826012|T102|strict|43791-3|LNC|Spine Lumbar X-ray oblique|Spine Lumbar X-ray oblique
C2826012|T102|strict|48749-6|LNC|Spine Thoracic X-ray oblique|Spine Thoracic X-ray oblique
C2826012|T102|strict|36749-0|LNC|Tibia - left and Fibula - left X-ray oblique|Tibia - left and Fibula - left X-ray oblique
C2826012|T102|strict|37817-4|LNC|Tibia - right and Fibula - right X-ray oblique|Tibia - right and Fibula - right X-ray oblique
C2826012|T102|strict|36894-4|LNC|Tibia and Fibula X-ray oblique|Tibia and Fibula X-ray oblique
C2826012|T102|strict|37544-4|LNC|Wrist - bilateral X-ray oblique|Wrist - bilateral X-ray oblique
C2826012|T102|strict|38839-7|LNC|Wrist - left X-ray oblique|Wrist - left X-ray oblique
C2826012|T102|strict|37643-4|LNC|Wrist - right X-ray oblique|Wrist - right X-ray oblique
C2826012|T102|strict|42398-8|LNC|Foot X-ray oblique and (AP and lateral) standing|Foot X-ray oblique and (AP and lateral) standing
C2826012|T102|strict|37139-3|LNC|Spine Cervical X-ray oblique and lateral W flexion and W extension|Spine Cervical X-ray oblique and lateral W flexion and W extension
C2826012|T102|strict|37154-2|LNC|Knee X-ray oblique and Sunrise|Knee X-ray oblique and Sunrise
C2826012|T102|strict|37155-9|LNC|Knee X-ray oblique and Sunrise and tunnel|Knee X-ray oblique and Sunrise and tunnel
C2826012|T102|strict|43469-6|LNC|Unspecified body region X-ray of foreign body|Unspecified body region X-ray of foreign body
C2826012|T102|strict|37063-5|LNC|Unspecified body region Fluoroscopy of foreign body|Unspecified body region Fluoroscopy of foreign body
C2826012|T102|strict|37546-9|LNC|Temporomandibular joint - bilateral X-ray open and closed mouth|Temporomandibular joint - bilateral X-ray open and closed mouth
C2826012|T102|strict|48491-5|LNC|Temporomandibular joint - left X-ray open and closed mouth|Temporomandibular joint - left X-ray open and closed mouth
C2826012|T102|strict|48490-7|LNC|Temporomandibular joint - right X-ray open and closed mouth|Temporomandibular joint - right X-ray open and closed mouth
C2826012|T102|strict|48699-3|LNC|Temporomandibular Joint - unilateral X-ray open and closed mouth|Temporomandibular Joint - unilateral X-ray open and closed mouth
C2826012|T102|strict|37152-6|LNC|Shoulder - bilateral X-ray outlet and Y|Shoulder - bilateral X-ray outlet and Y
C2826012|T102|strict|37140-1|LNC|Shoulder - left X-ray outlet and Y|Shoulder - left X-ray outlet and Y
C2826012|T102|strict|37804-2|LNC|Shoulder - right X-ray outlet and Y|Shoulder - right X-ray outlet and Y
C2826012|T102|strict|36750-8|LNC|Chest X-ray PA and AP lateral-decubitus|Chest X-ray PA and AP lateral-decubitus
C2826012|T102|strict|42272-5|LNC|Chest X-ray PA and lateral|Chest X-ray PA and lateral
C2826012|T102|strict|36751-6|LNC|Chest Fluoroscopy PA and lateral|Chest Fluoroscopy PA and lateral
C2826012|T102|strict|36752-4|LNC|Hand - bilateral X-ray PA and lateral|Hand - bilateral X-ray PA and lateral
C2826012|T102|strict|36753-2|LNC|Hand - left X-ray PA and lateral|Hand - left X-ray PA and lateral
C2826012|T102|strict|37713-5|LNC|Hand - right X-ray PA and lateral|Hand - right X-ray PA and lateral
C2826012|T102|strict|36754-0|LNC|Mandible X-ray PA and lateral|Mandible X-ray PA and lateral
C2826012|T102|strict|30721-5|LNC|Sinuses X-ray PA and lateral|Sinuses X-ray PA and lateral
C2826012|T102|strict|37547-7|LNC|Wrist - bilateral X-ray PA and lateral|Wrist - bilateral X-ray PA and lateral
C2826012|T102|strict|37548-5|LNC|Wrist - left X-ray PA and lateral|Wrist - left X-ray PA and lateral
C2826012|T102|strict|37835-6|LNC|Wrist - right X-ray PA and lateral|Wrist - right X-ray PA and lateral
C2826012|T102|strict|37143-5|LNC|Chest X-ray PA and lateral and AP lateral-decubitus|Chest X-ray PA and lateral and AP lateral-decubitus
C2826012|T102|strict|37144-3|LNC|Chest X-ray PA and lateral and AP left lateral-decubitus|Chest X-ray PA and lateral and AP left lateral-decubitus
C2826012|T102|strict|37145-0|LNC|Chest X-ray PA and lateral and AP right lateral-decubitus|Chest X-ray PA and lateral and AP right lateral-decubitus
C2826012|T102|strict|37142-7|LNC|Hand - bilateral X-ray PA and lateral and Ball Catcher|Hand - bilateral X-ray PA and lateral and Ball Catcher
C2826012|T102|strict|37860-4|LNC|Sinuses X-ray PA and lateral and Caldwell and Waters|Sinuses X-ray PA and lateral and Caldwell and Waters
C2826012|T102|strict|37146-8|LNC|Chest X-ray PA and lateral and left oblique|Chest X-ray PA and lateral and left oblique
C2826012|T102|strict|30741-3|LNC|Chest X-ray PA and lateral and lordotic upright|Chest X-ray PA and lateral and lordotic upright
C2826012|T102|strict|39078-1|LNC|Finger X-ray PA and lateral and oblique|Finger X-ray PA and lateral and oblique
C2826012|T102|strict|36755-7|LNC|Hand X-ray PA and lateral and oblique|Hand X-ray PA and lateral and oblique
C2826012|T102|strict|36756-5|LNC|Hand - bilateral X-ray PA and lateral and oblique|Hand - bilateral X-ray PA and lateral and oblique
C2826012|T102|strict|36757-3|LNC|Hand - left X-ray PA and lateral and oblique|Hand - left X-ray PA and lateral and oblique
C2826012|T102|strict|37715-0|LNC|Hand - right X-ray PA and lateral and oblique|Hand - right X-ray PA and lateral and oblique
C2826012|T102|strict|37884-4|LNC|Sternum X-ray PA and lateral and oblique|Sternum X-ray PA and lateral and oblique
C2826012|T102|strict|37549-3|LNC|Wrist - bilateral X-ray PA and lateral and oblique|Wrist - bilateral X-ray PA and lateral and oblique
C2826012|T102|strict|37550-1|LNC|Wrist - left X-ray PA and lateral and oblique|Wrist - left X-ray PA and lateral and oblique
C2826012|T102|strict|37836-4|LNC|Wrist - right X-ray PA and lateral and oblique|Wrist - right X-ray PA and lateral and oblique
C2826012|T102|strict|36758-1|LNC|Chest X-ray PA and lateral and oblique and lordotic|Chest X-ray PA and lateral and oblique and lordotic
C2826012|T102|strict|37148-4|LNC|Mandible X-ray PA and lateral and oblique and Towne|Mandible X-ray PA and lateral and oblique and Towne
C2826012|T102|strict|37147-6|LNC|Chest X-ray PA and lateral and right oblique|Chest X-ray PA and lateral and right oblique
C2826012|T102|strict|30742-1|LNC|Chest X-ray PA and lateral and right oblique and left oblique|Chest X-ray PA and lateral and right oblique and left oblique
C2826012|T102|strict|30743-9|LNC|Chest X-ray PA and lateral and right oblique and left oblique portable|Chest X-ray PA and lateral and right oblique and left oblique portable
C2826012|T102|strict|30744-7|LNC|Chest X-ray PA and lateral and right or-left oblique|Chest X-ray PA and lateral and right or-left oblique
C2826012|T102|strict|24643-9|LNC|Chest X-ray PA and lateral and right or-left oblique upright|Chest X-ray PA and lateral and right or-left oblique upright
C2826012|T102|strict|37149-2|LNC|Patella - left X-ray PA and lateral and Sunrise|Patella - left X-ray PA and lateral and Sunrise
C2826012|T102|strict|38790-2|LNC|Patella - right X-ray PA and lateral and Sunrise|Patella - right X-ray PA and lateral and Sunrise
C2826012|T102|strict|37859-6|LNC|Sinuses X-ray PA and lateral and Waters|Sinuses X-ray PA and lateral and Waters
C2826012|T102|strict|69271-5|LNC|Skull X-ray PA and lateral and Waters and Towne|Skull X-ray PA and lateral and Waters and Towne
C2826012|T102|strict|24647-0|LNC|Chest X-ray PA and lateral upright|Chest X-ray PA and lateral upright
C2826012|T102|strict|24644-7|LNC|Chest X-ray PA and lateral upright portable|Chest X-ray PA and lateral upright portable
C2826012|T102|strict|36759-9|LNC|Chest X-ray PA and lordotic|Chest X-ray PA and lordotic
C2826012|T102|strict|39079-9|LNC|Hand X-ray PA and oblique|Hand X-ray PA and oblique
C2826012|T102|strict|37141-9|LNC|Chest X-ray PA and right lateral|Chest X-ray PA and right lateral
C2826012|T102|strict|39519-4|LNC|Skull X-ray PA and right lateral and left lateral|Skull X-ray PA and right lateral and left lateral
C2826012|T102|strict|39521-0|LNC|Skull X-ray PA and right lateral and left lateral and Caldwell and Towne|Skull X-ray PA and right lateral and left lateral and Caldwell and Towne
C2826012|T102|strict|39520-2|LNC|Skull X-ray PA and right lateral and left lateral and Towne|Skull X-ray PA and right lateral and left lateral and Towne
C2826012|T102|strict|24646-2|LNC|Chest X-ray PA and right lateral and right oblique and left oblique upright|Chest X-ray PA and right lateral and right oblique and left oblique upright
C2826012|T102|strict|24645-4|LNC|Chest X-ray PA and right lateral and right oblique and left oblique upright portable|Chest X-ray PA and right lateral and right oblique and left oblique upright portable
C2826012|T102|strict|37150-0|LNC|Chest X-ray PA and right oblique and left oblique|Chest X-ray PA and right oblique and left oblique
C2826012|T102|strict|24635-5|LNC|Chest X-ray PA upright W inspiration and expiration|Chest X-ray PA upright W inspiration and expiration
C2826012|T102|strict|46378-6|LNC|Knee - bilateral X-ray PA standing and W flexion|Knee - bilateral X-ray PA standing and W flexion
C2826012|T102|strict|43660-0|LNC|Heart Scan perfusion qualitative at rest and W radionuclide IV|Heart Scan perfusion qualitative at rest and W radionuclide IV
C2826012|T102|strict|43661-8|LNC|Heart Scan perfusion quantitative at rest and W radionuclide IV|Heart Scan perfusion quantitative at rest and W radionuclide IV
C2826012|T102|strict|43658-4|LNC|Heart Scan perfusion quantitative|Heart Scan perfusion quantitative
C2826012|T102|strict|43656-8|LNC|Lung Scan perfusion quantitative|Lung Scan perfusion quantitative
C2826012|T102|strict|39719-0|LNC|Heart Scan perfusion at rest and W adenosine and W radionuclide IV|Heart Scan perfusion at rest and W adenosine and W radionuclide IV
C2826012|T102|strict|43777-2|LNC|Heart Scan perfusion at rest and W adenosine and W Tl-201 IV|Heart Scan perfusion at rest and W adenosine and W Tl-201 IV
C2826012|T102|strict|39722-4|LNC|Heart Scan perfusion at rest and W dipyridamole and W radionuclide IV|Heart Scan perfusion at rest and W dipyridamole and W radionuclide IV
C2826012|T102|strict|39720-8|LNC|Heart Scan perfusion at rest and W dipyridamole and W Tc-99m Sestamibi IV|Heart Scan perfusion at rest and W dipyridamole and W Tc-99m Sestamibi IV
C2826012|T102|strict|39728-1|LNC|Heart Scan perfusion at rest and W radionuclide IV|Heart Scan perfusion at rest and W radionuclide IV
C2826012|T102|strict|39726-5|LNC|Heart Scan perfusion at rest and W stress and W radionuclide IV|Heart Scan perfusion at rest and W stress and W radionuclide IV
C2826012|T102|strict|39727-3|LNC|Heart Scan perfusion at rest and W stress and W Tc-99m Sestamibi IV|Heart Scan perfusion at rest and W stress and W Tc-99m Sestamibi IV
C2826012|T102|strict|39699-4|LNC|Heart Scan perfusion at rest and W Tc-99m Sestamibi IV|Heart Scan perfusion at rest and W Tc-99m Sestamibi IV
C2826012|T102|strict|39701-8|LNC|Heart Scan perfusion W adenosine and W radionuclide IV|Heart Scan perfusion W adenosine and W radionuclide IV
C2826012|T102|strict|39731-5|LNC|Heart Scan perfusion W adenosine and W Tc-99m Sestamibi IV|Heart Scan perfusion W adenosine and W Tc-99m Sestamibi IV
C2826012|T102|strict|39735-6|LNC|Heart Scan perfusion W adenosine and W Tl-201 IV|Heart Scan perfusion W adenosine and W Tl-201 IV
C2826012|T102|strict|39708-3|LNC|Heart Scan perfusion W dipyridamole and W radionuclide IV|Heart Scan perfusion W dipyridamole and W radionuclide IV
C2826012|T102|strict|39709-1|LNC|Heart Scan perfusion W dipyridamole and W Tc-99m IV|Heart Scan perfusion W dipyridamole and W Tc-99m IV
C2826012|T102|strict|39705-9|LNC|Heart Scan perfusion W dipyridamole and W Tc-99m Sestamibi IV|Heart Scan perfusion W dipyridamole and W Tc-99m Sestamibi IV
C2826012|T102|strict|39707-5|LNC|Heart Scan perfusion W dipyridamole and W Tl-201 IV|Heart Scan perfusion W dipyridamole and W Tl-201 IV
C2826012|T102|strict|39703-4|LNC|Heart Scan perfusion W dobutamine and W radionuclide IV|Heart Scan perfusion W dobutamine and W radionuclide IV
C2826012|T102|strict|39702-6|LNC|Heart Scan perfusion W dobutamine and W Tc-99m Sestamibi IV|Heart Scan perfusion W dobutamine and W Tc-99m Sestamibi IV
C2826012|T102|strict|39733-1|LNC|Heart Scan perfusion W dobutamine and W Tl-201 IV|Heart Scan perfusion W dobutamine and W Tl-201 IV
C2826012|T102|strict|39941-0|LNC|Lung Scan perfusion W particulate radionuclide IV|Lung Scan perfusion W particulate radionuclide IV
C2826012|T102|strict|39833-9|LNC|Lung Scan perfusion W radionuclide gaseous inhaled|Lung Scan perfusion W radionuclide gaseous inhaled
C2826012|T102|strict|39716-6|LNC|Heart Scan perfusion|Heart Scan perfusion
C2826012|T102|strict|39697-8|LNC|Lung Scan perfusion|Lung Scan perfusion
C2826012|T102|strict|39730-7|LNC|Heart Scan perfusion W stress and W radionuclide IV|Heart Scan perfusion W stress and W radionuclide IV
C2826012|T102|strict|39732-3|LNC|Heart Scan perfusion W stress and W Tc-99m Sestamibi IV|Heart Scan perfusion W stress and W Tc-99m Sestamibi IV
C2826012|T102|strict|39715-8|LNC|Heart Scan perfusion W stress and W Tl-201 IV|Heart Scan perfusion W stress and W Tl-201 IV
C2826012|T102|strict|39704-2|LNC|Heart Scan perfusion W Tc-99m Sestamibi IV|Heart Scan perfusion W Tc-99m Sestamibi IV
C2826012|T102|strict|39714-1|LNC|Heart Scan perfusion W Tl-201 IV|Heart Scan perfusion W Tl-201 IV
C2826012|T102|strict|39713-3|LNC|Heart Scan perfusion W Tl-201 IV and Tc-99m Tetrofosmin IV|Heart Scan perfusion W Tl-201 IV and Tc-99m Tetrofosmin IV
C2826012|T102|strict|30765-2|LNC|Acetabulum X-ray portable|Acetabulum X-ray portable
C2826012|T102|strict|30764-5|LNC|Acetabulum - bilateral X-ray portable|Acetabulum - bilateral X-ray portable
C2826012|T102|strict|41823-6|LNC|Ankle - left X-ray portable|Ankle - left X-ray portable
C2826012|T102|strict|41782-4|LNC|Ankle - right X-ray portable|Ankle - right X-ray portable
C2826012|T102|strict|30746-2|LNC|Chest X-ray portable|Chest X-ray portable
C2826012|T102|strict|41827-7|LNC|Elbow - left X-ray portable|Elbow - left X-ray portable
C2826012|T102|strict|41786-5|LNC|Elbow - right X-ray portable|Elbow - right X-ray portable
C2826012|T102|strict|41773-3|LNC|Facial bones X-ray portable|Facial bones X-ray portable
C2826012|T102|strict|41818-6|LNC|Femur - left X-ray portable|Femur - left X-ray portable
C2826012|T102|strict|41778-2|LNC|Femur - right X-ray portable|Femur - right X-ray portable
C2826012|T102|strict|43570-1|LNC|Hand X-ray portable|Hand X-ray portable
C2826012|T102|strict|41829-3|LNC|Hand - left X-ray portable|Hand - left X-ray portable
C2826012|T102|strict|41788-1|LNC|Hand - right X-ray portable|Hand - right X-ray portable
C2826012|T102|strict|37168-2|LNC|Hip X-ray portable|Hip X-ray portable
C2826012|T102|strict|37169-0|LNC|Hip - left X-ray portable|Hip - left X-ray portable
C2826012|T102|strict|38796-9|LNC|Hip - right X-ray portable|Hip - right X-ray portable
C2826012|T102|strict|37170-8|LNC|Humerus X-ray portable|Humerus X-ray portable
C2826012|T102|strict|41825-1|LNC|Humerus - left X-ray portable|Humerus - left X-ray portable
C2826012|T102|strict|41784-0|LNC|Humerus - right X-ray portable|Humerus - right X-ray portable
C2826012|T102|strict|41820-2|LNC|Knee - left X-ray portable|Knee - left X-ray portable
C2826012|T102|strict|41779-0|LNC|Knee - right X-ray portable|Knee - right X-ray portable
C2826012|T102|strict|30792-6|LNC|Patella X-ray portable|Patella X-ray portable
C2826012|T102|strict|30772-8|LNC|Pelvis X-ray portable|Pelvis X-ray portable
C2826012|T102|strict|30747-0|LNC|Ribs X-ray portable|Ribs X-ray portable
C2826012|T102|strict|41831-9|LNC|Ribs - left X-ray portable|Ribs - left X-ray portable
C2826012|T102|strict|41791-5|LNC|Ribs - right X-ray portable|Ribs - right X-ray portable
C2826012|T102|strict|46391-9|LNC|Shoulder X-ray portable|Shoulder X-ray portable
C2826012|T102|strict|41824-4|LNC|Shoulder - left X-ray portable|Shoulder - left X-ray portable
C2826012|T102|strict|41783-2|LNC|Shoulder - right X-ray portable|Shoulder - right X-ray portable
C2826012|T102|strict|30723-1|LNC|Skull X-ray portable|Skull X-ray portable
C2826012|T102|strict|37171-6|LNC|Spine Cervical X-ray portable|Spine Cervical X-ray portable
C2826012|T102|strict|44203-8|LNC|Spine Cervical and Thoracic and Lumbar X-ray portable|Spine Cervical and Thoracic and Lumbar X-ray portable
C2826012|T102|strict|37172-4|LNC|Spine Lumbar X-ray portable|Spine Lumbar X-ray portable
C2826012|T102|strict|41828-5|LNC|Wrist - left X-ray portable|Wrist - left X-ray portable
C2826012|T102|strict|41787-3|LNC|Wrist - right X-ray portable|Wrist - right X-ray portable
C2826012|T102|strict|37151-8|LNC|Unspecified body region Fluoroscopy portable|Unspecified body region Fluoroscopy portable
C2826012|T102|strict|30731-4|LNC|Zygomatic arch X-ray portable|Zygomatic arch X-ray portable
C2826012|T102|strict|30730-6|LNC|Zygomatic arch - bilateral X-ray portable|Zygomatic arch - bilateral X-ray portable
C2826012|T102|strict|24634-8|LNC|Chest X-ray portable W inspiration and expiration|Chest X-ray portable W inspiration and expiration
C2826012|T102|strict|24824-5|LNC|Lung Scan portable|Lung Scan portable
C2826012|T102|strict|42402-8|LNC|Unspecified body region X-ray post mortem|Unspecified body region X-ray post mortem
C2826012|T102|strict|43657-6|LNC|Lung Scan quantitative|Lung Scan quantitative
C2826012|T102|strict|30733-0|LNC|Chest X-ray right and left oblique portable|Chest X-ray right and left oblique portable
C2826012|T102|strict|37131-0|LNC|Abdomen X-ray right lateral and left lateral|Abdomen X-ray right lateral and left lateral
C2826012|T102|strict|37138-5|LNC|Abdomen X-ray right oblique and left oblique|Abdomen X-ray right oblique and left oblique
C2826012|T102|strict|41792-3|LNC|Chest X-ray right oblique and left oblique|Chest X-ray right oblique and left oblique
C2826012|T102|strict|24651-2|LNC|Chest X-ray right oblique and left oblique upright|Chest X-ray right oblique and left oblique upright
C2826012|T102|strict|42414-3|LNC|Chest X-ray right oblique and left oblique W nipple markers|Chest X-ray right oblique and left oblique W nipple markers
C2826012|T102|strict|37016-3|LNC|Breast - bilateral Mammogram roll|Breast - bilateral Mammogram roll
C2826012|T102|strict|37017-1|LNC|Breast - left Mammogram roll|Breast - left Mammogram roll
C2826012|T102|strict|37775-4|LNC|Breast - right Mammogram roll|Breast - right Mammogram roll
C2826012|T102|strict|30740-5|LNC|Chest X-ray right or-left oblique|Chest X-ray right or-left oblique
C2826012|T102|strict|30739-7|LNC|Chest X-ray right or-left oblique portable|Chest X-ray right or-left oblique portable
C2826012|T102|strict|43479-5|LNC|Aorta abdominal Fluoroscopic angiogram runoff W contrast IA|Aorta abdominal Fluoroscopic angiogram runoff W contrast IA
C2826012|T102|strict|30838-7|LNC|Aorta and Femoral artery - bilateral Fluoroscopic angiogram runoff W contrast IA|Aorta and Femoral artery - bilateral Fluoroscopic angiogram runoff W contrast IA
C2826012|T102|strict|37364-7|LNC|Aorta and Femoral artery - left Fluoroscopic angiogram runoff W contrast IA|Aorta and Femoral artery - left Fluoroscopic angiogram runoff W contrast IA
C2826012|T102|strict|38799-3|LNC|Aorta and Femoral artery - right Fluoroscopic angiogram runoff W contrast IA|Aorta and Femoral artery - right Fluoroscopic angiogram runoff W contrast IA
C2826012|T102|strict|38107-9|LNC|Wrist X-ray scaphoid|Wrist X-ray scaphoid
C2826012|T102|strict|37304-3|LNC|Wrist - bilateral X-ray scaphoid|Wrist - bilateral X-ray scaphoid
C2826012|T102|strict|37302-7|LNC|Wrist - left X-ray scaphoid|Wrist - left X-ray scaphoid
C2826012|T102|strict|38115-2|LNC|Wrist - right X-ray scaphoid|Wrist - right X-ray scaphoid
C2826012|T102|strict|24930-0|LNC|Spine Thoracic and Lumbar X-ray scoliosis|Spine Thoracic and Lumbar X-ray scoliosis
C2826012|T102|strict|30715-7|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP and lateral|Spine Thoracic and Lumbar X-ray scoliosis AP and lateral
C2826012|T102|strict|42424-2|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP and lateral sitting|Spine Thoracic and Lumbar X-ray scoliosis AP and lateral sitting
C2826012|T102|strict|39367-8|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP and lateral standing|Spine Thoracic and Lumbar X-ray scoliosis AP and lateral standing
C2826012|T102|strict|42472-1|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP in traction|Spine Thoracic and Lumbar X-ray scoliosis AP in traction
C2826012|T102|strict|42425-9|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP standing and W right bending and W left bending and WO bending|Spine Thoracic and Lumbar X-ray scoliosis AP standing and W right bending and W left bending and WO bending
C2826012|T102|strict|43569-3|LNC|Spine Thoracic and Lumbar X-ray scoliosis AP upright and supine|Spine Thoracic and Lumbar X-ray scoliosis AP upright and supine
C2826012|T102|strict|30716-5|LNC|Spine Thoracic and Lumbar X-ray scoliosis lateral|Spine Thoracic and Lumbar X-ray scoliosis lateral
C2826012|T102|strict|30717-3|LNC|Spine Thoracic and Lumbar X-ray scoliosis standing|Spine Thoracic and Lumbar X-ray scoliosis standing
C2826012|T102|strict|24929-2|LNC|Spine Thoracic and Lumbar X-ray scoliosis W flexion and W extension|Spine Thoracic and Lumbar X-ray scoliosis W flexion and W extension
C2826012|T102|strict|24606-6|LNC|Breast Mammogram screening|Breast Mammogram screening
C2826012|T102|strict|39153-2|LNC|Breast FFD mammogram screening|Breast FFD mammogram screening
C2826012|T102|strict|69159-2|LNC|Breast implant X-ray screening|Breast implant X-ray screening
C2826012|T102|strict|48492-3|LNC|Breast implant - bilateral Mammogram screening|Breast implant - bilateral Mammogram screening
C2826012|T102|strict|26175-0|LNC|Breast - bilateral Mammogram screening|Breast - bilateral Mammogram screening
C2826012|T102|strict|42174-3|LNC|Breast - bilateral FFD mammogram screening|Breast - bilateral FFD mammogram screening
C2826012|T102|strict|26176-8|LNC|Breast - left Mammogram screening|Breast - left Mammogram screening
C2826012|T102|strict|46355-4|LNC|Breast - left FFD mammogram screening|Breast - left FFD mammogram screening
C2826012|T102|strict|26177-6|LNC|Breast - right Mammogram screening|Breast - right Mammogram screening
C2826012|T102|strict|46354-7|LNC|Breast - right FFD mammogram screening|Breast - right FFD mammogram screening
C2826012|T102|strict|46356-2|LNC|Breast - unilateral Mammogram screening|Breast - unilateral Mammogram screening
C2826012|T102|strict|37022-1|LNC|Calcaneus X-ray ski jump|Calcaneus X-ray ski jump
C2826012|T102|strict|37021-3|LNC|Calcaneus - bilateral X-ray ski jump|Calcaneus - bilateral X-ray ski jump
C2826012|T102|strict|37023-9|LNC|Calcaneus - left X-ray ski jump|Calcaneus - left X-ray ski jump
C2826012|T102|strict|38778-7|LNC|Calcaneus - right X-ray ski jump|Calcaneus - right X-ray ski jump
C2826012|T102|strict|37551-9|LNC|Breast Mammogram spot|Breast Mammogram spot
C2826012|T102|strict|37552-7|LNC|Breast - bilateral Mammogram spot|Breast - bilateral Mammogram spot
C2826012|T102|strict|38807-4|LNC|Breast - right Mammogram spot|Breast - right Mammogram spot
C2826012|T102|strict|37553-5|LNC|Breast - left Mammogram spot compression|Breast - left Mammogram spot compression
C2826012|T102|strict|43550-3|LNC|Brain Scan static and flow|Brain Scan static and flow
C2826012|T102|strict|39952-7|LNC|Scrotum and Testicle Scan static and flow|Scrotum and Testicle Scan static and flow
C2826012|T102|strict|39676-2|LNC|Scan static for infection W GA-67 IV|Scan static for infection W GA-67 IV
C2826012|T102|strict|39894-1|LNC|Heart Scan static for shunt detection|Heart Scan static for shunt detection
C2826012|T102|strict|39896-6|LNC|Scan static for tumor W GA-67 IV|Scan static for tumor W GA-67 IV
C2826012|T102|strict|39814-9|LNC|Bone Scan static limited|Bone Scan static limited
C2826012|T102|strict|39634-1|LNC|Brain Scan static limited|Brain Scan static limited
C2826012|T102|strict|39903-0|LNC|Bone Scan static multiple areas|Bone Scan static multiple areas
C2826012|T102|strict|39817-2|LNC|Bone Scan static whole body|Bone Scan static whole body
C2826012|T102|strict|39815-6|LNC|Bone Scan static|Bone Scan static
C2826012|T102|strict|39824-8|LNC|Bone marrow Scan static|Bone marrow Scan static
C2826012|T102|strict|39633-3|LNC|Brain Scan static|Brain Scan static
C2826012|T102|strict|39853-7|LNC|Kidney - bilateral Scan static|Kidney - bilateral Scan static
C2826012|T102|strict|39832-1|LNC|Liver Scan static|Liver Scan static
C2826012|T102|strict|39878-4|LNC|Liver and Spleen Scan static|Liver and Spleen Scan static
C2826012|T102|strict|39900-6|LNC|Salivary gland Scan static|Salivary gland Scan static
C2826012|T102|strict|39855-2|LNC|Scrotum and Testicle Scan static|Scrotum and Testicle Scan static
C2826012|T102|strict|43501-6|LNC|Vessel Scan static|Vessel Scan static
C2826012|T102|strict|44150-1|LNC|Brain Scan static W Tc-99m bicisate IV|Brain Scan static W Tc-99m bicisate IV
C2826012|T102|strict|39854-5|LNC|Kidney - bilateral Scan static W Tc-99m DMSA IV|Kidney - bilateral Scan static W Tc-99m DMSA IV
C2826012|T102|strict|37153-4|LNC|Mastoid X-ray Stenver and Arcelin|Mastoid X-ray Stenver and Arcelin
C2826012|T102|strict|69136-0|LNC|Knee X-ray Sunrise and tunnel|Knee X-ray Sunrise and tunnel
C2826012|T102|strict|37163-3|LNC|Knee - bilateral X-ray Sunrise and tunnel|Knee - bilateral X-ray Sunrise and tunnel
C2826012|T102|strict|37156-7|LNC|Knee - left X-ray Sunrise and tunnel|Knee - left X-ray Sunrise and tunnel
C2826012|T102|strict|37759-8|LNC|Knee - right X-ray Sunrise and tunnel|Knee - right X-ray Sunrise and tunnel
C2826012|T102|strict|39345-4|LNC|Knee - left X-ray Sunrise and tunnel standing|Knee - left X-ray Sunrise and tunnel standing
C2826012|T102|strict|69255-8|LNC|Knee - right X-ray Sunrise and tunnel standing|Knee - right X-ray Sunrise and tunnel standing
C2826012|T102|strict|38088-1|LNC|Knee - bilateral X-ray Sunrise 20 and 40 and 60 degrees|Knee - bilateral X-ray Sunrise 20 and 40 and 60 degrees
C2826012|T102|strict|38087-3|LNC|Knee - left X-ray Sunrise 20 and 40 and 60 degrees|Knee - left X-ray Sunrise 20 and 40 and 60 degrees
C2826012|T102|strict|38824-9|LNC|Knee - right X-ray Sunrise 20 and 40 and 60 degrees|Knee - right X-ray Sunrise 20 and 40 and 60 degrees
C2826012|T102|strict|24579-5|LNC|Bones long X-ray survey|Bones long X-ray survey
C2826012|T102|strict|43518-0|LNC|Bones X-ray survey|Bones X-ray survey
C2826012|T102|strict|37365-4|LNC|Bones X-ray survey for metastasis|Bones X-ray survey for metastasis
C2826012|T102|strict|39518-6|LNC|Bones long X-ray survey limited|Bones long X-ray survey limited
C2826012|T102|strict|43519-8|LNC|Bones X-ray survey limited|Bones X-ray survey limited
C2826012|T102|strict|38089-9|LNC|Bones X-ray survey limited for metastasis|Bones X-ray survey limited for metastasis
C2826012|T102|strict|37159-1|LNC|Foot - left X-ray tarsal|Foot - left X-ray tarsal
C2826012|T102|strict|38792-8|LNC|Foot - right X-ray tarsal|Foot - right X-ray tarsal
C2826012|T102|strict|43796-2|LNC|Wrist - bilateral X-ray tunnel.carpal|Wrist - bilateral X-ray tunnel.carpal
C2826012|T102|strict|69304-4|LNC|Wrist X-ray ulnar deviation|Wrist X-ray ulnar deviation
C2826012|T102|strict|69303-6|LNC|Wrist X-ray ulnar deviation and radial deviation|Wrist X-ray ulnar deviation and radial deviation
C2826012|T102|strict|69072-7|LNC|Wrist - bilateral X-ray ulnar deviation and radial deviation|Wrist - bilateral X-ray ulnar deviation and radial deviation
C2826012|T102|strict|37555-0|LNC|Wrist - left X-ray ulnar deviation and radial deviation|Wrist - left X-ray ulnar deviation and radial deviation
C2826012|T102|strict|38808-2|LNC|Wrist - right X-ray ulnar deviation and radial deviation|Wrist - right X-ray ulnar deviation and radial deviation
C2826012|T102|strict|43532-1|LNC|Chest and Abdomen X-ray upright and PA chest|Chest and Abdomen X-ray upright and PA chest
C2826012|T102|strict|39944-4|LNC|Lung Scan ventilation and equilibrium and washout W radionuclide inhaled|Lung Scan ventilation and equilibrium and washout W radionuclide inhaled
C2826012|T102|strict|39948-5|LNC|Lung Scan ventilation and equilibrium and washout W radionuclide inhaled single breath|Lung Scan ventilation and equilibrium and washout W radionuclide inhaled single breath
C2826012|T102|strict|39947-7|LNC|Lung Scan ventilation and equilibrium W radionuclide inhaled single breath|Lung Scan ventilation and equilibrium W radionuclide inhaled single breath
C2826012|T102|strict|39946-9|LNC|Lung Scan ventilation and perfusion and differential W radionuclide inhaled and W radionuclide IV|Lung Scan ventilation and perfusion and differential W radionuclide inhaled and W radionuclide IV
C2826012|T102|strict|39943-6|LNC|Lung Scan ventilation and perfusion W radionuclide inhaled and W particulate radionuclide IV|Lung Scan ventilation and perfusion W radionuclide inhaled and W particulate radionuclide IV
C2826012|T102|strict|30697-7|LNC|Pulmonary system Scan ventilation and perfusion W radionuclide inhaled and W radionuclide IV|Pulmonary system Scan ventilation and perfusion W radionuclide inhaled and W radionuclide IV
C2826012|T102|strict|39942-8|LNC|Lung Scan ventilation and perfusion W radionuclide inhaled single breath and W particulate radionuclide IV|Lung Scan ventilation and perfusion W radionuclide inhaled single breath and W particulate radionuclide IV
C2826012|T102|strict|24888-0|LNC|Pulmonary system Scan ventilation and perfusion W Xe-133 inhaled and W Tc-99m MAA IV|Pulmonary system Scan ventilation and perfusion W Xe-133 inhaled and W Tc-99m MAA IV
C2826012|T102|strict|39835-4|LNC|Lung Scan ventilation W radionuclide aerosol inhaled|Lung Scan ventilation W radionuclide aerosol inhaled
C2826012|T102|strict|39836-2|LNC|Lung Scan ventilation W radionuclide gaseous inhaled|Lung Scan ventilation W radionuclide gaseous inhaled
C2826012|T102|strict|39945-1|LNC|Lung Scan ventilation W radionuclide gaseous inhaled single breath|Lung Scan ventilation W radionuclide gaseous inhaled single breath
C2826012|T102|strict|39837-0|LNC|Lung Scan ventilation W radionuclide inhaled|Lung Scan ventilation W radionuclide inhaled
C2826012|T102|strict|39834-7|LNC|Lung Scan ventilation W Tc-99m DTPA aerosol inhaled|Lung Scan ventilation W Tc-99m DTPA aerosol inhaled
C2826012|T102|strict|46361-2|LNC|Lung Scan ventilation W Xe-133 inhaled|Lung Scan ventilation W Xe-133 inhaled
C2826012|T102|strict|39932-9|LNC|Heart Scan wall motion and ejection fraction|Heart Scan wall motion and ejection fraction
C2826012|T102|strict|39873-5|LNC|Heart Scan wall motion|Heart Scan wall motion
C2826012|T102|strict|39683-8|LNC|Scan whole body W GA-67 IV|Scan whole body W GA-67 IV
C2826012|T102|strict|39698-6|LNC|Scan whole body W I-131 MIBG IV|Scan whole body W I-131 MIBG IV
C2826012|T102|strict|39845-3|LNC|Scan whole body W In-111 Satumomab IV|Scan whole body W In-111 Satumomab IV
C2826012|T102|strict|42711-2|LNC|Scan whole body W In-111 tagged WBC IV|Scan whole body W In-111 tagged WBC IV
C2826012|T102|strict|42175-0|LNC|Scan whole body|Scan whole body
C2826012|T102|strict|39818-0|LNC|Bone Scan whole body|Bone Scan whole body
C2826012|T102|strict|39826-3|LNC|Bone marrow Scan whole body|Bone marrow Scan whole body
C2826012|T102|strict|39669-7|LNC|Scan whole body W Tc-99m Arcitumomab IV|Scan whole body W Tc-99m Arcitumomab IV
C2826012|T102|strict|24713-0|LNC|Gallbladder X-ray 48 hours post contrast PO|Gallbladder X-ray 48 hours post contrast PO
C2826012|T102|strict|39660-6|LNC|Heart Scan at rest and W dipyridamole and W radionuclide IV|Heart Scan at rest and W dipyridamole and W radionuclide IV
C2826012|T102|strict|39661-4|LNC|Heart Scan at rest and W dobutamine and W radionuclide IV|Heart Scan at rest and W dobutamine and W radionuclide IV
C2826012|T102|strict|39663-0|LNC|Heart Scan at rest and W stress and W radionuclide IV|Heart Scan at rest and W stress and W radionuclide IV
C2826012|T102|strict|42309-5|LNC|Heart Scan at rest and W stress and W Tl-201 IV|Heart Scan at rest and W stress and W Tl-201 IV
C2826012|T102|strict|24750-2|LNC|Heart Scan at rest and W Tl-201 IV|Heart Scan at rest and W Tl-201 IV
C2826012|T102|strict|43459-7|LNC|Brain Scan during electroconvulsive shock treatment|Brain Scan during electroconvulsive shock treatment
C2826012|T102|strict|24577-9|LNC|Bone X-ray during surgery|Bone X-ray during surgery
C2826012|T102|strict|47372-8|LNC|Hip X-ray during surgery|Hip X-ray during surgery
C2826012|T102|strict|25070-4|LNC|Unspecified body region Fluoroscopy during surgery|Unspecified body region Fluoroscopy during surgery
C2826012|T102|strict|24574-6|LNC|Biliary ducts and Gallbladder Fluoroscopy during surgery W contrast biliary duct|Biliary ducts and Gallbladder Fluoroscopy during surgery W contrast biliary duct
C2826012|T102|strict|46352-1|LNC|Breast duct Mammogram during surgery W contrast intra duct|Breast duct Mammogram during surgery W contrast intra duct
C2826012|T102|strict|43485-2|LNC|Kidney X-ray during surgery W contrast retrograde|Kidney X-ray during surgery W contrast retrograde
C2826012|T102|strict|39150-8|LNC|Breast FFD mammogram Post Localization|Breast FFD mammogram Post Localization
C2826012|T102|strict|69251-7|LNC|Breast Mammogram Post Wire Placement|Breast Mammogram Post Wire Placement
C2826012|T102|strict|42415-0|LNC|Breast - bilateral Mammogram Post Wire Placement|Breast - bilateral Mammogram Post Wire Placement
C2826012|T102|strict|42416-8|LNC|Breast - left Mammogram Post Wire Placement|Breast - left Mammogram Post Wire Placement
C2826012|T102|strict|37201-1|LNC|Ankle X-ray standing|Ankle X-ray standing
C2826012|T102|strict|37202-9|LNC|Ankle - bilateral X-ray standing|Ankle - bilateral X-ray standing
C2826012|T102|strict|37203-7|LNC|Ankle - left X-ray standing|Ankle - left X-ray standing
C2826012|T102|strict|37676-4|LNC|Ankle - right X-ray standing|Ankle - right X-ray standing
C2826012|T102|strict|37205-2|LNC|Calcaneus X-ray standing|Calcaneus X-ray standing
C2826012|T102|strict|37206-0|LNC|Calcaneus - left X-ray standing|Calcaneus - left X-ray standing
C2826012|T102|strict|37720-0|LNC|Calcaneus - right X-ray standing|Calcaneus - right X-ray standing
C2826012|T102|strict|38845-4|LNC|Femur - left X-ray standing|Femur - left X-ray standing
C2826012|T102|strict|37693-9|LNC|Femur - right X-ray standing|Femur - right X-ray standing
C2826012|T102|strict|24708-0|LNC|Foot X-ray standing|Foot X-ray standing
C2826012|T102|strict|26094-3|LNC|Foot - bilateral X-ray standing|Foot - bilateral X-ray standing
C2826012|T102|strict|26095-0|LNC|Foot - left X-ray standing|Foot - left X-ray standing
C2826012|T102|strict|26096-8|LNC|Foot - right X-ray standing|Foot - right X-ray standing
C2826012|T102|strict|37584-0|LNC|Great toe - left X-ray standing|Great toe - left X-ray standing
C2826012|T102|strict|38810-8|LNC|Great toe - right X-ray standing|Great toe - right X-ray standing
C2826012|T102|strict|24809-6|LNC|Knee X-ray standing|Knee X-ray standing
C2826012|T102|strict|26085-1|LNC|Knee - bilateral X-ray standing|Knee - bilateral X-ray standing
C2826012|T102|strict|26086-9|LNC|Knee - left X-ray standing|Knee - left X-ray standing
C2826012|T102|strict|26087-7|LNC|Knee - right X-ray standing|Knee - right X-ray standing
C2826012|T102|strict|37204-5|LNC|Lower extremity X-ray standing|Lower extremity X-ray standing
C2826012|T102|strict|69264-0|LNC|Sacrum X-ray standing|Sacrum X-ray standing
C2826012|T102|strict|37208-6|LNC|Spine Lumbar X-ray standing|Spine Lumbar X-ray standing
C2826012|T102|strict|69275-6|LNC|Spine Thoracic X-ray standing|Spine Thoracic X-ray standing
C2826012|T102|strict|38124-4|LNC|Spine Thoracic and Lumbar X-ray standing|Spine Thoracic and Lumbar X-ray standing
C2826012|T102|strict|37899-2|LNC|Tibia and Fibula X-ray standing|Tibia and Fibula X-ray standing
C2826012|T102|strict|37209-4|LNC|Toes - left X-ray standing|Toes - left X-ray standing
C2826012|T102|strict|37823-2|LNC|Toes - right X-ray standing|Toes - right X-ray standing
C2826012|T102|strict|44233-5|LNC|Kidney - bilateral Scan W and WO Tc-99m DTPA IV|Kidney - bilateral Scan W and WO Tc-99m DTPA IV
C2826012|T102|strict|44232-7|LNC|Kidney - bilateral Scan W and WO Tc-99m Mertiatide IV|Kidney - bilateral Scan W and WO Tc-99m Mertiatide IV
C2826012|T102|strict|37579-0|LNC|Acromioclavicular Joint X-ray W and WO weight|Acromioclavicular Joint X-ray W and WO weight
C2826012|T102|strict|37580-8|LNC|Acromioclavicular joint - bilateral X-ray W and WO weight|Acromioclavicular joint - bilateral X-ray W and WO weight
C2826012|T102|strict|37581-6|LNC|Acromioclavicular joint - left X-ray W and WO weight|Acromioclavicular joint - left X-ray W and WO weight
C2826012|T102|strict|37663-2|LNC|Acromioclavicular joint - right X-ray W and WO weight|Acromioclavicular joint - right X-ray W and WO weight
C2826012|T102|strict|39651-5|LNC|Heart Scan W adenosine and W Tl-201 IV|Heart Scan W adenosine and W Tl-201 IV
C2826012|T102|strict|38090-7|LNC|Breast - bilateral Mammogram W air|Breast - bilateral Mammogram W air
C2826012|T102|strict|38091-5|LNC|Breast - left Mammogram W air|Breast - left Mammogram W air
C2826012|T102|strict|39059-1|LNC|Gastrointestine upper Fluoroscopy W air and barium contrast PO|Gastrointestine upper Fluoroscopy W air and barium contrast PO
C2826012|T102|strict|24666-0|LNC|Colon Fluoroscopy W air and barium contrast PR|Colon Fluoroscopy W air and barium contrast PR
C2826012|T102|strict|46357-0|LNC|Colon Fluoroscopy W air contrast PR|Colon Fluoroscopy W air contrast PR
C2826012|T102|strict|30633-2|LNC|Esophagus Fluoroscopy W barium contrast PO|Esophagus Fluoroscopy W barium contrast PO
C2826012|T102|strict|42683-3|LNC|Gastrointestine upper Fluoroscopy W barium contrast PO|Gastrointestine upper Fluoroscopy W barium contrast PO
C2826012|T102|strict|43574-3|LNC|Upper Gastrointestine and Small bowel Fluoroscopy W barium contrast PO|Upper Gastrointestine and Small bowel Fluoroscopy W barium contrast PO
C2826012|T102|strict|44227-7|LNC|Colon Fluoroscopy W barium contrast PR|Colon Fluoroscopy W barium contrast PR
C2826012|T102|strict|37565-9|LNC|Unspecified body region Fluoroscopy W barium contrast via fistula|Unspecified body region Fluoroscopy W barium contrast via fistula
C2826012|T102|strict|38092-3|LNC|Urinary bladder Fluoroscopy W chain and contrast intra bladder|Urinary bladder Fluoroscopy W chain and contrast intra bladder
C2826012|T102|strict|41770-9|LNC|Gallbladder Scan W cholecystokinin and W radionuclide IV|Gallbladder Scan W cholecystokinin and W radionuclide IV
C2826012|T102|strict|43650-1|LNC|Liver and Biliary ducts and Gallbladder Scan W cholecystokinin and W radionuclide IV|Liver and Biliary ducts and Gallbladder Scan W cholecystokinin and W radionuclide IV
C2826012|T102|strict|30630-8|LNC|Head Cistern Fluoroscopy video W contrast|Head Cistern Fluoroscopy video W contrast
C2826012|T102|strict|30824-7|LNC|Intercranial vessel and Neck Vessel Fluoroscopic angiogram W contrast|Intercranial vessel and Neck Vessel Fluoroscopic angiogram W contrast
C2826012|T102|strict|37585-7|LNC|Jejunum Fluoroscopy W contrast|Jejunum Fluoroscopy W contrast
C2826012|T102|strict|38853-8|LNC|Lower extremity vessels - left Fluoroscopic angiogram W contrast|Lower extremity vessels - left Fluoroscopic angiogram W contrast
C2826012|T102|strict|37765-5|LNC|Lower extremity vessels - right Fluoroscopic angiogram W contrast|Lower extremity vessels - right Fluoroscopic angiogram W contrast
C2826012|T102|strict|37615-2|LNC|Pelvis vessels Fluoroscopic angiogram W contrast|Pelvis vessels Fluoroscopic angiogram W contrast
C2826012|T102|strict|37936-2|LNC|Peripheral vessels Fluoroscopic angiogram W contrast|Peripheral vessels Fluoroscopic angiogram W contrast
C2826012|T102|strict|37640-0|LNC|Renal vessels Fluoroscopic angiogram W contrast|Renal vessels Fluoroscopic angiogram W contrast
C2826012|T102|strict|64140-7|LNC|Renal vessels - left Fluoroscopic angiogram W contrast|Renal vessels - left Fluoroscopic angiogram W contrast
C2826012|T102|strict|64141-5|LNC|Renal vessels - right Fluoroscopic angiogram W contrast|Renal vessels - right Fluoroscopic angiogram W contrast
C2826012|T102|strict|38094-9|LNC|Spine.cavity Fluoroscopy W contrast|Spine.cavity Fluoroscopy W contrast
C2826012|T102|strict|37973-5|LNC|Testicle vessels Fluoroscopy W contrast|Testicle vessels Fluoroscopy W contrast
C2826012|T102|strict|25005-0|LNC|Three vessels Fluoroscopic angiogram W contrast|Three vessels Fluoroscopic angiogram W contrast
C2826012|T102|strict|25014-2|LNC|Two vessels Fluoroscopic angiogram W contrast|Two vessels Fluoroscopic angiogram W contrast
C2826012|T102|strict|37976-8|LNC|Upper extremity vessels Fluoroscopic angiogram W contrast|Upper extremity vessels Fluoroscopic angiogram W contrast
C2826012|T102|strict|42014-1|LNC|Urinary Bladder and Urethra Fluoroscopy W contrast|Urinary Bladder and Urethra Fluoroscopy W contrast
C2826012|T102|strict|37980-0|LNC|Vertebral vessels Fluoroscopic angiogram W contrast|Vertebral vessels Fluoroscopic angiogram W contrast
C2826012|T102|strict|37981-8|LNC|Visceral vessels Fluoroscopic angiogram W contrast|Visceral vessels Fluoroscopic angiogram W contrast
C2826012|T102|strict|37575-8|LNC|Gallbladder X-ray W contrast and fatty meal PO|Gallbladder X-ray W contrast and fatty meal PO
C2826012|T102|strict|38101-2|LNC|Kidney X-ray W contrast antegrade|Kidney X-ray W contrast antegrade
C2826012|T102|strict|46376-0|LNC|Kidney - bilateral Fluoroscopy W contrast antegrade|Kidney - bilateral Fluoroscopy W contrast antegrade
C2826012|T102|strict|38100-4|LNC|Urinary Bladder and Urethra Fluoroscopy W contrast antegrade|Urinary Bladder and Urethra Fluoroscopy W contrast antegrade
C2826012|T102|strict|38102-0|LNC|Kidney X-ray W contrast antegrade via pyelostomy|Kidney X-ray W contrast antegrade via pyelostomy
C2826012|T102|strict|25030-8|LNC|Abdominal Arteries Fluoroscopic angiogram W contrast IA|Abdominal Arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30832-0|LNC|Adrenal artery Fluoroscopic angiogram W contrast IA|Adrenal artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30831-2|LNC|Adrenal artery - bilateral Fluoroscopic angiogram W contrast IA|Adrenal artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37387-8|LNC|Adrenal artery - left Fluoroscopic angiogram W contrast IA|Adrenal artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37939-6|LNC|Adrenal artery - right Fluoroscopic angiogram W contrast IA|Adrenal artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|38861-1|LNC|Ankle arteries - left Fluoroscopic angiogram W contrast IA|Ankle arteries - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37941-2|LNC|Ankle arteries - right Fluoroscopic angiogram W contrast IA|Ankle arteries - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24658-7|LNC|Aorta Fluoroscopic angiogram W contrast IA|Aorta Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30837-9|LNC|Aorta abdominal Fluoroscopic angiogram W contrast IA|Aorta abdominal Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24546-4|LNC|Aorta arch and Neck Fluoroscopic angiogram W contrast IA|Aorta arch and Neck Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37366-2|LNC|Abdominal Aorta and Arteries Fluoroscopic angiogram W contrast IA|Abdominal Aorta and Arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|69054-5|LNC|Aortic arch Fluoroscopic angiogram W contrast IA|Aortic arch Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37380-3|LNC|Aortic arch and Brachial artery Fluoroscopic angiogram W contrast IA|Aortic arch and Brachial artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37381-1|LNC|Aortic arch and Carotid artery Fluoroscopic angiogram W contrast IA|Aortic arch and Carotid artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37587-3|LNC|Aortic arch and Carotid artery - bilateral and Vertebral artery - bilateral Fluoroscopic angiogram W contrast IA|Aortic arch and Carotid artery - bilateral and Vertebral artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37588-1|LNC|Aortic arch and Carotid artery.common - bilateral Fluoroscopic angiogram W contrast IA|Aortic arch and Carotid artery.common - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37589-9|LNC|Aortic arch and Carotid artery.common - left Fluoroscopic angiogram W contrast IA|Aortic arch and Carotid artery.common - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37590-7|LNC|Aortic arch and Carotid artery.common - right Fluoroscopic angiogram W contrast IA|Aortic arch and Carotid artery.common - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37591-5|LNC|Aortic arch and Carotid artery.external - bilateral Fluoroscopic angiogram W contrast IA|Aortic arch and Carotid artery.external - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37592-3|LNC|Aortic arch and Carotid artery.external - left Fluoroscopic angiogram W contrast IA|Aortic arch and Carotid artery.external - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37593-1|LNC|Aortic arch and Carotid artery.external - right Fluoroscopic angiogram W contrast IA|Aortic arch and Carotid artery.external - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37594-9|LNC|Aortic arch and Carotid artery and Vertebral artery Fluoroscopic angiogram W contrast IA|Aortic arch and Carotid artery and Vertebral artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37382-9|LNC|Aortic arch and Subclavian artery Fluoroscopic angiogram W contrast IA|Aortic arch and Subclavian artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37383-7|LNC|Aortic arch and Subclavian artery - left Fluoroscopic angiogram W contrast IA|Aortic arch and Subclavian artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|38800-9|LNC|Aortic arch and Subclavian artery - right Fluoroscopic angiogram W contrast IA|Aortic arch and Subclavian artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37379-5|LNC|Aortic arch and Upper Extremity artery Fluoroscopic angiogram W contrast IA|Aortic arch and Upper Extremity artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37384-5|LNC|Aortic arch and Vertebral artery Fluoroscopic angiogram W contrast IA|Aortic arch and Vertebral artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37385-2|LNC|Aortic arch and Vertebral artery - left Fluoroscopic angiogram W contrast IA|Aortic arch and Vertebral artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37386-0|LNC|Aortic arch and Vertebral artery - right Fluoroscopic angiogram W contrast IA|Aortic arch and Vertebral artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24551-4|LNC|AV fistula Fluoroscopic angiogram W contrast IA|AV fistula Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30828-8|LNC|Brachial artery Fluoroscopic angiogram W contrast IA|Brachial artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37388-6|LNC|Brachial artery - bilateral Fluoroscopic angiogram W contrast IA|Brachial artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24581-1|LNC|Brachial artery and Subclavian artery Fluoroscopic angiogram W contrast IA|Brachial artery and Subclavian artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|69077-6|LNC|Brachiocephalic artery Fluoroscopic angiogram W contrast IA|Brachiocephalic artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37389-4|LNC|Bronchial artery Fluoroscopic angiogram W contrast IA|Bronchial artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24617-3|LNC|Carotid artery Fluoroscopic angiogram W contrast IA|Carotid artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|26079-4|LNC|Carotid artery - bilateral Fluoroscopic angiogram W contrast IA|Carotid artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|39097-1|LNC|Carotid artery - bilateral and Cerebral artery - bilateral Fluoroscopic angiogram W contrast IA|Carotid artery - bilateral and Cerebral artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|39094-8|LNC|Carotid artery.cervical Fluoroscopic angiogram W contrast IA|Carotid artery.cervical Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|39098-9|LNC|Carotid artery.cervical - bilateral Fluoroscopic angiogram W contrast IA|Carotid artery.cervical - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|38863-7|LNC|Carotid artery.cervical - left Fluoroscopic angiogram W contrast IA|Carotid artery.cervical - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37945-3|LNC|Carotid artery.cervical - right Fluoroscopic angiogram W contrast IA|Carotid artery.cervical - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30821-3|LNC|Carotid artery.external Fluoroscopic angiogram W contrast IA|Carotid artery.external Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30820-5|LNC|Carotid artery.external - bilateral Fluoroscopic angiogram W contrast IA|Carotid artery.external - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37390-2|LNC|Carotid artery.external - left Fluoroscopic angiogram W contrast IA|Carotid artery.external - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37948-7|LNC|Carotid artery.external - right Fluoroscopic angiogram W contrast IA|Carotid artery.external - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|38864-5|LNC|Carotid artery.internal - left Fluoroscopic angiogram W contrast IA|Carotid artery.internal - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37952-9|LNC|Carotid artery.internal - right Fluoroscopic angiogram W contrast IA|Carotid artery.internal - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|26080-2|LNC|Carotid artery - left Fluoroscopic angiogram W contrast IA|Carotid artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|26081-0|LNC|Carotid artery - right Fluoroscopic angiogram W contrast IA|Carotid artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|39095-5|LNC|Carotid artery and Cerebral artery Fluoroscopic angiogram W contrast IA|Carotid artery and Cerebral artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|38865-2|LNC|Carotid artery and Cerebral artery internal - left Fluoroscopic angiogram W contrast IA|Carotid artery and Cerebral artery internal - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37953-7|LNC|Carotid artery and Cerebral artery internal - right Fluoroscopic angiogram W contrast IA|Carotid artery and Cerebral artery internal - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|38862-9|LNC|Carotid artery and Cerebral artery - left Fluoroscopic angiogram W contrast IA|Carotid artery and Cerebral artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37944-6|LNC|Carotid artery and Cerebral artery - right Fluoroscopic angiogram W contrast IA|Carotid artery and Cerebral artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37391-0|LNC|Carotid artery and Vertebral artery Fluoroscopic angiogram W contrast IA|Carotid artery and Vertebral artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37392-8|LNC|Carotid artery and Vertebral artery - bilateral Fluoroscopic angiogram W contrast IA|Carotid artery and Vertebral artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37393-6|LNC|Carotid artery+Vertebral artery - left Fluoroscopic angiogram W contrast IA|Carotid artery+Vertebral artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37943-8|LNC|Carotid artery+Vertebral artery - right Fluoroscopic angiogram W contrast IA|Carotid artery+Vertebral artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24622-3|LNC|Celiac artery Fluoroscopic angiogram W contrast IA|Celiac artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37403-3|LNC|Celiac artery and Gastric artery - left and Superior mesenteric artery Fluoroscopic angiogram W contrast IA|Celiac artery and Gastric artery - left and Superior mesenteric artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37394-4|LNC|Celiac artery and Superior mesenteric artery and Inferior mesenteric artery Fluoroscopic angiogram W contrast IA|Celiac artery and Superior mesenteric artery and Inferior mesenteric artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37173-2|LNC|Cerebral artery Fluoroscopic angiogram W contrast IA|Cerebral artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30891-6|LNC|Cervicocerebral artery Fluoroscopic angiogram W contrast IA|Cervicocerebral artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37174-0|LNC|Coronary arteries Fluoroscopic angiogram W contrast IA|Coronary arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37595-6|LNC|Coronary graft Fluoroscopic angiogram W contrast IA|Coronary graft Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30848-6|LNC|Extremity arteries Fluoroscopic angiogram W contrast IA|Extremity arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30849-4|LNC|Extremity arteries - bilateral Fluoroscopic angiogram W contrast IA|Extremity arteries - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37395-1|LNC|Extremity arteries - left Fluoroscopic angiogram W contrast IA|Extremity arteries - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37949-5|LNC|Extremity arteries - right Fluoroscopic angiogram W contrast IA|Extremity arteries - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37175-7|LNC|Femoral artery Fluoroscopic angiogram W contrast IA|Femoral artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37176-5|LNC|Femoral artery and Popliteal artery Fluoroscopic angiogram W contrast IA|Femoral artery and Popliteal artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37397-7|LNC|Gastric artery Fluoroscopic angiogram W contrast IA|Gastric artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37398-5|LNC|Gastric artery - left Fluoroscopic angiogram W contrast IA|Gastric artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|38801-7|LNC|Gastric artery - right Fluoroscopic angiogram W contrast IA|Gastric artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37399-3|LNC|Gastroduodenal artery Fluoroscopic angiogram W contrast IA|Gastroduodenal artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30822-1|LNC|Head artery - bilateral and Neck artery - bilateral Fluoroscopic angiogram W contrast IA|Head artery - bilateral and Neck artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|62448-6|LNC|Head artery.left+Neck artery.left Fluoroscopic angiogram W contrast IA|Head artery.left+Neck artery.left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|62449-4|LNC|Head artery.right+Neck artery.right Fluoroscopic angiogram W contrast IA|Head artery.right+Neck artery.right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30823-9|LNC|Head artery and Neck artery Fluoroscopic angiogram W contrast IA|Head artery and Neck artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|25076-1|LNC|Hepatic artery Fluoroscopic angiogram W contrast IA|Hepatic artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|43782-2|LNC|Iliac artery Fluoroscopic angiogram W contrast IA|Iliac artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37177-3|LNC|Iliac artery - bilateral Fluoroscopic angiogram W contrast IA|Iliac artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24862-5|LNC|Iliac artery Internal Fluoroscopic angiogram W contrast IA|Iliac artery Internal Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37178-1|LNC|Iliac artery - left Fluoroscopic angiogram W contrast IA|Iliac artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37739-0|LNC|Iliac artery - right Fluoroscopic angiogram W contrast IA|Iliac artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37179-9|LNC|Inferior mesenteric artery Fluoroscopic angiogram W contrast IA|Inferior mesenteric artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|25079-5|LNC|Kidney arteries Fluoroscopic angiogram W contrast IA|Kidney arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37487-6|LNC|Lower extremity arteries Fluoroscopic angiogram W contrast IA|Lower extremity arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|47986-5|LNC|Lower extremity arteries - left Fluoroscopic angiogram W contrast IA|Lower extremity arteries - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|47987-3|LNC|Lower extremity arteries - right Fluoroscopic angiogram W contrast IA|Lower extremity arteries - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30829-6|LNC|Internal mammary artery Fluoroscopic angiogram W contrast IA|Internal mammary artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|64995-4|LNC|Mammary artery.internal - left Fluoroscopic angiogram W contrast IA|Mammary artery.internal - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|65000-2|LNC|Mammary artery.internal - right Fluoroscopic angiogram W contrast IA|Mammary artery.internal - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37401-7|LNC|Maxillary artery.internal Fluoroscopic angiogram W contrast IA|Maxillary artery.internal Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24833-6|LNC|Mesenteric artery Fluoroscopic angiogram W contrast IA|Mesenteric artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24860-9|LNC|Pancreatic artery Fluoroscopic angiogram W contrast IA|Pancreatic artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30833-8|LNC|Pelvis arteries Fluoroscopic angiogram W contrast IA|Pelvis arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37935-4|LNC|Pelvis arteries and Lower extremity arteries - bilateral Fluoroscopic angiogram W contrast IA|Pelvis arteries and Lower extremity arteries - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24874-0|LNC|Peripheral arteries Fluoroscopic angiogram W contrast IA|Peripheral arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|44240-0|LNC|Peripheral arteries - bilateral Fluoroscopic angiogram W contrast IA|Peripheral arteries - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|69249-1|LNC|Popliteal artery Fluoroscopic angiogram W contrast IA|Popliteal artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37181-5|LNC|Popliteal artery - left Fluoroscopic angiogram W contrast IA|Popliteal artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37778-8|LNC|Popliteal artery - right Fluoroscopic angiogram W contrast IA|Popliteal artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37404-1|LNC|Pudendal artery.internal Fluoroscopic angiogram W contrast IA|Pudendal artery.internal Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|39057-5|LNC|Pulmonary artery Fluoroscopic angiogram W contrast IA|Pulmonary artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30830-4|LNC|Pulmonary artery - bilateral Fluoroscopic angiogram W contrast IA|Pulmonary artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37182-3|LNC|Pulmonary artery - left Fluoroscopic angiogram W contrast IA|Pulmonary artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37779-6|LNC|Pulmonary artery - right Fluoroscopic angiogram W contrast IA|Pulmonary artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|30834-6|LNC|Renal artery - bilateral Fluoroscopic angiogram W contrast IA|Renal artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|62446-0|LNC|Renal artery - left Fluoroscopic angiogram W contrast IA|Renal artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|62447-8|LNC|Renal artery - right Fluoroscopic angiogram W contrast IA|Renal artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24925-0|LNC|Spinal artery Fluoroscopic angiogram W contrast IA|Spinal artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|26082-8|LNC|Spinal artery - bilateral Fluoroscopic angiogram W contrast IA|Spinal artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|26083-6|LNC|Spinal artery - left Fluoroscopic angiogram W contrast IA|Spinal artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|26084-4|LNC|Spinal artery - right Fluoroscopic angiogram W contrast IA|Spinal artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24992-0|LNC|Splenic artery Fluoroscopic angiogram W contrast IA|Splenic artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24991-2|LNC|Splenic vein and Portal vein Fluoroscopic angiogram W contrast IA|Splenic vein and Portal vein Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37886-9|LNC|Subclavian artery Fluoroscopic angiogram W contrast IA|Subclavian artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37405-8|LNC|Subclavian artery - bilateral Fluoroscopic angiogram W contrast IA|Subclavian artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37406-6|LNC|Subclavian artery - left Fluoroscopic angiogram W contrast IA|Subclavian artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37966-9|LNC|Subclavian artery - right Fluoroscopic angiogram W contrast IA|Subclavian artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37180-7|LNC|Superior mesenteric artery Fluoroscopic angiogram W contrast IA|Superior mesenteric artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37402-5|LNC|Superior mesenteric artery and Inferior mesenteric artery Fluoroscopic angiogram W contrast IA|Superior mesenteric artery and Inferior mesenteric artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|38119-4|LNC|Thoracic artery Fluoroscopic angiogram W contrast IA|Thoracic artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37900-8|LNC|Tibial artery Fluoroscopic angiogram W contrast IA|Tibial artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37489-2|LNC|Tibioperoneal arteries Fluoroscopic angiogram W contrast IA|Tibioperoneal arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37977-6|LNC|Upper extremity arteries Fluoroscopic angiogram W contrast IA|Upper extremity arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37396-9|LNC|Upper extremity arteries - bilateral Fluoroscopic angiogram W contrast IA|Upper extremity arteries - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37488-4|LNC|Upper extremity arteries - left Fluoroscopic angiogram W contrast IA|Upper extremity arteries - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37967-7|LNC|Upper extremity arteries - right Fluoroscopic angiogram W contrast IA|Upper extremity arteries - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|24576-1|LNC|Urinary bladder arteries Fluoroscopic angiogram W contrast IA|Urinary bladder arteries Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37979-2|LNC|Uterine artery Fluoroscopic angiogram W contrast IA|Uterine artery Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37407-4|LNC|Vertebral artery - bilateral Fluoroscopic angiogram W contrast IA|Vertebral artery - bilateral Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37490-0|LNC|Vertebral artery - left Fluoroscopic angiogram W contrast IA|Vertebral artery - left Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|37968-5|LNC|Vertebral artery - right Fluoroscopic angiogram W contrast IA|Vertebral artery - right Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|42156-0|LNC|Vessels Fluoroscopic angiogram W contrast IA|Vessels Fluoroscopic angiogram W contrast IA
C2826012|T102|strict|25017-5|LNC|Urinary Bladder and Urethra Fluoroscopy W contrast intra bladder|Urinary Bladder and Urethra Fluoroscopy W contrast intra bladder
C2826012|T102|strict|43559-4|LNC|Urinary Bladder and Urethra Fluoroscopy W contrast intra bladder during voiding|Urinary Bladder and Urethra Fluoroscopy W contrast intra bladder during voiding
C2826012|T102|strict|37586-5|LNC|Penis Fluoroscopy W contrast intra corpus cavernosum|Penis Fluoroscopy W contrast intra corpus cavernosum
C2826012|T102|strict|39054-2|LNC|Breast duct Mammogram W contrast intra duct|Breast duct Mammogram W contrast intra duct
C2826012|T102|strict|38095-6|LNC|Breast duct - bilateral Mammogram W contrast intra duct|Breast duct - bilateral Mammogram W contrast intra duct
C2826012|T102|strict|38096-4|LNC|Breast duct - left Mammogram W contrast intra duct|Breast duct - left Mammogram W contrast intra duct
C2826012|T102|strict|38825-6|LNC|Breast duct - right Mammogram W contrast intra duct|Breast duct - right Mammogram W contrast intra duct
C2826012|T102|strict|30810-6|LNC|Lacrimal duct Fluoroscopy W contrast intra lacrimal duct|Lacrimal duct Fluoroscopy W contrast intra lacrimal duct
C2826012|T102|strict|38098-0|LNC|Lacrimal duct - bilateral Fluoroscopy W contrast intra lacrimal duct|Lacrimal duct - bilateral Fluoroscopy W contrast intra lacrimal duct
C2826012|T102|strict|38099-8|LNC|Lacrimal duct - left Fluoroscopy W contrast intra lacrimal duct|Lacrimal duct - left Fluoroscopy W contrast intra lacrimal duct
C2826012|T102|strict|38827-2|LNC|Lacrimal duct - right Fluoroscopy W contrast intra lacrimal duct|Lacrimal duct - right Fluoroscopy W contrast intra lacrimal duct
C2826012|T102|strict|24845-0|LNC|Neck Fluoroscopy W contrast intra larynx|Neck Fluoroscopy W contrast intra larynx
C2826012|T102|strict|30850-2|LNC|Extremity lymphatics Fluoroscopy W contrast intra lymphatic|Extremity lymphatics Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|30851-0|LNC|Extremity lymphatics - bilateral Fluoroscopy W contrast intra lymphatic|Extremity lymphatics - bilateral Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|37599-8|LNC|Extremity lymphatics - left Fluoroscopy W contrast intra lymphatic|Extremity lymphatics - left Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|38812-4|LNC|Extremity lymphatics - right Fluoroscopy W contrast intra lymphatic|Extremity lymphatics - right Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|24827-8|LNC|Lymphatics Fluoroscopy W contrast intra lymphatic|Lymphatics Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|30839-5|LNC|Lymphatics abdominal Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|30840-3|LNC|Lymphatics abdominal - bilateral Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal - bilateral Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|37597-2|LNC|Lymphatics abdominal and Lymphatics pelvic Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal and Lymphatics pelvic Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|37598-0|LNC|Lymphatics abdominal and Lymphatics pelvic - bilateral Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal and Lymphatics pelvic - bilateral Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|37596-4|LNC|Lymphatics abdominal and Lymphatics pelvic - left Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal and Lymphatics pelvic - left Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|38811-6|LNC|Lymphatics abdominal and Lymphatics pelvic - right Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal and Lymphatics pelvic - right Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|37600-4|LNC|Lymphatics - left Fluoroscopy W contrast intra lymphatic|Lymphatics - left Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|39510-3|LNC|Lymphatics pelvic Fluoroscopy W contrast intra lymphatic|Lymphatics pelvic Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|37601-2|LNC|Lymphatics pelvic - bilateral Fluoroscopy W contrast intra lymphatic|Lymphatics pelvic - bilateral Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|38813-2|LNC|Lymphatics - right Fluoroscopy W contrast intra lymphatic|Lymphatics - right Fluoroscopy W contrast intra lymphatic
C2826012|T102|strict|39148-2|LNC|Breast duct Mammogram W contrast intra multiple ducts|Breast duct Mammogram W contrast intra multiple ducts
C2826012|T102|strict|39146-6|LNC|Breast duct - bilateral Mammogram W contrast intra multiple ducts|Breast duct - bilateral Mammogram W contrast intra multiple ducts
C2826012|T102|strict|39145-8|LNC|Breast duct - left Mammogram W contrast intra multiple ducts|Breast duct - left Mammogram W contrast intra multiple ducts
C2826012|T102|strict|39147-4|LNC|Breast duct - right Mammogram W contrast intra multiple ducts|Breast duct - right Mammogram W contrast intra multiple ducts
C2826012|T102|strict|24661-1|LNC|Pleural space Fluoroscopy W contrast intra pleural space|Pleural space Fluoroscopy W contrast intra pleural space
C2826012|T102|strict|38116-0|LNC|Parotid gland Fluoroscopy W contrast intra salivary duct|Parotid gland Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|38097-2|LNC|Parotid gland - left Fluoroscopy W contrast intra salivary duct|Parotid gland - left Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|38826-4|LNC|Parotid gland - right Fluoroscopy W contrast intra salivary duct|Parotid gland - right Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|24902-9|LNC|Salivary gland Fluoroscopy W contrast intra salivary duct|Salivary gland Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|26067-9|LNC|Salivary gland - bilateral Fluoroscopy W contrast intra salivary duct|Salivary gland - bilateral Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|26068-7|LNC|Salivary gland - left Fluoroscopy W contrast intra salivary duct|Salivary gland - left Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|26069-5|LNC|Salivary gland - right Fluoroscopy W contrast intra salivary duct|Salivary gland - right Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|38153-3|LNC|Submandibular gland Fluoroscopy W contrast intra salivary duct|Submandibular gland Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|48698-5|LNC|Submandibular gland - bilateral Fluoroscopy W contrast intra salivary duct|Submandibular gland - bilateral Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|42460-6|LNC|Submandibular gland - left Fluoroscopy W contrast intra salivary duct|Submandibular gland - left Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|48696-9|LNC|Submandibular gland - right Fluoroscopy W contrast intra salivary duct|Submandibular gland - right Fluoroscopy W contrast intra salivary duct
C2826012|T102|strict|24912-8|LNC|Sinus tract Fluoroscopy W contrast intra sinus tract|Sinus tract Fluoroscopy W contrast intra sinus tract
C2826012|T102|strict|24552-2|LNC|Stent Fluoroscopy W contrast intra stent|Stent Fluoroscopy W contrast intra stent
C2826012|T102|strict|25016-7|LNC|Urethra Fluoroscopy W contrast intra urethra|Urethra Fluoroscopy W contrast intra urethra
C2826012|T102|strict|39151-6|LNC|Vas deferens Fluoroscopy W contrast intra vas deferens|Vas deferens Fluoroscopy W contrast intra vas deferens
C2826012|T102|strict|37183-1|LNC|Ankle Fluoroscopy W contrast intraarticular|Ankle Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37184-9|LNC|Ankle - bilateral Fluoroscopy W contrast intraarticular|Ankle - bilateral Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37185-6|LNC|Ankle - left Fluoroscopy W contrast intraarticular|Ankle - left Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37942-0|LNC|Ankle - right Fluoroscopy W contrast intraarticular|Ankle - right Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37186-4|LNC|Elbow Fluoroscopy W contrast intraarticular|Elbow Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37187-2|LNC|Elbow - bilateral Fluoroscopy W contrast intraarticular|Elbow - bilateral Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37188-0|LNC|Elbow - left Fluoroscopy W contrast intraarticular|Elbow - left Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37947-9|LNC|Elbow - right Fluoroscopy W contrast intraarticular|Elbow - right Fluoroscopy W contrast intraarticular
C2826012|T102|strict|24764-3|LNC|Hip Fluoroscopy W contrast intraarticular|Hip Fluoroscopy W contrast intraarticular
C2826012|T102|strict|26070-3|LNC|Hip - bilateral Fluoroscopy W contrast intraarticular|Hip - bilateral Fluoroscopy W contrast intraarticular
C2826012|T102|strict|26071-1|LNC|Hip - left Fluoroscopy W contrast intraarticular|Hip - left Fluoroscopy W contrast intraarticular
C2826012|T102|strict|26072-9|LNC|Hip - right Fluoroscopy W contrast intraarticular|Hip - right Fluoroscopy W contrast intraarticular
C2826012|T102|strict|24800-5|LNC|Knee Fluoroscopy W contrast intraarticular|Knee Fluoroscopy W contrast intraarticular
C2826012|T102|strict|26073-7|LNC|Knee - bilateral Fluoroscopy W contrast intraarticular|Knee - bilateral Fluoroscopy W contrast intraarticular
C2826012|T102|strict|26074-5|LNC|Knee - left Fluoroscopy W contrast intraarticular|Knee - left Fluoroscopy W contrast intraarticular
C2826012|T102|strict|26075-2|LNC|Knee - right Fluoroscopy W contrast intraarticular|Knee - right Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37647-5|LNC|Sacroiliac Joint Fluoroscopy W contrast intraarticular|Sacroiliac Joint Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37189-8|LNC|Sacroiliac joint - bilateral Fluoroscopy W contrast intraarticular|Sacroiliac joint - bilateral Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37190-6|LNC|Sacroiliac joint - left Fluoroscopy W contrast intraarticular|Sacroiliac joint - left Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37785-3|LNC|Sacroiliac joint - right Fluoroscopy W contrast intraarticular|Sacroiliac joint - right Fluoroscopy W contrast intraarticular
C2826012|T102|strict|24910-2|LNC|Shoulder Fluoroscopy W contrast intraarticular|Shoulder Fluoroscopy W contrast intraarticular
C2826012|T102|strict|26076-0|LNC|Shoulder - bilateral Fluoroscopy W contrast intraarticular|Shoulder - bilateral Fluoroscopy W contrast intraarticular
C2826012|T102|strict|26077-8|LNC|Shoulder - left Fluoroscopy W contrast intraarticular|Shoulder - left Fluoroscopy W contrast intraarticular
C2826012|T102|strict|26078-6|LNC|Shoulder - right Fluoroscopy W contrast intraarticular|Shoulder - right Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37901-6|LNC|Temporomandibular joint Fluoroscopy W contrast intraarticular|Temporomandibular joint Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37409-0|LNC|Temporomandibular joint - bilateral Fluoroscopy W contrast intraarticular|Temporomandibular joint - bilateral Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37410-8|LNC|Temporomandibular joint - left Fluoroscopy W contrast intraarticular|Temporomandibular joint - left Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37818-2|LNC|Temporomandibular joint - right Fluoroscopy W contrast intraarticular|Temporomandibular joint - right Fluoroscopy W contrast intraarticular
C2826012|T102|strict|25034-0|LNC|Wrist Fluoroscopy W contrast intraarticular|Wrist Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37570-9|LNC|Wrist - bilateral Fluoroscopy W contrast intraarticular|Wrist - bilateral Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37571-7|LNC|Wrist - left Fluoroscopy W contrast intraarticular|Wrist - left Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37641-8|LNC|Wrist - right Fluoroscopy W contrast intraarticular|Wrist - right Fluoroscopy W contrast intraarticular
C2826012|T102|strict|37191-4|LNC|Joint Fluoroscopy W contrast intraarticular|Joint Fluoroscopy W contrast intraarticular
C2826012|T102|strict|24825-2|LNC|Lung X-ray W contrast intrabronchial|Lung X-ray W contrast intrabronchial
C2826012|T102|strict|30813-0|LNC|Lung - bilateral X-ray W contrast intrabronchial|Lung - bilateral X-ray W contrast intrabronchial
C2826012|T102|strict|64996-2|LNC|Lung - left X-ray W contrast intrabronchial|Lung - left X-ray W contrast intrabronchial
C2826012|T102|strict|64997-0|LNC|Lung - right X-ray W contrast intrabronchial|Lung - right X-ray W contrast intrabronchial
C2826012|T102|strict|24927-6|LNC|Spine Fluoroscopy W contrast intradisc|Spine Fluoroscopy W contrast intradisc
C2826012|T102|strict|37192-2|LNC|Spine Cervical Fluoroscopy W contrast intradisc|Spine Cervical Fluoroscopy W contrast intradisc
C2826012|T102|strict|37193-0|LNC|Spine Lumbar Fluoroscopy W contrast intradisc|Spine Lumbar Fluoroscopy W contrast intradisc
C2826012|T102|strict|70933-7|LNC|Spine Thoracic Fluoroscopy W contrast intradisc|Spine Thoracic Fluoroscopy W contrast intradisc
C2826012|T102|strict|25022-5|LNC|Uterus and Fallopian tubes Fluoroscopy W contrast intrauterine|Uterus and Fallopian tubes Fluoroscopy W contrast intrauterine
C2826012|T102|strict|30811-4|LNC|Posterior fossa Fluoroscopy W contrast IT|Posterior fossa Fluoroscopy W contrast IT
C2826012|T102|strict|37572-5|LNC|Spine Fluoroscopy W contrast IT|Spine Fluoroscopy W contrast IT
C2826012|T102|strict|24947-4|LNC|Spine Cervical Fluoroscopy W contrast IT|Spine Cervical Fluoroscopy W contrast IT
C2826012|T102|strict|38103-8|LNC|Spine Cervical and Spine Lumbar Fluoroscopy W contrast IT|Spine Cervical and Spine Lumbar Fluoroscopy W contrast IT
C2826012|T102|strict|30808-0|LNC|Spine Cervical and Thoracic and Lumbar Fluoroscopy W contrast IT|Spine Cervical and Thoracic and Lumbar Fluoroscopy W contrast IT
C2826012|T102|strict|38104-6|LNC|Spine.epidural space Fluoroscopy W contrast IT|Spine.epidural space Fluoroscopy W contrast IT
C2826012|T102|strict|24974-8|LNC|Spine Lumbar Fluoroscopy W contrast IT|Spine Lumbar Fluoroscopy W contrast IT
C2826012|T102|strict|24985-4|LNC|Spine Thoracic Fluoroscopy W contrast IT|Spine Thoracic Fluoroscopy W contrast IT
C2826012|T102|strict|69066-9|LNC|Abdominal vessels Fluoroscopic angiogram W contrast IV|Abdominal vessels Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30843-7|LNC|Adrenal vein Fluoroscopic angiogram W contrast IV|Adrenal vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37602-0|LNC|Adrenal vein left Fluoroscopic angiogram W contrast IV|Adrenal vein left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30844-5|LNC|Adrenal vein - bilateral Fluoroscopic angiogram W contrast IV|Adrenal vein - bilateral Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37940-4|LNC|Adrenal vein - right Fluoroscopic angiogram W contrast IV|Adrenal vein - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|58746-9|LNC|AV fistula Fluoroscopic angiogram W contrast IV|AV fistula Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|24569-6|LNC|AV shunt Fluoroscopic angiogram W contrast IV|AV shunt Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37411-6|LNC|Azygos vein Fluoroscopic angiogram W contrast IV|Azygos vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|24573-8|LNC|Biliary ducts and Gallbladder X-ray W contrast IV|Biliary ducts and Gallbladder X-ray W contrast IV
C2826012|T102|strict|37195-5|LNC|Cerebral vein Fluoroscopic angiogram W contrast IV|Cerebral vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30819-7|LNC|Epidural veins Fluoroscopic angiogram W contrast IV|Epidural veins Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|39055-9|LNC|Extremity veins Fluoroscopic angiogram W contrast IV|Extremity veins Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37412-4|LNC|Extremity veins - bilateral Fluoroscopic angiogram W contrast IV|Extremity veins - bilateral Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37413-2|LNC|Extremity veins - left Fluoroscopic angiogram W contrast IV|Extremity veins - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37950-3|LNC|Extremity veins - right Fluoroscopic angiogram W contrast IV|Extremity veins - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|42157-8|LNC|Extremity vessels Fluoroscopic angiogram W contrast IV|Extremity vessels Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37416-5|LNC|Femoral vein Fluoroscopic angiogram W contrast IV|Femoral vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|39093-0|LNC|Hepatic veins Fluoroscopic angiogram W contrast IV|Hepatic veins Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37421-5|LNC|Inferior mesenteric vein Fluoroscopic angiogram W contrast IV|Inferior mesenteric vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37419-9|LNC|Intraosseous veins Fluoroscopic angiogram W contrast IV|Intraosseous veins Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37197-1|LNC|Jugular vein Fluoroscopic angiogram W contrast IV|Jugular vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37420-7|LNC|Jugular vein - left Fluoroscopic angiogram W contrast IV|Jugular vein - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37954-5|LNC|Jugular vein - right Fluoroscopic angiogram W contrast IV|Jugular vein - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37607-9|LNC|Kidney X-ray W contrast IV|Kidney X-ray W contrast IV
C2826012|T102|strict|24788-2|LNC|Kidney - bilateral X-ray W contrast IV|Kidney - bilateral X-ray W contrast IV
C2826012|T102|strict|37414-0|LNC|Lower extremity veins - bilateral Fluoroscopic angiogram W contrast IV|Lower extremity veins - bilateral Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37196-3|LNC|Lower extremity veins - left Fluoroscopic angiogram W contrast IV|Lower extremity veins - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37767-1|LNC|Lower extremity veins - right Fluoroscopic angiogram W contrast IV|Lower extremity veins - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37574-1|LNC|Lower extremity vessels Fluoroscopic angiogram W contrast IV|Lower extremity vessels Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30825-4|LNC|Orbit veins Fluoroscopic angiogram W contrast IV|Orbit veins Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37422-3|LNC|Orbit veins - left Fluoroscopic angiogram W contrast IV|Orbit veins - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37958-6|LNC|Orbit veins - right Fluoroscopic angiogram W contrast IV|Orbit veins - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30852-8|LNC|Peripheral veins - bilateral Fluoroscopic angiogram W contrast IV|Peripheral veins - bilateral Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|24685-0|LNC|Peripheral veins Fluoroscopic angiogram W contrast IV|Peripheral veins Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|69250-9|LNC|Portal vein Fluoroscopic angiogram W contrast IV|Portal vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30847-8|LNC|Renal vein Fluoroscopic angiogram W contrast IV|Renal vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30846-0|LNC|Renal vein - bilateral Fluoroscopic angiogram W contrast IV|Renal vein - bilateral Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37423-1|LNC|Renal vein - left Fluoroscopic angiogram W contrast IV|Renal vein - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37959-4|LNC|Renal vein - right Fluoroscopic angiogram W contrast IV|Renal vein - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30827-0|LNC|Sagittal sinus vein Fluoroscopic angiogram W contrast IV|Sagittal sinus vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|65803-9|LNC|Sagittal sinus vein - left Fluoroscopic angiogram W contrast IV|Sagittal sinus vein - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|65802-1|LNC|Sagittal sinus and Jugular veins - left Fluoroscopic angiogram W contrast IV|Sagittal sinus and Jugular veins - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|65804-7|LNC|Sagittal sinus vein - right Fluoroscopic angiogram W contrast IV|Sagittal sinus vein - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|65805-4|LNC|Sagittal sinus and Jugular veins - right Fluoroscopic angiogram W contrast IV|Sagittal sinus and Jugular veins - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30826-2|LNC|Sagittal sinus and Jugular veins Fluoroscopic angiogram W contrast IV|Sagittal sinus and Jugular veins Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37969-3|LNC|Sinus vein Fluoroscopic angiogram W contrast IV|Sinus vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37970-1|LNC|Splenic vein Fluoroscopic angiogram W contrast IV|Splenic vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37971-9|LNC|Subclavian vein Fluoroscopic angiogram W contrast IV|Subclavian vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37972-7|LNC|Superior mesenteric vein Fluoroscopic angiogram W contrast IV|Superior mesenteric vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|24550-6|LNC|Upper extremity veins Fluoroscopic angiogram W contrast IV|Upper extremity veins Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37415-7|LNC|Upper extremity veins - bilateral Fluoroscopic angiogram W contrast IV|Upper extremity veins - bilateral Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|38859-5|LNC|Upper extremity veins - left Fluoroscopic angiogram W contrast IV|Upper extremity veins - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|37824-0|LNC|Upper extremity veins - right Fluoroscopic angiogram W contrast IV|Upper extremity veins - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|25023-3|LNC|Vein Fluoroscopic angiogram W contrast IV|Vein Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|26064-6|LNC|Vein - bilateral Fluoroscopic angiogram W contrast IV|Vein - bilateral Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|26065-3|LNC|Vein - left Fluoroscopic angiogram W contrast IV|Vein - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|26066-1|LNC|Vein - right Fluoroscopic angiogram W contrast IV|Vein - right Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|25025-8|LNC|Vena cava Fluoroscopic angiogram W contrast IV|Vena cava Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30845-2|LNC|Inferior vena cava Fluoroscopic angiogram W contrast IV|Inferior vena cava Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|30645-6|LNC|Superior vena cava Fluoroscopic angiogram W contrast IV|Superior vena cava Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|43554-5|LNC|vessels - left Fluoroscopic angiogram W contrast IV|vessels - left Fluoroscopic angiogram W contrast IV
C2826012|T102|strict|39096-3|LNC|Hepatic veins Fluoroscopic angiogram W contrast IV and W hemodynamics|Hepatic veins Fluoroscopic angiogram W contrast IV and W hemodynamics
C2826012|T102|strict|43783-0|LNC|Renal vein Fluoroscopic angiogram W contrast IV and W renin sampling|Renal vein Fluoroscopic angiogram W contrast IV and W renin sampling
C2826012|T102|strict|25080-3|LNC|Renal vein - bilateral Fluoroscopic angiogram W contrast IV and W renin sampling|Renal vein - bilateral Fluoroscopic angiogram W contrast IV and W renin sampling
C2826012|T102|strict|30816-3|LNC|Peritoneum Fluoroscopic angiogram W contrast percutaneous|Peritoneum Fluoroscopic angiogram W contrast percutaneous
C2826012|T102|strict|24575-3|LNC|Biliary ducts and Gallbladder Fluoroscopy W contrast percutaneous transhepatic|Biliary ducts and Gallbladder Fluoroscopy W contrast percutaneous transhepatic
C2826012|T102|strict|37200-3|LNC|Chest X-ray W contrast PO|Chest X-ray W contrast PO
C2826012|T102|strict|37199-7|LNC|Chest Fluoroscopy W contrast PO|Chest Fluoroscopy W contrast PO
C2826012|T102|strict|37198-9|LNC|Esophagus X-ray W contrast PO|Esophagus X-ray W contrast PO
C2826012|T102|strict|24678-5|LNC|Esophagus Fluoroscopy W contrast PO|Esophagus Fluoroscopy W contrast PO
C2826012|T102|strict|24712-2|LNC|Gallbladder X-ray W contrast PO|Gallbladder X-ray W contrast PO
C2826012|T102|strict|42459-8|LNC|Gastrointestine upper Fluoroscopy W contrast PO|Gastrointestine upper Fluoroscopy W contrast PO
C2826012|T102|strict|24924-3|LNC|Small bowel Fluoroscopy W contrast PO|Small bowel Fluoroscopy W contrast PO
C2826012|T102|strict|24673-6|LNC|Duodenum Fluoroscopy W contrast PO and hypotonic agent per ng|Duodenum Fluoroscopy W contrast PO and hypotonic agent per ng
C2826012|T102|strict|24681-9|LNC|Esophagus and Hypopharynx Fluoroscopy video W contrast PO during swallowing|Esophagus and Hypopharynx Fluoroscopy video W contrast PO during swallowing
C2826012|T102|strict|24667-8|LNC|Colon Fluoroscopy W contrast PR|Colon Fluoroscopy W contrast PR
C2826012|T102|strict|24894-8|LNC|Rectum and Urinary bladder Fluoroscopy W contrast PR and intra bladder during defecation and voiding|Rectum and Urinary bladder Fluoroscopy W contrast PR and intra bladder during defecation and voiding
C2826012|T102|strict|39363-7|LNC|Fistula Fluoroscopy W contrast retrograde|Fistula Fluoroscopy W contrast retrograde
C2826012|T102|strict|38105-3|LNC|Kidney X-ray W contrast retrograde|Kidney X-ray W contrast retrograde
C2826012|T102|strict|39349-6|LNC|Kidney - bilateral Fluoroscopy W contrast retrograde|Kidney - bilateral Fluoroscopy W contrast retrograde
C2826012|T102|strict|30761-1|LNC|Kidney - bilateral Fluoroscopy W contrast retrograde via urethra|Kidney - bilateral Fluoroscopy W contrast retrograde via urethra
C2826012|T102|strict|38873-6|LNC|Kidney - left and Collecting system Fluoroscopy W contrast retrograde via urethra|Kidney - left and Collecting system Fluoroscopy W contrast retrograde via urethra
C2826012|T102|strict|38113-7|LNC|Kidney - right and Collecting system Fluoroscopy W contrast retrograde via urethra|Kidney - right and Collecting system Fluoroscopy W contrast retrograde via urethra
C2826012|T102|strict|25020-9|LNC|Urinary Bladder and Urethra Fluoroscopy W contrast retrograde via urethra|Urinary Bladder and Urethra Fluoroscopy W contrast retrograde via urethra
C2826012|T102|strict|30841-1|LNC|Portal vein Fluoroscopic angiogram W contrast transhepatic|Portal vein Fluoroscopic angiogram W contrast transhepatic
C2826012|T102|strict|30842-9|LNC|Portal vein Fluoroscopic angiogram W contrast transhepatic and W hemodynamics|Portal vein Fluoroscopic angiogram W contrast transhepatic and W hemodynamics
C2826012|T102|strict|37566-7|LNC|Unspecified body region Fluoroscopy W contrast via catheter|Unspecified body region Fluoroscopy W contrast via catheter
C2826012|T102|strict|37567-5|LNC|Colon Fluoroscopy W contrast via colostomy|Colon Fluoroscopy W contrast via colostomy
C2826012|T102|strict|37568-3|LNC|Unspecified body region Fluoroscopy W contrast via fistula|Unspecified body region Fluoroscopy W contrast via fistula
C2826012|T102|strict|69272-3|LNC|Small bowel Fluoroscopy W contrast via ileostomy|Small bowel Fluoroscopy W contrast via ileostomy
C2826012|T102|strict|24780-9|LNC|Kidney - bilateral Fluoroscopy W contrast via nephrostomy tube|Kidney - bilateral Fluoroscopy W contrast via nephrostomy tube
C2826012|T102|strict|38872-8|LNC|Kidney - left and Collecting system Fluoroscopy W contrast via nephrostomy tube|Kidney - left and Collecting system Fluoroscopy W contrast via nephrostomy tube
C2826012|T102|strict|38112-9|LNC|Kidney - right and Collecting system Fluoroscopy W contrast via nephrostomy tube|Kidney - right and Collecting system Fluoroscopy W contrast via nephrostomy tube
C2826012|T102|strict|37569-1|LNC|Urinary bladder Fluoroscopy W contrast via suprapubic tube|Urinary bladder Fluoroscopy W contrast via suprapubic tube
C2826012|T102|strict|30647-2|LNC|Biliary ducts and Gallbladder Fluoroscopy W contrast via T-tube|Biliary ducts and Gallbladder Fluoroscopy W contrast via T-tube
C2826012|T102|strict|39696-0|LNC|Lung Scan W depreotide and W radionuclide IV|Lung Scan W depreotide and W radionuclide IV
C2826012|T102|strict|42161-0|LNC|Heart Scan W dobutamine and W radionuclide IV|Heart Scan W dobutamine and W radionuclide IV
C2826012|T102|strict|39652-3|LNC|Heart Scan W dobutamine and W Tl-201 IV|Heart Scan W dobutamine and W Tl-201 IV
C2826012|T102|strict|42383-0|LNC|Gallbladder X-ray W double dose contrast PO|Gallbladder X-ray W double dose contrast PO
C2826012|T102|strict|42690-8|LNC|Spine X-ray W flexion and W extension|Spine X-ray W flexion and W extension
C2826012|T102|strict|24945-8|LNC|Spine Cervical X-ray W flexion and W extension|Spine Cervical X-ray W flexion and W extension
C2826012|T102|strict|24971-4|LNC|Spine Lumbar X-ray W flexion and W extension|Spine Lumbar X-ray W flexion and W extension
C2826012|T102|strict|43481-1|LNC|Joint X-ray W flexion and W extension|Joint X-ray W flexion and W extension
C2826012|T102|strict|30785-0|LNC|Foot X-ray W forced dorsiflexion|Foot X-ray W forced dorsiflexion
C2826012|T102|strict|43461-3|LNC|Kidney - bilateral Scan W furosemide and W radionuclide IV|Kidney - bilateral Scan W furosemide and W radionuclide IV
C2826012|T102|strict|39688-7|LNC|Scan W GA-67 IV|Scan W GA-67 IV
C2826012|T102|strict|24679-3|LNC|Esophagus Fluoroscopy W gastrografin PO|Esophagus Fluoroscopy W gastrografin PO
C2826012|T102|strict|42684-1|LNC|Gastrointestine upper Fluoroscopy W gastrografin PO|Gastrointestine upper Fluoroscopy W gastrografin PO
C2826012|T102|strict|42681-7|LNC|Colon Fluoroscopy W gastrografin PR|Colon Fluoroscopy W gastrografin PR
C2826012|T102|strict|37576-6|LNC|Unspecified body region Fluoroscopy W gastrografin via fistula|Unspecified body region Fluoroscopy W gastrografin via fistula
C2826012|T102|strict|39850-3|LNC|Kidney - bilateral Scan W I-131 IV|Kidney - bilateral Scan W I-131 IV
C2826012|T102|strict|25007-6|LNC|Thyroid Scan W I-131 IV|Thyroid Scan W I-131 IV
C2826012|T102|strict|39841-2|LNC|Scan W I-131 MIBG IV|Scan W I-131 MIBG IV
C2826012|T102|strict|39857-8|LNC|Adrenal gland Scan W I-131 MIBG IV|Adrenal gland Scan W I-131 MIBG IV
C2826012|T102|strict|39624-2|LNC|Adrenal gland Scan W I-131 NP59 IV|Adrenal gland Scan W I-131 NP59 IV
C2826012|T102|strict|24770-0|LNC|Joint Scan W In-111 intrajoint|Joint Scan W In-111 intrajoint
C2826012|T102|strict|39846-1|LNC|Scan W In-111 Satumomab IV|Scan W In-111 Satumomab IV
C2826012|T102|strict|39738-0|LNC|Abdomen Scan W In-111 Satumomab IV|Abdomen Scan W In-111 Satumomab IV
C2826012|T102|strict|25032-4|LNC|Bone Scan W In-111 tagged WBC IV|Bone Scan W In-111 tagged WBC IV
C2826012|T102|strict|42708-8|LNC|Scan W In-111 tiuxetan IV|Scan W In-111 tiuxetan IV
C2826012|T102|strict|30736-3|LNC|Chest X-ray W inspiration and expiration|Chest X-ray W inspiration and expiration
C2826012|T102|strict|24682-7|LNC|Esophagus and Hypopharynx Fluoroscopy video W liquid and paste contrast PO during swallowing|Esophagus and Hypopharynx Fluoroscopy video W liquid and paste contrast PO during swallowing
C2826012|T102|strict|37556-8|LNC|Ankle X-ray W manual stress|Ankle X-ray W manual stress
C2826012|T102|strict|37557-6|LNC|Ankle - bilateral X-ray W manual stress|Ankle - bilateral X-ray W manual stress
C2826012|T102|strict|37558-4|LNC|Ankle - left X-ray W manual stress|Ankle - left X-ray W manual stress
C2826012|T102|strict|37673-1|LNC|Ankle - right X-ray W manual stress|Ankle - right X-ray W manual stress
C2826012|T102|strict|37559-2|LNC|Foot - left X-ray W manual stress|Foot - left X-ray W manual stress
C2826012|T102|strict|37705-1|LNC|Foot - right X-ray W manual stress|Foot - right X-ray W manual stress
C2826012|T102|strict|37560-0|LNC|Knee X-ray W manual stress|Knee X-ray W manual stress
C2826012|T102|strict|37561-8|LNC|Knee - bilateral X-ray W manual stress|Knee - bilateral X-ray W manual stress
C2826012|T102|strict|37562-6|LNC|Knee - left X-ray W manual stress|Knee - left X-ray W manual stress
C2826012|T102|strict|37753-1|LNC|Knee - right X-ray W manual stress|Knee - right X-ray W manual stress
C2826012|T102|strict|37563-4|LNC|Thumb - bilateral X-ray W manual stress|Thumb - bilateral X-ray W manual stress
C2826012|T102|strict|37564-2|LNC|Thumb - left X-ray W manual stress|Thumb - left X-ray W manual stress
C2826012|T102|strict|37814-1|LNC|Thumb - right X-ray W manual stress|Thumb - right X-ray W manual stress
C2826012|T102|strict|39056-7|LNC|Unspecified body region X-ray W manual stress|Unspecified body region X-ray W manual stress
C2826012|T102|strict|38093-1|LNC|Chest X-ray W nipple markers|Chest X-ray W nipple markers
C2826012|T102|strict|39670-5|LNC|Lacrimal duct Scan W radionuclide intra lacrimal duct|Lacrimal duct Scan W radionuclide intra lacrimal duct
C2826012|T102|strict|64051-6|LNC|Breast lymphatics - left Scan W radionuclide intra lymphatic|Breast lymphatics - left Scan W radionuclide intra lymphatic
C2826012|T102|strict|64052-4|LNC|Breast lymphatics - right Scan W radionuclide intra lymphatic|Breast lymphatics - right Scan W radionuclide intra lymphatic
C2826012|T102|strict|24826-0|LNC|Lymphatics Scan W radionuclide intra lymphatic|Lymphatics Scan W radionuclide intra lymphatic
C2826012|T102|strict|24663-7|LNC|Head Cistern Scan W radionuclide IT|Head Cistern Scan W radionuclide IT
C2826012|T102|strict|42158-6|LNC|Adrenal gland Scan|Adrenal gland Scan
C2826012|T102|strict|42776-5|LNC|AV shunt Scan|AV shunt Scan
C2826012|T102|strict|25031-6|LNC|Bone Scan|Bone Scan
C2826012|T102|strict|24730-4|LNC|Brain Scan|Brain Scan
C2826012|T102|strict|39643-2|LNC|Brain veins Scan|Brain veins Scan
C2826012|T102|strict|39646-5|LNC|Breast Scan|Breast Scan
C2826012|T102|strict|39650-7|LNC|Heart Scan|Heart Scan
C2826012|T102|strict|24776-7|LNC|Kidney - bilateral Scan|Kidney - bilateral Scan
C2826012|T102|strict|30877-5|LNC|Kidney - bilateral and Renal vessels Scan|Kidney - bilateral and Renal vessels Scan
C2826012|T102|strict|24804-7|LNC|Knee Scan|Knee Scan
C2826012|T102|strict|26088-5|LNC|Knee - bilateral Scan|Knee - bilateral Scan
C2826012|T102|strict|26089-3|LNC|Knee - left Scan|Knee - left Scan
C2826012|T102|strict|26090-1|LNC|Knee - right Scan|Knee - right Scan
C2826012|T102|strict|39693-7|LNC|Liver Scan|Liver Scan
C2826012|T102|strict|39694-5|LNC|Liver transplant Scan|Liver transplant Scan
C2826012|T102|strict|43557-8|LNC|Liver and Biliary ducts and Gallbladder Scan|Liver and Biliary ducts and Gallbladder Scan
C2826012|T102|strict|39897-4|LNC|Liver and Lung Scan|Liver and Lung Scan
C2826012|T102|strict|39877-6|LNC|Liver and Spleen Scan|Liver and Spleen Scan
C2826012|T102|strict|39629-1|LNC|Meckels diverticulum Scan|Meckels diverticulum Scan
C2826012|T102|strict|39737-2|LNC|Neck Scan|Neck Scan
C2826012|T102|strict|39739-8|LNC|Pancreas Scan|Pancreas Scan
C2826012|T102|strict|39742-2|LNC|Parathyroid Scan|Parathyroid Scan
C2826012|T102|strict|39619-2|LNC|Pulmonary system Scan|Pulmonary system Scan
C2826012|T102|strict|43669-1|LNC|Renal vessels Scan|Renal vessels Scan
C2826012|T102|strict|39747-1|LNC|Salivary gland Scan|Salivary gland Scan
C2826012|T102|strict|30696-9|LNC|Scrotum and Testicle Scan|Scrotum and Testicle Scan
C2826012|T102|strict|39751-3|LNC|Spleen Scan|Spleen Scan
C2826012|T102|strict|30695-1|LNC|Thyroid Scan|Thyroid Scan
C2826012|T102|strict|25018-3|LNC|Urinary bladder Scan|Urinary bladder Scan
C2826012|T102|strict|39626-7|LNC|Vein - bilateral Scan|Vein - bilateral Scan
C2826012|T102|strict|49118-3|LNC|Unspecified body region Scan|Unspecified body region Scan
C2826012|T102|strict|39939-4|LNC|Joint Scan|Joint Scan
C2826012|T102|strict|39671-3|LNC|Rectum Scan W radionuclide PO|Rectum Scan W radionuclide PO
C2826012|T102|strict|39752-1|LNC|Spleen Scan W radionuclide tagged heat damaged RBC IV|Spleen Scan W radionuclide tagged heat damaged RBC IV
C2826012|T102|strict|24773-4|LNC|Kidney - bilateral Scan W radionuclide transplant scan|Kidney - bilateral Scan W radionuclide transplant scan
C2826012|T102|strict|30713-2|LNC|Spine X-ray W right bending and W left bending|Spine X-ray W right bending and W left bending
C2826012|T102|strict|42413-5|LNC|Spine Lumbar X-ray W right bending and W left bending|Spine Lumbar X-ray W right bending and W left bending
C2826012|T102|strict|43651-9|LNC|Liver and Biliary ducts and Gallbladder Scan W sincalide and W radionuclide IV|Liver and Biliary ducts and Gallbladder Scan W sincalide and W radionuclide IV
C2826012|T102|strict|39820-6|LNC|Bone Scan W SM153 IV|Bone Scan W SM153 IV
C2826012|T102|strict|39666-3|LNC|Heart Scan W stress and W 201 Th IV|Heart Scan W stress and W 201 Th IV
C2826012|T102|strict|39667-1|LNC|Heart Scan W stress and W radionuclide IV|Heart Scan W stress and W radionuclide IV
C2826012|T102|strict|69231-9|LNC|Heart Scan W stress and W Tc-99m IV|Heart Scan W stress and W Tc-99m IV
C2826012|T102|strict|69232-7|LNC|Heart Scan W stress and W Tc-99m Sestamibi IV|Heart Scan W stress and W Tc-99m Sestamibi IV
C2826012|T102|strict|24819-5|LNC|Liver and Spleen Scan W Tc-99m calcium colloid IV|Liver and Spleen Scan W Tc-99m calcium colloid IV
C2826012|T102|strict|39744-8|LNC|Prostate Scan W Tc-99m capromab pendatide IV|Prostate Scan W Tc-99m capromab pendatide IV
C2826012|T102|strict|39674-7|LNC|Gallbladder Scan W Tc-99m DISIDA IV|Gallbladder Scan W Tc-99m DISIDA IV
C2826012|T102|strict|41771-7|LNC|Kidney - bilateral Scan W Tc-99m DMSA IV|Kidney - bilateral Scan W Tc-99m DMSA IV
C2826012|T102|strict|39625-9|LNC|Artery Scan W Tc-99m DTPA IA|Artery Scan W Tc-99m DTPA IA
C2826012|T102|strict|39745-5|LNC|Kidney - bilateral Scan W Tc-99m DTPA IV|Kidney - bilateral Scan W Tc-99m DTPA IV
C2826012|T102|strict|43667-5|LNC|Kidney - bilateral and Renal vessels Scan W Tc-99m DTPA IV|Kidney - bilateral and Renal vessels Scan W Tc-99m DTPA IV
C2826012|T102|strict|39753-9|LNC|Scrotum and Testicle Scan W Tc-99m DTPA IV|Scrotum and Testicle Scan W Tc-99m DTPA IV
C2826012|T102|strict|39765-3|LNC|Vein Scan W Tc-99m DTPA IV|Vein Scan W Tc-99m DTPA IV
C2826012|T102|strict|39642-4|LNC|Brain Scan W Tc-99m glucoheptonate IV|Brain Scan W Tc-99m glucoheptonate IV
C2826012|T102|strict|44234-3|LNC|Kidney - bilateral Scan W Tc-99m glucoheptonate IV|Kidney - bilateral Scan W Tc-99m glucoheptonate IV
C2826012|T102|strict|39766-1|LNC|Vein Scan W Tc-99m HDP IV|Vein Scan W Tc-99m HDP IV
C2826012|T102|strict|39812-3|LNC|Bone Scan W Tc-99m HMPAO IV|Bone Scan W Tc-99m HMPAO IV
C2826012|T102|strict|39630-9|LNC|Brain Scan W Tc-99m HMPAO IV|Brain Scan W Tc-99m HMPAO IV
C2826012|T102|strict|39757-0|LNC|Thyroid Scan W Tc-99m IV|Thyroid Scan W Tc-99m IV
C2826012|T102|strict|24831-0|LNC|Meckels diverticulum Scan W Tc-99m M04 IV|Meckels diverticulum Scan W Tc-99m M04 IV
C2826012|T102|strict|44141-0|LNC|Liver and Spleen Scan W Tc-99m MAA IV|Liver and Spleen Scan W Tc-99m MAA IV
C2826012|T102|strict|44142-8|LNC|Bone Scan W Tc-99m medronate IV|Bone Scan W Tc-99m medronate IV
C2826012|T102|strict|39746-3|LNC|Kidney - bilateral Scan W Tc-99m Mertiatide IV|Kidney - bilateral Scan W Tc-99m Mertiatide IV
C2826012|T102|strict|69233-5|LNC|Parotid gland Scan W Tc-99m pertechnetate IV|Parotid gland Scan W Tc-99m pertechnetate IV
C2826012|T102|strict|25001-9|LNC|Scrotum and Testicle Scan W Tc-99m pertechnetate IV|Scrotum and Testicle Scan W Tc-99m pertechnetate IV
C2826012|T102|strict|26091-9|LNC|Scrotum and Testicle - bilateral Scan W Tc-99m pertechnetate IV|Scrotum and Testicle - bilateral Scan W Tc-99m pertechnetate IV
C2826012|T102|strict|26092-7|LNC|Scrotum and Testicle - left Scan W Tc-99m pertechnetate IV|Scrotum and Testicle - left Scan W Tc-99m pertechnetate IV
C2826012|T102|strict|26093-5|LNC|Scrotum and Testicle - right Scan W Tc-99m pertechnetate IV|Scrotum and Testicle - right Scan W Tc-99m pertechnetate IV
C2826012|T102|strict|44146-9|LNC|Bone marrow Scan W Tc-99m SC IV|Bone marrow Scan W Tc-99m SC IV
C2826012|T102|strict|39689-5|LNC|Gastrointestine Scan W Tc-99m SC IV|Gastrointestine Scan W Tc-99m SC IV
C2826012|T102|strict|69230-1|LNC|Liver Scan W Tc-99m SC IV|Liver Scan W Tc-99m SC IV
C2826012|T102|strict|39764-6|LNC|Vein Scan W Tc-99m SC IV|Vein Scan W Tc-99m SC IV
C2826012|T102|strict|24683-5|LNC|Esophagus and Stomach Scan W Tc-99m SC PO|Esophagus and Stomach Scan W Tc-99m SC PO
C2826012|T102|strict|44145-1|LNC|Parathyroid Scan W Tc-99m Sestamibi IV|Parathyroid Scan W Tc-99m Sestamibi IV
C2826012|T102|strict|39756-2|LNC|Thyroid Scan W Tc-99m Sestamibi IV|Thyroid Scan W Tc-99m Sestamibi IV
C2826012|T102|strict|24714-8|LNC|Gastrointestine Scan W Tc-99m tagged RBC IV|Gastrointestine Scan W Tc-99m tagged RBC IV
C2826012|T102|strict|44143-6|LNC|Heart Scan W Tc-99m tagged RBC IV|Heart Scan W Tc-99m tagged RBC IV
C2826012|T102|strict|39690-3|LNC|Liver Scan W Tc-99m tagged RBC IV|Liver Scan W Tc-99m tagged RBC IV
C2826012|T102|strict|42700-5|LNC|Bone Scan W Tc-99m tagged WBC IV|Bone Scan W Tc-99m tagged WBC IV
C2826012|T102|strict|24751-0|LNC|Parathyroid Scan W TI-201 subtraction Tc-99m IV|Parathyroid Scan W TI-201 subtraction Tc-99m IV
C2826012|T102|strict|39635-8|LNC|Brain Scan W Tl-201 IV|Brain Scan W Tl-201 IV
C2826012|T102|strict|51389-5|LNC|Breast Scan W Tl-201 IV|Breast Scan W Tl-201 IV
C2826012|T102|strict|42012-5|LNC|Gastrointestine upper Fluoroscopy W water soluble contrast PO|Gastrointestine upper Fluoroscopy W water soluble contrast PO
C2826012|T102|strict|24669-4|LNC|Colon Fluoroscopy W water soluble contrast PR|Colon Fluoroscopy W water soluble contrast PR
C2826012|T102|strict|37577-4|LNC|Acromioclavicular Joint X-ray W weight|Acromioclavicular Joint X-ray W weight
C2826012|T102|strict|37578-2|LNC|Acromioclavicular joint - bilateral X-ray W weight|Acromioclavicular joint - bilateral X-ray W weight
C2826012|T102|strict|44144-4|LNC|Liver Scan W Xe-133 inhaled|Liver Scan W Xe-133 inhaled
C2826012|T102|strict|37582-4|LNC|Acromioclavicular Joint X-ray WO weight|Acromioclavicular Joint X-ray WO weight
C2826012|T102|strict|69055-2|LNC|Acromioclavicular joint - bilateral X-ray WO weight|Acromioclavicular joint - bilateral X-ray WO weight
C2826012|T102|strict|52073-4|LNC|Vision attachment|Vision attachment
C2826012|T102|strict|28631-0|LNC|Visual acuity study|Visual acuity study
C2826012|T102|strict|46242-4|LNC|Fetal Document Vital signs measurements|Fetal Document Vital signs measurements
C2826012|T102|strict|52070-0|LNC|Workers compensation|Workers compensation
C2826012|T102|strict|74282-5|LNC|Individual counseling note|Individual counseling note
C2826012|T102|strict|71683-7|LNC|FDA package insert PMI - Stop taking and call your doctor section|FDA package insert PMI - Stop taking and call your doctor section
C2826012|T102|strict|71685-2|LNC|FDA package insert PMI - Tell your doctor before taking section|FDA package insert PMI - Tell your doctor before taking section
C2826012|T102|strict|34086-9|LNC|FDA package insert Abuse section|FDA package insert Abuse section
C2826012|T102|strict|60555-0|LNC|FDA package insert Accessories|FDA package insert Accessories
C2826012|T102|strict|34084-4|LNC|FDA package insert Adverse reactions section|FDA package insert Adverse reactions section
C2826012|T102|strict|69761-5|LNC|FDA package insert Alarms|FDA package insert Alarms
C2826012|T102|strict|70946-9|LNC|Ancillary eye tests Narrative|Ancillary eye tests Narrative
C2826012|T102|strict|34091-9|LNC|FDA package insert Animal pharmacology/toxicology section|FDA package insert Animal pharmacology/toxicology section
C2826012|T102|strict|48767-8|LNC|Annotation comment Narrative|Annotation comment Narrative
C2826012|T102|strict|60556-8|LNC|FDA package insert Assembly or installation instructions|FDA package insert Assembly or installation instructions
C2826012|T102|strict|35519-8|LNC|Clinical trial protocol Assessment of safety section|Clinical trial protocol Assessment of safety section
C2826012|T102|strict|35517-2|LNC|Clinical trial protocol Assessment section|Clinical trial protocol Assessment section
C2826012|T102|strict|35511-5|LNC|Clinical trial protocol Background information section|Clinical trial protocol Background information section
C2826012|T102|strict|34066-1|LNC|FDA package insert Boxed warning section|FDA package insert Boxed warning section
C2826012|T102|strict|60557-6|LNC|FDA package insert Calibration instructions|FDA package insert Calibration instructions
C2826012|T102|strict|72135-7|LNC|Cancer diagnosis Narrative|Cancer diagnosis Narrative
C2826012|T102|strict|34083-6|LNC|FDA package insert Carcinogenesis and mutagenesis and impairment of fertility section|FDA package insert Carcinogenesis and mutagenesis and impairment of fertility section
C2826012|T102|strict|60684-8|LNC|FDA product label Cellular therapy|FDA product label Cellular therapy
C2826012|T102|strict|60558-4|LNC|FDA package insert Cleaning, disinfecting, and sterilization instructions|FDA package insert Cleaning, disinfecting, and sterilization instructions
C2826012|T102|strict|34090-1|LNC|FDA package insert Clinical pharmacology section|FDA package insert Clinical pharmacology section
C2826012|T102|strict|34092-7|LNC|FDA package insert Clinical studies section|FDA package insert Clinical studies section
C2826012|T102|strict|35528-9|LNC|Clinical trial protocol Clinical trial protocol|Clinical trial protocol Clinical trial protocol
C2826012|T102|strict|69760-7|LNC|FDA package insert Compatible accessories|FDA package insert Compatible accessories
C2826012|T102|strict|60559-2|LNC|FDA package insert Components|FDA package insert Components
C2826012|T102|strict|70940-2|LNC|Confrontation visual field Narrative|Confrontation visual field Narrative
C2826012|T102|strict|34070-3|LNC|FDA package insert Contraindications section|FDA package insert Contraindications section
C2826012|T102|strict|34085-1|LNC|FDA package insert Controlled substance section|FDA package insert Controlled substance section
C2826012|T102|strict|57826-0|LNC|Co-payment amount Narrative|Co-payment amount Narrative
C2826012|T102|strict|57025-9|LNC|Data criteria Narrative|Data criteria Narrative
C2826012|T102|strict|35524-8|LNC|Clinical trial protocol Data handling and record keeping section|Clinical trial protocol Data handling and record keeping section
C2826012|T102|strict|34087-7|LNC|FDA package insert Dependence section|FDA package insert Dependence section
C2826012|T102|strict|34089-3|LNC|FDA package insert Description section|FDA package insert Description section
C2826012|T102|strict|69758-1|LNC|FDA package insert Diagram of device|FDA package insert Diagram of device
C2826012|T102|strict|35521-4|LNC|Clinical trial protocol Direct access to source data+documents section|Clinical trial protocol Direct access to source data+documents section
C2826012|T102|strict|69763-1|LNC|FDA package insert Disposal and waste handling|FDA package insert Disposal and waste handling
C2826012|T102|strict|34068-7|LNC|FDA package insert Dosage and administration section|FDA package insert Dosage and administration section
C2826012|T102|strict|43678-2|LNC|FDA package insert Dosage forms and strengths section|FDA package insert Dosage forms and strengths section
C2826012|T102|strict|34074-5|LNC|FDA package insert Drug/laboratory test interactions section|FDA package insert Drug/laboratory test interactions section
C2826012|T102|strict|42227-9|LNC|FDA package insert Drug abuse and dependence section|FDA package insert Drug abuse and dependence section
C2826012|T102|strict|34073-7|LNC|FDA package insert Drug interactions section|FDA package insert Drug interactions section
C2826012|T102|strict|35518-0|LNC|Clinical trial protocol Efficacy assessment section|Clinical trial protocol Efficacy assessment section
C2826012|T102|strict|35523-0|LNC|Clinical trial protocol Ethics section|Clinical trial protocol Ethics section
C2826012|T102|strict|61147-5|LNC|Expected outcomes Narrative|Expected outcomes Narrative
C2826012|T102|strict|70943-6|LNC|Eye anterior segment Narrative|Eye anterior segment Narrative
C2826012|T102|strict|70941-0|LNC|Eye external Narrative|Eye external Narrative
C2826012|T102|strict|70944-4|LNC|Eye posterior segment Narrative|Eye posterior segment Narrative
C2826012|T102|strict|35525-5|LNC|Clinical trial protocol Financing and insurance section|Clinical trial protocol Financing and insurance section
C2826012|T102|strict|35510-7|LNC|Clinical trial protocol General information section|Clinical trial protocol General information section
C2826012|T102|strict|34072-9|LNC|FDA package insert General precautions section|FDA package insert General precautions section
C2826012|T102|strict|71743-9|LNC|FDA product label Generic drug facility identification submission|FDA product label Generic drug facility identification submission
C2826012|T102|strict|34082-8|LNC|FDA package insert Geriatric use section|FDA package insert Geriatric use section
C2826012|T102|strict|61146-7|LNC|Goals Narrative|Goals Narrative
C2826012|T102|strict|71744-7|LNC|FDA package insert Health care provider letter|FDA package insert Health care provider letter
C2826012|T102|strict|69719-3|LNC|FDA product label Health claim section|FDA product label Health claim section
C2826012|T102|strict|69670-8|LNC|Health quality measure supplemental data Narrative|Health quality measure supplemental data Narrative
C2826012|T102|strict|34069-5|LNC|FDA package insert How supplied section|FDA package insert How supplied section
C2826012|T102|strict|72090-4|LNC|FDA product label Identification of CBER-regulated generic drug facility|FDA product label Identification of CBER-regulated generic drug facility
C2826012|T102|strict|64123-3|LNC|FDA package insert Indexing - adverse reaction|FDA package insert Indexing - adverse reaction
C2826012|T102|strict|71446-9|LNC|FDA package insert Indexing - billing unit|FDA package insert Indexing - billing unit
C2826012|T102|strict|60685-5|LNC|FDA package insert Indexing - pharmacologic class|FDA package insert Indexing - pharmacologic class
C2826012|T102|strict|73815-3|LNC|FDA package insert Indexing - product concept|FDA package insert Indexing - product concept
C2826012|T102|strict|64124-1|LNC|FDA package insert Indexing - substance|FDA package insert Indexing - substance
C2826012|T102|strict|34067-9|LNC|FDA package insert Indications and usage section|FDA package insert Indications and usage section
C2826012|T102|strict|34076-0|LNC|FDA package insert Information for patients section|FDA package insert Information for patients section
C2826012|T102|strict|69730-0|LNC|Instructions [Text] Narrative|Instructions [Text] Narrative
C2826012|T102|strict|59845-8|LNC|FDA package insert Instructions for use section|FDA package insert Instructions for use section
C2826012|T102|strict|60560-0|LNC|FDA package insert Intended use of the device|FDA package insert Intended use of the device
C2826012|T102|strict|62387-6|LNC|Interventions Narrative|Interventions Narrative
C2826012|T102|strict|34079-4|LNC|FDA package insert Labor and delivery section|FDA package insert Labor and delivery section
C2826012|T102|strict|34075-2|LNC|FDA package insert Laboratory tests section|FDA package insert Laboratory tests section
C2826012|T102|strict|70945-1|LNC|Lacrimal Narrative|Lacrimal Narrative
C2826012|T102|strict|70939-4|LNC|Lensometry measurements Narrative|Lensometry measurements Narrative
C2826012|T102|strict|66105-8|LNC|FDA package insert Lot distribution data|FDA package insert Lot distribution data
C2826012|T102|strict|74045-6|LNC|Measure description Narrative|Measure description Narrative
C2826012|T102|strict|57027-5|LNC|Measure observations Narrative|Measure observations Narrative
C2826012|T102|strict|43679-0|LNC|FDA package insert Mechanism of action section|FDA package insert Mechanism of action section
C2826012|T102|strict|49489-8|LNC|FDA package insert Microbiology section|FDA package insert Microbiology section
C2826012|T102|strict|43680-8|LNC|FDA package insert Nonclinical toxicology section|FDA package insert Nonclinical toxicology section
C2826012|T102|strict|34078-6|LNC|FDA package insert Nonteratogenic effects section|FDA package insert Nonteratogenic effects section
C2826012|T102|strict|34080-2|LNC|FDA package insert Nursing mothers section|FDA package insert Nursing mothers section
C2826012|T102|strict|61149-1|LNC|Objective Narrative|Objective Narrative
C2826012|T102|strict|70942-8|LNC|Ocular alignment and motility Narrative|Ocular alignment and motility Narrative
C2826012|T102|strict|70934-5|LNC|Ocular history Narrative|Ocular history Narrative
C2826012|T102|strict|70948-5|LNC|Ocular physical exam Narrative|Ocular physical exam Narrative
C2826012|T102|strict|70935-2|LNC|Ophthalmic medications Narrative|Ophthalmic medications Narrative
C2826012|T102|strict|60561-8|LNC|FDA package insert Other safety information|FDA package insert Other safety information
C2826012|T102|strict|34088-5|LNC|FDA package insert Overdosage section|FDA package insert Overdosage section
C2826012|T102|strict|51941-3|LNC|FDA product label Back panel of package|FDA product label Back panel of package
C2826012|T102|strict|51947-0|LNC|FDA product label Bottom panel of package|FDA product label Bottom panel of package
C2826012|T102|strict|51948-8|LNC|FDA product label Flap panel of package|FDA product label Flap panel of package
C2826012|T102|strict|51945-4|LNC|FDA product label Principal display panel of package|FDA product label Principal display panel of package
C2826012|T102|strict|51944-7|LNC|FDA product label Side panel of package|FDA product label Side panel of package
C2826012|T102|strict|51943-9|LNC|FDA product label Side panel of package Left|FDA product label Side panel of package Left
C2826012|T102|strict|51942-1|LNC|FDA product label Side panel of package Right|FDA product label Side panel of package Right
C2826012|T102|strict|51946-2|LNC|FDA product label Top panel of package|FDA product label Top panel of package
C2826012|T102|strict|34081-0|LNC|FDA package insert Pediatric use section|FDA package insert Pediatric use section
C2826012|T102|strict|43681-6|LNC|FDA package insert Pharmacodynamics section|FDA package insert Pharmacodynamics section
C2826012|T102|strict|66106-6|LNC|FDA package insert Pharmacogenomics section|FDA package insert Pharmacogenomics section
C2826012|T102|strict|43682-4|LNC|FDA package insert Pharmacokinetics section|FDA package insert Pharmacokinetics section
C2826012|T102|strict|59772-4|LNC|Planned procedure Narrative|Planned procedure Narrative
C2826012|T102|strict|60683-0|LNC|FDA product label Plasma derivative|FDA product label Plasma derivative
C2826012|T102|strict|71681-1|LNC|FDA package insert PMI - Common side effects section|FDA package insert PMI - Common side effects section
C2826012|T102|strict|71684-5|LNC|FDA package insert PMI - Directions for use section|FDA package insert PMI - Directions for use section
C2826012|T102|strict|71686-0|LNC|FDA package insert PMI - Do not take section|FDA package insert PMI - Do not take section
C2826012|T102|strict|71682-9|LNC|FDA package insert PMI - Get emergency medical help section|FDA package insert PMI - Get emergency medical help section
C2826012|T102|strict|71687-8|LNC|FDA package insert PMI - Important information section|FDA package insert PMI - Important information section
C2826012|T102|strict|71688-6|LNC|FDA package insert PMI - Uses section|FDA package insert PMI - Uses section
C2826012|T102|strict|57026-7|LNC|Population criteria Narrative|Population criteria Narrative
C2826012|T102|strict|69669-0|LNC|Population stratification description Narrative|Population stratification description Narrative
C2826012|T102|strict|59769-0|LNC|Postprocedure diagnosis Narrative|Postprocedure diagnosis Narrative
C2826012|T102|strict|42232-9|LNC|FDA package insert Precautions section|FDA package insert Precautions section
C2826012|T102|strict|42228-7|LNC|FDA package insert Pregnancy section|FDA package insert Pregnancy section
C2826012|T102|strict|57059-8|LNC|Pregnancy visit summary note Narrative|Pregnancy visit summary note Narrative
C2826012|T102|strict|59774-0|LNC|Procedure anesthesia Narrative|Procedure anesthesia Narrative
C2826012|T102|strict|59775-7|LNC|Procedure disposition Narrative|Procedure disposition Narrative
C2826012|T102|strict|59770-8|LNC|Procedure estimated blood loss Narrative|Procedure estimated blood loss Narrative
C2826012|T102|strict|59776-5|LNC|Procedure findings Narrative|Procedure findings Narrative
C2826012|T102|strict|59771-6|LNC|Procedure implants Narrative|Procedure implants Narrative
C2826012|T102|strict|59768-2|LNC|Procedure indications Narrative|Procedure indications Narrative
C2826012|T102|strict|59773-2|LNC|Procedure specimens taken Narrative|Procedure specimens taken Narrative
C2826012|T102|strict|35526-3|LNC|Clinical trial protocol Publication policy section|Clinical trial protocol Publication policy section
C2826012|T102|strict|35522-2|LNC|Clinical trial protocol Quality control and quality assurance section|Clinical trial protocol Quality control and quality assurance section
C2826012|T102|strict|57827-8|LNC|Reason for co-payment exemption Narrative|Reason for co-payment exemption Narrative
C2826012|T102|strict|43683-2|LNC|FDA package insert Recent major changes section|FDA package insert Recent major changes section
C2826012|T102|strict|34093-5|LNC|FDA package insert References section|FDA package insert References section
C2826012|T102|strict|70938-6|LNC|Refractive measurements Narrative|Refractive measurements Narrative
C2826012|T102|strict|69759-9|LNC|FDA package insert Risks|FDA package insert Risks
C2826012|T102|strict|48779-3|LNC|FDA package insert Structured product labelling indexing data elements section|FDA package insert Structured product labelling indexing data elements section
C2826012|T102|strict|48780-1|LNC|FDA package insert Structured product labelling listing data elements section|FDA package insert Structured product labelling listing data elements section
C2826012|T102|strict|42231-1|LNC|FDA package insert Structured product labelling medguide section|FDA package insert Structured product labelling medguide section
C2826012|T102|strict|42230-3|LNC|FDA package insert Structured product laballing patient package insert section|FDA package insert Structured product laballing patient package insert section
C2826012|T102|strict|38056-8|LNC|FDA package insert Structured product laballing supplemental patient material|FDA package insert Structured product laballing supplemental patient material
C2826012|T102|strict|42229-5|LNC|FDA package insert Structured patient labelling unclassified section|FDA package insert Structured patient labelling unclassified section
C2826012|T102|strict|69718-5|LNC|FDA product label Statement of identity section|FDA product label Statement of identity section
C2826012|T102|strict|35520-6|LNC|Clinical trial protocol Statistics section|Clinical trial protocol Statistics section
C2826012|T102|strict|44425-7|LNC|FDA package insert Storage and handling section|FDA package insert Storage and handling section
C2826012|T102|strict|35515-6|LNC|Clinical trial protocol Subject participation + epochs section|Clinical trial protocol Subject participation + epochs section
C2826012|T102|strict|35514-9|LNC|Clinical trial protocol Subject selection and withdrawal section|Clinical trial protocol Subject selection and withdrawal section
C2826012|T102|strict|61150-9|LNC|Subjective Narrative|Subjective Narrative
C2826012|T102|strict|35527-1|LNC|Clinical trial protocol Supplements section|Clinical trial protocol Supplements section
C2826012|T102|strict|55122-6|LNC|Surgical operation note implants Narrative|Surgical operation note implants Narrative
C2826012|T102|strict|34077-8|LNC|FDA package insert Teratogenic effects section|FDA package insert Teratogenic effects section
C2826012|T102|strict|35516-4|LNC|Clinical trial protocol Treatment of subjects + epochs section|Clinical trial protocol Treatment of subjects + epochs section
C2826012|T102|strict|35513-1|LNC|Clinical trial protocol Trial design section|Clinical trial protocol Trial design section
C2826012|T102|strict|42796-3|LNC|Clinical trial protocol Trial name|Clinical trial protocol Trial name
C2826012|T102|strict|35512-3|LNC|Clinical trial protocol Trial objectives and purpose section|Clinical trial protocol Trial objectives and purpose section
C2826012|T102|strict|69762-3|LNC|FDA package insert Troubleshooting|FDA package insert Troubleshooting
C2826012|T102|strict|43684-0|LNC|FDA package insert Use in specific populations section|FDA package insert Use in specific populations section
C2826012|T102|strict|54433-8|LNC|FDA package insert User safety warnings section|FDA package insert User safety warnings section
C2826012|T102|strict|70936-0|LNC|Vision testing Narrative|Vision testing Narrative
C2826012|T102|strict|43685-7|LNC|FDA package insert Warnings and precautions section|FDA package insert Warnings and precautions section
C2826012|T102|strict|34071-1|LNC|FDA package insert Warnings section|FDA package insert Warnings section
C2826012|T102|strict|74477-1|LNC|Clinical document Kind of document from LOINC Document Ontology|Clinical document Kind of document from LOINC Document Ontology
C2826012|T102|strict|74479-7|LNC|Clinical document Role from LOINC Document Ontology|Clinical document Role from LOINC Document Ontology
C2826012|T102|strict|74476-3|LNC|Clinical document Setting from LOINC Document Ontology|Clinical document Setting from LOINC Document Ontology
C2826012|T102|strict|74480-5|LNC|Clinical document Subject matter domain from LOINC Document Ontology|Clinical document Subject matter domain from LOINC Document Ontology
C2826012|T102|strict|74478-9|LNC|Clinical document Type of service from LOINC Document Ontology|Clinical document Type of service from LOINC Document Ontology
C2826012|T102|strict|42566-0|LNC|Contributing Factor communication/Documentation MERSTH|Contributing Factor communication/Documentation MERSTH
C2826012|T102|strict|21862-8|LNC|Source of document used to abstract Cancer|Source of document used to abstract Cancer
C2826012|T102|strict|69764-9|LNC|Document type|Document type
C2826012|T102|strict|48766-0|LNC|Information source|Information source
C2826012|T102|strict|70949-3|LNC|Pathology report.section heading|Pathology report.section heading
C2826012|T102|strict|60572-5|LNC|Report template ID|Report template ID
C2826012|T102|strict|60573-3|LNC|Report template source|Report template source
C2826012|T102|strict|60574-1|LNC|Report template version ID|Report template version ID
C2826012|T102|strict|73983-9|LNC|Report.section heading Unspecified body region|Report.section heading Unspecified body region
C2826012|T102|strict|40811-2|LNC|11-Deoxycorticosterone [Presence] in Serum or Plasma|11-Deoxycorticosterone [Presence] in Serum or Plasma
C2826012|T102|strict|29112-0|LNC|Photo documentation Eye - left|Photo documentation Eye - left
C2826012|T102|strict|29111-2|LNC|Photo documentation Eye - right|Photo documentation Eye - right
C2826012|T102|strict|72169-6|LNC|Permission to release immunization data from school record|Permission to release immunization data from school record
C2826012|T102|strict|44943-9|LNC|Self management|Self management
C2826012|T102|strict|11206-0|LNC|18-Hydroxydeoxycorticosterone [Mass/volume] in Serum or Plasma|18-Hydroxydeoxycorticosterone [Mass/volume] in Serum or Plasma
C2826012|T102|strict|26988-6|LNC|18-Hydroxydeoxycorticosterone [Mass/time] in 24 hour Urine|18-Hydroxydeoxycorticosterone [Mass/time] in 24 hour Urine
C2826012|T102|strict|50081-9|LNC|18-Hydroxydeoxycorticosterone [Moles/volume] in Serum or Plasma|18-Hydroxydeoxycorticosterone [Moles/volume] in Serum or Plasma
C2826012|T102|strict|57553-0|LNC|18-Hydroxydeoxycorticosterone [Moles/volume] in Serum or Plasma --1 hour post dose corticotropin|18-Hydroxydeoxycorticosterone [Moles/volume] in Serum or Plasma --1 hour post dose corticotropin
C2826012|T102|strict|57552-2|LNC|18-Hydroxydeoxycorticosterone [Moles/volume] in Serum or Plasma --30 minutes post dose corticotropin|18-Hydroxydeoxycorticosterone [Moles/volume] in Serum or Plasma --30 minutes post dose corticotropin
C2826012|T102|strict|57551-4|LNC|18-Hydroxydeoxycorticosterone [Moles/volume] in Serum or Plasma --pre dose corticotropin|18-Hydroxydeoxycorticosterone [Moles/volume] in Serum or Plasma --pre dose corticotropin
C2826012|T102|strict|53347-1|LNC|11-Deoxycorticosterone [Mass/volume] in Dried blood spot|11-Deoxycorticosterone [Mass/volume] in Dried blood spot
C2826012|T102|strict|1656-8|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma
C2826012|T102|strict|42855-7|LNC|11-Deoxycorticosterone [Mass/volume] in Urine|11-Deoxycorticosterone [Mass/volume] in Urine
C2826012|T102|strict|16110-9|LNC|11-Deoxycorticosterone [Mass/time] in 24 hour Urine|11-Deoxycorticosterone [Mass/time] in 24 hour Urine
C2826012|T102|strict|40818-7|LNC|11-Deoxycorticosterone [Moles/volume] in 24 hour Urine|11-Deoxycorticosterone [Moles/volume] in 24 hour Urine
C2826012|T102|strict|53348-9|LNC|11-Deoxycorticosterone [Moles/volume] in Dried blood spot|11-Deoxycorticosterone [Moles/volume] in Dried blood spot
C2826012|T102|strict|25561-2|LNC|11-Deoxycorticosterone [Moles/volume] in Serum or Plasma|11-Deoxycorticosterone [Moles/volume] in Serum or Plasma
C2826012|T102|strict|55808-0|LNC|11-Deoxycorticosterone [Moles/time] in 24 hour Urine|11-Deoxycorticosterone [Moles/time] in 24 hour Urine
C2826012|T102|strict|56611-7|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --1.5 hours post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --1.5 hours post XXX challenge
C2826012|T102|strict|56608-3|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --15 minutes post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --15 minutes post XXX challenge
C2826012|T102|strict|57493-9|LNC|11-Deoxycorticosterone [Moles/volume] in Serum or Plasma --1 hour post 250 ug corticotropin|11-Deoxycorticosterone [Moles/volume] in Serum or Plasma --1 hour post 250 ug corticotropin
C2826012|T102|strict|40816-1|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --1 hour post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --1 hour post XXX challenge
C2826012|T102|strict|56602-6|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --1st specimen post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --1st specimen post XXX challenge
C2826012|T102|strict|56613-3|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --2.5 hours post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --2.5 hours post XXX challenge
C2826012|T102|strict|56609-1|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --20 minutes post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --20 minutes post XXX challenge
C2826012|T102|strict|56612-5|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --2 hours post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --2 hours post XXX challenge
C2826012|T102|strict|56603-4|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --2nd specimen post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --2nd specimen post XXX challenge
C2826012|T102|strict|57492-1|LNC|11-Deoxycorticosterone [Moles/volume] in Serum or Plasma --30 minutes post 250 ug corticotropin|11-Deoxycorticosterone [Moles/volume] in Serum or Plasma --30 minutes post 250 ug corticotropin
C2826012|T102|strict|56556-4|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --30 minutes post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --30 minutes post XXX challenge
C2826012|T102|strict|56604-2|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --3rd specimen post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --3rd specimen post XXX challenge
C2826012|T102|strict|56610-9|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --40 minutes post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --40 minutes post XXX challenge
C2826012|T102|strict|56605-9|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --4th specimen post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --4th specimen post XXX challenge
C2826012|T102|strict|59987-8|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --5th specimen post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --5th specimen post XXX challenge
C2826012|T102|strict|59986-0|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --6th specimen post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --6th specimen post XXX challenge
C2826012|T102|strict|59985-2|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --7th specimen post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --7th specimen post XXX challenge
C2826012|T102|strict|59984-5|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --8th specimen post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --8th specimen post XXX challenge
C2826012|T102|strict|56555-6|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --baseline|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --baseline
C2826012|T102|strict|16294-1|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --post XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --post XXX challenge
C2826012|T102|strict|57491-3|LNC|11-Deoxycorticosterone [Moles/volume] in Serum or Plasma --pre 250 ug corticotropin|11-Deoxycorticosterone [Moles/volume] in Serum or Plasma --pre 250 ug corticotropin
C2826012|T102|strict|56606-7|LNC|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --pre XXX challenge|11-Deoxycorticosterone [Mass/volume] in Serum or Plasma --pre XXX challenge
C2826012|T102|strict|13480-9|LNC|18-Hydroxydeoxycortisol/Creatinine [Mass Ratio] in Urine|18-Hydroxydeoxycortisol/Creatinine [Mass Ratio] in Urine
C2826012|T102|strict|44729-2|LNC|Progesterone/11-Deoxycorticosterone [Mass Ratio] in Serum or Plasma|Progesterone/11-Deoxycorticosterone [Mass Ratio] in Serum or Plasma
C2826012|T102|strict|69799-5|LNC|21-Deoxycorticosterone [Moles/volume] in Serum or Plasma|21-Deoxycorticosterone [Moles/volume] in Serum or Plasma
C2826012|T102|strict|57562-1|LNC|21-Deoxycorticosterone [Moles/volume] in Serum or Plasma --1 hour post dose corticotropin|21-Deoxycorticosterone [Moles/volume] in Serum or Plasma --1 hour post dose corticotropin
C2826012|T102|strict|57561-3|LNC|21-Deoxycorticosterone [Moles/volume] in Serum or Plasma --30 minutes post dose corticotropin|21-Deoxycorticosterone [Moles/volume] in Serum or Plasma --30 minutes post dose corticotropin
C2826012|T102|strict|57560-5|LNC|21-Deoxycorticosterone [Moles/volume] in Serum or Plasma --pre dose corticotropin|21-Deoxycorticosterone [Moles/volume] in Serum or Plasma --pre dose corticotropin
C2826012|T102|strict|72510-1|LNC|Performance rate Reporting period population Calculated|Performance rate Reporting period population Calculated
C2826012|T102|strict|72509-3|LNC|Reporting rate Reporting period population Calculated|Reporting rate Reporting period population Calculated
C1547726|T102|strict|82242000|LNC|Hospital-children's|Hospital-children's
C1547726|T102|strict|225732001|LNC|Hospital-community|Hospital-community
C1547726|T102|strict|79993009|LNC|Hospital-government|Hospital-government
C1547726|T102|strict|32074000|LNC|Hospital-long term care|Hospital-long term care
C1547726|T102|strict|4322002|LNC|Hospital-military field|Hospital-military field
C1547726|T102|strict|224687002|LNC|Hospital-prison|Hospital-prison
C1547726|T102|strict|62480006|LNC|Hospital-psychiatric|Hospital-psychiatric
C1547726|T102|strict|80522000|LNC|Hospital-rehabilitation|Hospital-rehabilitation
C1547726|T102|strict|36125001|LNC|Hospital-trauma center|Hospital-trauma center
C1547726|T102|strict|48311003|LNC|Hospital-Veterans' Administration|Hospital-Veterans' Administration
C1547726|T102|strict|284546000|LNC|Hospice facility|Hospice facility
C1547726|T102|strict|42665001|LNC|Nursing home|Nursing home
C1547726|T102|strict|45618002|LNC|Skilled nursing facility|Skilled nursing facility
C1547726|T102|strict|418518002|LNC|Dialysis unit--hospital|Dialysis unit--hospital
C1547726|T102|strict|73770003|LNC|Emergency department--hospital|Emergency department--hospital
C1547726|T102|strict|69362002|LNC|Hospital ambulatory surgery facility|Hospital ambulatory surgery facility
C1547726|T102|strict|52668009|LNC|Hospital birthing center|Hospital birthing center
C1547726|T102|strict|360957003|LNC|Hospital outpatient allergy clinic|Hospital outpatient allergy clinic
C1547726|T102|strict|10206005|LNC|Hospital outpatient dental clinic|Hospital outpatient dental clinic
C1547726|T102|strict|37550003|LNC|Hospital outpatient dermatology clinic|Hospital outpatient dermatology clinic
C1547726|T102|strict|73644007|LNC|Hospital outpatient endocrinology clinic|Hospital outpatient endocrinology clinic
C1547726|T102|strict|31628002|LNC|Hospital outpatient family medicine clinic|Hospital outpatient family medicine clinic
C1547726|T102|strict|58482006|LNC|Hospital outpatient gastroenterology clinic|Hospital outpatient gastroenterology clinic
C1547726|T102|strict|90484001|LNC|Hospital outpatient general surgery clinic|Hospital outpatient general surgery clinic
C1547726|T102|strict|1814000|LNC|Hospital outpatient geriatric health center|Hospital outpatient geriatric health center
C1547726|T102|strict|22549003|LNC|Hospital outpatient gynecology clinic|Hospital outpatient gynecology clinic
C1547726|T102|strict|56293002|LNC|Hospital outpatient hematology clinic|Hospital outpatient hematology clinic
C1547726|T102|strict|360966004|LNC|Hospital outpatient immunology clinic|Hospital outpatient immunology clinic
C1547726|T102|strict|2849009|LNC|Hospital outpatient infectious disease clinic|Hospital outpatient infectious disease clinic
C1547726|T102|strict|14866005|LNC|Hospital outpatient mental health center|Hospital outpatient mental health center
C1547726|T102|strict|38238005|LNC|Hospital outpatient neurology clinic|Hospital outpatient neurology clinic
C1547726|T102|strict|56189001|LNC|Hospital outpatient obstetrical clinic|Hospital outpatient obstetrical clinic
C1547726|T102|strict|89972002|LNC|Hospital outpatient oncology clinic|Hospital outpatient oncology clinic
C1547726|T102|strict|78088001|LNC|Hospital outpatient ophthalmology clinic|Hospital outpatient ophthalmology clinic
C1547726|T102|strict|78001009|LNC|Hospital outpatient orthopedics clinic|Hospital outpatient orthopedics clinic
C1547726|T102|strict|23392004|LNC|Hospital outpatient otorhinolaryngology clinic|Hospital outpatient otorhinolaryngology clinic
C1547726|T102|strict|36293008|LNC|Hospital outpatient pain clinic|Hospital outpatient pain clinic
C1547726|T102|strict|3729002|LNC|Hospital outpatient pediatric clinic|Hospital outpatient pediatric clinic
C1547726|T102|strict|5584006|LNC|Hospital outpatient peripheral vascular clinic|Hospital outpatient peripheral vascular clinic
C1547726|T102|strict|37546005|LNC|Hospital outpatient rehabilitation clinic|Hospital outpatient rehabilitation clinic
C1547726|T102|strict|57159002|LNC|Hospital outpatient respiratory disease clinic|Hospital outpatient respiratory disease clinic
C1547726|T102|strict|331006|LNC|Hospital outpatient rheumatology clinic|Hospital outpatient rheumatology clinic
C1547726|T102|strict|50569004|LNC|Hospital outpatient urology clinic|Hospital outpatient urology clinic
C1547726|T102|strict|79491001|LNC|Hospital radiology facility|Hospital radiology facility
C1547726|T102|strict|33022008|LNC|Hospital-based outpatient clinic or department--OTHER-NOT LISTED|Hospital-based outpatient clinic or department--OTHER-NOT LISTED
C1547726|T102|strict|19602009|LNC|Fee-for-service private physicians' group office|Fee-for-service private physicians' group office
C1547726|T102|strict|39350007|LNC|Private physicians' group office|Private physicians' group office
C1547726|T102|strict|83891005|LNC|Solo practice private office|Solo practice private office
C1547726|T102|strict|394759007|LNC|Independent ambulatory care provider site--OTHER--NOT LISTED|Independent ambulatory care provider site--OTHER--NOT LISTED
C1547726|T102|strict|405607001|LNC|Ambulatory surgery center|Ambulatory surgery center
C1547726|T102|strict|309900005|LNC|Care of the elderly day hospital|Care of the elderly day hospital
C1547726|T102|strict|275576008|LNC|Elderly assessment clinic|Elderly assessment clinic
C1547726|T102|strict|10531005|LNC|Free-standing ambulatory surgery facility|Free-standing ambulatory surgery facility
C1547726|T102|strict|91154008|LNC|Free-standing birthing center|Free-standing birthing center
C1547726|T102|strict|41844007|LNC|Free-standing geriatric health center|Free-standing geriatric health center
C1547726|T102|strict|45899008|LNC|Free-standing laboratory facility|Free-standing laboratory facility
C1547726|T102|strict|51563005|LNC|Free-standing mental health center|Free-standing mental health center
C1547726|T102|strict|1773006|LNC|Free-standing radiology facility|Free-standing radiology facility
C1547726|T102|strict|72311000|LNC|Health maintenance organization|Health maintenance organization
C1547726|T102|strict|6827000|LNC|Local community health center|Local community health center
C1547726|T102|strict|309898008|LNC|Psychogeriatric day hospital|Psychogeriatric day hospital
C1547726|T102|strict|39913001|LNC|Residential school infirmary|Residential school infirmary
C1547726|T102|strict|77931003|LNC|Rural health center|Rural health center
C1547726|T102|strict|25681007|LNC|Sexually transmitted disease health center|Sexually transmitted disease health center
C1547726|T102|strict|20078004|LNC|Substance abuse treatment center|Substance abuse treatment center
C1547726|T102|strict|46224007|LNC|Vaccination clinic|Vaccination clinic
C1547726|T102|strict|81234003|LNC|Walk-in clinic|Walk-in clinic
C1547726|T102|strict|35971002|LNC|Ambulatory care site--OTHER--NOT LISTED|Ambulatory care site--OTHER--NOT LISTED
C1547726|T102|strict|11424001|LNC|Ambulance-based care|Ambulance-based care
C1547726|T102|strict|409519008|LNC|Contained casualty setting|Contained casualty setting
C1547726|T102|strict|901005|LNC|Helicopter-based care|Helicopter-based care
C1547726|T102|strict|2081004|LNC|Hospital ship|Hospital ship
C1547726|T102|strict|59374000|LNC|Traveler's aid clinic|Traveler's aid clinic
C1547726|T102|strict|413456002|LNC|Adult day care center|Adult day care center
C1547726|T102|strict|413817003|LNC|Child day care center|Child day care center
C1547726|T102|strict|310205006|LNC|Private residential home|Private residential home
C1547726|T102|strict|419955002|LNC|Residential institution|Residential institution
C1547726|T102|strict|272501009|LNC|Sports facility|Sports facility
C1547726|T102|strict|394777002|LNC|Health encounter site--NOT LISTED|Health encounter site--NOT LISTED
C1547726|T102|relax|82242000|LNC|children's Hospital|children's Hospital
C1547726|T102|relax|79993009|LNC|government hospital|government hospital
C1547726|T102|relax|32074000|LNC|long term care|long term care
C1547726|T102|relax|4322002|LNC|military Hospital|military Hospital
C1547726|T102|relax|224687002|LNC|Hospital prison|Hospital prison
C1547726|T102|relax|62480006|LNC|psychiatric Hospital|psychiatric Hospital
C1547726|T102|relax|80522000|LNC|rehabilitation Hospital|rehabilitation Hospital
C1547726|T102|relax|36125001|LNC|trauma center|trauma center
C1547726|T102|relax|48311003|LNC|Veterans Administration|Veterans Administration
C1547726|T102|relax|284546000|LNC|Hospice facility|Hospice facility
C1547726|T102|relax|42665001|LNC|Nursing home|Nursing home
C1547726|T102|relax|45618002|LNC|Skilled nursing facility|Skilled nursing facility
C1547726|T102|relax|418518002|LNC|Dialysis unit|Dialysis unit
C1547726|T102|relax|73770003|LNC|Emergency Department|Emergency Department
C1547726|T102|relax|69362002|LNC|surgical facility|surgical facility
C1547726|T102|relax|52668009|LNC|birthing center|birthing center
C1547726|T102|relax|360957003|LNC|allergy clinic|allergy clinic
C1547726|T102|relax|10206005|LNC|dental clinic|dental clinic
C1547726|T102|relax|37550003|LNC|dermatology clinic|dermatology clinic
C1547726|T102|relax|73644007|LNC|endocrinology clinic|endocrinology clinic
C1547726|T102|relax|31628002|LNC|family medicine clinic|family medicine clinic
C1547726|T102|relax|58482006|LNC|gastroenterology clinic|gastroenterology clinic
C1547726|T102|relax|90484001|LNC|general surgery clinic|general surgery clinic
C1547726|T102|relax|1814000|LNC|geriatric health center|geriatric health center
C1547726|T102|relax|22549003|LNC|gynecology clinic|gynecology clinic
C1547726|T102|relax|56293002|LNC|hematology clinic|hematology clinic
C1547726|T102|relax|360966004|LNC|immunology clinic|immunology clinic
C1547726|T102|relax|2849009|LNC|infectious disease clinic|infectious disease clinic
C1547726|T102|relax|14866005|LNC|mental health center|mental health center
C1547726|T102|relax|38238005|LNC|neurology clinic|neurology clinic
C1547726|T102|relax|56189001|LNC|obstetrical clinic|obstetrical clinic
C1547726|T102|relax|89972002|LNC|oncology clinic|oncology clinic
C1547726|T102|relax|78088001|LNC|ophthalmology clinic|ophthalmology clinic
C1547726|T102|relax|78001009|LNC|orthopedics clinic|orthopedics clinic
C1547726|T102|relax|23392004|LNC|otorhinolaryngology clinic|otorhinolaryngology clinic
C1547726|T102|relax|36293008|LNC|pain clinic|pain clinic
C1547726|T102|relax|3729002|LNC|pediatric clinic|pediatric clinic
C1547726|T102|relax|5584006|LNC|peripheral vascular clinic|peripheral vascular clinic
C1547726|T102|relax|37546005|LNC|rehabilitation clinic|rehabilitation clinic
C1547726|T102|relax|57159002|LNC|respiratory disease clinic|respiratory disease clinic
C1547726|T102|relax|331006|LNC|rheumatology clinic|rheumatology clinic
C1547726|T102|relax|50569004|LNC|urology clinic|urology clinic
C1547726|T102|relax|79491001|LNC|Hospital radiology|Hospital radiology
C1547726|T102|relax|33022008|LNC|Hospital outpatient|Hospital outpatient
C1547726|T102|relax|394759007|LNC|Independent ambulatory care provider|Independent ambulatory care provider
C1547726|T102|relax|405607001|LNC|Ambulatory surgery|Ambulatory surgery
C1547726|T102|relax|309900005|LNC|Care of the elderly day hospital|Care of the elderly day hospital
C1547726|T102|relax|275576008|LNC|Elderly assessment clinic|Elderly assessment clinic
C1547726|T102|relax|10531005|LNC|ambulatory surgery facility|ambulatory surgery facility
C1547726|T102|relax|91154008|LNC|birthing center|birthing center
C1547726|T102|relax|41844007|LNC|geriatric health center|geriatric health center
C1547726|T102|relax|45899008|LNC|laboratory facility|laboratory facility
C1547726|T102|relax|51563005|LNC|mental health center|mental health center
C1547726|T102|relax|1773006|LNC|radiology facility|radiology facility
C1547726|T102|relax|72311000|LNC|Health maintenance organization|Health maintenance organization
C1547726|T102|relax|6827000|LNC|Local community health center|Local community health center
C1547726|T102|relax|309898008|LNC|Psychogeriatric day hospital|Psychogeriatric day hospital
C1547726|T102|relax|39913001|LNC|Residential school infirmary|Residential school infirmary
C1547726|T102|relax|77931003|LNC|Rural health center|Rural health center
C1547726|T102|relax|46224007|LNC|Vaccination clinic|Vaccination clinic
C1547726|T102|relax|81234003|LNC|Walk-in clinic|Walk-in clinic
C1547726|T102|relax|35971002|LNC|Ambulatory care site|Ambulatory care site
C1547726|T102|relax|11424001|LNC|Ambulance based care|Ambulance based care
C1547726|T102|relax|409519008|LNC|Contained casualty setting|Contained casualty setting
C1547726|T102|relax|901005|LNC|Care in Helicopter|Care in Helicopter
C1547726|T102|relax|413456002|LNC|Adult day care|Adult day care
C1547726|T102|relax|413817003|LNC|Child day care|Child day care
C1547726|T102|relax|310205006|LNC|residential home|residential home
C1547726|T102|relax|419955002|LNC|Residential|Residential
C1547726|T102|relax|272501009|LNC|Sports facility|Sports facilityC0801762|T102|relax|24754-4|LNC|vasodilator catheter Vein|vasodilator catheter Vein
C0801762|T102|relax|26376-4|LNC|vasodilator catheter Vein bilateral|vasodilator catheter Vein bilateral
C0801762|T102|relax|26377-2|LNC|vasodilator catheter Vein left|vasodilator catheter Vein left
C0801762|T102|relax|26378-0|LNC|vasodilator catheter Vein right|vasodilator catheter Vein right
C0801762|T102|relax|30649-8|LNC|Peripheral artery Fluoroscopic angiogram Additional angioplasty W contrast IA|Peripheral artery Fluoroscopic angiogram Additional angioplasty W contrast IA
C0801762|T102|relax|30641-5|LNC|Vein Fluoroscopic angiogram Additional angioplasty W contrast IV|Vein Fluoroscopic angiogram Additional angioplasty W contrast IV
C0801762|T102|relax|36760-7|LNC|AV shunt Fluoroscopic angiogram Angioplasty W contrast|AV shunt Fluoroscopic angiogram Angioplasty W contrast
C0801762|T102|relax|36762-3|LNC|Extremity vessel Fluoroscopic angiogram Angioplasty W contrast|Extremity vessel Fluoroscopic angiogram Angioplasty W contrast
C0801762|T102|relax|69067-7|LNC|Unspecified body region Fluoroscopic angiogram Angioplasty W contrast|Unspecified body region Fluoroscopic angiogram Angioplasty W contrast
C0801762|T102|relax|24543-1|LNC|Aorta Fluoroscopic angiogram Angioplasty W contrast IA|Aorta Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|24580-3|LNC|Brachiocephalic artery Fluoroscopic angiogram Angioplasty W contrast IA|Brachiocephalic artery Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|26368-1|LNC|Brachiocephalic artery left Fluoroscopic angiogram Angioplasty W contrast IA|Brachiocephalic artery left Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|26369-9|LNC|Brachiocephalic artery right Fluoroscopic angiogram Angioplasty W contrast IA|Brachiocephalic artery right Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|24614-0|LNC|Carotid artery extracranial Fluoroscopic angiogram Angioplasty W contrast IA|Carotid artery extracranial Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|24615-7|LNC|Carotid artery intracranial Fluoroscopic angiogram Angioplasty W contrast IA|Carotid artery intracranial Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|35881-2|LNC|Extremity artery Fluoroscopic angiogram Angioplasty W contrast IA|Extremity artery Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|24698-3|LNC|Femoral artery Fluoroscopic angiogram Angioplasty W contrast IA|Femoral artery Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|36763-1|LNC|Femoral artery Popliteal artery Fluoroscopic angiogram Angioplasty W contrast IA|Femoral artery Popliteal artery Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|24766-8|LNC|Iliac artery Fluoroscopic angiogram Angioplasty W contrast IA|Iliac artery Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|26370-7|LNC|Iliac artery bilateral Fluoroscopic angiogram Angioplasty W contrast IA|Iliac artery bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|26371-5|LNC|Iliac artery left Fluoroscopic angiogram Angioplasty W contrast IA|Iliac artery left Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|26372-3|LNC|Iliac artery right Fluoroscopic angiogram Angioplasty W contrast IA|Iliac artery right Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|24832-8|LNC|Mesenteric artery Fluoroscopic angiogram Angioplasty W contrast IA|Mesenteric artery Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|30648-0|LNC|Peripheral artery Fluoroscopic angiogram Angioplasty W contrast IA|Peripheral artery Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|25081-1|LNC|Renal vessel Fluoroscopic angiogram Angioplasty W contrast IA|Renal vessel Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|25012-6|LNC|Tibial artery Fluoroscopic angiogram Angioplasty W contrast IA|Tibial artery Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|26373-1|LNC|Tibial artery bilateral Fluoroscopic angiogram Angioplasty W contrast IA|Tibial artery bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|26374-9|LNC|Tibial artery left Fluoroscopic angiogram Angioplasty W contrast IA|Tibial artery left Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|26375-6|LNC|Tibial artery right Fluoroscopic angiogram Angioplasty W contrast IA|Tibial artery right Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|43793-9|LNC|Tibioperoneal arteries Fluoroscopic angiogram Angioplasty W contrast IA|Tibioperoneal arteries Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|43794-7|LNC|Tibioperoneal arteries bilateral Fluoroscopic angiogram Angioplasty W contrast IA|Tibioperoneal arteries bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|43795-4|LNC|Tibioperoneal arteries left Fluoroscopic angiogram Angioplasty W contrast IA|Tibioperoneal arteries left Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|43792-1|LNC|Tibioperoneal arteries right Fluoroscopic angiogram Angioplasty W contrast IA|Tibioperoneal arteries right Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|25064-7|LNC|Vessel Fluoroscopic angiogram Angioplasty W contrast IA|Vessel Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|30836-1|LNC|Visceral artery Fluoroscopic angiogram Angioplasty W contrast IA|Visceral artery Fluoroscopic angiogram Angioplasty W contrast IA
C0801762|T102|relax|37426-4|LNC|Lower extremity vein Fluoroscopic angiogram Angioplasty W contrast IV|Lower extremity vein Fluoroscopic angiogram Angioplasty W contrast IV
C0801762|T102|relax|30640-7|LNC|Vein Fluoroscopic angiogram Angioplasty W contrast IV|Vein Fluoroscopic angiogram Angioplasty W contrast IV
C0801762|T102|relax|35882-0|LNC|Inferior vena cava Fluoroscopic angiogram Angioplasty W contrast IV|Inferior vena cava Fluoroscopic angiogram Angioplasty W contrast IV
C0801762|T102|relax|36764-9|LNC|Femoral vessel Popliteal artery Fluoroscopic angiogram Atherectomy W contrast|Femoral vessel Popliteal artery Fluoroscopic angiogram Atherectomy W contrast
C0801762|T102|relax|69135-2|LNC|Iliac artery Fluoroscopic angiogram Atherectomy W contrast|Iliac artery Fluoroscopic angiogram Atherectomy W contrast
C0801762|T102|relax|69253-3|LNC|Renal vessels Fluoroscopic angiogram Atherectomy W contrast|Renal vessels Fluoroscopic angiogram Atherectomy W contrast
C0801762|T102|relax|36765-6|LNC|Vessel Fluoroscopic angiogram Atherectomy W contrast|Vessel Fluoroscopic angiogram Atherectomy W contrast
C0801762|T102|relax|35883-8|LNC|Aorta Fluoroscopic angiogram Atherectomy W contrast IA|Aorta Fluoroscopic angiogram Atherectomy W contrast IA
C0801762|T102|relax|36766-4|LNC|Coronary arteries Fluoroscopic angiogram Atherectomy W contrast IA|Coronary arteries Fluoroscopic angiogram Atherectomy W contrast IA
C0801762|T102|relax|24568-8|LNC|AV fistula Fluoroscopic angiogram Atherectomy W contrast IV|AV fistula Fluoroscopic angiogram Atherectomy W contrast IV
C0801762|T102|relax|36761-5|LNC|Biliary ducts Fluoroscopy Balloon dilatation W contrast|Biliary ducts Fluoroscopy Balloon dilatation W contrast
C0801762|T102|relax|38268-9|LNC|Skeletal system DXA Bone density|Skeletal system DXA Bone density
C0801762|T102|relax|43562-8|LNC|Skeletal system axial Scan Bone density|Skeletal system axial Scan Bone density
C0801762|T102|relax|43563-6|LNC|Skeletal system peripheral Scan Bone density|Skeletal system peripheral Scan Bone density
C0801762|T102|relax|24631-4|LNC|Unspecified body region Fluoroscopy Central vein catheter placement check|Unspecified body region Fluoroscopy Central vein catheter placement check
C0801762|T102|relax|25062-1|LNC|Unspecified body region X-ray Comparison view|Unspecified body region X-ray Comparison view
C0801762|T102|relax|72555-6|LNC|Interventional radiology Consult note|Interventional radiology Consult note
C0801762|T102|relax|25038-1|LNC|Unspecified body region Courtesy consultation|Unspecified body region Courtesy consultation
C0801762|T102|relax|24684-3|LNC|Extracranial vessels Fluoroscopic angiogram Embolectomy W contrast IA|Extracranial vessels Fluoroscopic angiogram Embolectomy W contrast IA
C0801762|T102|relax|24887-2|LNC|Pulmonary artery Fluoroscopic angiogram Embolectomy W contrast IA|Pulmonary artery Fluoroscopic angiogram Embolectomy W contrast IA
C0801762|T102|relax|24553-0|LNC|Vessel intracranial Fluoroscopic angiogram Embolectomy W contrast IV|Vessel intracranial Fluoroscopic angiogram Embolectomy W contrast IV
C0801762|T102|relax|24554-8|LNC|Artery Fluoroscopic angiogram Embolization W contrast IA|Artery Fluoroscopic angiogram Embolization W contrast IA
C0801762|T102|relax|30600-1|LNC|Small bowel CT Views Enteroclysis W contrast PO via duodenal intubation|Small bowel CT Views Enteroclysis W contrast PO via duodenal intubation
C0801762|T102|relax|24923-5|LNC|Small bowel Fluoroscopy Views Enteroclysis W contrast PO via duodenal intubation|Small bowel Fluoroscopy Views Enteroclysis W contrast PO via duodenal intubation
C0801762|T102|relax|46365-3|LNC|CT Guided ablation tissue Celiac plexus|CT Guided ablation tissue Celiac plexus
C0801762|T102|relax|44228-5|LNC|CT Guided ablation tissue Kidney|CT Guided ablation tissue Kidney
C0801762|T102|relax|44156-8|LNC|US Guided ablation tissue Kidney|US Guided ablation tissue Kidney
C0801762|T102|relax|44101-4|LNC|CT Guided ablation tissue Liver|CT Guided ablation tissue Liver
C0801762|T102|relax|44155-0|LNC|US Guided ablation tissue Liver|US Guided ablation tissue Liver
C0801762|T102|relax|58747-7|LNC|CT Guided ablation tissue Unspecified body region|CT Guided ablation tissue Unspecified body region
C0801762|T102|relax|58743-6|LNC|US Guided ablation tissue Unspecified body region|US Guided ablation tissue Unspecified body region
C0801762|T102|relax|35884-6|LNC|CT Guided abscess drainage Abdomen|CT Guided abscess drainage Abdomen
C0801762|T102|relax|42280-8|LNC|CT Guided abscess drainage Appendix|CT Guided abscess drainage Appendix
C0801762|T102|relax|42705-4|LNC|US Guided abscess drainage Appendix|US Guided abscess drainage Appendix
C0801762|T102|relax|42281-6|LNC|CT Guided abscess drainage Chest|CT Guided abscess drainage Chest
C0801762|T102|relax|42285-7|LNC|CT Guided abscess drainage Kidney|CT Guided abscess drainage Kidney
C0801762|T102|relax|44167-5|LNC|US Guided abscess drainage Kidney|US Guided abscess drainage Kidney
C0801762|T102|relax|42282-4|LNC|CT Guided abscess drainage Liver|CT Guided abscess drainage Liver
C0801762|T102|relax|42133-9|LNC|US Guided abscess drainage Liver|US Guided abscess drainage Liver
C0801762|T102|relax|39361-1|LNC|Fluoroscopy Guided abscess drainage Liver|Fluoroscopy Guided abscess drainage Liver
C0801762|T102|relax|69120-4|LNC|Fluoroscopy Guided abscess drainage Neck|Fluoroscopy Guided abscess drainage Neck
C0801762|T102|relax|69122-0|LNC|Fluoroscopy Guided abscess drainage Pancreas|Fluoroscopy Guided abscess drainage Pancreas
C0801762|T102|relax|42286-5|LNC|CT Guided abscess drainage Pelvis|CT Guided abscess drainage Pelvis
C0801762|T102|relax|44168-3|LNC|US Guided abscess drainage Pelvis|US Guided abscess drainage Pelvis
C0801762|T102|relax|44169-1|LNC|US Guided abscess drainage Peritoneal space|US Guided abscess drainage Peritoneal space
C0801762|T102|relax|42284-0|LNC|CT Guided abscess drainage Pleural space|CT Guided abscess drainage Pleural space
C0801762|T102|relax|69123-8|LNC|Fluoroscopy Guided abscess drainage Pleural space|Fluoroscopy Guided abscess drainage Pleural space
C0801762|T102|relax|43502-4|LNC|CT Guided abscess drainage Subphrenic space|CT Guided abscess drainage Subphrenic space
C0801762|T102|relax|44166-7|LNC|US Guided abscess drainage Subphrenic space|US Guided abscess drainage Subphrenic space
C0801762|T102|relax|30578-9|LNC|CT Guided abscess drainage Unspecified body region|CT Guided abscess drainage Unspecified body region
C0801762|T102|relax|39451-0|LNC|US Guided abscess drainage Unspecified body region|US Guided abscess drainage Unspecified body region
C0801762|T102|relax|35885-3|LNC|Fluoroscopy Guided abscess drainage Unspecified body region|Fluoroscopy Guided abscess drainage Unspecified body region
C0801762|T102|relax|39620-0|LNC|Scan Guided abscess localization limited|Scan Guided abscess localization limited
C0801762|T102|relax|39623-4|LNC|Scan Guided abscess localization whole body|Scan Guided abscess localization whole body
C0801762|T102|relax|39622-6|LNC|SPECT Guided abscess localization whole body|SPECT Guided abscess localization whole body
C0801762|T102|relax|39621-8|LNC|SPECT Guided abscess localization|SPECT Guided abscess localization
C0801762|T102|relax|72533-3|LNC|US Guided ambulatory phlebectomy Extremity vein left|US Guided ambulatory phlebectomy Extremity vein left
C0801762|T102|relax|72532-5|LNC|US Guided ambulatory phlebectomy Extremity vein right|US Guided ambulatory phlebectomy Extremity vein right
C0801762|T102|relax|24623-1|LNC|CT Guided anesthetic block injection Celiac plexus|CT Guided anesthetic block injection Celiac plexus
C0801762|T102|relax|35886-1|LNC|CT Guided aspiration Breast|CT Guided aspiration Breast
C0801762|T102|relax|24598-5|LNC|Mammogram Guided aspiration Breast|Mammogram Guided aspiration Breast
C0801762|T102|relax|43756-6|LNC|US Guided aspiration Breast|US Guided aspiration Breast
C0801762|T102|relax|69278-0|LNC|US Guided aspiration Breast bilateral|US Guided aspiration Breast bilateral
C0801762|T102|relax|69292-1|LNC|US Guided aspiration Breast left|US Guided aspiration Breast left
C0801762|T102|relax|69296-2|LNC|US Guided aspiration Breast right|US Guided aspiration Breast right
C0801762|T102|relax|35888-7|LNC|Fluoroscopy Guided aspiration Hip|Fluoroscopy Guided aspiration Hip
C0801762|T102|relax|24771-8|LNC|Fluoroscopy Guided aspiration Joint space|Fluoroscopy Guided aspiration Joint space
C0801762|T102|relax|48434-5|LNC|US Guided aspiration Kidney|US Guided aspiration Kidney
C0801762|T102|relax|24811-2|LNC|CT Guided aspiration Liver|CT Guided aspiration Liver
C0801762|T102|relax|24822-9|LNC|CT Guided aspiration Lung|CT Guided aspiration Lung
C0801762|T102|relax|69287-1|LNC|US Guided aspiration Lymph node|US Guided aspiration Lymph node
C0801762|T102|relax|24837-7|LNC|CT Guided aspiration Neck|CT Guided aspiration Neck
C0801762|T102|relax|39452-8|LNC|US Guided aspiration Ovary|US Guided aspiration Ovary
C0801762|T102|relax|24856-7|LNC|CT Guided aspiration Pancreas|CT Guided aspiration Pancreas
C0801762|T102|relax|24863-3|LNC|CT Guided aspiration Pelvis|CT Guided aspiration Pelvis
C0801762|T102|relax|30703-3|LNC|US Guided aspiration Pericardial space|US Guided aspiration Pericardial space
C0801762|T102|relax|37491-8|LNC|CT Guided aspiration Pleural space|CT Guided aspiration Pleural space
C0801762|T102|relax|24662-9|LNC|US Guided aspiration Pleural space|US Guided aspiration Pleural space
C0801762|T102|relax|37887-7|LNC|Fluoroscopy Guided aspiration Pleural space|Fluoroscopy Guided aspiration Pleural space
C0801762|T102|relax|24973-0|LNC|Fluoroscopy Guided aspiration Spine Lumbar Space|Fluoroscopy Guided aspiration Spine Lumbar Space
C0801762|T102|relax|42134-7|LNC|US Guided aspiration Thyroid|US Guided aspiration Thyroid
C0801762|T102|relax|25043-1|LNC|CT Guided aspiration Unspecified body region|CT Guided aspiration Unspecified body region
C0801762|T102|relax|30878-3|LNC|US Guided aspiration Unspecified body region|US Guided aspiration Unspecified body region
C0801762|T102|relax|36926-4|LNC|CT Guided aspiration placement drainage tube Abdomen|CT Guided aspiration placement drainage tube Abdomen
C0801762|T102|relax|37210-2|LNC|CT Guided aspiration cyst Abdomen|CT Guided aspiration cyst Abdomen
C0801762|T102|relax|69306-9|LNC|Fluoroscopy Guided aspiration cyst Bone|Fluoroscopy Guided aspiration cyst Bone
C0801762|T102|relax|24594-4|LNC|Mammogram Guided aspiration cyst Breast|Mammogram Guided aspiration cyst Breast
C0801762|T102|relax|69192-3|LNC|MRI Guided aspiration cyst Breast|MRI Guided aspiration cyst Breast
C0801762|T102|relax|30653-0|LNC|US Guided aspiration cyst Breast|US Guided aspiration cyst Breast
C0801762|T102|relax|26343-4|LNC|Mammogram Guided aspiration cyst Breast bilateral|Mammogram Guided aspiration cyst Breast bilateral
C0801762|T102|relax|38012-1|LNC|US Guided aspiration cyst Breast bilateral|US Guided aspiration cyst Breast bilateral
C0801762|T102|relax|26344-2|LNC|Mammogram Guided aspiration cyst Breast left|Mammogram Guided aspiration cyst Breast left
C0801762|T102|relax|42450-7|LNC|US Guided aspiration cyst Breast left|US Guided aspiration cyst Breast left
C0801762|T102|relax|26345-9|LNC|Mammogram Guided aspiration cyst Breast right|Mammogram Guided aspiration cyst Breast right
C0801762|T102|relax|42458-0|LNC|US Guided aspiration cyst Breast right|US Guided aspiration cyst Breast right
C0801762|T102|relax|38126-9|LNC|US Guided aspiration cyst Kidney|US Guided aspiration cyst Kidney
C0801762|T102|relax|69121-2|LNC|Fluoroscopy Guided aspiration cyst Ovary|Fluoroscopy Guided aspiration cyst Ovary
C0801762|T102|relax|38133-5|LNC|US Guided aspiration cyst Pancreas|US Guided aspiration cyst Pancreas
C0801762|T102|relax|42447-3|LNC|US Guided aspiration cyst Thyroid|US Guided aspiration cyst Thyroid
C0801762|T102|relax|35887-9|LNC|CT Guided aspiration cyst Unspecified body region|CT Guided aspiration cyst Unspecified body region
C0801762|T102|relax|30698-5|LNC|US Guided aspiration cyst Unspecified body region|US Guided aspiration cyst Unspecified body region
C0801762|T102|relax|24671-0|LNC|Fluoroscopy Guided aspiration cyst Unspecified body region|Fluoroscopy Guided aspiration cyst Unspecified body region
C0801762|T102|relax|25042-3|LNC|CT Guided aspiration or biopsy Unspecified body region|CT Guided aspiration or biopsy Unspecified body region
C0801762|T102|relax|25041-5|LNC|CT Guided aspiration or biopsy Unspecified body region-- W contrast IV|CT Guided aspiration or biopsy Unspecified body region-- W contrast IV
C0801762|T102|relax|46281-2|LNC|CT Guided aspiration or injection cyst Unspecified body region|CT Guided aspiration or injection cyst Unspecified body region
C0801762|T102|relax|46282-0|LNC|US Guided aspiration or injection cyst Unspecified body region|US Guided aspiration or injection cyst Unspecified body region
C0801762|T102|relax|30602-7|LNC|CT Guided fine needle aspiration Abdomen|CT Guided fine needle aspiration Abdomen
C0801762|T102|relax|44107-1|LNC|CT Guided fine needle aspiration Abdomen retroperitoneum|CT Guided fine needle aspiration Abdomen retroperitoneum
C0801762|T102|relax|44108-9|LNC|CT Guided fine needle aspiration Adrenal gland|CT Guided fine needle aspiration Adrenal gland
C0801762|T102|relax|46387-7|LNC|Mammogram Guided fine needle aspiration Breast|Mammogram Guided fine needle aspiration Breast
C0801762|T102|relax|44160-0|LNC|US Guided fine needle aspiration Breast|US Guided fine needle aspiration Breast
C0801762|T102|relax|46284-6|LNC|Mammogram Guided fine needle aspiration Breast left|Mammogram Guided fine needle aspiration Breast left
C0801762|T102|relax|38026-1|LNC|US Guided fine needle aspiration Breast left|US Guided fine needle aspiration Breast left
C0801762|T102|relax|46283-8|LNC|Mammogram Guided fine needle aspiration Breast right|Mammogram Guided fine needle aspiration Breast right
C0801762|T102|relax|38033-7|LNC|US Guided fine needle aspiration Breast right|US Guided fine needle aspiration Breast right
C0801762|T102|relax|38135-0|LNC|US Guided fine needle aspiration Deep tissue|US Guided fine needle aspiration Deep tissue
C0801762|T102|relax|44221-0|LNC|Fluoroscopy Guided fine needle aspiration Deep tissue|Fluoroscopy Guided fine needle aspiration Deep tissue
C0801762|T102|relax|43757-4|LNC|CT Guided fine needle aspiration Kidney|CT Guided fine needle aspiration Kidney
C0801762|T102|relax|44159-2|LNC|US Guided fine needle aspiration Kidney|US Guided fine needle aspiration Kidney
C0801762|T102|relax|44217-8|LNC|Fluoroscopy Guided fine needle aspiration Kidney|Fluoroscopy Guided fine needle aspiration Kidney
C0801762|T102|relax|30608-4|LNC|CT Guided fine needle aspiration Kidney bilateral|CT Guided fine needle aspiration Kidney bilateral
C0801762|T102|relax|30603-5|LNC|CT Guided fine needle aspiration Liver|CT Guided fine needle aspiration Liver
C0801762|T102|relax|44158-4|LNC|US Guided fine needle aspiration Liver|US Guided fine needle aspiration Liver
C0801762|T102|relax|44220-2|LNC|Fluoroscopy Guided fine needle aspiration Liver|Fluoroscopy Guided fine needle aspiration Liver
C0801762|T102|relax|30595-3|LNC|CT Guided fine needle aspiration Lung|CT Guided fine needle aspiration Lung
C0801762|T102|relax|44103-0|LNC|CT Guided fine needle aspiration Lymph node|CT Guided fine needle aspiration Lymph node
C0801762|T102|relax|44219-4|LNC|Fluoroscopy Guided fine needle aspiration Lymph node|Fluoroscopy Guided fine needle aspiration Lymph node
C0801762|T102|relax|44104-8|LNC|CT Guided fine needle aspiration Mediastinum|CT Guided fine needle aspiration Mediastinum
C0801762|T102|relax|44105-5|LNC|CT Guided fine needle aspiration Muscle|CT Guided fine needle aspiration Muscle
C0801762|T102|relax|30605-0|LNC|CT Guided fine needle aspiration Pancreas|CT Guided fine needle aspiration Pancreas
C0801762|T102|relax|44157-6|LNC|US Guided fine needle aspiration Pancreas|US Guided fine needle aspiration Pancreas
C0801762|T102|relax|44218-6|LNC|Fluoroscopy Guided fine needle aspiration Pancreas|Fluoroscopy Guided fine needle aspiration Pancreas
C0801762|T102|relax|30606-8|LNC|CT Guided fine needle aspiration Pelvis|CT Guided fine needle aspiration Pelvis
C0801762|T102|relax|44106-3|LNC|CT Guided fine needle aspiration Prostate|CT Guided fine needle aspiration Prostate
C0801762|T102|relax|38017-0|LNC|US Guided fine needle aspiration Prostate|US Guided fine needle aspiration Prostate
C0801762|T102|relax|30610-0|LNC|CT Guided fine needle aspiration Spleen|CT Guided fine needle aspiration Spleen
C0801762|T102|relax|38136-8|LNC|US Guided fine needle aspiration Superficial tissue|US Guided fine needle aspiration Superficial tissue
C0801762|T102|relax|69124-6|LNC|Fluoroscopy Guided fine needle aspiration Superficial tissue|Fluoroscopy Guided fine needle aspiration Superficial tissue
C0801762|T102|relax|38019-6|LNC|US Guided fine needle aspiration Thyroid|US Guided fine needle aspiration Thyroid
C0801762|T102|relax|44216-0|LNC|Fluoroscopy Guided fine needle aspiration Thyroid|Fluoroscopy Guided fine needle aspiration Thyroid
C0801762|T102|relax|30580-5|LNC|CT Guided fine needle aspiration Unspecified body region|CT Guided fine needle aspiration Unspecified body region
C0801762|T102|relax|38018-8|LNC|US Guided fine needle aspiration Unspecified body region|US Guided fine needle aspiration Unspecified body region
C0801762|T102|relax|44215-2|LNC|Fluoroscopy Guided fine needle aspiration Unspecified body region|Fluoroscopy Guided fine needle aspiration Unspecified body region
C0801762|T102|relax|24755-1|LNC|Fluoroscopic angiogram Guided atherectomy Vein-- W contrast IV|Fluoroscopic angiogram Guided atherectomy Vein-- W contrast IV
C0801762|T102|relax|26298-0|LNC|Fluoroscopic angiogram Guided atherectomy Vein bilateral-- W contrast IV|Fluoroscopic angiogram Guided atherectomy Vein bilateral-- W contrast IV
C0801762|T102|relax|26299-8|LNC|Fluoroscopic angiogram Guided atherectomy Vein left-- W contrast IV|Fluoroscopic angiogram Guided atherectomy Vein left-- W contrast IV
C0801762|T102|relax|26300-4|LNC|Fluoroscopic angiogram Guided atherectomy Vein right-- W contrast IV|Fluoroscopic angiogram Guided atherectomy Vein right-- W contrast IV
C0801762|T102|relax|30601-9|LNC|CT Guided biopsy Abdomen|CT Guided biopsy Abdomen
C0801762|T102|relax|37913-1|LNC|US Guided biopsy Abdomen|US Guided biopsy Abdomen
C0801762|T102|relax|35890-3|LNC|Fluoroscopy Guided biopsy Abdomen|Fluoroscopy Guided biopsy Abdomen
C0801762|T102|relax|44117-0|LNC|CT Guided biopsy Abdomen retroperitoneum|CT Guided biopsy Abdomen retroperitoneum
C0801762|T102|relax|44162-6|LNC|US Guided biopsy Abdomen retroperitoneum|US Guided biopsy Abdomen retroperitoneum
C0801762|T102|relax|36767-2|LNC|CT Guided biopsy Adrenal gland|CT Guided biopsy Adrenal gland
C0801762|T102|relax|35891-1|LNC|CT Guided biopsy Bone|CT Guided biopsy Bone
C0801762|T102|relax|69076-8|LNC|Fluoroscopy Guided biopsy Bone|Fluoroscopy Guided biopsy Bone
C0801762|T102|relax|37211-0|LNC|CT Guided biopsy Bone marrow|CT Guided biopsy Bone marrow
C0801762|T102|relax|35893-7|LNC|CT Guided biopsy Breast|CT Guided biopsy Breast
C0801762|T102|relax|24602-5|LNC|Mammogram Guided biopsy Breast|Mammogram Guided biopsy Breast
C0801762|T102|relax|37914-9|LNC|US Guided biopsy Breast|US Guided biopsy Breast
C0801762|T102|relax|26337-6|LNC|Mammogram Guided biopsy Breast bilateral|Mammogram Guided biopsy Breast bilateral
C0801762|T102|relax|69169-1|LNC|MRI Guided biopsy Breast bilateral|MRI Guided biopsy Breast bilateral
C0801762|T102|relax|37912-3|LNC|US Guided biopsy Breast bilateral|US Guided biopsy Breast bilateral
C0801762|T102|relax|26338-4|LNC|Mammogram Guided biopsy Breast left|Mammogram Guided biopsy Breast left
C0801762|T102|relax|69203-8|LNC|MRI Guided biopsy Breast left|MRI Guided biopsy Breast left
C0801762|T102|relax|42449-9|LNC|US Guided biopsy Breast left|US Guided biopsy Breast left
C0801762|T102|relax|26339-2|LNC|Mammogram Guided biopsy Breast right|Mammogram Guided biopsy Breast right
C0801762|T102|relax|69213-7|LNC|MRI Guided biopsy Breast right|MRI Guided biopsy Breast right
C0801762|T102|relax|42457-2|LNC|US Guided biopsy Breast right|US Guided biopsy Breast right
C0801762|T102|relax|35895-2|LNC|CT Guided biopsy Chest|CT Guided biopsy Chest
C0801762|T102|relax|37915-6|LNC|US Guided biopsy Chest|US Guided biopsy Chest
C0801762|T102|relax|35894-5|LNC|Fluoroscopy Guided biopsy Chest|Fluoroscopy Guided biopsy Chest
C0801762|T102|relax|37492-6|LNC|CT Guided biopsy Chest pleura|CT Guided biopsy Chest pleura
C0801762|T102|relax|42333-5|LNC|US Guided biopsy Chest pleura|US Guided biopsy Chest pleura
C0801762|T102|relax|43567-7|LNC|CT Guided biopsy Deep bone|CT Guided biopsy Deep bone
C0801762|T102|relax|43565-1|LNC|US Guided biopsy Deep bone|US Guided biopsy Deep bone
C0801762|T102|relax|44109-7|LNC|CT Guided biopsy Deep muscle|CT Guided biopsy Deep muscle
C0801762|T102|relax|42463-0|LNC|US Guided biopsy Endomyocardium|US Guided biopsy Endomyocardium
C0801762|T102|relax|37212-8|LNC|CT Guided biopsy Epididymis|CT Guided biopsy Epididymis
C0801762|T102|relax|69387-9|LNC|US Guided biopsy Epididymis|US Guided biopsy Epididymis
C0801762|T102|relax|36927-2|LNC|CT Guided biopsy Facial bones Maxilla|CT Guided biopsy Facial bones Maxilla
C0801762|T102|relax|35892-9|LNC|CT Guided biopsy Head|CT Guided biopsy Head
C0801762|T102|relax|42136-2|LNC|CT Guided biopsy Heart|CT Guided biopsy Heart
C0801762|T102|relax|42279-0|LNC|CT Guided biopsy Kidney|CT Guided biopsy Kidney
C0801762|T102|relax|24772-6|LNC|US Guided biopsy Kidney|US Guided biopsy Kidney
C0801762|T102|relax|35899-4|LNC|Fluoroscopy Guided biopsy Kidney|Fluoroscopy Guided biopsy Kidney
C0801762|T102|relax|38766-2|LNC|US Guided biopsy Kidney transplant|US Guided biopsy Kidney transplant
C0801762|T102|relax|30607-6|LNC|CT Guided biopsy Kidney bilateral|CT Guided biopsy Kidney bilateral
C0801762|T102|relax|26340-0|LNC|US Guided biopsy Kidney bilateral|US Guided biopsy Kidney bilateral
C0801762|T102|relax|26341-8|LNC|US Guided biopsy Kidney left|US Guided biopsy Kidney left
C0801762|T102|relax|26342-6|LNC|US Guided biopsy Kidney right|US Guided biopsy Kidney right
C0801762|T102|relax|24812-0|LNC|CT Guided biopsy Liver|CT Guided biopsy Liver
C0801762|T102|relax|24816-1|LNC|US Guided biopsy Liver|US Guided biopsy Liver
C0801762|T102|relax|35900-0|LNC|Fluoroscopy Guided biopsy Liver|Fluoroscopy Guided biopsy Liver
C0801762|T102|relax|38765-4|LNC|US Guided biopsy Liver transplant|US Guided biopsy Liver transplant
C0801762|T102|relax|35896-0|LNC|CT Guided biopsy Lower extremity|CT Guided biopsy Lower extremity
C0801762|T102|relax|24823-7|LNC|CT Guided biopsy Lung|CT Guided biopsy Lung
C0801762|T102|relax|44161-8|LNC|US Guided biopsy Lung|US Guided biopsy Lung
C0801762|T102|relax|30634-0|LNC|Fluoroscopy Guided biopsy Lung|Fluoroscopy Guided biopsy Lung
C0801762|T102|relax|35901-8|LNC|CT Guided biopsy Lymph node|CT Guided biopsy Lymph node
C0801762|T102|relax|39522-8|LNC|US Guided biopsy Lymph node|US Guided biopsy Lymph node
C0801762|T102|relax|37213-6|LNC|CT Guided biopsy Mediastinum|CT Guided biopsy Mediastinum
C0801762|T102|relax|42137-0|LNC|US Guided biopsy Mediastinum|US Guided biopsy Mediastinum
C0801762|T102|relax|36768-0|LNC|CT Guided biopsy Muscle|CT Guided biopsy Muscle
C0801762|T102|relax|37917-2|LNC|US Guided biopsy Muscle|US Guided biopsy Muscle
C0801762|T102|relax|24838-5|LNC|CT Guided biopsy Neck|CT Guided biopsy Neck
C0801762|T102|relax|37918-0|LNC|US Guided biopsy Neck|US Guided biopsy Neck
C0801762|T102|relax|30604-3|LNC|CT Guided biopsy Pancreas|CT Guided biopsy Pancreas
C0801762|T102|relax|37919-8|LNC|US Guided biopsy Pancreas|US Guided biopsy Pancreas
C0801762|T102|relax|35902-6|LNC|Fluoroscopy Guided biopsy Pancreas|Fluoroscopy Guided biopsy Pancreas
C0801762|T102|relax|24864-1|LNC|CT Guided biopsy Pelvis|CT Guided biopsy Pelvis
C0801762|T102|relax|69074-3|LNC|Fluoroscopy Guided biopsy Pelvis|Fluoroscopy Guided biopsy Pelvis
C0801762|T102|relax|35903-4|LNC|CT Guided biopsy Prostate|CT Guided biopsy Prostate
C0801762|T102|relax|24883-1|LNC|US Guided biopsy Prostate|US Guided biopsy Prostate
C0801762|T102|relax|41802-0|LNC|Fluoroscopy Guided biopsy Prostate|Fluoroscopy Guided biopsy Prostate
C0801762|T102|relax|35898-6|LNC|CT Guided biopsy Salivary gland|CT Guided biopsy Salivary gland
C0801762|T102|relax|37920-6|LNC|US Guided biopsy Salivary gland|US Guided biopsy Salivary gland
C0801762|T102|relax|69075-0|LNC|Fluoroscopy Guided biopsy Salivary gland|Fluoroscopy Guided biopsy Salivary gland
C0801762|T102|relax|38132-7|LNC|US Guided biopsy Scrotum Testicle|US Guided biopsy Scrotum Testicle
C0801762|T102|relax|69396-0|LNC|US Guided biopsy Spinal cord|US Guided biopsy Spinal cord
C0801762|T102|relax|35904-2|LNC|CT Guided biopsy Spine Cervical|CT Guided biopsy Spine Cervical
C0801762|T102|relax|35905-9|LNC|CT Guided biopsy Spine Lumbar|CT Guided biopsy Spine Lumbar
C0801762|T102|relax|35906-7|LNC|CT Guided biopsy Spine Thoracic|CT Guided biopsy Spine Thoracic
C0801762|T102|relax|30609-2|LNC|CT Guided biopsy Spleen|CT Guided biopsy Spleen
C0801762|T102|relax|35907-5|LNC|Fluoroscopy Guided biopsy Spleen|Fluoroscopy Guided biopsy Spleen
C0801762|T102|relax|42265-9|LNC|CT Guided biopsy Superficial bone|CT Guided biopsy Superficial bone
C0801762|T102|relax|42135-4|LNC|US Guided biopsy Superficial bone|US Guided biopsy Superficial bone
C0801762|T102|relax|38154-1|LNC|Fluoroscopy Guided biopsy Superficial bone|Fluoroscopy Guided biopsy Superficial bone
C0801762|T102|relax|43797-0|LNC|US Guided biopsy Superficial lymph node|US Guided biopsy Superficial lymph node
C0801762|T102|relax|43564-4|LNC|US Guided biopsy Superficial muscle|US Guided biopsy Superficial muscle
C0801762|T102|relax|37214-4|LNC|CT Guided biopsy Superficial tissue|CT Guided biopsy Superficial tissue
C0801762|T102|relax|35908-3|LNC|CT Guided biopsy Thyroid|CT Guided biopsy Thyroid
C0801762|T102|relax|25009-2|LNC|US Guided biopsy Thyroid|US Guided biopsy Thyroid
C0801762|T102|relax|35897-8|LNC|CT Guided biopsy Upper extremity|CT Guided biopsy Upper extremity
C0801762|T102|relax|25044-9|LNC|CT Guided biopsy Unspecified body region|CT Guided biopsy Unspecified body region
C0801762|T102|relax|25059-7|LNC|US Guided biopsy Unspecified body region|US Guided biopsy Unspecified body region
C0801762|T102|relax|25069-6|LNC|Fluoroscopy Guided biopsy Unspecified body region|Fluoroscopy Guided biopsy Unspecified body region
C0801762|T102|relax|24670-2|LNC|US Guided biopsy cyst Unspecified body region|US Guided biopsy cyst Unspecified body region
C0801762|T102|relax|30651-4|LNC|US Guided core needle biopsy Breast|US Guided core needle biopsy Breast
C0801762|T102|relax|24813-8|LNC|CT Guided core needle biopsy Liver|CT Guided core needle biopsy Liver
C0801762|T102|relax|69279-8|LNC|US Guided core needle biopsy Lymph node|US Guided core needle biopsy Lymph node
C0801762|T102|relax|46285-3|LNC|US Guided core needle biopsy Thyroid|US Guided core needle biopsy Thyroid
C0801762|T102|relax|38024-6|LNC|US Guided core needle biopsy Unspecified body region|US Guided core needle biopsy Unspecified body region
C0801762|T102|relax|69073-5|LNC|Fluoroscopy Guided core needle biopsy Unspecified body region|Fluoroscopy Guided core needle biopsy Unspecified body region
C0801762|T102|relax|42448-1|LNC|US Guided excisional biopsy Breast|US Guided excisional biopsy Breast
C0801762|T102|relax|30652-2|LNC|US Guided fine needle biopsy Breast|US Guided fine needle biopsy Breast
C0801762|T102|relax|42288-1|LNC|CT Guided needle biopsy Abdomen|CT Guided needle biopsy Abdomen
C0801762|T102|relax|69224-4|LNC|Fluoroscopy Guided needle biopsy Abdomen|Fluoroscopy Guided needle biopsy Abdomen
C0801762|T102|relax|46367-9|LNC|CT Guided needle biopsy Adrenal gland|CT Guided needle biopsy Adrenal gland
C0801762|T102|relax|46368-7|LNC|CT Guided needle biopsy Breast|CT Guided needle biopsy Breast
C0801762|T102|relax|46286-1|LNC|Mammogram Guided needle biopsy Breast|Mammogram Guided needle biopsy Breast
C0801762|T102|relax|38028-7|LNC|US Guided needle biopsy Breast|US Guided needle biopsy Breast
C0801762|T102|relax|41803-8|LNC|Fluoroscopy Guided needle biopsy Breast|Fluoroscopy Guided needle biopsy Breast
C0801762|T102|relax|43462-1|LNC|US Guided needle biopsy Breast left|US Guided needle biopsy Breast left
C0801762|T102|relax|43447-2|LNC|Mammogram Guided needle biopsy Breast right|Mammogram Guided needle biopsy Breast right
C0801762|T102|relax|69290-5|LNC|US Guided needle biopsy Breast right|US Guided needle biopsy Breast right
C0801762|T102|relax|38029-5|LNC|US Guided needle biopsy Chest|US Guided needle biopsy Chest
C0801762|T102|relax|69225-1|LNC|Fluoroscopy Guided needle biopsy Chest|Fluoroscopy Guided needle biopsy Chest
C0801762|T102|relax|69099-0|LNC|CT Guided needle biopsy Chest pleura|CT Guided needle biopsy Chest pleura
C0801762|T102|relax|44171-7|LNC|US Guided needle biopsy Chest pleura|US Guided needle biopsy Chest pleura
C0801762|T102|relax|69127-9|LNC|Fluoroscopy Guided needle biopsy Chest pleura|Fluoroscopy Guided needle biopsy Chest pleura
C0801762|T102|relax|43568-5|LNC|CT Guided needle biopsy Deep bone|CT Guided needle biopsy Deep bone
C0801762|T102|relax|42289-9|LNC|CT Guided needle biopsy Kidney|CT Guided needle biopsy Kidney
C0801762|T102|relax|38027-9|LNC|US Guided needle biopsy Kidney bilateral|US Guided needle biopsy Kidney bilateral
C0801762|T102|relax|69097-4|LNC|CT Guided needle biopsy Liver|CT Guided needle biopsy Liver
C0801762|T102|relax|69197-2|LNC|MRI Guided needle biopsy Liver|MRI Guided needle biopsy Liver
C0801762|T102|relax|44170-9|LNC|US Guided needle biopsy Liver|US Guided needle biopsy Liver
C0801762|T102|relax|69125-3|LNC|Fluoroscopy Guided needle biopsy Liver|Fluoroscopy Guided needle biopsy Liver
C0801762|T102|relax|42267-5|LNC|CT Guided needle biopsy Lymph node|CT Guided needle biopsy Lymph node
C0801762|T102|relax|37916-4|LNC|US Guided needle biopsy Lymph node|US Guided needle biopsy Lymph node
C0801762|T102|relax|69098-2|LNC|CT Guided needle biopsy Muscle|CT Guided needle biopsy Muscle
C0801762|T102|relax|69198-0|LNC|MRI Guided needle biopsy Muscle|MRI Guided needle biopsy Muscle
C0801762|T102|relax|69288-9|LNC|US Guided needle biopsy Muscle|US Guided needle biopsy Muscle
C0801762|T102|relax|69226-9|LNC|Fluoroscopy Guided needle biopsy Muscle|Fluoroscopy Guided needle biopsy Muscle
C0801762|T102|relax|46369-5|LNC|US Guided needle biopsy Ovary|US Guided needle biopsy Ovary
C0801762|T102|relax|42290-7|LNC|CT Guided needle biopsy Pancreas|CT Guided needle biopsy Pancreas
C0801762|T102|relax|69199-8|LNC|MRI Guided needle biopsy Pancreas|MRI Guided needle biopsy Pancreas
C0801762|T102|relax|69289-7|LNC|US Guided needle biopsy Pancreas|US Guided needle biopsy Pancreas
C0801762|T102|relax|69126-1|LNC|Fluoroscopy Guided needle biopsy Pancreas|Fluoroscopy Guided needle biopsy Pancreas
C0801762|T102|relax|46370-3|LNC|US Guided needle biopsy Pelvis|US Guided needle biopsy Pelvis
C0801762|T102|relax|69200-4|LNC|MRI Guided needle biopsy Pleura|MRI Guided needle biopsy Pleura
C0801762|T102|relax|69227-7|LNC|Fluoroscopy Guided needle biopsy Pleura|Fluoroscopy Guided needle biopsy Pleura
C0801762|T102|relax|46288-7|LNC|US Guided needle biopsy Prostate|US Guided needle biopsy Prostate
C0801762|T102|relax|69228-5|LNC|Fluoroscopy Guided needle biopsy Prostate|Fluoroscopy Guided needle biopsy Prostate
C0801762|T102|relax|69100-6|LNC|CT Guided needle biopsy Salivary gland|CT Guided needle biopsy Salivary gland
C0801762|T102|relax|69201-2|LNC|MRI Guided needle biopsy Salivary gland|MRI Guided needle biopsy Salivary gland
C0801762|T102|relax|69291-3|LNC|US Guided needle biopsy Salivary gland|US Guided needle biopsy Salivary gland
C0801762|T102|relax|69128-7|LNC|Fluoroscopy Guided needle biopsy Salivary gland|Fluoroscopy Guided needle biopsy Salivary gland
C0801762|T102|relax|43571-9|LNC|CT Guided needle biopsy Soft bone|CT Guided needle biopsy Soft bone
C0801762|T102|relax|69401-8|LNC|US Guided needle biopsy Spinal cord|US Guided needle biopsy Spinal cord
C0801762|T102|relax|38030-3|LNC|US Guided needle biopsy Spleen|US Guided needle biopsy Spleen
C0801762|T102|relax|42266-7|LNC|CT Guided needle biopsy Superficial bone|CT Guided needle biopsy Superficial bone
C0801762|T102|relax|69101-4|LNC|CT Guided needle biopsy Thyroid|CT Guided needle biopsy Thyroid
C0801762|T102|relax|69202-0|LNC|MRI Guided needle biopsy Thyroid|MRI Guided needle biopsy Thyroid
C0801762|T102|relax|38031-1|LNC|US Guided needle biopsy Thyroid|US Guided needle biopsy Thyroid
C0801762|T102|relax|69129-5|LNC|Fluoroscopy Guided needle biopsy Thyroid|Fluoroscopy Guided needle biopsy Thyroid
C0801762|T102|relax|46287-9|LNC|CT Guided needle biopsy Unspecified body region|CT Guided needle biopsy Unspecified body region
C0801762|T102|relax|30700-9|LNC|US Guided needle biopsy Unspecified body region|US Guided needle biopsy Unspecified body region
C0801762|T102|relax|44225-1|LNC|Fluoroscopy Guided needle biopsy Liver-- W contrast IV|Fluoroscopy Guided needle biopsy Liver-- W contrast IV
C0801762|T102|relax|24718-9|LNC|Fluoroscopy Guided transjugular biopsy Liver-- W contrast IV|Fluoroscopy Guided transjugular biopsy Liver-- W contrast IV
C0801762|T102|relax|35910-9|LNC|CT Guided biopsy Chest-- W WO contrast IV|CT Guided biopsy Chest-- W WO contrast IV
C0801762|T102|relax|46289-5|LNC|CT Guided biopsy Unspecified body region-- W WO contrast IV|CT Guided biopsy Unspecified body region-- W WO contrast IV
C0801762|T102|relax|35909-1|LNC|CT Guided biopsy Chest-- W contrast IV|CT Guided biopsy Chest-- W contrast IV
C0801762|T102|relax|69093-3|LNC|CT Guided biopsy Pelvis-- W contrast IV|CT Guided biopsy Pelvis-- W contrast IV
C0801762|T102|relax|42260-0|LNC|CT Guided biopsy Unspecified body region-- W contrast IV|CT Guided biopsy Unspecified body region-- W contrast IV
C0801762|T102|relax|46366-1|LNC|SPECT Guided biopsy Bone|SPECT Guided biopsy Bone
C0801762|T102|relax|46384-4|LNC|SPECT Guided biopsy Superficial bone|SPECT Guided biopsy Superficial bone
C0801762|T102|relax|69083-4|LNC|CT Guided biopsy Abdomen-- WO contrast|CT Guided biopsy Abdomen-- WO contrast
C0801762|T102|relax|35911-7|LNC|CT Guided biopsy Chest-- WO contrast|CT Guided biopsy Chest-- WO contrast
C0801762|T102|relax|69092-5|LNC|CT Guided biopsy Liver-- WO contrast|CT Guided biopsy Liver-- WO contrast
C0801762|T102|relax|69094-1|LNC|CT Guided biopsy Pelvis-- WO contrast|CT Guided biopsy Pelvis-- WO contrast
C0801762|T102|relax|46290-3|LNC|CT Guided biopsy Unspecified body region-- WO contrast|CT Guided biopsy Unspecified body region-- WO contrast
C0801762|T102|relax|35889-5|LNC|Fluoroscopy Guided bronchoscopy Chest|Fluoroscopy Guided bronchoscopy Chest
C0801762|T102|relax|64998-8|LNC|Fluoroscopy Guided catheterization Fallopian tube left-- transcervical|Fluoroscopy Guided catheterization Fallopian tube left-- transcervical
C0801762|T102|relax|64999-6|LNC|Fluoroscopy Guided catheterization Fallopian tube -right-- transcervical|Fluoroscopy Guided catheterization Fallopian tube -right-- transcervical
C0801762|T102|relax|30818-9|LNC|Fluoroscopy Guided catheterization Fallopian tubes-- transcervical|Fluoroscopy Guided catheterization Fallopian tubes-- transcervical
C0801762|T102|relax|30892-4|LNC|Fluoroscopy Guided catheterization Biliary ducts Pancreatic duct-- W contrast retrograde|Fluoroscopy Guided catheterization Biliary ducts Pancreatic duct-- W contrast retrograde
C0801762|T102|relax|24624-9|LNC|Fluoroscopic angiogram Guided change central catheter in Central vein-- W contrast IV|Fluoroscopic angiogram Guided change central catheter in Central vein-- W contrast IV
C0801762|T102|relax|26331-9|LNC|Fluoroscopic angiogram Guided change central catheter in Central vein bilateral-- W contrast IV|Fluoroscopic angiogram Guided change central catheter in Central vein bilateral-- W contrast IV
C0801762|T102|relax|26332-7|LNC|Fluoroscopic angiogram Guided change central catheter in Central vein left-- W contrast IV|Fluoroscopic angiogram Guided change central catheter in Central vein left-- W contrast IV
C0801762|T102|relax|26333-5|LNC|Fluoroscopic angiogram Guided change central catheter in Central vein right-- W contrast IV|Fluoroscopic angiogram Guided change central catheter in Central vein right-- W contrast IV
C0801762|T102|relax|43558-6|LNC|Fluoroscopy Guided change dialysis catheter in Unspecified body region-- W contrast IV|Fluoroscopy Guided change dialysis catheter in Unspecified body region-- W contrast IV
C0801762|T102|relax|36769-8|LNC|CT Guided change nephrostomy tube in Kidney|CT Guided change nephrostomy tube in Kidney
C0801762|T102|relax|24781-7|LNC|Fluoroscopy Guided change percutaneous nephrostomy tube in Kidney bilateral-- W contrast|Fluoroscopy Guided change percutaneous nephrostomy tube in Kidney bilateral-- W contrast
C0801762|T102|relax|46371-1|LNC|X-ray Guided change percutaneous tube in Unspecified body region-- W contrast|X-ray Guided change percutaneous tube in Unspecified body region-- W contrast
C0801762|T102|relax|30646-4|LNC|Fluoroscopy Guided change tube in Sinus tract-- W contrast|Fluoroscopy Guided change tube in Sinus tract-- W contrast
C0801762|T102|relax|69400-0|LNC|US Guided chorionic villus sampling|US Guided chorionic villus sampling
C0801762|T102|relax|69391-1|LNC|US Guided cordocentesis|US Guided cordocentesis
C0801762|T102|relax|70915-4|LNC|US Guided CSF aspiration Spine Cervical|US Guided CSF aspiration Spine Cervical
C0801762|T102|relax|70916-2|LNC|US Guided CSF aspiration Spine Lumbar|US Guided CSF aspiration Spine Lumbar
C0801762|T102|relax|70917-0|LNC|US Guided CSF aspiration Spine Thoracic|US Guided CSF aspiration Spine Thoracic
C0801762|T102|relax|24680-1|LNC|Fluoroscopy Guided dilation Esophagus|Fluoroscopy Guided dilation Esophagus
C0801762|T102|relax|35913-3|LNC|CT Guided drainage Abdomen|CT Guided drainage Abdomen
C0801762|T102|relax|42287-3|LNC|CT Guided drainage Abdomen retroperitoneum|CT Guided drainage Abdomen retroperitoneum
C0801762|T102|relax|41809-5|LNC|US Guided drainage Abdomen retroperitoneum|US Guided drainage Abdomen retroperitoneum
C0801762|T102|relax|35914-1|LNC|CT Guided drainage Anus|CT Guided drainage Anus
C0801762|T102|relax|35915-8|LNC|CT Guided drainage Appendix|CT Guided drainage Appendix
C0801762|T102|relax|36770-6|LNC|CT Guided drainage Biliary ducts Gallbladder|CT Guided drainage Biliary ducts Gallbladder
C0801762|T102|relax|35916-6|LNC|CT Guided drainage Chest|CT Guided drainage Chest
C0801762|T102|relax|69078-4|LNC|Fluoroscopy Guided drainage Chest|Fluoroscopy Guided drainage Chest
C0801762|T102|relax|24692-6|LNC|US Guided drainage Extremity|US Guided drainage Extremity
C0801762|T102|relax|26325-1|LNC|US Guided drainage Extremity bilateral|US Guided drainage Extremity bilateral
C0801762|T102|relax|26326-9|LNC|US Guided drainage Extremity left|US Guided drainage Extremity left
C0801762|T102|relax|26327-7|LNC|US Guided drainage Extremity right|US Guided drainage Extremity right
C0801762|T102|relax|35917-4|LNC|CT Guided drainage Gallbladder|CT Guided drainage Gallbladder
C0801762|T102|relax|69133-7|LNC|Fluoroscopy Guided drainage Hip|Fluoroscopy Guided drainage Hip
C0801762|T102|relax|35918-2|LNC|CT Guided drainage Kidney|CT Guided drainage Kidney
C0801762|T102|relax|24896-3|LNC|US Guided drainage Kidney|US Guided drainage Kidney
C0801762|T102|relax|26328-5|LNC|US Guided drainage Kidney bilateral|US Guided drainage Kidney bilateral
C0801762|T102|relax|26329-3|LNC|US Guided drainage Kidney left|US Guided drainage Kidney left
C0801762|T102|relax|26330-1|LNC|US Guided drainage Kidney right|US Guided drainage Kidney right
C0801762|T102|relax|35919-0|LNC|CT Guided drainage Liver|CT Guided drainage Liver
C0801762|T102|relax|35920-8|LNC|CT Guided drainage Lymph node|CT Guided drainage Lymph node
C0801762|T102|relax|42283-2|LNC|CT Guided drainage Pancreas|CT Guided drainage Pancreas
C0801762|T102|relax|44172-5|LNC|US Guided drainage Pancreas|US Guided drainage Pancreas
C0801762|T102|relax|35921-6|LNC|CT Guided drainage Pelvis|CT Guided drainage Pelvis
C0801762|T102|relax|24868-2|LNC|US Guided drainage Pelvis|US Guided drainage Pelvis
C0801762|T102|relax|41800-4|LNC|Fluoroscopy Guided drainage Pharynx|Fluoroscopy Guided drainage Pharynx
C0801762|T102|relax|41798-0|LNC|US Guided drainage Prostate|US Guided drainage Prostate
C0801762|T102|relax|35922-4|LNC|CT Guided drainage Unspecified body region|CT Guided drainage Unspecified body region
C0801762|T102|relax|30699-3|LNC|US Guided drainage Unspecified body region|US Guided drainage Unspecified body region
C0801762|T102|relax|43537-0|LNC|Fluoroscopy Guided drainage Unspecified body region|Fluoroscopy Guided drainage Unspecified body region
C0801762|T102|relax|42478-8|LNC|US Guided drainage cyst Kidney|US Guided drainage cyst Kidney
C0801762|T102|relax|46291-1|LNC|CT Guided drainage Unspecified body region-- W WO contrast IV|CT Guided drainage Unspecified body region-- W WO contrast IV
C0801762|T102|relax|35923-2|LNC|CT Guided drainage Chest-- W contrast IV|CT Guided drainage Chest-- W contrast IV
C0801762|T102|relax|46292-9|LNC|CT Guided drainage Unspecified body region-- W contrast IV|CT Guided drainage Unspecified body region-- W contrast IV
C0801762|T102|relax|35924-0|LNC|CT Guided drainage Chest-- WO contrast|CT Guided drainage Chest-- WO contrast
C0801762|T102|relax|46293-7|LNC|CT Guided drainage Unspecified body region-- WO contrast|CT Guided drainage Unspecified body region-- WO contrast
C0801762|T102|relax|35925-7|LNC|Fluoroscopy Guided endoscopy Stomach|Fluoroscopy Guided endoscopy Stomach
C0801762|T102|relax|43478-7|LNC|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 1 5 hours post contrast retrograde|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 1 5 hours post contrast retrograde
C0801762|T102|relax|43474-6|LNC|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 15 minutes post contrast retrograde|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 15 minutes post contrast retrograde
C0801762|T102|relax|43477-9|LNC|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 1 hour post contrast retrograde|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 1 hour post contrast retrograde
C0801762|T102|relax|43473-8|LNC|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 2 hours post contrast retrograde|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 2 hours post contrast retrograde
C0801762|T102|relax|43475-3|LNC|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 30 minutes post contrast retrograde|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 30 minutes post contrast retrograde
C0801762|T102|relax|43476-1|LNC|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 45 minutes post contrast retrograde|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- 45 minutes post contrast retrograde
C0801762|T102|relax|72248-8|LNC|Abdomen MRCP with without contrast IV|Abdomen MRCP with without contrast IV
C0801762|T102|relax|44214-5|LNC|Fluoroscopy Guided endoscopy Biliary ducts-- W contrast retrograde|Fluoroscopy Guided endoscopy Biliary ducts-- W contrast retrograde
C0801762|T102|relax|30815-5|LNC|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- W contrast retrograde|Fluoroscopy Guided endoscopy Biliary ducts Pancreatic duct-- W contrast retrograde
C0801762|T102|relax|44213-7|LNC|Fluoroscopy Guided endoscopy Pancreatic duct-- W contrast retrograde|Fluoroscopy Guided endoscopy Pancreatic duct-- W contrast retrograde
C0801762|T102|relax|58740-2|LNC|Abdomen MRCP WO contrast|Abdomen MRCP WO contrast
C0801762|T102|relax|72541-6|LNC|Fluoroscopy Guided facet joint denervation Spine Cervical|Fluoroscopy Guided facet joint denervation Spine Cervical
C0801762|T102|relax|72542-4|LNC|Fluoroscopy Guided facet joint denervation Spine Lumbar|Fluoroscopy Guided facet joint denervation Spine Lumbar
C0801762|T102|relax|72540-8|LNC|Fluoroscopy Guided facet joint denervation Spine|Fluoroscopy Guided facet joint denervation Spine
C0801762|T102|relax|35926-5|LNC|Fluoroscopy Guided gastrostomy Stomach|Fluoroscopy Guided gastrostomy Stomach
C0801762|T102|relax|30638-1|LNC|Fluoroscopy Guided injection Hip|Fluoroscopy Guided injection Hip
C0801762|T102|relax|24769-2|LNC|CT Guided injection Joint space|CT Guided injection Joint space
C0801762|T102|relax|42334-3|LNC|Fluoroscopy Guided injection Mammary artery internal left|Fluoroscopy Guided injection Mammary artery internal left
C0801762|T102|relax|42706-2|LNC|US Guided injection Pleural space|US Guided injection Pleural space
C0801762|T102|relax|24901-1|LNC|CT Guided injection Sacroiliac Joint|CT Guided injection Sacroiliac Joint
C0801762|T102|relax|35927-3|LNC|Fluoroscopy Guided injection Sacroiliac Joint|Fluoroscopy Guided injection Sacroiliac Joint
C0801762|T102|relax|26319-4|LNC|CT Guided injection Sacroiliac joint bilateral|CT Guided injection Sacroiliac joint bilateral
C0801762|T102|relax|26320-2|LNC|CT Guided injection Sacroiliac joint left|CT Guided injection Sacroiliac joint left
C0801762|T102|relax|26321-0|LNC|CT Guided injection Sacroiliac joint right|CT Guided injection Sacroiliac joint right
C0801762|T102|relax|48435-2|LNC|Fluoroscopy Guided injection Salivary gland bilateral|Fluoroscopy Guided injection Salivary gland bilateral
C0801762|T102|relax|46392-7|LNC|Fluoroscopy Guided injection Sinuses|Fluoroscopy Guided injection Sinuses
C0801762|T102|relax|30579-7|LNC|CT Guided injection Spine facet joint|CT Guided injection Spine facet joint
C0801762|T102|relax|24931-8|LNC|Fluoroscopy Guided injection Spine facet joint|Fluoroscopy Guided injection Spine facet joint
C0801762|T102|relax|26322-8|LNC|Fluoroscopy Guided injection Spine facet joint bilateral|Fluoroscopy Guided injection Spine facet joint bilateral
C0801762|T102|relax|26323-6|LNC|Fluoroscopy Guided injection Spine facet joint left|Fluoroscopy Guided injection Spine facet joint left
C0801762|T102|relax|26324-4|LNC|Fluoroscopy Guided injection Spine facet joint right|Fluoroscopy Guided injection Spine facet joint right
C0801762|T102|relax|70918-8|LNC|Fluoroscopy Guided injection Spine Cervical|Fluoroscopy Guided injection Spine Cervical
C0801762|T102|relax|30812-2|LNC|Fluoroscopy Guided injection Spine Cervical Facet Joint|Fluoroscopy Guided injection Spine Cervical Facet Joint
C0801762|T102|relax|37493-4|LNC|CT Guided injection Spine disc cervical|CT Guided injection Spine disc cervical
C0801762|T102|relax|70919-6|LNC|Fluoroscopy Guided injection Spine Lumbar|Fluoroscopy Guided injection Spine Lumbar
C0801762|T102|relax|30817-1|LNC|Fluoroscopy Guided injection Spine Lumbar Facet Joint|Fluoroscopy Guided injection Spine Lumbar Facet Joint
C0801762|T102|relax|70920-4|LNC|Fluoroscopy Guided injection Spine Thoracic|Fluoroscopy Guided injection Spine Thoracic
C0801762|T102|relax|30814-8|LNC|Fluoroscopy Guided injection Spine Thoracic Facet Joint|Fluoroscopy Guided injection Spine Thoracic Facet Joint
C0801762|T102|relax|30702-5|LNC|US Guided injection Thyroid|US Guided injection Thyroid
C0801762|T102|relax|72530-9|LNC|US Guided injection Joint|US Guided injection Joint
C0801762|T102|relax|36771-4|LNC|Fluoroscopy Guided injection Joint|Fluoroscopy Guided injection Joint
C0801762|T102|relax|37494-2|LNC|Fluoroscopy Guided injection Tendon|Fluoroscopy Guided injection Tendon
C0801762|T102|relax|72537-4|LNC|US Guided injection sclerosing agent Extremity vein bilateral|US Guided injection sclerosing agent Extremity vein bilateral
C0801762|T102|relax|72645-5|LNC|US Guided injection sclerosing agent Extremity vein left|US Guided injection sclerosing agent Extremity vein left
C0801762|T102|relax|72644-8|LNC|US Guided injection sclerosing agent Extremity vein right|US Guided injection sclerosing agent Extremity vein right
C0801762|T102|relax|72536-6|LNC|US Guided injection sclerosing agent Extremity veins bilateral|US Guided injection sclerosing agent Extremity veins bilateral
C0801762|T102|relax|72643-0|LNC|US Guided injection sclerosing agent Extremity veins left|US Guided injection sclerosing agent Extremity veins left
C0801762|T102|relax|72642-2|LNC|US Guided injection sclerosing agent Extremity veins right|US Guided injection sclerosing agent Extremity veins right
C0801762|T102|relax|72543-2|LNC|Fluoroscopy Guided intercostal nerve devervation Spine Thoracic|Fluoroscopy Guided intercostal nerve devervation Spine Thoracic
C0801762|T102|relax|72552-3|LNC|Fluoroscopy Guided kyphoplasty Spine Lumbar|Fluoroscopy Guided kyphoplasty Spine Lumbar
C0801762|T102|relax|72553-1|LNC|Fluoroscopy Guided kyphoplasty Spine Thoracic|Fluoroscopy Guided kyphoplasty Spine Thoracic
C0801762|T102|relax|72535-8|LNC|US Guided laser ablation vein(s) Extremity vein left|US Guided laser ablation vein(s) Extremity vein left
C0801762|T102|relax|72534-1|LNC|US Guided laser ablation vein(s) Extremity vein right|US Guided laser ablation vein(s) Extremity vein right
C0801762|T102|relax|48735-5|LNC|Mammogram Guided localization Breast|Mammogram Guided localization Breast
C0801762|T102|relax|43759-0|LNC|US Guided localization Breast bilateral|US Guided localization Breast bilateral
C0801762|T102|relax|35928-1|LNC|CT Guided localization Breast left|CT Guided localization Breast left
C0801762|T102|relax|42296-4|LNC|Mammogram Guided localization Breast left|Mammogram Guided localization Breast left
C0801762|T102|relax|43758-2|LNC|US Guided localization Breast left|US Guided localization Breast left
C0801762|T102|relax|35929-9|LNC|CT Guided localization Breast right|CT Guided localization Breast right
C0801762|T102|relax|42297-2|LNC|Mammogram Guided localization Breast right|Mammogram Guided localization Breast right
C0801762|T102|relax|43760-8|LNC|US Guided localization Breast right|US Guided localization Breast right
C0801762|T102|relax|37608-7|LNC|US Guided localization foreign body Eye|US Guided localization foreign body Eye
C0801762|T102|relax|42701-3|LNC|CT Guided localization placenta Uterus|CT Guided localization placenta Uterus
C0801762|T102|relax|39760-4|LNC|Scan Guided localization tumor limited|Scan Guided localization tumor limited
C0801762|T102|relax|39759-6|LNC|SPECT Guided localization tumor limited|SPECT Guided localization tumor limited
C0801762|T102|relax|39761-2|LNC|Scan Guided localization tumor limited-- W Tc-99m Sestamibi IV|Scan Guided localization tumor limited-- W Tc-99m Sestamibi IV
C0801762|T102|relax|39953-5|LNC|Scan Guided localization tumor multiple areas|Scan Guided localization tumor multiple areas
C0801762|T102|relax|39763-8|LNC|Scan Guided localization tumor|Scan Guided localization tumor
C0801762|T102|relax|39762-0|LNC|SPECT Guided localization tumor|SPECT Guided localization tumor
C0801762|T102|relax|39758-8|LNC|Scan Guided localization tumor Breast|Scan Guided localization tumor Breast
C0801762|T102|relax|44110-5|LNC|CT Guided needle localization Breast|CT Guided needle localization Breast
C0801762|T102|relax|24600-9|LNC|US Guided needle localization Breast|US Guided needle localization Breast
C0801762|T102|relax|69068-5|LNC|Mammogram Guided needle localization Breast bilateral|Mammogram Guided needle localization Breast bilateral
C0801762|T102|relax|26313-7|LNC|US Guided needle localization Breast bilateral|US Guided needle localization Breast bilateral
C0801762|T102|relax|26314-5|LNC|US Guided needle localization Breast left|US Guided needle localization Breast left
C0801762|T102|relax|26318-6|LNC|US Guided needle localization Breast right|US Guided needle localization Breast right
C0801762|T102|relax|37921-4|LNC|US Guided needle localization Chest|US Guided needle localization Chest
C0801762|T102|relax|42021-6|LNC|CT Guided needle localization Spine Cervical|CT Guided needle localization Spine Cervical
C0801762|T102|relax|42020-8|LNC|CT Guided needle localization Spine Lumbar|CT Guided needle localization Spine Lumbar
C0801762|T102|relax|39026-0|LNC|CT Guided needle localization Unspecified body region|CT Guided needle localization Unspecified body region
C0801762|T102|relax|39028-6|LNC|MRI Guided needle localization Unspecified body region|MRI Guided needle localization Unspecified body region
C0801762|T102|relax|38032-9|LNC|US Guided needle localization Unspecified body region|US Guided needle localization Unspecified body region
C0801762|T102|relax|39027-8|LNC|Fluoroscopy Guided needle localization Unspecified body region|Fluoroscopy Guided needle localization Unspecified body region
C0801762|T102|relax|24595-1|LNC|Mammogram Guided needle localization mass Breast|Mammogram Guided needle localization mass Breast
C0801762|T102|relax|26315-2|LNC|Mammogram Guided needle localization mass Breast bilateral|Mammogram Guided needle localization mass Breast bilateral
C0801762|T102|relax|26316-0|LNC|Mammogram Guided needle localization mass Breast left|Mammogram Guided needle localization mass Breast left
C0801762|T102|relax|26317-8|LNC|Mammogram Guided needle localization mass Breast right|Mammogram Guided needle localization mass Breast right
C0801762|T102|relax|44118-8|LNC|CT Guided needle localization Breast-- W WO contrast IV|CT Guided needle localization Breast-- W WO contrast IV
C0801762|T102|relax|35930-7|LNC|CT Guided nerve block Abdomen|CT Guided nerve block Abdomen
C0801762|T102|relax|35931-5|LNC|CT Guided nerve block Pelvis|CT Guided nerve block Pelvis
C0801762|T102|relax|70921-2|LNC|CT Guided nerve block Spine Cervical|CT Guided nerve block Spine Cervical
C0801762|T102|relax|35932-3|LNC|CT Guided nerve block Spine Lumbar|CT Guided nerve block Spine Lumbar
C0801762|T102|relax|70922-0|LNC|CT Guided nerve block Spine Thoracic|CT Guided nerve block Spine Thoracic
C0801762|T102|relax|69240-0|LNC|Fluoroscopy Guided percutaneous biopsy Abdomen|Fluoroscopy Guided percutaneous biopsy Abdomen
C0801762|T102|relax|42139-6|LNC|US Guided percutaneous biopsy Muscle|US Guided percutaneous biopsy Muscle
C0801762|T102|relax|24609-0|LNC|Mammogram Guided core needle percutaneous biopsy Breast|Mammogram Guided core needle percutaneous biopsy Breast
C0801762|T102|relax|26334-3|LNC|Mammogram Guided core needle percutaneous biopsy Breast bilateral|Mammogram Guided core needle percutaneous biopsy Breast bilateral
C0801762|T102|relax|26335-0|LNC|Mammogram Guided core needle percutaneous biopsy Breast left|Mammogram Guided core needle percutaneous biopsy Breast left
C0801762|T102|relax|38023-8|LNC|US Guided core needle percutaneous biopsy Breast left|US Guided core needle percutaneous biopsy Breast left
C0801762|T102|relax|26336-8|LNC|Mammogram Guided core needle percutaneous biopsy Breast right|Mammogram Guided core needle percutaneous biopsy Breast right
C0801762|T102|relax|38025-3|LNC|US Guided core needle percutaneous biopsy Breast right|US Guided core needle percutaneous biopsy Breast right
C0801762|T102|relax|44121-2|LNC|Mammogram Guided percutaneous needle biopsy Breast|Mammogram Guided percutaneous needle biopsy Breast
C0801762|T102|relax|69245-9|LNC|Fluoroscopy Guided percutaneous needle biopsy Kidney|Fluoroscopy Guided percutaneous needle biopsy Kidney
C0801762|T102|relax|69246-7|LNC|Fluoroscopy Guided percutaneous needle biopsy Liver|Fluoroscopy Guided percutaneous needle biopsy Liver
C0801762|T102|relax|44204-6|LNC|Fluoroscopy Guided percutaneous needle biopsy Lung|Fluoroscopy Guided percutaneous needle biopsy Lung
C0801762|T102|relax|69247-5|LNC|Fluoroscopy Guided percutaneous needle biopsy Salivary gland|Fluoroscopy Guided percutaneous needle biopsy Salivary gland
C0801762|T102|relax|46372-9|LNC|Fluoroscopy Guided percutaneous drainage Biliary ducts|Fluoroscopy Guided percutaneous drainage Biliary ducts
C0801762|T102|relax|62494-0|LNC|US Guided percutaneous drainage Cavity|US Guided percutaneous drainage Cavity
C0801762|T102|relax|24621-5|LNC|Fluoroscopy Guided percutaneous drainage Cavity|Fluoroscopy Guided percutaneous drainage Cavity
C0801762|T102|relax|69241-8|LNC|Fluoroscopy Guided percutaneous drainage abscess Abdomen|Fluoroscopy Guided percutaneous drainage abscess Abdomen
C0801762|T102|relax|69242-6|LNC|Fluoroscopy Guided percutaneous drainage abscess Appendix|Fluoroscopy Guided percutaneous drainage abscess Appendix
C0801762|T102|relax|42422-6|LNC|Fluoroscopy Guided percutaneous drainage abscess Breast|Fluoroscopy Guided percutaneous drainage abscess Breast
C0801762|T102|relax|43444-9|LNC|CT Guided percutaneous drainage abscess Cavity|CT Guided percutaneous drainage abscess Cavity
C0801762|T102|relax|42423-4|LNC|Fluoroscopy Guided percutaneous drainage abscess Chest|Fluoroscopy Guided percutaneous drainage abscess Chest
C0801762|T102|relax|69243-4|LNC|Fluoroscopy Guided percutaneous drainage abscess Lung|Fluoroscopy Guided percutaneous drainage abscess Lung
C0801762|T102|relax|44223-6|LNC|Fluoroscopy Guided percutaneous drainage abscess Ovary|Fluoroscopy Guided percutaneous drainage abscess Ovary
C0801762|T102|relax|69244-2|LNC|Fluoroscopy Guided percutaneous drainage abscess Pelvis|Fluoroscopy Guided percutaneous drainage abscess Pelvis
C0801762|T102|relax|42421-8|LNC|Fluoroscopy Guided percutaneous drainage abscess Unspecified body region|Fluoroscopy Guided percutaneous drainage abscess Unspecified body region
C0801762|T102|relax|70923-8|LNC|Fluoroscopy Guided percutaneous vertebroplasty Spine Cervical|Fluoroscopy Guided percutaneous vertebroplasty Spine Cervical
C0801762|T102|relax|35934-9|LNC|CT Guided percutaneous vertebroplasty Spine Lumbar|CT Guided percutaneous vertebroplasty Spine Lumbar
C0801762|T102|relax|70924-6|LNC|Fluoroscopy Guided percutaneous vertebroplasty Spine Lumbar|Fluoroscopy Guided percutaneous vertebroplasty Spine Lumbar
C0801762|T102|relax|35935-6|LNC|CT Guided percutaneous vertebroplasty Spine Thoracic|CT Guided percutaneous vertebroplasty Spine Thoracic
C0801762|T102|relax|70925-3|LNC|Fluoroscopy Guided percutaneous vertebroplasty Spine Thoracic|Fluoroscopy Guided percutaneous vertebroplasty Spine Thoracic
C0801762|T102|relax|72539-0|LNC|Fluoroscopy Guided peripheral nerve denervation Unspecified body region|Fluoroscopy Guided peripheral nerve denervation Unspecified body region
C0801762|T102|relax|30643-1|LNC|US Guided placement catheter in Central vein|US Guided placement catheter in Central vein
C0801762|T102|relax|35912-5|LNC|Fluoroscopy Guided placement catheter in Unspecified body region|Fluoroscopy Guided placement catheter in Unspecified body region
C0801762|T102|relax|25028-2|LNC|Fluoroscopic angiogram Guided placement catheter adminstration thrombolytic in Vessel|Fluoroscopic angiogram Guided placement catheter adminstration thrombolytic in Vessel
C0801762|T102|relax|25029-0|LNC|Fluoroscopic angiogram Guided placement catheter vasoconstrictor infusion in Vessels|Fluoroscopic angiogram Guided placement catheter vasoconstrictor infusion in Vessels
C0801762|T102|relax|24613-2|LNC|Fluoroscopic angiogram Guided placement catheter in artery in Central cardiovascular artery|Fluoroscopic angiogram Guided placement catheter in artery in Central cardiovascular artery
C0801762|T102|relax|30644-9|LNC|US Guided placement catheter in Central vein-- Tunneled|US Guided placement catheter in Central vein-- Tunneled
C0801762|T102|relax|25077-9|LNC|Fluoroscopic angiogram Guided placement catheter in Hepatic artery-- W contrast IA|Fluoroscopic angiogram Guided placement catheter in Hepatic artery-- W contrast IA
C0801762|T102|relax|24625-6|LNC|Fluoroscopic angiogram Guided placement catheter in Central vein-- W contrast IV|Fluoroscopic angiogram Guided placement catheter in Central vein-- W contrast IV
C0801762|T102|relax|26310-3|LNC|Fluoroscopic angiogram Guided placement catheter in Central vein bilateral-- W contrast IV|Fluoroscopic angiogram Guided placement catheter in Central vein bilateral-- W contrast IV
C0801762|T102|relax|26311-1|LNC|Fluoroscopic angiogram Guided placement catheter in Central vein left-- W contrast IV|Fluoroscopic angiogram Guided placement catheter in Central vein left-- W contrast IV
C0801762|T102|relax|26312-9|LNC|Fluoroscopic angiogram Guided placement catheter in Central vein right-- W contrast IV|Fluoroscopic angiogram Guided placement catheter in Central vein right-- W contrast IV
C0801762|T102|relax|41801-2|LNC|Fluoroscopic angiogram Guided placement catheter in Portal vein-- W contrast IV|Fluoroscopic angiogram Guided placement catheter in Portal vein-- W contrast IV
C0801762|T102|relax|24716-3|LNC|Fluoroscopy Guided placement decompression tube in Gastrointestine|Fluoroscopy Guided placement decompression tube in Gastrointestine
C0801762|T102|relax|62491-6|LNC|Fluoroscopic angiogram Guided placement ilio-iliac tube endoprosthesis in Iliac artery left-- W contrast IA|Fluoroscopic angiogram Guided placement ilio-iliac tube endoprosthesis in Iliac artery left-- W contrast IA
C0801762|T102|relax|62492-4|LNC|Fluoroscopic angiogram Guided placement ilio-iliac tube endoprosthesis in Iliac artery right-- W contrast IA|Fluoroscopic angiogram Guided placement ilio-iliac tube endoprosthesis in Iliac artery right-- W contrast IA
C0801762|T102|relax|25072-0|LNC|Guided placement infusion port in Unspecified body region|Guided placement infusion port in Unspecified body region
C0801762|T102|relax|62450-2|LNC|Fluoroscopic angiogram Guided placement intraperitoneal catheter in Abdomen|Fluoroscopic angiogram Guided placement intraperitoneal catheter in Abdomen
C0801762|T102|relax|25026-6|LNC|Fluoroscopic angiogram Guided placement IVC filter in Inferior vena cava-- W contrast IV|Fluoroscopic angiogram Guided placement IVC filter in Inferior vena cava-- W contrast IV
C0801762|T102|relax|25027-4|LNC|Guided placement large bore catheter vessel in Central vein|Guided placement large bore catheter vessel in Central vein
C0801762|T102|relax|26307-9|LNC|Guided placement large bore catheter vessel in Central vein bilateral|Guided placement large bore catheter vessel in Central vein bilateral
C0801762|T102|relax|26308-7|LNC|Guided placement large bore catheter vessel in Central vein left|Guided placement large bore catheter vessel in Central vein left
C0801762|T102|relax|26309-5|LNC|Guided placement large bore catheter vessel in Central vein right|Guided placement large bore catheter vessel in Central vein right
C0801762|T102|relax|25024-1|LNC|Fluoroscopic angiogram Guided placement longterm peripheral catheter in Central vein|Fluoroscopic angiogram Guided placement longterm peripheral catheter in Central vein
C0801762|T102|relax|26304-6|LNC|Fluoroscopic angiogram Guided placement longterm peripheral catheter in Central vein bilateral|Fluoroscopic angiogram Guided placement longterm peripheral catheter in Central vein bilateral
C0801762|T102|relax|26305-3|LNC|Fluoroscopic angiogram Guided placement longterm peripheral catheter in Central vein left|Fluoroscopic angiogram Guided placement longterm peripheral catheter in Central vein left
C0801762|T102|relax|26306-1|LNC|Fluoroscopic angiogram Guided placement longterm peripheral catheter in Central vein right|Fluoroscopic angiogram Guided placement longterm peripheral catheter in Central vein right
C0801762|T102|relax|64993-9|LNC|US Guided placement needle in Unspecified body region|US Guided placement needle in Unspecified body region
C0801762|T102|relax|42456-4|LNC|US Guided placement needle wire in Breast|US Guided placement needle wire in Breast
C0801762|T102|relax|36772-2|LNC|CT Guided placement nephrostomy tube in Kidney|CT Guided placement nephrostomy tube in Kidney
C0801762|T102|relax|24779-1|LNC|Fluoroscopy Guided placement percutaneous nephrostomy in Kidney bilateral-- W contrast via tube|Fluoroscopy Guided placement percutaneous nephrostomy in Kidney bilateral-- W contrast via tube
C0801762|T102|relax|24782-5|LNC|Fluoroscopy Guided placement percutaneous nephroureteral stent in Kidney bilateral|Fluoroscopy Guided placement percutaneous nephroureteral stent in Kidney bilateral
C0801762|T102|relax|35937-2|LNC|CT Guided placement radiation therapy fields in Unspecified body region|CT Guided placement radiation therapy fields in Unspecified body region
C0801762|T102|relax|43487-8|LNC|US Guided placement radiation therapy fields in Unspecified body region|US Guided placement radiation therapy fields in Unspecified body region
C0801762|T102|relax|65797-3|LNC|Fluoroscopic angiogram Guided placement stent in Artery left|Fluoroscopic angiogram Guided placement stent in Artery left
C0801762|T102|relax|65798-1|LNC|Fluoroscopic angiogram Guided placement stent in Artery right|Fluoroscopic angiogram Guided placement stent in Artery right
C0801762|T102|relax|69134-5|LNC|Fluoroscopic angiogram Guided placement stent in Iliac artery|Fluoroscopic angiogram Guided placement stent in Iliac artery
C0801762|T102|relax|25078-7|LNC|Fluoroscopy Guided placement stent in Intrahepatic portal system|Fluoroscopy Guided placement stent in Intrahepatic portal system
C0801762|T102|relax|24756-9|LNC|Fluoroscopic angiogram Guided placement stent in Vein|Fluoroscopic angiogram Guided placement stent in Vein
C0801762|T102|relax|26301-2|LNC|Fluoroscopic angiogram Guided placement stent in Vein bilateral|Fluoroscopic angiogram Guided placement stent in Vein bilateral
C0801762|T102|relax|26302-0|LNC|Fluoroscopic angiogram Guided placement stent in Vein left|Fluoroscopic angiogram Guided placement stent in Vein left
C0801762|T102|relax|26303-8|LNC|Fluoroscopic angiogram Guided placement stent in Vein right|Fluoroscopic angiogram Guided placement stent in Vein right
C0801762|T102|relax|24555-5|LNC|Fluoroscopic angiogram Guided placement stent in Artery|Fluoroscopic angiogram Guided placement stent in Artery
C0801762|T102|relax|51391-1|LNC|Fluoroscopic angiogram Guided placement transjugular intrahepatic portosystemic shunt in Portal vein Hepatic vein|Fluoroscopic angiogram Guided placement transjugular intrahepatic portosystemic shunt in Portal vein Hepatic vein
C0801762|T102|relax|35938-0|LNC|CT Guided placement tube in Chest|CT Guided placement tube in Chest
C0801762|T102|relax|42140-4|LNC|US Guided placement tube in Chest|US Guided placement tube in Chest
C0801762|T102|relax|39362-9|LNC|Fluoroscopy Guided placement tube in Chest|Fluoroscopy Guided placement tube in Chest
C0801762|T102|relax|30637-3|LNC|Fluoroscopy Guided placement tube in Gastrointestine|Fluoroscopy Guided placement tube in Gastrointestine
C0801762|T102|relax|41799-8|LNC|Fluoroscopy Guided placement tube in Liver|Fluoroscopy Guided placement tube in Liver
C0801762|T102|relax|24995-3|LNC|Fluoroscopy Guided placement tube in Stomach|Fluoroscopy Guided placement tube in Stomach
C0801762|T102|relax|44224-4|LNC|Fluoroscopy Guided placement tube in Unspecified body region|Fluoroscopy Guided placement tube in Unspecified body region
C0801762|T102|relax|46373-7|LNC|SPECT Guided placement tube in Chest|SPECT Guided placement tube in Chest
C0801762|T102|relax|44102-2|LNC|CT Guided procedure Joint space|CT Guided procedure Joint space
C0801762|T102|relax|44222-8|LNC|Fluoroscopy Guided procedure Joint space|Fluoroscopy Guided procedure Joint space
C0801762|T102|relax|30629-0|LNC|Fluoroscopy Guided procedure Unspecified body region|Fluoroscopy Guided procedure Unspecified body region
C0801762|T102|relax|30581-3|LNC|CT Guided radiation treatment Unspecified body region-- W contrast IV|CT Guided radiation treatment Unspecified body region-- W contrast IV
C0801762|T102|relax|30664-7|LNC|MRI Guided radiation treatment Unspecified body region-- W contrast IV|MRI Guided radiation treatment Unspecified body region-- W contrast IV
C0801762|T102|relax|30582-1|LNC|CT Guided radiation treatment Unspecified body region-- WO contrast|CT Guided radiation treatment Unspecified body region-- WO contrast
C0801762|T102|relax|30665-4|LNC|MRI Guided radiation treatment Unspecified body region-- WO contrast|MRI Guided radiation treatment Unspecified body region-- WO contrast
C0801762|T102|relax|25053-0|LNC|CT Guided radiosurgery Unspecified body region|CT Guided radiosurgery Unspecified body region
C0801762|T102|relax|25054-8|LNC|CT Guided radiosurgery Unspecified body region-- W contrast IV|CT Guided radiosurgery Unspecified body region-- W contrast IV
C0801762|T102|relax|24537-3|LNC|US Guided removal amniotic fluid from Uterus|US Guided removal amniotic fluid from Uterus
C0801762|T102|relax|42141-2|LNC|US Guided removal catheter from Central vein-- Tunneled|US Guided removal catheter from Central vein-- Tunneled
C0801762|T102|relax|72549-9|LNC|Fluoroscopy Guided removal catheter from Central vein-- Tunneled|Fluoroscopy Guided removal catheter from Central vein-- Tunneled
C0801762|T102|relax|72548-1|LNC|Fluoroscopic angiogram Guided removal catheter from Central vein-- W contrast IV|Fluoroscopic angiogram Guided removal catheter from Central vein-- W contrast IV
C0801762|T102|relax|72547-3|LNC|Fluoroscopy Guided removal CVA device obstruction from Central vein|Fluoroscopy Guided removal CVA device obstruction from Central vein
C0801762|T102|relax|72546-5|LNC|Fluoroscopy Guided removal CVA lumen obstruction from Central vein|Fluoroscopy Guided removal CVA lumen obstruction from Central vein
C0801762|T102|relax|41810-3|LNC|CT Guided removal fluid from Abdomen|CT Guided removal fluid from Abdomen
C0801762|T102|relax|24559-7|LNC|US Guided removal fluid from Abdomen|US Guided removal fluid from Abdomen
C0801762|T102|relax|38142-6|LNC|US Guided removal fluid from Chest|US Guided removal fluid from Chest
C0801762|T102|relax|30628-2|LNC|Fluoroscopy Guided removal foreign body from Unspecified body region|Fluoroscopy Guided removal foreign body from Unspecified body region
C0801762|T102|relax|72538-2|LNC|Fluoroscopic angiogram Guided removal longterm peripheral catheter from Central vein|Fluoroscopic angiogram Guided removal longterm peripheral catheter from Central vein
C0801762|T102|relax|72544-0|LNC|Fluoroscopy Guided removal percutaneous nephrostomy tube from Kidney bilateral-- W contrast|Fluoroscopy Guided removal percutaneous nephrostomy tube from Kidney bilateral-- W contrast
C0801762|T102|relax|24885-6|LNC|US Guided repair Pseudoaneurysm/AV fistula|US Guided repair Pseudoaneurysm/AV fistula
C0801762|T102|relax|72550-7|LNC|Fluoroscopy Guided repair CVA catheter with port or pump Central vein|Fluoroscopy Guided repair CVA catheter with port or pump Central vein
C0801762|T102|relax|72551-5|LNC|Fluoroscopy Guided repair CVA catheter without port or pump Central vein|Fluoroscopy Guided repair CVA catheter without port or pump Central vein
C0801762|T102|relax|42017-4|LNC|Fluoroscopy Guided replacement percutaneous cholecystostomy in Abdomen|Fluoroscopy Guided replacement percutaneous cholecystostomy in Abdomen
C0801762|T102|relax|52790-3|LNC|CT Guided replacement percutaneous drainage tube in Abdomen|CT Guided replacement percutaneous drainage tube in Abdomen
C0801762|T102|relax|72545-7|LNC|Fluoroscopy Guided replacement percutaneous drainage tube in Biliary ducts Gallbladder|Fluoroscopy Guided replacement percutaneous drainage tube in Biliary ducts Gallbladder
C0801762|T102|relax|52791-1|LNC|CT Guided replacement percutaneous drainage tube in Pelvis|CT Guided replacement percutaneous drainage tube in Pelvis
C0801762|T102|relax|46294-5|LNC|Fluoroscopy Guided replacement percutaneous drainage tube in Stomach|Fluoroscopy Guided replacement percutaneous drainage tube in Stomach
C0801762|T102|relax|24996-1|LNC|Fluoroscopy Guided replacement percutaneous gastrostomy in Stomach|Fluoroscopy Guided replacement percutaneous gastrostomy in Stomach
C0801762|T102|relax|24626-4|LNC|Fluoroscopic angiogram Guided reposition catheter in Central vein-- W contrast IV|Fluoroscopic angiogram Guided reposition catheter in Central vein-- W contrast IV
C0801762|T102|relax|26295-6|LNC|Fluoroscopic angiogram Guided reposition catheter in Central vein bilateral-- W contrast IV|Fluoroscopic angiogram Guided reposition catheter in Central vein bilateral-- W contrast IV
C0801762|T102|relax|26296-4|LNC|Fluoroscopic angiogram Guided reposition catheter in Central vein left-- W contrast IV|Fluoroscopic angiogram Guided reposition catheter in Central vein left-- W contrast IV
C0801762|T102|relax|26297-2|LNC|Fluoroscopic angiogram Guided reposition catheter in Central vein right-- W contrast IV|Fluoroscopic angiogram Guided reposition catheter in Central vein right-- W contrast IV
C0801762|T102|relax|48740-5|LNC|Mammogram Guided sentinel lymph node injection Breast|Mammogram Guided sentinel lymph node injection Breast
C0801762|T102|relax|48736-3|LNC|Mammogram Guided sentinel lymph node injection Breast left|Mammogram Guided sentinel lymph node injection Breast left
C0801762|T102|relax|48739-7|LNC|Mammogram Guided sentinel lymph node injection Breast right|Mammogram Guided sentinel lymph node injection Breast right
C0801762|T102|relax|24570-4|LNC|Fluoroscopy Guided stone removal Biliary duct common-- W contrast intra biliary duct|Fluoroscopy Guided stone removal Biliary duct common-- W contrast intra biliary duct
C0801762|T102|relax|43763-2|LNC|Fluoroscopic angiogram Guided thrombectomy Vein-- W contrast IV|Fluoroscopic angiogram Guided thrombectomy Vein-- W contrast IV
C0801762|T102|relax|43761-6|LNC|Fluoroscopic angiogram Guided thrombectomy Vein bilateral-- W contrast IV|Fluoroscopic angiogram Guided thrombectomy Vein bilateral-- W contrast IV
C0801762|T102|relax|43762-4|LNC|Fluoroscopic angiogram Guided thrombectomy Vein left-- W contrast IV|Fluoroscopic angiogram Guided thrombectomy Vein left-- W contrast IV
C0801762|T102|relax|43764-0|LNC|Fluoroscopic angiogram Guided thrombectomy Vein right-- W contrast IV|Fluoroscopic angiogram Guided thrombectomy Vein right-- W contrast IV
C0801762|T102|relax|72554-9|LNC|Fluoroscopy Guided trigger point injection Muscle|Fluoroscopy Guided trigger point injection Muscle
C0801762|T102|relax|39138-3|LNC|Fluoroscopic angiogram Guided vascular access Vessel|Fluoroscopic angiogram Guided vascular access Vessel
C0801762|T102|relax|39139-1|LNC|US Guided vascular access Unspecified body region|US Guided vascular access Unspecified body region
C0801762|T102|relax|36936-3|LNC|MRI stereotactic biopsy Brain|MRI stereotactic biopsy Brain
C0801762|T102|relax|24603-3|LNC|Mammogram stereotactic biopsy Breast|Mammogram stereotactic biopsy Breast
C0801762|T102|relax|26292-3|LNC|Mammogram stereotactic biopsy Breast bilateral|Mammogram stereotactic biopsy Breast bilateral
C0801762|T102|relax|26293-1|LNC|Mammogram stereotactic biopsy Breast left|Mammogram stereotactic biopsy Breast left
C0801762|T102|relax|26294-9|LNC|Mammogram stereotactic biopsy Breast right|Mammogram stereotactic biopsy Breast right
C0801762|T102|relax|36928-0|LNC|CT stereotactic biopsy Head|CT stereotactic biopsy Head
C0801762|T102|relax|46296-0|LNC|Mammogram stereotactic core needle biopsy Breast|Mammogram stereotactic core needle biopsy Breast
C0801762|T102|relax|46295-2|LNC|Mammogram stereotactic core needle biopsy Breast left|Mammogram stereotactic core needle biopsy Breast left
C0801762|T102|relax|42433-3|LNC|Mammogram stereotactic core needle biopsy Breast right|Mammogram stereotactic core needle biopsy Breast right
C0801762|T102|relax|69160-0|LNC|Mammogram stereotactic needle biopsy Breast|Mammogram stereotactic needle biopsy Breast
C0801762|T102|relax|24585-2|LNC|CT stereotactic biopsy Head-- W contrast IV|CT stereotactic biopsy Head-- W contrast IV
C0801762|T102|relax|36929-8|LNC|CT stereotactic biopsy Head-- WO contrast|CT stereotactic biopsy Head-- WO contrast
C0801762|T102|relax|44122-0|LNC|MRI stereotactic localization in Brain-- W WO contrast IV|MRI stereotactic localization in Brain-- W WO contrast IV
C0801762|T102|relax|30656-3|LNC|MRI stereotactic localization in Brain-- W contrast IV|MRI stereotactic localization in Brain-- W contrast IV
C0801762|T102|relax|30800-7|LNC|MRI stereotactic localization in Brain-- WO contrast|MRI stereotactic localization in Brain-- WO contrast
C0801762|T102|relax|24655-3|LNC|Chest Fluoroscopy Image intensifier during surgery|Chest Fluoroscopy Image intensifier during surgery
C0801762|T102|relax|24717-1|LNC|Ileal conduit X-ray Loopogram|Ileal conduit X-ray Loopogram
C0801762|T102|relax|24672-8|LNC|Diaphragm US Motion|Diaphragm US Motion
C0801762|T102|relax|30632-4|LNC|Diaphragm Fluoroscopy Motion|Diaphragm Fluoroscopy Motion
C0801762|T102|relax|35990-1|LNC|Fetal MRI|Fetal MRI
C0801762|T102|relax|41806-1|LNC|Abdomen CT|Abdomen CT
C0801762|T102|relax|24556-3|LNC|Abdomen MRI|Abdomen MRI
C0801762|T102|relax|24558-9|LNC|Abdomen US|Abdomen US
C0801762|T102|relax|30762-9|LNC|Abdomen X-ray tomograph|Abdomen X-ray tomograph
C0801762|T102|relax|24566-2|LNC|Abdomen retroperitoneum CT|Abdomen retroperitoneum CT
C0801762|T102|relax|24531-6|LNC|Abdomen retroperitoneum US|Abdomen retroperitoneum US
C0801762|T102|relax|24532-4|LNC|Abdomen RUQ US|Abdomen RUQ US
C0801762|T102|relax|44115-4|LNC|Abdomen Pelvis CT|Abdomen Pelvis CT
C0801762|T102|relax|36781-3|LNC|Abdominal veins MRI angiogram|Abdominal veins MRI angiogram
C0801762|T102|relax|30864-3|LNC|Abdominal veins IVC MRI angiogram|Abdominal veins IVC MRI angiogram
C0801762|T102|relax|36791-2|LNC|Abdominal vessels MRI angiogram|Abdominal vessels MRI angiogram
C0801762|T102|relax|24534-0|LNC|Abdominal vessels US doppler|Abdominal vessels US doppler
C0801762|T102|relax|39494-0|LNC|Abdominal wall US|Abdominal wall US
C0801762|T102|relax|36930-6|LNC|Adrenal gland CT|Adrenal gland CT
C0801762|T102|relax|36931-4|LNC|Adrenal gland MRI|Adrenal gland MRI
C0801762|T102|relax|69277-2|LNC|Adrenal gland US|Adrenal gland US
C0801762|T102|relax|36792-0|LNC|Adrenal vessels MRI angiogram|Adrenal vessels MRI angiogram
C0801762|T102|relax|35940-6|LNC|Ankle CT|Ankle CT
C0801762|T102|relax|24538-1|LNC|Ankle MRI|Ankle MRI
C0801762|T102|relax|35939-8|LNC|Ankle X-ray tomograph|Ankle X-ray tomograph
C0801762|T102|relax|35941-4|LNC|Ankle bilateral CT|Ankle bilateral CT
C0801762|T102|relax|26208-9|LNC|Ankle bilateral MRI|Ankle bilateral MRI
C0801762|T102|relax|35942-2|LNC|Ankle left CT|Ankle left CT
C0801762|T102|relax|26209-7|LNC|Ankle left MRI|Ankle left MRI
C0801762|T102|relax|35943-0|LNC|Ankle left X-ray tomograph|Ankle left X-ray tomograph
C0801762|T102|relax|35944-8|LNC|Ankle right CT|Ankle right CT
C0801762|T102|relax|26210-5|LNC|Ankle right MRI|Ankle right MRI
C0801762|T102|relax|37674-9|LNC|Ankle right X-ray tomograph|Ankle right X-ray tomograph
C0801762|T102|relax|37222-7|LNC|Ankle Foot MRI|Ankle Foot MRI
C0801762|T102|relax|24542-3|LNC|Anus US|Anus US
C0801762|T102|relax|35945-5|LNC|Aorta CT|Aorta CT
C0801762|T102|relax|35947-1|LNC|Aorta MRI|Aorta MRI
C0801762|T102|relax|35946-3|LNC|Aorta MRI angiogram|Aorta MRI angiogram
C0801762|T102|relax|24547-2|LNC|Aorta US|Aorta US
C0801762|T102|relax|46388-5|LNC|Aorta US doppler|Aorta US doppler
C0801762|T102|relax|35948-9|LNC|Aorta abdominal CT|Aorta abdominal CT
C0801762|T102|relax|35949-7|LNC|Aorta abdominal MRI|Aorta abdominal MRI
C0801762|T102|relax|69276-4|LNC|Aorta abdominal US|Aorta abdominal US
C0801762|T102|relax|37216-9|LNC|Aorta endograft CT|Aorta endograft CT
C0801762|T102|relax|24544-9|LNC|Aorta thoracic CT|Aorta thoracic CT
C0801762|T102|relax|35950-5|LNC|Aorta thoracic MRI|Aorta thoracic MRI
C0801762|T102|relax|24660-3|LNC|Aorta thoracic MRI angiogram|Aorta thoracic MRI angiogram
C0801762|T102|relax|30863-5|LNC|Abdominal Aorta Arteries MRI angiogram|Abdominal Aorta Arteries MRI angiogram
C0801762|T102|relax|35951-3|LNC|Aortic arch MRI angiogram|Aortic arch MRI angiogram
C0801762|T102|relax|30861-9|LNC|Aortic arch Neck vessels MRI angiogram|Aortic arch Neck vessels MRI angiogram
C0801762|T102|relax|35952-1|LNC|Appendix CT|Appendix CT
C0801762|T102|relax|24548-0|LNC|Appendix US|Appendix US
C0801762|T102|relax|39040-1|LNC|AV fistula US|AV fistula US
C0801762|T102|relax|43508-1|LNC|Axilla left MRI|Axilla left MRI
C0801762|T102|relax|72529-1|LNC|Axilla left US|Axilla left US
C0801762|T102|relax|43510-7|LNC|Axilla right MRI|Axilla right MRI
C0801762|T102|relax|72528-3|LNC|Axilla right US|Axilla right US
C0801762|T102|relax|37219-3|LNC|Biliary ducts MRI|Biliary ducts MRI
C0801762|T102|relax|38021-2|LNC|Biliary ducts Gallbladder US|Biliary ducts Gallbladder US
C0801762|T102|relax|37220-1|LNC|Biliary ducts Pancreatic duct MRI|Biliary ducts Pancreatic duct MRI
C0801762|T102|relax|39039-3|LNC|Brachiocephalic artery US doppler|Brachiocephalic artery US doppler
C0801762|T102|relax|24590-2|LNC|Brain MRI|Brain MRI
C0801762|T102|relax|58748-5|LNC|Brain Functional MRI|Brain Functional MRI
C0801762|T102|relax|44138-6|LNC|Brain PET|Brain PET
C0801762|T102|relax|37217-7|LNC|Brain Stem Nerves cranial MRI|Brain Stem Nerves cranial MRI
C0801762|T102|relax|37218-5|LNC|Brain temporal MRI|Brain temporal MRI
C0801762|T102|relax|43772-3|LNC|Brain Internal auditory canal MRI|Brain Internal auditory canal MRI
C0801762|T102|relax|42385-5|LNC|Brain Pituitary Sella turcica MRI|Brain Pituitary Sella turcica MRI
C0801762|T102|relax|30794-2|LNC|Breast MRI|Breast MRI
C0801762|T102|relax|24601-7|LNC|Breast US|Breast US
C0801762|T102|relax|69165-9|LNC|Breast implant bilateral MRI|Breast implant bilateral MRI
C0801762|T102|relax|38057-6|LNC|Breast implant left MRI|Breast implant left MRI
C0801762|T102|relax|38058-4|LNC|Breast implant right MRI|Breast implant right MRI
C0801762|T102|relax|24596-9|LNC|Breast specimen US|Breast specimen US
C0801762|T102|relax|69397-8|LNC|Breast vessels US doppler|Breast vessels US doppler
C0801762|T102|relax|30795-9|LNC|Breast bilateral MRI|Breast bilateral MRI
C0801762|T102|relax|26214-7|LNC|Breast bilateral US|Breast bilateral US
C0801762|T102|relax|35954-7|LNC|Breast left MRI|Breast left MRI
C0801762|T102|relax|26215-4|LNC|Breast left US|Breast left US
C0801762|T102|relax|35955-4|LNC|Breast right MRI|Breast right MRI
C0801762|T102|relax|26216-2|LNC|Breast right US|Breast right US
C0801762|T102|relax|46299-4|LNC|Breast unilateral MRI|Breast unilateral MRI
C0801762|T102|relax|36010-7|LNC|Calcaneus CT|Calcaneus CT
C0801762|T102|relax|36011-5|LNC|Calcaneus X-ray tomograph|Calcaneus X-ray tomograph
C0801762|T102|relax|24616-5|LNC|Carotid artery US|Carotid artery US
C0801762|T102|relax|42146-1|LNC|Carotid artery US doppler|Carotid artery US doppler
C0801762|T102|relax|26217-0|LNC|Carotid artery bilateral US|Carotid artery bilateral US
C0801762|T102|relax|43765-7|LNC|Carotid artery bilateral US doppler|Carotid artery bilateral US doppler
C0801762|T102|relax|26218-8|LNC|Carotid artery left US|Carotid artery left US
C0801762|T102|relax|39427-0|LNC|Carotid artery left US doppler|Carotid artery left US doppler
C0801762|T102|relax|26219-6|LNC|Carotid artery right US|Carotid artery right US
C0801762|T102|relax|39437-9|LNC|Carotid artery right US doppler|Carotid artery right US doppler
C0801762|T102|relax|43552-9|LNC|Carotid artery unilateral US|Carotid artery unilateral US
C0801762|T102|relax|36793-8|LNC|Carotid vessel MRI angiogram|Carotid vessel MRI angiogram
C0801762|T102|relax|30859-3|LNC|Carotid vessels Neck Vessels MRI angiogram|Carotid vessels Neck Vessels MRI angiogram
C0801762|T102|relax|30865-0|LNC|Celiac vessels Superior mesenteric Vessels MRI angiogram|Celiac vessels Superior mesenteric Vessels MRI angiogram
C0801762|T102|relax|46374-5|LNC|Cerebral artery US|Cerebral artery US
C0801762|T102|relax|24627-2|LNC|Chest CT|Chest CT
C0801762|T102|relax|24629-8|LNC|Chest MRI|Chest MRI
C0801762|T102|relax|24630-6|LNC|Chest US|Chest US
C0801762|T102|relax|24657-9|LNC|Chest X-ray tomograph|Chest X-ray tomograph
C0801762|T102|relax|30862-7|LNC|Chest vessels MRI angiogram|Chest vessels MRI angiogram
C0801762|T102|relax|38016-2|LNC|Chest wall US|Chest wall US
C0801762|T102|relax|37235-9|LNC|Circle Willis MRI angiogram|Circle Willis MRI angiogram
C0801762|T102|relax|35960-4|LNC|Clavicle CT|Clavicle CT
C0801762|T102|relax|35961-2|LNC|Clavicle MRI|Clavicle MRI
C0801762|T102|relax|35959-6|LNC|Clavicle X-ray tomograph|Clavicle X-ray tomograph
C0801762|T102|relax|44120-4|LNC|Colon CT|Colon CT
C0801762|T102|relax|24757-7|LNC|Coronary arteries CT fast|Coronary arteries CT fast
C0801762|T102|relax|35962-0|LNC|Elbow CT|Elbow CT
C0801762|T102|relax|24674-4|LNC|Elbow MRI|Elbow MRI
C0801762|T102|relax|35963-8|LNC|Elbow X-ray tomograph|Elbow X-ray tomograph
C0801762|T102|relax|35965-3|LNC|Elbow bilateral CT|Elbow bilateral CT
C0801762|T102|relax|26220-4|LNC|Elbow bilateral MRI|Elbow bilateral MRI
C0801762|T102|relax|35964-6|LNC|Elbow bilateral X-ray tomograph|Elbow bilateral X-ray tomograph
C0801762|T102|relax|35966-1|LNC|Elbow left CT|Elbow left CT
C0801762|T102|relax|26221-2|LNC|Elbow left MRI|Elbow left MRI
C0801762|T102|relax|35967-9|LNC|Elbow left X-ray tomograph|Elbow left X-ray tomograph
C0801762|T102|relax|35968-7|LNC|Elbow right CT|Elbow right CT
C0801762|T102|relax|26222-0|LNC|Elbow right MRI|Elbow right MRI
C0801762|T102|relax|37688-9|LNC|Elbow right X-ray tomograph|Elbow right X-ray tomograph
C0801762|T102|relax|35969-5|LNC|Esophagus CT|Esophagus CT
C0801762|T102|relax|57823-7|LNC|Esophagus PET|Esophagus PET
C0801762|T102|relax|24690-0|LNC|Extremity CT|Extremity CT
C0801762|T102|relax|69193-1|LNC|Extremity MRI|Extremity MRI
C0801762|T102|relax|24693-4|LNC|Extremity US|Extremity US
C0801762|T102|relax|35970-3|LNC|Extremity X-ray tomograph|Extremity X-ray tomograph
C0801762|T102|relax|39042-7|LNC|Extremity artery US doppler|Extremity artery US doppler
C0801762|T102|relax|39031-0|LNC|Extremity artery bilateral US doppler|Extremity artery bilateral US doppler
C0801762|T102|relax|69293-9|LNC|Extremity artery left US|Extremity artery left US
C0801762|T102|relax|39428-8|LNC|Extremity artery left US doppler|Extremity artery left US doppler
C0801762|T102|relax|69297-0|LNC|Extremity artery right US|Extremity artery right US
C0801762|T102|relax|39439-5|LNC|Extremity artery right US doppler|Extremity artery right US doppler
C0801762|T102|relax|39449-4|LNC|Extremity vein US doppler|Extremity vein US doppler
C0801762|T102|relax|39418-9|LNC|Extremity vein bilateral US doppler|Extremity vein bilateral US doppler
C0801762|T102|relax|42145-3|LNC|Extremity vein left US|Extremity vein left US
C0801762|T102|relax|39429-6|LNC|Extremity vein left US doppler|Extremity vein left US doppler
C0801762|T102|relax|42144-6|LNC|Extremity vein right US|Extremity vein right US
C0801762|T102|relax|39440-3|LNC|Extremity vein right US doppler|Extremity vein right US doppler
C0801762|T102|relax|30876-7|LNC|Extremity veins MRI angiogram|Extremity veins MRI angiogram
C0801762|T102|relax|69283-0|LNC|Extremity veins bilateral US doppler|Extremity veins bilateral US doppler
C0801762|T102|relax|41835-0|LNC|Extremity veins left US|Extremity veins left US
C0801762|T102|relax|41816-0|LNC|Extremity veins right US|Extremity veins right US
C0801762|T102|relax|36794-6|LNC|Extremity vessels MRI angiogram|Extremity vessels MRI angiogram
C0801762|T102|relax|43771-5|LNC|Extremity vessels US doppler|Extremity vessels US doppler
C0801762|T102|relax|39495-7|LNC|Extremity vessels bilateral US doppler|Extremity vessels bilateral US doppler
C0801762|T102|relax|69398-6|LNC|Extremity vessels Left US doppler|Extremity vessels Left US doppler
C0801762|T102|relax|39503-8|LNC|Extremity vessels right US doppler|Extremity vessels right US doppler
C0801762|T102|relax|26224-6|LNC|Extremity bilateral CT|Extremity bilateral CT
C0801762|T102|relax|26223-8|LNC|Extremity bilateral US|Extremity bilateral US
C0801762|T102|relax|26226-1|LNC|Extremity left CT|Extremity left CT
C0801762|T102|relax|26225-3|LNC|Extremity left US|Extremity left US
C0801762|T102|relax|26231-1|LNC|Extremity right CT|Extremity right CT
C0801762|T102|relax|26230-3|LNC|Extremity right US|Extremity right US
C0801762|T102|relax|35953-9|LNC|Face MRI|Face MRI
C0801762|T102|relax|41808-7|LNC|Facial bones Maxilla CT|Facial bones Maxilla CT
C0801762|T102|relax|24696-7|LNC|Facial bones Sinuses CT|Facial bones Sinuses CT
C0801762|T102|relax|69389-5|LNC|Femoral artery Popliteal artery US|Femoral artery Popliteal artery US
C0801762|T102|relax|69399-4|LNC|Femoral vein Popliteal vein US|Femoral vein Popliteal vein US
C0801762|T102|relax|30871-8|LNC|Femoral vessels MRI angiogram|Femoral vessels MRI angiogram
C0801762|T102|relax|38134-3|LNC|Femoral vessels US|Femoral vessels US
C0801762|T102|relax|38128-5|LNC|Femoral vessels bilateral US|Femoral vessels bilateral US
C0801762|T102|relax|39498-1|LNC|Femoral vessels left US doppler|Femoral vessels left US doppler
C0801762|T102|relax|39504-6|LNC|Femoral vessels right US doppler|Femoral vessels right US doppler
C0801762|T102|relax|35984-4|LNC|Femur CT|Femur CT
C0801762|T102|relax|35985-1|LNC|Femur X-ray tomograph|Femur X-ray tomograph
C0801762|T102|relax|35986-9|LNC|Femur bilateral X-ray tomograph|Femur bilateral X-ray tomograph
C0801762|T102|relax|35987-7|LNC|Femur left CT|Femur left CT
C0801762|T102|relax|38037-8|LNC|Femur left US|Femur left US
C0801762|T102|relax|35988-5|LNC|Femur left X-ray tomograph|Femur left X-ray tomograph
C0801762|T102|relax|35989-3|LNC|Femur right CT|Femur right CT
C0801762|T102|relax|38048-5|LNC|Femur right US|Femur right US
C0801762|T102|relax|38768-8|LNC|Femur right X-ray tomograph|Femur right X-ray tomograph
C0801762|T102|relax|24705-6|LNC|Finger MRI|Finger MRI
C0801762|T102|relax|26238-6|LNC|Finger bilateral MRI|Finger bilateral MRI
C0801762|T102|relax|26239-4|LNC|Finger left MRI|Finger left MRI
C0801762|T102|relax|26240-2|LNC|Finger right MRI|Finger right MRI
C0801762|T102|relax|37221-9|LNC|Fistula CT|Fistula CT
C0801762|T102|relax|35991-9|LNC|Foot CT|Foot CT
C0801762|T102|relax|24707-2|LNC|Foot MRI|Foot MRI
C0801762|T102|relax|35992-7|LNC|Foot X-ray tomograph|Foot X-ray tomograph
C0801762|T102|relax|30872-6|LNC|Foot vessels MRI angiogram|Foot vessels MRI angiogram
C0801762|T102|relax|46362-0|LNC|Foot vessels US doppler|Foot vessels US doppler
C0801762|T102|relax|35993-5|LNC|Foot bilateral CT|Foot bilateral CT
C0801762|T102|relax|26241-0|LNC|Foot bilateral MRI|Foot bilateral MRI
C0801762|T102|relax|35994-3|LNC|Foot left CT|Foot left CT
C0801762|T102|relax|26242-8|LNC|Foot left MRI|Foot left MRI
C0801762|T102|relax|35995-0|LNC|Foot left X-ray tomograph|Foot left X-ray tomograph
C0801762|T102|relax|35996-8|LNC|Foot right CT|Foot right CT
C0801762|T102|relax|26243-6|LNC|Foot right MRI|Foot right MRI
C0801762|T102|relax|37706-9|LNC|Foot right X-ray tomograph|Foot right X-ray tomograph
C0801762|T102|relax|35997-6|LNC|Forearm CT|Forearm CT
C0801762|T102|relax|24710-6|LNC|Forearm MRI|Forearm MRI
C0801762|T102|relax|30873-4|LNC|Forearm vessels MRI angiogram|Forearm vessels MRI angiogram
C0801762|T102|relax|35998-4|LNC|Forearm bilateral CT|Forearm bilateral CT
C0801762|T102|relax|26244-4|LNC|Forearm bilateral MRI|Forearm bilateral MRI
C0801762|T102|relax|35999-2|LNC|Forearm left CT|Forearm left CT
C0801762|T102|relax|26245-1|LNC|Forearm left MRI|Forearm left MRI
C0801762|T102|relax|36000-8|LNC|Forearm right CT|Forearm right CT
C0801762|T102|relax|26246-9|LNC|Forearm right MRI|Forearm right MRI
C0801762|T102|relax|24711-4|LNC|Gallbladder US|Gallbladder US
C0801762|T102|relax|36001-6|LNC|Gallbladder X-ray tomograph|Gallbladder X-ray tomograph
C0801762|T102|relax|39415-5|LNC|Gastrointestine US|Gastrointestine US
C0801762|T102|relax|39416-3|LNC|Genitourinary system US|Genitourinary system US
C0801762|T102|relax|37236-7|LNC|Great vessel MRI|Great vessel MRI
C0801762|T102|relax|24719-7|LNC|Groin US|Groin US
C0801762|T102|relax|36002-4|LNC|Hand CT|Hand CT
C0801762|T102|relax|24720-5|LNC|Hand MRI|Hand MRI
C0801762|T102|relax|36003-2|LNC|Hand X-ray tomograph|Hand X-ray tomograph
C0801762|T102|relax|46382-8|LNC|Hand vessels US doppler|Hand vessels US doppler
C0801762|T102|relax|36004-0|LNC|Hand bilateral CT|Hand bilateral CT
C0801762|T102|relax|26247-7|LNC|Hand bilateral MRI|Hand bilateral MRI
C0801762|T102|relax|36005-7|LNC|Hand left CT|Hand left CT
C0801762|T102|relax|26248-5|LNC|Hand left MRI|Hand left MRI
C0801762|T102|relax|36006-5|LNC|Hand left X-ray tomograph|Hand left X-ray tomograph
C0801762|T102|relax|36007-3|LNC|Hand right CT|Hand right CT
C0801762|T102|relax|26249-3|LNC|Hand right MRI|Hand right MRI
C0801762|T102|relax|37717-6|LNC|Hand right X-ray tomograph|Hand right X-ray tomograph
C0801762|T102|relax|24725-4|LNC|Head CT|Head CT
C0801762|T102|relax|24728-8|LNC|Head CT cine|Head CT cine
C0801762|T102|relax|24731-2|LNC|Head US|Head US
C0801762|T102|relax|58741-0|LNC|Head to thigh PET|Head to thigh PET
C0801762|T102|relax|30858-5|LNC|Head veins MRI angiogram|Head veins MRI angiogram
C0801762|T102|relax|30856-9|LNC|Head vessels MRI angiogram|Head vessels MRI angiogram
C0801762|T102|relax|24733-8|LNC|Head vessels US doppler|Head vessels US doppler
C0801762|T102|relax|42304-6|LNC|Head vessels Neck vessels MRI angiogram|Head vessels Neck vessels MRI angiogram
C0801762|T102|relax|30880-9|LNC|Head vessels Neck vessels US doppler|Head vessels Neck vessels US doppler
C0801762|T102|relax|30655-5|LNC|Head Cistern MRI|Head Cistern MRI
C0801762|T102|relax|24746-0|LNC|Head Sagittal Sinus MRI|Head Sagittal Sinus MRI
C0801762|T102|relax|58742-8|LNC|Head Neck PET|Head Neck PET
C0801762|T102|relax|44164-2|LNC|Head Neck US|Head Neck US
C0801762|T102|relax|58744-4|LNC|Heart CT|Heart CT
C0801762|T102|relax|24748-6|LNC|Heart MRI|Heart MRI
C0801762|T102|relax|36009-9|LNC|Heart MRI angiogram|Heart MRI angiogram
C0801762|T102|relax|44137-8|LNC|Heart PET|Heart PET
C0801762|T102|relax|42148-7|LNC|Heart US|Heart US
C0801762|T102|relax|36014-9|LNC|Hip CT|Hip CT
C0801762|T102|relax|36013-1|LNC|Hip MRI|Hip MRI
C0801762|T102|relax|24760-1|LNC|Hip US|Hip US
C0801762|T102|relax|36012-3|LNC|Hip X-ray tomograph|Hip X-ray tomograph
C0801762|T102|relax|36016-4|LNC|Hip bilateral CT|Hip bilateral CT
C0801762|T102|relax|36017-2|LNC|Hip bilateral MRI|Hip bilateral MRI
C0801762|T102|relax|26250-1|LNC|Hip bilateral US|Hip bilateral US
C0801762|T102|relax|36015-6|LNC|Hip bilateral X-ray tomograph|Hip bilateral X-ray tomograph
C0801762|T102|relax|36018-0|LNC|Hip left CT|Hip left CT
C0801762|T102|relax|36020-6|LNC|Hip left MRI|Hip left MRI
C0801762|T102|relax|26251-9|LNC|Hip left US|Hip left US
C0801762|T102|relax|36019-8|LNC|Hip left X-ray tomograph|Hip left X-ray tomograph
C0801762|T102|relax|36021-4|LNC|Hip right CT|Hip right CT
C0801762|T102|relax|36022-2|LNC|Hip right MRI|Hip right MRI
C0801762|T102|relax|26252-7|LNC|Hip right US|Hip right US
C0801762|T102|relax|37735-8|LNC|Hip right X-ray tomograph|Hip right X-ray tomograph
C0801762|T102|relax|43566-9|LNC|Hip Thigh US|Hip Thigh US
C0801762|T102|relax|36024-8|LNC|Humerus X-ray tomograph|Humerus X-ray tomograph
C0801762|T102|relax|39425-4|LNC|Iliac artery US doppler|Iliac artery US doppler
C0801762|T102|relax|42147-9|LNC|Iliac graft US doppler|Iliac graft US doppler
C0801762|T102|relax|39497-3|LNC|Iliac vessels US doppler|Iliac vessels US doppler
C0801762|T102|relax|38129-3|LNC|Iliac vessels bilateral US|Iliac vessels bilateral US
C0801762|T102|relax|38137-6|LNC|Iliac vessels left US|Iliac vessels left US
C0801762|T102|relax|38141-8|LNC|Iliac vessels right US|Iliac vessels right US
C0801762|T102|relax|35958-8|LNC|Internal auditory canal CT|Internal auditory canal CT
C0801762|T102|relax|35956-2|LNC|Internal auditory canal MRI|Internal auditory canal MRI
C0801762|T102|relax|24767-6|LNC|Internal auditory canal X-ray tomograph|Internal auditory canal X-ray tomograph
C0801762|T102|relax|26253-5|LNC|Internal auditory canal bilateral X-ray tomograph|Internal auditory canal bilateral X-ray tomograph
C0801762|T102|relax|35957-0|LNC|Internal auditory canal left CT|Internal auditory canal left CT
C0801762|T102|relax|26254-3|LNC|Internal auditory canal left X-ray tomograph|Internal auditory canal left X-ray tomograph
C0801762|T102|relax|38767-0|LNC|Internal auditory canal right CT|Internal auditory canal right CT
C0801762|T102|relax|26255-0|LNC|Internal auditory canal right X-ray tomograph|Internal auditory canal right X-ray tomograph
C0801762|T102|relax|24735-3|LNC|Internal auditory canal Posterior fossa MRI|Internal auditory canal Posterior fossa MRI
C0801762|T102|relax|36033-9|LNC|Kidney MRI|Kidney MRI
C0801762|T102|relax|38036-0|LNC|Kidney US|Kidney US
C0801762|T102|relax|36032-1|LNC|Kidney X-ray tomograph|Kidney X-ray tomograph
C0801762|T102|relax|39032-8|LNC|Kidney transplant US|Kidney transplant US
C0801762|T102|relax|42477-0|LNC|Kidney vessels transplant US doppler|Kidney vessels transplant US doppler
C0801762|T102|relax|43767-3|LNC|Kidney bilateral CT|Kidney bilateral CT
C0801762|T102|relax|36034-7|LNC|Kidney bilateral MRI|Kidney bilateral MRI
C0801762|T102|relax|43774-9|LNC|Kidney bilateral US|Kidney bilateral US
C0801762|T102|relax|24789-0|LNC|Kidney bilateral X-ray tomograph|Kidney bilateral X-ray tomograph
C0801762|T102|relax|69402-6|LNC|Kidney Bilateral Bladder US|Kidney Bilateral Bladder US
C0801762|T102|relax|36035-4|LNC|Kidney left MRI|Kidney left MRI
C0801762|T102|relax|38038-6|LNC|Kidney left US|Kidney left US
C0801762|T102|relax|69113-9|LNC|Kidney right CT|Kidney right CT
C0801762|T102|relax|36036-2|LNC|Kidney right MRI|Kidney right MRI
C0801762|T102|relax|38049-3|LNC|Kidney right US|Kidney right US
C0801762|T102|relax|36037-0|LNC|Knee CT|Knee CT
C0801762|T102|relax|24802-1|LNC|Knee MRI|Knee MRI
C0801762|T102|relax|36038-8|LNC|Knee X-ray tomograph|Knee X-ray tomograph
C0801762|T102|relax|36799-5|LNC|Knee vessels MRI angiogram|Knee vessels MRI angiogram
C0801762|T102|relax|36800-1|LNC|Knee vessels left MRI angiogram|Knee vessels left MRI angiogram
C0801762|T102|relax|36801-9|LNC|Knee vessels right MRI angiogram|Knee vessels right MRI angiogram
C0801762|T102|relax|36040-4|LNC|Knee bilateral CT|Knee bilateral CT
C0801762|T102|relax|26256-8|LNC|Knee bilateral MRI|Knee bilateral MRI
C0801762|T102|relax|36039-6|LNC|Knee bilateral X-ray tomograph|Knee bilateral X-ray tomograph
C0801762|T102|relax|36041-2|LNC|Knee left CT|Knee left CT
C0801762|T102|relax|26257-6|LNC|Knee left MRI|Knee left MRI
C0801762|T102|relax|36042-0|LNC|Knee left X-ray tomograph|Knee left X-ray tomograph
C0801762|T102|relax|36043-8|LNC|Knee right CT|Knee right CT
C0801762|T102|relax|26258-4|LNC|Knee right MRI|Knee right MRI
C0801762|T102|relax|37760-6|LNC|Knee right X-ray tomograph|Knee right X-ray tomograph
C0801762|T102|relax|36045-3|LNC|Larynx MRI|Larynx MRI
C0801762|T102|relax|36044-6|LNC|Larynx X-ray tomograph|Larynx X-ray tomograph
C0801762|T102|relax|24814-6|LNC|Liver CT|Liver CT
C0801762|T102|relax|36046-1|LNC|Liver MRI|Liver MRI
C0801762|T102|relax|28614-6|LNC|Liver US|Liver US
C0801762|T102|relax|39454-4|LNC|Liver transplant US|Liver transplant US
C0801762|T102|relax|24818-7|LNC|Liver Diaphragm US|Liver Diaphragm US
C0801762|T102|relax|35971-1|LNC|Lower extremity CT|Lower extremity CT
C0801762|T102|relax|30692-8|LNC|Lower extremity MRI|Lower extremity MRI
C0801762|T102|relax|30709-0|LNC|Lower extremity US|Lower extremity US
C0801762|T102|relax|35972-9|LNC|Lower extremity X-ray tomograph|Lower extremity X-ray tomograph
C0801762|T102|relax|48693-6|LNC|Lower extremity artery US|Lower extremity artery US
C0801762|T102|relax|39434-6|LNC|Lower extremity artery US doppler|Lower extremity artery US doppler
C0801762|T102|relax|38130-1|LNC|Lower extremity artery bilateral US|Lower extremity artery bilateral US
C0801762|T102|relax|39421-3|LNC|Lower extremity artery bilateral US doppler|Lower extremity artery bilateral US doppler
C0801762|T102|relax|41834-3|LNC|Lower extremity artery left US|Lower extremity artery left US
C0801762|T102|relax|39499-9|LNC|Lower extremity artery left US doppler|Lower extremity artery left US doppler
C0801762|T102|relax|41815-2|LNC|Lower extremity artery right US|Lower extremity artery right US
C0801762|T102|relax|39505-3|LNC|Lower extremity artery right US doppler|Lower extremity artery right US doppler
C0801762|T102|relax|46363-8|LNC|Lower extremity vein US|Lower extremity vein US
C0801762|T102|relax|30881-7|LNC|Lower extremity vein US doppler|Lower extremity vein US doppler
C0801762|T102|relax|46364-6|LNC|Lower extremity vein bilateral US|Lower extremity vein bilateral US
C0801762|T102|relax|39420-5|LNC|Lower extremity vein bilateral US doppler|Lower extremity vein bilateral US doppler
C0801762|T102|relax|48692-8|LNC|Lower extremity vein left US|Lower extremity vein left US
C0801762|T102|relax|39432-0|LNC|Lower extremity vein left US doppler|Lower extremity vein left US doppler
C0801762|T102|relax|48691-0|LNC|Lower extremity vein right US|Lower extremity vein right US
C0801762|T102|relax|39443-7|LNC|Lower extremity vein right US doppler|Lower extremity vein right US doppler
C0801762|T102|relax|36079-2|LNC|Lower extremity veins MRI angiogram|Lower extremity veins MRI angiogram
C0801762|T102|relax|69385-3|LNC|Lower extremity veins bilateral US|Lower extremity veins bilateral US
C0801762|T102|relax|36784-7|LNC|Lower extremity veins left MRI angiogram|Lower extremity veins left MRI angiogram
C0801762|T102|relax|69392-9|LNC|Lower extremity veins left US|Lower extremity veins left US
C0801762|T102|relax|36785-4|LNC|Lower extremity veins right MRI angiogram|Lower extremity veins right MRI angiogram
C0801762|T102|relax|42461-4|LNC|Lower extremity vessel graft left US doppler|Lower extremity vessel graft left US doppler
C0801762|T102|relax|42462-2|LNC|Lower extremity vessel graft right US doppler|Lower extremity vessel graft right US doppler
C0801762|T102|relax|30874-2|LNC|Lower extremity vessels MRI angiogram|Lower extremity vessels MRI angiogram
C0801762|T102|relax|44174-1|LNC|Lower extremity vessels US doppler|Lower extremity vessels US doppler
C0801762|T102|relax|35974-5|LNC|Lower extremity vessels bilateral MRI angiogram|Lower extremity vessels bilateral MRI angiogram
C0801762|T102|relax|39422-1|LNC|Lower extremity vessels bilateral US doppler|Lower extremity vessels bilateral US doppler
C0801762|T102|relax|36795-3|LNC|Lower extremity vessels left MRI angiogram|Lower extremity vessels left MRI angiogram
C0801762|T102|relax|39431-2|LNC|Lower extremity vessels left US doppler|Lower extremity vessels left US doppler
C0801762|T102|relax|36796-1|LNC|Lower extremity vessels right MRI angiogram|Lower extremity vessels right MRI angiogram
C0801762|T102|relax|39442-9|LNC|Lower extremity vessels right US doppler|Lower extremity vessels right US doppler
C0801762|T102|relax|35973-7|LNC|Lower extremity bilateral CT|Lower extremity bilateral CT
C0801762|T102|relax|35975-2|LNC|Lower extremity bilateral MRI|Lower extremity bilateral MRI
C0801762|T102|relax|38013-9|LNC|Lower extremity bilateral US|Lower extremity bilateral US
C0801762|T102|relax|24687-6|LNC|Lower Extremity Joint MRI|Lower Extremity Joint MRI
C0801762|T102|relax|26227-9|LNC|Lower extremity joint bilateral MRI|Lower extremity joint bilateral MRI
C0801762|T102|relax|26228-7|LNC|Lower extremity joint left MRI|Lower extremity joint left MRI
C0801762|T102|relax|26229-5|LNC|Lower extremity joint right MRI|Lower extremity joint right MRI
C0801762|T102|relax|35976-0|LNC|Lower extremity left CT|Lower extremity left CT
C0801762|T102|relax|35978-6|LNC|Lower extremity left MRI|Lower extremity left MRI
C0801762|T102|relax|38040-2|LNC|Lower extremity left US|Lower extremity left US
C0801762|T102|relax|35977-8|LNC|Lower extremity left X-ray tomograph|Lower extremity left X-ray tomograph
C0801762|T102|relax|35979-4|LNC|Lower extremity right CT|Lower extremity right CT
C0801762|T102|relax|35980-2|LNC|Lower extremity right MRI|Lower extremity right MRI
C0801762|T102|relax|38051-9|LNC|Lower extremity right US|Lower extremity right US
C0801762|T102|relax|37766-3|LNC|Lower extremity right X-ray tomograph|Lower extremity right X-ray tomograph
C0801762|T102|relax|36074-3|LNC|Lower leg CT|Lower leg CT
C0801762|T102|relax|24821-1|LNC|Lower leg MRI|Lower leg MRI
C0801762|T102|relax|43513-1|LNC|Lower leg vessels left MRI angiogram|Lower leg vessels left MRI angiogram
C0801762|T102|relax|43556-0|LNC|Lower leg vessels right MRI angiogram|Lower leg vessels right MRI angiogram
C0801762|T102|relax|42696-5|LNC|Lower leg bilateral MRI|Lower leg bilateral MRI
C0801762|T102|relax|36075-0|LNC|Lower leg left MRI|Lower leg left MRI
C0801762|T102|relax|36076-8|LNC|Lower leg right MRI|Lower leg right MRI
C0801762|T102|relax|30866-8|LNC|Lumbar plexus MRI|Lumbar plexus MRI
C0801762|T102|relax|57822-9|LNC|Lung PET|Lung PET
C0801762|T102|relax|36047-9|LNC|Mandible CT|Mandible CT
C0801762|T102|relax|36048-7|LNC|Mandible X-ray tomograph|Mandible X-ray tomograph
C0801762|T102|relax|38043-6|LNC|Mastoid US|Mastoid US
C0801762|T102|relax|36776-3|LNC|Mastoid X-ray tomograph|Mastoid X-ray tomograph
C0801762|T102|relax|46298-6|LNC|Mastoid bilateral CT|Mastoid bilateral CT
C0801762|T102|relax|36050-3|LNC|Maxilla CT|Maxilla CT
C0801762|T102|relax|36049-5|LNC|Maxilla Mandible CT|Maxilla Mandible CT
C0801762|T102|relax|37234-2|LNC|Mediastinum MRI|Mediastinum MRI
C0801762|T102|relax|38044-4|LNC|Mediastinum US|Mediastinum US
C0801762|T102|relax|37233-4|LNC|Mediastinum X-ray tomograph|Mediastinum X-ray tomograph
C0801762|T102|relax|69394-5|LNC|Mesenteric artery US|Mesenteric artery US
C0801762|T102|relax|69211-1|LNC|Nasal bones MRI|Nasal bones MRI
C0801762|T102|relax|37606-1|LNC|Nasal bones X-ray tomograph|Nasal bones X-ray tomograph
C0801762|T102|relax|30860-1|LNC|Nasopharynx MRI|Nasopharynx MRI
C0801762|T102|relax|24835-1|LNC|Nasopharynx Neck CT|Nasopharynx Neck CT
C0801762|T102|relax|36051-1|LNC|Neck CT|Neck CT
C0801762|T102|relax|24839-3|LNC|Neck MRI|Neck MRI
C0801762|T102|relax|24842-7|LNC|Neck US|Neck US
C0801762|T102|relax|36788-8|LNC|Neck veins MRI angiogram|Neck veins MRI angiogram
C0801762|T102|relax|36085-9|LNC|Neck vessels MRI angiogram|Neck vessels MRI angiogram
C0801762|T102|relax|44175-8|LNC|Neck vessels US doppler|Neck vessels US doppler
C0801762|T102|relax|30857-7|LNC|Nerves cranial MRI|Nerves cranial MRI
C0801762|T102|relax|41807-9|LNC|Orbit CT|Orbit CT
C0801762|T102|relax|36777-1|LNC|Orbit MRI|Orbit MRI
C0801762|T102|relax|36802-7|LNC|Orbit vessels MRI angiogram|Orbit vessels MRI angiogram
C0801762|T102|relax|24848-4|LNC|Orbit bilateral CT|Orbit bilateral CT
C0801762|T102|relax|37611-1|LNC|Orbit bilateral X-ray tomograph|Orbit bilateral X-ray tomograph
C0801762|T102|relax|38836-3|LNC|Orbit left MRI|Orbit left MRI
C0801762|T102|relax|36778-9|LNC|Orbit right MRI|Orbit right MRI
C0801762|T102|relax|42303-8|LNC|Orbit Face MRI|Orbit Face MRI
C0801762|T102|relax|43530-5|LNC|Orbit Face Neck MRI|Orbit Face Neck MRI
C0801762|T102|relax|43455-5|LNC|Oropharynx MRI|Oropharynx MRI
C0801762|T102|relax|39502-0|LNC|Ovarian vessels US doppler|Ovarian vessels US doppler
C0801762|T102|relax|36779-7|LNC|Ovary MRI|Ovary MRI
C0801762|T102|relax|69390-3|LNC|Ovary US|Ovary US
C0801762|T102|relax|43506-5|LNC|Ovary bilateral MRI|Ovary bilateral MRI
C0801762|T102|relax|24857-5|LNC|Pancreas CT|Pancreas CT
C0801762|T102|relax|36052-9|LNC|Pancreas MRI|Pancreas MRI
C0801762|T102|relax|24859-1|LNC|Pancreas US|Pancreas US
C0801762|T102|relax|39509-5|LNC|Pancreas transplant US|Pancreas transplant US
C0801762|T102|relax|36053-7|LNC|Parathyroid MRI|Parathyroid MRI
C0801762|T102|relax|38045-1|LNC|Parathyroid US|Parathyroid US
C0801762|T102|relax|37223-5|LNC|Parotid gland CT|Parotid gland CT
C0801762|T102|relax|37224-3|LNC|Parotid gland MRI|Parotid gland MRI
C0801762|T102|relax|38138-4|LNC|Parotid gland US|Parotid gland US
C0801762|T102|relax|24865-8|LNC|Pelvis CT|Pelvis CT
C0801762|T102|relax|24867-4|LNC|Pelvis MRI|Pelvis MRI
C0801762|T102|relax|24869-0|LNC|Pelvis US|Pelvis US
C0801762|T102|relax|37632-7|LNC|Pelvis X-ray tomograph|Pelvis X-ray tomograph
C0801762|T102|relax|36789-6|LNC|Pelvis veins MRI angiogram|Pelvis veins MRI angiogram
C0801762|T102|relax|30867-6|LNC|Pelvis vessels MRI angiogram|Pelvis vessels MRI angiogram
C0801762|T102|relax|24870-8|LNC|Pelvis vessels US doppler|Pelvis vessels US doppler
C0801762|T102|relax|24872-4|LNC|Pelvis Hip MRI|Pelvis Hip MRI
C0801762|T102|relax|26259-2|LNC|Pelvis Hip bilateral MRI|Pelvis Hip bilateral MRI
C0801762|T102|relax|26260-0|LNC|Pelvis Hip left MRI|Pelvis Hip left MRI
C0801762|T102|relax|26261-8|LNC|Pelvis Hip right MRI|Pelvis Hip right MRI
C0801762|T102|relax|38140-0|LNC|Penis US|Penis US
C0801762|T102|relax|38139-2|LNC|Penis vessels US|Penis vessels US
C0801762|T102|relax|24877-3|LNC|Petrous bone CT|Petrous bone CT
C0801762|T102|relax|36932-2|LNC|Pituitary Sella turcica CT|Pituitary Sella turcica CT
C0801762|T102|relax|24880-7|LNC|Pituitary Sella turcica MRI|Pituitary Sella turcica MRI
C0801762|T102|relax|24881-5|LNC|Popliteal space US|Popliteal space US
C0801762|T102|relax|26262-6|LNC|Popliteal space bilateral US|Popliteal space bilateral US
C0801762|T102|relax|26263-4|LNC|Popliteal space left US|Popliteal space left US
C0801762|T102|relax|26264-2|LNC|Popliteal space right US|Popliteal space right US
C0801762|T102|relax|36077-6|LNC|Portal vein MRI angiogram|Portal vein MRI angiogram
C0801762|T102|relax|69284-8|LNC|Portal vein Hepatic vein US doppler|Portal vein Hepatic vein US doppler
C0801762|T102|relax|36055-2|LNC|Posterior fossa CT|Posterior fossa CT
C0801762|T102|relax|36056-0|LNC|Posterior fossa MRI|Posterior fossa MRI
C0801762|T102|relax|36057-8|LNC|Prostate CT|Prostate CT
C0801762|T102|relax|30675-3|LNC|Prostate MRI|Prostate MRI
C0801762|T102|relax|24884-9|LNC|Prostate US|Prostate US
C0801762|T102|relax|43445-6|LNC|Pulmonary system CT|Pulmonary system CT
C0801762|T102|relax|43454-8|LNC|Pulmonary system MRI|Pulmonary system MRI
C0801762|T102|relax|36803-5|LNC|Pulmonary vessels MRI angiogram|Pulmonary vessels MRI angiogram
C0801762|T102|relax|24892-2|LNC|Rectum US|Rectum US
C0801762|T102|relax|69294-7|LNC|Renal artery US|Renal artery US
C0801762|T102|relax|39435-3|LNC|Renal artery US doppler|Renal artery US doppler
C0801762|T102|relax|36078-4|LNC|Renal vein MRI angiogram|Renal vein MRI angiogram
C0801762|T102|relax|30868-4|LNC|Renal vessels MRI angiogram|Renal vessels MRI angiogram
C0801762|T102|relax|69295-4|LNC|Renal vessels US|Renal vessels US
C0801762|T102|relax|39426-2|LNC|Renal vessels US doppler|Renal vessels US doppler
C0801762|T102|relax|36804-3|LNC|Renal vessels bilateral MRI angiogram|Renal vessels bilateral MRI angiogram
C0801762|T102|relax|39419-7|LNC|Renal vessels bilateral US doppler|Renal vessels bilateral US doppler
C0801762|T102|relax|30619-1|LNC|Sacroiliac Joint CT|Sacroiliac Joint CT
C0801762|T102|relax|36031-3|LNC|Sacroiliac Joint MRI|Sacroiliac Joint MRI
C0801762|T102|relax|36058-6|LNC|Sacrum CT|Sacrum CT
C0801762|T102|relax|36059-4|LNC|Sacrum MRI|Sacrum MRI
C0801762|T102|relax|38053-5|LNC|Sacrum US|Sacrum US
C0801762|T102|relax|37653-3|LNC|Sacrum X-ray tomograph|Sacrum X-ray tomograph
C0801762|T102|relax|69116-2|LNC|Sacrum Coccyx CT|Sacrum Coccyx CT
C0801762|T102|relax|36060-2|LNC|Sacrum Coccyx MRI|Sacrum Coccyx MRI
C0801762|T102|relax|36933-0|LNC|Salivary gland MRI|Salivary gland MRI
C0801762|T102|relax|69298-8|LNC|Salivary gland US|Salivary gland US
C0801762|T102|relax|69117-0|LNC|Scapula CT|Scapula CT
C0801762|T102|relax|36061-0|LNC|Scapula MRI|Scapula MRI
C0801762|T102|relax|36073-5|LNC|Scrotum Testicle MRI|Scrotum Testicle MRI
C0801762|T102|relax|25002-7|LNC|Scrotum Testicle US|Scrotum Testicle US
C0801762|T102|relax|48742-1|LNC|Scrotum Testicle US doppler|Scrotum Testicle US doppler
C0801762|T102|relax|26271-7|LNC|Scrotum Testicle bilateral US|Scrotum Testicle bilateral US
C0801762|T102|relax|26272-5|LNC|Scrotum Testicle left US|Scrotum Testicle left US
C0801762|T102|relax|26273-3|LNC|Scrotum Testicle right US|Scrotum Testicle right US
C0801762|T102|relax|42437-4|LNC|Sella turcica X-ray tomograph|Sella turcica X-ray tomograph
C0801762|T102|relax|36062-8|LNC|Shoulder CT|Shoulder CT
C0801762|T102|relax|24905-2|LNC|Shoulder MRI|Shoulder MRI
C0801762|T102|relax|24907-8|LNC|Shoulder US|Shoulder US
C0801762|T102|relax|37850-5|LNC|Shoulder X-ray tomograph|Shoulder X-ray tomograph
C0801762|T102|relax|36805-0|LNC|Shoulder vessels MRI angiogram|Shoulder vessels MRI angiogram
C0801762|T102|relax|36806-8|LNC|Shoulder vessels left MRI angiogram|Shoulder vessels left MRI angiogram
C0801762|T102|relax|36807-6|LNC|Shoulder vessels right MRI angiogram|Shoulder vessels right MRI angiogram
C0801762|T102|relax|36063-6|LNC|Shoulder bilateral CT|Shoulder bilateral CT
C0801762|T102|relax|26266-7|LNC|Shoulder bilateral MRI|Shoulder bilateral MRI
C0801762|T102|relax|26265-9|LNC|Shoulder bilateral US|Shoulder bilateral US
C0801762|T102|relax|36064-4|LNC|Shoulder left CT|Shoulder left CT
C0801762|T102|relax|26268-3|LNC|Shoulder left MRI|Shoulder left MRI
C0801762|T102|relax|26267-5|LNC|Shoulder left US|Shoulder left US
C0801762|T102|relax|36065-1|LNC|Shoulder left X-ray tomograph|Shoulder left X-ray tomograph
C0801762|T102|relax|36066-9|LNC|Shoulder right CT|Shoulder right CT
C0801762|T102|relax|26270-9|LNC|Shoulder right MRI|Shoulder right MRI
C0801762|T102|relax|26269-1|LNC|Shoulder right US|Shoulder right US
C0801762|T102|relax|37811-7|LNC|Shoulder right X-ray tomograph|Shoulder right X-ray tomograph
C0801762|T102|relax|30588-8|LNC|Sinuses CT|Sinuses CT
C0801762|T102|relax|24914-4|LNC|Sinuses MRI|Sinuses MRI
C0801762|T102|relax|37866-1|LNC|Sinuses X-ray tomograph|Sinuses X-ray tomograph
C0801762|T102|relax|37874-5|LNC|Skull X-ray tomograph|Skull X-ray tomograph
C0801762|T102|relax|37495-9|LNC|Skull base CT|Skull base CT
C0801762|T102|relax|37497-5|LNC|Spine vessels MRI angiogram|Spine vessels MRI angiogram
C0801762|T102|relax|24932-6|LNC|Spine Cervical CT|Spine Cervical CT
C0801762|T102|relax|24935-9|LNC|Spine Cervical MRI|Spine Cervical MRI
C0801762|T102|relax|70926-1|LNC|Spine Cervical US|Spine Cervical US
C0801762|T102|relax|36068-5|LNC|Spine Cervical X-ray tomograph|Spine Cervical X-ray tomograph
C0801762|T102|relax|43457-1|LNC|Spine Cervical Spine Thoracic MRI|Spine Cervical Spine Thoracic MRI
C0801762|T102|relax|42698-1|LNC|Spine Cervical Thoracic Lumbar MRI|Spine Cervical Thoracic Lumbar MRI
C0801762|T102|relax|24963-1|LNC|Spine Lumbar CT|Spine Lumbar CT
C0801762|T102|relax|24968-0|LNC|Spine Lumbar MRI|Spine Lumbar MRI
C0801762|T102|relax|69393-7|LNC|Spine Lumbar US|Spine Lumbar US
C0801762|T102|relax|36069-3|LNC|Spine Lumbar X-ray tomograph|Spine Lumbar X-ray tomograph
C0801762|T102|relax|37232-6|LNC|Spine Lumbosacral Junction CT|Spine Lumbosacral Junction CT
C0801762|T102|relax|24978-9|LNC|Spine Thoracic CT|Spine Thoracic CT
C0801762|T102|relax|24980-5|LNC|Spine Thoracic MRI|Spine Thoracic MRI
C0801762|T102|relax|70927-9|LNC|Spine Thoracic US|Spine Thoracic US
C0801762|T102|relax|37911-5|LNC|Spine Thoracic X-ray tomograph|Spine Thoracic X-ray tomograph
C0801762|T102|relax|49565-5|LNC|Thoracic Spine vessels MRI angiogram|Thoracic Spine vessels MRI angiogram
C0801762|T102|relax|24988-8|LNC|Spleen CT|Spleen CT
C0801762|T102|relax|36070-1|LNC|Spleen MRI|Spleen MRI
C0801762|T102|relax|24990-4|LNC|Spleen US|Spleen US
C0801762|T102|relax|37225-0|LNC|Sternoclavicular Joint CT|Sternoclavicular Joint CT
C0801762|T102|relax|36071-9|LNC|Sternum CT|Sternum CT
C0801762|T102|relax|36072-7|LNC|Sternum MRI|Sternum MRI
C0801762|T102|relax|37885-1|LNC|Sternum X-ray tomograph|Sternum X-ray tomograph
C0801762|T102|relax|36782-1|LNC|Subclavian artery MRI angiogram|Subclavian artery MRI angiogram
C0801762|T102|relax|38131-9|LNC|Subclavian vessels bilateral US|Subclavian vessels bilateral US
C0801762|T102|relax|46359-6|LNC|Superior mesenteric vessels MRI angiogram|Superior mesenteric vessels MRI angiogram
C0801762|T102|relax|44235-0|LNC|Superior mesenteric vessels US doppler|Superior mesenteric vessels US doppler
C0801762|T102|relax|42468-9|LNC|Surgical specimen US|Surgical specimen US
C0801762|T102|relax|38059-2|LNC|Talus CT|Talus CT
C0801762|T102|relax|36773-0|LNC|Temporal bone CT|Temporal bone CT
C0801762|T102|relax|37226-8|LNC|Temporomandibular joint CT|Temporomandibular joint CT
C0801762|T102|relax|24999-5|LNC|Temporomandibular joint MRI|Temporomandibular joint MRI
C0801762|T102|relax|30719-9|LNC|Temporomandibular joint X-ray tomograph|Temporomandibular joint X-ray tomograph
C0801762|T102|relax|37228-4|LNC|Temporomandibular joint bilateral MRI|Temporomandibular joint bilateral MRI
C0801762|T102|relax|37227-6|LNC|Temporomandibular joint bilateral X-ray tomograph|Temporomandibular joint bilateral X-ray tomograph
C0801762|T102|relax|37230-0|LNC|Temporomandibular joint left MRI|Temporomandibular joint left MRI
C0801762|T102|relax|37229-2|LNC|Temporomandibular joint left X-ray tomograph|Temporomandibular joint left X-ray tomograph
C0801762|T102|relax|37231-8|LNC|Temporomandibular joint right MRI|Temporomandibular joint right MRI
C0801762|T102|relax|37819-0|LNC|Temporomandibular joint right X-ray tomograph|Temporomandibular joint right X-ray tomograph
C0801762|T102|relax|39446-0|LNC|Testicle vessels US doppler|Testicle vessels US doppler
C0801762|T102|relax|24702-3|LNC|Thigh MRI|Thigh MRI
C0801762|T102|relax|26235-2|LNC|Thigh bilateral MRI|Thigh bilateral MRI
C0801762|T102|relax|26236-0|LNC|Thigh left MRI|Thigh left MRI
C0801762|T102|relax|26237-8|LNC|Thigh right MRI|Thigh right MRI
C0801762|T102|relax|36054-5|LNC|Thoracic outlet CT|Thoracic outlet CT
C0801762|T102|relax|24582-9|LNC|Thoracic outlet MRI|Thoracic outlet MRI
C0801762|T102|relax|44163-4|LNC|Thoracic outlet US|Thoracic outlet US
C0801762|T102|relax|26211-3|LNC|Thoracic outlet bilateral MRI|Thoracic outlet bilateral MRI
C0801762|T102|relax|26212-1|LNC|Thoracic outlet left MRI|Thoracic outlet left MRI
C0801762|T102|relax|26213-9|LNC|Thoracic outlet right MRI|Thoracic outlet right MRI
C0801762|T102|relax|43507-3|LNC|Thymus gland MRI|Thymus gland MRI
C0801762|T102|relax|42300-4|LNC|Thyroid MRI|Thyroid MRI
C0801762|T102|relax|25010-0|LNC|Thyroid US|Thyroid US
C0801762|T102|relax|37898-4|LNC|Tibia Fibula X-ray tomograph|Tibia Fibula X-ray tomograph
C0801762|T102|relax|30888-2|LNC|Tibioperoneal vessels MRI angiogram|Tibioperoneal vessels MRI angiogram
C0801762|T102|relax|36780-5|LNC|Toe MRI|Toe MRI
C0801762|T102|relax|69285-5|LNC|Umbilical artery US doppler|Umbilical artery US doppler
C0801762|T102|relax|39508-7|LNC|Umbilical vessels US doppler|Umbilical vessels US doppler
C0801762|T102|relax|36023-0|LNC|Upper arm CT|Upper arm CT
C0801762|T102|relax|36025-5|LNC|Upper arm MRI|Upper arm MRI
C0801762|T102|relax|36026-3|LNC|Upper arm bilateral CT|Upper arm bilateral CT
C0801762|T102|relax|69180-8|LNC|Upper arm bilateral MRI|Upper arm bilateral MRI
C0801762|T102|relax|36027-1|LNC|Upper arm left CT|Upper arm left CT
C0801762|T102|relax|36028-9|LNC|Upper arm left MRI|Upper arm left MRI
C0801762|T102|relax|36029-7|LNC|Upper arm right CT|Upper arm right CT
C0801762|T102|relax|36030-5|LNC|Upper arm right MRI|Upper arm right MRI
C0801762|T102|relax|35981-0|LNC|Upper extremity CT|Upper extremity CT
C0801762|T102|relax|24688-4|LNC|Upper extremity MRI|Upper extremity MRI
C0801762|T102|relax|30710-8|LNC|Upper extremity US|Upper extremity US
C0801762|T102|relax|37923-0|LNC|Upper extremity X-ray tomograph|Upper extremity X-ray tomograph
C0801762|T102|relax|48448-5|LNC|Upper extremity artery US|Upper extremity artery US
C0801762|T102|relax|39447-8|LNC|Upper extremity artery US doppler|Upper extremity artery US doppler
C0801762|T102|relax|38014-7|LNC|Upper extremity artery bilateral US|Upper extremity artery bilateral US
C0801762|T102|relax|39423-9|LNC|Upper extremity artery bilateral US doppler|Upper extremity artery bilateral US doppler
C0801762|T102|relax|41833-5|LNC|Upper extremity artery left US|Upper extremity artery left US
C0801762|T102|relax|39500-4|LNC|Upper extremity artery left US doppler|Upper extremity artery left US doppler
C0801762|T102|relax|41814-5|LNC|Upper extremity artery right US|Upper extremity artery right US
C0801762|T102|relax|39506-1|LNC|Upper extremity artery right US doppler|Upper extremity artery right US doppler
C0801762|T102|relax|30882-5|LNC|Upper extremity vein US doppler|Upper extremity vein US doppler
C0801762|T102|relax|48690-2|LNC|Upper extremity vein bilateral US|Upper extremity vein bilateral US
C0801762|T102|relax|39496-5|LNC|Upper extremity vein bilateral US doppler|Upper extremity vein bilateral US doppler
C0801762|T102|relax|48689-4|LNC|Upper extremity vein left US|Upper extremity vein left US
C0801762|T102|relax|39501-2|LNC|Upper extremity vein left US doppler|Upper extremity vein left US doppler
C0801762|T102|relax|48688-6|LNC|Upper extremity vein right US|Upper extremity vein right US
C0801762|T102|relax|39507-9|LNC|Upper extremity vein right US doppler|Upper extremity vein right US doppler
C0801762|T102|relax|36080-0|LNC|Upper extremity veins MRI angiogram|Upper extremity veins MRI angiogram
C0801762|T102|relax|69395-2|LNC|Upper extremity veins US|Upper extremity veins US
C0801762|T102|relax|36786-2|LNC|Upper extremity veins left MRI angiogram|Upper extremity veins left MRI angiogram
C0801762|T102|relax|36787-0|LNC|Upper extremity veins right MRI angiogram|Upper extremity veins right MRI angiogram
C0801762|T102|relax|46385-1|LNC|Upper extremity vessel graft US doppler|Upper extremity vessel graft US doppler
C0801762|T102|relax|44236-8|LNC|Upper extremity vessel graft bilateral US doppler|Upper extremity vessel graft bilateral US doppler
C0801762|T102|relax|42475-4|LNC|Upper extremity vessel graft left US doppler|Upper extremity vessel graft left US doppler
C0801762|T102|relax|42476-2|LNC|Upper extremity vessel graft right US doppler|Upper extremity vessel graft right US doppler
C0801762|T102|relax|36084-2|LNC|Upper extremity vessels MRI angiogram|Upper extremity vessels MRI angiogram
C0801762|T102|relax|39448-6|LNC|Upper extremity vessels US doppler|Upper extremity vessels US doppler
C0801762|T102|relax|46379-4|LNC|Upper extremity vessels bilateral US doppler|Upper extremity vessels bilateral US doppler
C0801762|T102|relax|36797-9|LNC|Upper extremity vessels left MRI angiogram|Upper extremity vessels left MRI angiogram
C0801762|T102|relax|39433-8|LNC|Upper extremity vessels left US doppler|Upper extremity vessels left US doppler
C0801762|T102|relax|36798-7|LNC|Upper extremity vessels right MRI angiogram|Upper extremity vessels right MRI angiogram
C0801762|T102|relax|39444-5|LNC|Upper extremity vessels right US doppler|Upper extremity vessels right US doppler
C0801762|T102|relax|26232-9|LNC|Upper extremity bilateral MRI|Upper extremity bilateral MRI
C0801762|T102|relax|30875-9|LNC|Upper extremity  joint MRI|Upper extremity  joint MRI
C0801762|T102|relax|36774-8|LNC|Upper extremity joint left MRI|Upper extremity joint left MRI
C0801762|T102|relax|36775-5|LNC|Upper extremity joint right MRI|Upper extremity joint right MRI
C0801762|T102|relax|35982-8|LNC|Upper extremity left CT|Upper extremity left CT
C0801762|T102|relax|26233-7|LNC|Upper extremity left MRI|Upper extremity left MRI
C0801762|T102|relax|38041-0|LNC|Upper extremity left US|Upper extremity left US
C0801762|T102|relax|35983-6|LNC|Upper extremity right CT|Upper extremity right CT
C0801762|T102|relax|26234-5|LNC|Upper extremity right MRI|Upper extremity right MRI
C0801762|T102|relax|38052-7|LNC|Upper extremity right US|Upper extremity right US
C0801762|T102|relax|25019-1|LNC|Urinary bladder US|Urinary bladder US
C0801762|T102|relax|42301-2|LNC|Uterus MRI|Uterus MRI
C0801762|T102|relax|30705-8|LNC|Uterus Fallopian tubes US|Uterus Fallopian tubes US
C0801762|T102|relax|39036-9|LNC|Vein US|Vein US
C0801762|T102|relax|39525-1|LNC|Vein US doppler|Vein US doppler
C0801762|T102|relax|39030-2|LNC|Vein bilateral US|Vein bilateral US
C0801762|T102|relax|36783-9|LNC|Veins MRI angiogram|Veins MRI angiogram
C0801762|T102|relax|69222-8|LNC|Vena cava MRI|Vena cava MRI
C0801762|T102|relax|36081-8|LNC|Vena cava MRI angiogram|Vena cava MRI angiogram
C0801762|T102|relax|36083-4|LNC|Inferior vena cava MRI|Inferior vena cava MRI
C0801762|T102|relax|36082-6|LNC|Inferior vena cava MRI angiogram|Inferior vena cava MRI angiogram
C0801762|T102|relax|36790-4|LNC|Vena cava inferior Lower extremity veins MRI angiogram|Vena cava inferior Lower extremity veins MRI angiogram
C0801762|T102|relax|39445-2|LNC|Vessels US doppler|Vessels US doppler
C0801762|T102|relax|38054-3|LNC|Visceral artery US|Visceral artery US
C0801762|T102|relax|37428-0|LNC|Wrist CT|Wrist CT
C0801762|T102|relax|25033-2|LNC|Wrist MRI|Wrist MRI
C0801762|T102|relax|25036-5|LNC|Wrist US|Wrist US
C0801762|T102|relax|37932-1|LNC|Wrist X-ray tomograph|Wrist X-ray tomograph
C0801762|T102|relax|37430-6|LNC|Wrist bilateral CT|Wrist bilateral CT
C0801762|T102|relax|26277-4|LNC|Wrist bilateral MRI|Wrist bilateral MRI
C0801762|T102|relax|26278-2|LNC|Wrist bilateral US|Wrist bilateral US
C0801762|T102|relax|37429-8|LNC|Wrist bilateral X-ray tomograph|Wrist bilateral X-ray tomograph
C0801762|T102|relax|37431-4|LNC|Wrist left CT|Wrist left CT
C0801762|T102|relax|26279-0|LNC|Wrist left MRI|Wrist left MRI
C0801762|T102|relax|26280-8|LNC|Wrist left US|Wrist left US
C0801762|T102|relax|37432-2|LNC|Wrist left X-ray tomograph|Wrist left X-ray tomograph
C0801762|T102|relax|69209-5|LNC|Wrist left Hand left MRI|Wrist left Hand left MRI
C0801762|T102|relax|37433-0|LNC|Wrist right CT|Wrist right CT
C0801762|T102|relax|26281-6|LNC|Wrist right MRI|Wrist right MRI
C0801762|T102|relax|26282-4|LNC|Wrist right US|Wrist right US
C0801762|T102|relax|37644-2|LNC|Wrist right X-ray tomograph|Wrist right X-ray tomograph
C0801762|T102|relax|69219-4|LNC|Wrist right Hand right MRI|Wrist right Hand right MRI
C0801762|T102|relax|36008-1|LNC|Wrist Hand MRI|Wrist Hand MRI
C0801762|T102|relax|25045-6|LNC|Unspecified body region CT|Unspecified body region CT
C0801762|T102|relax|25040-7|LNC|Unspecified body region CT 3D|Unspecified body region CT 3D
C0801762|T102|relax|25056-3|LNC|Unspecified body region MRI|Unspecified body region MRI
C0801762|T102|relax|44136-0|LNC|Unspecified body region PET|Unspecified body region PET
C0801762|T102|relax|25061-3|LNC|Unspecified body region US|Unspecified body region US
C0801762|T102|relax|25071-2|LNC|Unspecified body region X-ray tomograph|Unspecified body region X-ray tomograph
C0801762|T102|relax|46375-2|LNC|Artery US|Artery US
C0801762|T102|relax|39523-6|LNC|Artery US doppler|Artery US doppler
C0801762|T102|relax|44229-3|LNC|Bones CT|Bones CT
C0801762|T102|relax|28576-7|LNC|Joint MRI|Joint MRI
C0801762|T102|relax|39453-6|LNC|Tendon US|Tendon US
C0801762|T102|relax|36957-9|LNC|Facial bones Maxilla CT 3D reconstruction|Facial bones Maxilla CT 3D reconstruction
C0801762|T102|relax|37294-6|LNC|Head CT 3D reconstruction|Head CT 3D reconstruction
C0801762|T102|relax|41804-6|LNC|Unspecified body region CT 3D reconstruction|Unspecified body region CT 3D reconstruction
C0801762|T102|relax|39043-5|LNC|Unspecified body region MRI 3D reconstruction|Unspecified body region MRI 3D reconstruction
C0801762|T102|relax|44165-9|LNC|Unspecified body region US 3D reconstruction|Unspecified body region US 3D reconstruction
C0801762|T102|relax|58745-1|LNC|Coronary arteries CT angiogram 3D reconstruction W contrast IV|Coronary arteries CT angiogram 3D reconstruction W contrast IV
C0801762|T102|relax|59255-0|LNC|Left atrium Pulmonary veins CT angiogram 3D reconstruction W contrast IV|Left atrium Pulmonary veins CT angiogram 3D reconstruction W contrast IV
C0801762|T102|relax|69082-6|LNC|Head CT 3D reconstruction WO contrast|Head CT 3D reconstruction WO contrast
C0801762|T102|relax|37295-3|LNC|Femur Hip CT anteversion measurement|Femur Hip CT anteversion measurement
C0801762|T102|relax|72830-3|LNC|Extremity arteries bilateral US doppler Multisection physiologic artery study|Extremity arteries bilateral US doppler Multisection physiologic artery study
C0801762|T102|relax|72832-9|LNC|Extremity arteries bilateral US doppler Multisection physiologic artery study at rest & W exercise|Extremity arteries bilateral US doppler Multisection physiologic artery study at rest & W exercise
C0801762|T102|relax|39879-2|LNC|Bone SPECT 1 phase|Bone SPECT 1 phase
C0801762|T102|relax|39881-8|LNC|Bone SPECT 3 phase whole body|Bone SPECT 3 phase whole body
C0801762|T102|relax|30760-3|LNC|Kidney bilateral X-ray tomograph 3 views W contrast IV|Kidney bilateral X-ray tomograph 3 views W contrast IV
C0801762|T102|relax|25055-5|LNC|Unspecified body region MRI additional sequence|Unspecified body region MRI additional sequence
C0801762|T102|relax|39408-0|LNC|Spine Thoracic X-ray tomograph AP|Spine Thoracic X-ray tomograph AP
C0801762|T102|relax|39862-8|LNC|Heart SPECT blood pool at rest W radionuclide IV|Heart SPECT blood pool at rest W radionuclide IV
C0801762|T102|relax|47378-5|LNC|Liver SPECT blood pool|Liver SPECT blood pool
C0801762|T102|relax|37435-5|LNC|Temporomandibular joint MRI cine|Temporomandibular joint MRI cine
C0801762|T102|relax|42693-2|LNC|Urinary Bladder Urethra MRI cine|Urinary Bladder Urethra MRI cine
C0801762|T102|relax|39140-9|LNC|Heart MRI cine blood flow velocity mapping|Heart MRI cine blood flow velocity mapping
C0801762|T102|relax|44126-1|LNC|Heart MRI cine blood flow velocity mapping W contrast IV|Heart MRI cine blood flow velocity mapping W contrast IV
C0801762|T102|relax|42386-3|LNC|Brain MRI cine CSF flow|Brain MRI cine CSF flow
C0801762|T102|relax|42387-1|LNC|Unspecified body region MRI cine CSF flow|Unspecified body region MRI cine CSF flow
C0801762|T102|relax|37434-8|LNC|Heart MRI cine function|Heart MRI cine function
C0801762|T102|relax|46300-0|LNC|Sinuses CT coronal|Sinuses CT coronal
C0801762|T102|relax|72139-9|LNC|Breast bilateral FFD mammogram-tomosynthesis diagnostic|Breast bilateral FFD mammogram-tomosynthesis diagnostic
C0801762|T102|relax|72138-1|LNC|Breast left FFD mammogram-tomosynthesis diagnostic|Breast left FFD mammogram-tomosynthesis diagnostic
C0801762|T102|relax|72137-3|LNC|Breast right FFD mammogram-tomosynthesis diagnostic|Breast right FFD mammogram-tomosynthesis diagnostic
C0801762|T102|relax|37436-3|LNC|Brain MRI diffusion weighted|Brain MRI diffusion weighted
C0801762|T102|relax|43555-2|LNC|Ankle left MRI dynamic W contrast IV|Ankle left MRI dynamic W contrast IV
C0801762|T102|relax|43449-8|LNC|Ankle right MRI dynamic W contrast IV|Ankle right MRI dynamic W contrast IV
C0801762|T102|relax|37437-1|LNC|Breast MRI dynamic W contrast IV|Breast MRI dynamic W contrast IV
C0801762|T102|relax|36114-7|LNC|Breast bilateral MRI dynamic W contrast IV|Breast bilateral MRI dynamic W contrast IV
C0801762|T102|relax|43450-6|LNC|Elbow left MRI dynamic W contrast IV|Elbow left MRI dynamic W contrast IV
C0801762|T102|relax|43451-4|LNC|Elbow right MRI dynamic W contrast IV|Elbow right MRI dynamic W contrast IV
C0801762|T102|relax|46394-3|LNC|Head CT dynamic W contrast IV|Head CT dynamic W contrast IV
C0801762|T102|relax|43452-2|LNC|Knee left MRI dynamic W contrast IV|Knee left MRI dynamic W contrast IV
C0801762|T102|relax|43453-0|LNC|Knee right MRI dynamic W contrast IV|Knee right MRI dynamic W contrast IV
C0801762|T102|relax|37438-9|LNC|Pituitary Sella turcica CT dynamic W contrast IV|Pituitary Sella turcica CT dynamic W contrast IV
C0801762|T102|relax|43527-1|LNC|Unspecified body region CT dynamic W contrast IV|Unspecified body region CT dynamic W contrast IV
C0801762|T102|relax|39637-4|LNC|Brain SPECT flow|Brain SPECT flow
C0801762|T102|relax|43655-0|LNC|Liver SPECT flow|Liver SPECT flow
C0801762|T102|relax|43652-7|LNC|Liver Spleen SPECT flow|Liver Spleen SPECT flow
C0801762|T102|relax|69235-0|LNC|Scrotum Testicle SPECT flow|Scrotum Testicle SPECT flow
C0801762|T102|relax|43670-9|LNC|Spleen SPECT flow|Spleen SPECT flow
C0801762|T102|relax|43673-3|LNC|Thyroid SPECT flow|Thyroid SPECT flow
C0801762|T102|relax|43662-6|LNC|Renal vessels SPECT flow W Tc-99m glucoheptonate IV|Renal vessels SPECT flow W Tc-99m glucoheptonate IV
C0801762|T102|relax|39684-6|LNC|SPECT abscess W GA-67 IV|SPECT abscess W GA-67 IV
C0801762|T102|relax|39811-5|LNC|SPECT abscess|SPECT abscess
C0801762|T102|relax|39141-7|LNC|Bone marrow MRI blood flow|Bone marrow MRI blood flow
C0801762|T102|relax|39656-4|LNC|Heart SPECT infarct|Heart SPECT infarct
C0801762|T102|relax|39654-9|LNC|Heart SPECT infarct W Tc-99m PYP IV|Heart SPECT infarct W Tc-99m PYP IV
C0801762|T102|relax|39655-6|LNC|Heart SPECT infarct W Tc-99m Sestamibi IV|Heart SPECT infarct W Tc-99m Sestamibi IV
C0801762|T102|relax|39675-4|LNC|SPECT infection W GA-67 IV|SPECT infection W GA-67 IV
C0801762|T102|relax|72251-2|LNC|Chest vessels CT Multisection pulmonary embolus|Chest vessels CT Multisection pulmonary embolus
C0801762|T102|relax|24889-8|LNC|Pylorus US pyloric stenosis|Pylorus US pyloric stenosis
C0801762|T102|relax|36934-8|LNC|Heart CT scoring|Heart CT scoring
C0801762|T102|relax|36935-5|LNC|Heart CT scoring W contrast IV|Heart CT scoring W contrast IV
C0801762|T102|relax|43446-4|LNC|CT tumor whole body|CT tumor whole body
C0801762|T102|relax|69237-6|LNC|SPECT tumor whole body|SPECT tumor whole body
C0801762|T102|relax|39678-8|LNC|SPECT tumor W GA-67 IV|SPECT tumor W GA-67 IV
C0801762|T102|relax|39748-9|LNC|SPECT tumor W Tc-99m Sestamibi IV|SPECT tumor W Tc-99m Sestamibi IV
C0801762|T102|relax|42292-3|LNC|SPECT tumor W Tl-201 IV|SPECT tumor W Tl-201 IV
C0801762|T102|relax|46395-0|LNC|Heart SPECT gated ejection fraction at rest W stress W radionuclide IV|Heart SPECT gated ejection fraction at rest W stress W radionuclide IV
C0801762|T102|relax|39913-9|LNC|Heart SPECT gated ejection fraction|Heart SPECT gated ejection fraction
C0801762|T102|relax|39918-8|LNC|Heart SPECT gated wall motion|Heart SPECT gated wall motion
C0801762|T102|relax|46396-8|LNC|Heart SPECT gated at rest W Tc-99m Sestamibi IV|Heart SPECT gated at rest W Tc-99m Sestamibi IV
C0801762|T102|relax|39916-2|LNC|Heart SPECT gated|Heart SPECT gated
C0801762|T102|relax|39930-3|LNC|Heart SPECT gated W stress W radionuclide IV|Heart SPECT gated W stress W radionuclide IV
C0801762|T102|relax|37439-7|LNC|Chest CT high resolution|Chest CT high resolution
C0801762|T102|relax|37440-5|LNC|Chest CT high resolution W contrast IV|Chest CT high resolution W contrast IV
C0801762|T102|relax|37441-3|LNC|Chest CT high resolution WO contrast|Chest CT high resolution WO contrast
C0801762|T102|relax|39409-8|LNC|Spine Thoracic X-ray tomograph lateral|Spine Thoracic X-ray tomograph lateral
C0801762|T102|relax|36086-7|LNC|Abdomen CT limited|Abdomen CT limited
C0801762|T102|relax|30704-1|LNC|Abdomen US limited|Abdomen US limited
C0801762|T102|relax|38047-7|LNC|Abdomen retroperitoneum US limited|Abdomen retroperitoneum US limited
C0801762|T102|relax|43572-7|LNC|Abdominal vessels US doppler limited|Abdominal vessels US doppler limited
C0801762|T102|relax|38011-3|LNC|Aorta US limited|Aorta US limited
C0801762|T102|relax|69280-6|LNC|Bladder US limited|Bladder US limited
C0801762|T102|relax|24599-3|LNC|Breast US limited|Breast US limited
C0801762|T102|relax|26286-5|LNC|Breast bilateral US limited|Breast bilateral US limited
C0801762|T102|relax|26288-1|LNC|Breast left US limited|Breast left US limited
C0801762|T102|relax|26290-7|LNC|Breast right US limited|Breast right US limited
C0801762|T102|relax|38015-4|LNC|Carotid artery US limited|Carotid artery US limited
C0801762|T102|relax|42149-5|LNC|Carotid artery left US limited|Carotid artery left US limited
C0801762|T102|relax|42151-1|LNC|Carotid artery right US limited|Carotid artery right US limited
C0801762|T102|relax|36089-1|LNC|Chest CT limited|Chest CT limited
C0801762|T102|relax|69281-4|LNC|Chest US limited|Chest US limited
C0801762|T102|relax|36090-9|LNC|Extremity CT limited|Extremity CT limited
C0801762|T102|relax|39526-9|LNC|Extremity US limited|Extremity US limited
C0801762|T102|relax|46301-8|LNC|Extremity vein bilateral US doppler limited|Extremity vein bilateral US doppler limited
C0801762|T102|relax|39424-7|LNC|Extremity vessels US doppler limited|Extremity vessels US doppler limited
C0801762|T102|relax|62451-0|LNC|Extremity left US limited|Extremity left US limited
C0801762|T102|relax|62452-8|LNC|Extremity right US limited|Extremity right US limited
C0801762|T102|relax|69286-3|LNC|Eye US limited|Eye US limited
C0801762|T102|relax|36937-1|LNC|Facial bones Maxilla CT limited|Facial bones Maxilla CT limited
C0801762|T102|relax|38020-4|LNC|Gallbladder US limited|Gallbladder US limited
C0801762|T102|relax|36087-5|LNC|Head CT limited|Head CT limited
C0801762|T102|relax|38034-5|LNC|Head US limited|Head US limited
C0801762|T102|relax|36808-4|LNC|Head vessels MRI angiogram limited|Head vessels MRI angiogram limited
C0801762|T102|relax|39044-3|LNC|Head vessels US doppler limited|Head vessels US doppler limited
C0801762|T102|relax|36091-7|LNC|Heart MRI limited|Heart MRI limited
C0801762|T102|relax|42707-0|LNC|Heart US limited|Heart US limited
C0801762|T102|relax|36092-5|LNC|Hip CT limited|Hip CT limited
C0801762|T102|relax|43776-4|LNC|Iliac artery US doppler limited|Iliac artery US doppler limited
C0801762|T102|relax|42150-3|LNC|Iliac graft US doppler limited|Iliac graft US doppler limited
C0801762|T102|relax|36088-3|LNC|Internal auditory canal MRI limited|Internal auditory canal MRI limited
C0801762|T102|relax|38035-2|LNC|Kidney US limited|Kidney US limited
C0801762|T102|relax|69300-2|LNC|Kidney transplant US limited|Kidney transplant US limited
C0801762|T102|relax|41812-9|LNC|Lower extremity artery US limited|Lower extremity artery US limited
C0801762|T102|relax|38042-8|LNC|Lower extremity artery US doppler limited|Lower extremity artery US doppler limited
C0801762|T102|relax|39430-4|LNC|Lower extremity vessels left US doppler limited|Lower extremity vessels left US doppler limited
C0801762|T102|relax|39441-1|LNC|Lower extremity vessels right US doppler limited|Lower extremity vessels right US doppler limited
C0801762|T102|relax|36093-3|LNC|Lower Extremity Joint MRI limited|Lower Extremity Joint MRI limited
C0801762|T102|relax|38039-4|LNC|Lower extremity left US limited|Lower extremity left US limited
C0801762|T102|relax|38050-1|LNC|Lower extremity right US limited|Lower extremity right US limited
C0801762|T102|relax|44116-2|LNC|Mandible CT limited|Mandible CT limited
C0801762|T102|relax|48461-8|LNC|Neck MRI limited|Neck MRI limited
C0801762|T102|relax|69212-9|LNC|Pelvis MRI limited|Pelvis MRI limited
C0801762|T102|relax|38046-9|LNC|Pelvis US limited|Pelvis US limited
C0801762|T102|relax|42152-9|LNC|Pelvis vessels US doppler limited|Pelvis vessels US doppler limited
C0801762|T102|relax|44173-3|LNC|Peripheral artery US limited|Peripheral artery US limited
C0801762|T102|relax|39436-1|LNC|Renal vessels US doppler limited|Renal vessels US doppler limited
C0801762|T102|relax|69299-6|LNC|Scrotum Testicle US limited|Scrotum Testicle US limited
C0801762|T102|relax|24913-6|LNC|Sinuses CT limited|Sinuses CT limited
C0801762|T102|relax|41813-7|LNC|Upper extremity artery US limited|Upper extremity artery US limited
C0801762|T102|relax|38143-4|LNC|Upper extremity artery US doppler limited|Upper extremity artery US doppler limited
C0801762|T102|relax|46302-6|LNC|Upper extremity artery bilateral US doppler limited|Upper extremity artery bilateral US doppler limited
C0801762|T102|relax|44237-6|LNC|Upper extremity vessel graft bilateral US doppler limited|Upper extremity vessel graft bilateral US doppler limited
C0801762|T102|relax|46303-4|LNC|Upper extremity vessels US doppler limited|Upper extremity vessels US doppler limited
C0801762|T102|relax|36094-1|LNC|Upper extremity  joint MRI limited|Upper extremity  joint MRI limited
C0801762|T102|relax|39045-0|LNC|Vein US limited|Vein US limited
C0801762|T102|relax|39524-4|LNC|Vein US doppler limited|Vein US doppler limited
C0801762|T102|relax|25039-9|LNC|Unspecified body region CT limited|Unspecified body region CT limited
C0801762|T102|relax|48460-0|LNC|Unspecified body region MRI limited|Unspecified body region MRI limited
C0801762|T102|relax|69282-2|LNC|Unspecified body region US doppler limited|Unspecified body region US doppler limited
C0801762|T102|relax|72831-1|LNC|Extremity arteries bilateral US doppler Multisection limited physiologic artery study|Extremity arteries bilateral US doppler Multisection limited physiologic artery study
C0801762|T102|relax|44127-9|LNC|Heart MRI limited cine function|Heart MRI limited cine function
C0801762|T102|relax|39046-8|LNC|Pelvis CT limited pelvimetry WO contrast|Pelvis CT limited pelvimetry WO contrast
C0801762|T102|relax|36102-2|LNC|Abdomen CT limited W WO contrast IV|Abdomen CT limited W WO contrast IV
C0801762|T102|relax|36095-8|LNC|Abdomen CT limited W contrast IV|Abdomen CT limited W contrast IV
C0801762|T102|relax|36096-6|LNC|Brain MRI limited W contrast IV|Brain MRI limited W contrast IV
C0801762|T102|relax|69096-6|LNC|Chest CT limited W contrast IV|Chest CT limited W contrast IV
C0801762|T102|relax|36098-2|LNC|Pelvis CT limited W contrast IV|Pelvis CT limited W contrast IV
C0801762|T102|relax|36099-0|LNC|Spine Cervical CT limited W contrast IV|Spine Cervical CT limited W contrast IV
C0801762|T102|relax|36100-6|LNC|Spine Lumbar MRI limited W contrast IV|Spine Lumbar MRI limited W contrast IV
C0801762|T102|relax|36101-4|LNC|Spine Thoracic MRI limited W contrast IV|Spine Thoracic MRI limited W contrast IV
C0801762|T102|relax|36097-4|LNC|Upper extremity CT limited W contrast IV|Upper extremity CT limited W contrast IV
C0801762|T102|relax|39681-2|LNC|SPECT limited W GA-67 IV|SPECT limited W GA-67 IV
C0801762|T102|relax|39813-1|LNC|Bone SPECT limited|Bone SPECT limited
C0801762|T102|relax|39821-4|LNC|Bone marrow SPECT limited|Bone marrow SPECT limited
C0801762|T102|relax|36103-0|LNC|Abdomen CT limited WO contrast|Abdomen CT limited WO contrast
C0801762|T102|relax|36105-5|LNC|Brain MRI limited WO contrast|Brain MRI limited WO contrast
C0801762|T102|relax|47366-0|LNC|Chest CT limited WO contrast|Chest CT limited WO contrast
C0801762|T102|relax|36938-9|LNC|Facial bones Maxilla CT limited WO contrast|Facial bones Maxilla CT limited WO contrast
C0801762|T102|relax|36104-8|LNC|Head CT limited WO contrast|Head CT limited WO contrast
C0801762|T102|relax|36106-3|LNC|Lower extremity CT limited WO contrast|Lower extremity CT limited WO contrast
C0801762|T102|relax|36107-1|LNC|Lower extremity joint left MRI limited WO contrast|Lower extremity joint left MRI limited WO contrast
C0801762|T102|relax|38769-6|LNC|Lower extremity joint right MRI limited WO contrast|Lower extremity joint right MRI limited WO contrast
C0801762|T102|relax|36108-9|LNC|Pelvis CT limited WO contrast|Pelvis CT limited WO contrast
C0801762|T102|relax|46304-2|LNC|Sinuses CT limited WO contrast|Sinuses CT limited WO contrast
C0801762|T102|relax|36109-7|LNC|Spine Cervical CT limited WO contrast|Spine Cervical CT limited WO contrast
C0801762|T102|relax|36110-5|LNC|Spine Lumbar CT limited WO contrast|Spine Lumbar CT limited WO contrast
C0801762|T102|relax|36111-3|LNC|Spine Lumbar MRI limited WO contrast|Spine Lumbar MRI limited WO contrast
C0801762|T102|relax|36112-1|LNC|Spine Thoracic MRI limited WO contrast|Spine Thoracic MRI limited WO contrast
C0801762|T102|relax|39905-5|LNC|Bone SPECT multiple areas|Bone SPECT multiple areas
C0801762|T102|relax|39906-3|LNC|Bone marrow SPECT multiple areas|Bone marrow SPECT multiple areas
C0801762|T102|relax|39527-7|LNC|Unspecified body region US foreign body|Unspecified body region US foreign body
C0801762|T102|relax|49569-7|LNC|Heart SPECT perfusion wall motion at rest W stress W Tl-201 IV W Tc-99m Sestamibi IV|Heart SPECT perfusion wall motion at rest W stress W Tl-201 IV W Tc-99m Sestamibi IV
C0801762|T102|relax|43659-2|LNC|Heart SPECT perfusion qualitative at rest W radionuclide IV|Heart SPECT perfusion qualitative at rest W radionuclide IV
C0801762|T102|relax|39725-7|LNC|Heart SPECT perfusion at rest W adenosine W Tl-201 IV|Heart SPECT perfusion at rest W adenosine W Tl-201 IV
C0801762|T102|relax|39718-2|LNC|Heart SPECT perfusion at rest W radionuclide IV|Heart SPECT perfusion at rest W radionuclide IV
C0801762|T102|relax|39724-0|LNC|Heart SPECT perfusion at rest W stress W radionuclide IV|Heart SPECT perfusion at rest W stress W radionuclide IV
C0801762|T102|relax|39723-2|LNC|Heart SPECT perfusion at rest W stress W Tl-201 IV|Heart SPECT perfusion at rest W stress W Tl-201 IV
C0801762|T102|relax|49568-9|LNC|Heart SPECT perfusion at rest W stress W Tl-201 IV W Tc-99m Sestamibi IV|Heart SPECT perfusion at rest W stress W Tl-201 IV W Tc-99m Sestamibi IV
C0801762|T102|relax|39729-9|LNC|Heart SPECT perfusion at rest W Tl-201 IV|Heart SPECT perfusion at rest W Tl-201 IV
C0801762|T102|relax|39700-0|LNC|Heart SPECT perfusion W adenosine W radionuclide IV|Heart SPECT perfusion W adenosine W radionuclide IV
C0801762|T102|relax|49567-1|LNC|Heart SPECT perfusion W adenosine W Tc-99m Sestamibi IV|Heart SPECT perfusion W adenosine W Tc-99m Sestamibi IV
C0801762|T102|relax|39142-5|LNC|Head CT perfusion W contrast IV|Head CT perfusion W contrast IV
C0801762|T102|relax|39712-5|LNC|Heart SPECT perfusion|Heart SPECT perfusion
C0801762|T102|relax|39734-9|LNC|Heart SPECT perfusion W stress W radionuclide IV|Heart SPECT perfusion W stress W radionuclide IV
C0801762|T102|relax|39736-4|LNC|Heart SPECT perfusion W stress W Tc-99m Sestamibi IV|Heart SPECT perfusion W stress W Tc-99m Sestamibi IV
C0801762|T102|relax|39710-9|LNC|Heart SPECT perfusion W Tc-99m Sestamibi IV|Heart SPECT perfusion W Tc-99m Sestamibi IV
C0801762|T102|relax|39711-7|LNC|Heart SPECT perfusion W Tl-201 IV|Heart SPECT perfusion W Tl-201 IV
C0801762|T102|relax|38060-0|LNC|Spine lumbosacral+Cervical+Thoracic MRI sagittal|Spine lumbosacral+Cervical+Thoracic MRI sagittal
C0801762|T102|relax|25052-2|LNC|Unspecified body region CT sagittal coronal|Unspecified body region CT sagittal coronal
C0801762|T102|relax|25050-6|LNC|Unspecified body region CT 3D sagittal coronal disarticulation|Unspecified body region CT 3D sagittal coronal disarticulation
C0801762|T102|relax|42132-1|LNC|Breast US screening|Breast US screening
C0801762|T102|relax|72142-3|LNC|Breast bilateral FFD mammogram-tomosynthesis screening|Breast bilateral FFD mammogram-tomosynthesis screening
C0801762|T102|relax|72141-5|LNC|Breast left FFD mammogram-tomosynthesis screening|Breast left FFD mammogram-tomosynthesis screening
C0801762|T102|relax|72140-7|LNC|Breast right FFD mammogram-tomosynthesis screening|Breast right FFD mammogram-tomosynthesis screening
C0801762|T102|relax|37442-1|LNC|Brain MRI spectroscopy|Brain MRI spectroscopy
C0801762|T102|relax|37443-9|LNC|Unspecified body region MRI spectroscopy|Unspecified body region MRI spectroscopy
C0801762|T102|relax|70929-5|LNC|Spine Cervical CT stereotactic|Spine Cervical CT stereotactic
C0801762|T102|relax|70928-7|LNC|Spine Lumbar CT stereotactic|Spine Lumbar CT stereotactic
C0801762|T102|relax|70930-3|LNC|Spine Thoracic CT stereotactic|Spine Thoracic CT stereotactic
C0801762|T102|relax|36940-5|LNC|Unspecified body region CT stereotactic|Unspecified body region CT stereotactic
C0801762|T102|relax|42455-6|LNC|Pelvis US transabdominal transvaginal|Pelvis US transabdominal transvaginal
C0801762|T102|relax|24677-7|LNC|Pelvis US transvaginal|Pelvis US transvaginal
C0801762|T102|relax|42390-5|LNC|Transvaginal MRI|Transvaginal MRI
C0801762|T102|relax|39838-8|LNC|Lung SPECT ventilation perfusion W radionuclide inhaled W radionuclide IV|Lung SPECT ventilation perfusion W radionuclide inhaled W radionuclide IV
C0801762|T102|relax|39898-2|LNC|Lung SPECT ventilation W radionuclide aerosol inhaled|Lung SPECT ventilation W radionuclide aerosol inhaled
C0801762|T102|relax|39872-7|LNC|Heart SPECT wall motion|Heart SPECT wall motion
C0801762|T102|relax|46305-9|LNC|CT whole body|CT whole body
C0801762|T102|relax|46358-8|LNC|MRI whole body|MRI whole body
C0801762|T102|relax|44139-4|LNC|PET whole body|PET whole body
C0801762|T102|relax|46306-7|LNC|CT whole body W contrast IV|CT whole body W contrast IV
C0801762|T102|relax|39680-4|LNC|SPECT whole body W GA-67 IV|SPECT whole body W GA-67 IV
C0801762|T102|relax|39816-4|LNC|Bone SPECT whole body|Bone SPECT whole body
C0801762|T102|relax|39825-5|LNC|Bone marrow SPECT whole body|Bone marrow SPECT whole body
C0801762|T102|relax|41837-6|LNC|SPECT whole body W Tc-99m Arcitumomab IV|SPECT whole body W Tc-99m Arcitumomab IV
C0801762|T102|relax|39658-0|LNC|Heart SPECT at rest W radionuclide IV|Heart SPECT at rest W radionuclide IV
C0801762|T102|relax|39662-2|LNC|Heart SPECT at rest W stress W Tc-99m Sestamibi IV|Heart SPECT at rest W stress W Tc-99m Sestamibi IV
C0801762|T102|relax|49566-3|LNC|Heart SPECT at rest W Tc-99m Sestamibi IV|Heart SPECT at rest W Tc-99m Sestamibi IV
C0801762|T102|relax|30711-6|LNC|Hip US developmental joint assessment|Hip US developmental joint assessment
C0801762|T102|relax|24732-0|LNC|Head US during surgery|Head US during surgery
C0801762|T102|relax|30706-6|LNC|Liver US during surgery|Liver US during surgery
C0801762|T102|relax|30701-7|LNC|Unspecified body region US during surgery|Unspecified body region US during surgery
C0801762|T102|relax|69388-7|LNC|Urinary bladder US post void|Urinary bladder US post void
C0801762|T102|relax|69086-7|LNC|Aorta CT W WO contrast|Aorta CT W WO contrast
C0801762|T102|relax|69108-9|LNC|Pulmonary vessels CT angiogram W WO contrast|Pulmonary vessels CT angiogram W WO contrast
C0801762|T102|relax|69085-9|LNC|Renal vessels CT angiogram W WO contrast|Renal vessels CT angiogram W WO contrast
C0801762|T102|relax|69207-9|LNC|Hip left MRI W WO contrast intraarticular|Hip left MRI W WO contrast intraarticular
C0801762|T102|relax|69217-8|LNC|Hip right MRI W WO contrast intraarticular|Hip right MRI W WO contrast intraarticular
C0801762|T102|relax|69208-7|LNC|Shoulder left MRI W WO contrast intraarticular|Shoulder left MRI W WO contrast intraarticular
C0801762|T102|relax|69218-6|LNC|Shoulder right MRI W WO contrast intraarticular|Shoulder right MRI W WO contrast intraarticular
C0801762|T102|relax|48450-1|LNC|Spine Cervical MRI W WO contrast IT|Spine Cervical MRI W WO contrast IT
C0801762|T102|relax|44114-7|LNC|Spine Lumbar CT W WO contrast IT|Spine Lumbar CT W WO contrast IT
C0801762|T102|relax|48452-7|LNC|Spine Lumbar MRI W WO contrast IT|Spine Lumbar MRI W WO contrast IT
C0801762|T102|relax|44113-9|LNC|Spine Thoracic CT W WO contrast IT|Spine Thoracic CT W WO contrast IT
C0801762|T102|relax|48441-0|LNC|Spine Thoracic MRI W WO contrast IT|Spine Thoracic MRI W WO contrast IT
C0801762|T102|relax|36267-3|LNC|Abdomen CT W WO contrast IV|Abdomen CT W WO contrast IV
C0801762|T102|relax|24557-1|LNC|Abdomen MRI W WO contrast IV|Abdomen MRI W WO contrast IV
C0801762|T102|relax|48743-9|LNC|Abdomen retroperitoneum CT W WO contrast IV|Abdomen retroperitoneum CT W WO contrast IV
C0801762|T102|relax|42274-1|LNC|Abdomen Pelvis CT W WO contrast IV|Abdomen Pelvis CT W WO contrast IV
C0801762|T102|relax|36846-4|LNC|Abdominal veins MRI angiogram W WO contrast IV|Abdominal veins MRI angiogram W WO contrast IV
C0801762|T102|relax|30805-6|LNC|Abdominal vessels CT angiogram W WO contrast IV|Abdominal vessels CT angiogram W WO contrast IV
C0801762|T102|relax|36855-5|LNC|Abdominal vessels MRI angiogram W WO contrast IV|Abdominal vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|36950-4|LNC|Adrenal gland CT W WO contrast IV|Adrenal gland CT W WO contrast IV
C0801762|T102|relax|36951-2|LNC|Adrenal gland MRI W WO contrast IV|Adrenal gland MRI W WO contrast IV
C0801762|T102|relax|36268-1|LNC|Ankle CT W WO contrast IV|Ankle CT W WO contrast IV
C0801762|T102|relax|24539-9|LNC|Ankle MRI W WO contrast IV|Ankle MRI W WO contrast IV
C0801762|T102|relax|26187-5|LNC|Ankle bilateral MRI W WO contrast IV|Ankle bilateral MRI W WO contrast IV
C0801762|T102|relax|36269-9|LNC|Ankle left CT W WO contrast IV|Ankle left CT W WO contrast IV
C0801762|T102|relax|26188-3|LNC|Ankle left MRI W WO contrast IV|Ankle left MRI W WO contrast IV
C0801762|T102|relax|36270-7|LNC|Ankle right CT W WO contrast IV|Ankle right CT W WO contrast IV
C0801762|T102|relax|26189-1|LNC|Ankle right MRI W WO contrast IV|Ankle right MRI W WO contrast IV
C0801762|T102|relax|44131-1|LNC|Aorta MRI angiogram W WO contrast IV|Aorta MRI angiogram W WO contrast IV
C0801762|T102|relax|36271-5|LNC|Aorta abdominal CT W WO contrast IV|Aorta abdominal CT W WO contrast IV
C0801762|T102|relax|36273-1|LNC|Aorta abdominal MRI W WO contrast IV|Aorta abdominal MRI W WO contrast IV
C0801762|T102|relax|36272-3|LNC|Aorta abdominal MRI angiogram W WO contrast IV|Aorta abdominal MRI angiogram W WO contrast IV
C0801762|T102|relax|36274-9|LNC|Aorta thoracic MRI angiogram W WO contrast IV|Aorta thoracic MRI angiogram W WO contrast IV
C0801762|T102|relax|30806-4|LNC|Aorta Femoral artery bilateral CT angiogram W WO contrast IV|Aorta Femoral artery bilateral CT angiogram W WO contrast IV
C0801762|T102|relax|46360-4|LNC|Aortic arch MRI angiogram W WO contrast IV|Aortic arch MRI angiogram W WO contrast IV
C0801762|T102|relax|43509-9|LNC|Axilla left MRI W WO contrast IV|Axilla left MRI W WO contrast IV
C0801762|T102|relax|43511-5|LNC|Axilla right MRI W WO contrast IV|Axilla right MRI W WO contrast IV
C0801762|T102|relax|36944-7|LNC|Biliary ducts Pancreatic duct MRI W WO contrast IV|Biliary ducts Pancreatic duct MRI W WO contrast IV
C0801762|T102|relax|24587-8|LNC|Brain MRI W WO contrast IV|Brain MRI W WO contrast IV
C0801762|T102|relax|48694-4|LNC|Brain temporal MRI W WO contrast IV|Brain temporal MRI W WO contrast IV
C0801762|T102|relax|43769-9|LNC|Brain Internal auditory canal MRI W WO contrast IV|Brain Internal auditory canal MRI W WO contrast IV
C0801762|T102|relax|42392-1|LNC|Brain Pituitary Sella turcica MRI W WO contrast IV|Brain Pituitary Sella turcica MRI W WO contrast IV
C0801762|T102|relax|36276-4|LNC|Breast MRI W WO contrast IV|Breast MRI W WO contrast IV
C0801762|T102|relax|69189-9|LNC|Breast implant MRI W WO contrast IV|Breast implant MRI W WO contrast IV
C0801762|T102|relax|69166-7|LNC|Breast implant bilateral MRI W WO contrast IV|Breast implant bilateral MRI W WO contrast IV
C0801762|T102|relax|38870-2|LNC|Breast implant left MRI W WO contrast IV|Breast implant left MRI W WO contrast IV
C0801762|T102|relax|38062-6|LNC|Breast implant right MRI W WO contrast IV|Breast implant right MRI W WO contrast IV
C0801762|T102|relax|36277-2|LNC|Breast bilateral MRI W WO contrast IV|Breast bilateral MRI W WO contrast IV
C0801762|T102|relax|36278-0|LNC|Breast left MRI W WO contrast IV|Breast left MRI W WO contrast IV
C0801762|T102|relax|36279-8|LNC|Breast right MRI W WO contrast IV|Breast right MRI W WO contrast IV
C0801762|T102|relax|43528-9|LNC|Breast unilateral MRI W WO contrast IV|Breast unilateral MRI W WO contrast IV
C0801762|T102|relax|36358-0|LNC|Calcaneus CT W WO contrast IV|Calcaneus CT W WO contrast IV
C0801762|T102|relax|36280-6|LNC|Calcaneus left CT W WO contrast IV|Calcaneus left CT W WO contrast IV
C0801762|T102|relax|36281-4|LNC|Calcaneus right CT W WO contrast IV|Calcaneus right CT W WO contrast IV
C0801762|T102|relax|36856-3|LNC|Carotid vessel MRI angiogram W WO contrast IV|Carotid vessel MRI angiogram W WO contrast IV
C0801762|T102|relax|30598-7|LNC|Chest CT W WO contrast IV|Chest CT W WO contrast IV
C0801762|T102|relax|36283-0|LNC|Chest MRI W WO contrast IV|Chest MRI W WO contrast IV
C0801762|T102|relax|36848-0|LNC|Chest veins MRI angiogram W WO contrast IV|Chest veins MRI angiogram W WO contrast IV
C0801762|T102|relax|30804-9|LNC|Chest vessels CT angiogram W WO contrast IV|Chest vessels CT angiogram W WO contrast IV
C0801762|T102|relax|36420-8|LNC|Chest vessels MRI angiogram W WO contrast IV|Chest vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|42277-4|LNC|Chest Abdomen CT W WO contrast IV|Chest Abdomen CT W WO contrast IV
C0801762|T102|relax|36284-8|LNC|Chest Abdomen MRI W WO contrast IV|Chest Abdomen MRI W WO contrast IV
C0801762|T102|relax|72252-0|LNC|Chest Abdomen Pelvis CT W WO contrast IV|Chest Abdomen Pelvis CT W WO contrast IV
C0801762|T102|relax|69161-8|LNC|Circle Willis MRI angiogram W WO contrast IV|Circle Willis MRI angiogram W WO contrast IV
C0801762|T102|relax|42299-8|LNC|Clavicle MRI W WO contrast IV|Clavicle MRI W WO contrast IV
C0801762|T102|relax|48455-0|LNC|Clavicle left MRI W WO contrast IV|Clavicle left MRI W WO contrast IV
C0801762|T102|relax|48454-3|LNC|Clavicle right MRI W WO contrast IV|Clavicle right MRI W WO contrast IV
C0801762|T102|relax|36285-5|LNC|Elbow CT W WO contrast IV|Elbow CT W WO contrast IV
C0801762|T102|relax|24675-1|LNC|Elbow MRI W WO contrast IV|Elbow MRI W WO contrast IV
C0801762|T102|relax|26193-3|LNC|Elbow bilateral MRI W WO contrast IV|Elbow bilateral MRI W WO contrast IV
C0801762|T102|relax|36286-3|LNC|Elbow left CT W WO contrast IV|Elbow left CT W WO contrast IV
C0801762|T102|relax|26194-1|LNC|Elbow left MRI W WO contrast IV|Elbow left MRI W WO contrast IV
C0801762|T102|relax|36287-1|LNC|Elbow right CT W WO contrast IV|Elbow right CT W WO contrast IV
C0801762|T102|relax|26195-8|LNC|Elbow right MRI W WO contrast IV|Elbow right MRI W WO contrast IV
C0801762|T102|relax|42268-3|LNC|Extremity CT W WO contrast IV|Extremity CT W WO contrast IV
C0801762|T102|relax|24694-2|LNC|Face MRI W WO contrast IV|Face MRI W WO contrast IV
C0801762|T102|relax|30803-1|LNC|Facial bones Maxilla CT W WO contrast IV|Facial bones Maxilla CT W WO contrast IV
C0801762|T102|relax|36338-2|LNC|Femur CT W WO contrast IV|Femur CT W WO contrast IV
C0801762|T102|relax|36339-0|LNC|Femur left CT W WO contrast IV|Femur left CT W WO contrast IV
C0801762|T102|relax|36340-8|LNC|Femur right CT W WO contrast IV|Femur right CT W WO contrast IV
C0801762|T102|relax|69194-9|LNC|Finger MRI W WO contrast IV|Finger MRI W WO contrast IV
C0801762|T102|relax|69204-6|LNC|Finger left MRI W WO contrast IV|Finger left MRI W WO contrast IV
C0801762|T102|relax|69214-5|LNC|Finger right MRI W WO contrast IV|Finger right MRI W WO contrast IV
C0801762|T102|relax|36341-6|LNC|Foot CT W WO contrast IV|Foot CT W WO contrast IV
C0801762|T102|relax|30682-9|LNC|Foot MRI W WO contrast IV|Foot MRI W WO contrast IV
C0801762|T102|relax|36342-4|LNC|Foot bilateral MRI W WO contrast IV|Foot bilateral MRI W WO contrast IV
C0801762|T102|relax|36343-2|LNC|Foot left CT W WO contrast IV|Foot left CT W WO contrast IV
C0801762|T102|relax|36344-0|LNC|Foot left MRI W WO contrast IV|Foot left MRI W WO contrast IV
C0801762|T102|relax|36345-7|LNC|Foot right CT W WO contrast IV|Foot right CT W WO contrast IV
C0801762|T102|relax|36346-5|LNC|Foot right MRI W WO contrast IV|Foot right MRI W WO contrast IV
C0801762|T102|relax|36347-3|LNC|Forearm CT W WO contrast IV|Forearm CT W WO contrast IV
C0801762|T102|relax|30684-5|LNC|Forearm MRI W WO contrast IV|Forearm MRI W WO contrast IV
C0801762|T102|relax|69174-1|LNC|Forearm bilateral MRI W WO contrast IV|Forearm bilateral MRI W WO contrast IV
C0801762|T102|relax|36348-1|LNC|Forearm left CT W WO contrast IV|Forearm left CT W WO contrast IV
C0801762|T102|relax|36349-9|LNC|Forearm left MRI W WO contrast IV|Forearm left MRI W WO contrast IV
C0801762|T102|relax|36350-7|LNC|Forearm right CT W WO contrast IV|Forearm right CT W WO contrast IV
C0801762|T102|relax|36351-5|LNC|Forearm right MRI W WO contrast IV|Forearm right MRI W WO contrast IV
C0801762|T102|relax|36352-3|LNC|Hand CT W WO contrast IV|Hand CT W WO contrast IV
C0801762|T102|relax|30686-0|LNC|Hand MRI W WO contrast IV|Hand MRI W WO contrast IV
C0801762|T102|relax|69177-4|LNC|Hand bilateral MRI W WO contrast IV|Hand bilateral MRI W WO contrast IV
C0801762|T102|relax|36353-1|LNC|Hand left CT W WO contrast IV|Hand left CT W WO contrast IV
C0801762|T102|relax|36354-9|LNC|Hand left MRI W WO contrast IV|Hand left MRI W WO contrast IV
C0801762|T102|relax|36355-6|LNC|Hand right CT W WO contrast IV|Hand right CT W WO contrast IV
C0801762|T102|relax|36356-4|LNC|Hand right MRI W WO contrast IV|Hand right MRI W WO contrast IV
C0801762|T102|relax|24726-2|LNC|Head CT W WO contrast IV|Head CT W WO contrast IV
C0801762|T102|relax|24729-6|LNC|Head CT cine W WO contrast IV|Head CT cine W WO contrast IV
C0801762|T102|relax|36847-2|LNC|Head veins MRI angiogram W WO contrast IV|Head veins MRI angiogram W WO contrast IV
C0801762|T102|relax|30593-8|LNC|Head vessels CT angiogram W WO contrast IV|Head vessels CT angiogram W WO contrast IV
C0801762|T102|relax|36857-1|LNC|Head vessels MRI angiogram W WO contrast IV|Head vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|36357-2|LNC|Heart MRI W WO contrast IV|Heart MRI W WO contrast IV
C0801762|T102|relax|36359-8|LNC|Hip CT W WO contrast IV|Hip CT W WO contrast IV
C0801762|T102|relax|30688-6|LNC|Hip MRI W WO contrast IV|Hip MRI W WO contrast IV
C0801762|T102|relax|36360-6|LNC|Hip bilateral CT W WO contrast IV|Hip bilateral CT W WO contrast IV
C0801762|T102|relax|36361-4|LNC|Hip bilateral MRI W WO contrast IV|Hip bilateral MRI W WO contrast IV
C0801762|T102|relax|36362-2|LNC|Hip left CT W WO contrast IV|Hip left CT W WO contrast IV
C0801762|T102|relax|36363-0|LNC|Hip left MRI W WO contrast IV|Hip left MRI W WO contrast IV
C0801762|T102|relax|36364-8|LNC|Hip right CT W WO contrast IV|Hip right CT W WO contrast IV
C0801762|T102|relax|36365-5|LNC|Hip right MRI W WO contrast IV|Hip right MRI W WO contrast IV
C0801762|T102|relax|36282-2|LNC|Internal auditory canal CT W WO contrast IV|Internal auditory canal CT W WO contrast IV
C0801762|T102|relax|30659-7|LNC|Internal auditory canal MRI W WO contrast IV|Internal auditory canal MRI W WO contrast IV
C0801762|T102|relax|24740-3|LNC|Internal auditory canal Posterior fossa MRI W WO contrast IV|Internal auditory canal Posterior fossa MRI W WO contrast IV
C0801762|T102|relax|43768-1|LNC|Kidney CT W WO contrast IV|Kidney CT W WO contrast IV
C0801762|T102|relax|43775-6|LNC|Kidney MRI W WO contrast IV|Kidney MRI W WO contrast IV
C0801762|T102|relax|36377-0|LNC|Kidney bilateral CT W WO contrast IV|Kidney bilateral CT W WO contrast IV
C0801762|T102|relax|36378-8|LNC|Kidney bilateral MRI W WO contrast IV|Kidney bilateral MRI W WO contrast IV
C0801762|T102|relax|24784-1|LNC|Kidney bilateral X-ray tomograph W WO contrast IV|Kidney bilateral X-ray tomograph W WO contrast IV
C0801762|T102|relax|36379-6|LNC|Knee CT W WO contrast IV|Knee CT W WO contrast IV
C0801762|T102|relax|24803-9|LNC|Knee MRI W WO contrast IV|Knee MRI W WO contrast IV
C0801762|T102|relax|38837-1|LNC|Knee vessels left MRI angiogram W WO contrast IV|Knee vessels left MRI angiogram W WO contrast IV
C0801762|T102|relax|36862-1|LNC|Knee vessels right MRI angiogram W WO contrast IV|Knee vessels right MRI angiogram W WO contrast IV
C0801762|T102|relax|26199-0|LNC|Knee bilateral MRI W WO contrast IV|Knee bilateral MRI W WO contrast IV
C0801762|T102|relax|36380-4|LNC|Knee left CT W WO contrast IV|Knee left CT W WO contrast IV
C0801762|T102|relax|26200-6|LNC|Knee left MRI W WO contrast IV|Knee left MRI W WO contrast IV
C0801762|T102|relax|36381-2|LNC|Knee right CT W WO contrast IV|Knee right CT W WO contrast IV
C0801762|T102|relax|26201-4|LNC|Knee right MRI W WO contrast IV|Knee right MRI W WO contrast IV
C0801762|T102|relax|36382-0|LNC|Larynx MRI W WO contrast IV|Larynx MRI W WO contrast IV
C0801762|T102|relax|30612-6|LNC|Liver CT W WO contrast IV|Liver CT W WO contrast IV
C0801762|T102|relax|30670-4|LNC|Liver MRI W WO contrast IV|Liver MRI W WO contrast IV
C0801762|T102|relax|36288-9|LNC|Lower extremity CT W WO contrast IV|Lower extremity CT W WO contrast IV
C0801762|T102|relax|39291-0|LNC|Lower extremity MRI W WO contrast IV|Lower extremity MRI W WO contrast IV
C0801762|T102|relax|36416-6|LNC|Lower extremity veins MRI angiogram W WO contrast IV|Lower extremity veins MRI angiogram W WO contrast IV
C0801762|T102|relax|36849-8|LNC|Lower extremity veins left MRI angiogram W WO contrast IV|Lower extremity veins left MRI angiogram W WO contrast IV
C0801762|T102|relax|36850-6|LNC|Lower extremity veins right MRI angiogram W WO contrast IV|Lower extremity veins right MRI angiogram W WO contrast IV
C0801762|T102|relax|30807-2|LNC|Lower extremity vessels CT angiogram W WO contrast IV|Lower extremity vessels CT angiogram W WO contrast IV
C0801762|T102|relax|44128-7|LNC|Lower extremity vessels MRI angiogram W WO contrast IV|Lower extremity vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|46308-3|LNC|Lower extremity vessels left CT angiogram W WO contrast IV|Lower extremity vessels left CT angiogram W WO contrast IV
C0801762|T102|relax|36858-9|LNC|Lower extremity vessels left MRI angiogram W WO contrast IV|Lower extremity vessels left MRI angiogram W WO contrast IV
C0801762|T102|relax|46307-5|LNC|Lower extremity vessels right CT angiogram W WO contrast IV|Lower extremity vessels right CT angiogram W WO contrast IV
C0801762|T102|relax|36859-7|LNC|Lower extremity vessels right MRI angiogram W WO contrast IV|Lower extremity vessels right MRI angiogram W WO contrast IV
C0801762|T102|relax|36289-7|LNC|Lower extremity bilateral MRI W WO contrast IV|Lower extremity bilateral MRI W WO contrast IV
C0801762|T102|relax|36371-3|LNC|Lower Extremity Joint MRI W WO contrast IV|Lower Extremity Joint MRI W WO contrast IV
C0801762|T102|relax|36372-1|LNC|Lower extremity joint left MRI W WO contrast IV|Lower extremity joint left MRI W WO contrast IV
C0801762|T102|relax|36373-9|LNC|Lower extremity joint right MRI W WO contrast IV|Lower extremity joint right MRI W WO contrast IV
C0801762|T102|relax|36290-5|LNC|Lower extremity left CT W WO contrast IV|Lower extremity left CT W WO contrast IV
C0801762|T102|relax|36291-3|LNC|Lower extremity left MRI W WO contrast IV|Lower extremity left MRI W WO contrast IV
C0801762|T102|relax|36292-1|LNC|Lower extremity right CT W WO contrast IV|Lower extremity right CT W WO contrast IV
C0801762|T102|relax|36333-3|LNC|Lower extremity right MRI W WO contrast IV|Lower extremity right MRI W WO contrast IV
C0801762|T102|relax|36408-3|LNC|Lower leg CT W WO contrast IV|Lower leg CT W WO contrast IV
C0801762|T102|relax|30870-0|LNC|Lower leg MRI W WO contrast IV|Lower leg MRI W WO contrast IV
C0801762|T102|relax|42697-3|LNC|Lower leg bilateral MRI W WO contrast IV|Lower leg bilateral MRI W WO contrast IV
C0801762|T102|relax|36409-1|LNC|Lower leg left CT W WO contrast IV|Lower leg left CT W WO contrast IV
C0801762|T102|relax|36410-9|LNC|Lower leg left MRI W WO contrast IV|Lower leg left MRI W WO contrast IV
C0801762|T102|relax|36411-7|LNC|Lower leg right CT W WO contrast IV|Lower leg right CT W WO contrast IV
C0801762|T102|relax|36412-5|LNC|Lower leg right MRI W WO contrast IV|Lower leg right MRI W WO contrast IV
C0801762|T102|relax|36383-8|LNC|Mandible CT W WO contrast IV|Mandible CT W WO contrast IV
C0801762|T102|relax|37272-2|LNC|Mediastinum MRI W WO contrast IV|Mediastinum MRI W WO contrast IV
C0801762|T102|relax|48443-6|LNC|Nasopharynx CT W WO contrast IV|Nasopharynx CT W WO contrast IV
C0801762|T102|relax|36384-6|LNC|Nasopharynx MRI W WO contrast IV|Nasopharynx MRI W WO contrast IV
C0801762|T102|relax|30586-2|LNC|Neck CT W WO contrast IV|Neck CT W WO contrast IV
C0801762|T102|relax|24840-1|LNC|Neck MRI W WO contrast IV|Neck MRI W WO contrast IV
C0801762|T102|relax|36853-0|LNC|Neck veins MRI angiogram W WO contrast IV|Neck veins MRI angiogram W WO contrast IV
C0801762|T102|relax|30594-6|LNC|Neck vessels CT angiogram W WO contrast IV|Neck vessels CT angiogram W WO contrast IV
C0801762|T102|relax|36423-2|LNC|Neck vessels MRI angiogram W WO contrast IV|Neck vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|48451-9|LNC|Orbit CT W WO contrast IV|Orbit CT W WO contrast IV
C0801762|T102|relax|36842-3|LNC|Orbit MRI W WO contrast IV|Orbit MRI W WO contrast IV
C0801762|T102|relax|43458-9|LNC|Orbit vessels MRI angiogram W WO contrast IV|Orbit vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|24849-2|LNC|Orbit bilateral CT W WO contrast IV|Orbit bilateral CT W WO contrast IV
C0801762|T102|relax|24851-8|LNC|Orbit bilateral MRI W WO contrast IV|Orbit bilateral MRI W WO contrast IV
C0801762|T102|relax|36843-1|LNC|Orbit left MRI W WO contrast IV|Orbit left MRI W WO contrast IV
C0801762|T102|relax|36844-9|LNC|Orbit right MRI W WO contrast IV|Orbit right MRI W WO contrast IV
C0801762|T102|relax|39029-4|LNC|Orbit Face MRI W WO contrast IV|Orbit Face MRI W WO contrast IV
C0801762|T102|relax|46310-9|LNC|Orbit Face Neck MRI W WO contrast IV|Orbit Face Neck MRI W WO contrast IV
C0801762|T102|relax|36845-6|LNC|Ovary MRI W WO contrast IV|Ovary MRI W WO contrast IV
C0801762|T102|relax|30614-2|LNC|Pancreas CT W WO contrast IV|Pancreas CT W WO contrast IV
C0801762|T102|relax|36385-3|LNC|Pancreas MRI W WO contrast IV|Pancreas MRI W WO contrast IV
C0801762|T102|relax|46311-7|LNC|Parotid gland CT W WO contrast IV|Parotid gland CT W WO contrast IV
C0801762|T102|relax|37265-6|LNC|Parotid gland MRI W WO contrast IV|Parotid gland MRI W WO contrast IV
C0801762|T102|relax|30616-7|LNC|Pelvis CT W WO contrast IV|Pelvis CT W WO contrast IV
C0801762|T102|relax|30674-6|LNC|Pelvis MRI W WO contrast IV|Pelvis MRI W WO contrast IV
C0801762|T102|relax|36854-8|LNC|Pelvis veins MRI angiogram W WO contrast IV|Pelvis veins MRI angiogram W WO contrast IV
C0801762|T102|relax|30623-3|LNC|Pelvis vessels CT angiogram W WO contrast IV|Pelvis vessels CT angiogram W WO contrast IV
C0801762|T102|relax|36863-9|LNC|Pelvis vessels MRI angiogram W WO contrast IV|Pelvis vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|30672-0|LNC|Pelvis Hip MRI W WO contrast IV|Pelvis Hip MRI W WO contrast IV
C0801762|T102|relax|36835-7|LNC|Petrous bone CT W WO contrast IV|Petrous bone CT W WO contrast IV
C0801762|T102|relax|24904-5|LNC|Pituitary Sella turcica CT W WO contrast IV|Pituitary Sella turcica CT W WO contrast IV
C0801762|T102|relax|24879-9|LNC|Pituitary Sella turcica MRI W WO contrast IV|Pituitary Sella turcica MRI W WO contrast IV
C0801762|T102|relax|36414-1|LNC|Portal vein MRI angiogram W WO contrast IV|Portal vein MRI angiogram W WO contrast IV
C0801762|T102|relax|36387-9|LNC|Posterior fossa CT W WO contrast IV|Posterior fossa CT W WO contrast IV
C0801762|T102|relax|36388-7|LNC|Posterior fossa MRI W WO contrast IV|Posterior fossa MRI W WO contrast IV
C0801762|T102|relax|36389-5|LNC|Prostate MRI W WO contrast IV|Prostate MRI W WO contrast IV
C0801762|T102|relax|36275-6|LNC|Renal artery MRI angiogram W WO contrast IV|Renal artery MRI angiogram W WO contrast IV
C0801762|T102|relax|36415-8|LNC|Renal vein MRI angiogram W WO contrast IV|Renal vein MRI angiogram W WO contrast IV
C0801762|T102|relax|44134-5|LNC|Renal vessels MRI angiogram W WO contrast IV|Renal vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|36375-4|LNC|Sacroiliac Joint CT W WO contrast IV|Sacroiliac Joint CT W WO contrast IV
C0801762|T102|relax|36376-2|LNC|Sacroiliac Joint MRI W WO contrast IV|Sacroiliac Joint MRI W WO contrast IV
C0801762|T102|relax|36390-3|LNC|Sacrum CT W WO contrast IV|Sacrum CT W WO contrast IV
C0801762|T102|relax|36391-1|LNC|Sacrum MRI W WO contrast IV|Sacrum MRI W WO contrast IV
C0801762|T102|relax|36392-9|LNC|Sacrum Coccyx MRI W WO contrast IV|Sacrum Coccyx MRI W WO contrast IV
C0801762|T102|relax|36393-7|LNC|Scapula left MRI W WO contrast IV|Scapula left MRI W WO contrast IV
C0801762|T102|relax|36394-5|LNC|Scapula right MRI W WO contrast IV|Scapula right MRI W WO contrast IV
C0801762|T102|relax|36406-7|LNC|Scrotum Testicle MRI W WO contrast IV|Scrotum Testicle MRI W WO contrast IV
C0801762|T102|relax|36395-2|LNC|Shoulder CT W WO contrast IV|Shoulder CT W WO contrast IV
C0801762|T102|relax|24906-0|LNC|Shoulder MRI W WO contrast IV|Shoulder MRI W WO contrast IV
C0801762|T102|relax|36864-7|LNC|Shoulder vessels left MRI angiogram W WO contrast IV|Shoulder vessels left MRI angiogram W WO contrast IV
C0801762|T102|relax|36865-4|LNC|Shoulder vessels right MRI angiogram W WO contrast IV|Shoulder vessels right MRI angiogram W WO contrast IV
C0801762|T102|relax|26202-2|LNC|Shoulder bilateral MRI W WO contrast IV|Shoulder bilateral MRI W WO contrast IV
C0801762|T102|relax|36396-0|LNC|Shoulder left CT W WO contrast IV|Shoulder left CT W WO contrast IV
C0801762|T102|relax|26203-0|LNC|Shoulder left MRI W WO contrast IV|Shoulder left MRI W WO contrast IV
C0801762|T102|relax|36397-8|LNC|Shoulder right CT W WO contrast IV|Shoulder right CT W WO contrast IV
C0801762|T102|relax|26204-8|LNC|Shoulder right MRI W WO contrast IV|Shoulder right MRI W WO contrast IV
C0801762|T102|relax|36398-6|LNC|Sinuses CT W WO contrast IV|Sinuses CT W WO contrast IV
C0801762|T102|relax|30663-9|LNC|Sinuses MRI W WO contrast IV|Sinuses MRI W WO contrast IV
C0801762|T102|relax|44111-3|LNC|Skull base CT W WO contrast IV|Skull base CT W WO contrast IV
C0801762|T102|relax|69220-2|LNC|Skull base MRI W WO contrast IV|Skull base MRI W WO contrast IV
C0801762|T102|relax|37277-1|LNC|Spinal vein MRI angiogram W WO contrast IV|Spinal vein MRI angiogram W WO contrast IV
C0801762|T102|relax|37505-5|LNC|Spine vessels MRI angiogram W WO contrast IV|Spine vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|36401-8|LNC|Spine Cervical CT W WO contrast IV|Spine Cervical CT W WO contrast IV
C0801762|T102|relax|24937-5|LNC|Spine Cervical MRI W WO contrast IV|Spine Cervical MRI W WO contrast IV
C0801762|T102|relax|37506-3|LNC|Cervical Spine vessels MRI angiogram W WO contrast IV|Cervical Spine vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|43456-3|LNC|Spine Cervical Spine Thoracic MRI W WO contrast IV|Spine Cervical Spine Thoracic MRI W WO contrast IV
C0801762|T102|relax|30855-1|LNC|Spine Cervical Thoracic Lumbar MRI W WO contrast IV|Spine Cervical Thoracic Lumbar MRI W WO contrast IV
C0801762|T102|relax|36402-6|LNC|Spine Lumbar CT W WO contrast IV|Spine Lumbar CT W WO contrast IV
C0801762|T102|relax|24967-2|LNC|Spine Lumbar MRI W WO contrast IV|Spine Lumbar MRI W WO contrast IV
C0801762|T102|relax|37507-1|LNC|Lumbar Spine vessels MRI angiogram W WO contrast IV|Lumbar Spine vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|36403-4|LNC|Spine Thoracic CT W WO contrast IV|Spine Thoracic CT W WO contrast IV
C0801762|T102|relax|24981-3|LNC|Spine Thoracic MRI W WO contrast IV|Spine Thoracic MRI W WO contrast IV
C0801762|T102|relax|37508-9|LNC|Thoracic Spine vessels MRI angiogram W WO contrast IV|Thoracic Spine vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|24989-6|LNC|Spleen CT W WO contrast IV|Spleen CT W WO contrast IV
C0801762|T102|relax|36404-2|LNC|Spleen MRI W WO contrast IV|Spleen MRI W WO contrast IV
C0801762|T102|relax|37266-4|LNC|Sternoclavicular Joint CT W WO contrast IV|Sternoclavicular Joint CT W WO contrast IV
C0801762|T102|relax|36405-9|LNC|Sternum CT W WO contrast IV|Sternum CT W WO contrast IV
C0801762|T102|relax|44231-9|LNC|Superior mesenteric vessels MRI angiogram W WO contrast IV|Superior mesenteric vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|36837-3|LNC|Temporal bone CT W WO contrast IV|Temporal bone CT W WO contrast IV
C0801762|T102|relax|37267-2|LNC|Temporomandibular joint CT W WO contrast IV|Temporomandibular joint CT W WO contrast IV
C0801762|T102|relax|37268-0|LNC|Temporomandibular joint MRI W WO contrast IV|Temporomandibular joint MRI W WO contrast IV
C0801762|T102|relax|37269-8|LNC|Temporomandibular joint bilateral MRI W WO contrast IV|Temporomandibular joint bilateral MRI W WO contrast IV
C0801762|T102|relax|37270-6|LNC|Temporomandibular joint left MRI W WO contrast IV|Temporomandibular joint left MRI W WO contrast IV
C0801762|T102|relax|37271-4|LNC|Temporomandibular joint right MRI W WO contrast IV|Temporomandibular joint right MRI W WO contrast IV
C0801762|T102|relax|24703-1|LNC|Thigh MRI W WO contrast IV|Thigh MRI W WO contrast IV
C0801762|T102|relax|26196-6|LNC|Thigh bilateral MRI W WO contrast IV|Thigh bilateral MRI W WO contrast IV
C0801762|T102|relax|26197-4|LNC|Thigh left MRI W WO contrast IV|Thigh left MRI W WO contrast IV
C0801762|T102|relax|26198-2|LNC|Thigh right MRI W WO contrast IV|Thigh right MRI W WO contrast IV
C0801762|T102|relax|24583-7|LNC|Thoracic outlet MRI W WO contrast IV|Thoracic outlet MRI W WO contrast IV
C0801762|T102|relax|26190-9|LNC|Thoracic outlet bilateral MRI W WO contrast IV|Thoracic outlet bilateral MRI W WO contrast IV
C0801762|T102|relax|26191-7|LNC|Thoracic outlet left MRI W WO contrast IV|Thoracic outlet left MRI W WO contrast IV
C0801762|T102|relax|26192-5|LNC|Thoracic outlet right MRI W WO contrast IV|Thoracic outlet right MRI W WO contrast IV
C0801762|T102|relax|36407-5|LNC|Thyroid MRI W WO contrast IV|Thyroid MRI W WO contrast IV
C0801762|T102|relax|72241-3|LNC|Toes left MRI W WO contrast IV|Toes left MRI W WO contrast IV
C0801762|T102|relax|72238-9|LNC|Toes right MRI W WO contrast IV|Toes right MRI W WO contrast IV
C0801762|T102|relax|36366-3|LNC|Upper arm CT W WO contrast IV|Upper arm CT W WO contrast IV
C0801762|T102|relax|30690-2|LNC|Upper arm MRI W WO contrast IV|Upper arm MRI W WO contrast IV
C0801762|T102|relax|69181-6|LNC|Upper arm bilateral MRI W WO contrast IV|Upper arm bilateral MRI W WO contrast IV
C0801762|T102|relax|36367-1|LNC|Upper arm left CT W WO contrast IV|Upper arm left CT W WO contrast IV
C0801762|T102|relax|36368-9|LNC|Upper arm left MRI W WO contrast IV|Upper arm left MRI W WO contrast IV
C0801762|T102|relax|36369-7|LNC|Upper arm right CT W WO contrast IV|Upper arm right CT W WO contrast IV
C0801762|T102|relax|36370-5|LNC|Upper arm right MRI W WO contrast IV|Upper arm right MRI W WO contrast IV
C0801762|T102|relax|36334-1|LNC|Upper extremity CT W WO contrast IV|Upper extremity CT W WO contrast IV
C0801762|T102|relax|39034-4|LNC|Upper extremity MRI W WO contrast IV|Upper extremity MRI W WO contrast IV
C0801762|T102|relax|36417-4|LNC|Upper extremity veins MRI angiogram W WO contrast IV|Upper extremity veins MRI angiogram W WO contrast IV
C0801762|T102|relax|36851-4|LNC|Upper extremity veins left MRI angiogram W WO contrast IV|Upper extremity veins left MRI angiogram W WO contrast IV
C0801762|T102|relax|36852-2|LNC|Upper extremity veins right MRI angiogram W WO contrast IV|Upper extremity veins right MRI angiogram W WO contrast IV
C0801762|T102|relax|36421-6|LNC|Upper extremity vessels CT angiogram W WO contrast IV|Upper extremity vessels CT angiogram W WO contrast IV
C0801762|T102|relax|36422-4|LNC|Upper extremity vessels MRI angiogram W WO contrast IV|Upper extremity vessels MRI angiogram W WO contrast IV
C0801762|T102|relax|46312-5|LNC|Upper extremity vessels left CT angiogram W WO contrast IV|Upper extremity vessels left CT angiogram W WO contrast IV
C0801762|T102|relax|36860-5|LNC|Upper extremity vessels left MRI angiogram W WO contrast IV|Upper extremity vessels left MRI angiogram W WO contrast IV
C0801762|T102|relax|46309-1|LNC|Upper extremity vessels right CT angiogram W WO contrast IV|Upper extremity vessels right CT angiogram W WO contrast IV
C0801762|T102|relax|36861-3|LNC|Upper extremity vessels right MRI angiogram W WO contrast IV|Upper extremity vessels right MRI angiogram W WO contrast IV
C0801762|T102|relax|69186-5|LNC|Upper extremity bilateral MRI W WO contrast IV|Upper extremity bilateral MRI W WO contrast IV
C0801762|T102|relax|36374-7|LNC|Upper extremity  joint MRI W WO contrast IV|Upper extremity  joint MRI W WO contrast IV
C0801762|T102|relax|36840-7|LNC|Upper extremity joint left MRI W WO contrast IV|Upper extremity joint left MRI W WO contrast IV
C0801762|T102|relax|36841-5|LNC|Upper extremity joint right MRI W WO contrast IV|Upper extremity joint right MRI W WO contrast IV
C0801762|T102|relax|36335-8|LNC|Upper extremity left CT W WO contrast IV|Upper extremity left CT W WO contrast IV
C0801762|T102|relax|38831-4|LNC|Upper extremity left MRI W WO contrast IV|Upper extremity left MRI W WO contrast IV
C0801762|T102|relax|36336-6|LNC|Upper extremity right CT W WO contrast IV|Upper extremity right CT W WO contrast IV
C0801762|T102|relax|36337-4|LNC|Upper extremity right MRI W WO contrast IV|Upper extremity right MRI W WO contrast IV
C0801762|T102|relax|36413-3|LNC|Uterus MRI W WO contrast IV|Uterus MRI W WO contrast IV
C0801762|T102|relax|36418-2|LNC|Inferior vena cava MRI W WO contrast IV|Inferior vena cava MRI W WO contrast IV
C0801762|T102|relax|36419-0|LNC|Superior vena cava MRI W WO contrast IV|Superior vena cava MRI W WO contrast IV
C0801762|T102|relax|37457-9|LNC|Wrist CT W WO contrast IV|Wrist CT W WO contrast IV
C0801762|T102|relax|25035-7|LNC|Wrist MRI W WO contrast IV|Wrist MRI W WO contrast IV
C0801762|T102|relax|26205-5|LNC|Wrist bilateral MRI W WO contrast IV|Wrist bilateral MRI W WO contrast IV
C0801762|T102|relax|37458-7|LNC|Wrist left CT W WO contrast IV|Wrist left CT W WO contrast IV
C0801762|T102|relax|26206-3|LNC|Wrist left MRI W WO contrast IV|Wrist left MRI W WO contrast IV
C0801762|T102|relax|38802-5|LNC|Wrist right CT W WO contrast IV|Wrist right CT W WO contrast IV
C0801762|T102|relax|26207-1|LNC|Wrist right MRI W WO contrast IV|Wrist right MRI W WO contrast IV
C0801762|T102|relax|42298-0|LNC|Unspecified body region MRI W WO contrast IV|Unspecified body region MRI W WO contrast IV
C0801762|T102|relax|24588-6|LNC|Brain MRI W WO contrast IV W anesthesia|Brain MRI W WO contrast IV W anesthesia
C0801762|T102|relax|72244-7|LNC|Pelvis MRI W WO contrast IV W endorectal coil|Pelvis MRI W WO contrast IV W endorectal coil
C0801762|T102|relax|43448-0|LNC|Liver MRI W WO ferumoxides IV|Liver MRI W WO ferumoxides IV
C0801762|T102|relax|46318-2|LNC|Abdomen CT W WO reduced contrast volume IV|Abdomen CT W WO reduced contrast volume IV
C0801762|T102|relax|46317-4|LNC|Chest CT W WO reduced contrast volume IV|Chest CT W WO reduced contrast volume IV
C0801762|T102|relax|46315-8|LNC|Facial bones Maxilla CT W WO reduced contrast volume IV|Facial bones Maxilla CT W WO reduced contrast volume IV
C0801762|T102|relax|46316-6|LNC|Head CT W WO reduced contrast volume IV|Head CT W WO reduced contrast volume IV
C0801762|T102|relax|46314-1|LNC|Internal auditory canal CT W WO reduced contrast volume IV|Internal auditory canal CT W WO reduced contrast volume IV
C0801762|T102|relax|46313-3|LNC|Pelvis CT W WO reduced contrast volume IV|Pelvis CT W WO reduced contrast volume IV
C0801762|T102|relax|60515-4|LNC|Rectum Colon CT 3D W air contrast PR|Rectum Colon CT 3D W air contrast PR
C0801762|T102|relax|24586-0|LNC|Brain MRI W anesthesia|Brain MRI W anesthesia
C0801762|T102|relax|24936-7|LNC|Spine Cervical MRI W anesthesia|Spine Cervical MRI W anesthesia
C0801762|T102|relax|24977-1|LNC|Spine Lumbar MRI W anesthesia|Spine Lumbar MRI W anesthesia
C0801762|T102|relax|25046-4|LNC|Unspecified body region CT W anesthesia|Unspecified body region CT W anesthesia
C0801762|T102|relax|38022-0|LNC|Gallbladder US W cholecystokinin|Gallbladder US W cholecystokinin
C0801762|T102|relax|25047-2|LNC|Unspecified body region CT W conscious sedation|Unspecified body region CT W conscious sedation
C0801762|T102|relax|25057-1|LNC|Unspecified body region MRI W conscious sedation|Unspecified body region MRI W conscious sedation
C0801762|T102|relax|30599-5|LNC|Abdomen CT W contrast|Abdomen CT W contrast
C0801762|T102|relax|24567-0|LNC|Abdomen retroperitoneum CT W contrast|Abdomen retroperitoneum CT W contrast
C0801762|T102|relax|38055-0|LNC|Unspecified body region US W contrast|Unspecified body region US W contrast
C0801762|T102|relax|36809-2|LNC|Hepatic artery CT angiogram W contrast IA|Hepatic artery CT angiogram W contrast IA
C0801762|T102|relax|69162-6|LNC|Pulmonary artery bilateral MRI angiogram W contrast IA|Pulmonary artery bilateral MRI angiogram W contrast IA
C0801762|T102|relax|69238-4|LNC|Urinary Bladder Urethra SPECT W contrast intra bladder during voiding|Urinary Bladder Urethra SPECT W contrast intra bladder during voiding
C0801762|T102|relax|30853-6|LNC|Breast duct US W contrast intra duct|Breast duct US W contrast intra duct
C0801762|T102|relax|36941-3|LNC|Salivary gland CT W contrast intra salivary duct|Salivary gland CT W contrast intra salivary duct
C0801762|T102|relax|37237-5|LNC|Sinus tract CT W contrast intra sinus tract|Sinus tract CT W contrast intra sinus tract
C0801762|T102|relax|36115-4|LNC|Ankle MRI W contrast intraarticular|Ankle MRI W contrast intraarticular
C0801762|T102|relax|69102-2|LNC|Ankle left CT W contrast intraarticular|Ankle left CT W contrast intraarticular
C0801762|T102|relax|36116-2|LNC|Ankle left MRI W contrast intraarticular|Ankle left MRI W contrast intraarticular
C0801762|T102|relax|69109-7|LNC|Ankle right CT W contrast intraarticular|Ankle right CT W contrast intraarticular
C0801762|T102|relax|36117-0|LNC|Ankle right MRI W contrast intraarticular|Ankle right MRI W contrast intraarticular
C0801762|T102|relax|46319-0|LNC|Elbow MRI W contrast intraarticular|Elbow MRI W contrast intraarticular
C0801762|T102|relax|69103-0|LNC|Elbow left CT W contrast intraarticular|Elbow left CT W contrast intraarticular
C0801762|T102|relax|36118-8|LNC|Elbow left MRI W contrast intraarticular|Elbow left MRI W contrast intraarticular
C0801762|T102|relax|69110-5|LNC|Elbow right CT W contrast intraarticular|Elbow right CT W contrast intraarticular
C0801762|T102|relax|36119-6|LNC|Elbow right MRI W contrast intraarticular|Elbow right MRI W contrast intraarticular
C0801762|T102|relax|36120-4|LNC|Hip MRI W contrast intraarticular|Hip MRI W contrast intraarticular
C0801762|T102|relax|69105-5|LNC|Hip left CT W contrast intraarticular|Hip left CT W contrast intraarticular
C0801762|T102|relax|36121-2|LNC|Hip left MRI W contrast intraarticular|Hip left MRI W contrast intraarticular
C0801762|T102|relax|69112-1|LNC|Hip right CT W contrast intraarticular|Hip right CT W contrast intraarticular
C0801762|T102|relax|36122-0|LNC|Hip right MRI W contrast intraarticular|Hip right MRI W contrast intraarticular
C0801762|T102|relax|36124-6|LNC|Knee CT W contrast intraarticular|Knee CT W contrast intraarticular
C0801762|T102|relax|36125-3|LNC|Knee MRI W contrast intraarticular|Knee MRI W contrast intraarticular
C0801762|T102|relax|69106-3|LNC|Knee left CT W contrast intraarticular|Knee left CT W contrast intraarticular
C0801762|T102|relax|36126-1|LNC|Knee left MRI W contrast intraarticular|Knee left MRI W contrast intraarticular
C0801762|T102|relax|69114-7|LNC|Knee right CT W contrast intraarticular|Knee right CT W contrast intraarticular
C0801762|T102|relax|36127-9|LNC|Knee right MRI W contrast intraarticular|Knee right MRI W contrast intraarticular
C0801762|T102|relax|37238-3|LNC|Lower Extremity Joint CT W contrast intraarticular|Lower Extremity Joint CT W contrast intraarticular
C0801762|T102|relax|69210-3|LNC|Lower Extremity Joint MRI W contrast intraarticular|Lower Extremity Joint MRI W contrast intraarticular
C0801762|T102|relax|36123-8|LNC|Sacroiliac Joint CT W contrast intraarticular|Sacroiliac Joint CT W contrast intraarticular
C0801762|T102|relax|36128-7|LNC|Shoulder CT W contrast intraarticular|Shoulder CT W contrast intraarticular
C0801762|T102|relax|36129-5|LNC|Shoulder MRI W contrast intraarticular|Shoulder MRI W contrast intraarticular
C0801762|T102|relax|38828-0|LNC|Shoulder left CT W contrast intraarticular|Shoulder left CT W contrast intraarticular
C0801762|T102|relax|36130-3|LNC|Shoulder left MRI W contrast intraarticular|Shoulder left MRI W contrast intraarticular
C0801762|T102|relax|36131-1|LNC|Shoulder right CT W contrast intraarticular|Shoulder right CT W contrast intraarticular
C0801762|T102|relax|36132-9|LNC|Shoulder right MRI W contrast intraarticular|Shoulder right MRI W contrast intraarticular
C0801762|T102|relax|36810-0|LNC|Upper Joint CT W contrast intraarticular|Upper Joint CT W contrast intraarticular
C0801762|T102|relax|37444-7|LNC|Wrist MRI W contrast intraarticular|Wrist MRI W contrast intraarticular
C0801762|T102|relax|69107-1|LNC|Wrist left CT W contrast intraarticular|Wrist left CT W contrast intraarticular
C0801762|T102|relax|37445-4|LNC|Wrist left MRI W contrast intraarticular|Wrist left MRI W contrast intraarticular
C0801762|T102|relax|69115-4|LNC|Wrist right CT W contrast intraarticular|Wrist right CT W contrast intraarticular
C0801762|T102|relax|37446-2|LNC|Wrist right MRI W contrast intraarticular|Wrist right MRI W contrast intraarticular
C0801762|T102|relax|36811-8|LNC|Joint CT W contrast intraarticular|Joint CT W contrast intraarticular
C0801762|T102|relax|36812-6|LNC|Joint MRI W contrast intraarticular|Joint MRI W contrast intraarticular
C0801762|T102|relax|37496-7|LNC|Spine Cervical CT W contrast intradisc|Spine Cervical CT W contrast intradisc
C0801762|T102|relax|37509-7|LNC|Spine Lumbar CT W contrast intradisc|Spine Lumbar CT W contrast intradisc
C0801762|T102|relax|70931-1|LNC|Spine Thoracic CT W contrast intradisc|Spine Thoracic CT W contrast intradisc
C0801762|T102|relax|24734-6|LNC|Head Cistern CT W contrast IT|Head Cistern CT W contrast IT
C0801762|T102|relax|24934-2|LNC|Spine Cervical CT W contrast IT|Spine Cervical CT W contrast IT
C0801762|T102|relax|48447-7|LNC|Spine Cervical MRI W contrast IT|Spine Cervical MRI W contrast IT
C0801762|T102|relax|24965-6|LNC|Spine Lumbar CT W contrast IT|Spine Lumbar CT W contrast IT
C0801762|T102|relax|48436-0|LNC|Spine Lumbar MRI W contrast IT|Spine Lumbar MRI W contrast IT
C0801762|T102|relax|30596-1|LNC|Spine Thoracic CT W contrast IT|Spine Thoracic CT W contrast IT
C0801762|T102|relax|48439-4|LNC|Spine Thoracic MRI W contrast IT|Spine Thoracic MRI W contrast IT
C0801762|T102|relax|36134-5|LNC|Abdomen MRI W contrast IV|Abdomen MRI W contrast IV
C0801762|T102|relax|36813-4|LNC|Abdomen Pelvis CT W contrast IV|Abdomen Pelvis CT W contrast IV
C0801762|T102|relax|36828-2|LNC|Abdominal vessels CT angiogram W contrast IV|Abdominal vessels CT angiogram W contrast IV
C0801762|T102|relax|24533-2|LNC|Abdominal vessels MRI angiogram W contrast IV|Abdominal vessels MRI angiogram W contrast IV
C0801762|T102|relax|69908-2|LNC|Abdominal vessels Pelvis vessels CT angiogram W contrast IV|Abdominal vessels Pelvis vessels CT angiogram W contrast IV
C0801762|T102|relax|36943-9|LNC|Adrenal gland CT W contrast IV|Adrenal gland CT W contrast IV
C0801762|T102|relax|44124-6|LNC|Adrenal gland MRI W contrast IV|Adrenal gland MRI W contrast IV
C0801762|T102|relax|36135-2|LNC|Ankle CT W contrast IV|Ankle CT W contrast IV
C0801762|T102|relax|36136-0|LNC|Ankle MRI W contrast IV|Ankle MRI W contrast IV
C0801762|T102|relax|69163-4|LNC|Ankle bilateral MRI W contrast IV|Ankle bilateral MRI W contrast IV
C0801762|T102|relax|36137-8|LNC|Ankle left CT W contrast IV|Ankle left CT W contrast IV
C0801762|T102|relax|36138-6|LNC|Ankle left MRI W contrast IV|Ankle left MRI W contrast IV
C0801762|T102|relax|36139-4|LNC|Ankle right CT W contrast IV|Ankle right CT W contrast IV
C0801762|T102|relax|36140-2|LNC|Ankle right MRI W contrast IV|Ankle right MRI W contrast IV
C0801762|T102|relax|36142-8|LNC|Aorta CT W contrast IV|Aorta CT W contrast IV
C0801762|T102|relax|36141-0|LNC|Aorta CT angiogram W contrast IV|Aorta CT angiogram W contrast IV
C0801762|T102|relax|36143-6|LNC|Aorta abdominal CT W contrast IV|Aorta abdominal CT W contrast IV
C0801762|T102|relax|24545-6|LNC|Aorta thoracic CT W contrast IV|Aorta thoracic CT W contrast IV
C0801762|T102|relax|72255-3|LNC|Aorta Femoral artery bilateral CT angiogram W contrast IV|Aorta Femoral artery bilateral CT angiogram W contrast IV
C0801762|T102|relax|43503-2|LNC|Aorta Lower extremity vessels CT angiogram W contrast IV|Aorta Lower extremity vessels CT angiogram W contrast IV
C0801762|T102|relax|36144-4|LNC|Aortic arch CT angiogram W contrast IV|Aortic arch CT angiogram W contrast IV
C0801762|T102|relax|37499-1|LNC|Aortic stent CT angiogram W contrast IV|Aortic stent CT angiogram W contrast IV
C0801762|T102|relax|36145-1|LNC|Appendix CT W contrast IV|Appendix CT W contrast IV
C0801762|T102|relax|43504-0|LNC|Axilla left MRI W contrast IV|Axilla left MRI W contrast IV
C0801762|T102|relax|43505-7|LNC|Axilla right MRI W contrast IV|Axilla right MRI W contrast IV
C0801762|T102|relax|44125-3|LNC|Biliary ducts Pancreatic duct MRI W contrast IV|Biliary ducts Pancreatic duct MRI W contrast IV
C0801762|T102|relax|69095-8|LNC|Bladder CT W contrast IV|Bladder CT W contrast IV
C0801762|T102|relax|24589-4|LNC|Brain MRI W contrast IV|Brain MRI W contrast IV
C0801762|T102|relax|48444-4|LNC|Brain temporal MRI W contrast IV|Brain temporal MRI W contrast IV
C0801762|T102|relax|37239-1|LNC|Brain Internal auditory canal MRI W contrast IV|Brain Internal auditory canal MRI W contrast IV
C0801762|T102|relax|37215-1|LNC|Brain Larynx MRI W contrast IV|Brain Larynx MRI W contrast IV
C0801762|T102|relax|42391-3|LNC|Brain Pituitary Sella turcica MRI W contrast IV|Brain Pituitary Sella turcica MRI W contrast IV
C0801762|T102|relax|36149-3|LNC|Breast MRI W contrast IV|Breast MRI W contrast IV
C0801762|T102|relax|69190-7|LNC|Breast implant MRI W contrast IV|Breast implant MRI W contrast IV
C0801762|T102|relax|69167-5|LNC|Breast implant bilateral MRI W contrast IV|Breast implant bilateral MRI W contrast IV
C0801762|T102|relax|36150-1|LNC|Breast bilateral MRI W contrast IV|Breast bilateral MRI W contrast IV
C0801762|T102|relax|36151-9|LNC|Breast left MRI W contrast IV|Breast left MRI W contrast IV
C0801762|T102|relax|36152-7|LNC|Breast right MRI W contrast IV|Breast right MRI W contrast IV
C0801762|T102|relax|46323-2|LNC|Breast unilateral MRI W contrast IV|Breast unilateral MRI W contrast IV
C0801762|T102|relax|36198-0|LNC|Calcaneus CT W contrast IV|Calcaneus CT W contrast IV
C0801762|T102|relax|36153-5|LNC|Calcaneus left CT W contrast IV|Calcaneus left CT W contrast IV
C0801762|T102|relax|36154-3|LNC|Calcaneus right CT W contrast IV|Calcaneus right CT W contrast IV
C0801762|T102|relax|36146-9|LNC|Carotid artery CT angiogram W contrast IV|Carotid artery CT angiogram W contrast IV
C0801762|T102|relax|36829-0|LNC|Carotid vessel MRI angiogram W contrast IV|Carotid vessel MRI angiogram W contrast IV
C0801762|T102|relax|24628-0|LNC|Chest CT W contrast IV|Chest CT W contrast IV
C0801762|T102|relax|36156-8|LNC|Chest MRI W contrast IV|Chest MRI W contrast IV
C0801762|T102|relax|36266-5|LNC|Chest vessels CT angiogram W contrast IV|Chest vessels CT angiogram W contrast IV
C0801762|T102|relax|24659-5|LNC|Chest vessels MRI angiogram W contrast IV|Chest vessels MRI angiogram W contrast IV
C0801762|T102|relax|42275-8|LNC|Chest Abdomen CT W contrast IV|Chest Abdomen CT W contrast IV
C0801762|T102|relax|36942-1|LNC|Chest Abdomen MRI W contrast IV|Chest Abdomen MRI W contrast IV
C0801762|T102|relax|72254-6|LNC|Chest Abdomen Pelvis CT W contrast IV|Chest Abdomen Pelvis CT W contrast IV
C0801762|T102|relax|37254-0|LNC|Circle Willis MRI angiogram W contrast IV|Circle Willis MRI angiogram W contrast IV
C0801762|T102|relax|42694-0|LNC|Clavicle MRI W contrast IV|Clavicle MRI W contrast IV
C0801762|T102|relax|48457-6|LNC|Clavicle left MRI W contrast IV|Clavicle left MRI W contrast IV
C0801762|T102|relax|48456-8|LNC|Clavicle right MRI W contrast IV|Clavicle right MRI W contrast IV
C0801762|T102|relax|36157-6|LNC|Elbow CT W contrast IV|Elbow CT W contrast IV
C0801762|T102|relax|36158-4|LNC|Elbow MRI W contrast IV|Elbow MRI W contrast IV
C0801762|T102|relax|69170-9|LNC|Elbow bilateral MRI W contrast IV|Elbow bilateral MRI W contrast IV
C0801762|T102|relax|36159-2|LNC|Elbow left CT W contrast IV|Elbow left CT W contrast IV
C0801762|T102|relax|36160-0|LNC|Elbow left MRI W contrast IV|Elbow left MRI W contrast IV
C0801762|T102|relax|36161-8|LNC|Elbow right CT W contrast IV|Elbow right CT W contrast IV
C0801762|T102|relax|36162-6|LNC|Elbow right MRI W contrast IV|Elbow right MRI W contrast IV
C0801762|T102|relax|24691-8|LNC|Extremity CT W contrast IV|Extremity CT W contrast IV
C0801762|T102|relax|26184-2|LNC|Extremity bilateral CT W contrast IV|Extremity bilateral CT W contrast IV
C0801762|T102|relax|26185-9|LNC|Extremity left CT W contrast IV|Extremity left CT W contrast IV
C0801762|T102|relax|26186-7|LNC|Extremity right CT W contrast IV|Extremity right CT W contrast IV
C0801762|T102|relax|36148-5|LNC|Face MRI W contrast IV|Face MRI W contrast IV
C0801762|T102|relax|30801-5|LNC|Facial bones Maxilla CT W contrast IV|Facial bones Maxilla CT W contrast IV
C0801762|T102|relax|24697-5|LNC|Facial bones Sinuses CT W contrast IV|Facial bones Sinuses CT W contrast IV
C0801762|T102|relax|36172-5|LNC|Femur CT W contrast IV|Femur CT W contrast IV
C0801762|T102|relax|69172-5|LNC|Femur bilateral MRI W contrast IV|Femur bilateral MRI W contrast IV
C0801762|T102|relax|36174-1|LNC|Femur left CT W contrast IV|Femur left CT W contrast IV
C0801762|T102|relax|36176-6|LNC|Femur right CT W contrast IV|Femur right CT W contrast IV
C0801762|T102|relax|69195-6|LNC|Finger MRI W contrast IV|Finger MRI W contrast IV
C0801762|T102|relax|69205-3|LNC|Finger left MRI W contrast IV|Finger left MRI W contrast IV
C0801762|T102|relax|69215-2|LNC|Finger right MRI W contrast IV|Finger right MRI W contrast IV
C0801762|T102|relax|36178-2|LNC|Foot CT W contrast IV|Foot CT W contrast IV
C0801762|T102|relax|36179-0|LNC|Foot MRI W contrast IV|Foot MRI W contrast IV
C0801762|T102|relax|36180-8|LNC|Foot bilateral MRI W contrast IV|Foot bilateral MRI W contrast IV
C0801762|T102|relax|36181-6|LNC|Foot left CT W contrast IV|Foot left CT W contrast IV
C0801762|T102|relax|36182-4|LNC|Foot left MRI W contrast IV|Foot left MRI W contrast IV
C0801762|T102|relax|36183-2|LNC|Foot right CT W contrast IV|Foot right CT W contrast IV
C0801762|T102|relax|36184-0|LNC|Foot right MRI W contrast IV|Foot right MRI W contrast IV
C0801762|T102|relax|36185-7|LNC|Forearm CT W contrast IV|Forearm CT W contrast IV
C0801762|T102|relax|36186-5|LNC|Forearm MRI W contrast IV|Forearm MRI W contrast IV
C0801762|T102|relax|69175-8|LNC|Forearm bilateral MRI W contrast IV|Forearm bilateral MRI W contrast IV
C0801762|T102|relax|36187-3|LNC|Forearm left CT W contrast IV|Forearm left CT W contrast IV
C0801762|T102|relax|36188-1|LNC|Forearm left MRI W contrast IV|Forearm left MRI W contrast IV
C0801762|T102|relax|36189-9|LNC|Forearm right CT W contrast IV|Forearm right CT W contrast IV
C0801762|T102|relax|36190-7|LNC|Forearm right MRI W contrast IV|Forearm right MRI W contrast IV
C0801762|T102|relax|36191-5|LNC|Hand CT W contrast IV|Hand CT W contrast IV
C0801762|T102|relax|36192-3|LNC|Hand MRI W contrast IV|Hand MRI W contrast IV
C0801762|T102|relax|69178-2|LNC|Hand bilateral MRI W contrast IV|Hand bilateral MRI W contrast IV
C0801762|T102|relax|36193-1|LNC|Hand left CT W contrast IV|Hand left CT W contrast IV
C0801762|T102|relax|36194-9|LNC|Hand left MRI W contrast IV|Hand left MRI W contrast IV
C0801762|T102|relax|36195-6|LNC|Hand right CT W contrast IV|Hand right CT W contrast IV
C0801762|T102|relax|36196-4|LNC|Hand right MRI W contrast IV|Hand right MRI W contrast IV
C0801762|T102|relax|24727-0|LNC|Head CT W contrast IV|Head CT W contrast IV
C0801762|T102|relax|36814-2|LNC|Head arteries CT angiogram W contrast IV|Head arteries CT angiogram W contrast IV
C0801762|T102|relax|36826-6|LNC|Head veins MRI angiogram W contrast IV|Head veins MRI angiogram W contrast IV
C0801762|T102|relax|36830-8|LNC|Head vessels CT angiogram W contrast IV|Head vessels CT angiogram W contrast IV
C0801762|T102|relax|24593-6|LNC|Head vessels MRI angiogram W contrast IV|Head vessels MRI angiogram W contrast IV
C0801762|T102|relax|37498-3|LNC|Head vessels Neck vessels CT angiogram W contrast IV|Head vessels Neck vessels CT angiogram W contrast IV
C0801762|T102|relax|24747-8|LNC|Head Sagittal Sinus MRI angiogram W contrast IV|Head Sagittal Sinus MRI angiogram W contrast IV
C0801762|T102|relax|36197-2|LNC|Heart MRI W contrast IV|Heart MRI W contrast IV
C0801762|T102|relax|36200-4|LNC|Hip CT W contrast IV|Hip CT W contrast IV
C0801762|T102|relax|36199-8|LNC|Hip MRI W contrast IV|Hip MRI W contrast IV
C0801762|T102|relax|36201-2|LNC|Hip bilateral CT W contrast IV|Hip bilateral CT W contrast IV
C0801762|T102|relax|36202-0|LNC|Hip bilateral MRI W contrast IV|Hip bilateral MRI W contrast IV
C0801762|T102|relax|36203-8|LNC|Hip left CT W contrast IV|Hip left CT W contrast IV
C0801762|T102|relax|36204-6|LNC|Hip left MRI W contrast IV|Hip left MRI W contrast IV
C0801762|T102|relax|36205-3|LNC|Hip right CT W contrast IV|Hip right CT W contrast IV
C0801762|T102|relax|36206-1|LNC|Hip right MRI W contrast IV|Hip right MRI W contrast IV
C0801762|T102|relax|30583-9|LNC|Internal auditory canal CT W contrast IV|Internal auditory canal CT W contrast IV
C0801762|T102|relax|36155-0|LNC|Internal auditory canal MRI W contrast IV|Internal auditory canal MRI W contrast IV
C0801762|T102|relax|46322-4|LNC|Kidney CT W contrast IV|Kidney CT W contrast IV
C0801762|T102|relax|36113-9|LNC|Kidney MRI W contrast IV|Kidney MRI W contrast IV
C0801762|T102|relax|43766-5|LNC|Kidney bilateral CT W contrast IV|Kidney bilateral CT W contrast IV
C0801762|T102|relax|36219-4|LNC|Kidney bilateral MRI W contrast IV|Kidney bilateral MRI W contrast IV
C0801762|T102|relax|24790-8|LNC|Kidney bilateral X-ray tomograph W contrast IV|Kidney bilateral X-ray tomograph W contrast IV
C0801762|T102|relax|36220-2|LNC|Kidney left MRI W contrast IV|Kidney left MRI W contrast IV
C0801762|T102|relax|36221-0|LNC|Kidney right MRI W contrast IV|Kidney right MRI W contrast IV
C0801762|T102|relax|36222-8|LNC|Knee CT W contrast IV|Knee CT W contrast IV
C0801762|T102|relax|36223-6|LNC|Knee MRI W contrast IV|Knee MRI W contrast IV
C0801762|T102|relax|69088-3|LNC|Knee bilateral CT W contrast IV|Knee bilateral CT W contrast IV
C0801762|T102|relax|36224-4|LNC|Knee bilateral MRI W contrast IV|Knee bilateral MRI W contrast IV
C0801762|T102|relax|36225-1|LNC|Knee left CT W contrast IV|Knee left CT W contrast IV
C0801762|T102|relax|36226-9|LNC|Knee left MRI W contrast IV|Knee left MRI W contrast IV
C0801762|T102|relax|36227-7|LNC|Knee right CT W contrast IV|Knee right CT W contrast IV
C0801762|T102|relax|36228-5|LNC|Knee right MRI W contrast IV|Knee right MRI W contrast IV
C0801762|T102|relax|36229-3|LNC|Larynx CT W contrast IV|Larynx CT W contrast IV
C0801762|T102|relax|36230-1|LNC|Larynx MRI W contrast IV|Larynx MRI W contrast IV
C0801762|T102|relax|24815-3|LNC|Liver CT W contrast IV|Liver CT W contrast IV
C0801762|T102|relax|36231-9|LNC|Liver MRI W contrast IV|Liver MRI W contrast IV
C0801762|T102|relax|30624-1|LNC|Lower extremity CT W contrast IV|Lower extremity CT W contrast IV
C0801762|T102|relax|39293-6|LNC|Lower extremity MRI W contrast IV|Lower extremity MRI W contrast IV
C0801762|T102|relax|36824-1|LNC|Lower extremity veins left CT W contrast IV|Lower extremity veins left CT W contrast IV
C0801762|T102|relax|36825-8|LNC|Lower extremity veins right CT W contrast IV|Lower extremity veins right CT W contrast IV
C0801762|T102|relax|36831-6|LNC|Lower extremity vessels CT angiogram W contrast IV|Lower extremity vessels CT angiogram W contrast IV
C0801762|T102|relax|46324-0|LNC|Lower extremity vessels MRI angiogram W contrast IV|Lower extremity vessels MRI angiogram W contrast IV
C0801762|T102|relax|44135-2|LNC|Lower extremity vessels bilateral MRI angiogram W contrast IV|Lower extremity vessels bilateral MRI angiogram W contrast IV
C0801762|T102|relax|50755-8|LNC|Lower extremity bilateral CT W contrast IV|Lower extremity bilateral CT W contrast IV
C0801762|T102|relax|36163-4|LNC|Lower extremity bilateral MRI W contrast IV|Lower extremity bilateral MRI W contrast IV
C0801762|T102|relax|36213-7|LNC|Lower Extremity Joint MRI W contrast IV|Lower Extremity Joint MRI W contrast IV
C0801762|T102|relax|36214-5|LNC|Lower extremity joint left MRI W contrast IV|Lower extremity joint left MRI W contrast IV
C0801762|T102|relax|36215-2|LNC|Lower extremity joint right MRI W contrast IV|Lower extremity joint right MRI W contrast IV
C0801762|T102|relax|36164-2|LNC|Lower extremity left CT W contrast IV|Lower extremity left CT W contrast IV
C0801762|T102|relax|36165-9|LNC|Lower extremity left MRI W contrast IV|Lower extremity left MRI W contrast IV
C0801762|T102|relax|36166-7|LNC|Lower extremity right CT W contrast IV|Lower extremity right CT W contrast IV
C0801762|T102|relax|36167-5|LNC|Lower extremity right MRI W contrast IV|Lower extremity right MRI W contrast IV
C0801762|T102|relax|36258-2|LNC|Lower leg CT W contrast IV|Lower leg CT W contrast IV
C0801762|T102|relax|36259-0|LNC|Lower leg MRI W contrast IV|Lower leg MRI W contrast IV
C0801762|T102|relax|24820-3|LNC|Lower leg vessels MRI angiogram W contrast IV|Lower leg vessels MRI angiogram W contrast IV
C0801762|T102|relax|43512-3|LNC|Lower leg vessels bilateral MRI angiogram W contrast IV|Lower leg vessels bilateral MRI angiogram W contrast IV
C0801762|T102|relax|42695-7|LNC|Lower leg bilateral MRI W contrast IV|Lower leg bilateral MRI W contrast IV
C0801762|T102|relax|36260-8|LNC|Lower leg left CT W contrast IV|Lower leg left CT W contrast IV
C0801762|T102|relax|36261-6|LNC|Lower leg left MRI W contrast IV|Lower leg left MRI W contrast IV
C0801762|T102|relax|36262-4|LNC|Lower leg right CT W contrast IV|Lower leg right CT W contrast IV
C0801762|T102|relax|36263-2|LNC|Lower leg right MRI W contrast IV|Lower leg right MRI W contrast IV
C0801762|T102|relax|36232-7|LNC|Mandible CT W contrast IV|Mandible CT W contrast IV
C0801762|T102|relax|48446-9|LNC|Nasopharynx CT W contrast IV|Nasopharynx CT W contrast IV
C0801762|T102|relax|36233-5|LNC|Nasopharynx MRI W contrast IV|Nasopharynx MRI W contrast IV
C0801762|T102|relax|24836-9|LNC|Nasopharynx Neck CT W contrast IV|Nasopharynx Neck CT W contrast IV
C0801762|T102|relax|36235-0|LNC|Neck CT W contrast IV|Neck CT W contrast IV
C0801762|T102|relax|24841-9|LNC|Neck MRI W contrast IV|Neck MRI W contrast IV
C0801762|T102|relax|36827-4|LNC|Neck veins MRI angiogram W contrast IV|Neck veins MRI angiogram W contrast IV
C0801762|T102|relax|36234-3|LNC|Neck vessels CT angiogram W contrast IV|Neck vessels CT angiogram W contrast IV
C0801762|T102|relax|24844-3|LNC|Neck vessels MRI angiogram W contrast IV|Neck vessels MRI angiogram W contrast IV
C0801762|T102|relax|48449-3|LNC|Orbit CT W contrast IV|Orbit CT W contrast IV
C0801762|T102|relax|36820-9|LNC|Orbit MRI W contrast IV|Orbit MRI W contrast IV
C0801762|T102|relax|36832-4|LNC|Orbit vessels MRI angiogram W contrast IV|Orbit vessels MRI angiogram W contrast IV
C0801762|T102|relax|24850-0|LNC|Orbit bilateral CT W contrast IV|Orbit bilateral CT W contrast IV
C0801762|T102|relax|24852-6|LNC|Orbit bilateral MRI W contrast IV|Orbit bilateral MRI W contrast IV
C0801762|T102|relax|36821-7|LNC|Orbit left MRI W contrast IV|Orbit left MRI W contrast IV
C0801762|T102|relax|36822-5|LNC|Orbit right MRI W contrast IV|Orbit right MRI W contrast IV
C0801762|T102|relax|46320-8|LNC|Orbit Face CT W contrast IV|Orbit Face CT W contrast IV
C0801762|T102|relax|39038-5|LNC|Orbit Face MRI W contrast IV|Orbit Face MRI W contrast IV
C0801762|T102|relax|46321-6|LNC|Orbit Face Neck MRI W contrast IV|Orbit Face Neck MRI W contrast IV
C0801762|T102|relax|36823-3|LNC|Ovary MRI W contrast IV|Ovary MRI W contrast IV
C0801762|T102|relax|24858-3|LNC|Pancreas CT W contrast IV|Pancreas CT W contrast IV
C0801762|T102|relax|36236-8|LNC|Pancreas MRI W contrast IV|Pancreas MRI W contrast IV
C0801762|T102|relax|37240-9|LNC|Parotid gland CT W contrast IV|Parotid gland CT W contrast IV
C0801762|T102|relax|37241-7|LNC|Parotid gland MRI W contrast IV|Parotid gland MRI W contrast IV
C0801762|T102|relax|24866-6|LNC|Pelvis CT W contrast IV|Pelvis CT W contrast IV
C0801762|T102|relax|36237-6|LNC|Pelvis MRI W contrast IV|Pelvis MRI W contrast IV
C0801762|T102|relax|42294-9|LNC|Pelvis vessels CT angiogram W contrast IV|Pelvis vessels CT angiogram W contrast IV
C0801762|T102|relax|24873-2|LNC|Pelvis vessels MRI angiogram W contrast IV|Pelvis vessels MRI angiogram W contrast IV
C0801762|T102|relax|24878-1|LNC|Petrous bone CT W contrast IV|Petrous bone CT W contrast IV
C0801762|T102|relax|30590-4|LNC|Pituitary Sella turcica CT W contrast IV|Pituitary Sella turcica CT W contrast IV
C0801762|T102|relax|36238-4|LNC|Pituitary Sella turcica MRI W contrast IV|Pituitary Sella turcica MRI W contrast IV
C0801762|T102|relax|36242-6|LNC|Posterior fossa CT W contrast IV|Posterior fossa CT W contrast IV
C0801762|T102|relax|36243-4|LNC|Posterior fossa MRI W contrast IV|Posterior fossa MRI W contrast IV
C0801762|T102|relax|36244-2|LNC|Prostate MRI W contrast IV|Prostate MRI W contrast IV
C0801762|T102|relax|36147-7|LNC|Pulmonary artery CT angiogram W contrast IV|Pulmonary artery CT angiogram W contrast IV
C0801762|T102|relax|36833-2|LNC|Renal vessels CT angiogram W contrast IV|Renal vessels CT angiogram W contrast IV
C0801762|T102|relax|30887-4|LNC|Renal vessels MRI angiogram W contrast IV|Renal vessels MRI angiogram W contrast IV
C0801762|T102|relax|36217-8|LNC|Sacroiliac Joint CT W contrast IV|Sacroiliac Joint CT W contrast IV
C0801762|T102|relax|36218-6|LNC|Sacroiliac Joint MRI W contrast IV|Sacroiliac Joint MRI W contrast IV
C0801762|T102|relax|36245-9|LNC|Sacrum CT W contrast IV|Sacrum CT W contrast IV
C0801762|T102|relax|36246-7|LNC|Sacrum MRI W contrast IV|Sacrum MRI W contrast IV
C0801762|T102|relax|36247-5|LNC|Sacrum Coccyx MRI W contrast IV|Sacrum Coccyx MRI W contrast IV
C0801762|T102|relax|36248-3|LNC|Scapula left MRI W contrast IV|Scapula left MRI W contrast IV
C0801762|T102|relax|36249-1|LNC|Scapula right MRI W contrast IV|Scapula right MRI W contrast IV
C0801762|T102|relax|69221-0|LNC|Scrotum Testicle MRI W contrast IV|Scrotum Testicle MRI W contrast IV
C0801762|T102|relax|36250-9|LNC|Shoulder CT W contrast IV|Shoulder CT W contrast IV
C0801762|T102|relax|36251-7|LNC|Shoulder MRI W contrast IV|Shoulder MRI W contrast IV
C0801762|T102|relax|69184-0|LNC|Shoulder bilateral MRI W contrast IV|Shoulder bilateral MRI W contrast IV
C0801762|T102|relax|36252-5|LNC|Shoulder left CT W contrast IV|Shoulder left CT W contrast IV
C0801762|T102|relax|38830-6|LNC|Shoulder left MRI W contrast IV|Shoulder left MRI W contrast IV
C0801762|T102|relax|36253-3|LNC|Shoulder right CT W contrast IV|Shoulder right CT W contrast IV
C0801762|T102|relax|36254-1|LNC|Shoulder right MRI W contrast IV|Shoulder right MRI W contrast IV
C0801762|T102|relax|36255-8|LNC|Sinuses CT W contrast IV|Sinuses CT W contrast IV
C0801762|T102|relax|24915-1|LNC|Sinuses MRI W contrast IV|Sinuses MRI W contrast IV
C0801762|T102|relax|48440-2|LNC|Skull base MRI W contrast IV|Skull base MRI W contrast IV
C0801762|T102|relax|37253-2|LNC|Soft tissue MRI W contrast IV|Soft tissue MRI W contrast IV
C0801762|T102|relax|37500-6|LNC|Spine vessels MRI angiogram W contrast IV|Spine vessels MRI angiogram W contrast IV
C0801762|T102|relax|24933-4|LNC|Spine Cervical CT W contrast IV|Spine Cervical CT W contrast IV
C0801762|T102|relax|24938-3|LNC|Spine Cervical MRI W contrast IV|Spine Cervical MRI W contrast IV
C0801762|T102|relax|37501-4|LNC|Cervical Spine vessels MRI angiogram W contrast IV|Cervical Spine vessels MRI angiogram W contrast IV
C0801762|T102|relax|38061-8|LNC|Spine Cervical Spine Thoracic Spine Lumbar Sacrum MRI W contrast IV|Spine Cervical Spine Thoracic Spine Lumbar Sacrum MRI W contrast IV
C0801762|T102|relax|24964-9|LNC|Spine Lumbar CT W contrast IV|Spine Lumbar CT W contrast IV
C0801762|T102|relax|30678-7|LNC|Spine Lumbar MRI W contrast IV|Spine Lumbar MRI W contrast IV
C0801762|T102|relax|37502-2|LNC|Lumbar Spine vessels MRI angiogram W contrast IV|Lumbar Spine vessels MRI angiogram W contrast IV
C0801762|T102|relax|24979-7|LNC|Spine Thoracic CT W contrast IV|Spine Thoracic CT W contrast IV
C0801762|T102|relax|24982-1|LNC|Spine Thoracic MRI W contrast IV|Spine Thoracic MRI W contrast IV
C0801762|T102|relax|37503-0|LNC|Thoracic Spine vessels MRI angiogram W contrast IV|Thoracic Spine vessels MRI angiogram W contrast IV
C0801762|T102|relax|30622-5|LNC|Spleen CT W contrast IV|Spleen CT W contrast IV
C0801762|T102|relax|37242-5|LNC|Sternoclavicular Joint CT W contrast IV|Sternoclavicular Joint CT W contrast IV
C0801762|T102|relax|36257-4|LNC|Sternum CT W contrast IV|Sternum CT W contrast IV
C0801762|T102|relax|36815-9|LNC|Temporal bone CT W contrast IV|Temporal bone CT W contrast IV
C0801762|T102|relax|38835-5|LNC|Temporal bone left CT W contrast IV|Temporal bone left CT W contrast IV
C0801762|T102|relax|36816-7|LNC|Temporal bone right CT W contrast IV|Temporal bone right CT W contrast IV
C0801762|T102|relax|37243-3|LNC|Temporomandibular joint CT W contrast IV|Temporomandibular joint CT W contrast IV
C0801762|T102|relax|37244-1|LNC|Temporomandibular joint MRI W contrast IV|Temporomandibular joint MRI W contrast IV
C0801762|T102|relax|37245-8|LNC|Temporomandibular joint bilateral MRI W contrast IV|Temporomandibular joint bilateral MRI W contrast IV
C0801762|T102|relax|37246-6|LNC|Temporomandibular joint left CT W contrast IV|Temporomandibular joint left CT W contrast IV
C0801762|T102|relax|37247-4|LNC|Temporomandibular joint left MRI W contrast IV|Temporomandibular joint left MRI W contrast IV
C0801762|T102|relax|37248-2|LNC|Temporomandibular joint right CT W contrast IV|Temporomandibular joint right CT W contrast IV
C0801762|T102|relax|37249-0|LNC|Temporomandibular joint right MRI W contrast IV|Temporomandibular joint right MRI W contrast IV
C0801762|T102|relax|36173-3|LNC|Thigh MRI W contrast IV|Thigh MRI W contrast IV
C0801762|T102|relax|25003-5|LNC|Thigh vessels MRI angiogram W contrast IV|Thigh vessels MRI angiogram W contrast IV
C0801762|T102|relax|36175-8|LNC|Thigh left MRI W contrast IV|Thigh left MRI W contrast IV
C0801762|T102|relax|36177-4|LNC|Thigh right MRI W contrast IV|Thigh right MRI W contrast IV
C0801762|T102|relax|36239-2|LNC|Thoracic outlet MRI W contrast IV|Thoracic outlet MRI W contrast IV
C0801762|T102|relax|24584-5|LNC|Thoracic outlet vessels MRI angiogram W contrast IV|Thoracic outlet vessels MRI angiogram W contrast IV
C0801762|T102|relax|26181-8|LNC|Thoracic outlet vessels bilateral MRI angiogram W contrast IV|Thoracic outlet vessels bilateral MRI angiogram W contrast IV
C0801762|T102|relax|26182-6|LNC|Thoracic outlet vessels left MRI angiogram W contrast IV|Thoracic outlet vessels left MRI angiogram W contrast IV
C0801762|T102|relax|26183-4|LNC|Thoracic outlet vessels right MRI angiogram W contrast IV|Thoracic outlet vessels right MRI angiogram W contrast IV
C0801762|T102|relax|36240-0|LNC|Thoracic outlet left MRI W contrast IV|Thoracic outlet left MRI W contrast IV
C0801762|T102|relax|36241-8|LNC|Thoracic outlet right MRI W contrast IV|Thoracic outlet right MRI W contrast IV
C0801762|T102|relax|72243-9|LNC|Toes left MRI W contrast IV|Toes left MRI W contrast IV
C0801762|T102|relax|72240-5|LNC|Toes right MRI W contrast IV|Toes right MRI W contrast IV
C0801762|T102|relax|36207-9|LNC|Upper arm CT W contrast IV|Upper arm CT W contrast IV
C0801762|T102|relax|36208-7|LNC|Upper arm MRI W contrast IV|Upper arm MRI W contrast IV
C0801762|T102|relax|69182-4|LNC|Upper arm bilateral MRI W contrast IV|Upper arm bilateral MRI W contrast IV
C0801762|T102|relax|36209-5|LNC|Upper arm left CT W contrast IV|Upper arm left CT W contrast IV
C0801762|T102|relax|36210-3|LNC|Upper arm left MRI W contrast IV|Upper arm left MRI W contrast IV
C0801762|T102|relax|36211-1|LNC|Upper arm right CT W contrast IV|Upper arm right CT W contrast IV
C0801762|T102|relax|36212-9|LNC|Upper arm right MRI W contrast IV|Upper arm right MRI W contrast IV
C0801762|T102|relax|30626-6|LNC|Upper extremity CT W contrast IV|Upper extremity CT W contrast IV
C0801762|T102|relax|39037-7|LNC|Upper extremity MRI W contrast IV|Upper extremity MRI W contrast IV
C0801762|T102|relax|42295-6|LNC|Upper extremity vessels CT angiogram W contrast IV|Upper extremity vessels CT angiogram W contrast IV
C0801762|T102|relax|24549-8|LNC|Upper extremity vessels MRI angiogram W contrast IV|Upper extremity vessels MRI angiogram W contrast IV
C0801762|T102|relax|36168-3|LNC|Upper extremity bilateral CT W contrast IV|Upper extremity bilateral CT W contrast IV
C0801762|T102|relax|69187-3|LNC|Upper extremity bilateral MRI W contrast IV|Upper extremity bilateral MRI W contrast IV
C0801762|T102|relax|36216-0|LNC|Upper extremity  joint MRI W contrast IV|Upper extremity  joint MRI W contrast IV
C0801762|T102|relax|36817-5|LNC|Upper extremity joint bilateral MRI W contrast IV|Upper extremity joint bilateral MRI W contrast IV
C0801762|T102|relax|36818-3|LNC|Upper extremity joint left MRI W contrast IV|Upper extremity joint left MRI W contrast IV
C0801762|T102|relax|36819-1|LNC|Upper extremity joint right MRI W contrast IV|Upper extremity joint right MRI W contrast IV
C0801762|T102|relax|36169-1|LNC|Upper extremity left CT W contrast IV|Upper extremity left CT W contrast IV
C0801762|T102|relax|38829-8|LNC|Upper extremity left MRI W contrast IV|Upper extremity left MRI W contrast IV
C0801762|T102|relax|36170-9|LNC|Upper extremity right CT W contrast IV|Upper extremity right CT W contrast IV
C0801762|T102|relax|36171-7|LNC|Upper extremity right MRI W contrast IV|Upper extremity right MRI W contrast IV
C0801762|T102|relax|36264-0|LNC|Uterus CT W contrast IV|Uterus CT W contrast IV
C0801762|T102|relax|36265-7|LNC|Uterus MRI W contrast IV|Uterus MRI W contrast IV
C0801762|T102|relax|36834-0|LNC|Vessel CT angiogram W contrast IV|Vessel CT angiogram W contrast IV
C0801762|T102|relax|37447-0|LNC|Wrist CT W contrast IV|Wrist CT W contrast IV
C0801762|T102|relax|37448-8|LNC|Wrist MRI W contrast IV|Wrist MRI W contrast IV
C0801762|T102|relax|69091-7|LNC|Wrist bilateral CT W contrast IV|Wrist bilateral CT W contrast IV
C0801762|T102|relax|37449-6|LNC|Wrist bilateral MRI W contrast IV|Wrist bilateral MRI W contrast IV
C0801762|T102|relax|37450-4|LNC|Wrist left CT W contrast IV|Wrist left CT W contrast IV
C0801762|T102|relax|37451-2|LNC|Wrist left MRI W contrast IV|Wrist left MRI W contrast IV
C0801762|T102|relax|37452-0|LNC|Wrist right CT W contrast IV|Wrist right CT W contrast IV
C0801762|T102|relax|37453-8|LNC|Wrist right MRI W contrast IV|Wrist right MRI W contrast IV
C0801762|T102|relax|24753-6|LNC|Unspecified body region CT W contrast IV|Unspecified body region CT W contrast IV
C0801762|T102|relax|49507-7|LNC|Unspecified body region MRI W contrast IV|Unspecified body region MRI W contrast IV
C0801762|T102|relax|25058-9|LNC|Unspecified body region MRI angiogram W contrast IV|Unspecified body region MRI angiogram W contrast IV
C0801762|T102|relax|72531-7|LNC|Rectum Colon CT 3D W contrast IV W air contrast PR|Rectum Colon CT 3D W contrast IV W air contrast PR
C0801762|T102|relax|39450-2|LNC|Gastrointestine US W contrast PO|Gastrointestine US W contrast PO
C0801762|T102|relax|72246-2|LNC|Abdomen Pelvis MRI W contrast PO W WO contrast IV|Abdomen Pelvis MRI W contrast PO W WO contrast IV
C0801762|T102|relax|72250-4|LNC|Abdomen Pelvis CT W contrast PO W contrast IV|Abdomen Pelvis CT W contrast PO W contrast IV
C0801762|T102|relax|72247-0|LNC|Abdomen Pelvis MRI W contrast PO WO contrast IV|Abdomen Pelvis MRI W contrast PO WO contrast IV
C0801762|T102|relax|72245-4|LNC|Pelvis MRI W contrast PR at rest maxmal sphincter contraction during straining defecation|Pelvis MRI W contrast PR at rest maxmal sphincter contraction during straining defecation
C0801762|T102|relax|39648-1|LNC|Heart SPECT W dipyridamole W radionuclide IV|Heart SPECT W dipyridamole W radionuclide IV
C0801762|T102|relax|44154-3|LNC|Heart SPECT W dipyridamole W Tc-99m Sestamibi IV|Heart SPECT W dipyridamole W Tc-99m Sestamibi IV
C0801762|T102|relax|42389-7|LNC|Pelvis MRI W endorectal coil|Pelvis MRI W endorectal coil
C0801762|T102|relax|42388-9|LNC|Prostate MRI W endorectal coil|Prostate MRI W endorectal coil
C0801762|T102|relax|42270-9|LNC|Spine Cervical MRI W flexion W extension|Spine Cervical MRI W flexion W extension
C0801762|T102|relax|39682-0|LNC|SPECT W GA-67 IV|SPECT W GA-67 IV
C0801762|T102|relax|39638-2|LNC|Brain SPECT W I-123 IV|Brain SPECT W I-123 IV
C0801762|T102|relax|39755-4|LNC|Thyroid SPECT W I-131 IV|Thyroid SPECT W I-131 IV
C0801762|T102|relax|39839-6|LNC|SPECT W I-131 MIBG IV|SPECT W I-131 MIBG IV
C0801762|T102|relax|39844-6|LNC|SPECT W In-111 Satumomab IV|SPECT W In-111 Satumomab IV
C0801762|T102|relax|41838-4|LNC|Prostate SPECT W In-111 Satumomab IV|Prostate SPECT W In-111 Satumomab IV
C0801762|T102|relax|41772-5|LNC|Bone SPECT W In-111 tagged WBC IV|Bone SPECT W In-111 tagged WBC IV
C0801762|T102|relax|46297-8|LNC|SPECT|SPECT
C0801762|T102|relax|39823-0|LNC|Bone marrow SPECT|Bone marrow SPECT
C0801762|T102|relax|24578-7|LNC|Bones SPECT|Bones SPECT
C0801762|T102|relax|39632-5|LNC|Brain SPECT|Brain SPECT
C0801762|T102|relax|39644-0|LNC|Breast SPECT|Breast SPECT
C0801762|T102|relax|39770-3|LNC|Gastrointestine SPECT|Gastrointestine SPECT
C0801762|T102|relax|39649-9|LNC|Heart SPECT|Heart SPECT
C0801762|T102|relax|42310-3|LNC|Kidney SPECT|Kidney SPECT
C0801762|T102|relax|39852-9|LNC|Kidney bilateral SPECT|Kidney bilateral SPECT
C0801762|T102|relax|39692-9|LNC|Liver SPECT|Liver SPECT
C0801762|T102|relax|39876-8|LNC|Liver Spleen SPECT|Liver Spleen SPECT
C0801762|T102|relax|39628-3|LNC|Meckels diverticulum SPECT|Meckels diverticulum SPECT
C0801762|T102|relax|39740-6|LNC|Parathyroid SPECT|Parathyroid SPECT
C0801762|T102|relax|43526-3|LNC|Unspecified body region SPECT|Unspecified body region SPECT
C0801762|T102|relax|39938-6|LNC|Joint SPECT|Joint SPECT
C0801762|T102|relax|46330-7|LNC|Abdomen CT W reduced contrast volume IV|Abdomen CT W reduced contrast volume IV
C0801762|T102|relax|46327-3|LNC|Chest CT W reduced contrast volume IV|Chest CT W reduced contrast volume IV
C0801762|T102|relax|46326-5|LNC|Facial bones Maxilla CT W reduced contrast volume IV|Facial bones Maxilla CT W reduced contrast volume IV
C0801762|T102|relax|46328-1|LNC|Head CT W reduced contrast volume IV|Head CT W reduced contrast volume IV
C0801762|T102|relax|46325-7|LNC|Internal auditory canal CT W reduced contrast volume IV|Internal auditory canal CT W reduced contrast volume IV
C0801762|T102|relax|46329-9|LNC|Pelvis CT W reduced contrast volume IV|Pelvis CT W reduced contrast volume IV
C0801762|T102|relax|42143-8|LNC|Uterus Fallopian tubes US W saline intrauterine|Uterus Fallopian tubes US W saline intrauterine
C0801762|T102|relax|58750-1|LNC|Heart MRI W stress|Heart MRI W stress
C0801762|T102|relax|58749-3|LNC|Heart MRI W stress W WO contrast IV|Heart MRI W stress W WO contrast IV
C0801762|T102|relax|39668-9|LNC|Heart SPECT W stress W radionuclide IV|Heart SPECT W stress W radionuclide IV
C0801762|T102|relax|44152-7|LNC|Brain SPECT W Tc-99m bicisate IV|Brain SPECT W Tc-99m bicisate IV
C0801762|T102|relax|39743-0|LNC|Prostate SPECT W Tc-99m capromab pendatide IV|Prostate SPECT W Tc-99m capromab pendatide IV
C0801762|T102|relax|39640-8|LNC|Brain SPECT W Tc-99m DTPA IV|Brain SPECT W Tc-99m DTPA IV
C0801762|T102|relax|39641-6|LNC|Brain SPECT W Tc-99m glucoheptonate IV|Brain SPECT W Tc-99m glucoheptonate IV
C0801762|T102|relax|44153-5|LNC|Kidney SPECT W Tc-99m glucoheptonate IV|Kidney SPECT W Tc-99m glucoheptonate IV
C0801762|T102|relax|39631-7|LNC|Brain SPECT W Tc-99m HMPAO IV|Brain SPECT W Tc-99m HMPAO IV
C0801762|T102|relax|24817-9|LNC|Liver SPECT W Tc-99m IV|Liver SPECT W Tc-99m IV
C0801762|T102|relax|39851-1|LNC|Kidney bilateral SPECT W Tc-99m Mertiatide IV|Kidney bilateral SPECT W Tc-99m Mertiatide IV
C0801762|T102|relax|69229-3|LNC|Liver SPECT W Tc-99m SC IV|Liver SPECT W Tc-99m SC IV
C0801762|T102|relax|44151-9|LNC|Heart SPECT W Tc-99m Sestamibi IV|Heart SPECT W Tc-99m Sestamibi IV
C0801762|T102|relax|39691-1|LNC|Liver SPECT W Tc-99m tagged RBC IV|Liver SPECT W Tc-99m tagged RBC IV
C0801762|T102|relax|69234-3|LNC|Spleen SPECT W Tc-99m tagged RBC IV|Spleen SPECT W Tc-99m tagged RBC IV
C0801762|T102|relax|39647-3|LNC|Heart SPECT W Tc-99m Tetrofosmin IV|Heart SPECT W Tc-99m Tetrofosmin IV
C0801762|T102|relax|39639-0|LNC|Brain SPECT W Tl-201 IV|Brain SPECT W Tl-201 IV
C0801762|T102|relax|42377-2|LNC|Brain CT W Xe-133 inhaled|Brain CT W Xe-133 inhaled
C0801762|T102|relax|46393-5|LNC|Liver CT W Xe-133 inhaled|Liver CT W Xe-133 inhaled
C0801762|T102|relax|42394-7|LNC|Pulmonary system CT W Xe-133 inhaled|Pulmonary system CT W Xe-133 inhaled
C0801762|T102|relax|36424-0|LNC|Abdomen CT WO contrast|Abdomen CT WO contrast
C0801762|T102|relax|30668-8|LNC|Abdomen MRI WO contrast|Abdomen MRI WO contrast
C0801762|T102|relax|42291-5|LNC|Abdomen retroperitoneum CT WO contrast|Abdomen retroperitoneum CT WO contrast
C0801762|T102|relax|36952-0|LNC|Abdomen Pelvis CT WO contrast|Abdomen Pelvis CT WO contrast
C0801762|T102|relax|36878-7|LNC|Abdominal vessels MRI angiogram WO contrast|Abdominal vessels MRI angiogram WO contrast
C0801762|T102|relax|36496-8|LNC|Acromioclavicular Joint MRI WO contrast|Acromioclavicular Joint MRI WO contrast
C0801762|T102|relax|36953-8|LNC|Adrenal gland CT WO contrast|Adrenal gland CT WO contrast
C0801762|T102|relax|36954-6|LNC|Adrenal gland MRI WO contrast|Adrenal gland MRI WO contrast
C0801762|T102|relax|36425-7|LNC|Ankle CT WO contrast|Ankle CT WO contrast
C0801762|T102|relax|30680-3|LNC|Ankle MRI WO contrast|Ankle MRI WO contrast
C0801762|T102|relax|36879-5|LNC|Ankle vessels MRI angiogram WO contrast|Ankle vessels MRI angiogram WO contrast
C0801762|T102|relax|69087-5|LNC|Ankle bilateral CT WO contrast|Ankle bilateral CT WO contrast
C0801762|T102|relax|69164-2|LNC|Ankle bilateral MRI WO contrast|Ankle bilateral MRI WO contrast
C0801762|T102|relax|36426-5|LNC|Ankle left CT WO contrast|Ankle left CT WO contrast
C0801762|T102|relax|36427-3|LNC|Ankle left MRI WO contrast|Ankle left MRI WO contrast
C0801762|T102|relax|36428-1|LNC|Ankle right CT WO contrast|Ankle right CT WO contrast
C0801762|T102|relax|36429-9|LNC|Ankle right MRI WO contrast|Ankle right MRI WO contrast
C0801762|T102|relax|36430-7|LNC|Aorta CT WO contrast|Aorta CT WO contrast
C0801762|T102|relax|44132-9|LNC|Aorta MRI angiogram WO contrast|Aorta MRI angiogram WO contrast
C0801762|T102|relax|36431-5|LNC|Aorta abdominal CT WO contrast|Aorta abdominal CT WO contrast
C0801762|T102|relax|36432-3|LNC|Aorta abdominal MRI angiogram WO contrast|Aorta abdominal MRI angiogram WO contrast
C0801762|T102|relax|69119-6|LNC|Aorta thoracic CT angiogram WO contrast|Aorta thoracic CT angiogram WO contrast
C0801762|T102|relax|36433-1|LNC|Aorta thoracic MRI angiogram WO contrast|Aorta thoracic MRI angiogram WO contrast
C0801762|T102|relax|44130-3|LNC|Aortic arch MRI angiogram WO contrast|Aortic arch MRI angiogram WO contrast
C0801762|T102|relax|36434-9|LNC|Appendix CT WO contrast|Appendix CT WO contrast
C0801762|T102|relax|44123-8|LNC|Biliary ducts Pancreatic duct MRI WO contrast|Biliary ducts Pancreatic duct MRI WO contrast
C0801762|T102|relax|30657-1|LNC|Brain MRI WO contrast|Brain MRI WO contrast
C0801762|T102|relax|48453-5|LNC|Brain temporal MRI WO contrast|Brain temporal MRI WO contrast
C0801762|T102|relax|37278-9|LNC|Brain Internal auditory canal MRI WO contrast|Brain Internal auditory canal MRI WO contrast
C0801762|T102|relax|37279-7|LNC|Brain Larynx MRI WO contrast|Brain Larynx MRI WO contrast
C0801762|T102|relax|42393-9|LNC|Brain Pituitary Sella turcica MRI WO contrast|Brain Pituitary Sella turcica MRI WO contrast
C0801762|T102|relax|36436-4|LNC|Breast MRI WO contrast|Breast MRI WO contrast
C0801762|T102|relax|69191-5|LNC|Breast implant MRI WO contrast|Breast implant MRI WO contrast
C0801762|T102|relax|69168-3|LNC|Breast implant bilateral MRI WO contrast|Breast implant bilateral MRI WO contrast
C0801762|T102|relax|38064-2|LNC|Breast implant left MRI WO contrast|Breast implant left MRI WO contrast
C0801762|T102|relax|38817-3|LNC|Breast implant right MRI WO contrast|Breast implant right MRI WO contrast
C0801762|T102|relax|44119-6|LNC|Breast bilateral CT WO contrast|Breast bilateral CT WO contrast
C0801762|T102|relax|36437-2|LNC|Breast bilateral MRI WO contrast|Breast bilateral MRI WO contrast
C0801762|T102|relax|36438-0|LNC|Breast left MRI WO contrast|Breast left MRI WO contrast
C0801762|T102|relax|36439-8|LNC|Breast right MRI WO contrast|Breast right MRI WO contrast
C0801762|T102|relax|46333-1|LNC|Breast unilateral MRI WO contrast|Breast unilateral MRI WO contrast
C0801762|T102|relax|36483-6|LNC|Calcaneus CT WO contrast|Calcaneus CT WO contrast
C0801762|T102|relax|36440-6|LNC|Calcaneus left CT WO contrast|Calcaneus left CT WO contrast
C0801762|T102|relax|36441-4|LNC|Calcaneus right CT WO contrast|Calcaneus right CT WO contrast
C0801762|T102|relax|36880-3|LNC|Carotid vessel MRI angiogram WO contrast|Carotid vessel MRI angiogram WO contrast
C0801762|T102|relax|29252-4|LNC|Chest CT WO contrast|Chest CT WO contrast
C0801762|T102|relax|36442-2|LNC|Chest MRI WO contrast|Chest MRI WO contrast
C0801762|T102|relax|69084-2|LNC|Chest vessels CT angiogram WO contrast|Chest vessels CT angiogram WO contrast
C0801762|T102|relax|36547-8|LNC|Chest vessels MRI angiogram WO contrast|Chest vessels MRI angiogram WO contrast
C0801762|T102|relax|42276-6|LNC|Chest Abdomen CT WO contrast|Chest Abdomen CT WO contrast
C0801762|T102|relax|72253-8|LNC|Chest Abdomen Pelvis CT WO contrast|Chest Abdomen Pelvis CT WO contrast
C0801762|T102|relax|42302-0|LNC|Clavicle MRI WO contrast|Clavicle MRI WO contrast
C0801762|T102|relax|48459-2|LNC|Clavicle left MRI WO contrast|Clavicle left MRI WO contrast
C0801762|T102|relax|48458-4|LNC|Clavicle right MRI WO contrast|Clavicle right MRI WO contrast
C0801762|T102|relax|36443-0|LNC|Elbow CT WO contrast|Elbow CT WO contrast
C0801762|T102|relax|30796-7|LNC|Elbow MRI WO contrast|Elbow MRI WO contrast
C0801762|T102|relax|36444-8|LNC|Elbow bilateral CT WO contrast|Elbow bilateral CT WO contrast
C0801762|T102|relax|69171-7|LNC|Elbow bilateral MRI WO contrast|Elbow bilateral MRI WO contrast
C0801762|T102|relax|36445-5|LNC|Elbow left CT WO contrast|Elbow left CT WO contrast
C0801762|T102|relax|36446-3|LNC|Elbow left MRI WO contrast|Elbow left MRI WO contrast
C0801762|T102|relax|36447-1|LNC|Elbow right CT WO contrast|Elbow right CT WO contrast
C0801762|T102|relax|36448-9|LNC|Elbow right MRI WO contrast|Elbow right MRI WO contrast
C0801762|T102|relax|42278-2|LNC|Extremity CT WO contrast|Extremity CT WO contrast
C0801762|T102|relax|69104-8|LNC|Extremity left CT WO contrast|Extremity left CT WO contrast
C0801762|T102|relax|69111-3|LNC|Extremity right CT WO contrast|Extremity right CT WO contrast
C0801762|T102|relax|36435-6|LNC|Face MRI WO contrast|Face MRI WO contrast
C0801762|T102|relax|30802-3|LNC|Facial bones Maxilla CT WO contrast|Facial bones Maxilla CT WO contrast
C0801762|T102|relax|72249-6|LNC|Facial bones Sinuses CT WO contrast|Facial bones Sinuses CT WO contrast
C0801762|T102|relax|36460-4|LNC|Femur CT WO contrast|Femur CT WO contrast
C0801762|T102|relax|69173-3|LNC|Femur bilateral MRI WO contrast|Femur bilateral MRI WO contrast
C0801762|T102|relax|36462-0|LNC|Femur left CT WO contrast|Femur left CT WO contrast
C0801762|T102|relax|36464-6|LNC|Femur right CT WO contrast|Femur right CT WO contrast
C0801762|T102|relax|69196-4|LNC|Finger MRI WO contrast|Finger MRI WO contrast
C0801762|T102|relax|69206-1|LNC|Finger left MRI WO contrast|Finger left MRI WO contrast
C0801762|T102|relax|69216-0|LNC|Finger right MRI WO contrast|Finger right MRI WO contrast
C0801762|T102|relax|36466-1|LNC|Foot CT WO contrast|Foot CT WO contrast
C0801762|T102|relax|30681-1|LNC|Foot MRI WO contrast|Foot MRI WO contrast
C0801762|T102|relax|36467-9|LNC|Foot bilateral MRI WO contrast|Foot bilateral MRI WO contrast
C0801762|T102|relax|36468-7|LNC|Foot left CT WO contrast|Foot left CT WO contrast
C0801762|T102|relax|36469-5|LNC|Foot left MRI WO contrast|Foot left MRI WO contrast
C0801762|T102|relax|36470-3|LNC|Foot right CT WO contrast|Foot right CT WO contrast
C0801762|T102|relax|36471-1|LNC|Foot right MRI WO contrast|Foot right MRI WO contrast
C0801762|T102|relax|36472-9|LNC|Forearm CT WO contrast|Forearm CT WO contrast
C0801762|T102|relax|30683-7|LNC|Forearm MRI WO contrast|Forearm MRI WO contrast
C0801762|T102|relax|69176-6|LNC|Forearm bilateral MRI WO contrast|Forearm bilateral MRI WO contrast
C0801762|T102|relax|36473-7|LNC|Forearm left CT WO contrast|Forearm left CT WO contrast
C0801762|T102|relax|36474-5|LNC|Forearm left MRI WO contrast|Forearm left MRI WO contrast
C0801762|T102|relax|36475-2|LNC|Forearm right CT WO contrast|Forearm right CT WO contrast
C0801762|T102|relax|36476-0|LNC|Forearm right MRI WO contrast|Forearm right MRI WO contrast
C0801762|T102|relax|36477-8|LNC|Hand CT WO contrast|Hand CT WO contrast
C0801762|T102|relax|30685-2|LNC|Hand MRI WO contrast|Hand MRI WO contrast
C0801762|T102|relax|69179-0|LNC|Hand bilateral MRI WO contrast|Hand bilateral MRI WO contrast
C0801762|T102|relax|36478-6|LNC|Hand left CT WO contrast|Hand left CT WO contrast
C0801762|T102|relax|36479-4|LNC|Hand left MRI WO contrast|Hand left MRI WO contrast
C0801762|T102|relax|36480-2|LNC|Hand right CT WO contrast|Hand right CT WO contrast
C0801762|T102|relax|36481-0|LNC|Hand right MRI WO contrast|Hand right MRI WO contrast
C0801762|T102|relax|30799-1|LNC|Head CT WO contrast|Head CT WO contrast
C0801762|T102|relax|36876-1|LNC|Head veins MRI angiogram WO contrast|Head veins MRI angiogram WO contrast
C0801762|T102|relax|42293-1|LNC|Head vessels CT angiogram WO contrast|Head vessels CT angiogram WO contrast
C0801762|T102|relax|36881-1|LNC|Head vessels MRI angiogram WO contrast|Head vessels MRI angiogram WO contrast
C0801762|T102|relax|36482-8|LNC|Heart MRI WO contrast|Heart MRI WO contrast
C0801762|T102|relax|36484-4|LNC|Hip CT WO contrast|Hip CT WO contrast
C0801762|T102|relax|30687-8|LNC|Hip MRI WO contrast|Hip MRI WO contrast
C0801762|T102|relax|36485-1|LNC|Hip bilateral CT WO contrast|Hip bilateral CT WO contrast
C0801762|T102|relax|36486-9|LNC|Hip bilateral MRI WO contrast|Hip bilateral MRI WO contrast
C0801762|T102|relax|36487-7|LNC|Hip left CT WO contrast|Hip left CT WO contrast
C0801762|T102|relax|36488-5|LNC|Hip left MRI WO contrast|Hip left MRI WO contrast
C0801762|T102|relax|36489-3|LNC|Hip right CT WO contrast|Hip right CT WO contrast
C0801762|T102|relax|36490-1|LNC|Hip right MRI WO contrast|Hip right MRI WO contrast
C0801762|T102|relax|30584-7|LNC|Internal auditory canal CT WO contrast|Internal auditory canal CT WO contrast
C0801762|T102|relax|30658-9|LNC|Internal auditory canal MRI WO contrast|Internal auditory canal MRI WO contrast
C0801762|T102|relax|43770-7|LNC|Kidney CT WO contrast|Kidney CT WO contrast
C0801762|T102|relax|43773-1|LNC|Kidney MRI WO contrast|Kidney MRI WO contrast
C0801762|T102|relax|36503-1|LNC|Kidney bilateral CT WO contrast|Kidney bilateral CT WO contrast
C0801762|T102|relax|36504-9|LNC|Kidney bilateral MRI WO contrast|Kidney bilateral MRI WO contrast
C0801762|T102|relax|39359-5|LNC|Kidney bilateral X-ray tomograph WO contrast|Kidney bilateral X-ray tomograph WO contrast
C0801762|T102|relax|36505-6|LNC|Knee CT WO contrast|Knee CT WO contrast
C0801762|T102|relax|30691-0|LNC|Knee MRI WO contrast|Knee MRI WO contrast
C0801762|T102|relax|69089-1|LNC|Knee bilateral CT WO contrast|Knee bilateral CT WO contrast
C0801762|T102|relax|36506-4|LNC|Knee bilateral MRI WO contrast|Knee bilateral MRI WO contrast
C0801762|T102|relax|36507-2|LNC|Knee left CT WO contrast|Knee left CT WO contrast
C0801762|T102|relax|36508-0|LNC|Knee left MRI WO contrast|Knee left MRI WO contrast
C0801762|T102|relax|36509-8|LNC|Knee right CT WO contrast|Knee right CT WO contrast
C0801762|T102|relax|36510-6|LNC|Knee right MRI WO contrast|Knee right MRI WO contrast
C0801762|T102|relax|36511-4|LNC|Larynx CT WO contrast|Larynx CT WO contrast
C0801762|T102|relax|48445-1|LNC|Larynx MRI WO contrast|Larynx MRI WO contrast
C0801762|T102|relax|30611-8|LNC|Liver CT WO contrast|Liver CT WO contrast
C0801762|T102|relax|30669-6|LNC|Liver MRI WO contrast|Liver MRI WO contrast
C0801762|T102|relax|30625-8|LNC|Lower extremity CT WO contrast|Lower extremity CT WO contrast
C0801762|T102|relax|39292-8|LNC|Lower extremity MRI WO contrast|Lower extremity MRI WO contrast
C0801762|T102|relax|44129-5|LNC|Lower extremity vessels MRI angiogram WO contrast|Lower extremity vessels MRI angiogram WO contrast
C0801762|T102|relax|36450-5|LNC|Lower extremity vessels bilateral MRI angiogram WO contrast|Lower extremity vessels bilateral MRI angiogram WO contrast
C0801762|T102|relax|36882-9|LNC|Lower extremity vessels left MRI angiogram WO contrast|Lower extremity vessels left MRI angiogram WO contrast
C0801762|T102|relax|38773-8|LNC|Lower extremity vessels right MRI angiogram WO contrast|Lower extremity vessels right MRI angiogram WO contrast
C0801762|T102|relax|36449-7|LNC|Lower extremity bilateral CT WO contrast|Lower extremity bilateral CT WO contrast
C0801762|T102|relax|36451-3|LNC|Lower extremity bilateral MRI WO contrast|Lower extremity bilateral MRI WO contrast
C0801762|T102|relax|36497-6|LNC|Lower Extremity Joint MRI WO contrast|Lower Extremity Joint MRI WO contrast
C0801762|T102|relax|36498-4|LNC|Lower extremity joint left MRI WO contrast|Lower extremity joint left MRI WO contrast
C0801762|T102|relax|36499-2|LNC|Lower extremity joint right MRI WO contrast|Lower extremity joint right MRI WO contrast
C0801762|T102|relax|36452-1|LNC|Lower extremity left CT WO contrast|Lower extremity left CT WO contrast
C0801762|T102|relax|36453-9|LNC|Lower extremity left MRI WO contrast|Lower extremity left MRI WO contrast
C0801762|T102|relax|36454-7|LNC|Lower extremity right CT WO contrast|Lower extremity right CT WO contrast
C0801762|T102|relax|36455-4|LNC|Lower extremity right MRI WO contrast|Lower extremity right MRI WO contrast
C0801762|T102|relax|36537-9|LNC|Lower leg CT WO contrast|Lower leg CT WO contrast
C0801762|T102|relax|30869-2|LNC|Lower leg MRI WO contrast|Lower leg MRI WO contrast
C0801762|T102|relax|69185-7|LNC|Lower leg bilateral MRI WO contrast|Lower leg bilateral MRI WO contrast
C0801762|T102|relax|36538-7|LNC|Lower leg left CT WO contrast|Lower leg left CT WO contrast
C0801762|T102|relax|36539-5|LNC|Lower leg left MRI WO contrast|Lower leg left MRI WO contrast
C0801762|T102|relax|36540-3|LNC|Lower leg right CT WO contrast|Lower leg right CT WO contrast
C0801762|T102|relax|36541-1|LNC|Lower leg right MRI WO contrast|Lower leg right MRI WO contrast
C0801762|T102|relax|36512-2|LNC|Mandible CT WO contrast|Mandible CT WO contrast
C0801762|T102|relax|36513-0|LNC|Nasopharynx MRI WO contrast|Nasopharynx MRI WO contrast
C0801762|T102|relax|30585-4|LNC|Nasopharynx Neck CT WO contrast|Nasopharynx Neck CT WO contrast
C0801762|T102|relax|36514-8|LNC|Neck CT WO contrast|Neck CT WO contrast
C0801762|T102|relax|30660-5|LNC|Neck MRI WO contrast|Neck MRI WO contrast
C0801762|T102|relax|36877-9|LNC|Neck veins MRI angiogram WO contrast|Neck veins MRI angiogram WO contrast
C0801762|T102|relax|36549-4|LNC|Neck vessels MRI angiogram WO contrast|Neck vessels MRI angiogram WO contrast
C0801762|T102|relax|46331-5|LNC|Orbit CT WO contrast|Orbit CT WO contrast
C0801762|T102|relax|36872-0|LNC|Orbit MRI WO contrast|Orbit MRI WO contrast
C0801762|T102|relax|30587-0|LNC|Orbit bilateral CT WO contrast|Orbit bilateral CT WO contrast
C0801762|T102|relax|30661-3|LNC|Orbit bilateral MRI WO contrast|Orbit bilateral MRI WO contrast
C0801762|T102|relax|36873-8|LNC|Orbit left MRI WO contrast|Orbit left MRI WO contrast
C0801762|T102|relax|36874-6|LNC|Orbit right MRI WO contrast|Orbit right MRI WO contrast
C0801762|T102|relax|36956-1|LNC|Orbit Face MRI WO contrast|Orbit Face MRI WO contrast
C0801762|T102|relax|46332-3|LNC|Orbit Face Neck MRI WO contrast|Orbit Face Neck MRI WO contrast
C0801762|T102|relax|36875-3|LNC|Ovary MRI WO contrast|Ovary MRI WO contrast
C0801762|T102|relax|30613-4|LNC|Pancreas CT WO contrast|Pancreas CT WO contrast
C0801762|T102|relax|36515-5|LNC|Pancreas MRI WO contrast|Pancreas MRI WO contrast
C0801762|T102|relax|37280-5|LNC|Parotid gland CT WO contrast|Parotid gland CT WO contrast
C0801762|T102|relax|37281-3|LNC|Parotid gland MRI WO contrast|Parotid gland MRI WO contrast
C0801762|T102|relax|30615-9|LNC|Pelvis CT WO contrast|Pelvis CT WO contrast
C0801762|T102|relax|30673-8|LNC|Pelvis MRI WO contrast|Pelvis MRI WO contrast
C0801762|T102|relax|36883-7|LNC|Pelvis vessels MRI angiogram WO contrast|Pelvis vessels MRI angiogram WO contrast
C0801762|T102|relax|30671-2|LNC|Pelvis Hip MRI WO contrast|Pelvis Hip MRI WO contrast
C0801762|T102|relax|30589-6|LNC|Petrous bone CT WO contrast|Petrous bone CT WO contrast
C0801762|T102|relax|30591-2|LNC|Pituitary Sella turcica CT WO contrast|Pituitary Sella turcica CT WO contrast
C0801762|T102|relax|30666-2|LNC|Pituitary Sella turcica MRI WO contrast|Pituitary Sella turcica MRI WO contrast
C0801762|T102|relax|36543-7|LNC|Portal vein MRI angiogram WO contrast|Portal vein MRI angiogram WO contrast
C0801762|T102|relax|36517-1|LNC|Posterior fossa CT WO contrast|Posterior fossa CT WO contrast
C0801762|T102|relax|36518-9|LNC|Posterior fossa MRI WO contrast|Posterior fossa MRI WO contrast
C0801762|T102|relax|36519-7|LNC|Prostate MRI WO contrast|Prostate MRI WO contrast
C0801762|T102|relax|36544-5|LNC|Renal vein MRI angiogram WO contrast|Renal vein MRI angiogram WO contrast
C0801762|T102|relax|44133-7|LNC|Renal vessels MRI angiogram WO contrast|Renal vessels MRI angiogram WO contrast
C0801762|T102|relax|36501-5|LNC|Sacroiliac Joint CT WO contrast|Sacroiliac Joint CT WO contrast
C0801762|T102|relax|36502-3|LNC|Sacroiliac Joint MRI WO contrast|Sacroiliac Joint MRI WO contrast
C0801762|T102|relax|36520-5|LNC|Sacrum CT WO contrast|Sacrum CT WO contrast
C0801762|T102|relax|36521-3|LNC|Sacrum MRI WO contrast|Sacrum MRI WO contrast
C0801762|T102|relax|36522-1|LNC|Sacrum Coccyx MRI WO contrast|Sacrum Coccyx MRI WO contrast
C0801762|T102|relax|69118-8|LNC|Scapula CT WO contrast|Scapula CT WO contrast
C0801762|T102|relax|36523-9|LNC|Scapula left MRI WO contrast|Scapula left MRI WO contrast
C0801762|T102|relax|38770-4|LNC|Scapula right MRI WO contrast|Scapula right MRI WO contrast
C0801762|T102|relax|36535-3|LNC|Scrotum Testicle MRI WO contrast|Scrotum Testicle MRI WO contrast
C0801762|T102|relax|36524-7|LNC|Shoulder CT WO contrast|Shoulder CT WO contrast
C0801762|T102|relax|30693-6|LNC|Shoulder MRI WO contrast|Shoulder MRI WO contrast
C0801762|T102|relax|69090-9|LNC|Shoulder bilateral CT WO contrast|Shoulder bilateral CT WO contrast
C0801762|T102|relax|36525-4|LNC|Shoulder bilateral MRI WO contrast|Shoulder bilateral MRI WO contrast
C0801762|T102|relax|36526-2|LNC|Shoulder left CT WO contrast|Shoulder left CT WO contrast
C0801762|T102|relax|38834-8|LNC|Shoulder left MRI WO contrast|Shoulder left MRI WO contrast
C0801762|T102|relax|36527-0|LNC|Shoulder right CT WO contrast|Shoulder right CT WO contrast
C0801762|T102|relax|36528-8|LNC|Shoulder right MRI WO contrast|Shoulder right MRI WO contrast
C0801762|T102|relax|36529-6|LNC|Sinuses CT WO contrast|Sinuses CT WO contrast
C0801762|T102|relax|30662-1|LNC|Sinuses MRI WO contrast|Sinuses MRI WO contrast
C0801762|T102|relax|44112-1|LNC|Skull base CT WO contrast|Skull base CT WO contrast
C0801762|T102|relax|48687-8|LNC|Skull base MRI WO contrast|Skull base MRI WO contrast
C0801762|T102|relax|37293-8|LNC|Soft tissue MRI WO contrast|Soft tissue MRI WO contrast
C0801762|T102|relax|37510-5|LNC|Spine vessels MRI angiogram WO contrast|Spine vessels MRI angiogram WO contrast
C0801762|T102|relax|30592-0|LNC|Spine Cervical CT WO contrast|Spine Cervical CT WO contrast
C0801762|T102|relax|30667-0|LNC|Spine Cervical MRI WO contrast|Spine Cervical MRI WO contrast
C0801762|T102|relax|37511-3|LNC|Cervical Spine vessels MRI angiogram WO contrast|Cervical Spine vessels MRI angiogram WO contrast
C0801762|T102|relax|30854-4|LNC|Spine Cervical Thoracic Lumbar MRI WO contrast|Spine Cervical Thoracic Lumbar MRI WO contrast
C0801762|T102|relax|30620-9|LNC|Spine Lumbar CT WO contrast|Spine Lumbar CT WO contrast
C0801762|T102|relax|30679-5|LNC|Spine Lumbar MRI WO contrast|Spine Lumbar MRI WO contrast
C0801762|T102|relax|37994-1|LNC|Lumbar Spine vessels MRI angiogram WO contrast|Lumbar Spine vessels MRI angiogram WO contrast
C0801762|T102|relax|37288-8|LNC|Spine Lumbosacral Junction CT WO contrast|Spine Lumbosacral Junction CT WO contrast
C0801762|T102|relax|30597-9|LNC|Spine Thoracic CT WO contrast|Spine Thoracic CT WO contrast
C0801762|T102|relax|36532-0|LNC|Spine Thoracic MRI WO contrast|Spine Thoracic MRI WO contrast
C0801762|T102|relax|37512-1|LNC|Thoracic Spine vessels MRI angiogram WO contrast|Thoracic Spine vessels MRI angiogram WO contrast
C0801762|T102|relax|30621-7|LNC|Spleen CT WO contrast|Spleen CT WO contrast
C0801762|T102|relax|36533-8|LNC|Spleen MRI WO contrast|Spleen MRI WO contrast
C0801762|T102|relax|37282-1|LNC|Sternoclavicular Joint CT WO contrast|Sternoclavicular Joint CT WO contrast
C0801762|T102|relax|36534-6|LNC|Sternum CT WO contrast|Sternum CT WO contrast
C0801762|T102|relax|44230-1|LNC|Superior mesenteric vessels MRI angiogram WO contrast|Superior mesenteric vessels MRI angiogram WO contrast
C0801762|T102|relax|36866-2|LNC|Temporal bone CT WO contrast|Temporal bone CT WO contrast
C0801762|T102|relax|36867-0|LNC|Temporal bone left CT WO contrast|Temporal bone left CT WO contrast
C0801762|T102|relax|36868-8|LNC|Temporal bone right CT WO contrast|Temporal bone right CT WO contrast
C0801762|T102|relax|37283-9|LNC|Temporomandibular joint CT WO contrast|Temporomandibular joint CT WO contrast
C0801762|T102|relax|37284-7|LNC|Temporomandibular joint MRI WO contrast|Temporomandibular joint MRI WO contrast
C0801762|T102|relax|37285-4|LNC|Temporomandibular joint bilateral MRI WO contrast|Temporomandibular joint bilateral MRI WO contrast
C0801762|T102|relax|37286-2|LNC|Temporomandibular joint left MRI WO contrast|Temporomandibular joint left MRI WO contrast
C0801762|T102|relax|37287-0|LNC|Temporomandibular joint right MRI WO contrast|Temporomandibular joint right MRI WO contrast
C0801762|T102|relax|36461-2|LNC|Thigh MRI WO contrast|Thigh MRI WO contrast
C0801762|T102|relax|43514-9|LNC|Thigh vessels left MRI angiogram WO contrast|Thigh vessels left MRI angiogram WO contrast
C0801762|T102|relax|43515-6|LNC|Thigh vessels right MRI angiogram WO contrast|Thigh vessels right MRI angiogram WO contrast
C0801762|T102|relax|36463-8|LNC|Thigh left MRI WO contrast|Thigh left MRI WO contrast
C0801762|T102|relax|36465-3|LNC|Thigh right MRI WO contrast|Thigh right MRI WO contrast
C0801762|T102|relax|30654-8|LNC|Thoracic outlet MRI WO contrast|Thoracic outlet MRI WO contrast
C0801762|T102|relax|38833-0|LNC|Thoracic outlet left MRI WO contrast|Thoracic outlet left MRI WO contrast
C0801762|T102|relax|36516-3|LNC|Thoracic outlet right MRI WO contrast|Thoracic outlet right MRI WO contrast
C0801762|T102|relax|36955-3|LNC|Thyroid CT WO contrast|Thyroid CT WO contrast
C0801762|T102|relax|36536-1|LNC|Thyroid MRI WO contrast|Thyroid MRI WO contrast
C0801762|T102|relax|72242-1|LNC|Toes left MRI WO contrast|Toes left MRI WO contrast
C0801762|T102|relax|72239-7|LNC|Toes right MRI WO contrast|Toes right MRI WO contrast
C0801762|T102|relax|36491-9|LNC|Upper arm CT WO contrast|Upper arm CT WO contrast
C0801762|T102|relax|30689-4|LNC|Upper arm MRI WO contrast|Upper arm MRI WO contrast
C0801762|T102|relax|69183-2|LNC|Upper arm bilateral MRI WO contrast|Upper arm bilateral MRI WO contrast
C0801762|T102|relax|36492-7|LNC|Upper arm left CT WO contrast|Upper arm left CT WO contrast
C0801762|T102|relax|36493-5|LNC|Upper arm left MRI WO contrast|Upper arm left MRI WO contrast
C0801762|T102|relax|36494-3|LNC|Upper arm right CT WO contrast|Upper arm right CT WO contrast
C0801762|T102|relax|36495-0|LNC|Upper arm right MRI WO contrast|Upper arm right MRI WO contrast
C0801762|T102|relax|30627-4|LNC|Upper extremity CT WO contrast|Upper extremity CT WO contrast
C0801762|T102|relax|39033-6|LNC|Upper extremity MRI WO contrast|Upper extremity MRI WO contrast
C0801762|T102|relax|36548-6|LNC|Upper extremity vessels MRI angiogram WO contrast|Upper extremity vessels MRI angiogram WO contrast
C0801762|T102|relax|36456-2|LNC|Upper extremity bilateral CT WO contrast|Upper extremity bilateral CT WO contrast
C0801762|T102|relax|69188-1|LNC|Upper extremity bilateral MRI WO contrast|Upper extremity bilateral MRI WO contrast
C0801762|T102|relax|36500-7|LNC|Upper extremity  joint MRI WO contrast|Upper extremity  joint MRI WO contrast
C0801762|T102|relax|36869-6|LNC|Upper extremity joint left MRI WO contrast|Upper extremity joint left MRI WO contrast
C0801762|T102|relax|36870-4|LNC|Upper extremity joint right MRI WO contrast|Upper extremity joint right MRI WO contrast
C0801762|T102|relax|36457-0|LNC|Upper extremity left CT WO contrast|Upper extremity left CT WO contrast
C0801762|T102|relax|38832-2|LNC|Upper extremity left MRI WO contrast|Upper extremity left MRI WO contrast
C0801762|T102|relax|36458-8|LNC|Upper extremity right CT WO contrast|Upper extremity right CT WO contrast
C0801762|T102|relax|36459-6|LNC|Upper extremity right MRI WO contrast|Upper extremity right MRI WO contrast
C0801762|T102|relax|36542-9|LNC|Uterus MRI WO contrast|Uterus MRI WO contrast
C0801762|T102|relax|36545-2|LNC|Inferior vena cava MRI WO contrast|Inferior vena cava MRI WO contrast
C0801762|T102|relax|36546-0|LNC|Superior vena cava MRI WO contrast|Superior vena cava MRI WO contrast
C0801762|T102|relax|37459-5|LNC|Wrist CT WO contrast|Wrist CT WO contrast
C0801762|T102|relax|37460-3|LNC|Wrist MRI WO contrast|Wrist MRI WO contrast
C0801762|T102|relax|43516-4|LNC|Wrist vessels left MRI angiogram WO contrast|Wrist vessels left MRI angiogram WO contrast
C0801762|T102|relax|43517-2|LNC|Wrist vessels right MRI angiogram WO contrast|Wrist vessels right MRI angiogram WO contrast
C0801762|T102|relax|37461-1|LNC|Wrist bilateral CT WO contrast|Wrist bilateral CT WO contrast
C0801762|T102|relax|37462-9|LNC|Wrist bilateral MRI WO contrast|Wrist bilateral MRI WO contrast
C0801762|T102|relax|37463-7|LNC|Wrist left CT WO contrast|Wrist left CT WO contrast
C0801762|T102|relax|37464-5|LNC|Wrist left MRI WO contrast|Wrist left MRI WO contrast
C0801762|T102|relax|37465-2|LNC|Wrist right CT WO contrast|Wrist right CT WO contrast
C0801762|T102|relax|37466-0|LNC|Wrist right MRI WO contrast|Wrist right MRI WO contrast
C0801762|T102|relax|43525-5|LNC|Unspecified body region CT WO contrast|Unspecified body region CT WO contrast
C0801762|T102|relax|69223-6|LNC|Unspecified body region MRI WO contrast|Unspecified body region MRI WO contrast
C0801762|T102|relax|36871-2|LNC|Joint MRI WO contrast|Joint MRI WO contrast
C0801762|T102|relax|24787-4|LNC|Kidney bilateral X-ray tomograph WO contrast 10M post contrast IV|Kidney bilateral X-ray tomograph WO contrast 10M post contrast IV
C0801762|T102|relax|30712-4|LNC|Hip US WO developmental joint assessment|Hip US WO developmental joint assessment
C0801762|T102|relax|25051-4|LNC|Unspecified body region CT Multisectional sagittal|Unspecified body region CT Multisectional sagittal
C0801762|T102|relax|25060-5|LNC|Unspecified body region US No charge|Unspecified body region US No charge
C0801762|T102|relax|24620-7|LNC|Catheter Fluoroscopy Patency check W contrast via catheter|Catheter Fluoroscopy Patency check W contrast via catheter
C0801762|T102|relax|24882-3|LNC|Popliteal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty vessel W contrast IA|Popliteal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty vessel W contrast IA
C0801762|T102|relax|69252-5|LNC|Pulmonary artery Fluoroscopic angiogram Percutaneous transluminal angioplasty vessel W contrast IA|Pulmonary artery Fluoroscopic angiogram Percutaneous transluminal angioplasty vessel W contrast IA
C0801762|T102|relax|69248-3|LNC|Renal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty vessel W contrast IA|Renal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty vessel W contrast IA
C0801762|T102|relax|69301-0|LNC|Upper extremity vein Fluoroscopic angiogram Percutaneous transluminal angioplasty vessel W contrast IV|Upper extremity vein Fluoroscopic angiogram Percutaneous transluminal angioplasty vessel W contrast IV
C0801762|T102|relax|24875-7|LNC|Peripheral vessel US doppler Peripheral plane|Peripheral vessel US doppler Peripheral plane
C0801762|T102|relax|24998-7|LNC|Placement check gastrostomy tube W contrast via GI tube|Placement check gastrostomy tube W contrast via GI tube
C0801762|T102|relax|44226-9|LNC|Colon Fluoroscopy Reduction W views W barium contrast PR|Colon Fluoroscopy Reduction W views W barium contrast PR
C0801762|T102|relax|30636-5|LNC|Colon Fluoroscopy Reduction W views W contrast PR|Colon Fluoroscopy Reduction W views W contrast PR
C0801762|T102|relax|25073-8|LNC|Vessel Fluoroscopic angiogram Removal foreign body from vascular space|Vessel Fluoroscopic angiogram Removal foreign body from vascular space
C0801762|T102|relax|25015-9|LNC|Upper GI tract Replacement percutaneous gastrojejunostomy|Upper GI tract Replacement percutaneous gastrojejunostomy
C0801762|T102|relax|29757-2|LNC|Colposcopy study|Colposcopy study
C0801762|T102|relax|18746-8|LNC|Colonoscopy study|Colonoscopy study
C0801762|T102|relax|18753-4|LNC|Flexible sigmoidoscopy study|Flexible sigmoidoscopy study
C0801762|T102|relax|11525-3|LNC|Obstetrical ultrasound study|Obstetrical ultrasound study
C0801762|T102|relax|18744-3|LNC|Bronchoscopy study|Bronchoscopy study
C0801762|T102|relax|38269-7|LNC|Study report Skeletal system DXA|Study report Skeletal system DXA
C0801762|T102|relax|17787-3|LNC|Thyroid Scan Study report|Thyroid Scan Study report
C0801762|T102|relax|18751-8|LNC|Endoscopy study|Endoscopy study
C0801762|T102|relax|18748-4|LNC|Diagnostic imaging study|Diagnostic imaging study
C0801762|T102|relax|24783-3|LNC|Kidney bilateral Fluoroscopy Urodynamics|Kidney bilateral Fluoroscopy Urodynamics
C0801762|T102|relax|25065-4|LNC|Unspecified body region Fluoroscopy 15 minutes|Unspecified body region Fluoroscopy 15 minutes
C0801762|T102|relax|25068-8|LNC|Unspecified body region Fluoroscopy 1 hour|Unspecified body region Fluoroscopy 1 hour
C0801762|T102|relax|43471-2|LNC|Unspecified body region Fluoroscopy 2 hour|Unspecified body region Fluoroscopy 2 hour
C0801762|T102|relax|25066-2|LNC|Unspecified body region Fluoroscopy 30 minutes|Unspecified body region Fluoroscopy 30 minutes
C0801762|T102|relax|25067-0|LNC|Unspecified body region Fluoroscopy 45 minutes|Unspecified body region Fluoroscopy 45 minutes
C0801762|T102|relax|43472-0|LNC|Unspecified body region Fluoroscopy 90 minutes|Unspecified body region Fluoroscopy 90 minutes
C0801762|T102|relax|42702-1|LNC|Unspecified body region Fluoroscopy Greater than 1 hour|Unspecified body region Fluoroscopy Greater than 1 hour
C0801762|T102|relax|42703-9|LNC|Unspecified body region Fluoroscopy Less than 1 hour|Unspecified body region Fluoroscopy Less than 1 hour
C0801762|T102|relax|36550-2|LNC|Abdomen X-ray Single view|Abdomen X-ray Single view
C0801762|T102|relax|36551-0|LNC|Ankle X-ray Single view|Ankle X-ray Single view
C0801762|T102|relax|69307-7|LNC|Ankle left X-ray Single view|Ankle left X-ray Single view
C0801762|T102|relax|69314-3|LNC|Ankle right X-ray Single view|Ankle right X-ray Single view
C0801762|T102|relax|46335-6|LNC|Breast bilateral Mammogram Single view|Breast bilateral Mammogram Single view
C0801762|T102|relax|46336-4|LNC|Breast left Mammogram Single view|Breast left Mammogram Single view
C0801762|T102|relax|46337-2|LNC|Breast right Mammogram Single view|Breast right Mammogram Single view
C0801762|T102|relax|46338-0|LNC|Breast unilateral Mammogram Single view|Breast unilateral Mammogram Single view
C0801762|T102|relax|36564-3|LNC|Calcaneus X-ray Single view|Calcaneus X-ray Single view
C0801762|T102|relax|69311-9|LNC|Calcaneus left X-ray Single view|Calcaneus left X-ray Single view
C0801762|T102|relax|69319-2|LNC|Calcaneus right X-ray Single view|Calcaneus right X-ray Single view
C0801762|T102|relax|36554-4|LNC|Chest X-ray Single view|Chest X-ray Single view
C0801762|T102|relax|42699-9|LNC|Chest Abdomen X-ray Single view|Chest Abdomen X-ray Single view
C0801762|T102|relax|36555-1|LNC|Clavicle X-ray Single view|Clavicle X-ray Single view
C0801762|T102|relax|36556-9|LNC|Elbow X-ray Single view|Elbow X-ray Single view
C0801762|T102|relax|69308-5|LNC|Elbow left X-ray Single view|Elbow left X-ray Single view
C0801762|T102|relax|69315-0|LNC|Elbow right X-ray Single view|Elbow right X-ray Single view
C0801762|T102|relax|42153-7|LNC|Extremity X-ray Single view|Extremity X-ray Single view
C0801762|T102|relax|36559-3|LNC|Femur X-ray Single view|Femur X-ray Single view
C0801762|T102|relax|36560-1|LNC|Femur left X-ray Single view|Femur left X-ray Single view
C0801762|T102|relax|37689-7|LNC|Femur right X-ray Single view|Femur right X-ray Single view
C0801762|T102|relax|36561-9|LNC|Foot X-ray Single view|Foot X-ray Single view
C0801762|T102|relax|69309-3|LNC|Foot left X-ray Single view|Foot left X-ray Single view
C0801762|T102|relax|69316-8|LNC|Foot right X-ray Single view|Foot right X-ray Single view
C0801762|T102|relax|36563-5|LNC|Hand X-ray Single view|Hand X-ray Single view
C0801762|T102|relax|69310-1|LNC|Hand left X-ray Single view|Hand left X-ray Single view
C0801762|T102|relax|69318-4|LNC|Hand right X-ray Single view|Hand right X-ray Single view
C0801762|T102|relax|24761-9|LNC|Hip X-ray Single view|Hip X-ray Single view
C0801762|T102|relax|26400-2|LNC|Hip bilateral X-ray Single view|Hip bilateral X-ray Single view
C0801762|T102|relax|26401-0|LNC|Hip left X-ray Single view|Hip left X-ray Single view
C0801762|T102|relax|26402-8|LNC|Hip right X-ray Single view|Hip right X-ray Single view
C0801762|T102|relax|36565-0|LNC|Humerus X-ray Single view|Humerus X-ray Single view
C0801762|T102|relax|69312-7|LNC|Humerus left X-ray Single view|Humerus left X-ray Single view
C0801762|T102|relax|69320-0|LNC|Humerus right X-ray Single view|Humerus right X-ray Single view
C0801762|T102|relax|36566-8|LNC|Knee bilateral X-ray Single view|Knee bilateral X-ray Single view
C0801762|T102|relax|36567-6|LNC|Knee left X-ray Single view|Knee left X-ray Single view
C0801762|T102|relax|37741-6|LNC|Knee right X-ray Single view|Knee right X-ray Single view
C0801762|T102|relax|36557-7|LNC|Lower extremity bilateral X-ray Single view|Lower extremity bilateral X-ray Single view
C0801762|T102|relax|36558-5|LNC|Lower extremity left X-ray Single view|Lower extremity left X-ray Single view
C0801762|T102|relax|37764-8|LNC|Lower extremity right X-ray Single view|Lower extremity right X-ray Single view
C0801762|T102|relax|37614-5|LNC|Patella X-ray Single view|Patella X-ray Single view
C0801762|T102|relax|69152-7|LNC|Patella left X-ray Single view|Patella left X-ray Single view
C0801762|T102|relax|69260-8|LNC|Patella right X-ray Single view|Patella right X-ray Single view
C0801762|T102|relax|37616-0|LNC|Pelvis X-ray Single view|Pelvis X-ray Single view
C0801762|T102|relax|69317-6|LNC|Radius right Ulna right X-ray Single view|Radius right Ulna right X-ray Single view
C0801762|T102|relax|42313-7|LNC|Ribs left X-ray Single view|Ribs left X-ray Single view
C0801762|T102|relax|42314-5|LNC|Ribs right X-ray Single view|Ribs right X-ray Single view
C0801762|T102|relax|37654-1|LNC|Scapula X-ray Single view|Scapula X-ray Single view
C0801762|T102|relax|30748-8|LNC|Shoulder X-ray Single view|Shoulder X-ray Single view
C0801762|T102|relax|36568-4|LNC|Shoulder bilateral X-ray Single view|Shoulder bilateral X-ray Single view
C0801762|T102|relax|36569-2|LNC|Shoulder left X-ray Single view|Shoulder left X-ray Single view
C0801762|T102|relax|37792-9|LNC|Shoulder right X-ray Single view|Shoulder right X-ray Single view
C0801762|T102|relax|37851-3|LNC|Sinuses X-ray Single view|Sinuses X-ray Single view
C0801762|T102|relax|24917-7|LNC|Skull X-ray Single view|Skull X-ray Single view
C0801762|T102|relax|48695-1|LNC|Skull base X-ray Single view|Skull base X-ray Single view
C0801762|T102|relax|24940-9|LNC|Spine Cervical X-ray Single view|Spine Cervical X-ray Single view
C0801762|T102|relax|30773-6|LNC|Spine Lumbar X-ray Single view|Spine Lumbar X-ray Single view
C0801762|T102|relax|37904-0|LNC|Spine Thoracic X-ray Single view|Spine Thoracic X-ray Single view
C0801762|T102|relax|38121-0|LNC|Spine Thoracic Lumbar X-ray Single view|Spine Thoracic Lumbar X-ray Single view
C0801762|T102|relax|69313-5|LNC|Tibia left Fibula left X-ray Single view|Tibia left Fibula left X-ray Single view
C0801762|T102|relax|69321-8|LNC|Tibia right Fibula right X-ray Single view|Tibia right Fibula right X-ray Single view
C0801762|T102|relax|37894-3|LNC|Tibia Fibula X-ray Single view|Tibia Fibula X-ray Single view
C0801762|T102|relax|37924-8|LNC|Wrist X-ray Single view|Wrist X-ray Single view
C0801762|T102|relax|42419-2|LNC|Wrist bilateral X-ray Single view|Wrist bilateral X-ray Single view
C0801762|T102|relax|36570-0|LNC|Wrist left X-ray Single view|Wrist left X-ray Single view
C0801762|T102|relax|37825-7|LNC|Wrist right X-ray Single view|Wrist right X-ray Single view
C0801762|T102|relax|30642-3|LNC|Unspecified body region Fluoroscopy Single view|Unspecified body region Fluoroscopy Single view
C0801762|T102|relax|30787-6|LNC|Joint X-ray Single view|Joint X-ray Single view
C0801762|T102|relax|44176-6|LNC|Hip X-ray Single view portable|Hip X-ray Single view portable
C0801762|T102|relax|41775-8|LNC|Pelvis X-ray Single view portable|Pelvis X-ray Single view portable
C0801762|T102|relax|30749-6|LNC|Shoulder X-ray Single view portable|Shoulder X-ray Single view portable
C0801762|T102|relax|30722-3|LNC|Skull X-ray Single view portable|Skull X-ray Single view portable
C0801762|T102|relax|30724-9|LNC|Spine Cervical X-ray Single view portable|Spine Cervical X-ray Single view portable
C0801762|T102|relax|30774-4|LNC|Spine Lumbar X-ray Single view portable|Spine Lumbar X-ray Single view portable
C0801762|T102|relax|70932-9|LNC|Spine Thoracic X-ray Single view portable|Spine Thoracic X-ray Single view portable
C0801762|T102|relax|25063-9|LNC|Vessel Fluoroscopic angiogram Single view W contrast IA|Vessel Fluoroscopic angiogram Single view W contrast IA
C0801762|T102|relax|69268-1|LNC|Breast duct Mammogram Single view W contrast intra duct|Breast duct Mammogram Single view W contrast intra duct
C0801762|T102|relax|49510-1|LNC|Breast duct left Mammogram Single view W contrast intra duct|Breast duct left Mammogram Single view W contrast intra duct
C0801762|T102|relax|49509-3|LNC|Breast duct right Mammogram Single view W contrast intra duct|Breast duct right Mammogram Single view W contrast intra duct
C0801762|T102|relax|24715-5|LNC|Gastrointestine upper Fluoroscopy Single view W contrast PO|Gastrointestine upper Fluoroscopy Single view W contrast PO
C0801762|T102|relax|37513-9|LNC|Tibia bilateral X-ray 10 degree caudal angle|Tibia bilateral X-ray 10 degree caudal angle
C0801762|T102|relax|37514-7|LNC|Tibia left X-ray 10 degree caudal angle|Tibia left X-ray 10 degree caudal angle
C0801762|T102|relax|38806-6|LNC|Tibia right X-ray 10 degree caudal angle|Tibia right X-ray 10 degree caudal angle
C0801762|T102|relax|37467-8|LNC|Acromioclavicular Joint X-ray 10 degree cephalic angle|Acromioclavicular Joint X-ray 10 degree cephalic angle
C0801762|T102|relax|37468-6|LNC|Shoulder bilateral X-ray 30 degree caudal angle|Shoulder bilateral X-ray 30 degree caudal angle
C0801762|T102|relax|42431-7|LNC|Knee right X-ray 30 degree standing|Knee right X-ray 30 degree standing
C0801762|T102|relax|69079-2|LNC|Clavicle X-ray 45 degree cephalic angle|Clavicle X-ray 45 degree cephalic angle
C0801762|T102|relax|37469-4|LNC|Clavicle bilateral X-ray 45 degree cephalic angle|Clavicle bilateral X-ray 45 degree cephalic angle
C0801762|T102|relax|37470-2|LNC|Clavicle left X-ray 45 degree cephalic angle|Clavicle left X-ray 45 degree cephalic angle
C0801762|T102|relax|38803-3|LNC|Clavicle right X-ray 45 degree cephalic angle|Clavicle right X-ray 45 degree cephalic angle
C0801762|T102|relax|24799-9|LNC|Abdomen X-ray AP single view|Abdomen X-ray AP single view
C0801762|T102|relax|36583-3|LNC|Acromioclavicular joint left X-ray AP single view|Acromioclavicular joint left X-ray AP single view
C0801762|T102|relax|37662-4|LNC|Acromioclavicular joint right X-ray AP single view|Acromioclavicular joint right X-ray AP single view
C0801762|T102|relax|36571-8|LNC|Ankle X-ray AP single view|Ankle X-ray AP single view
C0801762|T102|relax|36572-6|LNC|Chest X-ray AP single view|Chest X-ray AP single view
C0801762|T102|relax|36573-4|LNC|Clavicle X-ray AP single view|Clavicle X-ray AP single view
C0801762|T102|relax|36575-9|LNC|Femur X-ray AP single view|Femur X-ray AP single view
C0801762|T102|relax|36576-7|LNC|Finger fifth X-ray AP single view|Finger fifth X-ray AP single view
C0801762|T102|relax|36577-5|LNC|Finger fourth X-ray AP single view|Finger fourth X-ray AP single view
C0801762|T102|relax|36578-3|LNC|Finger third X-ray AP single view|Finger third X-ray AP single view
C0801762|T102|relax|36579-1|LNC|Foot X-ray AP single view|Foot X-ray AP single view
C0801762|T102|relax|36580-9|LNC|Foot bilateral X-ray AP single view|Foot bilateral X-ray AP single view
C0801762|T102|relax|36581-7|LNC|Hip X-ray AP single view|Hip X-ray AP single view
C0801762|T102|relax|36582-5|LNC|Hip left X-ray AP single view|Hip left X-ray AP single view
C0801762|T102|relax|37726-7|LNC|Hip right X-ray AP single view|Hip right X-ray AP single view
C0801762|T102|relax|36584-1|LNC|Knee X-ray AP single view|Knee X-ray AP single view
C0801762|T102|relax|36585-8|LNC|Knee bilateral X-ray AP single view|Knee bilateral X-ray AP single view
C0801762|T102|relax|48462-6|LNC|Knee left X-ray AP single view|Knee left X-ray AP single view
C0801762|T102|relax|48463-4|LNC|Knee right X-ray AP single view|Knee right X-ray AP single view
C0801762|T102|relax|36574-2|LNC|Lower extremity X-ray AP single view|Lower extremity X-ray AP single view
C0801762|T102|relax|42439-0|LNC|Neck X-ray AP single view|Neck X-ray AP single view
C0801762|T102|relax|37622-8|LNC|Pelvis X-ray AP single view|Pelvis X-ray AP single view
C0801762|T102|relax|39050-0|LNC|Ribs X-ray AP single view|Ribs X-ray AP single view
C0801762|T102|relax|36958-7|LNC|Ribs bilateral X-ray AP single view|Ribs bilateral X-ray AP single view
C0801762|T102|relax|36959-5|LNC|Ribs left X-ray AP single view|Ribs left X-ray AP single view
C0801762|T102|relax|37783-8|LNC|Ribs right X-ray AP single view|Ribs right X-ray AP single view
C0801762|T102|relax|39048-4|LNC|Scapula X-ray AP single view|Scapula X-ray AP single view
C0801762|T102|relax|37842-2|LNC|Shoulder X-ray AP single view|Shoulder X-ray AP single view
C0801762|T102|relax|36586-6|LNC|Shoulder bilateral X-ray AP single view|Shoulder bilateral X-ray AP single view
C0801762|T102|relax|36587-4|LNC|Shoulder left X-ray AP single view|Shoulder left X-ray AP single view
C0801762|T102|relax|37798-6|LNC|Shoulder right X-ray AP single view|Shoulder right X-ray AP single view
C0801762|T102|relax|69269-9|LNC|Skull X-ray AP single view|Skull X-ray AP single view
C0801762|T102|relax|30725-6|LNC|Spine Cervical X-ray AP single view|Spine Cervical X-ray AP single view
C0801762|T102|relax|24948-2|LNC|Spine Cervical Odontoid Cervical axis X-ray AP single view|Spine Cervical Odontoid Cervical axis X-ray AP single view
C0801762|T102|relax|30777-7|LNC|Spine Lumbar X-ray AP single view|Spine Lumbar X-ray AP single view
C0801762|T102|relax|30752-0|LNC|Spine Thoracic X-ray AP single view|Spine Thoracic X-ray AP single view
C0801762|T102|relax|39049-2|LNC|Spine Thoracic Lumbar X-ray AP single view|Spine Thoracic Lumbar X-ray AP single view
C0801762|T102|relax|37880-2|LNC|Sternoclavicular Joint X-ray AP single view|Sternoclavicular Joint X-ray AP single view
C0801762|T102|relax|37890-1|LNC|Thumb X-ray AP single view|Thumb X-ray AP single view
C0801762|T102|relax|37897-6|LNC|Tibia Fibula X-ray AP single view|Tibia Fibula X-ray AP single view
C0801762|T102|relax|39402-3|LNC|Shoulder X-ray AP (W internal rotation W external rotation)|Shoulder X-ray AP (W internal rotation W external rotation)
C0801762|T102|relax|37634-3|LNC|Pelvis X-ray AP 20 degree cephalic angle|Pelvis X-ray AP 20 degree cephalic angle
C0801762|T102|relax|30734-8|LNC|Chest X-ray AP lateral-decubitus|Chest X-ray AP lateral-decubitus
C0801762|T102|relax|30735-5|LNC|Chest X-ray AP lateral-decubitus portable|Chest X-ray AP lateral-decubitus portable
C0801762|T102|relax|24561-3|LNC|Abdomen X-ray AP left lateral-decubitus|Abdomen X-ray AP left lateral-decubitus
C0801762|T102|relax|24637-1|LNC|Chest X-ray AP left lateral-decubitus|Chest X-ray AP left lateral-decubitus
C0801762|T102|relax|24560-5|LNC|Abdomen X-ray AP left lateral-decubitus portable|Abdomen X-ray AP left lateral-decubitus portable
C0801762|T102|relax|24636-3|LNC|Chest X-ray AP left lateral-decubitus portable|Chest X-ray AP left lateral-decubitus portable
C0801762|T102|relax|36588-2|LNC|Abdomen X-ray AP portable single view|Abdomen X-ray AP portable single view
C0801762|T102|relax|36589-0|LNC|Chest X-ray AP portable single view|Chest X-ray AP portable single view
C0801762|T102|relax|30727-2|LNC|Spine Cervical X-ray AP portable single view|Spine Cervical X-ray AP portable single view
C0801762|T102|relax|30729-8|LNC|Spine Cervical Odontoid Cervical axis X-ray AP portable single view|Spine Cervical Odontoid Cervical axis X-ray AP portable single view
C0801762|T102|relax|30755-3|LNC|Spine Thoracic X-ray AP portable single view|Spine Thoracic X-ray AP portable single view
C0801762|T102|relax|24563-9|LNC|Abdomen X-ray AP right lateral-decubitus|Abdomen X-ray AP right lateral-decubitus
C0801762|T102|relax|43466-2|LNC|Chest X-ray AP right lateral-decubitus|Chest X-ray AP right lateral-decubitus
C0801762|T102|relax|24652-0|LNC|Chest X-ray AP right lateral-decubitus portable|Chest X-ray AP right lateral-decubitus portable
C0801762|T102|relax|43778-0|LNC|Chest X-ray AP supine portable|Chest X-ray AP supine portable
C0801762|T102|relax|24564-7|LNC|Abdomen X-ray AP upright portable|Abdomen X-ray AP upright portable
C0801762|T102|relax|36960-3|LNC|Chest X-ray AP upright portable|Chest X-ray AP upright portable
C0801762|T102|relax|24807-0|LNC|Knee X-ray AP single view standing|Knee X-ray AP single view standing
C0801762|T102|relax|26358-2|LNC|Knee bilateral X-ray AP single view standing|Knee bilateral X-ray AP single view standing
C0801762|T102|relax|26359-0|LNC|Knee left X-ray AP single view standing|Knee left X-ray AP single view standing
C0801762|T102|relax|26360-8|LNC|Knee right X-ray AP single view standing|Knee right X-ray AP single view standing
C0801762|T102|relax|44177-4|LNC|Lower extremity bilateral X-ray AP single view standing|Lower extremity bilateral X-ray AP single view standing
C0801762|T102|relax|38849-6|LNC|Lower extremity left X-ray AP single view standing|Lower extremity left X-ray AP single view standing
C0801762|T102|relax|37733-3|LNC|Lower extremity right X-ray AP single view standing|Lower extremity right X-ray AP single view standing
C0801762|T102|relax|42420-0|LNC|Pelvis X-ray AP single view standing|Pelvis X-ray AP single view standing
C0801762|T102|relax|42378-0|LNC|Spine Lumbar X-ray AP single view W left bending|Spine Lumbar X-ray AP single view W left bending
C0801762|T102|relax|39410-6|LNC|Spine Thoracic X-ray AP single view W left bending|Spine Thoracic X-ray AP single view W left bending
C0801762|T102|relax|42379-8|LNC|Spine Lumbar X-ray AP single view W right bending|Spine Lumbar X-ray AP single view W right bending
C0801762|T102|relax|39411-4|LNC|Spine Thoracic X-ray AP single view W right bending|Spine Thoracic X-ray AP single view W right bending
C0801762|T102|relax|24723-9|LNC|Hand X-ray arthritis|Hand X-ray arthritis
C0801762|T102|relax|26355-8|LNC|Hand bilateral X-ray arthritis|Hand bilateral X-ray arthritis
C0801762|T102|relax|26356-6|LNC|Hand left X-ray arthritis|Hand left X-ray arthritis
C0801762|T102|relax|26357-4|LNC|Hand right X-ray arthritis|Hand right X-ray arthritis
C0801762|T102|relax|42395-4|LNC|Foot sesamoid bones bilateral X-ray axial|Foot sesamoid bones bilateral X-ray axial
C0801762|T102|relax|42396-2|LNC|Foot sesamoid bones left X-ray axial|Foot sesamoid bones left X-ray axial
C0801762|T102|relax|36962-9|LNC|Breast Mammogram axillary|Breast Mammogram axillary
C0801762|T102|relax|37849-7|LNC|Shoulder X-ray axillary|Shoulder X-ray axillary
C0801762|T102|relax|36963-7|LNC|Shoulder bilateral X-ray axillary|Shoulder bilateral X-ray axillary
C0801762|T102|relax|36964-5|LNC|Shoulder left X-ray axillary|Shoulder left X-ray axillary
C0801762|T102|relax|37800-0|LNC|Shoulder right X-ray axillary|Shoulder right X-ray axillary
C0801762|T102|relax|36965-2|LNC|Hand X-ray Ball Catcher|Hand X-ray Ball Catcher
C0801762|T102|relax|37471-0|LNC|Hand bilateral X-ray Bora|Hand bilateral X-ray Bora
C0801762|T102|relax|37472-8|LNC|Hand left X-ray Bora|Hand left X-ray Bora
C0801762|T102|relax|38804-1|LNC|Hand right X-ray Bora|Hand right X-ray Bora
C0801762|T102|relax|36966-0|LNC|Hand bilateral X-ray Brewerton|Hand bilateral X-ray Brewerton
C0801762|T102|relax|36967-8|LNC|Hand left X-ray Brewerton|Hand left X-ray Brewerton
C0801762|T102|relax|38775-3|LNC|Hand right X-ray Brewerton|Hand right X-ray Brewerton
C0801762|T102|relax|37928-9|LNC|Wrist X-ray Brewerton|Wrist X-ray Brewerton
C0801762|T102|relax|37857-0|LNC|Sinuses X-ray Caldwell|Sinuses X-ray Caldwell
C0801762|T102|relax|69132-9|LNC|Hip X-ray Danelius Miller|Hip X-ray Danelius Miller
C0801762|T102|relax|69141-0|LNC|Hip left X-ray Danelius Miller|Hip left X-ray Danelius Miller
C0801762|T102|relax|39514-5|LNC|Hip right X-ray Danelius Miller|Hip right X-ray Danelius Miller
C0801762|T102|relax|37625-1|LNC|Pelvis X-ray Ferguson|Pelvis X-ray Ferguson
C0801762|T102|relax|37650-9|LNC|Sacroiliac Joint X-ray Ferguson|Sacroiliac Joint X-ray Ferguson
C0801762|T102|relax|65799-9|LNC|Kidney bilateral Fluoroscopy View cyst examination|Kidney bilateral Fluoroscopy View cyst examination
C0801762|T102|relax|65800-5|LNC|Kidney left Fluoroscopy View cyst examination|Kidney left Fluoroscopy View cyst examination
C0801762|T102|relax|65801-3|LNC|Kidney right Fluoroscopy View cyst examination|Kidney right Fluoroscopy View cyst examination
C0801762|T102|relax|37297-9|LNC|Abdomen Fetus X-ray View fetal age|Abdomen Fetus X-ray View fetal age
C0801762|T102|relax|39149-0|LNC|Gastrointestinal system Respiratory system X-ray foreign body|Gastrointestinal system Respiratory system X-ray foreign body
C0801762|T102|relax|36973-6|LNC|Hip X-ray Friedman|Hip X-ray Friedman
C0801762|T102|relax|37843-0|LNC|Shoulder X-ray Garth|Shoulder X-ray Garth
C0801762|T102|relax|36974-4|LNC|Shoulder left X-ray Garth|Shoulder left X-ray Garth
C0801762|T102|relax|37801-8|LNC|Shoulder right X-ray Garth|Shoulder right X-ray Garth
C0801762|T102|relax|37844-8|LNC|Shoulder X-ray Grashey|Shoulder X-ray Grashey
C0801762|T102|relax|37035-3|LNC|Shoulder bilateral X-ray Grashey|Shoulder bilateral X-ray Grashey
C0801762|T102|relax|37473-6|LNC|Shoulder left X-ray Grashey|Shoulder left X-ray Grashey
C0801762|T102|relax|38805-8|LNC|Shoulder right X-ray Grashey|Shoulder right X-ray Grashey
C0801762|T102|relax|36975-1|LNC|Calcaneus bilateral X-ray Harris|Calcaneus bilateral X-ray Harris
C0801762|T102|relax|36977-7|LNC|Calcaneus left X-ray Harris|Calcaneus left X-ray Harris
C0801762|T102|relax|38776-1|LNC|Calcaneus right X-ray Harris|Calcaneus right X-ray Harris
C0801762|T102|relax|36976-9|LNC|Foot X-ray Harris|Foot X-ray Harris
C0801762|T102|relax|36978-5|LNC|Knee X-ray Holmblad|Knee X-ray Holmblad
C0801762|T102|relax|37628-5|LNC|Pelvis X-ray inlet|Pelvis X-ray inlet
C0801762|T102|relax|36979-3|LNC|Elbow X-ray Jones|Elbow X-ray Jones
C0801762|T102|relax|36980-1|LNC|Elbow left X-ray Jones|Elbow left X-ray Jones
C0801762|T102|relax|38777-9|LNC|Elbow right X-ray Jones|Elbow right X-ray Jones
C0801762|T102|relax|36981-9|LNC|Hip X-ray Judet|Hip X-ray Judet
C0801762|T102|relax|36982-7|LNC|Hip bilateral X-ray Judet|Hip bilateral X-ray Judet
C0801762|T102|relax|36983-5|LNC|Hip left X-ray Judet|Hip left X-ray Judet
C0801762|T102|relax|37732-5|LNC|Hip right X-ray Judet|Hip right X-ray Judet
C0801762|T102|relax|36620-3|LNC|Chest X-ray left anterior oblique|Chest X-ray left anterior oblique
C0801762|T102|relax|36591-6|LNC|Abdomen X-ray lateral|Abdomen X-ray lateral
C0801762|T102|relax|36592-4|LNC|Ankle X-ray lateral|Ankle X-ray lateral
C0801762|T102|relax|39051-8|LNC|Chest X-ray lateral|Chest X-ray lateral
C0801762|T102|relax|36593-2|LNC|Femur X-ray lateral|Femur X-ray lateral
C0801762|T102|relax|36594-0|LNC|Finger fifth X-ray lateral|Finger fifth X-ray lateral
C0801762|T102|relax|36595-7|LNC|Finger fourth X-ray lateral|Finger fourth X-ray lateral
C0801762|T102|relax|36596-5|LNC|Finger second X-ray lateral|Finger second X-ray lateral
C0801762|T102|relax|36597-3|LNC|Finger third X-ray lateral|Finger third X-ray lateral
C0801762|T102|relax|36598-1|LNC|Foot left X-ray lateral|Foot left X-ray lateral
C0801762|T102|relax|37703-6|LNC|Foot right X-ray lateral|Foot right X-ray lateral
C0801762|T102|relax|36599-9|LNC|Hand X-ray lateral|Hand X-ray lateral
C0801762|T102|relax|36600-5|LNC|Hand bilateral X-ray lateral|Hand bilateral X-ray lateral
C0801762|T102|relax|36601-3|LNC|Hand left X-ray lateral|Hand left X-ray lateral
C0801762|T102|relax|37712-7|LNC|Hand right X-ray lateral|Hand right X-ray lateral
C0801762|T102|relax|36602-1|LNC|Hip X-ray lateral|Hip X-ray lateral
C0801762|T102|relax|36603-9|LNC|Hip left X-ray lateral|Hip left X-ray lateral
C0801762|T102|relax|37730-9|LNC|Hip right X-ray lateral|Hip right X-ray lateral
C0801762|T102|relax|36604-7|LNC|Knee X-ray lateral|Knee X-ray lateral
C0801762|T102|relax|36605-4|LNC|Knee bilateral X-ray lateral|Knee bilateral X-ray lateral
C0801762|T102|relax|36606-2|LNC|Knee left X-ray lateral|Knee left X-ray lateral
C0801762|T102|relax|37751-5|LNC|Knee right X-ray lateral|Knee right X-ray lateral
C0801762|T102|relax|24843-5|LNC|Neck X-ray lateral|Neck X-ray lateral
C0801762|T102|relax|37629-3|LNC|Pelvis X-ray lateral|Pelvis X-ray lateral
C0801762|T102|relax|39053-4|LNC|Ribs X-ray lateral|Ribs X-ray lateral
C0801762|T102|relax|38857-9|LNC|Ribs left X-ray lateral|Ribs left X-ray lateral
C0801762|T102|relax|37784-6|LNC|Ribs right X-ray lateral|Ribs right X-ray lateral
C0801762|T102|relax|37858-8|LNC|Sinuses X-ray lateral|Sinuses X-ray lateral
C0801762|T102|relax|24920-1|LNC|Skull X-ray lateral|Skull X-ray lateral
C0801762|T102|relax|24943-3|LNC|Spine Cervical X-ray lateral|Spine Cervical X-ray lateral
C0801762|T102|relax|24969-8|LNC|Spine Lumbar X-ray lateral|Spine Lumbar X-ray lateral
C0801762|T102|relax|30756-1|LNC|Spine Thoracic X-ray lateral|Spine Thoracic X-ray lateral
C0801762|T102|relax|37891-9|LNC|Thumb X-ray lateral|Thumb X-ray lateral
C0801762|T102|relax|37893-5|LNC|Tibia Fibula X-ray lateral|Tibia Fibula X-ray lateral
C0801762|T102|relax|37930-5|LNC|Wrist X-ray lateral|Wrist X-ray lateral
C0801762|T102|relax|36984-3|LNC|Abdomen X-ray lateral crosstable|Abdomen X-ray lateral crosstable
C0801762|T102|relax|36985-0|LNC|Hip X-ray lateral crosstable|Hip X-ray lateral crosstable
C0801762|T102|relax|36986-8|LNC|Hip bilateral X-ray lateral crosstable|Hip bilateral X-ray lateral crosstable
C0801762|T102|relax|36987-6|LNC|Hip left X-ray lateral crosstable|Hip left X-ray lateral crosstable
C0801762|T102|relax|37727-5|LNC|Hip right X-ray lateral crosstable|Hip right X-ray lateral crosstable
C0801762|T102|relax|36988-4|LNC|Knee X-ray lateral crosstable|Knee X-ray lateral crosstable
C0801762|T102|relax|37872-9|LNC|Skull X-ray lateral crosstable|Skull X-ray lateral crosstable
C0801762|T102|relax|36989-2|LNC|Spine Cervical X-ray lateral crosstable|Spine Cervical X-ray lateral crosstable
C0801762|T102|relax|36990-0|LNC|Spine Lumbar X-ray lateral crosstable|Spine Lumbar X-ray lateral crosstable
C0801762|T102|relax|37903-2|LNC|Spine Thoracic X-ray lateral crosstable|Spine Thoracic X-ray lateral crosstable
C0801762|T102|relax|36991-8|LNC|Spine Cervical X-ray lateral crosstable portable|Spine Cervical X-ray lateral crosstable portable
C0801762|T102|relax|36992-6|LNC|Spine Lumbar X-ray lateral crosstable portable|Spine Lumbar X-ray lateral crosstable portable
C0801762|T102|relax|30786-8|LNC|Hip X-ray lateral frog|Hip X-ray lateral frog
C0801762|T102|relax|36993-4|LNC|Hip bilateral X-ray lateral frog|Hip bilateral X-ray lateral frog
C0801762|T102|relax|36994-2|LNC|Hip left X-ray lateral frog|Hip left X-ray lateral frog
C0801762|T102|relax|37729-1|LNC|Hip right X-ray lateral frog|Hip right X-ray lateral frog
C0801762|T102|relax|37626-9|LNC|Pelvis X-ray lateral frog|Pelvis X-ray lateral frog
C0801762|T102|relax|36999-1|LNC|Knee bilateral X-ray lateral hyperextension|Knee bilateral X-ray lateral hyperextension
C0801762|T102|relax|37000-7|LNC|Knee left X-ray lateral hyperextension|Knee left X-ray lateral hyperextension
C0801762|T102|relax|37750-7|LNC|Knee right X-ray lateral hyperextension|Knee right X-ray lateral hyperextension
C0801762|T102|relax|37909-9|LNC|Spine Thoracic X-ray lateral hyperextension|Spine Thoracic X-ray lateral hyperextension
C0801762|T102|relax|41774-1|LNC|Neck X-ray lateral portable|Neck X-ray lateral portable
C0801762|T102|relax|30757-9|LNC|Spine Thoracic X-ray lateral portable|Spine Thoracic X-ray lateral portable
C0801762|T102|relax|37515-4|LNC|Spine Lumbosacral Junction X-ray lateral spot|Spine Lumbosacral Junction X-ray lateral spot
C0801762|T102|relax|37516-2|LNC|Spine Lumbosacral Junction X-ray lateral spot standing|Spine Lumbosacral Junction X-ray lateral spot standing
C0801762|T102|relax|38066-7|LNC|Hip left X-ray lateral during surgery|Hip left X-ray lateral during surgery
C0801762|T102|relax|38819-9|LNC|Hip right X-ray lateral during surgery|Hip right X-ray lateral during surgery
C0801762|T102|relax|37001-5|LNC|Foot X-ray lateral standing|Foot X-ray lateral standing
C0801762|T102|relax|37002-3|LNC|Knee left X-ray lateral standing|Knee left X-ray lateral standing
C0801762|T102|relax|37754-9|LNC|Knee right X-ray lateral standing|Knee right X-ray lateral standing
C0801762|T102|relax|37003-1|LNC|Spine Lumbar X-ray lateral standing|Spine Lumbar X-ray lateral standing
C0801762|T102|relax|37910-7|LNC|Spine Thoracic X-ray lateral standing|Spine Thoracic X-ray lateral standing
C0801762|T102|relax|36997-5|LNC|Spine Cervical X-ray lateral W extension|Spine Cervical X-ray lateral W extension
C0801762|T102|relax|36971-0|LNC|Wrist left X-ray lateral W extension|Wrist left X-ray lateral W extension
C0801762|T102|relax|37833-1|LNC|Wrist right X-ray lateral W extension|Wrist right X-ray lateral W extension
C0801762|T102|relax|36998-3|LNC|Spine Cervical X-ray lateral W flexion|Spine Cervical X-ray lateral W flexion
C0801762|T102|relax|36972-8|LNC|Wrist left X-ray lateral W flexion|Wrist left X-ray lateral W flexion
C0801762|T102|relax|37834-9|LNC|Wrist right X-ray lateral W flexion|Wrist right X-ray lateral W flexion
C0801762|T102|relax|37004-9|LNC|Knee X-ray Laurin|Knee X-ray Laurin
C0801762|T102|relax|36995-9|LNC|Abdomen X-ray left lateral|Abdomen X-ray left lateral
C0801762|T102|relax|30737-1|LNC|Chest X-ray left lateral|Chest X-ray left lateral
C0801762|T102|relax|30738-9|LNC|Chest X-ray left lateral portable|Chest X-ray left lateral portable
C0801762|T102|relax|24639-7|LNC|Chest X-ray left lateral upright|Chest X-ray left lateral upright
C0801762|T102|relax|24638-9|LNC|Chest X-ray left lateral upright portable|Chest X-ray left lateral upright portable
C0801762|T102|relax|37008-0|LNC|Chest X-ray left oblique|Chest X-ray left oblique
C0801762|T102|relax|37009-8|LNC|Spine Lumbar X-ray left oblique|Spine Lumbar X-ray left oblique
C0801762|T102|relax|24641-3|LNC|Chest X-ray left oblique portable|Chest X-ray left oblique portable
C0801762|T102|relax|24640-5|LNC|Chest X-ray lordotic|Chest X-ray lordotic
C0801762|T102|relax|38069-1|LNC|Abdomen X-ray left posterior oblique|Abdomen X-ray left posterior oblique
C0801762|T102|relax|37005-6|LNC|Breast left Mammogram magnification|Breast left Mammogram magnification
C0801762|T102|relax|37773-9|LNC|Breast right Mammogram magnification|Breast right Mammogram magnification
C0801762|T102|relax|42441-6|LNC|Neck X-ray magnification|Neck X-ray magnification
C0801762|T102|relax|24801-3|LNC|Knee X-ray Merchants|Knee X-ray Merchants
C0801762|T102|relax|26283-2|LNC|Knee bilateral X-ray Merchants|Knee bilateral X-ray Merchants
C0801762|T102|relax|26284-0|LNC|Knee left X-ray Merchants|Knee left X-ray Merchants
C0801762|T102|relax|26285-7|LNC|Knee right X-ray Merchants|Knee right X-ray Merchants
C0801762|T102|relax|37006-4|LNC|Breast bilateral Mammogram MLO|Breast bilateral Mammogram MLO
C0801762|T102|relax|37007-2|LNC|Ankle X-ray Mortise|Ankle X-ray Mortise
C0801762|T102|relax|37475-1|LNC|Ankle left X-ray Mortise W manual stress|Ankle left X-ray Mortise W manual stress
C0801762|T102|relax|37671-5|LNC|Ankle right X-ray Mortise W manual stress|Ankle right X-ray Mortise W manual stress
C0801762|T102|relax|38067-5|LNC|Breast bilateral Mammogram nipple profile|Breast bilateral Mammogram nipple profile
C0801762|T102|relax|36607-0|LNC|Abdomen X-ray oblique single view|Abdomen X-ray oblique single view
C0801762|T102|relax|36609-6|LNC|Femur X-ray oblique single view|Femur X-ray oblique single view
C0801762|T102|relax|36610-4|LNC|Finger fifth X-ray oblique single view|Finger fifth X-ray oblique single view
C0801762|T102|relax|36611-2|LNC|Finger fourth X-ray oblique single view|Finger fourth X-ray oblique single view
C0801762|T102|relax|36612-0|LNC|Finger second X-ray oblique single view|Finger second X-ray oblique single view
C0801762|T102|relax|36613-8|LNC|Finger third X-ray oblique single view|Finger third X-ray oblique single view
C0801762|T102|relax|36614-6|LNC|Foot X-ray oblique single view|Foot X-ray oblique single view
C0801762|T102|relax|36615-3|LNC|Foot left X-ray oblique single view|Foot left X-ray oblique single view
C0801762|T102|relax|37704-4|LNC|Foot right X-ray oblique single view|Foot right X-ray oblique single view
C0801762|T102|relax|36616-1|LNC|Hand X-ray oblique single view|Hand X-ray oblique single view
C0801762|T102|relax|36617-9|LNC|Hip X-ray oblique single view|Hip X-ray oblique single view
C0801762|T102|relax|36618-7|LNC|Hip bilateral X-ray oblique single view|Hip bilateral X-ray oblique single view
C0801762|T102|relax|30778-5|LNC|Spine Lumbar X-ray oblique single view|Spine Lumbar X-ray oblique single view
C0801762|T102|relax|30758-7|LNC|Spine Thoracic X-ray oblique single view|Spine Thoracic X-ray oblique single view
C0801762|T102|relax|37892-7|LNC|Thumb X-ray oblique single view|Thumb X-ray oblique single view
C0801762|T102|relax|44178-2|LNC|Spine Lumbar X-ray oblique view (views W right bending W left bending)|Spine Lumbar X-ray oblique view (views W right bending W left bending)
C0801762|T102|relax|37545-1|LNC|Hip left X-ray oblique crosstable|Hip left X-ray oblique crosstable
C0801762|T102|relax|37728-3|LNC|Hip right X-ray oblique crosstable|Hip right X-ray oblique crosstable
C0801762|T102|relax|30759-5|LNC|Spine Thoracic X-ray oblique portable|Spine Thoracic X-ray oblique portable
C0801762|T102|relax|37631-9|LNC|Pelvis X-ray outlet|Pelvis X-ray outlet
C0801762|T102|relax|37845-5|LNC|Shoulder X-ray outlet|Shoulder X-ray outlet
C0801762|T102|relax|37012-2|LNC|Shoulder bilateral X-ray outlet|Shoulder bilateral X-ray outlet
C0801762|T102|relax|37013-0|LNC|Shoulder left X-ray outlet|Shoulder left X-ray outlet
C0801762|T102|relax|37802-6|LNC|Shoulder right X-ray outlet|Shoulder right X-ray outlet
C0801762|T102|relax|36621-1|LNC|Hand X-ray PA|Hand X-ray PA
C0801762|T102|relax|36622-9|LNC|Hand bilateral X-ray PA|Hand bilateral X-ray PA
C0801762|T102|relax|36623-7|LNC|Hand left X-ray PA|Hand left X-ray PA
C0801762|T102|relax|37714-3|LNC|Hand right X-ray PA|Hand right X-ray PA
C0801762|T102|relax|69270-7|LNC|Skull X-ray PA|Skull X-ray PA
C0801762|T102|relax|37931-3|LNC|Wrist X-ray PA|Wrist X-ray PA
C0801762|T102|relax|36624-5|LNC|Wrist bilateral X-ray PA|Wrist bilateral X-ray PA
C0801762|T102|relax|37015-5|LNC|Abdomen X-ray PA prone|Abdomen X-ray PA prone
C0801762|T102|relax|24648-8|LNC|Chest X-ray PA upright|Chest X-ray PA upright
C0801762|T102|relax|37014-8|LNC|Knee left X-ray PA standing|Knee left X-ray PA standing
C0801762|T102|relax|37755-6|LNC|Knee right X-ray PA standing|Knee right X-ray PA standing
C0801762|T102|relax|37477-7|LNC|Knee X-ray PA standing W 45 degree flexion|Knee X-ray PA standing W 45 degree flexion
C0801762|T102|relax|37476-9|LNC|Knee X-ray PA W 45 degree flexion|Knee X-ray PA W 45 degree flexion
C0801762|T102|relax|39324-9|LNC|Wrist left X-ray PA W clenched fist|Wrist left X-ray PA W clenched fist
C0801762|T102|relax|69263-2|LNC|Wrist right X-ray PA W clenched fist|Wrist right X-ray PA W clenched fist
C0801762|T102|relax|24828-6|LNC|Mandible X-ray panorex|Mandible X-ray panorex
C0801762|T102|relax|24871-6|LNC|Pelvis X-ray pelvimetry|Pelvis X-ray pelvimetry
C0801762|T102|relax|37998-2|LNC|Elbow X-ray radial head capitellar|Elbow X-ray radial head capitellar
C0801762|T102|relax|37999-0|LNC|Elbow bilateral X-ray radial head capitellar|Elbow bilateral X-ray radial head capitellar
C0801762|T102|relax|38000-6|LNC|Elbow left X-ray radial head capitellar|Elbow left X-ray radial head capitellar
C0801762|T102|relax|38006-3|LNC|Elbow right X-ray radial head capitellar|Elbow right X-ray radial head capitellar
C0801762|T102|relax|38068-3|LNC|Chest X-ray right anterior oblique|Chest X-ray right anterior oblique
C0801762|T102|relax|36996-7|LNC|Abdomen X-ray right lateral|Abdomen X-ray right lateral
C0801762|T102|relax|37010-6|LNC|Chest X-ray right oblique|Chest X-ray right oblique
C0801762|T102|relax|37011-4|LNC|Spine Lumbar X-ray right oblique|Spine Lumbar X-ray right oblique
C0801762|T102|relax|37018-9|LNC|Knee X-ray Rosenberg standing|Knee X-ray Rosenberg standing
C0801762|T102|relax|37020-5|LNC|Knee bilateral X-ray Rosenberg standing|Knee bilateral X-ray Rosenberg standing
C0801762|T102|relax|37019-7|LNC|Knee left X-ray Rosenberg standing|Knee left X-ray Rosenberg standing
C0801762|T102|relax|37752-3|LNC|Knee right X-ray Rosenberg standing|Knee right X-ray Rosenberg standing
C0801762|T102|relax|39323-1|LNC|Abdomen X-ray right posterior oblique|Abdomen X-ray right posterior oblique
C0801762|T102|relax|49511-9|LNC|Femoral artery Fluoroscopic angiogram runoff W WO contrast IA|Femoral artery Fluoroscopic angiogram runoff W WO contrast IA
C0801762|T102|relax|24699-1|LNC|Femoral artery Fluoroscopic angiogram runoff W contrast IA|Femoral artery Fluoroscopic angiogram runoff W contrast IA
C0801762|T102|relax|26178-4|LNC|Femoral artery bilateral Fluoroscopic angiogram runoff W contrast IA|Femoral artery bilateral Fluoroscopic angiogram runoff W contrast IA
C0801762|T102|relax|26179-2|LNC|Femoral artery left Fluoroscopic angiogram runoff W contrast IA|Femoral artery left Fluoroscopic angiogram runoff W contrast IA
C0801762|T102|relax|26180-0|LNC|Femoral artery right Fluoroscopic angiogram runoff W contrast IA|Femoral artery right Fluoroscopic angiogram runoff W contrast IA
C0801762|T102|relax|42812-8|LNC|Wrist X-ray scaphoid single view|Wrist X-ray scaphoid single view
C0801762|T102|relax|42813-6|LNC|Wrist bilateral X-ray scaphoid single view|Wrist bilateral X-ray scaphoid single view
C0801762|T102|relax|42814-4|LNC|Wrist left X-ray scaphoid single view|Wrist left X-ray scaphoid single view
C0801762|T102|relax|42811-0|LNC|Wrist right X-ray scaphoid single view|Wrist right X-ray scaphoid single view
C0801762|T102|relax|44206-1|LNC|Spine Thoracic Lumbar X-ray scoliosis single view|Spine Thoracic Lumbar X-ray scoliosis single view
C0801762|T102|relax|30714-0|LNC|Spine Thoracic Lumbar X-ray scoliosis AP|Spine Thoracic Lumbar X-ray scoliosis AP
C0801762|T102|relax|42426-7|LNC|Spine Thoracic Lumbar X-ray scoliosis AP sitting|Spine Thoracic Lumbar X-ray scoliosis AP sitting
C0801762|T102|relax|37659-0|LNC|Spine Thoracic Lumbar X-ray scoliosis AP standing|Spine Thoracic Lumbar X-ray scoliosis AP standing
C0801762|T102|relax|42428-3|LNC|Spine Thoracic Lumbar X-ray scoliosis AP standing in brace|Spine Thoracic Lumbar X-ray scoliosis AP standing in brace
C0801762|T102|relax|42429-1|LNC|Spine Thoracic Lumbar X-ray scoliosis AP standing W right bending|Spine Thoracic Lumbar X-ray scoliosis AP standing W right bending
C0801762|T102|relax|42427-5|LNC|Spine Thoracic Lumbar X-ray scoliosis lateral sitting|Spine Thoracic Lumbar X-ray scoliosis lateral sitting
C0801762|T102|relax|37660-8|LNC|Spine Thoracic Lumbar X-ray scoliosis lateral standing|Spine Thoracic Lumbar X-ray scoliosis lateral standing
C0801762|T102|relax|37846-3|LNC|Sternoclavicular Joint X-ray Serendipity|Sternoclavicular Joint X-ray Serendipity
C0801762|T102|relax|37298-7|LNC|Sternoclavicular joint bilateral X-ray Serendipity|Sternoclavicular joint bilateral X-ray Serendipity
C0801762|T102|relax|37299-5|LNC|Sternoclavicular joint left X-ray Serendipity|Sternoclavicular joint left X-ray Serendipity
C0801762|T102|relax|37808-3|LNC|Sternoclavicular joint right X-ray Serendipity|Sternoclavicular joint right X-ray Serendipity
C0801762|T102|relax|43671-7|LNC|Thyroid Scan spot|Thyroid Scan spot
C0801762|T102|relax|42471-3|LNC|Pelvis X-ray stereo|Pelvis X-ray stereo
C0801762|T102|relax|42474-7|LNC|Skull X-ray stereo|Skull X-ray stereo
C0801762|T102|relax|39516-0|LNC|Shoulder X-ray Stryker Notch|Shoulder X-ray Stryker Notch
C0801762|T102|relax|37024-7|LNC|Shoulder bilateral X-ray Stryker Notch|Shoulder bilateral X-ray Stryker Notch
C0801762|T102|relax|37025-4|LNC|Shoulder left X-ray Stryker Notch|Shoulder left X-ray Stryker Notch
C0801762|T102|relax|37791-1|LNC|Shoulder right X-ray Stryker Notch|Shoulder right X-ray Stryker Notch
C0801762|T102|relax|39517-8|LNC|Shoulder X-ray Stryker Notch West Point|Shoulder X-ray Stryker Notch West Point
C0801762|T102|relax|37861-2|LNC|Sinuses X-ray submentovertex|Sinuses X-ray submentovertex
C0801762|T102|relax|37026-2|LNC|Skull X-ray submentovertex|Skull X-ray submentovertex
C0801762|T102|relax|43780-6|LNC|Knee X-ray Sunrise|Knee X-ray Sunrise
C0801762|T102|relax|37027-0|LNC|Knee bilateral X-ray Sunrise|Knee bilateral X-ray Sunrise
C0801762|T102|relax|43779-8|LNC|Knee left X-ray Sunrise|Knee left X-ray Sunrise
C0801762|T102|relax|69256-6|LNC|Knee right X-ray Sunrise|Knee right X-ray Sunrise
C0801762|T102|relax|69239-2|LNC|Patella X-ray Sunrise|Patella X-ray Sunrise
C0801762|T102|relax|69069-3|LNC|Patella bilateral X-ray Sunrise|Patella bilateral X-ray Sunrise
C0801762|T102|relax|69064-4|LNC|Knee bilateral X-ray Sunrise (views standing)|Knee bilateral X-ray Sunrise (views standing)
C0801762|T102|relax|69149-3|LNC|Knee left X-ray Sunrise (views standing)|Knee left X-ray Sunrise (views standing)
C0801762|T102|relax|42432-5|LNC|Knee right X-ray Sunrise (views standing)|Knee right X-ray Sunrise (views standing)
C0801762|T102|relax|24944-1|LNC|Spine Cervical X-ray Swimmers|Spine Cervical X-ray Swimmers
C0801762|T102|relax|37028-8|LNC|Breast Mammogram tangential|Breast Mammogram tangential
C0801762|T102|relax|37029-6|LNC|Breast bilateral Mammogram tangential|Breast bilateral Mammogram tangential
C0801762|T102|relax|37030-4|LNC|Breast left Mammogram tangential|Breast left Mammogram tangential
C0801762|T102|relax|37770-5|LNC|Breast right Mammogram tangential|Breast right Mammogram tangential
C0801762|T102|relax|37870-3|LNC|Skull X-ray Towne|Skull X-ray Towne
C0801762|T102|relax|24668-6|LNC|Colon Fluoroscopy transit Post solid contrast|Colon Fluoroscopy transit Post solid contrast
C0801762|T102|relax|37031-2|LNC|Humerus X-ray transthoracic|Humerus X-ray transthoracic
C0801762|T102|relax|37032-0|LNC|Humerus bilateral X-ray transthoracic|Humerus bilateral X-ray transthoracic
C0801762|T102|relax|37033-8|LNC|Humerus left X-ray transthoracic|Humerus left X-ray transthoracic
C0801762|T102|relax|38007-1|LNC|Humerus right X-ray transthoracic|Humerus right X-ray transthoracic
C0801762|T102|relax|37034-6|LNC|Shoulder left X-ray transthoracic|Shoulder left X-ray transthoracic
C0801762|T102|relax|38779-5|LNC|Shoulder right X-ray transthoracic|Shoulder right X-ray transthoracic
C0801762|T102|relax|37300-1|LNC|Spine Lumbosacral Junction X-ray true AP|Spine Lumbosacral Junction X-ray true AP
C0801762|T102|relax|37037-9|LNC|Breast Mammogram true lateral|Breast Mammogram true lateral
C0801762|T102|relax|37038-7|LNC|Breast bilateral Mammogram true lateral|Breast bilateral Mammogram true lateral
C0801762|T102|relax|38855-3|LNC|Breast left Mammogram true lateral|Breast left Mammogram true lateral
C0801762|T102|relax|37771-3|LNC|Breast right Mammogram true lateral|Breast right Mammogram true lateral
C0801762|T102|relax|37039-5|LNC|Hip X-ray true lateral|Hip X-ray true lateral
C0801762|T102|relax|37040-3|LNC|Hip left X-ray true lateral|Hip left X-ray true lateral
C0801762|T102|relax|38772-0|LNC|Hip right X-ray true lateral|Hip right X-ray true lateral
C0801762|T102|relax|30790-0|LNC|Knee X-ray tunnel|Knee X-ray tunnel
C0801762|T102|relax|37041-1|LNC|Knee bilateral X-ray tunnel|Knee bilateral X-ray tunnel
C0801762|T102|relax|37042-9|LNC|Knee left X-ray tunnel|Knee left X-ray tunnel
C0801762|T102|relax|37761-4|LNC|Knee right X-ray tunnel|Knee right X-ray tunnel
C0801762|T102|relax|38842-1|LNC|Wrist left X-ray tunnel carpal|Wrist left X-ray tunnel carpal
C0801762|T102|relax|37677-2|LNC|Wrist right X-ray tunnel carpal|Wrist right X-ray tunnel carpal
C0801762|T102|relax|37043-7|LNC|Knee left X-ray tunnel standing|Knee left X-ray tunnel standing
C0801762|T102|relax|37756-4|LNC|Knee right X-ray tunnel standing|Knee right X-ray tunnel standing
C0801762|T102|relax|37044-5|LNC|Wrist left X-ray ulnar deviation|Wrist left X-ray ulnar deviation
C0801762|T102|relax|37645-9|LNC|Wrist right X-ray ulnar deviation|Wrist right X-ray ulnar deviation
C0801762|T102|relax|37045-2|LNC|Wrist bilateral X-ray ulnar variance|Wrist bilateral X-ray ulnar variance
C0801762|T102|relax|37046-0|LNC|Abdomen X-ray upright|Abdomen X-ray upright
C0801762|T102|relax|37047-8|LNC|Shoulder bilateral X-ray Velpeau axillary|Shoulder bilateral X-ray Velpeau axillary
C0801762|T102|relax|37048-6|LNC|Shoulder left X-ray Velpeau axillary|Shoulder left X-ray Velpeau axillary
C0801762|T102|relax|38780-3|LNC|Shoulder right X-ray Velpeau axillary|Shoulder right X-ray Velpeau axillary
C0801762|T102|relax|37049-4|LNC|Hip X-ray Von rossen|Hip X-ray Von rossen
C0801762|T102|relax|37613-7|LNC|Orbit bilateral X-ray Waters|Orbit bilateral X-ray Waters
C0801762|T102|relax|37863-8|LNC|Sinuses X-ray Waters|Sinuses X-ray Waters
C0801762|T102|relax|24921-9|LNC|Skull X-ray Waters|Skull X-ray Waters
C0801762|T102|relax|42473-9|LNC|Sinuses X-ray Waters stereo|Sinuses X-ray Waters stereo
C0801762|T102|relax|38117-8|LNC|Sinuses X-ray Waters upright|Sinuses X-ray Waters upright
C0801762|T102|relax|30751-2|LNC|Shoulder X-ray West Point|Shoulder X-ray West Point
C0801762|T102|relax|37050-2|LNC|Shoulder bilateral X-ray West Point|Shoulder bilateral X-ray West Point
C0801762|T102|relax|37051-0|LNC|Shoulder left X-ray West Point|Shoulder left X-ray West Point
C0801762|T102|relax|37809-1|LNC|Shoulder right X-ray West Point|Shoulder right X-ray West Point
C0801762|T102|relax|42680-9|LNC|Breast Mammogram XCCL|Breast Mammogram XCCL
C0801762|T102|relax|37052-8|LNC|Breast bilateral Mammogram XCCL|Breast bilateral Mammogram XCCL
C0801762|T102|relax|37053-6|LNC|Breast left Mammogram XCCL|Breast left Mammogram XCCL
C0801762|T102|relax|37772-1|LNC|Breast right Mammogram XCCL|Breast right Mammogram XCCL
C0801762|T102|relax|37656-6|LNC|Scapula X-ray Y|Scapula X-ray Y
C0801762|T102|relax|37055-1|LNC|Scapula bilateral X-ray Y|Scapula bilateral X-ray Y
C0801762|T102|relax|37054-4|LNC|Scapula left X-ray Y|Scapula left X-ray Y
C0801762|T102|relax|37790-3|LNC|Scapula right X-ray Y|Scapula right X-ray Y
C0801762|T102|relax|37847-1|LNC|Shoulder X-ray Y|Shoulder X-ray Y
C0801762|T102|relax|38858-7|LNC|Shoulder left X-ray Y|Shoulder left X-ray Y
C0801762|T102|relax|37805-9|LNC|Shoulder right X-ray Y|Shoulder right X-ray Y
C0801762|T102|relax|37848-9|LNC|Acromioclavicular Joint X-ray Zanca|Acromioclavicular Joint X-ray Zanca
C0801762|T102|relax|37056-9|LNC|Acromioclavicular joint bilateral X-ray Zanca|Acromioclavicular joint bilateral X-ray Zanca
C0801762|T102|relax|37057-7|LNC|Acromioclavicular joint left X-ray Zanca|Acromioclavicular joint left X-ray Zanca
C0801762|T102|relax|37810-9|LNC|Acromioclavicular joint right X-ray Zanca|Acromioclavicular joint right X-ray Zanca
C0801762|T102|relax|41793-1|LNC|Abdomen X-ray during surgery|Abdomen X-ray during surgery
C0801762|T102|relax|41790-7|LNC|Chest X-ray during surgery|Chest X-ray during surgery
C0801762|T102|relax|24656-1|LNC|Chest Fluoroscopy during surgery|Chest Fluoroscopy during surgery
C0801762|T102|relax|39047-6|LNC|Hip Fluoroscopy during surgery|Hip Fluoroscopy during surgery
C0801762|T102|relax|38065-9|LNC|Hip left X-ray during surgery|Hip left X-ray during surgery
C0801762|T102|relax|38818-1|LNC|Hip right X-ray during surgery|Hip right X-ray during surgery
C0801762|T102|relax|42008-3|LNC|Humerus X-ray during surgery|Humerus X-ray during surgery
C0801762|T102|relax|24893-0|LNC|Rectum Fluoroscopy post contrast PR during defecation|Rectum Fluoroscopy post contrast PR during defecation
C0801762|T102|relax|37058-5|LNC|Calcaneus bilateral X-ray standing|Calcaneus bilateral X-ray standing
C0801762|T102|relax|37059-3|LNC|Hip bilateral X-ray standing|Hip bilateral X-ray standing
C0801762|T102|relax|37207-8|LNC|Hip left X-ray standing|Hip left X-ray standing
C0801762|T102|relax|37731-7|LNC|Hip right X-ray standing|Hip right X-ray standing
C0801762|T102|relax|44205-3|LNC|Lower extremity bilateral X-ray standing|Lower extremity bilateral X-ray standing
C0801762|T102|relax|38850-4|LNC|Lower extremity left X-ray standing|Lower extremity left X-ray standing
C0801762|T102|relax|37734-1|LNC|Lower extremity right X-ray standing|Lower extremity right X-ray standing
C0801762|T102|relax|37633-5|LNC|Pelvis X-ray standing|Pelvis X-ray standing
C0801762|T102|relax|39144-1|LNC|Gastrointestine upper Fluoroscopy W air contrast PO|Gastrointestine upper Fluoroscopy W air contrast PO
C0801762|T102|relax|69302-8|LNC|Wrist X-ray W clenched fist|Wrist X-ray W clenched fist
C0801762|T102|relax|36968-6|LNC|Wrist bilateral X-ray W clenched fist|Wrist bilateral X-ray W clenched fist
C0801762|T102|relax|30639-9|LNC|Vessel Fluoroscopic angiogram W contrast|Vessel Fluoroscopic angiogram W contrast
C0801762|T102|relax|42470-5|LNC|Gastrointestine upper Gallbladder Fluoroscopy W contrast PO|Gastrointestine upper Gallbladder Fluoroscopy W contrast PO
C0801762|T102|relax|30809-8|LNC|Upper Gastrointestine Small bowel Fluoroscopy W contrast PO|Upper Gastrointestine Small bowel Fluoroscopy W contrast PO
C0801762|T102|relax|42469-7|LNC|Gastrointestine upper Small bowel Gallbladder Fluoroscopy W contrast PO|Gastrointestine upper Small bowel Gallbladder Fluoroscopy W contrast PO
C0801762|T102|relax|38001-4|LNC|Chest X-ray W expiration|Chest X-ray W expiration
C0801762|T102|relax|38002-2|LNC|Chest X-ray W inspiration|Chest X-ray W inspiration
C0801762|T102|relax|37060-1|LNC|Fetal X-ray|Fetal X-ray
C0801762|T102|relax|37636-8|LNC|Abdomen X-ray|Abdomen X-ray
C0801762|T102|relax|46341-4|LNC|Abdomen Fluoroscopy|Abdomen Fluoroscopy
C0801762|T102|relax|24535-7|LNC|Acetabulum X-ray|Acetabulum X-ray
C0801762|T102|relax|26133-9|LNC|Acetabulum bilateral X-ray|Acetabulum bilateral X-ray
C0801762|T102|relax|26134-7|LNC|Acetabulum left X-ray|Acetabulum left X-ray
C0801762|T102|relax|26135-4|LNC|Acetabulum right X-ray|Acetabulum right X-ray
C0801762|T102|relax|24536-5|LNC|Acromioclavicular Joint X-ray|Acromioclavicular Joint X-ray
C0801762|T102|relax|26136-2|LNC|Acromioclavicular joint bilateral X-ray|Acromioclavicular joint bilateral X-ray
C0801762|T102|relax|26137-0|LNC|Acromioclavicular joint left X-ray|Acromioclavicular joint left X-ray
C0801762|T102|relax|26138-8|LNC|Acromioclavicular joint right X-ray|Acromioclavicular joint right X-ray
C0801762|T102|relax|24541-5|LNC|Ankle X-ray|Ankle X-ray
C0801762|T102|relax|26097-6|LNC|Ankle bilateral X-ray|Ankle bilateral X-ray
C0801762|T102|relax|26098-4|LNC|Ankle left X-ray|Ankle left X-ray
C0801762|T102|relax|51395-2|LNC|Ankle left Foot left X-ray|Ankle left Foot left X-ray
C0801762|T102|relax|26099-2|LNC|Ankle right X-ray|Ankle right X-ray
C0801762|T102|relax|51394-5|LNC|Ankle right Foot right X-ray|Ankle right Foot right X-ray
C0801762|T102|relax|36625-2|LNC|Breast Mammogram|Breast Mammogram
C0801762|T102|relax|46342-2|LNC|Breast FFD mammogram|Breast FFD mammogram
C0801762|T102|relax|38070-9|LNC|Breast implant Mammogram|Breast implant Mammogram
C0801762|T102|relax|38071-7|LNC|Breast implant bilateral Mammogram|Breast implant bilateral Mammogram
C0801762|T102|relax|38072-5|LNC|Breast implant left Mammogram|Breast implant left Mammogram
C0801762|T102|relax|38820-7|LNC|Breast implant right Mammogram|Breast implant right Mammogram
C0801762|T102|relax|46380-2|LNC|Breast Implant unilateral Mammogram|Breast Implant unilateral Mammogram
C0801762|T102|relax|24597-7|LNC|Breast specimen Mammogram|Breast specimen Mammogram
C0801762|T102|relax|38079-0|LNC|Breast specimen bilateral Mammogram|Breast specimen bilateral Mammogram
C0801762|T102|relax|38080-8|LNC|Breast specimen left Mammogram|Breast specimen left Mammogram
C0801762|T102|relax|38821-5|LNC|Breast specimen right Mammogram|Breast specimen right Mammogram
C0801762|T102|relax|36626-0|LNC|Breast bilateral Mammogram|Breast bilateral Mammogram
C0801762|T102|relax|36627-8|LNC|Breast left Mammogram|Breast left Mammogram
C0801762|T102|relax|37774-7|LNC|Breast right Mammogram|Breast right Mammogram
C0801762|T102|relax|46339-8|LNC|Breast unilateral Mammogram|Breast unilateral Mammogram
C0801762|T102|relax|24612-4|LNC|Calcaneus X-ray|Calcaneus X-ray
C0801762|T102|relax|26100-8|LNC|Calcaneus bilateral X-ray|Calcaneus bilateral X-ray
C0801762|T102|relax|26101-6|LNC|Calcaneus left X-ray|Calcaneus left X-ray
C0801762|T102|relax|26102-4|LNC|Calcaneus right X-ray|Calcaneus right X-ray
C0801762|T102|relax|30745-4|LNC|Chest X-ray|Chest X-ray
C0801762|T102|relax|30631-6|LNC|Chest Fluoroscopy|Chest Fluoroscopy
C0801762|T102|relax|42269-1|LNC|Chest Abdomen X-ray|Chest Abdomen X-ray
C0801762|T102|relax|24664-5|LNC|Clavicle X-ray|Clavicle X-ray
C0801762|T102|relax|26106-5|LNC|Clavicle bilateral X-ray|Clavicle bilateral X-ray
C0801762|T102|relax|26107-3|LNC|Clavicle left X-ray|Clavicle left X-ray
C0801762|T102|relax|26108-1|LNC|Clavicle right X-ray|Clavicle right X-ray
C0801762|T102|relax|30883-3|LNC|Coccyx X-ray|Coccyx X-ray
C0801762|T102|relax|24676-9|LNC|Elbow X-ray|Elbow X-ray
C0801762|T102|relax|26109-9|LNC|Elbow bilateral X-ray|Elbow bilateral X-ray
C0801762|T102|relax|26110-7|LNC|Elbow left X-ray|Elbow left X-ray
C0801762|T102|relax|26111-5|LNC|Elbow right X-ray|Elbow right X-ray
C0801762|T102|relax|46381-0|LNC|Elbow+Radius+Ulna X-ray|Elbow+Radius+Ulna X-ray
C0801762|T102|relax|37637-6|LNC|Extremity X-ray|Extremity X-ray
C0801762|T102|relax|24695-9|LNC|Facial bones X-ray|Facial bones X-ray
C0801762|T102|relax|37303-5|LNC|Facial bones Zygomatic arch X-ray|Facial bones Zygomatic arch X-ray
C0801762|T102|relax|24704-9|LNC|Femur X-ray|Femur X-ray
C0801762|T102|relax|26118-0|LNC|Femur bilateral X-ray|Femur bilateral X-ray
C0801762|T102|relax|26120-6|LNC|Femur left X-ray|Femur left X-ray
C0801762|T102|relax|26122-2|LNC|Femur right X-ray|Femur right X-ray
C0801762|T102|relax|24706-4|LNC|Finger X-ray|Finger X-ray
C0801762|T102|relax|26124-8|LNC|Finger bilateral X-ray|Finger bilateral X-ray
C0801762|T102|relax|30783-5|LNC|Finger fifth X-ray|Finger fifth X-ray
C0801762|T102|relax|37517-0|LNC|Finger fifth bilateral X-ray|Finger fifth bilateral X-ray
C0801762|T102|relax|37518-8|LNC|Finger fifth left X-ray|Finger fifth left X-ray
C0801762|T102|relax|38147-5|LNC|Finger fifth right X-ray|Finger fifth right X-ray
C0801762|T102|relax|30782-7|LNC|Finger fourth X-ray|Finger fourth X-ray
C0801762|T102|relax|37519-6|LNC|Finger fourth bilateral X-ray|Finger fourth bilateral X-ray
C0801762|T102|relax|37520-4|LNC|Finger fourth left X-ray|Finger fourth left X-ray
C0801762|T102|relax|38146-7|LNC|Finger fourth right X-ray|Finger fourth right X-ray
C0801762|T102|relax|26125-5|LNC|Finger left X-ray|Finger left X-ray
C0801762|T102|relax|26126-3|LNC|Finger right X-ray|Finger right X-ray
C0801762|T102|relax|30780-1|LNC|Finger second X-ray|Finger second X-ray
C0801762|T102|relax|37521-2|LNC|Finger second bilateral X-ray|Finger second bilateral X-ray
C0801762|T102|relax|37522-0|LNC|Finger second left X-ray|Finger second left X-ray
C0801762|T102|relax|38144-2|LNC|Finger second right X-ray|Finger second right X-ray
C0801762|T102|relax|30781-9|LNC|Finger third X-ray|Finger third X-ray
C0801762|T102|relax|37523-8|LNC|Finger third bilateral X-ray|Finger third bilateral X-ray
C0801762|T102|relax|37524-6|LNC|Finger third left X-ray|Finger third left X-ray
C0801762|T102|relax|38145-9|LNC|Finger third right X-ray|Finger third right X-ray
C0801762|T102|relax|24709-8|LNC|Foot X-ray|Foot X-ray
C0801762|T102|relax|26127-1|LNC|Foot bilateral X-ray|Foot bilateral X-ray
C0801762|T102|relax|26128-9|LNC|Foot left X-ray|Foot left X-ray
C0801762|T102|relax|26129-7|LNC|Foot right X-ray|Foot right X-ray
C0801762|T102|relax|42399-6|LNC|Foot sesamoid bones X-ray|Foot sesamoid bones X-ray
C0801762|T102|relax|42400-2|LNC|Foot sesamoid bones bilateral X-ray|Foot sesamoid bones bilateral X-ray
C0801762|T102|relax|43641-0|LNC|Foot sesamoid bones left X-ray|Foot sesamoid bones left X-ray
C0801762|T102|relax|42434-1|LNC|Foot sesamoid bones right X-ray|Foot sesamoid bones right X-ray
C0801762|T102|relax|37532-9|LNC|Great toe bilateral X-ray|Great toe bilateral X-ray
C0801762|T102|relax|37533-7|LNC|Great toe left X-ray|Great toe left X-ray
C0801762|T102|relax|38152-5|LNC|Great toe right X-ray|Great toe right X-ray
C0801762|T102|relax|28582-5|LNC|Hand X-ray|Hand X-ray
C0801762|T102|relax|36629-4|LNC|Hand bilateral X-ray|Hand bilateral X-ray
C0801762|T102|relax|36630-2|LNC|Hand left X-ray|Hand left X-ray
C0801762|T102|relax|37716-8|LNC|Hand right X-ray|Hand right X-ray
C0801762|T102|relax|24752-8|LNC|Heart Fluoroscopy video|Heart Fluoroscopy video
C0801762|T102|relax|24762-7|LNC|Hip X-ray|Hip X-ray
C0801762|T102|relax|26130-5|LNC|Hip bilateral X-ray|Hip bilateral X-ray
C0801762|T102|relax|26131-3|LNC|Hip left X-ray|Hip left X-ray
C0801762|T102|relax|26132-1|LNC|Hip right X-ray|Hip right X-ray
C0801762|T102|relax|28567-6|LNC|Humerus X-ray|Humerus X-ray
C0801762|T102|relax|37319-1|LNC|Humerus bicipital groove X-ray|Humerus bicipital groove X-ray
C0801762|T102|relax|37321-7|LNC|Humerus bicipital groove bilateral X-ray|Humerus bicipital groove bilateral X-ray
C0801762|T102|relax|37320-9|LNC|Humerus bicipital groove left X-ray|Humerus bicipital groove left X-ray
C0801762|T102|relax|38797-7|LNC|Humerus bicipital groove right X-ray|Humerus bicipital groove right X-ray
C0801762|T102|relax|37062-7|LNC|Humerus bilateral X-ray|Humerus bilateral X-ray
C0801762|T102|relax|36632-8|LNC|Humerus left X-ray|Humerus left X-ray
C0801762|T102|relax|37738-2|LNC|Humerus right X-ray|Humerus right X-ray
C0801762|T102|relax|36628-6|LNC|Internal auditory canal X-ray|Internal auditory canal X-ray
C0801762|T102|relax|28565-0|LNC|Knee X-ray|Knee X-ray
C0801762|T102|relax|36635-1|LNC|Knee bilateral X-ray|Knee bilateral X-ray
C0801762|T102|relax|36636-9|LNC|Knee left X-ray|Knee left X-ray
C0801762|T102|relax|37758-0|LNC|Knee right X-ray|Knee right X-ray
C0801762|T102|relax|48465-9|LNC|Larynx Fluoroscopy|Larynx Fluoroscopy
C0801762|T102|relax|24686-8|LNC|Lower extremity X-ray|Lower extremity X-ray
C0801762|T102|relax|26112-3|LNC|Lower extremity bilateral X-ray|Lower extremity bilateral X-ray
C0801762|T102|relax|26113-1|LNC|Lower extremity left X-ray|Lower extremity left X-ray
C0801762|T102|relax|26114-9|LNC|Lower extremity right X-ray|Lower extremity right X-ray
C0801762|T102|relax|24829-4|LNC|Mandible X-ray|Mandible X-ray
C0801762|T102|relax|48745-4|LNC|Mandible left X-ray|Mandible left X-ray
C0801762|T102|relax|43533-9|LNC|Mandible right X-ray|Mandible right X-ray
C0801762|T102|relax|24830-2|LNC|Mastoid X-ray|Mastoid X-ray
C0801762|T102|relax|26139-6|LNC|Mastoid bilateral X-ray|Mastoid bilateral X-ray
C0801762|T102|relax|26140-4|LNC|Mastoid left X-ray|Mastoid left X-ray
C0801762|T102|relax|26141-2|LNC|Mastoid right X-ray|Mastoid right X-ray
C0801762|T102|relax|36637-7|LNC|Maxilla X-ray|Maxilla X-ray
C0801762|T102|relax|24834-4|LNC|Nasal bones X-ray|Nasal bones X-ray
C0801762|T102|relax|37639-2|LNC|Neck X-ray|Neck X-ray
C0801762|T102|relax|37332-4|LNC|Olecranon left X-ray|Olecranon left X-ray
C0801762|T102|relax|38798-5|LNC|Olecranon right X-ray|Olecranon right X-ray
C0801762|T102|relax|24846-8|LNC|Optic foramen X-ray|Optic foramen X-ray
C0801762|T102|relax|26142-0|LNC|Optic foramen bilateral X-ray|Optic foramen bilateral X-ray
C0801762|T102|relax|26143-8|LNC|Optic foramen left X-ray|Optic foramen left X-ray
C0801762|T102|relax|26144-6|LNC|Optic foramen right X-ray|Optic foramen right X-ray
C0801762|T102|relax|36886-0|LNC|Orbit X-ray|Orbit X-ray
C0801762|T102|relax|24854-2|LNC|Orbit bilateral X-ray|Orbit bilateral X-ray
C0801762|T102|relax|36887-8|LNC|Orbit left X-ray|Orbit left X-ray
C0801762|T102|relax|38774-6|LNC|Orbit right X-ray|Orbit right X-ray
C0801762|T102|relax|43529-7|LNC|Orbit + Facial bones X-ray|Orbit + Facial bones X-ray
C0801762|T102|relax|24855-9|LNC|Oropharynx Fluoroscopy video|Oropharynx Fluoroscopy video
C0801762|T102|relax|30791-8|LNC|Patella X-ray|Patella X-ray
C0801762|T102|relax|36638-5|LNC|Patella bilateral X-ray|Patella bilateral X-ray
C0801762|T102|relax|36639-3|LNC|Patella left X-ray|Patella left X-ray
C0801762|T102|relax|37777-0|LNC|Patella right X-ray|Patella right X-ray
C0801762|T102|relax|28561-9|LNC|Pelvis X-ray|Pelvis X-ray
C0801762|T102|relax|30885-8|LNC|Pelvis symphysis pubis X-ray|Pelvis symphysis pubis X-ray
C0801762|T102|relax|30767-8|LNC|Pelvis Hip X-ray|Pelvis Hip X-ray
C0801762|T102|relax|30768-6|LNC|Pelvis Hip bilateral X-ray|Pelvis Hip bilateral X-ray
C0801762|T102|relax|36631-0|LNC|Pelvis Hip left X-ray|Pelvis Hip left X-ray
C0801762|T102|relax|38771-2|LNC|Pelvis Hip right X-ray|Pelvis Hip right X-ray
C0801762|T102|relax|47984-0|LNC|Pelvis Spine Lumbar X-ray|Pelvis Spine Lumbar X-ray
C0801762|T102|relax|24745-2|LNC|Petrous bone X-ray|Petrous bone X-ray
C0801762|T102|relax|26146-1|LNC|Radius bilateral Ulna bilateral X-ray|Radius bilateral Ulna bilateral X-ray
C0801762|T102|relax|26148-7|LNC|Radius left Ulna left X-ray|Radius left Ulna left X-ray
C0801762|T102|relax|26150-3|LNC|Radius right Ulna right X-ray|Radius right Ulna right X-ray
C0801762|T102|relax|24891-4|LNC|Radius Ulna X-ray|Radius Ulna X-ray
C0801762|T102|relax|24899-7|LNC|Ribs X-ray|Ribs X-ray
C0801762|T102|relax|37937-0|LNC|Ribs anterior X-ray|Ribs anterior X-ray
C0801762|T102|relax|38073-3|LNC|Ribs anterior bilateral X-ray|Ribs anterior bilateral X-ray
C0801762|T102|relax|38074-1|LNC|Ribs anterior left X-ray|Ribs anterior left X-ray
C0801762|T102|relax|37963-6|LNC|Ribs anterior right X-ray|Ribs anterior right X-ray
C0801762|T102|relax|38868-6|LNC|Ribs anterior posterior left X-ray|Ribs anterior posterior left X-ray
C0801762|T102|relax|37962-8|LNC|Ribs anterior posterior right X-ray|Ribs anterior posterior right X-ray
C0801762|T102|relax|26151-1|LNC|Ribs bilateral X-ray|Ribs bilateral X-ray
C0801762|T102|relax|69071-9|LNC|Ribs bilateral Chest X-ray|Ribs bilateral Chest X-ray
C0801762|T102|relax|26152-9|LNC|Ribs left X-ray|Ribs left X-ray
C0801762|T102|relax|39326-4|LNC|Ribs left Chest X-ray|Ribs left Chest X-ray
C0801762|T102|relax|38866-0|LNC|Ribs lower left X-ray|Ribs lower left X-ray
C0801762|T102|relax|39489-0|LNC|Ribs lower posterior X-ray|Ribs lower posterior X-ray
C0801762|T102|relax|42381-4|LNC|Ribs lower posterior left X-ray|Ribs lower posterior left X-ray
C0801762|T102|relax|39493-2|LNC|Ribs lower posterior right X-ray|Ribs lower posterior right X-ray
C0801762|T102|relax|37960-2|LNC|Ribs lower right X-ray|Ribs lower right X-ray
C0801762|T102|relax|37938-8|LNC|Ribs posterior X-ray|Ribs posterior X-ray
C0801762|T102|relax|39352-0|LNC|Ribs posterior bilateral X-ray|Ribs posterior bilateral X-ray
C0801762|T102|relax|38869-4|LNC|Ribs posterior left X-ray|Ribs posterior left X-ray
C0801762|T102|relax|37964-4|LNC|Ribs posterior right X-ray|Ribs posterior right X-ray
C0801762|T102|relax|26153-7|LNC|Ribs right X-ray|Ribs right X-ray
C0801762|T102|relax|39351-2|LNC|Ribs upper anterior posterior left X-ray|Ribs upper anterior posterior left X-ray
C0801762|T102|relax|39491-6|LNC|Ribs upper anterior posterior right X-ray|Ribs upper anterior posterior right X-ray
C0801762|T102|relax|38867-8|LNC|Ribs upper left X-ray|Ribs upper left X-ray
C0801762|T102|relax|39353-8|LNC|Ribs upper posterior left X-ray|Ribs upper posterior left X-ray
C0801762|T102|relax|39492-4|LNC|Ribs upper posterior right X-ray|Ribs upper posterior right X-ray
C0801762|T102|relax|37961-0|LNC|Ribs upper right X-ray|Ribs upper right X-ray
C0801762|T102|relax|24900-3|LNC|Sacroiliac Joint X-ray|Sacroiliac Joint X-ray
C0801762|T102|relax|36633-6|LNC|Sacroiliac joint bilateral X-ray|Sacroiliac joint bilateral X-ray
C0801762|T102|relax|36634-4|LNC|Sacroiliac joint left X-ray|Sacroiliac joint left X-ray
C0801762|T102|relax|37786-1|LNC|Sacroiliac joint right X-ray|Sacroiliac joint right X-ray
C0801762|T102|relax|30884-1|LNC|Sacrum X-ray|Sacrum X-ray
C0801762|T102|relax|24665-2|LNC|Sacrum Coccyx X-ray|Sacrum Coccyx X-ray
C0801762|T102|relax|39058-3|LNC|Salivary gland X-ray|Salivary gland X-ray
C0801762|T102|relax|24903-7|LNC|Scapula X-ray|Scapula X-ray
C0801762|T102|relax|26154-5|LNC|Scapula bilateral X-ray|Scapula bilateral X-ray
C0801762|T102|relax|26155-2|LNC|Scapula left X-ray|Scapula left X-ray
C0801762|T102|relax|26156-0|LNC|Scapula right X-ray|Scapula right X-ray
C0801762|T102|relax|42159-4|LNC|Sella turcica X-ray|Sella turcica X-ray
C0801762|T102|relax|24909-4|LNC|Shoulder X-ray|Shoulder X-ray
C0801762|T102|relax|26157-8|LNC|Shoulder bilateral X-ray|Shoulder bilateral X-ray
C0801762|T102|relax|26158-6|LNC|Shoulder left X-ray|Shoulder left X-ray
C0801762|T102|relax|26159-4|LNC|Shoulder right X-ray|Shoulder right X-ray
C0801762|T102|relax|42160-2|LNC|Shunt X-ray|Shunt X-ray
C0801762|T102|relax|24911-0|LNC|Shunt Fluoroscopy|Shunt Fluoroscopy
C0801762|T102|relax|24916-9|LNC|Sinuses X-ray|Sinuses X-ray
C0801762|T102|relax|28564-3|LNC|Skull X-ray|Skull X-ray
C0801762|T102|relax|48697-7|LNC|Skull base X-ray|Skull base X-ray
C0801762|T102|relax|37338-1|LNC|Skull Facial bones Mandible X-ray|Skull Facial bones Mandible X-ray
C0801762|T102|relax|24946-6|LNC|Spine Cervical X-ray|Spine Cervical X-ray
C0801762|T102|relax|36640-1|LNC|Spine Cervical Fluoroscopy|Spine Cervical Fluoroscopy
C0801762|T102|relax|43538-8|LNC|Spine Cervical Fluoroscopy video|Spine Cervical Fluoroscopy video
C0801762|T102|relax|37481-9|LNC|Spine Cervical Spine Thoracic X-ray|Spine Cervical Spine Thoracic X-ray
C0801762|T102|relax|38008-9|LNC|Spine Cervical Thoracic Lumbar X-ray|Spine Cervical Thoracic Lumbar X-ray
C0801762|T102|relax|43781-4|LNC|Spine Cervicothoracic Junction X-ray|Spine Cervicothoracic Junction X-ray
C0801762|T102|relax|24972-2|LNC|Spine Lumbar X-ray|Spine Lumbar X-ray
C0801762|T102|relax|43536-2|LNC|Spine Lumbar Fluoroscopy video|Spine Lumbar Fluoroscopy video
C0801762|T102|relax|24975-5|LNC|Spine lumbar Sacroiliac joint bilateral X-ray|Spine lumbar Sacroiliac joint bilateral X-ray
C0801762|T102|relax|37340-7|LNC|Spine Lumbar Sacrum X-ray|Spine Lumbar Sacrum X-ray
C0801762|T102|relax|37341-5|LNC|Spine Lumbar Sacrum Coccyx X-ray|Spine Lumbar Sacrum Coccyx X-ray
C0801762|T102|relax|37342-3|LNC|Spine Lumbar Sacrum Sacroiliac Joint Coccyx X-ray|Spine Lumbar Sacrum Sacroiliac Joint Coccyx X-ray
C0801762|T102|relax|46340-6|LNC|Spine Lumbosacral Junction X-ray|Spine Lumbosacral Junction X-ray
C0801762|T102|relax|24983-9|LNC|Spine Thoracic X-ray|Spine Thoracic X-ray
C0801762|T102|relax|42692-4|LNC|Spine Thoracic Lumbar X-ray|Spine Thoracic Lumbar X-ray
C0801762|T102|relax|37975-0|LNC|Spine Thoracolumbar Junction X-ray|Spine Thoracolumbar Junction X-ray
C0801762|T102|relax|37323-3|LNC|Sternoclavicular joint bilateral X-ray|Sternoclavicular joint bilateral X-ray
C0801762|T102|relax|37324-1|LNC|Sternoclavicular joint left X-ray|Sternoclavicular joint left X-ray
C0801762|T102|relax|37965-1|LNC|Sternoclavicular joint right X-ray|Sternoclavicular joint right X-ray
C0801762|T102|relax|24993-8|LNC|Sternoclavicular Joints X-ray|Sternoclavicular Joints X-ray
C0801762|T102|relax|24994-6|LNC|Sternum X-ray|Sternum X-ray
C0801762|T102|relax|72876-6|LNC|Surgical specimen X-ray|Surgical specimen X-ray
C0801762|T102|relax|25000-1|LNC|Temporomandibular joint X-ray|Temporomandibular joint X-ray
C0801762|T102|relax|37325-8|LNC|Temporomandibular joint bilateral X-ray|Temporomandibular joint bilateral X-ray
C0801762|T102|relax|30889-0|LNC|Temporomandibular joint left X-ray|Temporomandibular joint left X-ray
C0801762|T102|relax|30890-8|LNC|Temporomandibular joint right X-ray|Temporomandibular joint right X-ray
C0801762|T102|relax|25006-8|LNC|Thumb X-ray|Thumb X-ray
C0801762|T102|relax|26160-2|LNC|Thumb bilateral X-ray|Thumb bilateral X-ray
C0801762|T102|relax|26161-0|LNC|Thumb left X-ray|Thumb left X-ray
C0801762|T102|relax|26162-8|LNC|Thumb right X-ray|Thumb right X-ray
C0801762|T102|relax|26163-6|LNC|Tibia bilateral Fibula bilateral X-ray|Tibia bilateral Fibula bilateral X-ray
C0801762|T102|relax|26164-4|LNC|Tibia left Fibula left X-ray|Tibia left Fibula left X-ray
C0801762|T102|relax|26165-1|LNC|Tibia right Fibula right X-ray|Tibia right Fibula right X-ray
C0801762|T102|relax|25011-8|LNC|Tibia Fibula X-ray|Tibia Fibula X-ray
C0801762|T102|relax|37530-3|LNC|Toe fifth left X-ray|Toe fifth left X-ray
C0801762|T102|relax|38151-7|LNC|Toe fifth right X-ray|Toe fifth right X-ray
C0801762|T102|relax|37531-1|LNC|Toe fourth left X-ray|Toe fourth left X-ray
C0801762|T102|relax|38150-9|LNC|Toe fourth right X-ray|Toe fourth right X-ray
C0801762|T102|relax|37534-5|LNC|Toe second left X-ray|Toe second left X-ray
C0801762|T102|relax|38148-3|LNC|Toe second right X-ray|Toe second right X-ray
C0801762|T102|relax|37535-2|LNC|Toe third left X-ray|Toe third left X-ray
C0801762|T102|relax|38149-1|LNC|Toe third right X-ray|Toe third right X-ray
C0801762|T102|relax|25013-4|LNC|Toes X-ray|Toes X-ray
C0801762|T102|relax|26166-9|LNC|Toes bilateral X-ray|Toes bilateral X-ray
C0801762|T102|relax|26167-7|LNC|Toes left X-ray|Toes left X-ray
C0801762|T102|relax|26168-5|LNC|Toes right X-ray|Toes right X-ray
C0801762|T102|relax|48464-2|LNC|Trachea Fluoroscopy|Trachea Fluoroscopy
C0801762|T102|relax|24689-2|LNC|Upper extremity X-ray|Upper extremity X-ray
C0801762|T102|relax|26115-6|LNC|Upper extremity bilateral X-ray|Upper extremity bilateral X-ray
C0801762|T102|relax|26116-4|LNC|Upper extremity left X-ray|Upper extremity left X-ray
C0801762|T102|relax|26117-2|LNC|Upper extremity right X-ray|Upper extremity right X-ray
C0801762|T102|relax|24619-9|LNC|Wrist X-ray|Wrist X-ray
C0801762|T102|relax|26169-3|LNC|Wrist bilateral X-ray|Wrist bilateral X-ray
C0801762|T102|relax|26170-1|LNC|Wrist left X-ray|Wrist left X-ray
C0801762|T102|relax|51392-9|LNC|Wrist left Hand left X-ray|Wrist left Hand left X-ray
C0801762|T102|relax|26171-9|LNC|Wrist right X-ray|Wrist right X-ray
C0801762|T102|relax|51388-7|LNC|Wrist right Hand right X-ray|Wrist right Hand right X-ray
C0801762|T102|relax|43468-8|LNC|Unspecified body region X-ray|Unspecified body region X-ray
C0801762|T102|relax|49512-7|LNC|Unspecified body region Fluoroscopy|Unspecified body region Fluoroscopy
C0801762|T102|relax|25074-6|LNC|Zygomatic arch X-ray|Zygomatic arch X-ray
C0801762|T102|relax|26172-7|LNC|Zygomatic arch bilateral X-ray|Zygomatic arch bilateral X-ray
C0801762|T102|relax|26173-5|LNC|Zygomatic arch left X-ray|Zygomatic arch left X-ray
C0801762|T102|relax|26174-3|LNC|Zygomatic arch right X-ray|Zygomatic arch right X-ray
C0801762|T102|relax|51387-9|LNC|Knee bilateral X-ray (AP view standing)|Knee bilateral X-ray (AP view standing)
C0801762|T102|relax|39370-2|LNC|Ankle right X-ray (view W manual stress)|Ankle right X-ray (view W manual stress)
C0801762|T102|relax|30635-7|LNC|Gastrointestine upper Fluoroscopy AP W contrast PO|Gastrointestine upper Fluoroscopy AP W contrast PO
C0801762|T102|relax|42162-8|LNC|Gastrointestine upper Fluoroscopy AP W water soluble contrast PO|Gastrointestine upper Fluoroscopy AP W water soluble contrast PO
C0801762|T102|relax|39400-7|LNC|Wrist right X-ray carpal tunnel|Wrist right X-ray carpal tunnel
C0801762|T102|relax|69131-1|LNC|Hip X-ray Danelius Miller|Hip X-ray Danelius Miller
C0801762|T102|relax|69140-2|LNC|Hip left X-ray Danelius Miller|Hip left X-ray Danelius Miller
C0801762|T102|relax|39513-7|LNC|Hip right X-ray Danelius Miller|Hip right X-ray Danelius Miller
C0801762|T102|relax|39360-3|LNC|Pelvis X-ray inlet outlet|Pelvis X-ray inlet outlet
C0801762|T102|relax|69059-4|LNC|Hip bilateral X-ray lateral crosstable|Hip bilateral X-ray lateral crosstable
C0801762|T102|relax|69139-4|LNC|Hip left X-ray lateral crosstable|Hip left X-ray lateral crosstable
C0801762|T102|relax|39377-7|LNC|Hip right X-ray lateral crosstable|Hip right X-ray lateral crosstable
C0801762|T102|relax|37583-2|LNC|Pelvis Hip bilateral X-ray lateral frog|Pelvis Hip bilateral X-ray lateral frog
C0801762|T102|relax|39372-8|LNC|Ankle right X-ray Mortise|Ankle right X-ray Mortise
C0801762|T102|relax|39373-6|LNC|Elbow right X-ray oblique|Elbow right X-ray oblique
C0801762|T102|relax|39390-0|LNC|Knee right X-ray oblique|Knee right X-ray oblique
C0801762|T102|relax|39511-1|LNC|Pelvis X-ray oblique|Pelvis X-ray oblique
C0801762|T102|relax|39376-9|LNC|Radius right Ulna right X-ray oblique|Radius right Ulna right X-ray oblique
C0801762|T102|relax|42164-4|LNC|Spine Cervical X-ray oblique|Spine Cervical X-ray oblique
C0801762|T102|relax|42163-6|LNC|Spine Lumbar X-ray oblique|Spine Lumbar X-ray oblique
C0801762|T102|relax|39414-8|LNC|Spine Thoracic X-ray oblique|Spine Thoracic X-ray oblique
C0801762|T102|relax|39398-3|LNC|Tibia right Fibula right X-ray oblique|Tibia right Fibula right X-ray oblique
C0801762|T102|relax|69056-0|LNC|Elbow bilateral X-ray obliques|Elbow bilateral X-ray obliques
C0801762|T102|relax|41811-1|LNC|Ribs bilateral Chest X-ray PA chest|Ribs bilateral Chest X-ray PA chest
C0801762|T102|relax|41832-7|LNC|Ribs left Chest X-ray PA chest|Ribs left Chest X-ray PA chest
C0801762|T102|relax|42010-9|LNC|Ribs right Chest X-ray PA chest|Ribs right Chest X-ray PA chest
C0801762|T102|relax|42165-1|LNC|Ribs Chest X-ray PA chest|Ribs Chest X-ray PA chest
C0801762|T102|relax|46389-3|LNC|Elbow bilateral X-ray radial head capitellar|Elbow bilateral X-ray radial head capitellar
C0801762|T102|relax|39391-8|LNC|Knee right X-ray Sunrise|Knee right X-ray Sunrise
C0801762|T102|relax|39412-2|LNC|Spine Thoracic X-ray Swimmers|Spine Thoracic X-ray Swimmers
C0801762|T102|relax|69148-5|LNC|Knee left X-ray tunnel|Knee left X-ray tunnel
C0801762|T102|relax|39389-2|LNC|Knee right X-ray tunnel|Knee right X-ray tunnel
C0801762|T102|relax|30694-4|LNC|Thyroid Scan uptake single|Thyroid Scan uptake single
C0801762|T102|relax|42271-7|LNC|Thyroid Scan uptake W I-123 IV|Thyroid Scan uptake W I-123 IV
C0801762|T102|relax|60527-9|LNC|Thyroid Scan uptake W I-123 PO|Thyroid Scan uptake W I-123 PO
C0801762|T102|relax|25008-4|LNC|Thyroid Scan uptake W I-131 IV|Thyroid Scan uptake W I-131 IV
C0801762|T102|relax|69236-8|LNC|Thyroid Scan uptake W I-131 PO|Thyroid Scan uptake W I-131 PO
C0801762|T102|relax|43672-5|LNC|Thyroid Scan uptake|Thyroid Scan uptake
C0801762|T102|relax|44147-7|LNC|Thyroid Scan uptake W Tc-99m pertechnetate IV|Thyroid Scan uptake W Tc-99m pertechnetate IV
C0801762|T102|relax|42405-1|LNC|Knee X-ray (AP^standing) (lateral^W hyperextension)|Knee X-ray (AP^standing) (lateral^W hyperextension)
C0801762|T102|relax|42401-0|LNC|Spine Lumbar X-ray (AP W R-bending W L-bending WO bending) Lateral|Spine Lumbar X-ray (AP W R-bending W L-bending WO bending) Lateral
C0801762|T102|relax|42411-9|LNC|Spine Lumbar X-ray (AP^W R-bending W L-bending) (lateral^W flexion W extension)|Spine Lumbar X-ray (AP^W R-bending W L-bending) (lateral^W flexion W extension)
C0801762|T102|relax|39392-6|LNC|Shoulder right X-ray (W internal rotation W external rotation) axillary|Shoulder right X-ray (W internal rotation W external rotation) axillary
C0801762|T102|relax|44199-8|LNC|Facial bones X-ray 1 or 2 views|Facial bones X-ray 1 or 2 views
C0801762|T102|relax|44198-0|LNC|Knee X-ray 1 or 2 views|Knee X-ray 1 or 2 views
C0801762|T102|relax|47373-6|LNC|Knee left X-ray 1 or 2 views|Knee left X-ray 1 or 2 views
C0801762|T102|relax|47375-1|LNC|Knee right X-ray 1 or 2 views|Knee right X-ray 1 or 2 views
C0801762|T102|relax|43521-4|LNC|Mandible X-ray 1 or 2 views|Mandible X-ray 1 or 2 views
C0801762|T102|relax|47983-2|LNC|Mastoid bilateral X-ray 1 or 2 views|Mastoid bilateral X-ray 1 or 2 views
C0801762|T102|relax|48489-9|LNC|Mastoid left X-ray 1 or 2 views|Mastoid left X-ray 1 or 2 views
C0801762|T102|relax|48488-1|LNC|Mastoid right X-ray 1 or 2 views|Mastoid right X-ray 1 or 2 views
C0801762|T102|relax|43522-2|LNC|Pelvis X-ray 1 or 2 views|Pelvis X-ray 1 or 2 views
C0801762|T102|relax|48467-5|LNC|Sacroiliac Joint X-ray 1 or 2 views|Sacroiliac Joint X-ray 1 or 2 views
C0801762|T102|relax|43523-0|LNC|Sinuses X-ray 1 or 2 views|Sinuses X-ray 1 or 2 views
C0801762|T102|relax|44202-0|LNC|Knee X-ray 1 or 2 views portable|Knee X-ray 1 or 2 views portable
C0801762|T102|relax|44201-2|LNC|Pelvis X-ray 1 or 2 views portable|Pelvis X-ray 1 or 2 views portable
C0801762|T102|relax|36641-9|LNC|Abdomen X-ray 2 views|Abdomen X-ray 2 views
C0801762|T102|relax|37064-3|LNC|Acetabulum left X-ray 2 views|Acetabulum left X-ray 2 views
C0801762|T102|relax|37664-0|LNC|Acetabulum right X-ray 2 views|Acetabulum right X-ray 2 views
C0801762|T102|relax|36665-8|LNC|Acromioclavicular joint left X-ray 2 views|Acromioclavicular joint left X-ray 2 views
C0801762|T102|relax|37661-6|LNC|Acromioclavicular joint right X-ray 2 views|Acromioclavicular joint right X-ray 2 views
C0801762|T102|relax|24540-7|LNC|Ankle X-ray 2 views|Ankle X-ray 2 views
C0801762|T102|relax|26385-5|LNC|Ankle bilateral X-ray 2 views|Ankle bilateral X-ray 2 views
C0801762|T102|relax|26386-3|LNC|Ankle left X-ray 2 views|Ankle left X-ray 2 views
C0801762|T102|relax|26387-1|LNC|Ankle right X-ray 2 views|Ankle right X-ray 2 views
C0801762|T102|relax|36642-7|LNC|Breast left Mammogram 2 views|Breast left Mammogram 2 views
C0801762|T102|relax|37768-9|LNC|Breast right Mammogram 2 views|Breast right Mammogram 2 views
C0801762|T102|relax|36661-7|LNC|Calcaneus X-ray 2 views|Calcaneus X-ray 2 views
C0801762|T102|relax|48433-7|LNC|Calcaneus bilateral X-ray 2 views|Calcaneus bilateral X-ray 2 views
C0801762|T102|relax|36662-5|LNC|Calcaneus left X-ray 2 views|Calcaneus left X-ray 2 views
C0801762|T102|relax|37718-4|LNC|Calcaneus right X-ray 2 views|Calcaneus right X-ray 2 views
C0801762|T102|relax|36643-5|LNC|Chest X-ray 2 views|Chest X-ray 2 views
C0801762|T102|relax|36644-3|LNC|Chest Fluoroscopy 2 views|Chest Fluoroscopy 2 views
C0801762|T102|relax|36645-0|LNC|Clavicle X-ray 2 views|Clavicle X-ray 2 views
C0801762|T102|relax|36646-8|LNC|Clavicle left X-ray 2 views|Clavicle left X-ray 2 views
C0801762|T102|relax|37679-8|LNC|Clavicle right X-ray 2 views|Clavicle right X-ray 2 views
C0801762|T102|relax|36647-6|LNC|Coccyx X-ray 2 views|Coccyx X-ray 2 views
C0801762|T102|relax|36648-4|LNC|Elbow X-ray 2 views|Elbow X-ray 2 views
C0801762|T102|relax|36649-2|LNC|Elbow bilateral X-ray 2 views|Elbow bilateral X-ray 2 views
C0801762|T102|relax|36650-0|LNC|Elbow left X-ray 2 views|Elbow left X-ray 2 views
C0801762|T102|relax|37681-4|LNC|Elbow right X-ray 2 views|Elbow right X-ray 2 views
C0801762|T102|relax|36652-6|LNC|Femur X-ray 2 views|Femur X-ray 2 views
C0801762|T102|relax|36653-4|LNC|Femur bilateral X-ray 2 views|Femur bilateral X-ray 2 views
C0801762|T102|relax|36654-2|LNC|Femur left X-ray 2 views|Femur left X-ray 2 views
C0801762|T102|relax|37690-5|LNC|Femur right X-ray 2 views|Femur right X-ray 2 views
C0801762|T102|relax|36655-9|LNC|Finger X-ray 2 views|Finger X-ray 2 views
C0801762|T102|relax|36656-7|LNC|Finger left X-ray 2 views|Finger left X-ray 2 views
C0801762|T102|relax|37694-7|LNC|Finger right X-ray 2 views|Finger right X-ray 2 views
C0801762|T102|relax|30784-3|LNC|Foot X-ray 2 views|Foot X-ray 2 views
C0801762|T102|relax|36657-5|LNC|Foot bilateral X-ray 2 views|Foot bilateral X-ray 2 views
C0801762|T102|relax|38846-2|LNC|Foot left X-ray 2 views|Foot left X-ray 2 views
C0801762|T102|relax|37697-0|LNC|Foot right X-ray 2 views|Foot right X-ray 2 views
C0801762|T102|relax|24721-3|LNC|Hand X-ray 2 views|Hand X-ray 2 views
C0801762|T102|relax|26388-9|LNC|Hand bilateral X-ray 2 views|Hand bilateral X-ray 2 views
C0801762|T102|relax|26389-7|LNC|Hand left X-ray 2 views|Hand left X-ray 2 views
C0801762|T102|relax|26390-5|LNC|Hand right X-ray 2 views|Hand right X-ray 2 views
C0801762|T102|relax|36663-3|LNC|Hip X-ray 2 views|Hip X-ray 2 views
C0801762|T102|relax|69058-6|LNC|Hip bilateral X-ray 2 views|Hip bilateral X-ray 2 views
C0801762|T102|relax|36664-1|LNC|Hip left X-ray 2 views|Hip left X-ray 2 views
C0801762|T102|relax|37721-8|LNC|Hip right X-ray 2 views|Hip right X-ray 2 views
C0801762|T102|relax|24765-0|LNC|Humerus X-ray 2 views|Humerus X-ray 2 views
C0801762|T102|relax|26391-3|LNC|Humerus bilateral X-ray 2 views|Humerus bilateral X-ray 2 views
C0801762|T102|relax|26392-1|LNC|Humerus left X-ray 2 views|Humerus left X-ray 2 views
C0801762|T102|relax|26393-9|LNC|Humerus right X-ray 2 views|Humerus right X-ray 2 views
C0801762|T102|relax|24806-2|LNC|Knee X-ray 2 views|Knee X-ray 2 views
C0801762|T102|relax|26394-7|LNC|Knee bilateral X-ray 2 views|Knee bilateral X-ray 2 views
C0801762|T102|relax|26395-4|LNC|Knee left X-ray 2 views|Knee left X-ray 2 views
C0801762|T102|relax|26396-2|LNC|Knee right X-ray 2 views|Knee right X-ray 2 views
C0801762|T102|relax|36651-8|LNC|Lower extremity X-ray 2 views|Lower extremity X-ray 2 views
C0801762|T102|relax|69257-4|LNC|Lower extremity right X-ray 2 views|Lower extremity right X-ray 2 views
C0801762|T102|relax|24861-7|LNC|Patella X-ray 2 views|Patella X-ray 2 views
C0801762|T102|relax|26397-0|LNC|Patella bilateral X-ray 2 views|Patella bilateral X-ray 2 views
C0801762|T102|relax|26398-8|LNC|Patella left X-ray 2 views|Patella left X-ray 2 views
C0801762|T102|relax|26399-6|LNC|Patella right X-ray 2 views|Patella right X-ray 2 views
C0801762|T102|relax|37617-8|LNC|Pelvis X-ray 2 views|Pelvis X-ray 2 views
C0801762|T102|relax|42685-8|LNC|Pelvis Hip left X-ray 2 views|Pelvis Hip left X-ray 2 views
C0801762|T102|relax|42686-6|LNC|Pelvis Hip right X-ray 2 views|Pelvis Hip right X-ray 2 views
C0801762|T102|relax|36659-1|LNC|Radius bilateral Ulna bilateral X-ray 2 views|Radius bilateral Ulna bilateral X-ray 2 views
C0801762|T102|relax|36660-9|LNC|Radius left Ulna left X-ray 2 views|Radius left Ulna left X-ray 2 views
C0801762|T102|relax|37707-7|LNC|Radius right Ulna right X-ray 2 views|Radius right Ulna right X-ray 2 views
C0801762|T102|relax|36658-3|LNC|Radius Ulna X-ray 2 views|Radius Ulna X-ray 2 views
C0801762|T102|relax|39060-9|LNC|Ribs X-ray 2 views|Ribs X-ray 2 views
C0801762|T102|relax|42687-4|LNC|Ribs bilateral X-ray 2 views|Ribs bilateral X-ray 2 views
C0801762|T102|relax|37066-8|LNC|Ribs left X-ray 2 views|Ribs left X-ray 2 views
C0801762|T102|relax|37780-4|LNC|Ribs right X-ray 2 views|Ribs right X-ray 2 views
C0801762|T102|relax|37651-7|LNC|Sacrum X-ray 2 views|Sacrum X-ray 2 views
C0801762|T102|relax|44179-0|LNC|Sacrum Coccyx X-ray 2 views|Sacrum Coccyx X-ray 2 views
C0801762|T102|relax|37655-8|LNC|Scapula X-ray 2 views|Scapula X-ray 2 views
C0801762|T102|relax|36666-6|LNC|Scapula left X-ray 2 views|Scapula left X-ray 2 views
C0801762|T102|relax|37787-9|LNC|Scapula right X-ray 2 views|Scapula right X-ray 2 views
C0801762|T102|relax|42435-8|LNC|Sella turcica X-ray 2 views|Sella turcica X-ray 2 views
C0801762|T102|relax|37840-6|LNC|Shoulder X-ray 2 views|Shoulder X-ray 2 views
C0801762|T102|relax|36667-4|LNC|Shoulder bilateral X-ray 2 views|Shoulder bilateral X-ray 2 views
C0801762|T102|relax|36668-2|LNC|Shoulder left X-ray 2 views|Shoulder left X-ray 2 views
C0801762|T102|relax|37793-7|LNC|Shoulder right X-ray 2 views|Shoulder right X-ray 2 views
C0801762|T102|relax|37853-9|LNC|Sinuses X-ray 2 views|Sinuses X-ray 2 views
C0801762|T102|relax|37867-9|LNC|Skull X-ray 2 views|Skull X-ray 2 views
C0801762|T102|relax|36669-0|LNC|Spine Cervical X-ray 2 views|Spine Cervical X-ray 2 views
C0801762|T102|relax|43784-8|LNC|Spine Cervical Thoracic Lumbar X-ray 2 views|Spine Cervical Thoracic Lumbar X-ray 2 views
C0801762|T102|relax|36670-8|LNC|Spine Lumbar X-ray 2 views|Spine Lumbar X-ray 2 views
C0801762|T102|relax|37905-7|LNC|Spine Thoracic X-ray 2 views|Spine Thoracic X-ray 2 views
C0801762|T102|relax|24984-7|LNC|Spine Thoracic Lumbar X-ray 2 views|Spine Thoracic Lumbar X-ray 2 views
C0801762|T102|relax|69273-1|LNC|Spine Thoracolumbar Junction X-ray 2 views|Spine Thoracolumbar Junction X-ray 2 views
C0801762|T102|relax|37883-6|LNC|Sternum X-ray 2 views|Sternum X-ray 2 views
C0801762|T102|relax|36671-6|LNC|Tibia bilateral Fibula bilateral X-ray 2 views|Tibia bilateral Fibula bilateral X-ray 2 views
C0801762|T102|relax|36672-4|LNC|Tibia left Fibula left X-ray 2 views|Tibia left Fibula left X-ray 2 views
C0801762|T102|relax|37815-8|LNC|Tibia right Fibula right X-ray 2 views|Tibia right Fibula right X-ray 2 views
C0801762|T102|relax|37895-0|LNC|Tibia Fibula X-ray 2 views|Tibia Fibula X-ray 2 views
C0801762|T102|relax|37902-4|LNC|Toes X-ray 2 views|Toes X-ray 2 views
C0801762|T102|relax|37348-0|LNC|Toes bilateral X-ray 2 views|Toes bilateral X-ray 2 views
C0801762|T102|relax|36673-2|LNC|Toes left X-ray 2 views|Toes left X-ray 2 views
C0801762|T102|relax|37821-6|LNC|Toes right X-ray 2 views|Toes right X-ray 2 views
C0801762|T102|relax|37922-2|LNC|Upper extremity X-ray 2 views|Upper extremity X-ray 2 views
C0801762|T102|relax|37925-5|LNC|Wrist X-ray 2 views|Wrist X-ray 2 views
C0801762|T102|relax|37482-7|LNC|Wrist bilateral X-ray 2 views|Wrist bilateral X-ray 2 views
C0801762|T102|relax|37483-5|LNC|Wrist left X-ray 2 views|Wrist left X-ray 2 views
C0801762|T102|relax|37826-5|LNC|Wrist right X-ray 2 views|Wrist right X-ray 2 views
C0801762|T102|relax|69305-1|LNC|Zygomatic arch X-ray 2 views|Zygomatic arch X-ray 2 views
C0801762|T102|relax|42430-9|LNC|Knee right X-ray 2 views (views standing)|Knee right X-ray 2 views (views standing)
C0801762|T102|relax|42009-1|LNC|Chest X-ray 2 views apical|Chest X-ray 2 views apical
C0801762|T102|relax|39378-5|LNC|Knee right X-ray 2 views oblique|Knee right X-ray 2 views oblique
C0801762|T102|relax|48468-3|LNC|Ribs bilateral Chest X-ray 2 views PA chest|Ribs bilateral Chest X-ray 2 views PA chest
C0801762|T102|relax|43467-0|LNC|Chest X-ray 2 views right oblique left oblique|Chest X-ray 2 views right oblique left oblique
C0801762|T102|relax|69060-2|LNC|Knee bilateral X-ray 2 views Sunrise|Knee bilateral X-ray 2 views Sunrise
C0801762|T102|relax|69142-8|LNC|Knee left X-ray 2 views Sunrise|Knee left X-ray 2 views Sunrise
C0801762|T102|relax|39379-3|LNC|Knee right X-ray 2 views Sunrise|Knee right X-ray 2 views Sunrise
C0801762|T102|relax|39380-1|LNC|Knee right X-ray 2 views Sunrise tunnel|Knee right X-ray 2 views Sunrise tunnel
C0801762|T102|relax|69061-0|LNC|Knee bilateral X-ray 2 views tunnel|Knee bilateral X-ray 2 views tunnel
C0801762|T102|relax|41819-4|LNC|Knee left X-ray 2 views tunnel|Knee left X-ray 2 views tunnel
C0801762|T102|relax|39381-9|LNC|Knee right X-ray 2 views tunnel|Knee right X-ray 2 views tunnel
C0801762|T102|relax|69143-6|LNC|Knee left X-ray 2 views tunnel standing|Knee left X-ray 2 views tunnel standing
C0801762|T102|relax|39382-7|LNC|Knee right X-ray 2 views tunnel standing|Knee right X-ray 2 views tunnel standing
C0801762|T102|relax|38118-6|LNC|Neck X-ray 2 views lateral|Neck X-ray 2 views lateral
C0801762|T102|relax|38844-7|LNC|Elbow left X-ray 2 views Oblique|Elbow left X-ray 2 views Oblique
C0801762|T102|relax|37686-3|LNC|Elbow right X-ray 2 views Oblique|Elbow right X-ray 2 views Oblique
C0801762|T102|relax|38871-0|LNC|Knee left X-ray 2 views Oblique|Knee left X-ray 2 views Oblique
C0801762|T102|relax|38108-7|LNC|Knee right X-ray 2 views Oblique|Knee right X-ray 2 views Oblique
C0801762|T102|relax|38874-4|LNC|Tibia left Fibula left X-ray 2 views Oblique|Tibia left Fibula left X-ray 2 views Oblique
C0801762|T102|relax|38114-5|LNC|Tibia right Fibula right X-ray 2 views Oblique|Tibia right Fibula right X-ray 2 views Oblique
C0801762|T102|relax|44181-6|LNC|Sacroiliac Joint X-ray 2 or 3 views|Sacroiliac Joint X-ray 2 or 3 views
C0801762|T102|relax|43539-6|LNC|Spine Cervical X-ray 2 or 3 views|Spine Cervical X-ray 2 or 3 views
C0801762|T102|relax|48469-1|LNC|Spine Lumbar X-ray 2 or 3 views|Spine Lumbar X-ray 2 or 3 views
C0801762|T102|relax|39880-0|LNC|Bone Scan 2 views phase|Bone Scan 2 views phase
C0801762|T102|relax|44184-0|LNC|Elbow X-ray 2 views portable|Elbow X-ray 2 views portable
C0801762|T102|relax|44182-4|LNC|Hand X-ray 2 views portable|Hand X-ray 2 views portable
C0801762|T102|relax|44183-2|LNC|Radius Ulna X-ray 2 views portable|Radius Ulna X-ray 2 views portable
C0801762|T102|relax|36674-0|LNC|Spine Lumbar X-ray 2 views portable|Spine Lumbar X-ray 2 views portable
C0801762|T102|relax|37658-2|LNC|Spine Thoracic Lumbar X-ray 2 views scoliosis|Spine Thoracic Lumbar X-ray 2 views scoliosis
C0801762|T102|relax|38843-9|LNC|Wrist left X-ray 2 views tunnel carpal|Wrist left X-ray 2 views tunnel carpal
C0801762|T102|relax|37678-0|LNC|Wrist right X-ray 2 views tunnel carpal|Wrist right X-ray 2 views tunnel carpal
C0801762|T102|relax|42166-9|LNC|Heart Scan 2 views at rest W Tl-201 IV|Heart Scan 2 views at rest W Tl-201 IV
C0801762|T102|relax|38841-3|LNC|Ankle left X-ray 2 views standing|Ankle left X-ray 2 views standing
C0801762|T102|relax|37675-6|LNC|Ankle right X-ray 2 views standing|Ankle right X-ray 2 views standing
C0801762|T102|relax|37068-4|LNC|Foot bilateral X-ray 2 views standing|Foot bilateral X-ray 2 views standing
C0801762|T102|relax|37069-2|LNC|Foot left X-ray 2 views standing|Foot left X-ray 2 views standing
C0801762|T102|relax|37698-8|LNC|Foot right X-ray 2 views standing|Foot right X-ray 2 views standing
C0801762|T102|relax|36945-4|LNC|Knee bilateral X-ray 2 views standing|Knee bilateral X-ray 2 views standing
C0801762|T102|relax|38851-2|LNC|Knee left X-ray 2 views standing|Knee left X-ray 2 views standing
C0801762|T102|relax|37762-2|LNC|Knee right X-ray 2 views standing|Knee right X-ray 2 views standing
C0801762|T102|relax|36946-2|LNC|Spine Lumbar X-ray 2 views standing|Spine Lumbar X-ray 2 views standing
C0801762|T102|relax|69274-9|LNC|Spine Thoracic X-ray 2 views standing|Spine Thoracic X-ray 2 views standing
C0801762|T102|relax|38840-5|LNC|Ankle left X-ray 2 views W manual stress|Ankle left X-ray 2 views W manual stress
C0801762|T102|relax|37672-3|LNC|Ankle right X-ray 2 views W manual stress|Ankle right X-ray 2 views W manual stress
C0801762|T102|relax|37067-6|LNC|Chest X-ray 2 views W nipple markers|Chest X-ray 2 views W nipple markers
C0801762|T102|relax|36293-9|LNC|Abdomen X-ray 3 views|Abdomen X-ray 3 views
C0801762|T102|relax|37635-0|LNC|Acetabulum X-ray 3 views|Acetabulum X-ray 3 views
C0801762|T102|relax|36294-7|LNC|Ankle X-ray 3 views|Ankle X-ray 3 views
C0801762|T102|relax|36295-4|LNC|Ankle bilateral X-ray 3 views|Ankle bilateral X-ray 3 views
C0801762|T102|relax|36296-2|LNC|Ankle left X-ray 3 views|Ankle left X-ray 3 views
C0801762|T102|relax|37665-7|LNC|Ankle right X-ray 3 views|Ankle right X-ray 3 views
C0801762|T102|relax|36298-8|LNC|Chest X-ray 3 views|Chest X-ray 3 views
C0801762|T102|relax|36299-6|LNC|Elbow X-ray 3 views|Elbow X-ray 3 views
C0801762|T102|relax|36300-2|LNC|Elbow bilateral X-ray 3 views|Elbow bilateral X-ray 3 views
C0801762|T102|relax|36301-0|LNC|Elbow left X-ray 3 views|Elbow left X-ray 3 views
C0801762|T102|relax|37682-2|LNC|Elbow right X-ray 3 views|Elbow right X-ray 3 views
C0801762|T102|relax|36297-0|LNC|Facial bones X-ray 3 views|Facial bones X-ray 3 views
C0801762|T102|relax|36302-8|LNC|Femur X-ray 3 views|Femur X-ray 3 views
C0801762|T102|relax|36303-6|LNC|Finger X-ray 3 views|Finger X-ray 3 views
C0801762|T102|relax|36304-4|LNC|Finger left X-ray 3 views|Finger left X-ray 3 views
C0801762|T102|relax|37695-4|LNC|Finger right X-ray 3 views|Finger right X-ray 3 views
C0801762|T102|relax|36305-1|LNC|Foot X-ray 3 views|Foot X-ray 3 views
C0801762|T102|relax|36306-9|LNC|Foot bilateral X-ray 3 views|Foot bilateral X-ray 3 views
C0801762|T102|relax|36307-7|LNC|Foot left X-ray 3 views|Foot left X-ray 3 views
C0801762|T102|relax|37699-6|LNC|Foot right X-ray 3 views|Foot right X-ray 3 views
C0801762|T102|relax|24722-1|LNC|Hand X-ray 3 views|Hand X-ray 3 views
C0801762|T102|relax|26379-8|LNC|Hand bilateral X-ray 3 views|Hand bilateral X-ray 3 views
C0801762|T102|relax|26380-6|LNC|Hand left X-ray 3 views|Hand left X-ray 3 views
C0801762|T102|relax|26381-4|LNC|Hand right X-ray 3 views|Hand right X-ray 3 views
C0801762|T102|relax|36308-5|LNC|Hip bilateral X-ray 3 views|Hip bilateral X-ray 3 views
C0801762|T102|relax|36309-3|LNC|Hip left X-ray 3 views|Hip left X-ray 3 views
C0801762|T102|relax|37722-6|LNC|Hip right X-ray 3 views|Hip right X-ray 3 views
C0801762|T102|relax|30788-4|LNC|Knee X-ray 3 views|Knee X-ray 3 views
C0801762|T102|relax|36310-1|LNC|Knee bilateral X-ray 3 views|Knee bilateral X-ray 3 views
C0801762|T102|relax|36311-9|LNC|Knee left X-ray 3 views|Knee left X-ray 3 views
C0801762|T102|relax|37742-4|LNC|Knee right X-ray 3 views|Knee right X-ray 3 views
C0801762|T102|relax|36312-7|LNC|Mandible X-ray 3 views|Mandible X-ray 3 views
C0801762|T102|relax|36838-1|LNC|Mastoid X-ray 3 views|Mastoid X-ray 3 views
C0801762|T102|relax|48470-9|LNC|Mastoid left X-ray 3 views|Mastoid left X-ray 3 views
C0801762|T102|relax|48471-7|LNC|Mastoid right X-ray 3 views|Mastoid right X-ray 3 views
C0801762|T102|relax|37604-6|LNC|Nasal bones X-ray 3 views|Nasal bones X-ray 3 views
C0801762|T102|relax|69261-6|LNC|Patella right X-ray 3 views|Patella right X-ray 3 views
C0801762|T102|relax|30766-0|LNC|Pelvis X-ray 3 views|Pelvis X-ray 3 views
C0801762|T102|relax|37256-5|LNC|Pelvis Spine Lumbar X-ray 3 views|Pelvis Spine Lumbar X-ray 3 views
C0801762|T102|relax|39062-5|LNC|Ribs X-ray 3 views|Ribs X-ray 3 views
C0801762|T102|relax|36313-5|LNC|Ribs bilateral X-ray 3 views|Ribs bilateral X-ray 3 views
C0801762|T102|relax|36314-3|LNC|Ribs left X-ray 3 views|Ribs left X-ray 3 views
C0801762|T102|relax|37781-2|LNC|Ribs right X-ray 3 views|Ribs right X-ray 3 views
C0801762|T102|relax|37648-3|LNC|Sacroiliac Joint X-ray 3 views|Sacroiliac Joint X-ray 3 views
C0801762|T102|relax|39061-7|LNC|Sacrum Coccyx X-ray 3 views|Sacrum Coccyx X-ray 3 views
C0801762|T102|relax|24908-6|LNC|Shoulder X-ray 3 views|Shoulder X-ray 3 views
C0801762|T102|relax|26382-2|LNC|Shoulder bilateral X-ray 3 views|Shoulder bilateral X-ray 3 views
C0801762|T102|relax|26383-0|LNC|Shoulder left X-ray 3 views|Shoulder left X-ray 3 views
C0801762|T102|relax|26384-8|LNC|Shoulder right X-ray 3 views|Shoulder right X-ray 3 views
C0801762|T102|relax|37854-7|LNC|Sinuses X-ray 3 views|Sinuses X-ray 3 views
C0801762|T102|relax|24918-5|LNC|Skull X-ray 3 views|Skull X-ray 3 views
C0801762|T102|relax|24941-7|LNC|Spine Cervical X-ray 3 views|Spine Cervical X-ray 3 views
C0801762|T102|relax|30775-1|LNC|Spine Lumbar X-ray 3 views|Spine Lumbar X-ray 3 views
C0801762|T102|relax|37257-3|LNC|Spine Lumbar Sacroiliac Joint X-ray 3 views|Spine Lumbar Sacroiliac Joint X-ray 3 views
C0801762|T102|relax|37259-9|LNC|Spine Lumbar Sacrum X-ray 3 views|Spine Lumbar Sacrum X-ray 3 views
C0801762|T102|relax|37260-7|LNC|Spine Lumbar Sacrum Coccyx X-ray 3 views|Spine Lumbar Sacrum Coccyx X-ray 3 views
C0801762|T102|relax|37261-5|LNC|Spine Lumbar Sacrum Sacroiliac Joint Coccyx X-ray 3 views|Spine Lumbar Sacrum Sacroiliac Joint Coccyx X-ray 3 views
C0801762|T102|relax|37906-5|LNC|Spine Thoracic X-ray 3 views|Spine Thoracic X-ray 3 views
C0801762|T102|relax|37881-0|LNC|Sternoclavicular Joint X-ray 3 views|Sternoclavicular Joint X-ray 3 views
C0801762|T102|relax|37888-5|LNC|Thumb X-ray 3 views|Thumb X-ray 3 views
C0801762|T102|relax|36315-0|LNC|Thumb left X-ray 3 views|Thumb left X-ray 3 views
C0801762|T102|relax|37812-5|LNC|Thumb right X-ray 3 views|Thumb right X-ray 3 views
C0801762|T102|relax|36316-8|LNC|Toes left X-ray 3 views|Toes left X-ray 3 views
C0801762|T102|relax|37820-8|LNC|Toes right X-ray 3 views|Toes right X-ray 3 views
C0801762|T102|relax|37926-3|LNC|Wrist X-ray 3 views|Wrist X-ray 3 views
C0801762|T102|relax|37454-6|LNC|Wrist bilateral X-ray 3 views|Wrist bilateral X-ray 3 views
C0801762|T102|relax|48738-9|LNC|Wrist bilateral Hand bilateral X-ray 3 views|Wrist bilateral Hand bilateral X-ray 3 views
C0801762|T102|relax|37455-3|LNC|Wrist left X-ray 3 views|Wrist left X-ray 3 views
C0801762|T102|relax|37827-3|LNC|Wrist right X-ray 3 views|Wrist right X-ray 3 views
C0801762|T102|relax|48737-1|LNC|Wrist Hand X-ray 3 views|Wrist Hand X-ray 3 views
C0801762|T102|relax|37933-9|LNC|Zygomatic arch X-ray 3 views|Zygomatic arch X-ray 3 views
C0801762|T102|relax|69154-3|LNC|Shoulder left X-ray 3 views axillary|Shoulder left X-ray 3 views axillary
C0801762|T102|relax|39393-4|LNC|Shoulder right X-ray 3 views axillary|Shoulder right X-ray 3 views axillary
C0801762|T102|relax|39399-1|LNC|Wrist right X-ray 3 views carpal tunnel|Wrist right X-ray 3 views carpal tunnel
C0801762|T102|relax|39364-5|LNC|Wrist right X-ray 3 views radial deviation|Wrist right X-ray 3 views radial deviation
C0801762|T102|relax|39404-9|LNC|Sinuses X-ray 3 views submentovertex|Sinuses X-ray 3 views submentovertex
C0801762|T102|relax|39383-5|LNC|Knee right X-ray 3 views Sunrise|Knee right X-ray 3 views Sunrise
C0801762|T102|relax|48472-5|LNC|Spine Thoracic X-ray 3 views Swimmers|Spine Thoracic X-ray 3 views Swimmers
C0801762|T102|relax|39365-2|LNC|Wrist right X-ray 3 views ulnar deviation|Wrist right X-ray 3 views ulnar deviation
C0801762|T102|relax|69155-0|LNC|Shoulder left X-ray 3 views Y|Shoulder left X-ray 3 views Y
C0801762|T102|relax|39394-2|LNC|Shoulder right X-ray 3 views Y|Shoulder right X-ray 3 views Y
C0801762|T102|relax|43499-3|LNC|Foot left X-ray 3 or 4 views|Foot left X-ray 3 or 4 views
C0801762|T102|relax|43483-7|LNC|Foot right X-ray 3 or 4 views|Foot right X-ray 3 or 4 views
C0801762|T102|relax|39901-4|LNC|Bone Scan 3 views phase multiple areas|Bone Scan 3 views phase multiple areas
C0801762|T102|relax|39902-2|LNC|Bone Scan 3 views phase single area|Bone Scan 3 views phase single area
C0801762|T102|relax|39882-6|LNC|Bone Scan 3 views phase whole body|Bone Scan 3 views phase whole body
C0801762|T102|relax|39883-4|LNC|Bone Scan 3 views phase|Bone Scan 3 views phase
C0801762|T102|relax|30776-9|LNC|Spine Lumbar X-ray 3 views portable|Spine Lumbar X-ray 3 views portable
C0801762|T102|relax|69151-9|LNC|Wrist left X-ray 3 views scaphoid|Wrist left X-ray 3 views scaphoid
C0801762|T102|relax|24778-3|LNC|Kidney bilateral X-ray 3 views serial W WO contrast IV|Kidney bilateral X-ray 3 views serial W WO contrast IV
C0801762|T102|relax|69138-6|LNC|Ankle left X-ray 3 views standing|Ankle left X-ray 3 views standing
C0801762|T102|relax|69254-1|LNC|Ankle right X-ray 3 views standing|Ankle right X-ray 3 views standing
C0801762|T102|relax|36947-0|LNC|Foot bilateral X-ray 3 views standing|Foot bilateral X-ray 3 views standing
C0801762|T102|relax|36948-8|LNC|Foot left X-ray 3 views standing|Foot left X-ray 3 views standing
C0801762|T102|relax|37700-2|LNC|Foot right X-ray 3 views standing|Foot right X-ray 3 views standing
C0801762|T102|relax|36949-6|LNC|Spine Lumbar X-ray 3 views standing|Spine Lumbar X-ray 3 views standing
C0801762|T102|relax|42443-2|LNC|Spine Thoracic X-ray 3 views standing|Spine Thoracic X-ray 3 views standing
C0801762|T102|relax|36317-6|LNC|Ankle X-ray 4 views|Ankle X-ray 4 views
C0801762|T102|relax|36319-2|LNC|Breast Mammogram 4 views|Breast Mammogram 4 views
C0801762|T102|relax|36320-0|LNC|Chest X-ray 4 views|Chest X-ray 4 views
C0801762|T102|relax|36321-8|LNC|Chest Fluoroscopy 4 views|Chest Fluoroscopy 4 views
C0801762|T102|relax|36322-6|LNC|Elbow bilateral X-ray 4 views|Elbow bilateral X-ray 4 views
C0801762|T102|relax|36323-4|LNC|Elbow left X-ray 4 views|Elbow left X-ray 4 views
C0801762|T102|relax|37683-0|LNC|Elbow right X-ray 4 views|Elbow right X-ray 4 views
C0801762|T102|relax|36318-4|LNC|Facial bones X-ray 4 views|Facial bones X-ray 4 views
C0801762|T102|relax|36324-2|LNC|Femur left X-ray 4 views|Femur left X-ray 4 views
C0801762|T102|relax|37691-3|LNC|Femur right X-ray 4 views|Femur right X-ray 4 views
C0801762|T102|relax|30789-2|LNC|Knee X-ray 4 views|Knee X-ray 4 views
C0801762|T102|relax|36325-9|LNC|Knee bilateral X-ray 4 views|Knee bilateral X-ray 4 views
C0801762|T102|relax|36326-7|LNC|Knee left X-ray 4 views|Knee left X-ray 4 views
C0801762|T102|relax|37743-2|LNC|Knee right X-ray 4 views|Knee right X-ray 4 views
C0801762|T102|relax|36327-5|LNC|Mandible X-ray 4 views|Mandible X-ray 4 views
C0801762|T102|relax|43534-7|LNC|Mandible left X-ray 4 views|Mandible left X-ray 4 views
C0801762|T102|relax|43535-4|LNC|Mandible right X-ray 4 views|Mandible right X-ray 4 views
C0801762|T102|relax|36839-9|LNC|Mastoid X-ray 4 views|Mastoid X-ray 4 views
C0801762|T102|relax|37609-5|LNC|Optic foramen X-ray 4 views|Optic foramen X-ray 4 views
C0801762|T102|relax|37612-9|LNC|Orbit bilateral X-ray 4 views|Orbit bilateral X-ray 4 views
C0801762|T102|relax|36328-3|LNC|Ribs bilateral X-ray 4 views|Ribs bilateral X-ray 4 views
C0801762|T102|relax|69265-7|LNC|Shoulder X-ray 4 views|Shoulder X-ray 4 views
C0801762|T102|relax|36329-1|LNC|Shoulder bilateral X-ray 4 views|Shoulder bilateral X-ray 4 views
C0801762|T102|relax|36330-9|LNC|Shoulder left X-ray 4 views|Shoulder left X-ray 4 views
C0801762|T102|relax|37794-5|LNC|Shoulder right X-ray 4 views|Shoulder right X-ray 4 views
C0801762|T102|relax|37855-4|LNC|Sinuses X-ray 4 views|Sinuses X-ray 4 views
C0801762|T102|relax|37868-7|LNC|Skull X-ray 4 views|Skull X-ray 4 views
C0801762|T102|relax|36331-7|LNC|Spine Cervical X-ray 4 views|Spine Cervical X-ray 4 views
C0801762|T102|relax|36332-5|LNC|Spine Lumbar X-ray 4 views|Spine Lumbar X-ray 4 views
C0801762|T102|relax|48473-3|LNC|Spine Lumbar Sacrum X-ray 4 views|Spine Lumbar Sacrum X-ray 4 views
C0801762|T102|relax|37907-3|LNC|Spine Thoracic X-ray 4 views|Spine Thoracic X-ray 4 views
C0801762|T102|relax|37882-8|LNC|Sternoclavicular Joint X-ray 4 views|Sternoclavicular Joint X-ray 4 views
C0801762|T102|relax|38155-8|LNC|Wrist X-ray 4 views|Wrist X-ray 4 views
C0801762|T102|relax|37070-0|LNC|Wrist bilateral X-ray 4 views|Wrist bilateral X-ray 4 views
C0801762|T102|relax|37071-8|LNC|Wrist left X-ray 4 views|Wrist left X-ray 4 views
C0801762|T102|relax|37828-1|LNC|Wrist right X-ray 4 views|Wrist right X-ray 4 views
C0801762|T102|relax|37934-7|LNC|Zygomatic arch X-ray 4 views|Zygomatic arch X-ray 4 views
C0801762|T102|relax|69144-4|LNC|Knee left X-ray 4 views AP standing|Knee left X-ray 4 views AP standing
C0801762|T102|relax|39384-3|LNC|Knee right X-ray 4 views AP standing|Knee right X-ray 4 views AP standing
C0801762|T102|relax|39385-0|LNC|Knee right X-ray 4 views oblique|Knee right X-ray 4 views oblique
C0801762|T102|relax|39413-0|LNC|Spine Thoracic X-ray 4 views oblique|Spine Thoracic X-ray 4 views oblique
C0801762|T102|relax|39099-7|LNC|Ribs bilateral Chest X-ray 4 views PA chest|Ribs bilateral Chest X-ray 4 views PA chest
C0801762|T102|relax|69063-6|LNC|Knee bilateral X-ray 4 views Sunrise tunnel|Knee bilateral X-ray 4 views Sunrise tunnel
C0801762|T102|relax|39387-6|LNC|Knee right X-ray 4 views Sunrise tunnel|Knee right X-ray 4 views Sunrise tunnel
C0801762|T102|relax|69145-1|LNC|Knee left X-ray 4 views tunnel|Knee left X-ray 4 views tunnel
C0801762|T102|relax|39386-8|LNC|Knee right X-ray 4 views tunnel|Knee right X-ray 4 views tunnel
C0801762|T102|relax|69062-8|LNC|Knee bilateral X-ray 4 views standing|Knee bilateral X-ray 4 views standing
C0801762|T102|relax|38852-0|LNC|Knee left X-ray 4 views standing|Knee left X-ray 4 views standing
C0801762|T102|relax|37763-0|LNC|Knee right X-ray 4 views standing|Knee right X-ray 4 views standing
C0801762|T102|relax|36675-7|LNC|Facial bones X-ray 5 views|Facial bones X-ray 5 views
C0801762|T102|relax|36676-5|LNC|Knee left X-ray 5 views|Knee left X-ray 5 views
C0801762|T102|relax|37744-0|LNC|Knee right X-ray 5 views|Knee right X-ray 5 views
C0801762|T102|relax|36890-2|LNC|Mastoid X-ray 5 views|Mastoid X-ray 5 views
C0801762|T102|relax|37351-4|LNC|Pelvis Spine Lumbar X-ray 5 views|Pelvis Spine Lumbar X-ray 5 views
C0801762|T102|relax|30750-4|LNC|Shoulder X-ray 5 views|Shoulder X-ray 5 views
C0801762|T102|relax|36677-3|LNC|Shoulder left X-ray 5 views|Shoulder left X-ray 5 views
C0801762|T102|relax|37795-2|LNC|Shoulder right X-ray 5 views|Shoulder right X-ray 5 views
C0801762|T102|relax|37856-2|LNC|Sinuses X-ray 5 views|Sinuses X-ray 5 views
C0801762|T102|relax|24922-7|LNC|Skull X-ray 5 views|Skull X-ray 5 views
C0801762|T102|relax|24939-1|LNC|Spine Cervical X-ray 5 views|Spine Cervical X-ray 5 views
C0801762|T102|relax|30797-5|LNC|Spine Lumbar X-ray 5 views|Spine Lumbar X-ray 5 views
C0801762|T102|relax|37353-0|LNC|Spine Lumbar Sacroiliac Joint X-ray 5 views|Spine Lumbar Sacroiliac Joint X-ray 5 views
C0801762|T102|relax|37355-5|LNC|Spine Lumbar Sacrum X-ray 5 views|Spine Lumbar Sacrum X-ray 5 views
C0801762|T102|relax|37356-3|LNC|Spine Lumbar Sacrum Coccyx X-ray 5 views|Spine Lumbar Sacrum Coccyx X-ray 5 views
C0801762|T102|relax|37357-1|LNC|Spine Lumbar Sacrum Sacroiliac Joint Coccyx X-ray 5 views|Spine Lumbar Sacrum Sacroiliac Joint Coccyx X-ray 5 views
C0801762|T102|relax|37350-6|LNC|Temporomandibular joint bilateral X-ray 5 views|Temporomandibular joint bilateral X-ray 5 views
C0801762|T102|relax|37072-6|LNC|Wrist left X-ray 5 views|Wrist left X-ray 5 views
C0801762|T102|relax|37829-9|LNC|Wrist right X-ray 5 views|Wrist right X-ray 5 views
C0801762|T102|relax|39407-2|LNC|Spine Thoracic X-ray 5 views oblique|Spine Thoracic X-ray 5 views oblique
C0801762|T102|relax|69081-8|LNC|Spine Cervical X-ray 5 views Swimmers|Spine Cervical X-ray 5 views Swimmers
C0801762|T102|relax|37073-4|LNC|Spine Lumbar X-ray 5 views standing|Spine Lumbar X-ray 5 views standing
C0801762|T102|relax|69080-0|LNC|Spine Cervical X-ray 5 views W flexion W extension|Spine Cervical X-ray 5 views W flexion W extension
C0801762|T102|relax|39063-3|LNC|Spine Lumbar X-ray 5 views W flexion W extension|Spine Lumbar X-ray 5 views W flexion W extension
C0801762|T102|relax|42273-3|LNC|Ankle bilateral X-ray 6 views|Ankle bilateral X-ray 6 views
C0801762|T102|relax|36678-1|LNC|Knee bilateral X-ray 6 views|Knee bilateral X-ray 6 views
C0801762|T102|relax|36679-9|LNC|Shoulder left X-ray 6 views|Shoulder left X-ray 6 views
C0801762|T102|relax|37796-0|LNC|Shoulder right X-ray 6 views|Shoulder right X-ray 6 views
C0801762|T102|relax|42691-6|LNC|Spine Cervical X-ray 6 views|Spine Cervical X-ray 6 views
C0801762|T102|relax|38156-6|LNC|Wrist X-ray 6 views|Wrist X-ray 6 views
C0801762|T102|relax|37074-2|LNC|Wrist left X-ray 6 views|Wrist left X-ray 6 views
C0801762|T102|relax|37830-7|LNC|Wrist right X-ray 6 views|Wrist right X-ray 6 views
C0801762|T102|relax|36680-7|LNC|Spine Cervical X-ray 7 views|Spine Cervical X-ray 7 views
C0801762|T102|relax|36681-5|LNC|Spine Lumbar X-ray 7 views|Spine Lumbar X-ray 7 views
C0801762|T102|relax|36682-3|LNC|Knee bilateral X-ray 8 views|Knee bilateral X-ray 8 views
C0801762|T102|relax|36683-1|LNC|Wrist left X-ray 8 views|Wrist left X-ray 8 views
C0801762|T102|relax|37831-5|LNC|Wrist right X-ray 8 views|Wrist right X-ray 8 views
C0801762|T102|relax|42412-7|LNC|Shoulder left X-ray 90 degree abduction|Shoulder left X-ray 90 degree abduction
C0801762|T102|relax|39064-1|LNC|Ribs X-ray anterior lateral|Ribs X-ray anterior lateral
C0801762|T102|relax|69070-1|LNC|Ribs bilateral X-ray anterior lateral|Ribs bilateral X-ray anterior lateral
C0801762|T102|relax|38856-1|LNC|Ribs left X-ray anterior lateral|Ribs left X-ray anterior lateral
C0801762|T102|relax|37782-0|LNC|Ribs right X-ray anterior lateral|Ribs right X-ray anterior lateral
C0801762|T102|relax|24796-5|LNC|Abdomen X-ray AP AP left lateral-decubitus|Abdomen X-ray AP AP left lateral-decubitus
C0801762|T102|relax|24792-4|LNC|Abdomen X-ray AP AP left lateral-decubitus portable|Abdomen X-ray AP AP left lateral-decubitus portable
C0801762|T102|relax|24653-8|LNC|Chest X-ray AP AP right lateral-decubitus|Chest X-ray AP AP right lateral-decubitus
C0801762|T102|relax|24654-6|LNC|Chest X-ray AP AP right lateral-decubitus portable|Chest X-ray AP AP right lateral-decubitus portable
C0801762|T102|relax|37080-9|LNC|Shoulder bilateral X-ray AP axillary|Shoulder bilateral X-ray AP axillary
C0801762|T102|relax|37081-7|LNC|Shoulder bilateral X-ray AP axillary outlet|Shoulder bilateral X-ray AP axillary outlet
C0801762|T102|relax|37082-5|LNC|Shoulder left X-ray AP axillary outlet|Shoulder left X-ray AP axillary outlet
C0801762|T102|relax|38781-1|LNC|Shoulder right X-ray AP axillary outlet|Shoulder right X-ray AP axillary outlet
C0801762|T102|relax|39339-7|LNC|Shoulder bilateral X-ray AP axillary outlet 30 degree caudal angle|Shoulder bilateral X-ray AP axillary outlet 30 degree caudal angle
C0801762|T102|relax|37083-3|LNC|Shoulder left X-ray AP axillary outlet Zanca|Shoulder left X-ray AP axillary outlet Zanca
C0801762|T102|relax|38782-9|LNC|Shoulder right X-ray AP axillary outlet Zanca|Shoulder right X-ray AP axillary outlet Zanca
C0801762|T102|relax|37126-0|LNC|Shoulder bilateral X-ray AP axillary Y|Shoulder bilateral X-ray AP axillary Y
C0801762|T102|relax|37084-1|LNC|Shoulder left X-ray AP axillary Y|Shoulder left X-ray AP axillary Y
C0801762|T102|relax|38783-7|LNC|Shoulder right X-ray AP axillary Y|Shoulder right X-ray AP axillary Y
C0801762|T102|relax|39512-9|LNC|Hip right X-ray AP Danelius Miller|Hip right X-ray AP Danelius Miller
C0801762|T102|relax|39401-5|LNC|Shoulder X-ray AP Grashey axillary|Shoulder X-ray AP Grashey axillary
C0801762|T102|relax|69153-5|LNC|Shoulder left X-ray AP Grashey axillary|Shoulder left X-ray AP Grashey axillary
C0801762|T102|relax|69262-4|LNC|Shoulder right X-ray AP Grashey axillary|Shoulder right X-ray AP Grashey axillary
C0801762|T102|relax|37618-6|LNC|Pelvis X-ray AP inlet|Pelvis X-ray AP inlet
C0801762|T102|relax|37623-6|LNC|Pelvis X-ray AP inlet outlet|Pelvis X-ray AP inlet outlet
C0801762|T102|relax|39065-8|LNC|Pelvis X-ray AP inlet outlet oblique|Pelvis X-ray AP inlet outlet oblique
C0801762|T102|relax|37619-4|LNC|Pelvis X-ray AP Judet|Pelvis X-ray AP Judet
C0801762|T102|relax|24794-0|LNC|Abdomen X-ray AP lateral|Abdomen X-ray AP lateral
C0801762|T102|relax|30779-3|LNC|Ankle X-ray AP lateral|Ankle X-ray AP lateral
C0801762|T102|relax|36684-9|LNC|Ankle bilateral X-ray AP lateral|Ankle bilateral X-ray AP lateral
C0801762|T102|relax|36685-6|LNC|Ankle left X-ray AP lateral|Ankle left X-ray AP lateral
C0801762|T102|relax|37667-3|LNC|Ankle right X-ray AP lateral|Ankle right X-ray AP lateral
C0801762|T102|relax|36686-4|LNC|Calcaneus bilateral X-ray AP lateral|Calcaneus bilateral X-ray AP lateral
C0801762|T102|relax|36701-1|LNC|Calcaneus left X-ray AP lateral|Calcaneus left X-ray AP lateral
C0801762|T102|relax|37719-2|LNC|Calcaneus right X-ray AP lateral|Calcaneus right X-ray AP lateral
C0801762|T102|relax|36687-2|LNC|Chest X-ray AP lateral|Chest X-ray AP lateral
C0801762|T102|relax|39066-6|LNC|Chest Fluoroscopy AP lateral|Chest Fluoroscopy AP lateral
C0801762|T102|relax|36688-0|LNC|Coccyx X-ray AP lateral|Coccyx X-ray AP lateral
C0801762|T102|relax|36689-8|LNC|Elbow X-ray AP lateral|Elbow X-ray AP lateral
C0801762|T102|relax|36690-6|LNC|Elbow bilateral X-ray AP lateral|Elbow bilateral X-ray AP lateral
C0801762|T102|relax|36691-4|LNC|Elbow left X-ray AP lateral|Elbow left X-ray AP lateral
C0801762|T102|relax|37684-8|LNC|Elbow right X-ray AP lateral|Elbow right X-ray AP lateral
C0801762|T102|relax|36693-0|LNC|Femur X-ray AP lateral|Femur X-ray AP lateral
C0801762|T102|relax|36694-8|LNC|Femur bilateral X-ray AP lateral|Femur bilateral X-ray AP lateral
C0801762|T102|relax|36695-5|LNC|Femur left X-ray AP lateral|Femur left X-ray AP lateral
C0801762|T102|relax|37692-1|LNC|Femur right X-ray AP lateral|Femur right X-ray AP lateral
C0801762|T102|relax|39069-0|LNC|Foot X-ray AP lateral|Foot X-ray AP lateral
C0801762|T102|relax|36696-3|LNC|Foot bilateral X-ray AP lateral|Foot bilateral X-ray AP lateral
C0801762|T102|relax|36697-1|LNC|Foot left X-ray AP lateral|Foot left X-ray AP lateral
C0801762|T102|relax|37701-0|LNC|Foot right X-ray AP lateral|Foot right X-ray AP lateral
C0801762|T102|relax|42409-3|LNC|Foot sesamoid bones X-ray AP lateral|Foot sesamoid bones X-ray AP lateral
C0801762|T102|relax|69130-3|LNC|Hand X-ray AP lateral|Hand X-ray AP lateral
C0801762|T102|relax|48474-1|LNC|Hand bilateral X-ray AP lateral|Hand bilateral X-ray AP lateral
C0801762|T102|relax|38847-0|LNC|Hand left X-ray AP lateral|Hand left X-ray AP lateral
C0801762|T102|relax|37710-1|LNC|Hand right X-ray AP lateral|Hand right X-ray AP lateral
C0801762|T102|relax|36702-9|LNC|Hip X-ray AP lateral|Hip X-ray AP lateral
C0801762|T102|relax|36703-7|LNC|Hip bilateral X-ray AP lateral|Hip bilateral X-ray AP lateral
C0801762|T102|relax|36704-5|LNC|Hip left X-ray AP lateral|Hip left X-ray AP lateral
C0801762|T102|relax|37725-9|LNC|Hip right X-ray AP lateral|Hip right X-ray AP lateral
C0801762|T102|relax|36706-0|LNC|Humerus X-ray AP lateral|Humerus X-ray AP lateral
C0801762|T102|relax|36707-8|LNC|Humerus bilateral X-ray AP lateral|Humerus bilateral X-ray AP lateral
C0801762|T102|relax|36708-6|LNC|Humerus left X-ray AP lateral|Humerus left X-ray AP lateral
C0801762|T102|relax|37736-6|LNC|Humerus right X-ray AP lateral|Humerus right X-ray AP lateral
C0801762|T102|relax|36709-4|LNC|Knee X-ray AP lateral|Knee X-ray AP lateral
C0801762|T102|relax|36590-8|LNC|Knee bilateral X-ray AP lateral|Knee bilateral X-ray AP lateral
C0801762|T102|relax|36710-2|LNC|Knee left X-ray AP lateral|Knee left X-ray AP lateral
C0801762|T102|relax|37745-7|LNC|Knee right X-ray AP lateral|Knee right X-ray AP lateral
C0801762|T102|relax|36692-2|LNC|Lower extremity X-ray AP lateral|Lower extremity X-ray AP lateral
C0801762|T102|relax|69258-2|LNC|Lower extremity right X-ray AP lateral|Lower extremity right X-ray AP lateral
C0801762|T102|relax|36711-0|LNC|Mandible X-ray AP lateral|Mandible X-ray AP lateral
C0801762|T102|relax|42438-2|LNC|Neck X-ray AP lateral|Neck X-ray AP lateral
C0801762|T102|relax|36712-8|LNC|Patella bilateral X-ray AP lateral|Patella bilateral X-ray AP lateral
C0801762|T102|relax|36713-6|LNC|Patella left X-ray AP lateral|Patella left X-ray AP lateral
C0801762|T102|relax|37776-2|LNC|Patella right X-ray AP lateral|Patella right X-ray AP lateral
C0801762|T102|relax|37620-2|LNC|Pelvis X-ray AP lateral|Pelvis X-ray AP lateral
C0801762|T102|relax|36705-2|LNC|Pelvis Hip X-ray AP lateral|Pelvis Hip X-ray AP lateral
C0801762|T102|relax|36699-7|LNC|Radius bilateral Ulna bilateral X-ray AP lateral|Radius bilateral Ulna bilateral X-ray AP lateral
C0801762|T102|relax|36700-3|LNC|Radius left Ulna left X-ray AP lateral|Radius left Ulna left X-ray AP lateral
C0801762|T102|relax|37708-5|LNC|Radius right Ulna right X-ray AP lateral|Radius right Ulna right X-ray AP lateral
C0801762|T102|relax|36698-9|LNC|Radius Ulna X-ray AP lateral|Radius Ulna X-ray AP lateral
C0801762|T102|relax|37652-5|LNC|Sacrum X-ray AP lateral|Sacrum X-ray AP lateral
C0801762|T102|relax|36714-4|LNC|Scapula bilateral X-ray AP lateral|Scapula bilateral X-ray AP lateral
C0801762|T102|relax|36715-1|LNC|Scapula left X-ray AP lateral|Scapula left X-ray AP lateral
C0801762|T102|relax|37788-7|LNC|Scapula right X-ray AP lateral|Scapula right X-ray AP lateral
C0801762|T102|relax|37841-4|LNC|Shoulder X-ray AP lateral|Shoulder X-ray AP lateral
C0801762|T102|relax|36716-9|LNC|Shoulder bilateral X-ray AP lateral|Shoulder bilateral X-ray AP lateral
C0801762|T102|relax|24919-3|LNC|Skull X-ray AP lateral|Skull X-ray AP lateral
C0801762|T102|relax|24942-5|LNC|Spine Cervical X-ray AP lateral|Spine Cervical X-ray AP lateral
C0801762|T102|relax|37361-3|LNC|Spine Cervical Spine Thoracic X-ray AP lateral|Spine Cervical Spine Thoracic X-ray AP lateral
C0801762|T102|relax|39067-4|LNC|Spine Cervical Thoracic Lumbar X-ray AP lateral|Spine Cervical Thoracic Lumbar X-ray AP lateral
C0801762|T102|relax|43785-5|LNC|Spine Cervicothoracic Junction X-ray AP lateral|Spine Cervicothoracic Junction X-ray AP lateral
C0801762|T102|relax|24970-6|LNC|Spine Lumbar X-ray AP lateral|Spine Lumbar X-ray AP lateral
C0801762|T102|relax|30753-8|LNC|Spine Thoracic X-ray AP lateral|Spine Thoracic X-ray AP lateral
C0801762|T102|relax|38123-6|LNC|Spine Thoracic Lumbar X-ray AP lateral|Spine Thoracic Lumbar X-ray AP lateral
C0801762|T102|relax|37974-3|LNC|Spine Thoracolumbar Junction X-ray AP lateral|Spine Thoracolumbar Junction X-ray AP lateral
C0801762|T102|relax|37889-3|LNC|Thumb X-ray AP lateral|Thumb X-ray AP lateral
C0801762|T102|relax|36717-7|LNC|Tibia bilateral Fibula bilateral X-ray AP lateral|Tibia bilateral Fibula bilateral X-ray AP lateral
C0801762|T102|relax|36718-5|LNC|Tibia left Fibula left X-ray AP lateral|Tibia left Fibula left X-ray AP lateral
C0801762|T102|relax|37816-6|LNC|Tibia right Fibula right X-ray AP lateral|Tibia right Fibula right X-ray AP lateral
C0801762|T102|relax|37896-8|LNC|Tibia Fibula X-ray AP lateral|Tibia Fibula X-ray AP lateral
C0801762|T102|relax|36719-3|LNC|Toes left X-ray AP lateral|Toes left X-ray AP lateral
C0801762|T102|relax|37822-4|LNC|Toes right X-ray AP lateral|Toes right X-ray AP lateral
C0801762|T102|relax|30793-4|LNC|Wrist X-ray AP lateral|Wrist X-ray AP lateral
C0801762|T102|relax|38860-3|LNC|Wrist left X-ray AP lateral|Wrist left X-ray AP lateral
C0801762|T102|relax|37832-3|LNC|Wrist right X-ray AP lateral|Wrist right X-ray AP lateral
C0801762|T102|relax|37839-8|LNC|Shoulder X-ray AP lateral axillary|Shoulder X-ray AP lateral axillary
C0801762|T102|relax|39070-8|LNC|Chest X-ray AP lateral lordotic|Chest X-ray AP lateral lordotic
C0801762|T102|relax|42404-4|LNC|Hip left X-ray AP lateral measurement|Hip left X-ray AP lateral measurement
C0801762|T102|relax|39071-6|LNC|Knee X-ray AP lateral Merchants|Knee X-ray AP lateral Merchants
C0801762|T102|relax|37095-7|LNC|Ankle X-ray AP lateral Mortise|Ankle X-ray AP lateral Mortise
C0801762|T102|relax|37096-5|LNC|Ankle bilateral X-ray AP lateral Mortise|Ankle bilateral X-ray AP lateral Mortise
C0801762|T102|relax|37097-3|LNC|Ankle left X-ray AP lateral Mortise|Ankle left X-ray AP lateral Mortise
C0801762|T102|relax|37666-5|LNC|Ankle right X-ray AP lateral Mortise|Ankle right X-ray AP lateral Mortise
C0801762|T102|relax|39072-4|LNC|Ankle X-ray AP lateral oblique|Ankle X-ray AP lateral oblique
C0801762|T102|relax|36720-1|LNC|Ankle bilateral X-ray AP lateral oblique|Ankle bilateral X-ray AP lateral oblique
C0801762|T102|relax|36721-9|LNC|Ankle left X-ray AP lateral oblique|Ankle left X-ray AP lateral oblique
C0801762|T102|relax|37668-1|LNC|Ankle right X-ray AP lateral oblique|Ankle right X-ray AP lateral oblique
C0801762|T102|relax|36731-8|LNC|Calcaneus X-ray AP lateral oblique|Calcaneus X-ray AP lateral oblique
C0801762|T102|relax|36722-7|LNC|Elbow X-ray AP lateral oblique|Elbow X-ray AP lateral oblique
C0801762|T102|relax|36723-5|LNC|Elbow bilateral X-ray AP lateral oblique|Elbow bilateral X-ray AP lateral oblique
C0801762|T102|relax|36724-3|LNC|Elbow left X-ray AP lateral oblique|Elbow left X-ray AP lateral oblique
C0801762|T102|relax|37685-5|LNC|Elbow right X-ray AP lateral oblique|Elbow right X-ray AP lateral oblique
C0801762|T102|relax|36725-0|LNC|Finger X-ray AP lateral oblique|Finger X-ray AP lateral oblique
C0801762|T102|relax|36726-8|LNC|Finger bilateral X-ray AP lateral oblique|Finger bilateral X-ray AP lateral oblique
C0801762|T102|relax|36727-6|LNC|Finger left X-ray AP lateral oblique|Finger left X-ray AP lateral oblique
C0801762|T102|relax|37696-2|LNC|Finger right X-ray AP lateral oblique|Finger right X-ray AP lateral oblique
C0801762|T102|relax|36728-4|LNC|Foot X-ray AP lateral oblique|Foot X-ray AP lateral oblique
C0801762|T102|relax|36729-2|LNC|Foot bilateral X-ray AP lateral oblique|Foot bilateral X-ray AP lateral oblique
C0801762|T102|relax|36730-0|LNC|Foot left X-ray AP lateral oblique|Foot left X-ray AP lateral oblique
C0801762|T102|relax|37702-8|LNC|Foot right X-ray AP lateral oblique|Foot right X-ray AP lateral oblique
C0801762|T102|relax|69057-8|LNC|Hand bilateral X-ray AP lateral oblique|Hand bilateral X-ray AP lateral oblique
C0801762|T102|relax|38848-8|LNC|Hand left X-ray AP lateral oblique|Hand left X-ray AP lateral oblique
C0801762|T102|relax|37711-9|LNC|Hand right X-ray AP lateral oblique|Hand right X-ray AP lateral oblique
C0801762|T102|relax|36732-6|LNC|Knee bilateral X-ray AP lateral oblique|Knee bilateral X-ray AP lateral oblique
C0801762|T102|relax|36733-4|LNC|Knee left X-ray AP lateral oblique|Knee left X-ray AP lateral oblique
C0801762|T102|relax|37748-1|LNC|Knee right X-ray AP lateral oblique|Knee right X-ray AP lateral oblique
C0801762|T102|relax|37624-4|LNC|Pelvis X-ray AP lateral oblique|Pelvis X-ray AP lateral oblique
C0801762|T102|relax|36734-2|LNC|Spine Cervical X-ray AP lateral oblique|Spine Cervical X-ray AP lateral oblique
C0801762|T102|relax|36735-9|LNC|Spine Lumbar X-ray AP lateral oblique|Spine Lumbar X-ray AP lateral oblique
C0801762|T102|relax|37908-1|LNC|Spine Thoracic X-ray AP lateral oblique|Spine Thoracic X-ray AP lateral oblique
C0801762|T102|relax|36736-7|LNC|Thumb left X-ray AP lateral oblique|Thumb left X-ray AP lateral oblique
C0801762|T102|relax|37813-3|LNC|Thumb right X-ray AP lateral oblique|Thumb right X-ray AP lateral oblique
C0801762|T102|relax|37927-1|LNC|Wrist X-ray AP lateral oblique|Wrist X-ray AP lateral oblique
C0801762|T102|relax|37099-9|LNC|Spine Cervical X-ray AP lateral oblique odontoid|Spine Cervical X-ray AP lateral oblique odontoid
C0801762|T102|relax|38083-2|LNC|Spine Cervical X-ray AP lateral oblique odontoid swimmer|Spine Cervical X-ray AP lateral oblique odontoid swimmer
C0801762|T102|relax|37101-3|LNC|Spine Lumbar X-ray AP lateral oblique spot|Spine Lumbar X-ray AP lateral oblique spot
C0801762|T102|relax|42410-1|LNC|Spine Lumbar X-ray AP lateral oblique spot standing|Spine Lumbar X-ray AP lateral oblique spot standing
C0801762|T102|relax|37102-1|LNC|Knee bilateral X-ray AP lateral oblique Sunrise|Knee bilateral X-ray AP lateral oblique Sunrise
C0801762|T102|relax|37118-7|LNC|Knee bilateral X-ray AP lateral oblique Sunrise tunnel|Knee bilateral X-ray AP lateral oblique Sunrise tunnel
C0801762|T102|relax|37115-3|LNC|Knee X-ray AP lateral oblique tunnel|Knee X-ray AP lateral oblique tunnel
C0801762|T102|relax|69137-8|LNC|Ankle left X-ray AP lateral oblique standing|Ankle left X-ray AP lateral oblique standing
C0801762|T102|relax|39371-0|LNC|Ankle right X-ray AP lateral oblique standing|Ankle right X-ray AP lateral oblique standing
C0801762|T102|relax|39334-8|LNC|Foot left X-ray AP lateral oblique standing|Foot left X-ray AP lateral oblique standing
C0801762|T102|relax|39375-1|LNC|Foot right X-ray AP lateral oblique standing|Foot right X-ray AP lateral oblique standing
C0801762|T102|relax|42417-6|LNC|Ankle bilateral X-ray AP lateral oblique W manual stress|Ankle bilateral X-ray AP lateral oblique W manual stress
C0801762|T102|relax|42418-4|LNC|Ankle left X-ray AP lateral oblique W manual stress|Ankle left X-ray AP lateral oblique W manual stress
C0801762|T102|relax|39369-4|LNC|Ankle right X-ray AP lateral oblique W manual stress|Ankle right X-ray AP lateral oblique W manual stress
C0801762|T102|relax|37103-9|LNC|Spine Cervical X-ray AP lateral odontoid|Spine Cervical X-ray AP lateral odontoid
C0801762|T102|relax|37079-1|LNC|Spine Cervical X-ray AP lateral odontoid portable|Spine Cervical X-ray AP lateral odontoid portable
C0801762|T102|relax|39074-0|LNC|Chest X-ray AP lateral right oblique left oblique|Chest X-ray AP lateral right oblique left oblique
C0801762|T102|relax|39073-2|LNC|Knee X-ray AP lateral right oblique left oblique|Knee X-ray AP lateral right oblique left oblique
C0801762|T102|relax|69147-7|LNC|Knee left X-ray AP lateral right oblique left oblique|Knee left X-ray AP lateral right oblique left oblique
C0801762|T102|relax|39388-4|LNC|Knee right X-ray AP lateral right oblique left oblique|Knee right X-ray AP lateral right oblique left oblique
C0801762|T102|relax|37105-4|LNC|Spine Lumbar X-ray AP lateral spot|Spine Lumbar X-ray AP lateral spot
C0801762|T102|relax|37106-2|LNC|Knee X-ray AP lateral Sunrise|Knee X-ray AP lateral Sunrise
C0801762|T102|relax|37107-0|LNC|Knee bilateral X-ray AP lateral Sunrise|Knee bilateral X-ray AP lateral Sunrise
C0801762|T102|relax|37108-8|LNC|Knee left X-ray AP lateral Sunrise|Knee left X-ray AP lateral Sunrise
C0801762|T102|relax|37749-9|LNC|Knee right X-ray AP lateral Sunrise|Knee right X-ray AP lateral Sunrise
C0801762|T102|relax|37109-6|LNC|Patella bilateral X-ray AP lateral Sunrise|Patella bilateral X-ray AP lateral Sunrise
C0801762|T102|relax|37110-4|LNC|Patella left X-ray AP lateral Sunrise|Patella left X-ray AP lateral Sunrise
C0801762|T102|relax|38786-0|LNC|Patella right X-ray AP lateral Sunrise|Patella right X-ray AP lateral Sunrise
C0801762|T102|relax|37111-2|LNC|Knee X-ray AP lateral Sunrise tunnel|Knee X-ray AP lateral Sunrise tunnel
C0801762|T102|relax|37116-1|LNC|Knee bilateral X-ray AP lateral Sunrise tunnel|Knee bilateral X-ray AP lateral Sunrise tunnel
C0801762|T102|relax|37117-9|LNC|Knee left X-ray AP lateral Sunrise tunnel|Knee left X-ray AP lateral Sunrise tunnel
C0801762|T102|relax|37740-8|LNC|Knee right X-ray AP lateral Sunrise tunnel|Knee right X-ray AP lateral Sunrise tunnel
C0801762|T102|relax|38009-7|LNC|Spine Thoracic X-ray AP lateral Swimmers|Spine Thoracic X-ray AP lateral Swimmers
C0801762|T102|relax|37112-0|LNC|Knee X-ray AP lateral tunnel|Knee X-ray AP lateral tunnel
C0801762|T102|relax|37113-8|LNC|Knee bilateral X-ray AP lateral tunnel|Knee bilateral X-ray AP lateral tunnel
C0801762|T102|relax|37114-6|LNC|Knee left X-ray AP lateral tunnel|Knee left X-ray AP lateral tunnel
C0801762|T102|relax|37747-3|LNC|Knee right X-ray AP lateral tunnel|Knee right X-ray AP lateral tunnel
C0801762|T102|relax|69065-1|LNC|Abdomen X-ray AP lateral crosstable|Abdomen X-ray AP lateral crosstable
C0801762|T102|relax|37086-6|LNC|Hip X-ray AP lateral crosstable|Hip X-ray AP lateral crosstable
C0801762|T102|relax|37087-4|LNC|Hip left X-ray AP lateral crosstable|Hip left X-ray AP lateral crosstable
C0801762|T102|relax|37723-4|LNC|Hip right X-ray AP lateral crosstable|Hip right X-ray AP lateral crosstable
C0801762|T102|relax|37090-8|LNC|Knee X-ray AP lateral crosstable|Knee X-ray AP lateral crosstable
C0801762|T102|relax|69146-9|LNC|Knee left X-ray AP lateral crosstable|Knee left X-ray AP lateral crosstable
C0801762|T102|relax|37089-0|LNC|Pelvis Hip X-ray AP lateral crosstable|Pelvis Hip X-ray AP lateral crosstable
C0801762|T102|relax|37088-2|LNC|Pelvis Hip left X-ray AP lateral crosstable|Pelvis Hip left X-ray AP lateral crosstable
C0801762|T102|relax|38784-5|LNC|Pelvis Hip right X-ray AP lateral crosstable|Pelvis Hip right X-ray AP lateral crosstable
C0801762|T102|relax|30763-7|LNC|Abdomen X-ray AP lateral crosstable portable|Abdomen X-ray AP lateral crosstable portable
C0801762|T102|relax|37077-5|LNC|Hip X-ray AP lateral crosstable portable|Hip X-ray AP lateral crosstable portable
C0801762|T102|relax|37091-6|LNC|Hip X-ray AP lateral frog|Hip X-ray AP lateral frog
C0801762|T102|relax|37092-4|LNC|Hip bilateral X-ray AP lateral frog|Hip bilateral X-ray AP lateral frog
C0801762|T102|relax|37093-2|LNC|Hip left X-ray AP lateral frog|Hip left X-ray AP lateral frog
C0801762|T102|relax|37724-2|LNC|Hip right X-ray AP lateral frog|Hip right X-ray AP lateral frog
C0801762|T102|relax|30770-2|LNC|Pelvis Hip X-ray AP lateral frog|Pelvis Hip X-ray AP lateral frog
C0801762|T102|relax|42167-7|LNC|Pelvis Hip bilateral X-ray AP lateral frog|Pelvis Hip bilateral X-ray AP lateral frog
C0801762|T102|relax|37094-0|LNC|Pelvis Hip left X-ray AP lateral frog|Pelvis Hip left X-ray AP lateral frog
C0801762|T102|relax|38785-2|LNC|Pelvis Hip right X-ray AP lateral frog|Pelvis Hip right X-ray AP lateral frog
C0801762|T102|relax|41776-6|LNC|Pelvis Hip right X-ray AP lateral frog portable|Pelvis Hip right X-ray AP lateral frog portable
C0801762|T102|relax|24793-2|LNC|Abdomen X-ray AP lateral portable|Abdomen X-ray AP lateral portable
C0801762|T102|relax|44185-7|LNC|Femur X-ray AP lateral portable|Femur X-ray AP lateral portable
C0801762|T102|relax|44186-5|LNC|Foot X-ray AP lateral portable|Foot X-ray AP lateral portable
C0801762|T102|relax|41817-8|LNC|Hip left X-ray AP lateral portable|Hip left X-ray AP lateral portable
C0801762|T102|relax|41777-4|LNC|Hip right X-ray AP lateral portable|Hip right X-ray AP lateral portable
C0801762|T102|relax|30726-4|LNC|Spine Cervical X-ray AP lateral portable|Spine Cervical X-ray AP lateral portable
C0801762|T102|relax|37078-3|LNC|Spine Lumbar X-ray AP lateral portable|Spine Lumbar X-ray AP lateral portable
C0801762|T102|relax|30754-6|LNC|Spine Thoracic X-ray AP lateral portable|Spine Thoracic X-ray AP lateral portable
C0801762|T102|relax|39330-6|LNC|Ankle bilateral X-ray AP lateral standing|Ankle bilateral X-ray AP lateral standing
C0801762|T102|relax|42380-6|LNC|Ankle left X-ray AP lateral standing|Ankle left X-ray AP lateral standing
C0801762|T102|relax|39368-6|LNC|Ankle right X-ray AP lateral standing|Ankle right X-ray AP lateral standing
C0801762|T102|relax|39068-2|LNC|Foot X-ray AP lateral standing|Foot X-ray AP lateral standing
C0801762|T102|relax|39331-4|LNC|Foot bilateral X-ray AP lateral standing|Foot bilateral X-ray AP lateral standing
C0801762|T102|relax|39332-2|LNC|Foot left X-ray AP lateral standing|Foot left X-ray AP lateral standing
C0801762|T102|relax|39374-4|LNC|Foot right X-ray AP lateral standing|Foot right X-ray AP lateral standing
C0801762|T102|relax|24805-4|LNC|Knee X-ray AP lateral standing|Knee X-ray AP lateral standing
C0801762|T102|relax|26364-0|LNC|Knee bilateral X-ray AP lateral standing|Knee bilateral X-ray AP lateral standing
C0801762|T102|relax|26365-7|LNC|Knee left X-ray AP lateral standing|Knee left X-ray AP lateral standing
C0801762|T102|relax|26366-5|LNC|Knee right X-ray AP lateral standing|Knee right X-ray AP lateral standing
C0801762|T102|relax|39333-0|LNC|Spine Lumbar X-ray AP lateral standing|Spine Lumbar X-ray AP lateral standing
C0801762|T102|relax|38084-0|LNC|Abdomen X-ray AP left posterior oblique|Abdomen X-ray AP left posterior oblique
C0801762|T102|relax|37119-5|LNC|Abdomen X-ray AP oblique|Abdomen X-ray AP oblique
C0801762|T102|relax|39076-5|LNC|Foot X-ray AP oblique|Foot X-ray AP oblique
C0801762|T102|relax|37621-0|LNC|Pelvis X-ray AP oblique|Pelvis X-ray AP oblique
C0801762|T102|relax|37649-1|LNC|Sacroiliac Joint X-ray AP oblique|Sacroiliac Joint X-ray AP oblique
C0801762|T102|relax|39075-7|LNC|Toes X-ray AP oblique|Toes X-ray AP oblique
C0801762|T102|relax|37098-1|LNC|Spine Cervical X-ray AP oblique lateral W flexion W extension|Spine Cervical X-ray AP oblique lateral W flexion W extension
C0801762|T102|relax|44187-3|LNC|Spine Cervical X-ray AP oblique odontoid lateral portable W flexion W extension|Spine Cervical X-ray AP oblique odontoid lateral portable W flexion W extension
C0801762|T102|relax|37100-5|LNC|Spine Cervical X-ray AP oblique odontoid lateral W flexion W extension|Spine Cervical X-ray AP oblique odontoid lateral W flexion W extension
C0801762|T102|relax|24797-3|LNC|Abdomen X-ray AP oblique prone|Abdomen X-ray AP oblique prone
C0801762|T102|relax|37120-3|LNC|Spine Cervical X-ray AP odontoid lateral crosstable|Spine Cervical X-ray AP odontoid lateral crosstable
C0801762|T102|relax|37104-7|LNC|Spine Cervical X-ray AP odontoid lateral W flexion W extension|Spine Cervical X-ray AP odontoid lateral W flexion W extension
C0801762|T102|relax|42011-7|LNC|Chest Abdomen X-ray AP PA chest|Chest Abdomen X-ray AP PA chest
C0801762|T102|relax|24642-1|LNC|Chest X-ray AP PA upright|Chest X-ray AP PA upright
C0801762|T102|relax|24808-8|LNC|Knee X-ray AP PA standing|Knee X-ray AP PA standing
C0801762|T102|relax|26361-6|LNC|Knee bilateral X-ray AP PA standing|Knee bilateral X-ray AP PA standing
C0801762|T102|relax|26362-4|LNC|Knee left X-ray AP PA standing|Knee left X-ray AP PA standing
C0801762|T102|relax|26363-2|LNC|Knee right X-ray AP PA standing|Knee right X-ray AP PA standing
C0801762|T102|relax|37121-1|LNC|Clavicle left X-ray AP Serendipity|Clavicle left X-ray AP Serendipity
C0801762|T102|relax|37680-6|LNC|Clavicle right X-ray AP Serendipity|Clavicle right X-ray AP Serendipity
C0801762|T102|relax|37122-9|LNC|Shoulder left X-ray AP Stryker Notch|Shoulder left X-ray AP Stryker Notch
C0801762|T102|relax|37797-8|LNC|Shoulder right X-ray AP Stryker Notch|Shoulder right X-ray AP Stryker Notch
C0801762|T102|relax|37485-0|LNC|Humerus X-ray AP transthoracic|Humerus X-ray AP transthoracic
C0801762|T102|relax|39077-3|LNC|Shoulder X-ray AP transthoracic|Shoulder X-ray AP transthoracic
C0801762|T102|relax|46349-7|LNC|Shoulder bilateral X-ray AP transthoracic|Shoulder bilateral X-ray AP transthoracic
C0801762|T102|relax|38082-4|LNC|Shoulder left X-ray AP transthoracic|Shoulder left X-ray AP transthoracic
C0801762|T102|relax|38822-3|LNC|Shoulder right X-ray AP transthoracic|Shoulder right X-ray AP transthoracic
C0801762|T102|relax|37123-7|LNC|Shoulder left X-ray AP West Point|Shoulder left X-ray AP West Point
C0801762|T102|relax|38787-8|LNC|Shoulder right X-ray AP West Point|Shoulder right X-ray AP West Point
C0801762|T102|relax|36961-1|LNC|Shoulder left X-ray AP West Point outlet|Shoulder left X-ray AP West Point outlet
C0801762|T102|relax|37799-4|LNC|Shoulder right X-ray AP West Point outlet|Shoulder right X-ray AP West Point outlet
C0801762|T102|relax|37124-5|LNC|Scapula left X-ray AP Y|Scapula left X-ray AP Y
C0801762|T102|relax|37789-5|LNC|Scapula right X-ray AP Y|Scapula right X-ray AP Y
C0801762|T102|relax|69266-5|LNC|Shoulder X-ray AP Y|Shoulder X-ray AP Y
C0801762|T102|relax|37125-2|LNC|Shoulder left X-ray AP Y|Shoulder left X-ray AP Y
C0801762|T102|relax|38788-6|LNC|Shoulder right X-ray AP Y|Shoulder right X-ray AP Y
C0801762|T102|relax|24562-1|LNC|Abdomen X-ray AP (left lateral-decubitus right lateral-decubitus)|Abdomen X-ray AP (left lateral-decubitus right lateral-decubitus)
C0801762|T102|relax|24650-4|LNC|Chest X-ray AP (right lateral-decubitus left lateral-decubitus)|Chest X-ray AP (right lateral-decubitus left lateral-decubitus)
C0801762|T102|relax|24649-6|LNC|Chest X-ray AP (right lateral-decubitus left lateral-decubitus) portable|Chest X-ray AP (right lateral-decubitus left lateral-decubitus) portable
C0801762|T102|relax|37085-8|LNC|Abdomen X-ray AP (supine lateral-decubitus)|Abdomen X-ray AP (supine lateral-decubitus)
C0801762|T102|relax|37076-7|LNC|Abdomen X-ray AP (supine lateral-decubitus) portable|Abdomen X-ray AP (supine lateral-decubitus) portable
C0801762|T102|relax|24798-1|LNC|Abdomen X-ray AP (supine upright)|Abdomen X-ray AP (supine upright)
C0801762|T102|relax|43463-9|LNC|Chest Abdomen X-ray AP (supine upright) PA chest|Chest Abdomen X-ray AP (supine upright) PA chest
C0801762|T102|relax|24795-7|LNC|Abdomen X-ray AP (supine upright) portable|Abdomen X-ray AP (supine upright) portable
C0801762|T102|relax|42019-0|LNC|Abdomen X-ray AP (upright left lateral decubitus)|Abdomen X-ray AP (upright left lateral decubitus)
C0801762|T102|relax|39329-8|LNC|Shoulder bilateral X-ray AP (W internal rotation W external rotation)|Shoulder bilateral X-ray AP (W internal rotation W external rotation)
C0801762|T102|relax|39328-0|LNC|Shoulder left X-ray AP (W internal rotation W external rotation)|Shoulder left X-ray AP (W internal rotation W external rotation)
C0801762|T102|relax|39395-9|LNC|Shoulder right X-ray AP (W internal rotation W external rotation)|Shoulder right X-ray AP (W internal rotation W external rotation)
C0801762|T102|relax|39321-5|LNC|Shoulder X-ray AP (W internal rotation W external rotation) axillary|Shoulder X-ray AP (W internal rotation W external rotation) axillary
C0801762|T102|relax|39336-3|LNC|Shoulder bilateral X-ray AP (W internal rotation W external rotation) axillary|Shoulder bilateral X-ray AP (W internal rotation W external rotation) axillary
C0801762|T102|relax|39335-5|LNC|Shoulder left X-ray AP (W internal rotation W external rotation) axillary|Shoulder left X-ray AP (W internal rotation W external rotation) axillary
C0801762|T102|relax|39337-1|LNC|Shoulder bilateral X-ray AP (W internal rotation W external rotation) axillary outlet|Shoulder bilateral X-ray AP (W internal rotation W external rotation) axillary outlet
C0801762|T102|relax|39344-7|LNC|Shoulder bilateral X-ray AP (W internal rotation W external rotation) axillary Y|Shoulder bilateral X-ray AP (W internal rotation W external rotation) axillary Y
C0801762|T102|relax|39338-9|LNC|Shoulder left X-ray AP (W internal rotation W external rotation) axillary Y|Shoulder left X-ray AP (W internal rotation W external rotation) axillary Y
C0801762|T102|relax|39397-5|LNC|Shoulder right X-ray AP (W internal rotation W external rotation) West Point|Shoulder right X-ray AP (W internal rotation W external rotation) West Point
C0801762|T102|relax|39343-9|LNC|Shoulder bilateral X-ray AP (W internal rotation W external rotation) Y|Shoulder bilateral X-ray AP (W internal rotation W external rotation) Y
C0801762|T102|relax|39348-8|LNC|Shoulder left X-ray AP (W internal rotation W external rotation) Y|Shoulder left X-ray AP (W internal rotation W external rotation) Y
C0801762|T102|relax|39325-6|LNC|Shoulder left X-ray AP (W internal rotation) Grashey axillary outlet|Shoulder left X-ray AP (W internal rotation) Grashey axillary outlet
C0801762|T102|relax|39346-2|LNC|Shoulder bilateral X-ray AP (W internal rotation) West Point|Shoulder bilateral X-ray AP (W internal rotation) West Point
C0801762|T102|relax|39347-0|LNC|Shoulder left X-ray AP (W internal rotation) West Point|Shoulder left X-ray AP (W internal rotation) West Point
C0801762|T102|relax|39396-7|LNC|Shoulder right X-ray AP (W internal rotation) West Point|Shoulder right X-ray AP (W internal rotation) West Point
C0801762|T102|relax|24632-2|LNC|Chest X-ray AP portable|Chest X-ray AP portable
C0801762|T102|relax|37075-9|LNC|Hip X-ray AP portable|Hip X-ray AP portable
C0801762|T102|relax|43561-0|LNC|Chest Abdomen X-ray AP upright AP chest|Chest Abdomen X-ray AP upright AP chest
C0801762|T102|relax|38003-0|LNC|Foot left X-ray AP standing|Foot left X-ray AP standing
C0801762|T102|relax|38815-7|LNC|Foot right X-ray AP standing|Foot right X-ray AP standing
C0801762|T102|relax|42406-9|LNC|Spine Lumbar X-ray AP W WO left bending|Spine Lumbar X-ray AP W WO left bending
C0801762|T102|relax|42407-7|LNC|Spine Lumbar X-ray AP W WO right bending|Spine Lumbar X-ray AP W WO right bending
C0801762|T102|relax|42445-7|LNC|Spine Thoracic X-ray AP W left bending WO bending|Spine Thoracic X-ray AP W left bending WO bending
C0801762|T102|relax|37484-3|LNC|Knee left X-ray AP W manual stress|Knee left X-ray AP W manual stress
C0801762|T102|relax|37746-5|LNC|Knee right X-ray AP W manual stress|Knee right X-ray AP W manual stress
C0801762|T102|relax|42403-6|LNC|Spine Lumbar X-ray AP W right bending W left bending|Spine Lumbar X-ray AP W right bending W left bending
C0801762|T102|relax|42408-5|LNC|Spine Lumbar X-ray AP W right bending W left bending WO bending|Spine Lumbar X-ray AP W right bending W left bending WO bending
C0801762|T102|relax|42444-0|LNC|Spine Thoracic X-ray AP W right bending W left bending WO bending|Spine Thoracic X-ray AP W right bending W left bending WO bending
C0801762|T102|relax|42446-5|LNC|Spine Thoracic X-ray AP W right bending WO bending|Spine Thoracic X-ray AP W right bending WO bending
C0801762|T102|relax|39403-1|LNC|Shoulder X-ray axillary transcapular|Shoulder X-ray axillary transcapular
C0801762|T102|relax|37127-8|LNC|Shoulder bilateral X-ray axillary Y|Shoulder bilateral X-ray axillary Y
C0801762|T102|relax|37128-6|LNC|Shoulder left X-ray axillary Y|Shoulder left X-ray axillary Y
C0801762|T102|relax|37807-5|LNC|Shoulder right X-ray axillary Y|Shoulder right X-ray axillary Y
C0801762|T102|relax|46386-9|LNC|Teeth X-ray bitewing|Teeth X-ray bitewing
C0801762|T102|relax|39884-2|LNC|Bone Scan blood pool|Bone Scan blood pool
C0801762|T102|relax|39861-0|LNC|Heart Scan blood pool|Heart Scan blood pool
C0801762|T102|relax|42709-6|LNC|Liver Scan blood pool|Liver Scan blood pool
C0801762|T102|relax|39860-2|LNC|Heart Scan blood pool W stress W radionuclide IV|Heart Scan blood pool W stress W radionuclide IV
C0801762|T102|relax|26352-5|LNC|Wrist bilateral Hand bilateral X-ray bone age|Wrist bilateral Hand bilateral X-ray bone age
C0801762|T102|relax|26353-3|LNC|Wrist left Hand left X-ray bone age|Wrist left Hand left X-ray bone age
C0801762|T102|relax|26354-1|LNC|Wrist right Hand right X-ray bone age|Wrist right Hand right X-ray bone age
C0801762|T102|relax|24724-7|LNC|Wrist Hand X-ray bone age|Wrist Hand X-ray bone age
C0801762|T102|relax|37362-1|LNC|Bones X-ray bone age|Bones X-ray bone age
C0801762|T102|relax|24591-0|LNC|Brain Scan brain death protocol W Tc-99m HMPAO IV|Brain Scan brain death protocol W Tc-99m HMPAO IV
C0801762|T102|relax|37996-6|LNC|Calcaneus X-ray Broden|Calcaneus X-ray Broden
C0801762|T102|relax|37995-8|LNC|Calcaneus bilateral X-ray Broden|Calcaneus bilateral X-ray Broden
C0801762|T102|relax|37997-4|LNC|Calcaneus left X-ray Broden|Calcaneus left X-ray Broden
C0801762|T102|relax|38814-0|LNC|Calcaneus right X-ray Broden|Calcaneus right X-ray Broden
C0801762|T102|relax|37486-8|LNC|Ankle X-ray Broden W manual stress|Ankle X-ray Broden W manual stress
C0801762|T102|relax|37852-1|LNC|Sinuses X-ray Caldwell Waters|Sinuses X-ray Caldwell Waters
C0801762|T102|relax|39859-4|LNC|Brain Scan delayed static|Brain Scan delayed static
C0801762|T102|relax|39875-0|LNC|Scan delayed W GA-67 IV|Scan delayed W GA-67 IV
C0801762|T102|relax|39840-4|LNC|Scan delayed W I-131 MIBG IV|Scan delayed W I-131 MIBG IV
C0801762|T102|relax|39842-0|LNC|Scan delayed W In-111 Satumomab IV|Scan delayed W In-111 Satumomab IV
C0801762|T102|relax|39874-3|LNC|Head Cistern Scan delayed W radionuclide IT|Head Cistern Scan delayed W radionuclide IT
C0801762|T102|relax|39819-8|LNC|Bone Scan delayed|Bone Scan delayed
C0801762|T102|relax|39741-4|LNC|Parathyroid Scan delayed|Parathyroid Scan delayed
C0801762|T102|relax|24605-8|LNC|Breast Mammogram diagnostic|Breast Mammogram diagnostic
C0801762|T102|relax|39152-4|LNC|Breast FFD mammogram diagnostic|Breast FFD mammogram diagnostic
C0801762|T102|relax|69158-4|LNC|Breast implant X-ray diagnostic|Breast implant X-ray diagnostic
C0801762|T102|relax|48475-8|LNC|Breast implant bilateral Mammogram diagnostic|Breast implant bilateral Mammogram diagnostic
C0801762|T102|relax|69150-1|LNC|Breast implant left Mammogram diagnostic|Breast implant left Mammogram diagnostic
C0801762|T102|relax|69259-0|LNC|Breast implant right Mammogram diagnostic|Breast implant right Mammogram diagnostic
C0801762|T102|relax|26346-7|LNC|Breast bilateral Mammogram diagnostic|Breast bilateral Mammogram diagnostic
C0801762|T102|relax|39154-0|LNC|Breast bilateral FFD mammogram diagnostic|Breast bilateral FFD mammogram diagnostic
C0801762|T102|relax|26347-5|LNC|Breast left Mammogram diagnostic|Breast left Mammogram diagnostic
C0801762|T102|relax|42169-3|LNC|Breast left FFD mammogram diagnostic|Breast left FFD mammogram diagnostic
C0801762|T102|relax|26348-3|LNC|Breast right Mammogram diagnostic|Breast right Mammogram diagnostic
C0801762|T102|relax|42168-5|LNC|Breast right FFD mammogram diagnostic|Breast right FFD mammogram diagnostic
C0801762|T102|relax|46350-5|LNC|Breast unilateral Mammogram diagnostic|Breast unilateral Mammogram diagnostic
C0801762|T102|relax|24604-1|LNC|Breast Mammogram diagnostic limited|Breast Mammogram diagnostic limited
C0801762|T102|relax|26349-1|LNC|Breast bilateral Mammogram diagnostic limited|Breast bilateral Mammogram diagnostic limited
C0801762|T102|relax|26350-9|LNC|Breast left Mammogram diagnostic limited|Breast left Mammogram diagnostic limited
C0801762|T102|relax|26351-7|LNC|Breast right Mammogram diagnostic limited|Breast right Mammogram diagnostic limited
C0801762|T102|relax|46351-3|LNC|Breast implant bilateral Mammogram displacement|Breast implant bilateral Mammogram displacement
C0801762|T102|relax|39895-8|LNC|Gallbladder Scan ejection fraction W Tc-99m DISIDA IV|Gallbladder Scan ejection fraction W Tc-99m DISIDA IV
C0801762|T102|relax|39887-5|LNC|Heart Scan first pass ejection fraction at rest W radionuclide IV|Heart Scan first pass ejection fraction at rest W radionuclide IV
C0801762|T102|relax|39889-1|LNC|Heart Scan first pass ejection fraction|Heart Scan first pass ejection fraction
C0801762|T102|relax|39885-9|LNC|Heart Scan first pass ventricular volume|Heart Scan first pass ventricular volume
C0801762|T102|relax|39910-5|LNC|Heart Scan first pass wall motion ejection fraction|Heart Scan first pass wall motion ejection fraction
C0801762|T102|relax|39912-1|LNC|Heart Scan first pass wall motion ventricular volume ejection fraction|Heart Scan first pass wall motion ventricular volume ejection fraction
C0801762|T102|relax|39909-7|LNC|Heart Scan first pass wall motion ventricular volume ejection fraction W stress W radionuclide IV|Heart Scan first pass wall motion ventricular volume ejection fraction W stress W radionuclide IV
C0801762|T102|relax|39908-9|LNC|Heart Scan first pass wall motion ventricular volume W stress W radionuclide IV|Heart Scan first pass wall motion ventricular volume W stress W radionuclide IV
C0801762|T102|relax|39886-7|LNC|Heart Scan first pass wall motion at rest W radionuclide IV|Heart Scan first pass wall motion at rest W radionuclide IV
C0801762|T102|relax|39890-9|LNC|Heart Scan first pass wall motion|Heart Scan first pass wall motion
C0801762|T102|relax|39888-3|LNC|Heart Scan first pass wall motion W stress W radionuclide IV|Heart Scan first pass wall motion W stress W radionuclide IV
C0801762|T102|relax|39867-7|LNC|Heart Scan first pass at rest W radionuclide IV|Heart Scan first pass at rest W radionuclide IV
C0801762|T102|relax|39863-6|LNC|Heart Scan first pass at rest W stress W radionuclide IV|Heart Scan first pass at rest W stress W radionuclide IV
C0801762|T102|relax|39866-9|LNC|Heart Scan first pass at rest W Tc-99m Sestamibi IV|Heart Scan first pass at rest W Tc-99m Sestamibi IV
C0801762|T102|relax|39864-4|LNC|Heart Scan first pass|Heart Scan first pass
C0801762|T102|relax|39865-1|LNC|Left ventricle Scan first pass|Left ventricle Scan first pass
C0801762|T102|relax|39869-3|LNC|Heart Scan first pass W stress W radionuclide IV|Heart Scan first pass W stress W radionuclide IV
C0801762|T102|relax|39868-5|LNC|Heart Scan first pass W stress W Tc-99m Sestamibi IV|Heart Scan first pass W stress W Tc-99m Sestamibi IV
C0801762|T102|relax|39893-3|LNC|Heart Scan flow shunt detection|Heart Scan flow shunt detection
C0801762|T102|relax|43644-4|LNC|Brain Scan flow limited|Brain Scan flow limited
C0801762|T102|relax|39858-6|LNC|Bone Scan flow|Bone Scan flow
C0801762|T102|relax|39636-6|LNC|Brain Scan flow|Brain Scan flow
C0801762|T102|relax|39871-9|LNC|Heart Scan flow|Heart Scan flow
C0801762|T102|relax|42261-8|LNC|Kidney bilateral Scan flow|Kidney bilateral Scan flow
C0801762|T102|relax|42262-6|LNC|Liver Scan flow|Liver Scan flow
C0801762|T102|relax|43653-5|LNC|Liver Spleen Scan flow|Liver Spleen Scan flow
C0801762|T102|relax|39847-9|LNC|Parotid gland Scan flow|Parotid gland Scan flow
C0801762|T102|relax|39899-0|LNC|Salivary gland Scan flow|Salivary gland Scan flow
C0801762|T102|relax|42308-7|LNC|Scrotum Testicle Scan flow|Scrotum Testicle Scan flow
C0801762|T102|relax|42263-4|LNC|Spleen Scan flow|Spleen Scan flow
C0801762|T102|relax|39856-0|LNC|Thyroid Scan flow|Thyroid Scan flow
C0801762|T102|relax|43500-8|LNC|Vessel Scan flow|Vessel Scan flow
C0801762|T102|relax|44148-5|LNC|Brain Scan flow W Tc-99m bicisate IV|Brain Scan flow W Tc-99m bicisate IV
C0801762|T102|relax|43642-8|LNC|Brain Scan flow W Tc-99m DTPA IV|Brain Scan flow W Tc-99m DTPA IV
C0801762|T102|relax|43664-2|LNC|Renal vessels Scan flow W Tc-99m DTPA IV|Renal vessels Scan flow W Tc-99m DTPA IV
C0801762|T102|relax|43643-6|LNC|Brain Scan flow W Tc-99m glucoheptonate IV|Brain Scan flow W Tc-99m glucoheptonate IV
C0801762|T102|relax|43666-7|LNC|Kidney bilateral Renal vessels Scan flow W Tc-99m glucoheptonate IV|Kidney bilateral Renal vessels Scan flow W Tc-99m glucoheptonate IV
C0801762|T102|relax|43663-4|LNC|Renal vessels Scan flow W Tc-99m glucoheptonate IV|Renal vessels Scan flow W Tc-99m glucoheptonate IV
C0801762|T102|relax|43665-9|LNC|Renal vessels Scan flow W Tc-99m Mertiatide IV|Renal vessels Scan flow W Tc-99m Mertiatide IV
C0801762|T102|relax|39870-1|LNC|Heart Scan flow W Tc-99m pertechnetate IV|Heart Scan flow W Tc-99m pertechnetate IV
C0801762|T102|relax|43654-3|LNC|Liver Scan flow W Tc-99m tagged RBC IV|Liver Scan flow W Tc-99m tagged RBC IV
C0801762|T102|relax|39685-3|LNC|Scan abscess W GA-67 IV|Scan abscess W GA-67 IV
C0801762|T102|relax|39940-2|LNC|Lung Scan Clearance W Tc-99m DTPA aerosol inhaled|Lung Scan Clearance W Tc-99m DTPA aerosol inhaled
C0801762|T102|relax|43787-1|LNC|Skull Facial bones Mandible X-ray dental measurement|Skull Facial bones Mandible X-ray dental measurement
C0801762|T102|relax|43648-5|LNC|Scan endocrine tumor multiple areas W I-131 MIBG IV|Scan endocrine tumor multiple areas W I-131 MIBG IV
C0801762|T102|relax|43649-3|LNC|Scan endocrine tumor multiple areas W In-111 pentetreotide IV|Scan endocrine tumor multiple areas W In-111 pentetreotide IV
C0801762|T102|relax|39827-1|LNC|Scan endocrine tumor whole body W I-131 MIBG IV|Scan endocrine tumor whole body W I-131 MIBG IV
C0801762|T102|relax|39828-9|LNC|Scan endocrine tumor whole body W In-111 pentetreotide IV|Scan endocrine tumor whole body W In-111 pentetreotide IV
C0801762|T102|relax|39327-2|LNC|Abdomen Fetus X-ray fetal age|Abdomen Fetus X-ray fetal age
C0801762|T102|relax|44208-7|LNC|Orbit X-ray foreign body|Orbit X-ray foreign body
C0801762|T102|relax|30720-7|LNC|Orbit bilateral X-ray foreign body|Orbit bilateral X-ray foreign body
C0801762|T102|relax|42311-1|LNC|Orbit left X-ray foreign body|Orbit left X-ray foreign body
C0801762|T102|relax|42312-9|LNC|Orbit right X-ray foreign body|Orbit right X-ray foreign body
C0801762|T102|relax|39768-7|LNC|Stomach Scan gastric emptying W Tc-99m SC PO|Stomach Scan gastric emptying W Tc-99m SC PO
C0801762|T102|relax|39767-9|LNC|Stomach Scan gastric emptying liquid phase W radionuclide PO|Stomach Scan gastric emptying liquid phase W radionuclide PO
C0801762|T102|relax|24997-9|LNC|Stomach Scan gastric emptying solid phase W Tc-99m SC PO|Stomach Scan gastric emptying solid phase W Tc-99m SC PO
C0801762|T102|relax|39769-5|LNC|Stomach Scan gastric emptying W radionuclide PO|Stomach Scan gastric emptying W radionuclide PO
C0801762|T102|relax|39892-5|LNC|Heart Scan infarct first pass|Heart Scan infarct first pass
C0801762|T102|relax|39891-7|LNC|Heart Scan infarct first pass W Tc-99m PYP IV|Heart Scan infarct first pass W Tc-99m PYP IV
C0801762|T102|relax|43646-9|LNC|Heart Scan infarct qualitative quantitative|Heart Scan infarct qualitative quantitative
C0801762|T102|relax|43645-1|LNC|Heart Scan infarct qualitative|Heart Scan infarct qualitative
C0801762|T102|relax|43647-7|LNC|Heart Scan infarct quantitative|Heart Scan infarct quantitative
C0801762|T102|relax|39653-1|LNC|Heart Scan infarct|Heart Scan infarct
C0801762|T102|relax|39657-2|LNC|Heart Scan infarct W Tc-99m PYP IV|Heart Scan infarct W Tc-99m PYP IV
C0801762|T102|relax|39933-7|LNC|Scan infection multiple areas W GA-67 IV|Scan infection multiple areas W GA-67 IV
C0801762|T102|relax|39830-5|LNC|Scan infection whole body W GA-67 IV|Scan infection whole body W GA-67 IV
C0801762|T102|relax|39677-0|LNC|Scan infection W GA-67 IV|Scan infection W GA-67 IV
C0801762|T102|relax|39490-8|LNC|Femur right Tibia right X-ray leg length|Femur right Tibia right X-ray leg length
C0801762|T102|relax|24700-7|LNC|Femur Tibia X-ray leg length|Femur Tibia X-ray leg length
C0801762|T102|relax|39686-1|LNC|Scan lymphoma W GA-67 IV|Scan lymphoma W GA-67 IV
C0801762|T102|relax|42170-1|LNC|Scan lymphoma|Scan lymphoma
C0801762|T102|relax|39672-1|LNC|Esophagus Scan motility W radionuclide PO|Esophagus Scan motility W radionuclide PO
C0801762|T102|relax|72256-1|LNC|Abdomen X-ray motility with radioopaque markers|Abdomen X-ray motility with radioopaque markers
C0801762|T102|relax|24571-2|LNC|Biliary ducts Gallbladder Scan patency biliary structures ejection fraction W sincalide W radionuclide IV|Biliary ducts Gallbladder Scan patency biliary structures ejection fraction W sincalide W radionuclide IV
C0801762|T102|relax|24572-0|LNC|Biliary ducts Gallbladder Scan patency biliary structures W Tc-99m IV|Biliary ducts Gallbladder Scan patency biliary structures W Tc-99m IV
C0801762|T102|relax|43788-9|LNC|Tube Fluoroscopy patency W contrast via tube|Tube Fluoroscopy patency W contrast via tube
C0801762|T102|relax|43789-7|LNC|Liver Biliary ducts Gallbladder Scan patency W Tc-99m IV|Liver Biliary ducts Gallbladder Scan patency W Tc-99m IV
C0801762|T102|relax|39673-9|LNC|Esophagus Scan reflux W radionuclide PO|Esophagus Scan reflux W radionuclide PO
C0801762|T102|relax|30650-6|LNC|Unspecified body region Fluoroscopy shunt|Unspecified body region Fluoroscopy shunt
C0801762|T102|relax|39665-5|LNC|Heart Scan shunt detection|Heart Scan shunt detection
C0801762|T102|relax|39664-8|LNC|Heart Scan shunt detection W Tc-99m MAA IV|Heart Scan shunt detection W Tc-99m MAA IV
C0801762|T102|relax|39848-7|LNC|Peritoneovenous shunt Scan patency W In-111 IT|Peritoneovenous shunt Scan patency W In-111 IT
C0801762|T102|relax|39849-5|LNC|Peritoneovenous shunt Scan patency W radionuclide IT|Peritoneovenous shunt Scan patency W radionuclide IT
C0801762|T102|relax|24876-5|LNC|Peritoneovenous shunt Scan patency W Tc-99m DTPA IT|Peritoneovenous shunt Scan patency W Tc-99m DTPA IT
C0801762|T102|relax|44149-3|LNC|Peritoneovenous shunt Scan patency W Tc-99m MAA inj|Peritoneovenous shunt Scan patency W Tc-99m MAA inj
C0801762|T102|relax|39954-3|LNC|Vein Scan thrombosis|Vein Scan thrombosis
C0801762|T102|relax|44140-2|LNC|Abdomen Pelvis Scan tumor|Abdomen Pelvis Scan tumor
C0801762|T102|relax|39831-3|LNC|Scan tumor limited W GA-67 IV|Scan tumor limited W GA-67 IV
C0801762|T102|relax|39951-9|LNC|Scan tumor multiple area W Tc-99m Sestamibi IV|Scan tumor multiple area W Tc-99m Sestamibi IV
C0801762|T102|relax|39934-5|LNC|Scan tumor multiple areas W GA-67 IV|Scan tumor multiple areas W GA-67 IV
C0801762|T102|relax|39829-7|LNC|Scan tumor whole body W GA-67 IV|Scan tumor whole body W GA-67 IV
C0801762|T102|relax|42171-9|LNC|Scan tumor whole body|Scan tumor whole body
C0801762|T102|relax|39749-7|LNC|Scan tumor whole body W Tc-99m Sestamibi IV|Scan tumor whole body W Tc-99m Sestamibi IV
C0801762|T102|relax|39679-6|LNC|Scan tumor W GA-67 IV|Scan tumor W GA-67 IV
C0801762|T102|relax|39750-5|LNC|Scan tumor W Tc-99m Sestamibi IV|Scan tumor W Tc-99m Sestamibi IV
C0801762|T102|relax|42305-3|LNC|Scan tumor W Tl-201 IV|Scan tumor W Tl-201 IV
C0801762|T102|relax|42397-0|LNC|Chest X-ray frontal stereo|Chest X-ray frontal stereo
C0801762|T102|relax|39923-8|LNC|Heart Scan gated ejection fraction at rest W radionuclide IV|Heart Scan gated ejection fraction at rest W radionuclide IV
C0801762|T102|relax|39917-0|LNC|Heart Scan gated ejection fraction|Heart Scan gated ejection fraction
C0801762|T102|relax|39919-6|LNC|Heart Scan gated first pass|Heart Scan gated first pass
C0801762|T102|relax|39925-3|LNC|Heart Scan gated wall motion ejection fraction at rest W radionuclide IV|Heart Scan gated wall motion ejection fraction at rest W radionuclide IV
C0801762|T102|relax|39931-1|LNC|Heart Scan gated wall motion ejection fraction|Heart Scan gated wall motion ejection fraction
C0801762|T102|relax|42306-1|LNC|Heart Scan gated wall motion|Heart Scan gated wall motion
C0801762|T102|relax|39929-5|LNC|Heart Scan gated wall motion W stress W radionuclide IV|Heart Scan gated wall motion W stress W radionuclide IV
C0801762|T102|relax|39921-2|LNC|Heart Scan gated at rest W radionuclide IV|Heart Scan gated at rest W radionuclide IV
C0801762|T102|relax|39924-6|LNC|Heart Scan gated at rest W stress W radionuclide IV|Heart Scan gated at rest W stress W radionuclide IV
C0801762|T102|relax|39922-0|LNC|Heart Scan gated at rest W Tc-99m pertechnetate IV|Heart Scan gated at rest W Tc-99m pertechnetate IV
C0801762|T102|relax|39920-4|LNC|Heart Scan gated at rest W Tc-99m Sestamibi IV|Heart Scan gated at rest W Tc-99m Sestamibi IV
C0801762|T102|relax|39915-4|LNC|Heart Scan gated|Heart Scan gated
C0801762|T102|relax|39928-7|LNC|Heart Scan gated W stress W radionuclide IV|Heart Scan gated W stress W radionuclide IV
C0801762|T102|relax|39927-9|LNC|Heart Scan gated W stress W Tc-99m pertechnetate IV|Heart Scan gated W stress W Tc-99m pertechnetate IV
C0801762|T102|relax|39914-7|LNC|Heart Scan gated W Tc-99m Sestamibi IV|Heart Scan gated W Tc-99m Sestamibi IV
C0801762|T102|relax|46348-9|LNC|Chest X-ray GE 2 PA Lateral views|Chest X-ray GE 2 PA Lateral views
C0801762|T102|relax|44210-3|LNC|Ankle X-ray GE 3 views|Ankle X-ray GE 3 views
C0801762|T102|relax|48480-8|LNC|Ankle bilateral X-ray GE 3 views|Ankle bilateral X-ray GE 3 views
C0801762|T102|relax|46390-1|LNC|Ankle left X-ray GE 3 views|Ankle left X-ray GE 3 views
C0801762|T102|relax|46347-1|LNC|Ankle right X-ray GE 3 views|Ankle right X-ray GE 3 views
C0801762|T102|relax|48481-6|LNC|Elbow bilateral X-ray GE 3 views|Elbow bilateral X-ray GE 3 views
C0801762|T102|relax|46344-8|LNC|Elbow left X-ray GE 3 views|Elbow left X-ray GE 3 views
C0801762|T102|relax|46345-5|LNC|Elbow right X-ray GE 3 views|Elbow right X-ray GE 3 views
C0801762|T102|relax|48479-0|LNC|Facial bones X-ray GE 3 views|Facial bones X-ray GE 3 views
C0801762|T102|relax|43492-8|LNC|Finger fifth left X-ray GE 3 views|Finger fifth left X-ray GE 3 views
C0801762|T102|relax|43497-7|LNC|Finger fifth right X-ray GE 3 views|Finger fifth right X-ray GE 3 views
C0801762|T102|relax|43491-0|LNC|Finger fourth left X-ray GE 3 views|Finger fourth left X-ray GE 3 views
C0801762|T102|relax|43496-9|LNC|Finger fourth right X-ray GE 3 views|Finger fourth right X-ray GE 3 views
C0801762|T102|relax|43489-4|LNC|Finger second left X-ray GE 3 views|Finger second left X-ray GE 3 views
C0801762|T102|relax|43494-4|LNC|Finger second right X-ray GE 3 views|Finger second right X-ray GE 3 views
C0801762|T102|relax|43490-2|LNC|Finger third left X-ray GE 3 views|Finger third left X-ray GE 3 views
C0801762|T102|relax|43495-1|LNC|Finger third right X-ray GE 3 views|Finger third right X-ray GE 3 views
C0801762|T102|relax|44188-1|LNC|Foot X-ray GE 3 views|Foot X-ray GE 3 views
C0801762|T102|relax|48478-2|LNC|Foot bilateral X-ray GE 3 views|Foot bilateral X-ray GE 3 views
C0801762|T102|relax|48477-4|LNC|Foot left X-ray GE 3 views|Foot left X-ray GE 3 views
C0801762|T102|relax|48476-6|LNC|Foot right X-ray GE 3 views|Foot right X-ray GE 3 views
C0801762|T102|relax|47370-2|LNC|Hand left X-ray GE 3 views|Hand left X-ray GE 3 views
C0801762|T102|relax|47371-0|LNC|Hand right X-ray GE 3 views|Hand right X-ray GE 3 views
C0801762|T102|relax|43498-5|LNC|Knee left X-ray GE 3 views|Knee left X-ray GE 3 views
C0801762|T102|relax|43482-9|LNC|Knee right X-ray GE 3 views|Knee right X-ray GE 3 views
C0801762|T102|relax|47381-9|LNC|Mastoid X-ray GE 3 views|Mastoid X-ray GE 3 views
C0801762|T102|relax|43543-8|LNC|Pelvis X-ray GE 3 views|Pelvis X-ray GE 3 views
C0801762|T102|relax|44189-9|LNC|Sacroiliac Joint X-ray GE 3 views|Sacroiliac Joint X-ray GE 3 views
C0801762|T102|relax|48746-2|LNC|Sacroiliac joint bilateral X-ray GE 3 views|Sacroiliac joint bilateral X-ray GE 3 views
C0801762|T102|relax|43486-0|LNC|Sinuses X-ray GE 3 views|Sinuses X-ray GE 3 views
C0801762|T102|relax|46377-8|LNC|Skull X-ray GE 3 views|Skull X-ray GE 3 views
C0801762|T102|relax|48482-4|LNC|Sternoclavicular Joints X-ray GE 3 views|Sternoclavicular Joints X-ray GE 3 views
C0801762|T102|relax|43488-6|LNC|Thumb left X-ray GE 3 views|Thumb left X-ray GE 3 views
C0801762|T102|relax|43493-6|LNC|Thumb right X-ray GE 3 views|Thumb right X-ray GE 3 views
C0801762|T102|relax|44190-7|LNC|Wrist X-ray GE 3 views|Wrist X-ray GE 3 views
C0801762|T102|relax|48483-2|LNC|Wrist bilateral X-ray GE 3 views|Wrist bilateral X-ray GE 3 views
C0801762|T102|relax|46346-3|LNC|Wrist left X-ray GE 3 views|Wrist left X-ray GE 3 views
C0801762|T102|relax|46343-0|LNC|Wrist right X-ray GE 3 views|Wrist right X-ray GE 3 views
C0801762|T102|relax|48485-7|LNC|Ribs bilateral Chest X-ray GE 3 PA Chest views|Ribs bilateral Chest X-ray GE 3 PA Chest views
C0801762|T102|relax|48486-5|LNC|Ribs left Chest X-ray GE 3 PA Chest views|Ribs left Chest X-ray GE 3 PA Chest views
C0801762|T102|relax|48484-0|LNC|Ribs right Chest X-ray GE 3 PA Chest views|Ribs right Chest X-ray GE 3 PA Chest views
C0801762|T102|relax|44191-5|LNC|Ribs Chest X-ray GE 3 PA Chest views|Ribs Chest X-ray GE 3 PA Chest views
C0801762|T102|relax|44239-2|LNC|Ribs unilateral Chest X-ray Ge 3 PA Chest Portable views|Ribs unilateral Chest X-ray Ge 3 PA Chest Portable views
C0801762|T102|relax|44193-1|LNC|Hand X-ray GE 3 Portable views|Hand X-ray GE 3 Portable views
C0801762|T102|relax|44192-3|LNC|Pelvis X-ray GE 3 Portable views|Pelvis X-ray GE 3 Portable views
C0801762|T102|relax|44211-1|LNC|Chest X-ray GE 4 views|Chest X-ray GE 4 views
C0801762|T102|relax|47367-8|LNC|Chest Fluoroscopy GE 4 views|Chest Fluoroscopy GE 4 views
C0801762|T102|relax|47374-4|LNC|Knee left X-ray GE 4 views|Knee left X-ray GE 4 views
C0801762|T102|relax|47376-9|LNC|Knee right X-ray GE 4 views|Knee right X-ray GE 4 views
C0801762|T102|relax|47379-3|LNC|Mandible X-ray GE 4 views|Mandible X-ray GE 4 views
C0801762|T102|relax|48747-0|LNC|Orbit bilateral X-ray GE 4 views|Orbit bilateral X-ray GE 4 views
C0801762|T102|relax|48487-3|LNC|Skull X-ray GE 4 views|Skull X-ray GE 4 views
C0801762|T102|relax|44212-9|LNC|Spine Cervical X-ray GE 4 views|Spine Cervical X-ray GE 4 views
C0801762|T102|relax|47382-7|LNC|Spine Lumbar X-ray GE 4 views|Spine Lumbar X-ray GE 4 views
C0801762|T102|relax|47368-6|LNC|Chest X-ray GE 4 Pa Lateral views|Chest X-ray GE 4 Pa Lateral views
C0801762|T102|relax|44194-9|LNC|Spine X-ray GE 4 views W right bending W left bending|Spine X-ray GE 4 views W right bending W left bending
C0801762|T102|relax|44195-6|LNC|Knee X-ray GE 5 views|Knee X-ray GE 5 views
C0801762|T102|relax|43524-8|LNC|Skull X-ray GE 5 views|Skull X-ray GE 5 views
C0801762|T102|relax|44197-2|LNC|Knee bilateral X-ray GE 5 views standing|Knee bilateral X-ray GE 5 views standing
C0801762|T102|relax|44196-4|LNC|Spine Lumbar X-ray GE 5 views W right bending W left bending|Spine Lumbar X-ray GE 5 views W right bending W left bending
C0801762|T102|relax|49570-5|LNC|Ankle bilateral X-ray GE 6 views|Ankle bilateral X-ray GE 6 views
C0801762|T102|relax|37160-9|LNC|Shoulder left X-ray Grashey axillary|Shoulder left X-ray Grashey axillary
C0801762|T102|relax|38793-6|LNC|Shoulder right X-ray Grashey axillary|Shoulder right X-ray Grashey axillary
C0801762|T102|relax|37158-3|LNC|Shoulder left X-ray Grashey axillary outlet|Shoulder left X-ray Grashey axillary outlet
C0801762|T102|relax|37806-7|LNC|Shoulder right X-ray Grashey axillary outlet|Shoulder right X-ray Grashey axillary outlet
C0801762|T102|relax|37161-7|LNC|Shoulder bilateral X-ray Grashey axillary outlet Zanca|Shoulder bilateral X-ray Grashey axillary outlet Zanca
C0801762|T102|relax|69267-3|LNC|Shoulder X-ray Grashey axillary Y|Shoulder X-ray Grashey axillary Y
C0801762|T102|relax|37538-6|LNC|Shoulder left X-ray Grashey axillary Y|Shoulder left X-ray Grashey axillary Y
C0801762|T102|relax|38789-4|LNC|Shoulder right X-ray Grashey axillary Y|Shoulder right X-ray Grashey axillary Y
C0801762|T102|relax|37157-5|LNC|Shoulder left X-ray Grashey outlet|Shoulder left X-ray Grashey outlet
C0801762|T102|relax|38791-0|LNC|Shoulder right X-ray Grashey outlet|Shoulder right X-ray Grashey outlet
C0801762|T102|relax|39350-4|LNC|Shoulder bilateral X-ray Grashey outlet Serendipity|Shoulder bilateral X-ray Grashey outlet Serendipity
C0801762|T102|relax|37162-5|LNC|Shoulder left X-ray Grashey outlet Serendipity|Shoulder left X-ray Grashey outlet Serendipity
C0801762|T102|relax|38794-4|LNC|Shoulder right X-ray Grashey outlet Serendipity|Shoulder right X-ray Grashey outlet Serendipity
C0801762|T102|relax|37167-4|LNC|Shoulder left X-ray Grashey West Point|Shoulder left X-ray Grashey West Point
C0801762|T102|relax|38795-1|LNC|Shoulder right X-ray Grashey West Point|Shoulder right X-ray Grashey West Point
C0801762|T102|relax|69156-8|LNC|Shoulder left X-ray Grashey Y|Shoulder left X-ray Grashey Y
C0801762|T102|relax|43790-5|LNC|Shoulder right X-ray Grashey Y|Shoulder right X-ray Grashey Y
C0801762|T102|relax|38004-8|LNC|Shoulder left X-ray Grashey W WO weight|Shoulder left X-ray Grashey W WO weight
C0801762|T102|relax|38816-5|LNC|Shoulder right X-ray Grashey W WO weight|Shoulder right X-ray Grashey W WO weight
C0801762|T102|relax|37539-4|LNC|Breast Mammogram grid|Breast Mammogram grid
C0801762|T102|relax|37540-2|LNC|Knee bilateral X-ray Holmblad standing|Knee bilateral X-ray Holmblad standing
C0801762|T102|relax|30771-0|LNC|Pelvis X-ray inlet outlet|Pelvis X-ray inlet outlet
C0801762|T102|relax|37627-7|LNC|Pelvis X-ray inlet outlet oblique|Pelvis X-ray inlet outlet oblique
C0801762|T102|relax|37164-1|LNC|Facial bones X-ray lateral Caldwell Waters|Facial bones X-ray lateral Caldwell Waters
C0801762|T102|relax|37864-6|LNC|Sinuses X-ray lateral Caldwell Waters|Sinuses X-ray lateral Caldwell Waters
C0801762|T102|relax|37165-8|LNC|Facial bones X-ray lateral Caldwell Waters submentovertex|Facial bones X-ray lateral Caldwell Waters submentovertex
C0801762|T102|relax|37166-6|LNC|Facial bones X-ray lateral Caldwell Waters submentovertex Towne|Facial bones X-ray lateral Caldwell Waters submentovertex Towne
C0801762|T102|relax|37871-1|LNC|Skull X-ray lateral Caldwell Waters Towne|Skull X-ray lateral Caldwell Waters Towne
C0801762|T102|relax|37134-4|LNC|Ankle bilateral X-ray lateral Mortise|Ankle bilateral X-ray lateral Mortise
C0801762|T102|relax|37135-1|LNC|Ankle left X-ray lateral Mortise|Ankle left X-ray lateral Mortise
C0801762|T102|relax|37670-7|LNC|Ankle right X-ray lateral Mortise|Ankle right X-ray lateral Mortise
C0801762|T102|relax|42382-2|LNC|Ankle left X-ray lateral Mortise Broden W manual stress|Ankle left X-ray lateral Mortise Broden W manual stress
C0801762|T102|relax|39366-0|LNC|Scapula X-ray lateral outlet|Scapula X-ray lateral outlet
C0801762|T102|relax|43464-7|LNC|Ribs bilateral Chest X-ray lateral PA chest|Ribs bilateral Chest X-ray lateral PA chest
C0801762|T102|relax|37603-8|LNC|Ribs left Chest X-ray lateral PA chest|Ribs left Chest X-ray lateral PA chest
C0801762|T102|relax|39100-3|LNC|Ribs right Chest X-ray lateral PA chest|Ribs right Chest X-ray lateral PA chest
C0801762|T102|relax|39101-1|LNC|Ribs Chest X-ray lateral PA chest|Ribs Chest X-ray lateral PA chest
C0801762|T102|relax|39341-3|LNC|Chest X-ray lateral PA W inspiration expiration|Chest X-ray lateral PA W inspiration expiration
C0801762|T102|relax|39406-4|LNC|Sternum X-ray lateral right anterior oblique|Sternum X-ray lateral right anterior oblique
C0801762|T102|relax|39405-6|LNC|Sternum X-ray lateral right oblique left oblique|Sternum X-ray lateral right oblique left oblique
C0801762|T102|relax|42436-6|LNC|Sella turcica X-ray lateral Towne|Sella turcica X-ray lateral Towne
C0801762|T102|relax|37869-5|LNC|Skull X-ray lateral Towne|Skull X-ray lateral Towne
C0801762|T102|relax|37605-3|LNC|Nasal bones X-ray lateral Waters|Nasal bones X-ray lateral Waters
C0801762|T102|relax|37862-0|LNC|Sinuses X-ray lateral Waters|Sinuses X-ray lateral Waters
C0801762|T102|relax|37136-9|LNC|Shoulder left X-ray lateral Y|Shoulder left X-ray lateral Y
C0801762|T102|relax|37803-4|LNC|Shoulder right X-ray lateral Y|Shoulder right X-ray lateral Y
C0801762|T102|relax|39340-5|LNC|Spine Lumbar X-ray lateral standing W flexion W extension|Spine Lumbar X-ray lateral standing W flexion W extension
C0801762|T102|relax|37133-6|LNC|Spine Cervical X-ray lateral W flexion W extension|Spine Cervical X-ray lateral W flexion W extension
C0801762|T102|relax|37132-8|LNC|Spine Lumbar X-ray lateral W flexion W extension|Spine Lumbar X-ray lateral W flexion W extension
C0801762|T102|relax|38010-5|LNC|Spine Thoracic X-ray lateral W flexion W extension|Spine Thoracic X-ray lateral W flexion W extension
C0801762|T102|relax|37929-7|LNC|Wrist X-ray lateral W flexion W extension|Wrist X-ray lateral W flexion W extension
C0801762|T102|relax|69157-6|LNC|Wrist left X-ray lateral W flexion W extension|Wrist left X-ray lateral W flexion W extension
C0801762|T102|relax|39515-2|LNC|Wrist right X-ray lateral W flexion W extension|Wrist right X-ray lateral W flexion W extension
C0801762|T102|relax|37474-4|LNC|Ankle left X-ray lateral W manual stress|Ankle left X-ray lateral W manual stress
C0801762|T102|relax|37669-9|LNC|Ankle right X-ray lateral W manual stress|Ankle right X-ray lateral W manual stress
C0801762|T102|relax|43480-3|LNC|Joint X-ray lateral W manual stress|Joint X-ray lateral W manual stress
C0801762|T102|relax|37541-0|LNC|Mastoid bilateral X-ray law Mayer Stenver Towne|Mastoid bilateral X-ray law Mayer Stenver Towne
C0801762|T102|relax|47380-1|LNC|Mandible X-ray LE 3 views|Mandible X-ray LE 3 views
C0801762|T102|relax|43470-4|LNC|Skull X-ray LE 3 views|Skull X-ray LE 3 views
C0801762|T102|relax|47377-7|LNC|Knee right X-ray LE 4 views|Knee right X-ray LE 4 views
C0801762|T102|relax|24610-8|LNC|Breast Mammogram limited|Breast Mammogram limited
C0801762|T102|relax|26287-3|LNC|Breast bilateral Mammogram limited|Breast bilateral Mammogram limited
C0801762|T102|relax|26289-9|LNC|Breast left Mammogram limited|Breast left Mammogram limited
C0801762|T102|relax|26291-5|LNC|Breast right Mammogram limited|Breast right Mammogram limited
C0801762|T102|relax|41826-9|LNC|Elbow left X-ray limited|Elbow left X-ray limited
C0801762|T102|relax|41785-7|LNC|Elbow right X-ray limited|Elbow right X-ray limited
C0801762|T102|relax|36737-5|LNC|Facial bones X-ray limited|Facial bones X-ray limited
C0801762|T102|relax|41830-1|LNC|Hand left X-ray limited|Hand left X-ray limited
C0801762|T102|relax|41789-9|LNC|Hand right X-ray limited|Hand right X-ray limited
C0801762|T102|relax|36738-3|LNC|Mandible X-ray limited|Mandible X-ray limited
C0801762|T102|relax|36893-6|LNC|Mastoid X-ray limited|Mastoid X-ray limited
C0801762|T102|relax|42007-5|LNC|Mastoid bilateral X-ray limited|Mastoid bilateral X-ray limited
C0801762|T102|relax|37646-7|LNC|Sacroiliac Joint X-ray limited|Sacroiliac Joint X-ray limited
C0801762|T102|relax|44209-5|LNC|Sinuses X-ray limited|Sinuses X-ray limited
C0801762|T102|relax|48466-7|LNC|Skull X-ray limited|Skull X-ray limited
C0801762|T102|relax|42710-4|LNC|Spine Cervical X-ray limited|Spine Cervical X-ray limited
C0801762|T102|relax|36739-1|LNC|Wrist bilateral X-ray limited|Wrist bilateral X-ray limited
C0801762|T102|relax|38838-9|LNC|Wrist left X-ray limited|Wrist left X-ray limited
C0801762|T102|relax|37642-6|LNC|Wrist right X-ray limited|Wrist right X-ray limited
C0801762|T102|relax|41797-2|LNC|Colon Fluoroscopy limited W air barium contrast PR|Colon Fluoroscopy limited W air barium contrast PR
C0801762|T102|relax|42335-0|LNC|Spine Cervical Fluoroscopy limited W contrast IT|Spine Cervical Fluoroscopy limited W contrast IT
C0801762|T102|relax|38125-1|LNC|Spine Cervical Thoracic Lumbar Fluoroscopy limited W contrast IT|Spine Cervical Thoracic Lumbar Fluoroscopy limited W contrast IT
C0801762|T102|relax|38120-2|LNC|Spine Thoracic Fluoroscopy limited W contrast IT|Spine Thoracic Fluoroscopy limited W contrast IT
C0801762|T102|relax|37137-7|LNC|Kidney X-ray limited W contrast IV|Kidney X-ray limited W contrast IV
C0801762|T102|relax|39687-9|LNC|Scan limited W GA-67 IV|Scan limited W GA-67 IV
C0801762|T102|relax|39754-7|LNC|Thyroid Scan limited W I-131 IV|Thyroid Scan limited W I-131 IV
C0801762|T102|relax|49571-3|LNC|Scan limited W I-131 MIBG IV|Scan limited W I-131 MIBG IV
C0801762|T102|relax|39843-8|LNC|Scan limited W In-111 Satumomab IV|Scan limited W In-111 Satumomab IV
C0801762|T102|relax|41836-8|LNC|Bone Scan limited W In-111 tagged WBC IV|Bone Scan limited W In-111 tagged WBC IV
C0801762|T102|relax|39627-5|LNC|Bone Scan limited|Bone Scan limited
C0801762|T102|relax|39822-2|LNC|Bone marrow Scan limited|Bone marrow Scan limited
C0801762|T102|relax|39645-7|LNC|Breast Scan limited|Breast Scan limited
C0801762|T102|relax|39695-2|LNC|Lung Scan limited|Lung Scan limited
C0801762|T102|relax|39936-0|LNC|Joint Scan limited|Joint Scan limited
C0801762|T102|relax|37542-8|LNC|Breast Mammogram magnification|Breast Mammogram magnification
C0801762|T102|relax|37543-6|LNC|Breast bilateral Mammogram magnification|Breast bilateral Mammogram magnification
C0801762|T102|relax|37554-3|LNC|Breast bilateral Mammogram magnification spot|Breast bilateral Mammogram magnification spot
C0801762|T102|relax|38854-6|LNC|Breast left Mammogram magnification spot|Breast left Mammogram magnification spot
C0801762|T102|relax|37769-7|LNC|Breast right Mammogram magnification spot|Breast right Mammogram magnification spot
C0801762|T102|relax|30769-4|LNC|Pelvis Hip bilateral X-ray max abduction|Pelvis Hip bilateral X-ray max abduction
C0801762|T102|relax|38086-5|LNC|Knee X-ray Merchants 30 45 60 degrees|Knee X-ray Merchants 30 45 60 degrees
C0801762|T102|relax|39935-2|LNC|Scan multiple areas W GA-67 IV|Scan multiple areas W GA-67 IV
C0801762|T102|relax|39949-3|LNC|Scan multiple areas W In-111 Satumomab IV|Scan multiple areas W In-111 Satumomab IV
C0801762|T102|relax|39904-8|LNC|Bone Scan multiple areas|Bone Scan multiple areas
C0801762|T102|relax|39907-1|LNC|Bone marrow Scan multiple areas|Bone marrow Scan multiple areas
C0801762|T102|relax|39937-8|LNC|Joint Scan multiple areas|Joint Scan multiple areas
C0801762|T102|relax|39950-1|LNC|Prostate Scan multiple areas W Tc-99m capromab pendatide IV|Prostate Scan multiple areas W Tc-99m capromab pendatide IV
C0801762|T102|relax|36608-8|LNC|Elbow X-ray oblique|Elbow X-ray oblique
C0801762|T102|relax|36740-9|LNC|Elbow bilateral X-ray oblique|Elbow bilateral X-ray oblique
C0801762|T102|relax|36741-7|LNC|Elbow left X-ray oblique|Elbow left X-ray oblique
C0801762|T102|relax|37687-1|LNC|Elbow right X-ray oblique|Elbow right X-ray oblique
C0801762|T102|relax|36744-1|LNC|Humerus left X-ray oblique|Humerus left X-ray oblique
C0801762|T102|relax|37737-4|LNC|Humerus right X-ray oblique|Humerus right X-ray oblique
C0801762|T102|relax|36619-5|LNC|Knee X-ray oblique|Knee X-ray oblique
C0801762|T102|relax|36745-8|LNC|Knee bilateral X-ray oblique|Knee bilateral X-ray oblique
C0801762|T102|relax|36746-6|LNC|Knee left X-ray oblique|Knee left X-ray oblique
C0801762|T102|relax|37757-2|LNC|Knee right X-ray oblique|Knee right X-ray oblique
C0801762|T102|relax|36747-4|LNC|Mandible X-ray oblique|Mandible X-ray oblique
C0801762|T102|relax|37630-1|LNC|Pelvis X-ray oblique|Pelvis X-ray oblique
C0801762|T102|relax|36742-5|LNC|Radius bilateral Ulna bilateral X-ray oblique|Radius bilateral Ulna bilateral X-ray oblique
C0801762|T102|relax|36743-3|LNC|Radius left Ulna left X-ray oblique|Radius left Ulna left X-ray oblique
C0801762|T102|relax|37709-3|LNC|Radius right Ulna right X-ray oblique|Radius right Ulna right X-ray oblique
C0801762|T102|relax|36748-2|LNC|Spine Cervical X-ray oblique|Spine Cervical X-ray oblique
C0801762|T102|relax|43791-3|LNC|Spine Lumbar X-ray oblique|Spine Lumbar X-ray oblique
C0801762|T102|relax|48749-6|LNC|Spine Thoracic X-ray oblique|Spine Thoracic X-ray oblique
C0801762|T102|relax|36749-0|LNC|Tibia left Fibula left X-ray oblique|Tibia left Fibula left X-ray oblique
C0801762|T102|relax|37817-4|LNC|Tibia right Fibula right X-ray oblique|Tibia right Fibula right X-ray oblique
C0801762|T102|relax|36894-4|LNC|Tibia Fibula X-ray oblique|Tibia Fibula X-ray oblique
C0801762|T102|relax|37544-4|LNC|Wrist bilateral X-ray oblique|Wrist bilateral X-ray oblique
C0801762|T102|relax|38839-7|LNC|Wrist left X-ray oblique|Wrist left X-ray oblique
C0801762|T102|relax|37643-4|LNC|Wrist right X-ray oblique|Wrist right X-ray oblique
C0801762|T102|relax|42398-8|LNC|Foot X-ray oblique (AP lateral) standing|Foot X-ray oblique (AP lateral) standing
C0801762|T102|relax|37139-3|LNC|Spine Cervical X-ray oblique lateral W flexion W extension|Spine Cervical X-ray oblique lateral W flexion W extension
C0801762|T102|relax|37154-2|LNC|Knee X-ray oblique Sunrise|Knee X-ray oblique Sunrise
C0801762|T102|relax|37155-9|LNC|Knee X-ray oblique Sunrise tunnel|Knee X-ray oblique Sunrise tunnel
C0801762|T102|relax|43469-6|LNC|Unspecified body region X-ray foreign body|Unspecified body region X-ray foreign body
C0801762|T102|relax|37063-5|LNC|Unspecified body region Fluoroscopy foreign body|Unspecified body region Fluoroscopy foreign body
C0801762|T102|relax|37546-9|LNC|Temporomandibular joint bilateral X-ray open closed mouth|Temporomandibular joint bilateral X-ray open closed mouth
C0801762|T102|relax|48491-5|LNC|Temporomandibular joint left X-ray open closed mouth|Temporomandibular joint left X-ray open closed mouth
C0801762|T102|relax|48490-7|LNC|Temporomandibular joint right X-ray open closed mouth|Temporomandibular joint right X-ray open closed mouth
C0801762|T102|relax|48699-3|LNC|Temporomandibular Joint unilateral X-ray open closed mouth|Temporomandibular Joint unilateral X-ray open closed mouth
C0801762|T102|relax|37152-6|LNC|Shoulder bilateral X-ray outlet Y|Shoulder bilateral X-ray outlet Y
C0801762|T102|relax|37140-1|LNC|Shoulder left X-ray outlet Y|Shoulder left X-ray outlet Y
C0801762|T102|relax|37804-2|LNC|Shoulder right X-ray outlet Y|Shoulder right X-ray outlet Y
C0801762|T102|relax|36750-8|LNC|Chest X-ray PA AP lateral-decubitus|Chest X-ray PA AP lateral-decubitus
C0801762|T102|relax|42272-5|LNC|Chest X-ray PA lateral|Chest X-ray PA lateral
C0801762|T102|relax|36751-6|LNC|Chest Fluoroscopy PA lateral|Chest Fluoroscopy PA lateral
C0801762|T102|relax|36752-4|LNC|Hand bilateral X-ray PA lateral|Hand bilateral X-ray PA lateral
C0801762|T102|relax|36753-2|LNC|Hand left X-ray PA lateral|Hand left X-ray PA lateral
C0801762|T102|relax|37713-5|LNC|Hand right X-ray PA lateral|Hand right X-ray PA lateral
C0801762|T102|relax|36754-0|LNC|Mandible X-ray PA lateral|Mandible X-ray PA lateral
C0801762|T102|relax|30721-5|LNC|Sinuses X-ray PA lateral|Sinuses X-ray PA lateral
C0801762|T102|relax|37547-7|LNC|Wrist bilateral X-ray PA lateral|Wrist bilateral X-ray PA lateral
C0801762|T102|relax|37548-5|LNC|Wrist left X-ray PA lateral|Wrist left X-ray PA lateral
C0801762|T102|relax|37835-6|LNC|Wrist right X-ray PA lateral|Wrist right X-ray PA lateral
C0801762|T102|relax|37143-5|LNC|Chest X-ray PA lateral AP lateral-decubitus|Chest X-ray PA lateral AP lateral-decubitus
C0801762|T102|relax|37144-3|LNC|Chest X-ray PA lateral AP left lateral-decubitus|Chest X-ray PA lateral AP left lateral-decubitus
C0801762|T102|relax|37145-0|LNC|Chest X-ray PA lateral AP right lateral-decubitus|Chest X-ray PA lateral AP right lateral-decubitus
C0801762|T102|relax|37142-7|LNC|Hand bilateral X-ray PA lateral Ball Catcher|Hand bilateral X-ray PA lateral Ball Catcher
C0801762|T102|relax|37860-4|LNC|Sinuses X-ray PA lateral Caldwell Waters|Sinuses X-ray PA lateral Caldwell Waters
C0801762|T102|relax|37146-8|LNC|Chest X-ray PA lateral left oblique|Chest X-ray PA lateral left oblique
C0801762|T102|relax|30741-3|LNC|Chest X-ray PA lateral lordotic upright|Chest X-ray PA lateral lordotic upright
C0801762|T102|relax|39078-1|LNC|Finger X-ray PA lateral oblique|Finger X-ray PA lateral oblique
C0801762|T102|relax|36755-7|LNC|Hand X-ray PA lateral oblique|Hand X-ray PA lateral oblique
C0801762|T102|relax|36756-5|LNC|Hand bilateral X-ray PA lateral oblique|Hand bilateral X-ray PA lateral oblique
C0801762|T102|relax|36757-3|LNC|Hand left X-ray PA lateral oblique|Hand left X-ray PA lateral oblique
C0801762|T102|relax|37715-0|LNC|Hand right X-ray PA lateral oblique|Hand right X-ray PA lateral oblique
C0801762|T102|relax|37884-4|LNC|Sternum X-ray PA lateral oblique|Sternum X-ray PA lateral oblique
C0801762|T102|relax|37549-3|LNC|Wrist bilateral X-ray PA lateral oblique|Wrist bilateral X-ray PA lateral oblique
C0801762|T102|relax|37550-1|LNC|Wrist left X-ray PA lateral oblique|Wrist left X-ray PA lateral oblique
C0801762|T102|relax|37836-4|LNC|Wrist right X-ray PA lateral oblique|Wrist right X-ray PA lateral oblique
C0801762|T102|relax|36758-1|LNC|Chest X-ray PA lateral oblique lordotic|Chest X-ray PA lateral oblique lordotic
C0801762|T102|relax|37148-4|LNC|Mandible X-ray PA lateral oblique Towne|Mandible X-ray PA lateral oblique Towne
C0801762|T102|relax|37147-6|LNC|Chest X-ray PA lateral right oblique|Chest X-ray PA lateral right oblique
C0801762|T102|relax|30742-1|LNC|Chest X-ray PA lateral right oblique left oblique|Chest X-ray PA lateral right oblique left oblique
C0801762|T102|relax|30743-9|LNC|Chest X-ray PA lateral right oblique left oblique portable|Chest X-ray PA lateral right oblique left oblique portable
C0801762|T102|relax|30744-7|LNC|Chest X-ray PA lateral right or-left oblique|Chest X-ray PA lateral right or-left oblique
C0801762|T102|relax|24643-9|LNC|Chest X-ray PA lateral right or-left oblique upright|Chest X-ray PA lateral right or-left oblique upright
C0801762|T102|relax|37149-2|LNC|Patella left X-ray PA lateral Sunrise|Patella left X-ray PA lateral Sunrise
C0801762|T102|relax|38790-2|LNC|Patella right X-ray PA lateral Sunrise|Patella right X-ray PA lateral Sunrise
C0801762|T102|relax|37859-6|LNC|Sinuses X-ray PA lateral Waters|Sinuses X-ray PA lateral Waters
C0801762|T102|relax|69271-5|LNC|Skull X-ray PA lateral Waters Towne|Skull X-ray PA lateral Waters Towne
C0801762|T102|relax|24647-0|LNC|Chest X-ray PA lateral upright|Chest X-ray PA lateral upright
C0801762|T102|relax|24644-7|LNC|Chest X-ray PA lateral upright portable|Chest X-ray PA lateral upright portable
C0801762|T102|relax|36759-9|LNC|Chest X-ray PA lordotic|Chest X-ray PA lordotic
C0801762|T102|relax|39079-9|LNC|Hand X-ray PA oblique|Hand X-ray PA oblique
C0801762|T102|relax|37141-9|LNC|Chest X-ray PA right lateral|Chest X-ray PA right lateral
C0801762|T102|relax|39519-4|LNC|Skull X-ray PA right lateral left lateral|Skull X-ray PA right lateral left lateral
C0801762|T102|relax|39521-0|LNC|Skull X-ray PA right lateral left lateral Caldwell Towne|Skull X-ray PA right lateral left lateral Caldwell Towne
C0801762|T102|relax|39520-2|LNC|Skull X-ray PA right lateral left lateral Towne|Skull X-ray PA right lateral left lateral Towne
C0801762|T102|relax|24646-2|LNC|Chest X-ray PA right lateral right oblique left oblique upright|Chest X-ray PA right lateral right oblique left oblique upright
C0801762|T102|relax|24645-4|LNC|Chest X-ray PA right lateral right oblique left oblique upright portable|Chest X-ray PA right lateral right oblique left oblique upright portable
C0801762|T102|relax|37150-0|LNC|Chest X-ray PA right oblique left oblique|Chest X-ray PA right oblique left oblique
C0801762|T102|relax|24635-5|LNC|Chest X-ray PA upright W inspiration expiration|Chest X-ray PA upright W inspiration expiration
C0801762|T102|relax|46378-6|LNC|Knee bilateral X-ray PA standing W flexion|Knee bilateral X-ray PA standing W flexion
C0801762|T102|relax|43660-0|LNC|Heart Scan perfusion qualitative at rest W radionuclide IV|Heart Scan perfusion qualitative at rest W radionuclide IV
C0801762|T102|relax|43661-8|LNC|Heart Scan perfusion quantitative at rest W radionuclide IV|Heart Scan perfusion quantitative at rest W radionuclide IV
C0801762|T102|relax|43658-4|LNC|Heart Scan perfusion quantitative|Heart Scan perfusion quantitative
C0801762|T102|relax|43656-8|LNC|Lung Scan perfusion quantitative|Lung Scan perfusion quantitative
C0801762|T102|relax|39719-0|LNC|Heart Scan perfusion at rest W adenosine W radionuclide IV|Heart Scan perfusion at rest W adenosine W radionuclide IV
C0801762|T102|relax|43777-2|LNC|Heart Scan perfusion at rest W adenosine W Tl-201 IV|Heart Scan perfusion at rest W adenosine W Tl-201 IV
C0801762|T102|relax|39722-4|LNC|Heart Scan perfusion at rest W dipyridamole W radionuclide IV|Heart Scan perfusion at rest W dipyridamole W radionuclide IV
C0801762|T102|relax|39720-8|LNC|Heart Scan perfusion at rest W dipyridamole W Tc-99m Sestamibi IV|Heart Scan perfusion at rest W dipyridamole W Tc-99m Sestamibi IV
C0801762|T102|relax|39728-1|LNC|Heart Scan perfusion at rest W radionuclide IV|Heart Scan perfusion at rest W radionuclide IV
C0801762|T102|relax|39726-5|LNC|Heart Scan perfusion at rest W stress W radionuclide IV|Heart Scan perfusion at rest W stress W radionuclide IV
C0801762|T102|relax|39727-3|LNC|Heart Scan perfusion at rest W stress W Tc-99m Sestamibi IV|Heart Scan perfusion at rest W stress W Tc-99m Sestamibi IV
C0801762|T102|relax|39699-4|LNC|Heart Scan perfusion at rest W Tc-99m Sestamibi IV|Heart Scan perfusion at rest W Tc-99m Sestamibi IV
C0801762|T102|relax|39701-8|LNC|Heart Scan perfusion W adenosine W radionuclide IV|Heart Scan perfusion W adenosine W radionuclide IV
C0801762|T102|relax|39731-5|LNC|Heart Scan perfusion W adenosine W Tc-99m Sestamibi IV|Heart Scan perfusion W adenosine W Tc-99m Sestamibi IV
C0801762|T102|relax|39735-6|LNC|Heart Scan perfusion W adenosine W Tl-201 IV|Heart Scan perfusion W adenosine W Tl-201 IV
C0801762|T102|relax|39708-3|LNC|Heart Scan perfusion W dipyridamole W radionuclide IV|Heart Scan perfusion W dipyridamole W radionuclide IV
C0801762|T102|relax|39709-1|LNC|Heart Scan perfusion W dipyridamole W Tc-99m IV|Heart Scan perfusion W dipyridamole W Tc-99m IV
C0801762|T102|relax|39705-9|LNC|Heart Scan perfusion W dipyridamole W Tc-99m Sestamibi IV|Heart Scan perfusion W dipyridamole W Tc-99m Sestamibi IV
C0801762|T102|relax|39707-5|LNC|Heart Scan perfusion W dipyridamole W Tl-201 IV|Heart Scan perfusion W dipyridamole W Tl-201 IV
C0801762|T102|relax|39703-4|LNC|Heart Scan perfusion W dobutamine W radionuclide IV|Heart Scan perfusion W dobutamine W radionuclide IV
C0801762|T102|relax|39702-6|LNC|Heart Scan perfusion W dobutamine W Tc-99m Sestamibi IV|Heart Scan perfusion W dobutamine W Tc-99m Sestamibi IV
C0801762|T102|relax|39733-1|LNC|Heart Scan perfusion W dobutamine W Tl-201 IV|Heart Scan perfusion W dobutamine W Tl-201 IV
C0801762|T102|relax|39941-0|LNC|Lung Scan perfusion W particulate radionuclide IV|Lung Scan perfusion W particulate radionuclide IV
C0801762|T102|relax|39833-9|LNC|Lung Scan perfusion W radionuclide gaseous inhaled|Lung Scan perfusion W radionuclide gaseous inhaled
C0801762|T102|relax|39716-6|LNC|Heart Scan perfusion|Heart Scan perfusion
C0801762|T102|relax|39697-8|LNC|Lung Scan perfusion|Lung Scan perfusion
C0801762|T102|relax|39730-7|LNC|Heart Scan perfusion W stress W radionuclide IV|Heart Scan perfusion W stress W radionuclide IV
C0801762|T102|relax|39732-3|LNC|Heart Scan perfusion W stress W Tc-99m Sestamibi IV|Heart Scan perfusion W stress W Tc-99m Sestamibi IV
C0801762|T102|relax|39715-8|LNC|Heart Scan perfusion W stress W Tl-201 IV|Heart Scan perfusion W stress W Tl-201 IV
C0801762|T102|relax|39704-2|LNC|Heart Scan perfusion W Tc-99m Sestamibi IV|Heart Scan perfusion W Tc-99m Sestamibi IV
C0801762|T102|relax|39714-1|LNC|Heart Scan perfusion W Tl-201 IV|Heart Scan perfusion W Tl-201 IV
C0801762|T102|relax|39713-3|LNC|Heart Scan perfusion W Tl-201 IV Tc-99m Tetrofosmin IV|Heart Scan perfusion W Tl-201 IV Tc-99m Tetrofosmin IV
C0801762|T102|relax|30765-2|LNC|Acetabulum X-ray portable|Acetabulum X-ray portable
C0801762|T102|relax|30764-5|LNC|Acetabulum bilateral X-ray portable|Acetabulum bilateral X-ray portable
C0801762|T102|relax|41823-6|LNC|Ankle left X-ray portable|Ankle left X-ray portable
C0801762|T102|relax|41782-4|LNC|Ankle right X-ray portable|Ankle right X-ray portable
C0801762|T102|relax|30746-2|LNC|Chest X-ray portable|Chest X-ray portable
C0801762|T102|relax|41827-7|LNC|Elbow left X-ray portable|Elbow left X-ray portable
C0801762|T102|relax|41786-5|LNC|Elbow right X-ray portable|Elbow right X-ray portable
C0801762|T102|relax|41773-3|LNC|Facial bones X-ray portable|Facial bones X-ray portable
C0801762|T102|relax|41818-6|LNC|Femur left X-ray portable|Femur left X-ray portable
C0801762|T102|relax|41778-2|LNC|Femur right X-ray portable|Femur right X-ray portable
C0801762|T102|relax|43570-1|LNC|Hand X-ray portable|Hand X-ray portable
C0801762|T102|relax|41829-3|LNC|Hand left X-ray portable|Hand left X-ray portable
C0801762|T102|relax|41788-1|LNC|Hand right X-ray portable|Hand right X-ray portable
C0801762|T102|relax|37168-2|LNC|Hip X-ray portable|Hip X-ray portable
C0801762|T102|relax|37169-0|LNC|Hip left X-ray portable|Hip left X-ray portable
C0801762|T102|relax|38796-9|LNC|Hip right X-ray portable|Hip right X-ray portable
C0801762|T102|relax|37170-8|LNC|Humerus X-ray portable|Humerus X-ray portable
C0801762|T102|relax|41825-1|LNC|Humerus left X-ray portable|Humerus left X-ray portable
C0801762|T102|relax|41784-0|LNC|Humerus right X-ray portable|Humerus right X-ray portable
C0801762|T102|relax|41820-2|LNC|Knee left X-ray portable|Knee left X-ray portable
C0801762|T102|relax|41779-0|LNC|Knee right X-ray portable|Knee right X-ray portable
C0801762|T102|relax|30792-6|LNC|Patella X-ray portable|Patella X-ray portable
C0801762|T102|relax|30772-8|LNC|Pelvis X-ray portable|Pelvis X-ray portable
C0801762|T102|relax|30747-0|LNC|Ribs X-ray portable|Ribs X-ray portable
C0801762|T102|relax|41831-9|LNC|Ribs left X-ray portable|Ribs left X-ray portable
C0801762|T102|relax|41791-5|LNC|Ribs right X-ray portable|Ribs right X-ray portable
C0801762|T102|relax|46391-9|LNC|Shoulder X-ray portable|Shoulder X-ray portable
C0801762|T102|relax|41824-4|LNC|Shoulder left X-ray portable|Shoulder left X-ray portable
C0801762|T102|relax|41783-2|LNC|Shoulder right X-ray portable|Shoulder right X-ray portable
C0801762|T102|relax|30723-1|LNC|Skull X-ray portable|Skull X-ray portable
C0801762|T102|relax|37171-6|LNC|Spine Cervical X-ray portable|Spine Cervical X-ray portable
C0801762|T102|relax|44203-8|LNC|Spine Cervical Thoracic Lumbar X-ray portable|Spine Cervical Thoracic Lumbar X-ray portable
C0801762|T102|relax|37172-4|LNC|Spine Lumbar X-ray portable|Spine Lumbar X-ray portable
C0801762|T102|relax|41828-5|LNC|Wrist left X-ray portable|Wrist left X-ray portable
C0801762|T102|relax|41787-3|LNC|Wrist right X-ray portable|Wrist right X-ray portable
C0801762|T102|relax|37151-8|LNC|Unspecified body region Fluoroscopy portable|Unspecified body region Fluoroscopy portable
C0801762|T102|relax|30731-4|LNC|Zygomatic arch X-ray portable|Zygomatic arch X-ray portable
C0801762|T102|relax|30730-6|LNC|Zygomatic arch bilateral X-ray portable|Zygomatic arch bilateral X-ray portable
C0801762|T102|relax|24634-8|LNC|Chest X-ray portable W inspiration expiration|Chest X-ray portable W inspiration expiration
C0801762|T102|relax|24824-5|LNC|Lung Scan portable|Lung Scan portable
C0801762|T102|relax|42402-8|LNC|Unspecified body region X-ray post mortem|Unspecified body region X-ray post mortem
C0801762|T102|relax|43657-6|LNC|Lung Scan quantitative|Lung Scan quantitative
C0801762|T102|relax|30733-0|LNC|Chest X-ray right left oblique portable|Chest X-ray right left oblique portable
C0801762|T102|relax|37131-0|LNC|Abdomen X-ray right lateral left lateral|Abdomen X-ray right lateral left lateral
C0801762|T102|relax|37138-5|LNC|Abdomen X-ray right oblique left oblique|Abdomen X-ray right oblique left oblique
C0801762|T102|relax|41792-3|LNC|Chest X-ray right oblique left oblique|Chest X-ray right oblique left oblique
C0801762|T102|relax|24651-2|LNC|Chest X-ray right oblique left oblique upright|Chest X-ray right oblique left oblique upright
C0801762|T102|relax|42414-3|LNC|Chest X-ray right oblique left oblique W nipple markers|Chest X-ray right oblique left oblique W nipple markers
C0801762|T102|relax|37016-3|LNC|Breast bilateral Mammogram roll|Breast bilateral Mammogram roll
C0801762|T102|relax|37017-1|LNC|Breast left Mammogram roll|Breast left Mammogram roll
C0801762|T102|relax|37775-4|LNC|Breast right Mammogram roll|Breast right Mammogram roll
C0801762|T102|relax|30740-5|LNC|Chest X-ray right or-left oblique|Chest X-ray right or-left oblique
C0801762|T102|relax|30739-7|LNC|Chest X-ray right or-left oblique portable|Chest X-ray right or-left oblique portable
C0801762|T102|relax|43479-5|LNC|Aorta abdominal Fluoroscopic angiogram runoff W contrast IA|Aorta abdominal Fluoroscopic angiogram runoff W contrast IA
C0801762|T102|relax|30838-7|LNC|Aorta Femoral artery bilateral Fluoroscopic angiogram runoff W contrast IA|Aorta Femoral artery bilateral Fluoroscopic angiogram runoff W contrast IA
C0801762|T102|relax|37364-7|LNC|Aorta Femoral artery left Fluoroscopic angiogram runoff W contrast IA|Aorta Femoral artery left Fluoroscopic angiogram runoff W contrast IA
C0801762|T102|relax|38799-3|LNC|Aorta Femoral artery right Fluoroscopic angiogram runoff W contrast IA|Aorta Femoral artery right Fluoroscopic angiogram runoff W contrast IA
C0801762|T102|relax|38107-9|LNC|Wrist X-ray scaphoid|Wrist X-ray scaphoid
C0801762|T102|relax|37304-3|LNC|Wrist bilateral X-ray scaphoid|Wrist bilateral X-ray scaphoid
C0801762|T102|relax|37302-7|LNC|Wrist left X-ray scaphoid|Wrist left X-ray scaphoid
C0801762|T102|relax|38115-2|LNC|Wrist right X-ray scaphoid|Wrist right X-ray scaphoid
C0801762|T102|relax|24930-0|LNC|Spine Thoracic Lumbar X-ray scoliosis|Spine Thoracic Lumbar X-ray scoliosis
C0801762|T102|relax|30715-7|LNC|Spine Thoracic Lumbar X-ray scoliosis AP lateral|Spine Thoracic Lumbar X-ray scoliosis AP lateral
C0801762|T102|relax|42424-2|LNC|Spine Thoracic Lumbar X-ray scoliosis AP lateral sitting|Spine Thoracic Lumbar X-ray scoliosis AP lateral sitting
C0801762|T102|relax|39367-8|LNC|Spine Thoracic Lumbar X-ray scoliosis AP lateral standing|Spine Thoracic Lumbar X-ray scoliosis AP lateral standing
C0801762|T102|relax|42472-1|LNC|Spine Thoracic Lumbar X-ray scoliosis AP in traction|Spine Thoracic Lumbar X-ray scoliosis AP in traction
C0801762|T102|relax|42425-9|LNC|Spine Thoracic Lumbar X-ray scoliosis AP standing W right bending W left bending WO bending|Spine Thoracic Lumbar X-ray scoliosis AP standing W right bending W left bending WO bending
C0801762|T102|relax|43569-3|LNC|Spine Thoracic Lumbar X-ray scoliosis AP upright supine|Spine Thoracic Lumbar X-ray scoliosis AP upright supine
C0801762|T102|relax|30716-5|LNC|Spine Thoracic Lumbar X-ray scoliosis lateral|Spine Thoracic Lumbar X-ray scoliosis lateral
C0801762|T102|relax|30717-3|LNC|Spine Thoracic Lumbar X-ray scoliosis standing|Spine Thoracic Lumbar X-ray scoliosis standing
C0801762|T102|relax|24929-2|LNC|Spine Thoracic Lumbar X-ray scoliosis W flexion W extension|Spine Thoracic Lumbar X-ray scoliosis W flexion W extension
C0801762|T102|relax|24606-6|LNC|Breast Mammogram screening|Breast Mammogram screening
C0801762|T102|relax|39153-2|LNC|Breast FFD mammogram screening|Breast FFD mammogram screening
C0801762|T102|relax|69159-2|LNC|Breast implant X-ray screening|Breast implant X-ray screening
C0801762|T102|relax|48492-3|LNC|Breast implant bilateral Mammogram screening|Breast implant bilateral Mammogram screening
C0801762|T102|relax|26175-0|LNC|Breast bilateral Mammogram screening|Breast bilateral Mammogram screening
C0801762|T102|relax|42174-3|LNC|Breast bilateral FFD mammogram screening|Breast bilateral FFD mammogram screening
C0801762|T102|relax|26176-8|LNC|Breast left Mammogram screening|Breast left Mammogram screening
C0801762|T102|relax|46355-4|LNC|Breast left FFD mammogram screening|Breast left FFD mammogram screening
C0801762|T102|relax|26177-6|LNC|Breast right Mammogram screening|Breast right Mammogram screening
C0801762|T102|relax|46354-7|LNC|Breast right FFD mammogram screening|Breast right FFD mammogram screening
C0801762|T102|relax|46356-2|LNC|Breast unilateral Mammogram screening|Breast unilateral Mammogram screening
C0801762|T102|relax|37022-1|LNC|Calcaneus X-ray ski jump|Calcaneus X-ray ski jump
C0801762|T102|relax|37021-3|LNC|Calcaneus bilateral X-ray ski jump|Calcaneus bilateral X-ray ski jump
C0801762|T102|relax|37023-9|LNC|Calcaneus left X-ray ski jump|Calcaneus left X-ray ski jump
C0801762|T102|relax|38778-7|LNC|Calcaneus right X-ray ski jump|Calcaneus right X-ray ski jump
C0801762|T102|relax|37551-9|LNC|Breast Mammogram spot|Breast Mammogram spot
C0801762|T102|relax|37552-7|LNC|Breast bilateral Mammogram spot|Breast bilateral Mammogram spot
C0801762|T102|relax|38807-4|LNC|Breast right Mammogram spot|Breast right Mammogram spot
C0801762|T102|relax|37553-5|LNC|Breast left Mammogram spot compression|Breast left Mammogram spot compression
C0801762|T102|relax|43550-3|LNC|Brain Scan static flow|Brain Scan static flow
C0801762|T102|relax|39952-7|LNC|Scrotum Testicle Scan static flow|Scrotum Testicle Scan static flow
C0801762|T102|relax|39676-2|LNC|Scan static infection W GA-67 IV|Scan static infection W GA-67 IV
C0801762|T102|relax|39894-1|LNC|Heart Scan static shunt detection|Heart Scan static shunt detection
C0801762|T102|relax|39896-6|LNC|Scan static tumor W GA-67 IV|Scan static tumor W GA-67 IV
C0801762|T102|relax|39814-9|LNC|Bone Scan static limited|Bone Scan static limited
C0801762|T102|relax|39634-1|LNC|Brain Scan static limited|Brain Scan static limited
C0801762|T102|relax|39903-0|LNC|Bone Scan static multiple areas|Bone Scan static multiple areas
C0801762|T102|relax|39817-2|LNC|Bone Scan static whole body|Bone Scan static whole body
C0801762|T102|relax|39815-6|LNC|Bone Scan static|Bone Scan static
C0801762|T102|relax|39824-8|LNC|Bone marrow Scan static|Bone marrow Scan static
C0801762|T102|relax|39633-3|LNC|Brain Scan static|Brain Scan static
C0801762|T102|relax|39853-7|LNC|Kidney bilateral Scan static|Kidney bilateral Scan static
C0801762|T102|relax|39832-1|LNC|Liver Scan static|Liver Scan static
C0801762|T102|relax|39878-4|LNC|Liver Spleen Scan static|Liver Spleen Scan static
C0801762|T102|relax|39900-6|LNC|Salivary gland Scan static|Salivary gland Scan static
C0801762|T102|relax|39855-2|LNC|Scrotum Testicle Scan static|Scrotum Testicle Scan static
C0801762|T102|relax|43501-6|LNC|Vessel Scan static|Vessel Scan static
C0801762|T102|relax|44150-1|LNC|Brain Scan static W Tc-99m bicisate IV|Brain Scan static W Tc-99m bicisate IV
C0801762|T102|relax|39854-5|LNC|Kidney bilateral Scan static W Tc-99m DMSA IV|Kidney bilateral Scan static W Tc-99m DMSA IV
C0801762|T102|relax|37153-4|LNC|Mastoid X-ray Stenver Arcelin|Mastoid X-ray Stenver Arcelin
C0801762|T102|relax|69136-0|LNC|Knee X-ray Sunrise tunnel|Knee X-ray Sunrise tunnel
C0801762|T102|relax|37163-3|LNC|Knee bilateral X-ray Sunrise tunnel|Knee bilateral X-ray Sunrise tunnel
C0801762|T102|relax|37156-7|LNC|Knee left X-ray Sunrise tunnel|Knee left X-ray Sunrise tunnel
C0801762|T102|relax|37759-8|LNC|Knee right X-ray Sunrise tunnel|Knee right X-ray Sunrise tunnel
C0801762|T102|relax|39345-4|LNC|Knee left X-ray Sunrise tunnel standing|Knee left X-ray Sunrise tunnel standing
C0801762|T102|relax|69255-8|LNC|Knee right X-ray Sunrise tunnel standing|Knee right X-ray Sunrise tunnel standing
C0801762|T102|relax|38088-1|LNC|Knee bilateral X-ray Sunrise 20 40 60 degrees|Knee bilateral X-ray Sunrise 20 40 60 degrees
C0801762|T102|relax|38087-3|LNC|Knee left X-ray Sunrise 20 40 60 degrees|Knee left X-ray Sunrise 20 40 60 degrees
C0801762|T102|relax|38824-9|LNC|Knee right X-ray Sunrise 20 40 60 degrees|Knee right X-ray Sunrise 20 40 60 degrees
C0801762|T102|relax|24579-5|LNC|Bones long X-ray survey|Bones long X-ray survey
C0801762|T102|relax|43518-0|LNC|Bones X-ray survey|Bones X-ray survey
C0801762|T102|relax|37365-4|LNC|Bones X-ray survey metastasis|Bones X-ray survey metastasis
C0801762|T102|relax|39518-6|LNC|Bones long X-ray survey limited|Bones long X-ray survey limited
C0801762|T102|relax|43519-8|LNC|Bones X-ray survey limited|Bones X-ray survey limited
C0801762|T102|relax|38089-9|LNC|Bones X-ray survey limited metastasis|Bones X-ray survey limited metastasis
C0801762|T102|relax|37159-1|LNC|Foot left X-ray tarsal|Foot left X-ray tarsal
C0801762|T102|relax|38792-8|LNC|Foot right X-ray tarsal|Foot right X-ray tarsal
C0801762|T102|relax|43796-2|LNC|Wrist bilateral X-ray tunnel carpal|Wrist bilateral X-ray tunnel carpal
C0801762|T102|relax|69304-4|LNC|Wrist X-ray ulnar deviation|Wrist X-ray ulnar deviation
C0801762|T102|relax|69303-6|LNC|Wrist X-ray ulnar deviation radial deviation|Wrist X-ray ulnar deviation radial deviation
C0801762|T102|relax|69072-7|LNC|Wrist bilateral X-ray ulnar deviation radial deviation|Wrist bilateral X-ray ulnar deviation radial deviation
C0801762|T102|relax|37555-0|LNC|Wrist left X-ray ulnar deviation radial deviation|Wrist left X-ray ulnar deviation radial deviation
C0801762|T102|relax|38808-2|LNC|Wrist right X-ray ulnar deviation radial deviation|Wrist right X-ray ulnar deviation radial deviation
C0801762|T102|relax|43532-1|LNC|Chest Abdomen X-ray upright PA chest|Chest Abdomen X-ray upright PA chest
C0801762|T102|relax|39944-4|LNC|Lung Scan ventilation equilibrium washout W radionuclide inhaled|Lung Scan ventilation equilibrium washout W radionuclide inhaled
C0801762|T102|relax|39948-5|LNC|Lung Scan ventilation equilibrium washout W radionuclide inhaled single breath|Lung Scan ventilation equilibrium washout W radionuclide inhaled single breath
C0801762|T102|relax|39947-7|LNC|Lung Scan ventilation equilibrium W radionuclide inhaled single breath|Lung Scan ventilation equilibrium W radionuclide inhaled single breath
C0801762|T102|relax|39946-9|LNC|Lung Scan ventilation perfusion differential W radionuclide inhaled W radionuclide IV|Lung Scan ventilation perfusion differential W radionuclide inhaled W radionuclide IV
C0801762|T102|relax|39943-6|LNC|Lung Scan ventilation perfusion W radionuclide inhaled W particulate radionuclide IV|Lung Scan ventilation perfusion W radionuclide inhaled W particulate radionuclide IV
C0801762|T102|relax|30697-7|LNC|Pulmonary system Scan ventilation perfusion W radionuclide inhaled W radionuclide IV|Pulmonary system Scan ventilation perfusion W radionuclide inhaled W radionuclide IV
C0801762|T102|relax|39942-8|LNC|Lung Scan ventilation perfusion W radionuclide inhaled single breath W particulate radionuclide IV|Lung Scan ventilation perfusion W radionuclide inhaled single breath W particulate radionuclide IV
C0801762|T102|relax|24888-0|LNC|Pulmonary system Scan ventilation perfusion W Xe-133 inhaled W Tc-99m MAA IV|Pulmonary system Scan ventilation perfusion W Xe-133 inhaled W Tc-99m MAA IV
C0801762|T102|relax|39835-4|LNC|Lung Scan ventilation W radionuclide aerosol inhaled|Lung Scan ventilation W radionuclide aerosol inhaled
C0801762|T102|relax|39836-2|LNC|Lung Scan ventilation W radionuclide gaseous inhaled|Lung Scan ventilation W radionuclide gaseous inhaled
C0801762|T102|relax|39945-1|LNC|Lung Scan ventilation W radionuclide gaseous inhaled single breath|Lung Scan ventilation W radionuclide gaseous inhaled single breath
C0801762|T102|relax|39837-0|LNC|Lung Scan ventilation W radionuclide inhaled|Lung Scan ventilation W radionuclide inhaled
C0801762|T102|relax|39834-7|LNC|Lung Scan ventilation W Tc-99m DTPA aerosol inhaled|Lung Scan ventilation W Tc-99m DTPA aerosol inhaled
C0801762|T102|relax|46361-2|LNC|Lung Scan ventilation W Xe-133 inhaled|Lung Scan ventilation W Xe-133 inhaled
C0801762|T102|relax|39932-9|LNC|Heart Scan wall motion ejection fraction|Heart Scan wall motion ejection fraction
C0801762|T102|relax|39873-5|LNC|Heart Scan wall motion|Heart Scan wall motion
C0801762|T102|relax|39683-8|LNC|Scan whole body W GA-67 IV|Scan whole body W GA-67 IV
C0801762|T102|relax|39698-6|LNC|Scan whole body W I-131 MIBG IV|Scan whole body W I-131 MIBG IV
C0801762|T102|relax|39845-3|LNC|Scan whole body W In-111 Satumomab IV|Scan whole body W In-111 Satumomab IV
C0801762|T102|relax|42711-2|LNC|Scan whole body W In-111 tagged WBC IV|Scan whole body W In-111 tagged WBC IV
C0801762|T102|relax|42175-0|LNC|Scan whole body|Scan whole body
C0801762|T102|relax|39818-0|LNC|Bone Scan whole body|Bone Scan whole body
C0801762|T102|relax|39826-3|LNC|Bone marrow Scan whole body|Bone marrow Scan whole body
C0801762|T102|relax|39669-7|LNC|Scan whole body W Tc-99m Arcitumomab IV|Scan whole body W Tc-99m Arcitumomab IV
C0801762|T102|relax|24713-0|LNC|Gallbladder X-ray 48 hours post contrast PO|Gallbladder X-ray 48 hours post contrast PO
C0801762|T102|relax|39660-6|LNC|Heart Scan at rest W dipyridamole W radionuclide IV|Heart Scan at rest W dipyridamole W radionuclide IV
C0801762|T102|relax|39661-4|LNC|Heart Scan at rest W dobutamine W radionuclide IV|Heart Scan at rest W dobutamine W radionuclide IV
C0801762|T102|relax|39663-0|LNC|Heart Scan at rest W stress W radionuclide IV|Heart Scan at rest W stress W radionuclide IV
C0801762|T102|relax|42309-5|LNC|Heart Scan at rest W stress W Tl-201 IV|Heart Scan at rest W stress W Tl-201 IV
C0801762|T102|relax|24750-2|LNC|Heart Scan at rest W Tl-201 IV|Heart Scan at rest W Tl-201 IV
C0801762|T102|relax|43459-7|LNC|Brain Scan during electroconvulsive shock treatment|Brain Scan during electroconvulsive shock treatment
C0801762|T102|relax|24577-9|LNC|Bone X-ray during surgery|Bone X-ray during surgery
C0801762|T102|relax|47372-8|LNC|Hip X-ray during surgery|Hip X-ray during surgery
C0801762|T102|relax|25070-4|LNC|Unspecified body region Fluoroscopy during surgery|Unspecified body region Fluoroscopy during surgery
C0801762|T102|relax|24574-6|LNC|Biliary ducts Gallbladder Fluoroscopy during surgery W contrast biliary duct|Biliary ducts Gallbladder Fluoroscopy during surgery W contrast biliary duct
C0801762|T102|relax|46352-1|LNC|Breast duct Mammogram during surgery W contrast intra duct|Breast duct Mammogram during surgery W contrast intra duct
C0801762|T102|relax|43485-2|LNC|Kidney X-ray during surgery W contrast retrograde|Kidney X-ray during surgery W contrast retrograde
C0801762|T102|relax|39150-8|LNC|Breast FFD mammogram Post Localization|Breast FFD mammogram Post Localization
C0801762|T102|relax|69251-7|LNC|Breast Mammogram Post Wire Placement|Breast Mammogram Post Wire Placement
C0801762|T102|relax|42415-0|LNC|Breast bilateral Mammogram Post Wire Placement|Breast bilateral Mammogram Post Wire Placement
C0801762|T102|relax|42416-8|LNC|Breast left Mammogram Post Wire Placement|Breast left Mammogram Post Wire Placement
C0801762|T102|relax|37201-1|LNC|Ankle X-ray standing|Ankle X-ray standing
C0801762|T102|relax|37202-9|LNC|Ankle bilateral X-ray standing|Ankle bilateral X-ray standing
C0801762|T102|relax|37203-7|LNC|Ankle left X-ray standing|Ankle left X-ray standing
C0801762|T102|relax|37676-4|LNC|Ankle right X-ray standing|Ankle right X-ray standing
C0801762|T102|relax|37205-2|LNC|Calcaneus X-ray standing|Calcaneus X-ray standing
C0801762|T102|relax|37206-0|LNC|Calcaneus left X-ray standing|Calcaneus left X-ray standing
C0801762|T102|relax|37720-0|LNC|Calcaneus right X-ray standing|Calcaneus right X-ray standing
C0801762|T102|relax|38845-4|LNC|Femur left X-ray standing|Femur left X-ray standing
C0801762|T102|relax|37693-9|LNC|Femur right X-ray standing|Femur right X-ray standing
C0801762|T102|relax|24708-0|LNC|Foot X-ray standing|Foot X-ray standing
C0801762|T102|relax|26094-3|LNC|Foot bilateral X-ray standing|Foot bilateral X-ray standing
C0801762|T102|relax|26095-0|LNC|Foot left X-ray standing|Foot left X-ray standing
C0801762|T102|relax|26096-8|LNC|Foot right X-ray standing|Foot right X-ray standing
C0801762|T102|relax|37584-0|LNC|Great toe left X-ray standing|Great toe left X-ray standing
C0801762|T102|relax|38810-8|LNC|Great toe right X-ray standing|Great toe right X-ray standing
C0801762|T102|relax|24809-6|LNC|Knee X-ray standing|Knee X-ray standing
C0801762|T102|relax|26085-1|LNC|Knee bilateral X-ray standing|Knee bilateral X-ray standing
C0801762|T102|relax|26086-9|LNC|Knee left X-ray standing|Knee left X-ray standing
C0801762|T102|relax|26087-7|LNC|Knee right X-ray standing|Knee right X-ray standing
C0801762|T102|relax|37204-5|LNC|Lower extremity X-ray standing|Lower extremity X-ray standing
C0801762|T102|relax|69264-0|LNC|Sacrum X-ray standing|Sacrum X-ray standing
C0801762|T102|relax|37208-6|LNC|Spine Lumbar X-ray standing|Spine Lumbar X-ray standing
C0801762|T102|relax|69275-6|LNC|Spine Thoracic X-ray standing|Spine Thoracic X-ray standing
C0801762|T102|relax|38124-4|LNC|Spine Thoracic Lumbar X-ray standing|Spine Thoracic Lumbar X-ray standing
C0801762|T102|relax|37899-2|LNC|Tibia Fibula X-ray standing|Tibia Fibula X-ray standing
C0801762|T102|relax|37209-4|LNC|Toes left X-ray standing|Toes left X-ray standing
C0801762|T102|relax|37823-2|LNC|Toes right X-ray standing|Toes right X-ray standing
C0801762|T102|relax|44233-5|LNC|Kidney bilateral Scan W WO Tc-99m DTPA IV|Kidney bilateral Scan W WO Tc-99m DTPA IV
C0801762|T102|relax|44232-7|LNC|Kidney bilateral Scan W WO Tc-99m Mertiatide IV|Kidney bilateral Scan W WO Tc-99m Mertiatide IV
C0801762|T102|relax|37579-0|LNC|Acromioclavicular Joint X-ray W WO weight|Acromioclavicular Joint X-ray W WO weight
C0801762|T102|relax|37580-8|LNC|Acromioclavicular joint bilateral X-ray W WO weight|Acromioclavicular joint bilateral X-ray W WO weight
C0801762|T102|relax|37581-6|LNC|Acromioclavicular joint left X-ray W WO weight|Acromioclavicular joint left X-ray W WO weight
C0801762|T102|relax|37663-2|LNC|Acromioclavicular joint right X-ray W WO weight|Acromioclavicular joint right X-ray W WO weight
C0801762|T102|relax|39651-5|LNC|Heart Scan W adenosine W Tl-201 IV|Heart Scan W adenosine W Tl-201 IV
C0801762|T102|relax|38090-7|LNC|Breast bilateral Mammogram W air|Breast bilateral Mammogram W air
C0801762|T102|relax|38091-5|LNC|Breast left Mammogram W air|Breast left Mammogram W air
C0801762|T102|relax|39059-1|LNC|Gastrointestine upper Fluoroscopy W air barium contrast PO|Gastrointestine upper Fluoroscopy W air barium contrast PO
C0801762|T102|relax|24666-0|LNC|Colon Fluoroscopy W air barium contrast PR|Colon Fluoroscopy W air barium contrast PR
C0801762|T102|relax|46357-0|LNC|Colon Fluoroscopy W air contrast PR|Colon Fluoroscopy W air contrast PR
C0801762|T102|relax|30633-2|LNC|Esophagus Fluoroscopy W barium contrast PO|Esophagus Fluoroscopy W barium contrast PO
C0801762|T102|relax|42683-3|LNC|Gastrointestine upper Fluoroscopy W barium contrast PO|Gastrointestine upper Fluoroscopy W barium contrast PO
C0801762|T102|relax|43574-3|LNC|Upper Gastrointestine Small bowel Fluoroscopy W barium contrast PO|Upper Gastrointestine Small bowel Fluoroscopy W barium contrast PO
C0801762|T102|relax|44227-7|LNC|Colon Fluoroscopy W barium contrast PR|Colon Fluoroscopy W barium contrast PR
C0801762|T102|relax|37565-9|LNC|Unspecified body region Fluoroscopy W barium contrast via fistula|Unspecified body region Fluoroscopy W barium contrast via fistula
C0801762|T102|relax|38092-3|LNC|Urinary bladder Fluoroscopy W chain contrast intra bladder|Urinary bladder Fluoroscopy W chain contrast intra bladder
C0801762|T102|relax|41770-9|LNC|Gallbladder Scan W cholecystokinin W radionuclide IV|Gallbladder Scan W cholecystokinin W radionuclide IV
C0801762|T102|relax|43650-1|LNC|Liver Biliary ducts Gallbladder Scan W cholecystokinin W radionuclide IV|Liver Biliary ducts Gallbladder Scan W cholecystokinin W radionuclide IV
C0801762|T102|relax|30630-8|LNC|Head Cistern Fluoroscopy video W contrast|Head Cistern Fluoroscopy video W contrast
C0801762|T102|relax|30824-7|LNC|Intercranial vessel Neck Vessel Fluoroscopic angiogram W contrast|Intercranial vessel Neck Vessel Fluoroscopic angiogram W contrast
C0801762|T102|relax|37585-7|LNC|Jejunum Fluoroscopy W contrast|Jejunum Fluoroscopy W contrast
C0801762|T102|relax|38853-8|LNC|Lower extremity vessels left Fluoroscopic angiogram W contrast|Lower extremity vessels left Fluoroscopic angiogram W contrast
C0801762|T102|relax|37765-5|LNC|Lower extremity vessels right Fluoroscopic angiogram W contrast|Lower extremity vessels right Fluoroscopic angiogram W contrast
C0801762|T102|relax|37615-2|LNC|Pelvis vessels Fluoroscopic angiogram W contrast|Pelvis vessels Fluoroscopic angiogram W contrast
C0801762|T102|relax|37936-2|LNC|Peripheral vessels Fluoroscopic angiogram W contrast|Peripheral vessels Fluoroscopic angiogram W contrast
C0801762|T102|relax|37640-0|LNC|Renal vessels Fluoroscopic angiogram W contrast|Renal vessels Fluoroscopic angiogram W contrast
C0801762|T102|relax|64140-7|LNC|Renal vessels left Fluoroscopic angiogram W contrast|Renal vessels left Fluoroscopic angiogram W contrast
C0801762|T102|relax|64141-5|LNC|Renal vessels right Fluoroscopic angiogram W contrast|Renal vessels right Fluoroscopic angiogram W contrast
C0801762|T102|relax|38094-9|LNC|Spine cavity Fluoroscopy W contrast|Spine cavity Fluoroscopy W contrast
C0801762|T102|relax|37973-5|LNC|Testicle vessels Fluoroscopy W contrast|Testicle vessels Fluoroscopy W contrast
C0801762|T102|relax|37976-8|LNC|Upper extremity vessels Fluoroscopic angiogram W contrast|Upper extremity vessels Fluoroscopic angiogram W contrast
C0801762|T102|relax|42014-1|LNC|Urinary Bladder Urethra Fluoroscopy W contrast|Urinary Bladder Urethra Fluoroscopy W contrast
C0801762|T102|relax|37980-0|LNC|Vertebral vessels Fluoroscopic angiogram W contrast|Vertebral vessels Fluoroscopic angiogram W contrast
C0801762|T102|relax|37981-8|LNC|Visceral vessels Fluoroscopic angiogram W contrast|Visceral vessels Fluoroscopic angiogram W contrast
C0801762|T102|relax|37575-8|LNC|Gallbladder X-ray W contrast fatty meal PO|Gallbladder X-ray W contrast fatty meal PO
C0801762|T102|relax|38101-2|LNC|Kidney X-ray W contrast antegrade|Kidney X-ray W contrast antegrade
C0801762|T102|relax|46376-0|LNC|Kidney bilateral Fluoroscopy W contrast antegrade|Kidney bilateral Fluoroscopy W contrast antegrade
C0801762|T102|relax|38100-4|LNC|Urinary Bladder Urethra Fluoroscopy W contrast antegrade|Urinary Bladder Urethra Fluoroscopy W contrast antegrade
C0801762|T102|relax|38102-0|LNC|Kidney X-ray W contrast antegrade via pyelostomy|Kidney X-ray W contrast antegrade via pyelostomy
C0801762|T102|relax|25030-8|LNC|Abdominal Artieries Fluoroscopic angiogram W contrast IA|Abdominal Artieries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30832-0|LNC|Adrenal artery Fluoroscopic angiogram W contrast IA|Adrenal artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30831-2|LNC|Adrenal artery bilateral Fluoroscopic angiogram W contrast IA|Adrenal artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37387-8|LNC|Adrenal artery left Fluoroscopic angiogram W contrast IA|Adrenal artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37939-6|LNC|Adrenal artery right Fluoroscopic angiogram W contrast IA|Adrenal artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|38861-1|LNC|Ankle arteries left Fluoroscopic angiogram W contrast IA|Ankle arteries left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37941-2|LNC|Ankle arteries right Fluoroscopic angiogram W contrast IA|Ankle arteries right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24658-7|LNC|Aorta Fluoroscopic angiogram W contrast IA|Aorta Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30837-9|LNC|Aorta abdominal Fluoroscopic angiogram W contrast IA|Aorta abdominal Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24546-4|LNC|Aorta arch Neck Fluoroscopic angiogram W contrast IA|Aorta arch Neck Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37366-2|LNC|Abdominal Aorta Arteries Fluoroscopic angiogram W contrast IA|Abdominal Aorta Arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|69054-5|LNC|Aortic arch Fluoroscopic angiogram W contrast IA|Aortic arch Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37380-3|LNC|Aortic arch Brachial artery Fluoroscopic angiogram W contrast IA|Aortic arch Brachial artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37381-1|LNC|Aortic arch Carotid artery Fluoroscopic angiogram W contrast IA|Aortic arch Carotid artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37587-3|LNC|Aortic arch Carotid artery bilateral Vertebral artery bilateral Fluoroscopic angiogram W contrast IA|Aortic arch Carotid artery bilateral Vertebral artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37588-1|LNC|Aortic arch Carotid artery common bilateral Fluoroscopic angiogram W contrast IA|Aortic arch Carotid artery common bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37589-9|LNC|Aortic arch Carotid artery common left Fluoroscopic angiogram W contrast IA|Aortic arch Carotid artery common left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37590-7|LNC|Aortic arch Carotid artery common right Fluoroscopic angiogram W contrast IA|Aortic arch Carotid artery common right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37591-5|LNC|Aortic arch Carotid artery external bilateral Fluoroscopic angiogram W contrast IA|Aortic arch Carotid artery external bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37592-3|LNC|Aortic arch Carotid artery external left Fluoroscopic angiogram W contrast IA|Aortic arch Carotid artery external left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37593-1|LNC|Aortic arch Carotid artery external right Fluoroscopic angiogram W contrast IA|Aortic arch Carotid artery external right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37594-9|LNC|Aortic arch Carotid artery Vertebral artery Fluoroscopic angiogram W contrast IA|Aortic arch Carotid artery Vertebral artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37382-9|LNC|Aortic arch Subclavian artery Fluoroscopic angiogram W contrast IA|Aortic arch Subclavian artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37383-7|LNC|Aortic arch Subclavian artery left Fluoroscopic angiogram W contrast IA|Aortic arch Subclavian artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|38800-9|LNC|Aortic arch Subclavian artery right Fluoroscopic angiogram W contrast IA|Aortic arch Subclavian artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37379-5|LNC|Aortic arch Upper Extremity artery Fluoroscopic angiogram W contrast IA|Aortic arch Upper Extremity artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37384-5|LNC|Aortic arch Vertebral artery Fluoroscopic angiogram W contrast IA|Aortic arch Vertebral artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37385-2|LNC|Aortic arch Vertebral artery left Fluoroscopic angiogram W contrast IA|Aortic arch Vertebral artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37386-0|LNC|Aortic arch Vertebral artery right Fluoroscopic angiogram W contrast IA|Aortic arch Vertebral artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24551-4|LNC|AV fistula Fluoroscopic angiogram W contrast IA|AV fistula Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30828-8|LNC|Brachial artery Fluoroscopic angiogram W contrast IA|Brachial artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37388-6|LNC|Brachial artery bilateral Fluoroscopic angiogram W contrast IA|Brachial artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24581-1|LNC|Brachial artery Subclavian artery Fluoroscopic angiogram W contrast IA|Brachial artery Subclavian artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|69077-6|LNC|Brachiocephalic artery Fluoroscopic angiogram W contrast IA|Brachiocephalic artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37389-4|LNC|Bronchial artery Fluoroscopic angiogram W contrast IA|Bronchial artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24617-3|LNC|Carotid artery Fluoroscopic angiogram W contrast IA|Carotid artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|26079-4|LNC|Carotid artery bilateral Fluoroscopic angiogram W contrast IA|Carotid artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|39097-1|LNC|Carotid artery bilateral Cerebral artery bilateral Fluoroscopic angiogram W contrast IA|Carotid artery bilateral Cerebral artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|39094-8|LNC|Carotid artery cervical Fluoroscopic angiogram W contrast IA|Carotid artery cervical Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|39098-9|LNC|Carotid artery cervical bilateral Fluoroscopic angiogram W contrast IA|Carotid artery cervical bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|38863-7|LNC|Carotid artery cervical left Fluoroscopic angiogram W contrast IA|Carotid artery cervical left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37945-3|LNC|Carotid artery cervical right Fluoroscopic angiogram W contrast IA|Carotid artery cervical right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30821-3|LNC|Carotid artery external Fluoroscopic angiogram W contrast IA|Carotid artery external Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30820-5|LNC|Carotid artery external bilateral Fluoroscopic angiogram W contrast IA|Carotid artery external bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37390-2|LNC|Carotid artery external left Fluoroscopic angiogram W contrast IA|Carotid artery external left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37948-7|LNC|Carotid artery external right Fluoroscopic angiogram W contrast IA|Carotid artery external right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|38864-5|LNC|Carotid artery internal left Fluoroscopic angiogram W contrast IA|Carotid artery internal left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37952-9|LNC|Carotid artery internal right Fluoroscopic angiogram W contrast IA|Carotid artery internal right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|26080-2|LNC|Carotid artery left Fluoroscopic angiogram W contrast IA|Carotid artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|26081-0|LNC|Carotid artery right Fluoroscopic angiogram W contrast IA|Carotid artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|39095-5|LNC|Carotid artery Cerebral artery Fluoroscopic angiogram W contrast IA|Carotid artery Cerebral artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|38865-2|LNC|Carotid artery Cerebral artery internal left Fluoroscopic angiogram W contrast IA|Carotid artery Cerebral artery internal left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37953-7|LNC|Carotid artery Cerebral artery internal right Fluoroscopic angiogram W contrast IA|Carotid artery Cerebral artery internal right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|38862-9|LNC|Carotid artery Cerebral artery left Fluoroscopic angiogram W contrast IA|Carotid artery Cerebral artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37944-6|LNC|Carotid artery Cerebral artery right Fluoroscopic angiogram W contrast IA|Carotid artery Cerebral artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37391-0|LNC|Carotid artery Vertebral artery Fluoroscopic angiogram W contrast IA|Carotid artery Vertebral artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37392-8|LNC|Carotid artery Vertebral artery bilateral Fluoroscopic angiogram W contrast IA|Carotid artery Vertebral artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37393-6|LNC|Carotid artery+Vertebral artery left Fluoroscopic angiogram W contrast IA|Carotid artery+Vertebral artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37943-8|LNC|Carotid artery+Vertebral artery right Fluoroscopic angiogram W contrast IA|Carotid artery+Vertebral artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24622-3|LNC|Celiac artery Fluoroscopic angiogram W contrast IA|Celiac artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37403-3|LNC|Celiac artery Gastric artery left Superior mesenteric artery Fluoroscopic angiogram W contrast IA|Celiac artery Gastric artery left Superior mesenteric artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37394-4|LNC|Celiac artery Superior mesenteric artery Inferior mesenteric artery Fluoroscopic angiogram W contrast IA|Celiac artery Superior mesenteric artery Inferior mesenteric artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37173-2|LNC|Cerebral artery Fluoroscopic angiogram W contrast IA|Cerebral artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30891-6|LNC|Cervicocerebral artery Fluoroscopic angiogram W contrast IA|Cervicocerebral artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37174-0|LNC|Coronary arteries Fluoroscopic angiogram W contrast IA|Coronary arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37595-6|LNC|Coronary graft Fluoroscopic angiogram W contrast IA|Coronary graft Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30848-6|LNC|Extremity arteries Fluoroscopic angiogram W contrast IA|Extremity arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30849-4|LNC|Extremity arteries bilateral Fluoroscopic angiogram W contrast IA|Extremity arteries bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37395-1|LNC|Extremity arteries left Fluoroscopic angiogram W contrast IA|Extremity arteries left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37949-5|LNC|Extremity arteries right Fluoroscopic angiogram W contrast IA|Extremity arteries right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37175-7|LNC|Femoral artery Fluoroscopic angiogram W contrast IA|Femoral artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37176-5|LNC|Femoral artery Popliteal artery Fluoroscopic angiogram W contrast IA|Femoral artery Popliteal artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37397-7|LNC|Gastric artery Fluoroscopic angiogram W contrast IA|Gastric artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37398-5|LNC|Gastric artery left Fluoroscopic angiogram W contrast IA|Gastric artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|38801-7|LNC|Gastric artery right Fluoroscopic angiogram W contrast IA|Gastric artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37399-3|LNC|Gastroduodenal artery Fluoroscopic angiogram W contrast IA|Gastroduodenal artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30822-1|LNC|Head artery bilateral Neck artery bilateral Fluoroscopic angiogram W contrast IA|Head artery bilateral Neck artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|62448-6|LNC|Head artery left+Neck artery left Fluoroscopic angiogram W contrast IA|Head artery left+Neck artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|62449-4|LNC|Head artery right+Neck artery right Fluoroscopic angiogram W contrast IA|Head artery right+Neck artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30823-9|LNC|Head artery Neck artery Fluoroscopic angiogram W contrast IA|Head artery Neck artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|25076-1|LNC|Hepatic artery Fluoroscopic angiogram W contrast IA|Hepatic artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|43782-2|LNC|Iliac artery Fluoroscopic angiogram W contrast IA|Iliac artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37177-3|LNC|Iliac artery bilateral Fluoroscopic angiogram W contrast IA|Iliac artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24862-5|LNC|Iliac artery Internal Fluoroscopic angiogram W contrast IA|Iliac artery Internal Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37178-1|LNC|Iliac artery left Fluoroscopic angiogram W contrast IA|Iliac artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37739-0|LNC|Iliac artery right Fluoroscopic angiogram W contrast IA|Iliac artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37179-9|LNC|Inferior mesenteric artery Fluoroscopic angiogram W contrast IA|Inferior mesenteric artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|25079-5|LNC|Kidney arteries Fluoroscopic angiogram W contrast IA|Kidney arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37487-6|LNC|Lower extremity arteries Fluoroscopic angiogram W contrast IA|Lower extremity arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|47986-5|LNC|Lower extremity arteries left Fluoroscopic angiogram W contrast IA|Lower extremity arteries left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|47987-3|LNC|Lower extremity arteries right Fluoroscopic angiogram W contrast IA|Lower extremity arteries right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30829-6|LNC|Internal mammary artery Fluoroscopic angiogram W contrast IA|Internal mammary artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|64995-4|LNC|Mammary artery internal left Fluoroscopic angiogram W contrast IA|Mammary artery internal left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|65000-2|LNC|Mammary artery internal right Fluoroscopic angiogram W contrast IA|Mammary artery internal right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37401-7|LNC|Maxillary artery internal Fluoroscopic angiogram W contrast IA|Maxillary artery internal Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24833-6|LNC|Mesenteric artery Fluoroscopic angiogram W contrast IA|Mesenteric artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24860-9|LNC|Pancreatic artery Fluoroscopic angiogram W contrast IA|Pancreatic artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30833-8|LNC|Pelvis arteries Fluoroscopic angiogram W contrast IA|Pelvis arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37935-4|LNC|Pelvis arteries Lower extremity arteries bilateral Fluoroscopic angiogram W contrast IA|Pelvis arteries Lower extremity arteries bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24874-0|LNC|Peripheral arteries Fluoroscopic angiogram W contrast IA|Peripheral arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|44240-0|LNC|Peripheral arteries bilateral Fluoroscopic angiogram W contrast IA|Peripheral arteries bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|69249-1|LNC|Popliteal artery Fluoroscopic angiogram W contrast IA|Popliteal artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37181-5|LNC|Popliteal artery left Fluoroscopic angiogram W contrast IA|Popliteal artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37778-8|LNC|Popliteal artery right Fluoroscopic angiogram W contrast IA|Popliteal artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37404-1|LNC|Pudendal artery internal Fluoroscopic angiogram W contrast IA|Pudendal artery internal Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|39057-5|LNC|Pulmonary artery Fluoroscopic angiogram W contrast IA|Pulmonary artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30830-4|LNC|Pulmonary artery bilateral Fluoroscopic angiogram W contrast IA|Pulmonary artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37182-3|LNC|Pulmonary artery left Fluoroscopic angiogram W contrast IA|Pulmonary artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37779-6|LNC|Pulmonary artery right Fluoroscopic angiogram W contrast IA|Pulmonary artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|30834-6|LNC|Renal artery bilateral Fluoroscopic angiogram W contrast IA|Renal artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|62446-0|LNC|Renal artery left Fluoroscopic angiogram W contrast IA|Renal artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|62447-8|LNC|Renal artery right Fluoroscopic angiogram W contrast IA|Renal artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24925-0|LNC|Spinal artery Fluoroscopic angiogram W contrast IA|Spinal artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|26082-8|LNC|Spinal artery bilateral Fluoroscopic angiogram W contrast IA|Spinal artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|26083-6|LNC|Spinal artery left Fluoroscopic angiogram W contrast IA|Spinal artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|26084-4|LNC|Spinal artery right Fluoroscopic angiogram W contrast IA|Spinal artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24992-0|LNC|Splenic artery Fluoroscopic angiogram W contrast IA|Splenic artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24991-2|LNC|Splenic vein Portal vein Fluoroscopic angiogram W contrast IA|Splenic vein Portal vein Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37886-9|LNC|Subclavian artery Fluoroscopic angiogram W contrast IA|Subclavian artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37405-8|LNC|Subclavian artery bilateral Fluoroscopic angiogram W contrast IA|Subclavian artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37406-6|LNC|Subclavian artery left Fluoroscopic angiogram W contrast IA|Subclavian artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37966-9|LNC|Subclavian artery right Fluoroscopic angiogram W contrast IA|Subclavian artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37180-7|LNC|Superior mesenteric artery Fluoroscopic angiogram W contrast IA|Superior mesenteric artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37402-5|LNC|Superior mesenteric artery Inferior mesenteric artery Fluoroscopic angiogram W contrast IA|Superior mesenteric artery Inferior mesenteric artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|38119-4|LNC|Thoracic artery Fluoroscopic angiogram W contrast IA|Thoracic artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37900-8|LNC|Tibial artery Fluoroscopic angiogram W contrast IA|Tibial artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37489-2|LNC|Tibioperoneal arteries Fluoroscopic angiogram W contrast IA|Tibioperoneal arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37977-6|LNC|Upper extremity arteries Fluoroscopic angiogram W contrast IA|Upper extremity arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37396-9|LNC|Upper extremity arteries bilateral Fluoroscopic angiogram W contrast IA|Upper extremity arteries bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37488-4|LNC|Upper extremity arteries left Fluoroscopic angiogram W contrast IA|Upper extremity arteries left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37967-7|LNC|Upper extremity arteries right Fluoroscopic angiogram W contrast IA|Upper extremity arteries right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|24576-1|LNC|Urinary bladder arteries Fluoroscopic angiogram W contrast IA|Urinary bladder arteries Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37979-2|LNC|Uterine artery Fluoroscopic angiogram W contrast IA|Uterine artery Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37407-4|LNC|Vertebral artery bilateral Fluoroscopic angiogram W contrast IA|Vertebral artery bilateral Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37490-0|LNC|Vertebral artery left Fluoroscopic angiogram W contrast IA|Vertebral artery left Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|37968-5|LNC|Vertebral artery right Fluoroscopic angiogram W contrast IA|Vertebral artery right Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|42156-0|LNC|Vessels Fluoroscopic angiogram W contrast IA|Vessels Fluoroscopic angiogram W contrast IA
C0801762|T102|relax|25017-5|LNC|Urinary Bladder Urethra Fluoroscopy W contrast intra bladder|Urinary Bladder Urethra Fluoroscopy W contrast intra bladder
C0801762|T102|relax|43559-4|LNC|Urinary Bladder Urethra Fluoroscopy W contrast intra bladder during voiding|Urinary Bladder Urethra Fluoroscopy W contrast intra bladder during voiding
C0801762|T102|relax|37586-5|LNC|Penis Fluoroscopy W contrast intra corpus cavernosum|Penis Fluoroscopy W contrast intra corpus cavernosum
C0801762|T102|relax|39054-2|LNC|Breast duct Mammogram W contrast intra duct|Breast duct Mammogram W contrast intra duct
C0801762|T102|relax|38095-6|LNC|Breast duct bilateral Mammogram W contrast intra duct|Breast duct bilateral Mammogram W contrast intra duct
C0801762|T102|relax|38096-4|LNC|Breast duct left Mammogram W contrast intra duct|Breast duct left Mammogram W contrast intra duct
C0801762|T102|relax|38825-6|LNC|Breast duct right Mammogram W contrast intra duct|Breast duct right Mammogram W contrast intra duct
C0801762|T102|relax|30810-6|LNC|Lacrimal duct Fluoroscopy W contrast intra lacrimal duct|Lacrimal duct Fluoroscopy W contrast intra lacrimal duct
C0801762|T102|relax|38098-0|LNC|Lacrimal duct bilateral Fluoroscopy W contrast intra lacrimal duct|Lacrimal duct bilateral Fluoroscopy W contrast intra lacrimal duct
C0801762|T102|relax|38099-8|LNC|Lacrimal duct left Fluoroscopy W contrast intra lacrimal duct|Lacrimal duct left Fluoroscopy W contrast intra lacrimal duct
C0801762|T102|relax|38827-2|LNC|Lacrimal duct right Fluoroscopy W contrast intra lacrimal duct|Lacrimal duct right Fluoroscopy W contrast intra lacrimal duct
C0801762|T102|relax|24845-0|LNC|Neck Fluoroscopy W contrast intra larynx|Neck Fluoroscopy W contrast intra larynx
C0801762|T102|relax|30850-2|LNC|Extremity lymphatics Fluoroscopy W contrast intra lymphatic|Extremity lymphatics Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|30851-0|LNC|Extremity lymphatics bilateral Fluoroscopy W contrast intra lymphatic|Extremity lymphatics bilateral Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|37599-8|LNC|Extremity lymphatics left Fluoroscopy W contrast intra lymphatic|Extremity lymphatics left Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|38812-4|LNC|Extremity lymphatics right Fluoroscopy W contrast intra lymphatic|Extremity lymphatics right Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|24827-8|LNC|Lymphatics Fluoroscopy W contrast intra lymphatic|Lymphatics Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|30839-5|LNC|Lymphatics abdominal Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|30840-3|LNC|Lymphatics abdominal bilateral Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal bilateral Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|37597-2|LNC|Lymphatics abdominal Lymphatics pelvic Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal Lymphatics pelvic Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|37598-0|LNC|Lymphatics abdominal Lymphatics pelvic bilateral Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal Lymphatics pelvic bilateral Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|37596-4|LNC|Lymphatics abdominal Lymphatics pelvic left Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal Lymphatics pelvic left Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|38811-6|LNC|Lymphatics abdominal Lymphatics pelvic right Fluoroscopy W contrast intra lymphatic|Lymphatics abdominal Lymphatics pelvic right Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|37600-4|LNC|Lymphatics left Fluoroscopy W contrast intra lymphatic|Lymphatics left Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|39510-3|LNC|Lymphatics pelvic Fluoroscopy W contrast intra lymphatic|Lymphatics pelvic Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|37601-2|LNC|Lymphatics pelvic bilateral Fluoroscopy W contrast intra lymphatic|Lymphatics pelvic bilateral Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|38813-2|LNC|Lymphatics right Fluoroscopy W contrast intra lymphatic|Lymphatics right Fluoroscopy W contrast intra lymphatic
C0801762|T102|relax|39148-2|LNC|Breast duct Mammogram W contrast intra multiple ducts|Breast duct Mammogram W contrast intra multiple ducts
C0801762|T102|relax|39146-6|LNC|Breast duct bilateral Mammogram W contrast intra multiple ducts|Breast duct bilateral Mammogram W contrast intra multiple ducts
C0801762|T102|relax|39145-8|LNC|Breast duct left Mammogram W contrast intra multiple ducts|Breast duct left Mammogram W contrast intra multiple ducts
C0801762|T102|relax|39147-4|LNC|Breast duct right Mammogram W contrast intra multiple ducts|Breast duct right Mammogram W contrast intra multiple ducts
C0801762|T102|relax|24661-1|LNC|Pleural space Fluoroscopy W contrast intra pleural space|Pleural space Fluoroscopy W contrast intra pleural space
C0801762|T102|relax|38116-0|LNC|Parotid gland Fluoroscopy W contrast intra salivary duct|Parotid gland Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|38097-2|LNC|Parotid gland left Fluoroscopy W contrast intra salivary duct|Parotid gland left Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|38826-4|LNC|Parotid gland right Fluoroscopy W contrast intra salivary duct|Parotid gland right Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|24902-9|LNC|Salivary gland Fluoroscopy W contrast intra salivary duct|Salivary gland Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|26067-9|LNC|Salivary gland bilateral Fluoroscopy W contrast intra salivary duct|Salivary gland bilateral Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|26068-7|LNC|Salivary gland left Fluoroscopy W contrast intra salivary duct|Salivary gland left Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|26069-5|LNC|Salivary gland right Fluoroscopy W contrast intra salivary duct|Salivary gland right Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|38153-3|LNC|Submandibular gland Fluoroscopy W contrast intra salivary duct|Submandibular gland Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|48698-5|LNC|Submandibular gland bilateral Fluoroscopy W contrast intra salivary duct|Submandibular gland bilateral Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|42460-6|LNC|Submandibular gland left Fluoroscopy W contrast intra salivary duct|Submandibular gland left Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|48696-9|LNC|Submandibular gland right Fluoroscopy W contrast intra salivary duct|Submandibular gland right Fluoroscopy W contrast intra salivary duct
C0801762|T102|relax|24912-8|LNC|Sinus tract Fluoroscopy W contrast intra sinus tract|Sinus tract Fluoroscopy W contrast intra sinus tract
C0801762|T102|relax|24552-2|LNC|Stent Fluoroscopy W contrast intra stent|Stent Fluoroscopy W contrast intra stent
C0801762|T102|relax|25016-7|LNC|Urethra Fluoroscopy W contrast intra urethra|Urethra Fluoroscopy W contrast intra urethra
C0801762|T102|relax|39151-6|LNC|Vas deferens Fluoroscopy W contrast intra vas deferens|Vas deferens Fluoroscopy W contrast intra vas deferens
C0801762|T102|relax|37183-1|LNC|Ankle Fluoroscopy W contrast intraarticular|Ankle Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37184-9|LNC|Ankle bilateral Fluoroscopy W contrast intraarticular|Ankle bilateral Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37185-6|LNC|Ankle left Fluoroscopy W contrast intraarticular|Ankle left Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37942-0|LNC|Ankle right Fluoroscopy W contrast intraarticular|Ankle right Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37186-4|LNC|Elbow Fluoroscopy W contrast intraarticular|Elbow Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37187-2|LNC|Elbow bilateral Fluoroscopy W contrast intraarticular|Elbow bilateral Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37188-0|LNC|Elbow left Fluoroscopy W contrast intraarticular|Elbow left Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37947-9|LNC|Elbow right Fluoroscopy W contrast intraarticular|Elbow right Fluoroscopy W contrast intraarticular
C0801762|T102|relax|24764-3|LNC|Hip Fluoroscopy W contrast intraarticular|Hip Fluoroscopy W contrast intraarticular
C0801762|T102|relax|26070-3|LNC|Hip bilateral Fluoroscopy W contrast intraarticular|Hip bilateral Fluoroscopy W contrast intraarticular
C0801762|T102|relax|26071-1|LNC|Hip left Fluoroscopy W contrast intraarticular|Hip left Fluoroscopy W contrast intraarticular
C0801762|T102|relax|26072-9|LNC|Hip right Fluoroscopy W contrast intraarticular|Hip right Fluoroscopy W contrast intraarticular
C0801762|T102|relax|24800-5|LNC|Knee Fluoroscopy W contrast intraarticular|Knee Fluoroscopy W contrast intraarticular
C0801762|T102|relax|26073-7|LNC|Knee bilateral Fluoroscopy W contrast intraarticular|Knee bilateral Fluoroscopy W contrast intraarticular
C0801762|T102|relax|26074-5|LNC|Knee left Fluoroscopy W contrast intraarticular|Knee left Fluoroscopy W contrast intraarticular
C0801762|T102|relax|26075-2|LNC|Knee right Fluoroscopy W contrast intraarticular|Knee right Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37647-5|LNC|Sacroiliac Joint Fluoroscopy W contrast intraarticular|Sacroiliac Joint Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37189-8|LNC|Sacroiliac joint bilateral Fluoroscopy W contrast intraarticular|Sacroiliac joint bilateral Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37190-6|LNC|Sacroiliac joint left Fluoroscopy W contrast intraarticular|Sacroiliac joint left Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37785-3|LNC|Sacroiliac joint right Fluoroscopy W contrast intraarticular|Sacroiliac joint right Fluoroscopy W contrast intraarticular
C0801762|T102|relax|24910-2|LNC|Shoulder Fluoroscopy W contrast intraarticular|Shoulder Fluoroscopy W contrast intraarticular
C0801762|T102|relax|26076-0|LNC|Shoulder bilateral Fluoroscopy W contrast intraarticular|Shoulder bilateral Fluoroscopy W contrast intraarticular
C0801762|T102|relax|26077-8|LNC|Shoulder left Fluoroscopy W contrast intraarticular|Shoulder left Fluoroscopy W contrast intraarticular
C0801762|T102|relax|26078-6|LNC|Shoulder right Fluoroscopy W contrast intraarticular|Shoulder right Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37901-6|LNC|Temporomandibular joint Fluoroscopy W contrast intraarticular|Temporomandibular joint Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37409-0|LNC|Temporomandibular joint bilateral Fluoroscopy W contrast intraarticular|Temporomandibular joint bilateral Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37410-8|LNC|Temporomandibular joint left Fluoroscopy W contrast intraarticular|Temporomandibular joint left Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37818-2|LNC|Temporomandibular joint right Fluoroscopy W contrast intraarticular|Temporomandibular joint right Fluoroscopy W contrast intraarticular
C0801762|T102|relax|25034-0|LNC|Wrist Fluoroscopy W contrast intraarticular|Wrist Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37570-9|LNC|Wrist bilateral Fluoroscopy W contrast intraarticular|Wrist bilateral Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37571-7|LNC|Wrist left Fluoroscopy W contrast intraarticular|Wrist left Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37641-8|LNC|Wrist right Fluoroscopy W contrast intraarticular|Wrist right Fluoroscopy W contrast intraarticular
C0801762|T102|relax|37191-4|LNC|Joint Fluoroscopy W contrast intraarticular|Joint Fluoroscopy W contrast intraarticular
C0801762|T102|relax|24825-2|LNC|Lung X-ray W contrast intrabronchial|Lung X-ray W contrast intrabronchial
C0801762|T102|relax|30813-0|LNC|Lung bilateral X-ray W contrast intrabronchial|Lung bilateral X-ray W contrast intrabronchial
C0801762|T102|relax|64996-2|LNC|Lung left X-ray W contrast intrabronchial|Lung left X-ray W contrast intrabronchial
C0801762|T102|relax|64997-0|LNC|Lung right X-ray W contrast intrabronchial|Lung right X-ray W contrast intrabronchial
C0801762|T102|relax|37192-2|LNC|Spine Cervical Fluoroscopy W contrast intradisc|Spine Cervical Fluoroscopy W contrast intradisc
C0801762|T102|relax|37193-0|LNC|Spine Lumbar Fluoroscopy W contrast intradisc|Spine Lumbar Fluoroscopy W contrast intradisc
C0801762|T102|relax|70933-7|LNC|Spine Thoracic Fluoroscopy W contrast intradisc|Spine Thoracic Fluoroscopy W contrast intradisc
C0801762|T102|relax|25022-5|LNC|Uterus Fallopian tubes Fluoroscopy W contrast intrauterine|Uterus Fallopian tubes Fluoroscopy W contrast intrauterine
C0801762|T102|relax|30811-4|LNC|Posterior fossa Fluoroscopy W contrast IT|Posterior fossa Fluoroscopy W contrast IT
C0801762|T102|relax|24947-4|LNC|Spine Cervical Fluoroscopy W contrast IT|Spine Cervical Fluoroscopy W contrast IT
C0801762|T102|relax|38103-8|LNC|Spine Cervical Spine Lumbar Fluoroscopy W contrast IT|Spine Cervical Spine Lumbar Fluoroscopy W contrast IT
C0801762|T102|relax|30808-0|LNC|Spine Cervical Thoracic Lumbar Fluoroscopy W contrast IT|Spine Cervical Thoracic Lumbar Fluoroscopy W contrast IT
C0801762|T102|relax|38104-6|LNC|Spine epidural space Fluoroscopy W contrast IT|Spine epidural space Fluoroscopy W contrast IT
C0801762|T102|relax|24974-8|LNC|Spine Lumbar Fluoroscopy W contrast IT|Spine Lumbar Fluoroscopy W contrast IT
C0801762|T102|relax|24985-4|LNC|Spine Thoracic Fluoroscopy W contrast IT|Spine Thoracic Fluoroscopy W contrast IT
C0801762|T102|relax|69066-9|LNC|Abdominal vessels Fluoroscopic angiogram W contrast IV|Abdominal vessels Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30843-7|LNC|Adrenal vein Fluoroscopic angiogram W contrast IV|Adrenal vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37602-0|LNC|Adrenal vein left Fluoroscopic angiogram W contrast IV|Adrenal vein left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30844-5|LNC|Adrenal vein bilateral Fluoroscopic angiogram W contrast IV|Adrenal vein bilateral Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37940-4|LNC|Adrenal vein right Fluoroscopic angiogram W contrast IV|Adrenal vein right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|58746-9|LNC|AV fistula Fluoroscopic angiogram W contrast IV|AV fistula Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|24569-6|LNC|AV shunt Fluoroscopic angiogram W contrast IV|AV shunt Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37411-6|LNC|Azygos vein Fluoroscopic angiogram W contrast IV|Azygos vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|24573-8|LNC|Biliary ducts Gallbladder X-ray W contrast IV|Biliary ducts Gallbladder X-ray W contrast IV
C0801762|T102|relax|37195-5|LNC|Cerebral vein Fluoroscopic angiogram W contrast IV|Cerebral vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30819-7|LNC|Epidural veins Fluoroscopic angiogram W contrast IV|Epidural veins Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|39055-9|LNC|Extremity veins Fluoroscopic angiogram W contrast IV|Extremity veins Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37412-4|LNC|Extremity veins bilateral Fluoroscopic angiogram W contrast IV|Extremity veins bilateral Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37413-2|LNC|Extremity veins left Fluoroscopic angiogram W contrast IV|Extremity veins left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37950-3|LNC|Extremity veins right Fluoroscopic angiogram W contrast IV|Extremity veins right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|42157-8|LNC|Extremity vessels Fluoroscopic angiogram W contrast IV|Extremity vessels Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37416-5|LNC|Femoral vein Fluoroscopic angiogram W contrast IV|Femoral vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|39093-0|LNC|Hepatic veins Fluoroscopic angiogram W contrast IV|Hepatic veins Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37421-5|LNC|Inferior mesenteric vein Fluoroscopic angiogram W contrast IV|Inferior mesenteric vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37419-9|LNC|Intraosseous veins Fluoroscopic angiogram W contrast IV|Intraosseous veins Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37197-1|LNC|Jugular vein Fluoroscopic angiogram W contrast IV|Jugular vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37420-7|LNC|Jugular vein left Fluoroscopic angiogram W contrast IV|Jugular vein left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37954-5|LNC|Jugular vein right Fluoroscopic angiogram W contrast IV|Jugular vein right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37607-9|LNC|Kidney X-ray W contrast IV|Kidney X-ray W contrast IV
C0801762|T102|relax|24788-2|LNC|Kidney bilateral X-ray W contrast IV|Kidney bilateral X-ray W contrast IV
C0801762|T102|relax|37414-0|LNC|Lower extremity veins bilateral Fluoroscopic angiogram W contrast IV|Lower extremity veins bilateral Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37196-3|LNC|Lower extremity veins left Fluoroscopic angiogram W contrast IV|Lower extremity veins left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37767-1|LNC|Lower extremity veins right Fluoroscopic angiogram W contrast IV|Lower extremity veins right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37574-1|LNC|Lower extremity vessels Fluoroscopic angiogram W contrast IV|Lower extremity vessels Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30825-4|LNC|Orbit veins Fluoroscopic angiogram W contrast IV|Orbit veins Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37422-3|LNC|Orbit veins left Fluoroscopic angiogram W contrast IV|Orbit veins left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37958-6|LNC|Orbit veins right Fluoroscopic angiogram W contrast IV|Orbit veins right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30852-8|LNC|Peripheral veins bilateral Fluoroscopic angiogram W contrast IV|Peripheral veins bilateral Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|24685-0|LNC|Peripheral veins Fluoroscopic angiogram W contrast IV|Peripheral veins Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|69250-9|LNC|Portal vein Fluoroscopic angiogram W contrast IV|Portal vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30847-8|LNC|Renal vein Fluoroscopic angiogram W contrast IV|Renal vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30846-0|LNC|Renal vein bilateral Fluoroscopic angiogram W contrast IV|Renal vein bilateral Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37423-1|LNC|Renal vein left Fluoroscopic angiogram W contrast IV|Renal vein left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37959-4|LNC|Renal vein right Fluoroscopic angiogram W contrast IV|Renal vein right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30827-0|LNC|Sagittal sinus vein Fluoroscopic angiogram W contrast IV|Sagittal sinus vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|65803-9|LNC|Sagittal sinus vein left Fluoroscopic angiogram W contrast IV|Sagittal sinus vein left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|65802-1|LNC|Sagittal sinus Jugular veins left Fluoroscopic angiogram W contrast IV|Sagittal sinus Jugular veins left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|65804-7|LNC|Sagittal sinus vein right Fluoroscopic angiogram W contrast IV|Sagittal sinus vein right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|65805-4|LNC|Sagittal sinus Jugular veins right Fluoroscopic angiogram W contrast IV|Sagittal sinus Jugular veins right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30826-2|LNC|Sagittal sinus Jugular veins Fluoroscopic angiogram W contrast IV|Sagittal sinus Jugular veins Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37969-3|LNC|Sinus vein Fluoroscopic angiogram W contrast IV|Sinus vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37970-1|LNC|Splenic vein Fluoroscopic angiogram W contrast IV|Splenic vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37971-9|LNC|Subclavian vein Fluoroscopic angiogram W contrast IV|Subclavian vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37972-7|LNC|Superior mesenteric vein Fluoroscopic angiogram W contrast IV|Superior mesenteric vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|24550-6|LNC|Upper extremity veins Fluoroscopic angiogram W contrast IV|Upper extremity veins Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37415-7|LNC|Upper extremity veins bilateral Fluoroscopic angiogram W contrast IV|Upper extremity veins bilateral Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|38859-5|LNC|Upper extremity veins left Fluoroscopic angiogram W contrast IV|Upper extremity veins left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|37824-0|LNC|Upper extremity veins right Fluoroscopic angiogram W contrast IV|Upper extremity veins right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|25023-3|LNC|Vein Fluoroscopic angiogram W contrast IV|Vein Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|26064-6|LNC|Vein bilateral Fluoroscopic angiogram W contrast IV|Vein bilateral Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|26065-3|LNC|Vein left Fluoroscopic angiogram W contrast IV|Vein left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|26066-1|LNC|Vein right Fluoroscopic angiogram W contrast IV|Vein right Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|25025-8|LNC|Vena cava Fluoroscopic angiogram W contrast IV|Vena cava Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30845-2|LNC|Inferior vena cava Fluoroscopic angiogram W contrast IV|Inferior vena cava Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|30645-6|LNC|Superior vena cava Fluoroscopic angiogram W contrast IV|Superior vena cava Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|43554-5|LNC|vessels left Fluoroscopic angiogram W contrast IV|vessels left Fluoroscopic angiogram W contrast IV
C0801762|T102|relax|39096-3|LNC|Hepatic veins Fluoroscopic angiogram W contrast IV W hemodynamics|Hepatic veins Fluoroscopic angiogram W contrast IV W hemodynamics
C0801762|T102|relax|43783-0|LNC|Renal vein Fluoroscopic angiogram W contrast IV W renin sampling|Renal vein Fluoroscopic angiogram W contrast IV W renin sampling
C0801762|T102|relax|25080-3|LNC|Renal vein bilateral Fluoroscopic angiogram W contrast IV W renin sampling|Renal vein bilateral Fluoroscopic angiogram W contrast IV W renin sampling
C0801762|T102|relax|30816-3|LNC|Peritoneum Fluoroscopic angiogram W contrast percutaneous|Peritoneum Fluoroscopic angiogram W contrast percutaneous
C0801762|T102|relax|24575-3|LNC|Biliary ducts Gallbladder Fluoroscopy W contrast percutaneous transhepatic|Biliary ducts Gallbladder Fluoroscopy W contrast percutaneous transhepatic
C0801762|T102|relax|37200-3|LNC|Chest X-ray W contrast PO|Chest X-ray W contrast PO
C0801762|T102|relax|37199-7|LNC|Chest Fluoroscopy W contrast PO|Chest Fluoroscopy W contrast PO
C0801762|T102|relax|37198-9|LNC|Esophagus X-ray W contrast PO|Esophagus X-ray W contrast PO
C0801762|T102|relax|24678-5|LNC|Esophagus Fluoroscopy W contrast PO|Esophagus Fluoroscopy W contrast PO
C0801762|T102|relax|24712-2|LNC|Gallbladder X-ray W contrast PO|Gallbladder X-ray W contrast PO
C0801762|T102|relax|42459-8|LNC|Gastrointestine upper Fluoroscopy W contrast PO|Gastrointestine upper Fluoroscopy W contrast PO
C0801762|T102|relax|24924-3|LNC|Small bowel Fluoroscopy W contrast PO|Small bowel Fluoroscopy W contrast PO
C0801762|T102|relax|24673-6|LNC|Duodenum Fluoroscopy W contrast PO hypotonic agent per ng|Duodenum Fluoroscopy W contrast PO hypotonic agent per ng
C0801762|T102|relax|24681-9|LNC|Esophagus Hypopharynx Fluoroscopy video W contrast PO during swallowing|Esophagus Hypopharynx Fluoroscopy video W contrast PO during swallowing
C0801762|T102|relax|24667-8|LNC|Colon Fluoroscopy W contrast PR|Colon Fluoroscopy W contrast PR
C0801762|T102|relax|24894-8|LNC|Rectum Urinary bladder Fluoroscopy W contrast PR intra bladder during defecation voiding|Rectum Urinary bladder Fluoroscopy W contrast PR intra bladder during defecation voiding
C0801762|T102|relax|39363-7|LNC|Fistula Fluoroscopy W contrast retrograde|Fistula Fluoroscopy W contrast retrograde
C0801762|T102|relax|38105-3|LNC|Kidney X-ray W contrast retrograde|Kidney X-ray W contrast retrograde
C0801762|T102|relax|39349-6|LNC|Kidney bilateral Fluoroscopy W contrast retrograde|Kidney bilateral Fluoroscopy W contrast retrograde
C0801762|T102|relax|30761-1|LNC|Kidney bilateral Fluoroscopy W contrast retrograde via urethra|Kidney bilateral Fluoroscopy W contrast retrograde via urethra
C0801762|T102|relax|38873-6|LNC|Kidney left Collecting system Fluoroscopy W contrast retrograde via urethra|Kidney left Collecting system Fluoroscopy W contrast retrograde via urethra
C0801762|T102|relax|38113-7|LNC|Kidney right Collecting system Fluoroscopy W contrast retrograde via urethra|Kidney right Collecting system Fluoroscopy W contrast retrograde via urethra
C0801762|T102|relax|25020-9|LNC|Urinary Bladder Urethra Fluoroscopy W contrast retrograde via urethra|Urinary Bladder Urethra Fluoroscopy W contrast retrograde via urethra
C0801762|T102|relax|30841-1|LNC|Portal vein Fluoroscopic angiogram W contrast transhepatic|Portal vein Fluoroscopic angiogram W contrast transhepatic
C0801762|T102|relax|30842-9|LNC|Portal vein Fluoroscopic angiogram W contrast transhepatic W hemodynamics|Portal vein Fluoroscopic angiogram W contrast transhepatic W hemodynamics
C0801762|T102|relax|37566-7|LNC|Unspecified body region Fluoroscopy W contrast via catheter|Unspecified body region Fluoroscopy W contrast via catheter
C0801762|T102|relax|37567-5|LNC|Colon Fluoroscopy W contrast via colostomy|Colon Fluoroscopy W contrast via colostomy
C0801762|T102|relax|37568-3|LNC|Unspecified body region Fluoroscopy W contrast via fistula|Unspecified body region Fluoroscopy W contrast via fistula
C0801762|T102|relax|69272-3|LNC|Small bowel Fluoroscopy W contrast via ileostomy|Small bowel Fluoroscopy W contrast via ileostomy
C0801762|T102|relax|24780-9|LNC|Kidney bilateral Fluoroscopy W contrast via nephrostomy tube|Kidney bilateral Fluoroscopy W contrast via nephrostomy tube
C0801762|T102|relax|38872-8|LNC|Kidney left Collecting system Fluoroscopy W contrast via nephrostomy tube|Kidney left Collecting system Fluoroscopy W contrast via nephrostomy tube
C0801762|T102|relax|38112-9|LNC|Kidney right Collecting system Fluoroscopy W contrast via nephrostomy tube|Kidney right Collecting system Fluoroscopy W contrast via nephrostomy tube
C0801762|T102|relax|37569-1|LNC|Urinary bladder Fluoroscopy W contrast via suprapubic tube|Urinary bladder Fluoroscopy W contrast via suprapubic tube
C0801762|T102|relax|30647-2|LNC|Biliary ducts Gallbladder Fluoroscopy W contrast via T-tube|Biliary ducts Gallbladder Fluoroscopy W contrast via T-tube
C0801762|T102|relax|39696-0|LNC|Lung Scan W depreotide W radionuclide IV|Lung Scan W depreotide W radionuclide IV
C0801762|T102|relax|42161-0|LNC|Heart Scan W dobutamine W radionuclide IV|Heart Scan W dobutamine W radionuclide IV
C0801762|T102|relax|39652-3|LNC|Heart Scan W dobutamine W Tl-201 IV|Heart Scan W dobutamine W Tl-201 IV
C0801762|T102|relax|42383-0|LNC|Gallbladder X-ray W double dose contrast PO|Gallbladder X-ray W double dose contrast PO
C0801762|T102|relax|42690-8|LNC|Spine X-ray W flexion W extension|Spine X-ray W flexion W extension
C0801762|T102|relax|24945-8|LNC|Spine Cervical X-ray W flexion W extension|Spine Cervical X-ray W flexion W extension
C0801762|T102|relax|24971-4|LNC|Spine Lumbar X-ray W flexion W extension|Spine Lumbar X-ray W flexion W extension
C0801762|T102|relax|43481-1|LNC|Joint X-ray W flexion W extension|Joint X-ray W flexion W extension
C0801762|T102|relax|30785-0|LNC|Foot X-ray W forced dorsiflexion|Foot X-ray W forced dorsiflexion
C0801762|T102|relax|43461-3|LNC|Kidney bilateral Scan W furosemide W radionuclide IV|Kidney bilateral Scan W furosemide W radionuclide IV
C0801762|T102|relax|39688-7|LNC|Scan W GA-67 IV|Scan W GA-67 IV
C0801762|T102|relax|24679-3|LNC|Esophagus Fluoroscopy W gastrografin PO|Esophagus Fluoroscopy W gastrografin PO
C0801762|T102|relax|42684-1|LNC|Gastrointestine upper Fluoroscopy W gastrografin PO|Gastrointestine upper Fluoroscopy W gastrografin PO
C0801762|T102|relax|42681-7|LNC|Colon Fluoroscopy W gastrografin PR|Colon Fluoroscopy W gastrografin PR
C0801762|T102|relax|37576-6|LNC|Unspecified body region Fluoroscopy W gastrografin via fistula|Unspecified body region Fluoroscopy W gastrografin via fistula
C0801762|T102|relax|39850-3|LNC|Kidney bilateral Scan W I-131 IV|Kidney bilateral Scan W I-131 IV
C0801762|T102|relax|25007-6|LNC|Thyroid Scan W I-131 IV|Thyroid Scan W I-131 IV
C0801762|T102|relax|39841-2|LNC|Scan W I-131 MIBG IV|Scan W I-131 MIBG IV
C0801762|T102|relax|39857-8|LNC|Adrenal gland Scan W I-131 MIBG IV|Adrenal gland Scan W I-131 MIBG IV
C0801762|T102|relax|39624-2|LNC|Adrenal gland Scan W I-131 NP59 IV|Adrenal gland Scan W I-131 NP59 IV
C0801762|T102|relax|24770-0|LNC|Joint Scan W In-111 intrajoint|Joint Scan W In-111 intrajoint
C0801762|T102|relax|39846-1|LNC|Scan W In-111 Satumomab IV|Scan W In-111 Satumomab IV
C0801762|T102|relax|39738-0|LNC|Abdomen Scan W In-111 Satumomab IV|Abdomen Scan W In-111 Satumomab IV
C0801762|T102|relax|25032-4|LNC|Bone Scan W In-111 tagged WBC IV|Bone Scan W In-111 tagged WBC IV
C0801762|T102|relax|42708-8|LNC|Scan W In-111 tiuxetan IV|Scan W In-111 tiuxetan IV
C0801762|T102|relax|30736-3|LNC|Chest X-ray W inspiration expiration|Chest X-ray W inspiration expiration
C0801762|T102|relax|24682-7|LNC|Esophagus Hypopharynx Fluoroscopy video W liquid paste contrast PO during swallowing|Esophagus Hypopharynx Fluoroscopy video W liquid paste contrast PO during swallowing
C0801762|T102|relax|37556-8|LNC|Ankle X-ray W manual stress|Ankle X-ray W manual stress
C0801762|T102|relax|37557-6|LNC|Ankle bilateral X-ray W manual stress|Ankle bilateral X-ray W manual stress
C0801762|T102|relax|37558-4|LNC|Ankle left X-ray W manual stress|Ankle left X-ray W manual stress
C0801762|T102|relax|37673-1|LNC|Ankle right X-ray W manual stress|Ankle right X-ray W manual stress
C0801762|T102|relax|37559-2|LNC|Foot left X-ray W manual stress|Foot left X-ray W manual stress
C0801762|T102|relax|37705-1|LNC|Foot right X-ray W manual stress|Foot right X-ray W manual stress
C0801762|T102|relax|37560-0|LNC|Knee X-ray W manual stress|Knee X-ray W manual stress
C0801762|T102|relax|37561-8|LNC|Knee bilateral X-ray W manual stress|Knee bilateral X-ray W manual stress
C0801762|T102|relax|37562-6|LNC|Knee left X-ray W manual stress|Knee left X-ray W manual stress
C0801762|T102|relax|37753-1|LNC|Knee right X-ray W manual stress|Knee right X-ray W manual stress
C0801762|T102|relax|37563-4|LNC|Thumb bilateral X-ray W manual stress|Thumb bilateral X-ray W manual stress
C0801762|T102|relax|37564-2|LNC|Thumb left X-ray W manual stress|Thumb left X-ray W manual stress
C0801762|T102|relax|37814-1|LNC|Thumb right X-ray W manual stress|Thumb right X-ray W manual stress
C0801762|T102|relax|39056-7|LNC|Unspecified body region X-ray W manual stress|Unspecified body region X-ray W manual stress
C0801762|T102|relax|38093-1|LNC|Chest X-ray W nipple markers|Chest X-ray W nipple markers
C0801762|T102|relax|39670-5|LNC|Lacrimal duct Scan W radionuclide intra lacrimal duct|Lacrimal duct Scan W radionuclide intra lacrimal duct
C0801762|T102|relax|64051-6|LNC|Breast lymphatics left Scan W radionuclide intra lymphatic|Breast lymphatics left Scan W radionuclide intra lymphatic
C0801762|T102|relax|64052-4|LNC|Breast lymphatics right Scan W radionuclide intra lymphatic|Breast lymphatics right Scan W radionuclide intra lymphatic
C0801762|T102|relax|24826-0|LNC|Lymphatics Scan W radionuclide intra lymphatic|Lymphatics Scan W radionuclide intra lymphatic
C0801762|T102|relax|24663-7|LNC|Head Cistern Scan W radionuclide IT|Head Cistern Scan W radionuclide IT
C0801762|T102|relax|42158-6|LNC|Adrenal gland Scan|Adrenal gland Scan
C0801762|T102|relax|42776-5|LNC|AV shunt Scan|AV shunt Scan
C0801762|T102|relax|25031-6|LNC|Bone Scan|Bone Scan
C0801762|T102|relax|24730-4|LNC|Brain Scan|Brain Scan
C0801762|T102|relax|39643-2|LNC|Brain veins Scan|Brain veins Scan
C0801762|T102|relax|39646-5|LNC|Breast Scan|Breast Scan
C0801762|T102|relax|39650-7|LNC|Heart Scan|Heart Scan
C0801762|T102|relax|24776-7|LNC|Kidney bilateral Scan|Kidney bilateral Scan
C0801762|T102|relax|30877-5|LNC|Kidney bilateral Renal vessels Scan|Kidney bilateral Renal vessels Scan
C0801762|T102|relax|24804-7|LNC|Knee Scan|Knee Scan
C0801762|T102|relax|26088-5|LNC|Knee bilateral Scan|Knee bilateral Scan
C0801762|T102|relax|26089-3|LNC|Knee left Scan|Knee left Scan
C0801762|T102|relax|26090-1|LNC|Knee right Scan|Knee right Scan
C0801762|T102|relax|39693-7|LNC|Liver Scan|Liver Scan
C0801762|T102|relax|39694-5|LNC|Liver transplant Scan|Liver transplant Scan
C0801762|T102|relax|43557-8|LNC|Liver Biliary ducts Gallbladder Scan|Liver Biliary ducts Gallbladder Scan
C0801762|T102|relax|39897-4|LNC|Liver Lung Scan|Liver Lung Scan
C0801762|T102|relax|39877-6|LNC|Liver Spleen Scan|Liver Spleen Scan
C0801762|T102|relax|39629-1|LNC|Meckels diverticulum Scan|Meckels diverticulum Scan
C0801762|T102|relax|39737-2|LNC|Neck Scan|Neck Scan
C0801762|T102|relax|39739-8|LNC|Pancreas Scan|Pancreas Scan
C0801762|T102|relax|39742-2|LNC|Parathyroid Scan|Parathyroid Scan
C0801762|T102|relax|39619-2|LNC|Pulmonary system Scan|Pulmonary system Scan
C0801762|T102|relax|43669-1|LNC|Renal vessels Scan|Renal vessels Scan
C0801762|T102|relax|39747-1|LNC|Salivary gland Scan|Salivary gland Scan
C0801762|T102|relax|30696-9|LNC|Scrotum Testicle Scan|Scrotum Testicle Scan
C0801762|T102|relax|39751-3|LNC|Spleen Scan|Spleen Scan
C0801762|T102|relax|30695-1|LNC|Thyroid Scan|Thyroid Scan
C0801762|T102|relax|25018-3|LNC|Urinary bladder Scan|Urinary bladder Scan
C0801762|T102|relax|39626-7|LNC|Vein bilateral Scan|Vein bilateral Scan
C0801762|T102|relax|49118-3|LNC|Unspecified body region Scan|Unspecified body region Scan
C0801762|T102|relax|39939-4|LNC|Joint Scan|Joint Scan
C0801762|T102|relax|39671-3|LNC|Rectum Scan W radionuclide PO|Rectum Scan W radionuclide PO
C0801762|T102|relax|39752-1|LNC|Spleen Scan W radionuclide tagged heat damaged RBC IV|Spleen Scan W radionuclide tagged heat damaged RBC IV
C0801762|T102|relax|24773-4|LNC|Kidney bilateral Scan W radionuclide transplant scan|Kidney bilateral Scan W radionuclide transplant scan
C0801762|T102|relax|30713-2|LNC|Spine X-ray W right bending W left bending|Spine X-ray W right bending W left bending
C0801762|T102|relax|42413-5|LNC|Spine Lumbar X-ray W right bending W left bending|Spine Lumbar X-ray W right bending W left bending
C0801762|T102|relax|43651-9|LNC|Liver Biliary ducts Gallbladder Scan W sincalide W radionuclide IV|Liver Biliary ducts Gallbladder Scan W sincalide W radionuclide IV
C0801762|T102|relax|39820-6|LNC|Bone Scan W SM153 IV|Bone Scan W SM153 IV
C0801762|T102|relax|39666-3|LNC|Heart Scan W stress W 201 Th IV|Heart Scan W stress W 201 Th IV
C0801762|T102|relax|39667-1|LNC|Heart Scan W stress W radionuclide IV|Heart Scan W stress W radionuclide IV
C0801762|T102|relax|69231-9|LNC|Heart Scan W stress W Tc-99m IV|Heart Scan W stress W Tc-99m IV
C0801762|T102|relax|69232-7|LNC|Heart Scan W stress W Tc-99m Sestamibi IV|Heart Scan W stress W Tc-99m Sestamibi IV
C0801762|T102|relax|24819-5|LNC|Liver Spleen Scan W Tc-99m calcium colloid IV|Liver Spleen Scan W Tc-99m calcium colloid IV
C0801762|T102|relax|39744-8|LNC|Prostate Scan W Tc-99m capromab pendatide IV|Prostate Scan W Tc-99m capromab pendatide IV
C0801762|T102|relax|39674-7|LNC|Gallbladder Scan W Tc-99m DISIDA IV|Gallbladder Scan W Tc-99m DISIDA IV
C0801762|T102|relax|41771-7|LNC|Kidney bilateral Scan W Tc-99m DMSA IV|Kidney bilateral Scan W Tc-99m DMSA IV
C0801762|T102|relax|39625-9|LNC|Artery Scan W Tc-99m DTPA IA|Artery Scan W Tc-99m DTPA IA
C0801762|T102|relax|39745-5|LNC|Kidney bilateral Scan W Tc-99m DTPA IV|Kidney bilateral Scan W Tc-99m DTPA IV
C0801762|T102|relax|43667-5|LNC|Kidney bilateral Renal vessels Scan W Tc-99m DTPA IV|Kidney bilateral Renal vessels Scan W Tc-99m DTPA IV
C0801762|T102|relax|39753-9|LNC|Scrotum Testicle Scan W Tc-99m DTPA IV|Scrotum Testicle Scan W Tc-99m DTPA IV
C0801762|T102|relax|39765-3|LNC|Vein Scan W Tc-99m DTPA IV|Vein Scan W Tc-99m DTPA IV
C0801762|T102|relax|39642-4|LNC|Brain Scan W Tc-99m glucoheptonate IV|Brain Scan W Tc-99m glucoheptonate IV
C0801762|T102|relax|44234-3|LNC|Kidney bilateral Scan W Tc-99m glucoheptonate IV|Kidney bilateral Scan W Tc-99m glucoheptonate IV
C0801762|T102|relax|39766-1|LNC|Vein Scan W Tc-99m HDP IV|Vein Scan W Tc-99m HDP IV
C0801762|T102|relax|39812-3|LNC|Bone Scan W Tc-99m HMPAO IV|Bone Scan W Tc-99m HMPAO IV
C0801762|T102|relax|39630-9|LNC|Brain Scan W Tc-99m HMPAO IV|Brain Scan W Tc-99m HMPAO IV
C0801762|T102|relax|39757-0|LNC|Thyroid Scan W Tc-99m IV|Thyroid Scan W Tc-99m IV
C0801762|T102|relax|24831-0|LNC|Meckels diverticulum Scan W Tc-99m M04 IV|Meckels diverticulum Scan W Tc-99m M04 IV
C0801762|T102|relax|44141-0|LNC|Liver Spleen Scan W Tc-99m MAA IV|Liver Spleen Scan W Tc-99m MAA IV
C0801762|T102|relax|44142-8|LNC|Bone Scan W Tc-99m medronate IV|Bone Scan W Tc-99m medronate IV
C0801762|T102|relax|39746-3|LNC|Kidney bilateral Scan W Tc-99m Mertiatide IV|Kidney bilateral Scan W Tc-99m Mertiatide IV
C0801762|T102|relax|69233-5|LNC|Parotid gland Scan W Tc-99m pertechnetate IV|Parotid gland Scan W Tc-99m pertechnetate IV
C0801762|T102|relax|25001-9|LNC|Scrotum Testicle Scan W Tc-99m pertechnetate IV|Scrotum Testicle Scan W Tc-99m pertechnetate IV
C0801762|T102|relax|26091-9|LNC|Scrotum Testicle bilateral Scan W Tc-99m pertechnetate IV|Scrotum Testicle bilateral Scan W Tc-99m pertechnetate IV
C0801762|T102|relax|26092-7|LNC|Scrotum Testicle left Scan W Tc-99m pertechnetate IV|Scrotum Testicle left Scan W Tc-99m pertechnetate IV
C0801762|T102|relax|26093-5|LNC|Scrotum Testicle right Scan W Tc-99m pertechnetate IV|Scrotum Testicle right Scan W Tc-99m pertechnetate IV
C0801762|T102|relax|44146-9|LNC|Bone marrow Scan W Tc-99m SC IV|Bone marrow Scan W Tc-99m SC IV
C0801762|T102|relax|39689-5|LNC|Gastrointestine Scan W Tc-99m SC IV|Gastrointestine Scan W Tc-99m SC IV
C0801762|T102|relax|69230-1|LNC|Liver Scan W Tc-99m SC IV|Liver Scan W Tc-99m SC IV
C0801762|T102|relax|39764-6|LNC|Vein Scan W Tc-99m SC IV|Vein Scan W Tc-99m SC IV
C0801762|T102|relax|24683-5|LNC|Esophagus Stomach Scan W Tc-99m SC PO|Esophagus Stomach Scan W Tc-99m SC PO
C0801762|T102|relax|44145-1|LNC|Parathyroid Scan W Tc-99m Sestamibi IV|Parathyroid Scan W Tc-99m Sestamibi IV
C0801762|T102|relax|39756-2|LNC|Thyroid Scan W Tc-99m Sestamibi IV|Thyroid Scan W Tc-99m Sestamibi IV
C0801762|T102|relax|24714-8|LNC|Gastrointestine Scan W Tc-99m tagged RBC IV|Gastrointestine Scan W Tc-99m tagged RBC IV
C0801762|T102|relax|44143-6|LNC|Heart Scan W Tc-99m tagged RBC IV|Heart Scan W Tc-99m tagged RBC IV
C0801762|T102|relax|39690-3|LNC|Liver Scan W Tc-99m tagged RBC IV|Liver Scan W Tc-99m tagged RBC IV
C0801762|T102|relax|42700-5|LNC|Bone Scan W Tc-99m tagged WBC IV|Bone Scan W Tc-99m tagged WBC IV
C0801762|T102|relax|24751-0|LNC|Parathyroid Scan W TI-201 subtraction Tc-99m IV|Parathyroid Scan W TI-201 subtraction Tc-99m IV
C0801762|T102|relax|39635-8|LNC|Brain Scan W Tl-201 IV|Brain Scan W Tl-201 IV
C0801762|T102|relax|51389-5|LNC|Breast Scan W Tl-201 IV|Breast Scan W Tl-201 IV
C0801762|T102|relax|42012-5|LNC|Gastrointestine upper Fluoroscopy W water soluble contrast PO|Gastrointestine upper Fluoroscopy W water soluble contrast PO
C0801762|T102|relax|24669-4|LNC|Colon Fluoroscopy W water soluble contrast PR|Colon Fluoroscopy W water soluble contrast PR
C0801762|T102|relax|37577-4|LNC|Acromioclavicular Joint X-ray W weight|Acromioclavicular Joint X-ray W weight
C0801762|T102|relax|37578-2|LNC|Acromioclavicular joint bilateral X-ray W weight|Acromioclavicular joint bilateral X-ray W weight
C0801762|T102|relax|44144-4|LNC|Liver Scan W Xe-133 inhaled|Liver Scan W Xe-133 inhaled
C0801762|T102|relax|37582-4|LNC|Acromioclavicular Joint X-ray WO weight|Acromioclavicular Joint X-ray WO weight
C0801762|T102|relax|69055-2|LNC|Acromioclavicular joint bilateral X-ray WO weight|Acromioclavicular joint bilateral X-ray WO weight