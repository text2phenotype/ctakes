C0024808|T053|228997001|SNOMEDCT_US|SMOKES WEED|MARIHUANA
C0024808|T053|228997001|SNOMEDCT_US|WEED SMOKER|MARIHUANA
C0024808|T053|228997001|SNOMEDCT_US|MARIJUANA SMOKER|MARIHUANA
C0024808|T053|228997001|SNOMEDCT_US|SMOKES MARIJUANA|MARIHUANA
C0024808|T053|228997001|SNOMEDCT_US|MARIHUANA|MARIHUANA
C0024809|T053||SNOMEDCT_US|MARIJUANA ABUSE
C0678449|T053|398705004|SNOMEDCT_US|CANNABIS SUBSTANCE|CANNABIS
C0936079|T053|22924007|SNOMEDCT_US|CANNABIS|CANNABIS (ORGANISM)
C0936079|T053|22924007|SNOMEDCT_US|CANNABIS SMOKER|CANNABIS (ORGANISM)
C0936079|T053|22924007|SNOMEDCT_US|SMOKES CANNABIS|CANNABIS (ORGANISM)
C1547291|T053||SNOMEDCT_US|MARIJUANA RECREATIONAL DRUG USE CODE
C0024808|T053|228997001|SNOMEDCT_US|MARIHUANA|MARIHUANA
C0024808|T053|228997001|SNOMEDCT_US|MARIJUANA|MARIHUANA
C0024808|T053|228997001|SNOMEDCT_US|CANNABIS|MARIHUANA
C0024808|T053|228997001|SNOMEDCT_US|MARIJUANAS|MARIHUANA
C0024808|T053|228997001|SNOMEDCT_US|MARIHUANAS|MARIHUANA
C0024808|T053|228997001|SNOMEDCT_US|MARIJUANA [VA PRODUCT]|MARIHUANA
C0024809|T053||SNOMEDCT_US|ABUSE, MARIHUANA
C0024809|T053||SNOMEDCT_US|ABUSE, MARIJUANA
C0024809|T053||SNOMEDCT_US|MARIJUANA ABUSE
C0024809|T053||SNOMEDCT_US|MARIJUANA
C0024809|T053||SNOMEDCT_US|MARIHUANA ABUSE
C0024809|T053||SNOMEDCT_US|MARIJUANA ABUSE [DISEASE/FINDING]
C0024809|T053||SNOMEDCT_US|ABUSE;DRUG(S);MARIJUANA
C0024809|T053||SNOMEDCT_US|CANNABIS
# C0024809|T053||SNOMEDCT_US|HASH
# C0024809|T053||SNOMEDCT_US|WEED
# C0024809|T053||SNOMEDCT_US|POT
C0024809|T053||SNOMEDCT_US|HASH USER 
C0024809|T053||SNOMEDCT_US|WEED USER 
C0024809|T053||SNOMEDCT_US|POT USER
C0024809|T053||SNOMEDCT_US|USES HASH
C0024809|T053||SNOMEDCT_US|USES WEED
C0024809|T053||SNOMEDCT_US|USES POT
C0024809|T053||SNOMEDCT_US|ABUSE; MARIHUANA
C0024809|T053||SNOMEDCT_US|MARIHUANA; ABUSE
C0018614|T053||SNOMEDCT_US|ABUSE, HASHISH
C0018614|T053||SNOMEDCT_US|HASHISH; ABUSE
C0018614|T053||SNOMEDCT_US|ABUSE; HASHISH
C0018614|T053||SNOMEDCT_US|HASHISH ABUSE
C0017089|T053||SNOMEDCT_US|GANJAS
C0017089|T053||SNOMEDCT_US|GANJA
C0018210|T053|422304003|SNOMEDCT_US|GRAMINEAE|FAMILY POACEAE
C0018210|T053|422304003|SNOMEDCT_US|POACEAE|FAMILY POACEAE
C0006863|T053|96223000|SNOMEDCT_US|CANNABIDIOL|CANNABIDIOL (SUBSTANCE)
C0006863|T053|96223000|SNOMEDCT_US|1,3-BENZENEDIOL, 2-(3-METHYL-6-(1-METHYLETHENYL)-2-CYCLOHEXEN-1-YL)-5-PENTYL-, (1R-TRANS)-|CANNABIDIOL (SUBSTANCE)
C0006863|T053|96223000|SNOMEDCT_US|CANNABIDIOL [CHEMICAL/INGREDIENT]|CANNABIDIOL (SUBSTANCE)
C0006863|T053|96223000|SNOMEDCT_US|CBD|CANNABIDIOL (SUBSTANCE)
C0006863|T053|96223000|SNOMEDCT_US|CANNABIDIOL |CANNABIDIOL (SUBSTANCE)
C0006865|T053|96222005|SNOMEDCT_US|CANNABINOL|CANNABINOL (SUBSTANCE)
C0006865|T053|96222005|SNOMEDCT_US|6H-DIBENZO(B,D)PYRAN-1-OL, 6,6,9-TRIMETHYL-3-PENTYL-|CANNABINOL (SUBSTANCE)
C0006865|T053|96222005|SNOMEDCT_US|3-AMYL-1-HYDROXY-6,6,9-TRIMETHYL-6H-DIBENZO(B,D)PYRAN|CANNABINOL (SUBSTANCE)
C0006865|T053|96222005|SNOMEDCT_US|CANNABINOL [CHEMICAL/INGREDIENT]|CANNABINOL (SUBSTANCE)
C0006865|T053|96222005|SNOMEDCT_US|6,6,9-TRIMETHYL-3-PENTYL-6H-DIBENZO(B,D)PYRAN-1-OL|CANNABINOL (SUBSTANCE)
C0006865|T053|96222005|SNOMEDCT_US|CBN|CANNABINOL (SUBSTANCE)
C0006865|T053|96222005|SNOMEDCT_US|CANNABINOL |CANNABINOL (SUBSTANCE)
C0556618|T053|229001002|SNOMEDCT_US|CANNABIS GRASS - NON-PHARMACEUTICAL|CANNABIS GRASS - NON-PHARMACEUTICAL (SUBSTANCE)
C0556618|T053|229001002|SNOMEDCT_US|MARIJUANA GRASS|CANNABIS GRASS - NON-PHARMACEUTICAL (SUBSTANCE)
C0556618|T053|229001002|SNOMEDCT_US|MARIHUANA GRASS|CANNABIS GRASS - NON-PHARMACEUTICAL (SUBSTANCE)
C0556618|T053|229001002|SNOMEDCT_US|CANNABIS GRASS - NON-PHARMACEUTICAL |CANNABIS GRASS - NON-PHARMACEUTICAL (SUBSTANCE)
C0700258|T053|228998006|SNOMEDCT_US|MARIJUANA LEAF|CANNABIS LEAVES - NON-PHARMACEUTICAL (SUBSTANCE)
C0700258|T053|228998006|SNOMEDCT_US|CANNABIS LEAVES - NON-PHARMACEUTICAL|CANNABIS LEAVES - NON-PHARMACEUTICAL (SUBSTANCE)
C0700258|T053|228998006|SNOMEDCT_US|MARIHUANA LEAF|CANNABIS LEAVES - NON-PHARMACEUTICAL (SUBSTANCE)
C0700258|T053|228998006|SNOMEDCT_US|CANNABIS LEAVES - NON-PHARMACEUTICAL |CANNABIS LEAVES - NON-PHARMACEUTICAL (SUBSTANCE)
C0556617|T053|229000001|SNOMEDCT_US|CANNABIS OIL - NON-PHARMACEUTICAL|CANNABIS OIL - NON-PHARMACEUTICAL (SUBSTANCE)
C0556617|T053|229000001|SNOMEDCT_US|MARIJUANA OIL|CANNABIS OIL - NON-PHARMACEUTICAL (SUBSTANCE)
C0556617|T053|229000001|SNOMEDCT_US|MARIHUANA OIL|CANNABIS OIL - NON-PHARMACEUTICAL (SUBSTANCE)
C0556617|T053|229000001|SNOMEDCT_US|CANNABIS OIL - NON-PHARMACEUTICAL |CANNABIS OIL - NON-PHARMACEUTICAL (SUBSTANCE)
C0018613|T053|228999003|SNOMEDCT_US|HASHISH|CANNABIS RESIN - NON-PHARMACEUTICAL (SUBSTANCE)
C0018613|T053|228999003|SNOMEDCT_US|HASHISHS|CANNABIS RESIN - NON-PHARMACEUTICAL (SUBSTANCE)
C0018613|T053|228999003|SNOMEDCT_US|CANNABIS RESIN - NON-PHARMACEUTICAL|CANNABIS RESIN - NON-PHARMACEUTICAL (SUBSTANCE)
C0018613|T053|228999003|SNOMEDCT_US|MARIJUANA RESIN|CANNABIS RESIN - NON-PHARMACEUTICAL (SUBSTANCE)
C0018613|T053|228999003|SNOMEDCT_US|MARIHUANA RESIN|CANNABIS RESIN - NON-PHARMACEUTICAL (SUBSTANCE)
C0018613|T053|228999003|SNOMEDCT_US|CANNABIS RESIN - NON-PHARMACEUTICAL |CANNABIS RESIN - NON-PHARMACEUTICAL (SUBSTANCE)
C0005337|T053||SNOMEDCT_US|BHANGS
C0005337|T053||SNOMEDCT_US|BHANG
C0700268|T053|10083006|SNOMEDCT_US|MARIJUANA|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|CANNABIS SATIVA|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|CANNABIS SATIVA PLANT|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|SATIVAS, CANNABIS|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|CANNABIS SATIVAS|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|SATIVA, CANNABIS|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|CANNABIS SATIVA L.|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|CANNABIS|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|CANNABIS SATIVA WHOLE|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|MARIHUANA|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|INDIAN HEMP|CANNABIS SATIVA (ORGANISM)
C0700268|T053|10083006|SNOMEDCT_US|CANNABIS SATIVA |CANNABIS SATIVA (ORGANISM)
C0949248|T053||SNOMEDCT_US|INDICA, CANNABIS
C0949248|T053||SNOMEDCT_US|INDICAS, CANNABIS
C0949248|T053||SNOMEDCT_US|CANNABIS INDICAS
C0949248|T053||SNOMEDCT_US|CANNABIS INDICA
C0936079|T053|22924007|SNOMEDCT_US|CANNABIS|CANNABIS (ORGANISM)
C0936079|T053|22924007|SNOMEDCT_US|CANNABI|CANNABIS (ORGANISM)
C0936079|T053|22924007|SNOMEDCT_US|CANNABIS L., 1753|CANNABIS (ORGANISM)
C0936079|T053|22924007|SNOMEDCT_US|HEMP PLANT|CANNABIS (ORGANISM)
C0936079|T053|22924007|SNOMEDCT_US|CANNABIS |CANNABIS (ORGANISM)
C0936079|T053|22924007|SNOMEDCT_US|CANNABIS, NOS|CANNABIS (ORGANISM)
C0936079|T053|22924007|SNOMEDCT_US|HEMP (CANNABIS)|CANNABIS (ORGANISM)