C1531491|T053|413473000|SNOMEDCT_US|ALCOHOL CONSUMPTION COUNSELING|COUNSELING ABOUT ALCOHOL CONSUMPTION (PROCEDURE)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL ABUSE|ETHANOL ABUSE (FINDING)
C0560219|T053|160592001|SNOMEDCT_US|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS (FINDING)
0679277|T053||SNOMEDCT_US|ALCOHOL USE DISORDER CLASSIFICATION
C0687132|T053||SNOMEDCT_US|HEAVY DRINKING
C0740870|T053||SNOMEDCT_US|ALCOHOL USE FOR SLEEP
C1387092|T053||SNOMEDCT_US|ALCOHOL; HARMFUL USE
C2136082|T053||SNOMEDCT_US|ALCOHOL USE INTERFERING WITH SCHOOL
C2136085|T053||SNOMEDCT_US|ALCOHOL USE CAUSING HAZARD
C2215686|T053||SNOMEDCT_US|ALCOHOL USE DURING PREGNANCY
C2215687|T053||SNOMEDCT_US|ALCOHOL USE INTERFERING WITH WORK
C3837075|T053||SNOMEDCT_US|INTERVENTION FOR ALCOHOL USE
C3838370|T053||SNOMEDCT_US|BRIEF INTERVENTION FOR ALCOHOL USE
C0038586|T053||SNOMEDCT_US|SUBSTANCE USE DISORDERS
C0687725|T053|228281002|SNOMEDCT_US|ALCOHOLICS|PROBLEM DRINKER (LIFE STYLE)
C0337678|T053|86933000|SNOMEDCT_US|ALCOHOLIC BEVERAGE HEAVY DRINKER|HEAVY DRINKER (LIFE STYLE)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL ABUSE|ETHANOL ABUSE (FINDING)
C0001956|T053||SNOMEDCT_US|ALCOHOL USE DISORDER
C0001969|T053|231464007|SNOMEDCT_US|ALCOHOLIC INTOXICATION|INEBRIETY NOS (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLIC INTOXICATION, CHRONIC|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0683991|T053||SNOMEDCT_US|EX-ALCOHOLIC
C2366975|T053||SNOMEDCT_US|COUNSELING ABOUT RISK OF ALCOHOL CONSUMPTION
C2366975|T053||SNOMEDCT_US|COUNSELING ABOUT RISK OF ALCOHOL CONSUMPTION 
C2366975|T053||SNOMEDCT_US|EDUCATION PERFORMED ABOUT RISK OF ALCOHOL CONSUMPTION
C1531492|T053|413474006|SNOMEDCT_US|ALCOHOL COUNSELLING BY OTHER AGENCIES |COUNSELING ABOUT ALCOHOL BY OTHER AGENCIES (PROCEDURE)
C1531492|T053|413474006|SNOMEDCT_US|COUNSELLING ABOUT ALCOHOL BY OTHER AGENCIES|COUNSELING ABOUT ALCOHOL BY OTHER AGENCIES (PROCEDURE)
C1531492|T053|413474006|SNOMEDCT_US|COUNSELING ABOUT ALCOHOL BY OTHER AGENCIES |COUNSELING ABOUT ALCOHOL BY OTHER AGENCIES (PROCEDURE)
C1531492|T053|413474006|SNOMEDCT_US|ALCOHOL COUNSELING BY OTHER AGENCIES|COUNSELING ABOUT ALCOHOL BY OTHER AGENCIES (PROCEDURE)
C1531492|T053|413474006|SNOMEDCT_US|ALCOHOL COUNSELLING BY OTHER AGENCIES|COUNSELING ABOUT ALCOHOL BY OTHER AGENCIES (PROCEDURE)
C1531492|T053|413474006|SNOMEDCT_US|COUNSELING ABOUT ALCOHOL BY OTHER AGENCIES|COUNSELING ABOUT ALCOHOL BY OTHER AGENCIES (PROCEDURE)
C1531492|T053|413474006|SNOMEDCT_US|ALCOHOL COUNSELLING BY OTHER AGENCIES (REGIME/THERAPY)|COUNSELING ABOUT ALCOHOL BY OTHER AGENCIES (PROCEDURE)
C3494740|T053|429291000124102|SNOMEDCT_US|ALCOHOL BRIEF INTERVENTION|ALCOHOL BRIEF INTERVENTION (PROCEDURE)
C3494740|T053|429291000124102|SNOMEDCT_US|ALCOHOL BRIEF INTERVENTION |ALCOHOL BRIEF INTERVENTION (PROCEDURE)
C3165324|T053||SNOMEDCT_US|COUNSELING ABOUT ALCOHOL USE
C3165324|T053||SNOMEDCT_US|COUNSELLING ABOUT ALCOHOL USE
C0418859|T053|281078001|SNOMEDCT_US|ADVICE ON ALCOHOL CONSUMPTION|EDUCATION ABOUT ALCOHOL CONSUMPTION (PROCEDURE)
C0418859|T053|281078001|SNOMEDCT_US|ADVICE RELATING TO ALCOHOL CONSUMPTION|EDUCATION ABOUT ALCOHOL CONSUMPTION (PROCEDURE)
C0418859|T053|281078001|SNOMEDCT_US|EDUCATION ABOUT ALCOHOL CONSUMPTION|EDUCATION ABOUT ALCOHOL CONSUMPTION (PROCEDURE)
C0418859|T053|281078001|SNOMEDCT_US|EDUCATION ABOUT ALCOHOL CONSUMPTION |EDUCATION ABOUT ALCOHOL CONSUMPTION (PROCEDURE)
C0418859|T053|281078001|SNOMEDCT_US|ADVICE RELATING TO ALCOHOL CONSUMPTION |EDUCATION ABOUT ALCOHOL CONSUMPTION (PROCEDURE)
C0418859|T053|281078001|SNOMEDCT_US|ADVICE ON ALCOHOL CONSUMPTION |EDUCATION ABOUT ALCOHOL CONSUMPTION (PROCEDURE)
C0418859|T053|281078001|SNOMEDCT_US|ADVICE ON ALCOHOL CONSUMPTION (REGIME/THERAPY)|EDUCATION ABOUT ALCOHOL CONSUMPTION (PROCEDURE)
C0085762|T053|304606004|SNOMEDCT_US|ABUSE, ALCOHOL|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL ABUSE|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL ABUSE |ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ETHANOL ABUSE|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ETOH ABUSE|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL ABUSE-UNSPEC|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|RNDX ALCOHOL ABUSE|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|RNDX ALCOHOL ABUSE |ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL ABUSE, UNSPECIFIED|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL ABUSE, UNSPECIFIED DRINKING BEHAVIOR|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ETHANOL ABUSE |ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL ABUSE, UNSPECIFIED DRINKING BEHAVIOUR|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|AA - ALCOHOL ABUSE|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL ABUSE |ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ABUSE; ALCOHOL|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL; ABUSE|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|PROBLEM; ALCOHOL USE|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|ALCOHOL; USE, PROBLEM|ETHANOL ABUSE (FINDING)
C0085762|T053|304606004|SNOMEDCT_US|PROBLEM DRINKING|ETHANOL ABUSE (FINDING)
C2874370|T053||SNOMEDCT_US|ALCOHOL ABUSE, UNCOMPLICATED
C2874370|T053||SNOMEDCT_US|ALCOHOL ABUSE - UNCOMPLICATED
C2874370|T053||SNOMEDCT_US|ALCOHOL ABUSE - UNCOMPLICATED 
C2874371|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH INTOXICATION
C2874371|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH INTOXICATION, UNSPECIFIED
C2874371|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH INTOXICATION 
C2874377|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED MOOD DISORDER
C2874377|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2874377|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER
C2874377|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER, UNSP
C2874377|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED MOOD DISORDER 
C2874377|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER 
C2874381|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH OTHER ALCOHOL-INDUCED DISORDERS
C2874381|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH OTHER ALCOHOL-INDUCED DISORDER
C2874382|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH UNSPECIFIED ALCOHOL-INDUCED DISORDER
C1812624|T053||SNOMEDCT_US|ALCOHOL ABUSE, CONTINUOUS DRINKING BEHAVIOR
C1812624|T053||SNOMEDCT_US|CONTINUOUS ALCOHOL ABUSE 
C1812624|T053||SNOMEDCT_US|CONTINUOUS ALCOHOL ABUSE
C1812624|T053||SNOMEDCT_US|CONTINUOUS ETOH ABUSE
C1812624|T053||SNOMEDCT_US|CONTINUOUS ETHANOL ABUSE
C1812624|T053||SNOMEDCT_US|ALCOHOL ABUSE-CONTINUOUS
C1812624|T053||SNOMEDCT_US|ALCOHOL ABUSE, CONTINUOUS
C0154515|T053||SNOMEDCT_US|EPISODIC ALCOHOL ABUSE
C0154515|T053||SNOMEDCT_US|EPISODIC ALCOHOL ABUSE 
C0154515|T053||SNOMEDCT_US|ALCOHOL ABUSE, EPISODIC DRINKING BEHAVIOR
C0154515|T053||SNOMEDCT_US|EPISODIC ETHANOL ABUSE
C0154515|T053||SNOMEDCT_US|EPISODIC ETOH ABUSE
C0154515|T053||SNOMEDCT_US|ALCOHOL ABUSE-EPISODIC
C0154515|T053||SNOMEDCT_US|ALCOHOL ABUSE, EPISODIC
C0154515|T053||SNOMEDCT_US|ALCOHOL ABUSE, EPISODIC DRINKING BEHAVIOUR
C0154516|T053||SNOMEDCT_US|ALCOHOL ABUSE IN REMISSION
C0154516|T053||SNOMEDCT_US|ALCOHOL ABUSE IN REMISSION 
C0154516|T053||SNOMEDCT_US|ALCOHOL ABUSE, IN REMISSION
C0154516|T053||SNOMEDCT_US|ETOH ABUSE IN REMISSION
C0154516|T053||SNOMEDCT_US|ETHANOL ABUSE IN REMISSION
C0154516|T053||SNOMEDCT_US|ALCOHOL ABUSE-IN REMISS
C2874372|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH INTOXICATION, UNCOMPLICATED
C2874372|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH INTOXICATION - UNCOMPLICATED
C2874372|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH INTOXICATION - UNCOMPLICATED 
C2874373|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH INTOXICATION DELIRIUM
C2874373|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH INTOXICATION DELIRIUM 
C2874375|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS
C2874375|T053||SNOMEDCT_US|ALCOHOL ABUSE W ALCOH-INDUCE PSYCHOTIC DISORDER W DELUSIONS
C2874375|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS 
C2874376|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS
C2874376|T053||SNOMEDCT_US|ALCOHOL ABUSE W ALCOH-INDUCE PSYCHOTIC DISORDER W HALLUCIN
C2874376|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS 
C3509160|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED DISORDER 
C3509160|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED DISORDER
C2874378|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED ANXIETY DISORDER
C2874378|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED ANXIETY DISORDER 
C2874379|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED SEXUAL DYSFUNCTION
C2874379|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED SEXUAL DYSFUNCTION 
C2874380|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED SLEEP DISORDER
C2874380|T053||SNOMEDCT_US|ALCOHOL ABUSE WITH ALCOHOL-INDUCED SLEEP DISORDER 
C0338709|T053|191881009|SNOMEDCT_US|NONDEPENDENT ALCOHOL ABUSE|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|ALCOHOL ABUSE -NON DEP.|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED |NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|NONDEPENDENT ALCOHOL ABUSE NOS|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|NONDEPENDENT ALCOHOL ABUSE NOS |NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|NON-DEPENDENT ABUSE OF ALCOHOL|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|ALCOHOL ABUSE NONDEPENDENT|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|NONDEPENDENT ALCOHOL ABUSE |NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|NONDEPENDENT ABUSE OF ALCOHOL|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|NONDEPENDENT ALCOHOL ABUSE |NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|ALCOHOL; USE, HARMFUL (NON-DEPENDENT)|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0338709|T053|191881009|SNOMEDCT_US|USE; ALCOHOL, HARMFUL (NON-DEPENDENT)|NONDEPENDENT ALCOHOL ABUSE, UNSPECIFIED (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLISM|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|DIPSOMANIA|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOLIC INTOXICATION|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|INTOXICATION, CHRONIC ALCOHOLIC|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL, DEPENDENCE SYNDROME|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF ALCOHOL, DEPENDENCE SYNDROME|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL DEPENDENCE|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLIC INTOX CHRONIC|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ETOHISM|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ETOH DEPENDENCE|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ADDICTED TO ALCOHOL|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL DEPENDENCE |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLISM [DISEASE/FINDING]|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLIC INTOXICATION, CHRONIC|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ABUSE;ALCOHOL;CHRONIC|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ADDICTION;ALCOHOL|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|INTOXICATION;ALCOHOL;CHRONIC|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|DEPENDENCE;ALCOHOL|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLISM;CHRONIC|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLISM/ALCOHOL ABUSE|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ADDICTION, ALCOHOL|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|DEPENDENCE, ALCOHOL|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|UNSPECIFIED CHRONIC ALCOHOLISM |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL PROBLEM DRINKING|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|[X]MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF ALCOHOL: DEPENDENCE SYNDROME|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOLISM |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOLISM (& [DIPSOMANIA])|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: DEPENDENCE SYNDROME|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOLISM|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA])|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL DEPENDENCE SYNDROME NOS|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOLISM NOS |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|[X]ALCOHOL ADDICTION|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOLISM NOS|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|[X]DIPSOMANIA|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|(ALCOHOL DEPENDENCE SYNDROME [INCLUDING ALCOHOLISM]) OR (ALCOHOL PROBLEM DRINKING) |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL DEPENDENCE SYNDROME|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL DEPENDENCE SYNDROME NOS |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOLISM (& [DIPSOMANIA]) |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|(ALCOHOL DEPENDENCE SYNDROME [INCLUDING ALCOHOLISM]) OR (ALCOHOL PROBLEM DRINKING)|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|UNSPECIFIED CHRONIC ALCOHOLISM|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|DIPSOMANIA |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: DEPENDENCE SYNDROME |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|[X]CHRONIC ALCOHOLISM|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL ABUSE - PERSISTENT|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL ABUSE - PERSISTENT |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL ADDICTION|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL DEPENDENCY|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLISM AND ALCOHOL ABUSE|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL ABUSE CHRONIC|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL ABUSE, CONTINUOUS DRINKING BEHAVIOUR|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL ABUSE, CONTINUOUS DRINKING BEHAVIOR|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOL ABUSE|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|PERSISTENT ALCOHOL ABUSE|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL DEPENDENCE |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLISM |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|PERSISTENT ALCOHOL ABUSE |ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC; DRUNKENNESS|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|DEPENDENCE; ALCOHOL|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|DRUNKENNESS; CHRONIC|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ADDICTION; ALCOHOL|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL; ADDICTION|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOL; DEPENDENCE|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ALCOHOLISM, NOS|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOLISM [AMBIGUOUS]|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|DEPENDENCE; ETHYL ALCOHOL|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|ETHYL ALCOHOL; DEPENDENCE|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0001973|T053|154908007|SNOMEDCT_US|CHRONIC ALCOHOL INTOXICATION|ALCOHOL DEPENDENCE SYNDROME (& [DIPSOMANIA]) (DISORDER)
C0349269|T053|192481004|SNOMEDCT_US|ABUSE OF NON-DEPENDENCE-PRODUCING SUBSTANCES|[X]ABUSE OF NON-DEPENDENCE-PRODUCING SUBSTANCES
C0349269|T053|192481004|SNOMEDCT_US|[X]ABUSE OF NON-DEPENDENCE-PRODUCING SUBSTANCES|[X]ABUSE OF NON-DEPENDENCE-PRODUCING SUBSTANCES
C0349269|T053|192481004|SNOMEDCT_US|ABUSE OF NON-DEPENDENCE-PRODUCING SUBSTANCES |[X]ABUSE OF NON-DEPENDENCE-PRODUCING SUBSTANCES
C0582513|T053|304605000|SNOMEDCT_US|METHANOL ABUSE|METHANOL ABUSE (DISORDER)
C0582513|T053|304605000|SNOMEDCT_US|METHANOL ABUSE |METHANOL ABUSE (DISORDER)
C0582513|T053|304605000|SNOMEDCT_US|UNSPECIFIED PSYCH SUBSTANCE ABUSE METHANOL|METHANOL ABUSE (DISORDER)
C0582513|T053|304605000|SNOMEDCT_US|METHANOL ABUSE |METHANOL ABUSE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|MARCHIAFAVA-BIGNAMI DISEASE|MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|MARCHIAFAVA BIGNAMI DISEASE|MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|MARCHIAFAVA BIGNAMI SYNDROME|MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|MARCHIAFAVA-BIGNAMI DISEASE |MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|MARCHIAFAVA-BIGNAMI SYNDROME|MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|MARCHIAFAVA-BIGNAMI DISEASE [DISEASE/FINDING]|MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|MARCHIAFAVA DISEASE|MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|MARCHIAFAVA-BIGNAMI DISEASE |MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|CENTRAL DEMYELINATION OF CORPUS CALLOSUM |MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|MARCHIAFAVA|MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0238265|T053|386766007|SNOMEDCT_US|ENCEPHALOPATHY; DEMYELINATING CALLOSAL|MARCHIAFAVA-BIGNAMI DISEASE (DISORDER)
C0556330|T053|228310006|SNOMEDCT_US|DRINKS IN MORNING TO GET RID OF HANGOVER|DRINKS IN MORNING TO GET RID OF HANGOVER (FINDING)
C0556330|T053|228310006|SNOMEDCT_US|DRINKS IN MORNING TO GET RID OF HANGOVER |DRINKS IN MORNING TO GET RID OF HANGOVER (FINDING)
C0556343|T053|228323004|SNOMEDCT_US|DRINKING BOUT|DRINKING BOUT (FINDING)
C0556343|T053|228323004|SNOMEDCT_US|DRINKING BOUT |DRINKING BOUT (FINDING)
C0556383|T053|228363003|SNOMEDCT_US|FEELS DRINKING IS OUT OF CONTROL|FEELS DRINKING IS OUT OF CONTROL (FINDING)
C0556383|T053|228363003|SNOMEDCT_US|FEELS DRINKING IS OUT OF CONTROL |FEELS DRINKING IS OUT OF CONTROL (FINDING)
C0556364|T053|228344004|SNOMEDCT_US|UNABLE TO STOP DRINKING BEFORE INTOXICATION|UNABLE TO STOP DRINKING BEFORE INTOXICATION (FINDING)
C0556364|T053|228344004|SNOMEDCT_US|UNABLE TO STOP DRINKING BEFORE INTOXICATION |UNABLE TO STOP DRINKING BEFORE INTOXICATION (FINDING)
C0560219|T053|160592001|SNOMEDCT_US|EXCESSIVE ALCOHOL USE|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS (FINDING)
C0560219|T053|160592001|SNOMEDCT_US|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS (FINDING)
C0560219|T053|160592001|SNOMEDCT_US|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS |ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS (FINDING)
C0560219|T053|160592001|SNOMEDCT_US|EXCESSIVE ALCOHOL CONSUMPTION|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS (FINDING)
C0560219|T053|160592001|SNOMEDCT_US|XS - EXCESSIVE ALCOHOL CONSUMPTION|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS (FINDING)
C0560219|T053|160592001|SNOMEDCT_US|XS - EXCESSIVE ETHANOL CONSUMPTION|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS (FINDING)
C0560219|T053|160592001|SNOMEDCT_US|EXCESSIVE ETHANOL CONSUMPTION|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS (FINDING)
C0560219|T053|160592001|SNOMEDCT_US|EXCESSIVE DRINKING OF ALCOHOL NOS|ALCOHOL INTAKE ABOVE RECOMMENDED SENSIBLE LIMITS (FINDING)
C0556337|T053|228317009|SNOMEDCT_US|ALCOHOLIC BINGES EXCEEDING SAFE AMOUNTS|ALCOHOLIC BINGES EXCEEDING SAFE AMOUNTS (FINDING)
C0556337|T053|228317009|SNOMEDCT_US|ALCOHOLIC BINGES EXCEEDING SAFE AMOUNTS |ALCOHOLIC BINGES EXCEEDING SAFE AMOUNTS (FINDING)
C0556336|T053|228316000|SNOMEDCT_US|ALCOHOLIC BINGES EXCEEDING SENSIBLE AMOUNTS|ALCOHOLIC BINGES EXCEEDING SENSIBLE AMOUNTS (FINDING)
C0556336|T053|228316000|SNOMEDCT_US|ALCOHOLIC BINGES EXCEEDING SENSIBLE AMOUNTS |ALCOHOLIC BINGES EXCEEDING SENSIBLE AMOUNTS (FINDING)
C0556346|T053|228326007|SNOMEDCT_US|BINGE DRINKING|DRINKING BINGE (FINDING)
C0556346|T053|228326007|SNOMEDCT_US|DRINKING, BINGE|DRINKING BINGE (FINDING)
C0556346|T053|228326007|SNOMEDCT_US|BINGE DRINKING [DISEASE/FINDING]|DRINKING BINGE (FINDING)
C0556346|T053|228326007|SNOMEDCT_US|ALCOHOL BINGE|DRINKING BINGE (FINDING)
C0556346|T053|228326007|SNOMEDCT_US|DRINKING BINGE|DRINKING BINGE (FINDING)
C0556346|T053|228326007|SNOMEDCT_US|DRINKING BINGE |DRINKING BINGE (FINDING)
C0556335|T053|228315001|SNOMEDCT_US|BINGE DRINKER|BINGE DRINKER (FINDING)
C0556335|T053|228315001|SNOMEDCT_US|BOUT DRINKER|BINGE DRINKER (FINDING)
C0556335|T053|228315001|SNOMEDCT_US|EPISODIC DRINKER|BINGE DRINKER (FINDING)
C0556335|T053|228315001|SNOMEDCT_US|BINGE DRINKER |BINGE DRINKER (FINDING)
C0556363|T053|228343005|SNOMEDCT_US|UNABLE TO CONTROL SPONTANEOUS DRINKING BOUTS|UNABLE TO CONTROL SPONTANEOUS DRINKING BOUTS (FINDING)
C0556363|T053|228343005|SNOMEDCT_US|UNABLE TO CONTROL SPONTANEOUS DRINKING BOUTS |UNABLE TO CONTROL SPONTANEOUS DRINKING BOUTS (FINDING)
C2106524|T053||SNOMEDCT_US|COMBINED DRUG AND ALCOHOL ABUSE 
C2106524|T053||SNOMEDCT_US|COMBINED DRUG AND ALCOHOL ABUSE
C2181572|T053||SNOMEDCT_US|A BREATHALYZER FOR BLOOD ALCOHOL CONTENT SHOWED AN EXCESSIVE BLOOD ALCOHOL LEVEL
C2181572|T053||SNOMEDCT_US|BREATHALYZER FOR BLOOD ALCOHOL CONTENT EXCESSIVE BLOOD ALCOHOL LEVEL
C2181572|T053||SNOMEDCT_US|BREATHALYZER FOR BLOOD ALCOHOL CONTENT: EXCESSIVE BLOOD ALCOHOL LEVEL 
C2181572|T053||SNOMEDCT_US|BREATHALYZER FOR BLOOD ALCOHOL CONTENT: EXCESSIVE BLOOD ALCOHOL LEVEL
C1387092|T053||SNOMEDCT_US|HARMFUL; USE, ALCOHOL
C1387092|T053||SNOMEDCT_US|ALCOHOL; HARMFUL USE
C2136086|T053||SNOMEDCT_US|ALCOHOL USE CAUSING HAZARD AT WORK 
C2136086|T053||SNOMEDCT_US|ALCOHOL USE CAUSING HAZARD AT WORK
C2136087|T053||SNOMEDCT_US|ALCOHOL USE CAUSING HAZARD WHILE DRIVING
C2136087|T053||SNOMEDCT_US|ALCOHOL USE CAUSING HAZARD WHILE DRIVING 
C1959897|T053|427013000|SNOMEDCT_US|ALCOHOL CONSUMPTION DURING PREGNANCY|ALCOHOL CONSUMPTION DURING PREGNANCY (FINDING)
C1959897|T053|427013000|SNOMEDCT_US|ALCOHOL CONSUMPTION DURING PREGNANCY |ALCOHOL CONSUMPTION DURING PREGNANCY (FINDING)
C3838370|T053||SNOMEDCT_US|BRIEF INTERVENTION FOR ALCOHOL USE 
C3838370|T053||SNOMEDCT_US|BRIEF INTERVENTION FOR ALCOHOL USE
C3838370|T053||SNOMEDCT_US|INTERVENTION FOR ALCOHOL USE BRIEF
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL RELATED DISORDERS|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL-RELATED DISORDER|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL-RELATED DISORDERS|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|DISORDER, ALCOHOL-RELATED|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|DISORDERS, ALCOHOL-RELATED|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL RELATED DIS|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL-RELATED DISORDERS [DISEASE/FINDING]|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL-RELATED DISORDERS |ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL DISORDERS|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER |ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER, NOS|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL-RELATED DISORDER, NOS|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0236664|T053|29212009|SNOMEDCT_US|ALCOHOL-RELATED DISORDER NOS|ALCOHOL-INDUCED ORGANIC MENTAL DISORDER (DISORDER)
C0687725|T053|228281002|SNOMEDCT_US|ALCOHOLIC|PROBLEM DRINKER (LIFE STYLE)
C0687725|T053|228281002|SNOMEDCT_US|ALCOHOLICS|PROBLEM DRINKER (LIFE STYLE)
C0687725|T053|228281002|SNOMEDCT_US|BOOZER|PROBLEM DRINKER (LIFE STYLE)
C0687725|T053|228281002|SNOMEDCT_US|DEPENDENT DRINKER|PROBLEM DRINKER (LIFE STYLE)
C0687725|T053|228281002|SNOMEDCT_US|PROBLEM DRINKER|PROBLEM DRINKER (LIFE STYLE)
C0687725|T053|228281002|SNOMEDCT_US|PROBLEM DRINKER |PROBLEM DRINKER (LIFE STYLE)
C0687725|T053|228281002|SNOMEDCT_US|PROBLEM DRINKER |PROBLEM DRINKER (LIFE STYLE)
C0037263|T053||SNOMEDCT_US|ALCOHOLIC, SKID ROW
C0037263|T053||SNOMEDCT_US|ALCOHOLICS, SKID ROW
C0037263|T053||SNOMEDCT_US|SKID ROW ALCOHOLICS
C0037263|T053||SNOMEDCT_US|SKID ROW ALCOHOLIC
C2030272|T053||SNOMEDCT_US|HEAVY ALCOHOL CONSUMPTION
C2030272|T053||SNOMEDCT_US|HEAVY ALCOHOL CONSUMPTION 
C0337678|T053|86933000|SNOMEDCT_US|ALCOHOLIC BEVERAGE HEAVY DRINKER|HEAVY DRINKER (LIFE STYLE)
C0337678|T053|86933000|SNOMEDCT_US|HEAVY DRINKER |HEAVY DRINKER (LIFE STYLE)
C0337678|T053|86933000|SNOMEDCT_US|HEAVY DRINKER|HEAVY DRINKER (LIFE STYLE)
C0337678|T053|86933000|SNOMEDCT_US|DRINKS HEAVILY|HEAVY DRINKER (LIFE STYLE)
C0337678|T053|86933000|SNOMEDCT_US|HEAVY DRINKER |HEAVY DRINKER (LIFE STYLE)
C0425319|T053|160577002|SNOMEDCT_US|HEAVY DRINKER - 7-9U/DAY|HEAVY DRINKER - 7-9U/DAY (LIFE STYLE)
C0425319|T053|160577002|SNOMEDCT_US|HEAVY DRINKER - 7-9U/DAY |HEAVY DRINKER - 7-9U/DAY (LIFE STYLE)
C0425319|T053|160577002|SNOMEDCT_US|HEAVY DRINKER - 7-9U/DAY |HEAVY DRINKER - 7-9U/DAY (LIFE STYLE)
C0496556|T053||SNOMEDCT_US|MILD ALCOHOL INTOXICATION
C0496557|T053||SNOMEDCT_US|MODERATE ALCOHOL INTOXICATION
C0496558|T053||SNOMEDCT_US|SEVERE ALCOHOL INTOXICATION
C0496559|T053||SNOMEDCT_US|VERY SEVERE ALCOHOL INTOXICATION
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|AC ALCOHOL INTOX-UNSPEC|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE DRUNKENNESS (IN ALCOHOLISM)|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM, UNSPECIFIED|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM, UNSPECIFIED DRINKING BEHAVIOR|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM |ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM NOS|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM NOS |ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOL INTOXICATION IN ALCOHOLISM|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ALCOHOL INTOXICATION - ACUTE IN ALCOHOLISM|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOL INTOXICATION IN ALCOHOLISM |ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM, UNSPECIFIED DRINKING BEHAVIOUR|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ACUTE ALCOHOLIC INTOXICATION|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM |ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|DRUNKENNESS; ACUTE IN ALCOHOLISM|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE; DRUNKENNESS IN ALCOHOLISM|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED DRINKING BEHAVIOR|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0812429|T053|191803009|SNOMEDCT_US|ACUTE DRUNKENNESS IN ALCOHOLISM|ACUTE ALCOHOLIC INTOXICATION, UNSPECIFIED, IN ALCOHOLISM (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|ACUTE ALCOHOLIC INTOXICATION|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL, ACUTE INTOXICATION|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF ALCOHOL, ACUTE INTOXICATION|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|INTOXICATION;ALCOHOL;ACUTE|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|[X]MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION |[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|ALCOHOL INTOXICATION ACUTE|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|ALCOHOL INTOXICATION, ACUTE|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0394996|T053|192207001|SNOMEDCT_US|ACUTE ALCOHOL INTOXICATION|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: ACUTE INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|IDIOSYNCRATIC ALCOHOL INTOXICATION|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|ALCOHOL IDIOSYNCRATIC INTOXICATION |IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|ALCOHOL IDIOSYNCRATIC INTOXICATION|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|PATHOLOGIC ALCOHOL INTOX|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|ALCOHOL INTOXICATION - PATHOLOGICAL |IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|ALCOHOL INTOXICATION - PATHOLOGICAL|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|PATHOLOGICAL ALCOHOL INTOXICATION|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|PATHOLOGICAL DRUNKENNESS|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|PATHOLOGICAL INTOXICATION|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|EXTREME SENSITIVITY TO ALCOHOL SYNDROME|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|IDIOSYNCRATIC INTOXICATION|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|DRUNKENNESS - PATHOLOGICAL|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|IDIOSYNCRATIC INTOXICATION |IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|PATHOLOGICAL ALCOHOL INTOXICATION |IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|DRUNKENNESS; PATHOLOGICAL|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|INTOXICATION; ALCOHOL, IDIOSYNCRATIC|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|INTOXICATION; ALCOHOL, PATHOLOGICAL|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|INTOXICATION; PATHOLOGIC|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|PATHOLOGIC; INTOXICATION|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|PATHOLOGICAL; DRUNKENNESS|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|ALCOHOL; INTOXICATION, IDIOSYNCRATIC|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|ALCOHOL; INTOXICATION, PATHOLOGICAL|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|PATHOLOGIC ALCOHOL INTOXICATION|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001950|T053|21000000|SNOMEDCT_US|PATHOLOGIC DRUNKENNESS|IDIOSYNCRATIC INTOXICATION (DISORDER)
C0001969|T053|231464007|SNOMEDCT_US|ABUSE;ALCOHOL;ACUTE|INEBRIETY NOS (DISORDER)
C0001969|T053|231464007|SNOMEDCT_US|ADDICTION;ALCOHOL;ACUTE|INEBRIETY NOS (DISORDER)
C2104528|T053||SNOMEDCT_US|CONTINUOUS ALCOHOL INTOXICATION 
C2104528|T053||SNOMEDCT_US|CONTINUOUS ALCOHOL INTOXICATION
C2104529|T053||SNOMEDCT_US|EPISODIC ALCOHOL INTOXICATION
C2104529|T053||SNOMEDCT_US|EPISODIC ALCOHOL INTOXICATION 
C2104530|T053||SNOMEDCT_US|ALCOHOL INTOXICATION IN REMISSION 
C2104530|T053||SNOMEDCT_US|ALCOHOL INTOXICATION IN REMISSION
C3650362|T053||SNOMEDCT_US|ALCOHOL INTOXICATION - UNCOMPLICATED
C0236654|T053|18653004|SNOMEDCT_US|ALCOHOL INTOXICATION DELIRIUM|ALCOHOL INTOXICATION DELIRIUM (DISORDER)
C0236654|T053|18653004|SNOMEDCT_US|ALCOHOL INTOXICATION DELIRIUM |ALCOHOL INTOXICATION DELIRIUM (DISORDER)
C0236654|T053|18653004|SNOMEDCT_US|ALCOHOL INTOXICATION DELIRIUM |ALCOHOL INTOXICATION DELIRIUM (DISORDER)
C0236654|T053|18653004|SNOMEDCT_US|INTOXICATION; ALCOHOL, DELIRIUM|ALCOHOL INTOXICATION DELIRIUM (DISORDER)
C0236654|T053|18653004|SNOMEDCT_US|ALCOHOL; DELIRIUM, INTOXICATION|ALCOHOL INTOXICATION DELIRIUM (DISORDER)
C0236654|T053|18653004|SNOMEDCT_US|ALCOHOL; INTOXICATION, DELIRIUM|ALCOHOL INTOXICATION DELIRIUM (DISORDER)
C0033936|T053|192212000|SNOMEDCT_US|PSYCHOSES, ALCOHOLIC|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOLIC PSYCHOSES|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOLIC PSYCHOSIS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL, PSYCHOTIC DISORDER|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF ALCOHOL, PSYCHOTIC DISORDER|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOL-INDUCED PSYCHOTIC DISORDER|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOL-INDUCED PSYCHOTIC DISORDER |[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOL MENTAL DISOR NOS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|PSYCHOSES, ALCOHOLIC [DISEASE/FINDING]|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|PSYCHOSIS;ALCOHOLIC|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOL INDUCED PSYCHOSIS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|[X]ALCOHOLIC PSYCHOSIS NOS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOLIC PSYCHOSES |[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: PSYCHOTIC DISORDER|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|[X]MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF ALCOHOL: PSYCHOTIC DISORDER|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOLIC PSYCHOSIS NOS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOLIC PSYCHOSIS NOS |[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: PSYCHOTIC DISORDER |[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOLIC PSYCHOSIS, UNSPECIFIED|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|UNSPECIFIED ALCOHOLIC PSYCHOSIS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|PSYCHOSIS ALCOHOLIC|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOL-INDUCED PSYCHOSIS |[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOL-INDUCED PSYCHOSIS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|DISORDER; PSYCHOTIC, ALCOHOL (DUE TO), ALCOHOLIC|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOLISM; PSYCHOSIS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|PSYCHOSIS; ALCOHOLIC|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|PSYCHOTIC; DISORDER, ALCOHOL (DUE TO), ALCOHOLIC|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOL-INDUCED PSYCHOSIS, NOS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOLIC PSYCHOSIS, NOS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|ALCOHOLISM WITH PSYCHOSIS|[X]ALCOHOLIC PSYCHOSIS NOS
C0033936|T053|192212000|SNOMEDCT_US|UNSPECIFIED ALCOHOL-INDUCED MENTAL DISORDERS|[X]ALCOHOLIC PSYCHOSIS NOS
C0392621|T053|212809004|SNOMEDCT_US|METHANOL POISONING|METHYL ALCOHOL POISONING
C0392621|T053|212809004|SNOMEDCT_US|POISONING BY METHYL ALCOHOL|METHYL ALCOHOL POISONING
C0392621|T053|212809004|SNOMEDCT_US|POISONING BY METHYL ALCOHOL |METHYL ALCOHOL POISONING
C0392621|T053|212809004|SNOMEDCT_US|METHYL ALCOHOL POISONING|METHYL ALCOHOL POISONING
C0556374|T053|228354000|SNOMEDCT_US|ALCOHOL INFLUENCED DRIVING|DRUNK DRIVING (FINDING)
C0556374|T053|228354000|SNOMEDCT_US|DRUNK DRIVING|DRUNK DRIVING (FINDING)
C0556374|T053|228354000|SNOMEDCT_US|DRIVING WHILE INTOXICATED|DRUNK DRIVING (FINDING)
C0556374|T053|228354000|SNOMEDCT_US|DRINK DRIVING|DRUNK DRIVING (FINDING)
C0556374|T053|228354000|SNOMEDCT_US|DRUNK DRIVING |DRUNK DRIVING (FINDING)
C0556374|T053|228354000|SNOMEDCT_US|DRINK DRIVING |DRUNK DRIVING (FINDING)
C0338785|T053|191811004|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH CONTINUOUS DRINKING BEHAVIOR|CONTINUOUS CHRONIC ALCOHOLISM (DISORDER)
C0338785|T053|191811004|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH CONTINUOUS DRINKING BEHAVIOR |CONTINUOUS CHRONIC ALCOHOLISM (DISORDER)
C0338785|T053|191811004|SNOMEDCT_US|CONTINUOUS CHRONIC ALCOHOLISM|CONTINUOUS CHRONIC ALCOHOLISM (DISORDER)
C0338785|T053|191811004|SNOMEDCT_US|CONTINUOUS CHRONIC ALCOHOLISM |CONTINUOUS CHRONIC ALCOHOLISM (DISORDER)
C2874383|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE, UNCOMPLICATED
C2874383|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE UNCOMPLICATED 
C2874383|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE UNCOMPLICATED
C2197979|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE IN REMISSION 
C2197979|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE IN REMISSION
C2197979|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE, IN REMISSION
C2874387|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH INTOXICATION
C2874387|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH INTOXICATION, UNSPECIFIED
C2874387|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH INTOXICATION 
C2874392|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL
C2874392|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL, UNSPECIFIED
C2874392|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL 
C2874393|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED MOOD DISORDER
C2874393|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED MOOD DISORDER 
C2874397|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER
C2874397|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER, UNSPECIFIED
C2874397|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE W ALCOH-INDUCE PSYCHOTIC DISORDER, UNSP
C2874397|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER 
C2874398|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PERSISTING AMNESTIC DISORDER
C2874398|T053||SNOMEDCT_US|ALCOHOL DEPEND W ALCOH-INDUCE PERSISTING AMNESTIC DISORDER
C2874399|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PERSISTING DEMENTIA
C2874403|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH OTHER ALCOHOL-INDUCED DISORDER
C2874403|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH OTHER ALCOHOL-INDUCED DISORDERS
C2874404|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH UNSPECIFIED ALCOHOL-INDUCED DISORDER
C2048484|T053||SNOMEDCT_US|INABILITY TO QUIT DRINKING ALCOHOL 
C2048484|T053||SNOMEDCT_US|INABILITY TO QUIT DRINKING ALCOHOL
C0338784|T053|191812006|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH EPISODIC DRINKING BEHAVIOR|EPISODIC CHRONIC ALCOHOLISM (DISORDER)
C0338784|T053|191812006|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH EPISODIC DRINKING BEHAVIOR |EPISODIC CHRONIC ALCOHOLISM (DISORDER)
C0338784|T053|191812006|SNOMEDCT_US|EPISODIC CHRONIC ALCOHOLISM|EPISODIC CHRONIC ALCOHOLISM (DISORDER)
C0338784|T053|191812006|SNOMEDCT_US|EPISODIC CHRONIC ALCOHOLISM |EPISODIC CHRONIC ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOL-INDUCED PERSISTENT DEMENTIA |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOL-INDUCED PERSISTENT DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH DEMENTIA |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOL INDUCED PERSISTING DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOL PERSIST DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|DEMENTIA;ALCOHOLIC|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOLIC DEMENTIA NOS|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|[X]ALCOHOLIC DEMENTIA NOS|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|[X]CHRONIC ALCOHOLIC BRAIN SYNDROME|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOLIC DEMENTIA NOS |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|CHRONIC ORGANIC MENTAL DISORDER ALCOHOLIC BRAIN SYNDROME|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|CHRONIC ALCOHOLIC BRAIN SYNDROME|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|CHRONIC ALCOHOLIC BRAIN SYNDROME |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|DEMENTIA ASSOCIATED WITH ALCOHOLISM|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOL-INDUCED PERSISTING DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOLIC DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|CHRONIC ALCOHOLIC BRAIN SYNDROME |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|DEMENTIA ASSOCIATED WITH ALCOHOLISM |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|BRAIN; SYNDROME, ALCOHOLIC (CHRONIC)|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|DEMENTIA; ALCOHOLIC|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|DEMENTIA; ALCOHOL|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOL; DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|SYNDROME; BRAIN, ALCOHOLIC (CHRONIC)|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T053|281004|SNOMEDCT_US|ALCOHOLISM ASSOCIATED WITH DEMENTIA NOS|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C2874389|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL, UNCOMPLICATED
C2874389|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL - UNCOMPLICATED 
C2874389|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL - UNCOMPLICATED
C2874390|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL DELIRIUM
C2874390|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL DELIRIUM 
C2874391|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL WITH PERCEPTUAL DISTURBANCE
C2874391|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE W WITHDRAWAL WITH PERCEPTUAL DISTURBANCE
C2874391|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH WITHDRAWAL WITH PERCEPTUAL DISTURBANCE 
C2874395|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS
C2874395|T053||SNOMEDCT_US|ALCOHOL DEPEND W ALCOH-INDUCE PSYCHOTIC DISORDER W DELUSIONS
C2874395|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH DELUSIONS 
C2874396|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS
C2874396|T053||SNOMEDCT_US|ALCOHOL DEPEND W ALCOH-INDUCE PSYCHOTIC DISORDER W HALLUCIN
C2874396|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PSYCHOTIC DISORDER WITH HALLUCINATIONS 
C3509162|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PERSISTNG AMNESTIC DISORDER
C3509162|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PERSISTNG AMNESTIC DISORDER 
C3509163|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PERSISTNG DEMENTIA
C3509163|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED PERSISTNG DEMENTIA 
C3509161|T053|288031000119105|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED DISORDER|ALCOHOL INDUCED DISORDER CO-OCCURRENT AND DUE TO ALCOHOL DEPENDENCE (DISORDER)
C3509161|T053|288031000119105|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED DISORDER |ALCOHOL INDUCED DISORDER CO-OCCURRENT AND DUE TO ALCOHOL DEPENDENCE (DISORDER)
C2874400|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED ANXIETY DISORDER
C2874400|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED ANXIETY DISORDER 
C2874401|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED SEXUAL DYSFUNCTION
C2874401|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED SEXUAL DYSFUNCTION 
C2874402|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED SLEEP DISORDER
C2874402|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH ALCOHOL-INDUCED SLEEP DISORDER 
C2874386|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH INTOXICATION DELIRIUM
C2874386|T053||SNOMEDCT_US|ALCOHOL DEPENDENCE WITH INTOXICATION DELIRIUM 
C0023896|T053|41309000|SNOMEDCT_US|LIVER DISEASE, ALCOHOLIC|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|LIVER DISEASES, ALCOHOLIC|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALCOHOLIC LIVER DISEASE|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALCOHOLIC LIVER DISEASE, UNSPECIFIED|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|LIVER DIS ALCOHOLIC|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALCOHOLIC LIVER DIS|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALCOHOL INDUCED LIVER DISORDER|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|LIVER DISEASES, ALCOHOLIC [DISEASE/FINDING]|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALCOHOLIC LIVER DISEASES|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALCOHOLIC LIVER DISEASE |ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALCOHOLIC LIVER DISEASE NOS|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|HEPATOPATHY ALCOHOLIC|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALD - ALCOHOLIC LIVER DISEASE|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|DISEASE (OR DISORDER); LIVER, ALCOHOLIC|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|LIVER; ALCOHOL|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|LIVER; DISEASE, ALCOHOLIC|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALCOHOL; LIVER|ALD - ALCOHOLIC LIVER DISEASE
C0023896|T053|41309000|SNOMEDCT_US|ALCOHOLIC LIVER DISEASE, NOS|ALD - ALCOHOLIC LIVER DISEASE
C0272023|T053|86325007|SNOMEDCT_US|NON MEGALOBLASTIC ANEMIA DUE TO ALCOHOLISM|NON MEGALOBLASTIC ANEMIA DUE TO ALCOHOLISM (DISORDER)
C0272023|T053|86325007|SNOMEDCT_US|NON MEGALOBLASTIC ANAEMIA DUE TO ALCOHOLISM|NON MEGALOBLASTIC ANEMIA DUE TO ALCOHOLISM (DISORDER)
C0272023|T053|86325007|SNOMEDCT_US|NON MEGALOBLASTIC ANEMIA DUE TO ALCOHOLISM |NON MEGALOBLASTIC ANEMIA DUE TO ALCOHOLISM (DISORDER)
C3839769|T053|10755041000119100|SNOMEDCT_US|ALCOHOL DEPENDENCE IN CHILDBIRTH |ALCOHOL DEPENDENCE IN CHILDBIRTH (DISORDER)
C3839769|T053|10755041000119100|SNOMEDCT_US|ALCOHOL DEPENDENCE IN CHILDBIRTH|ALCOHOL DEPENDENCE IN CHILDBIRTH (DISORDER)
C1411379|T053|10741871000119101|SNOMEDCT_US|ALCOHOL DEPENDENCE IN PREGNANCY |ALCOHOL DEPENDENCE IN PREGNANCY (DISORDER)
C1411379|T053|10741871000119101|SNOMEDCT_US|ALCOHOL DEPENDENCE IN PREGNANCY|ALCOHOL DEPENDENCE IN PREGNANCY (DISORDER)
C1411379|T053|10741871000119101|SNOMEDCT_US|PREGNANCY; ALCOHOL DEPENDENCE|ALCOHOL DEPENDENCE IN PREGNANCY (DISORDER)
C4075901|T053|713583005|SNOMEDCT_US|MILD ALCOHOL DEPENDENCE |MILD ALCOHOL DEPENDENCE (DISORDER)
C4075901|T053|713583005|SNOMEDCT_US|MILD ALCOHOL DEPENDENCE|MILD ALCOHOL DEPENDENCE (DISORDER)
C4075720|T053|713862009|SNOMEDCT_US|SEVERE ALCOHOL DEPENDENCE |SEVERE ALCOHOL DEPENDENCE (DISORDER)
C4075720|T053|713862009|SNOMEDCT_US|SEVERE ALCOHOL DEPENDENCE|SEVERE ALCOHOL DEPENDENCE (DISORDER)
C4075073|T053|714829008|SNOMEDCT_US|MODERATE ALCOHOL DEPENDENCE |MODERATE ALCOHOL DEPENDENCE (DISORDER)
C4075073|T053|714829008|SNOMEDCT_US|MODERATE ALCOHOL DEPENDENCE|MODERATE ALCOHOL DEPENDENCE (DISORDER)
C4076151|T053|97571000119109|SNOMEDCT_US|THROMBOCYTOPAENIA CO-OCCURRENT AND DUE TO ALCOHOLISM|THROMBOCYTOPENIA CO-OCCURRENT AND DUE TO ALCOHOLISM (DISORDER)
C4076151|T053|97571000119109|SNOMEDCT_US|THROMBOCYTOPENIA CO-OCCURRENT AND DUE TO ALCOHOLISM|THROMBOCYTOPENIA CO-OCCURRENT AND DUE TO ALCOHOLISM (DISORDER)
C4076151|T053|97571000119109|SNOMEDCT_US|THROMBOCYTOPENIA CO-OCCURRENT AND DUE TO ALCOHOLISM |THROMBOCYTOPENIA CO-OCCURRENT AND DUE TO ALCOHOLISM (DISORDER)
C0338783|T053|191813001|SNOMEDCT_US|CHRONIC ALCOHOLISM IN REMISSION|CHRONIC ALCOHOLISM IN REMISSION (DISORDER)
C0338783|T053|191813001|SNOMEDCT_US|CHRONIC ALCOHOLISM IN REMISSION |CHRONIC ALCOHOLISM IN REMISSION (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOLIC LIVER DAMAGE|ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOLIC LIVER DAMAGE |ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOL LIVER DAMAGE NOS|ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOLIC LIVER DAMAGE UNSPECIFIED |ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOLIC LIVER DAMAGE NOS |ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOLIC LIVER DAMAGE NOS|ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOLIC LIVER DAMAGE UNSPECIFIED|ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOLIC LIVER DAMAGE, UNSPECIFIED|ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOLIC LIVER DAMAGE |ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|DAMAGE; LIVER, ALCOHOLIC|ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|LIVER; DAMAGE, ALCOHOLIC|ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1442981|T053|197282000|SNOMEDCT_US|ALCOHOLIC LIVER DAMAGE, NOS|ALCOHOLIC LIVER DAMAGE UNSPECIFIED (DISORDER)
C1386568|T053||SNOMEDCT_US|DEPENDENCE; METHYLATED SPIRIT
C1386568|T053||SNOMEDCT_US|METHYLATED SPIRIT; DEPENDENCE
C1386585|T053||SNOMEDCT_US|DEPENDENCE; METHYL ALCOHOL
C1386585|T053||SNOMEDCT_US|METHYL ALCOHOL; DEPENDENCE
C1387095|T053||SNOMEDCT_US|POISONING; ALCOHOL, WITH DEPENDENCE
C1387095|T053||SNOMEDCT_US|ALCOHOL; POISONING, WITH DEPENDENCE
C1395804|T053||SNOMEDCT_US|DRINKING; EXCESS, HABIT (CONTINUAL)
C1395804|T053||SNOMEDCT_US|DRINKING; EXCESSIVE, HABIT (CONTINUAL)
C1395804|T053||SNOMEDCT_US|EXCESS; DRINKING, HABIT (CONTINUAL)
C1395804|T053||SNOMEDCT_US|EXCESSIVE; DRINKING, HABIT (CONTINUAL)
C1395805|T053||SNOMEDCT_US|DRINKING; HABITUAL
C1395805|T053||SNOMEDCT_US|HABITUAL; DRINKING
C0014984|T053||SNOMEDCT_US|ETHANOLISM
C0392620|T053|82782008|SNOMEDCT_US|ALCOHOL POISONING|ETHANOL POISONING
C0392620|T053|82782008|SNOMEDCT_US|POISONING BY ETHYL ALCOHOL |ETHANOL POISONING
C0392620|T053|82782008|SNOMEDCT_US|POISONING BY ALCOHOL|ETHANOL POISONING
C0392620|T053|82782008|SNOMEDCT_US|POISONING BY ALCOHOL |ETHANOL POISONING
C0392620|T053|82782008|SNOMEDCT_US|POISONING BY ETHYL ALCOHOL|ETHANOL POISONING
C0392620|T053|82782008|SNOMEDCT_US|ETHANOL POISONING|ETHANOL POISONING
C0392620|T053|82782008|SNOMEDCT_US|ETHYL ALCOHOL POISONING|ETHANOL POISONING
C0392620|T053|82782008|SNOMEDCT_US|ETHYLISM|ETHANOL POISONING
C0392620|T053|82782008|SNOMEDCT_US|POISONING; ALCOHOL|ETHANOL POISONING
C0392620|T053|82782008|SNOMEDCT_US|ALCOHOL; POISONING|ETHANOL POISONING
C0338787|T053|191804003|SNOMEDCT_US|CONTINUOUS ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM|CONTINUOUS ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM (DISORDER)
C0338787|T053|191804003|SNOMEDCT_US|CONTINUOUS ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM |CONTINUOUS ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM (DISORDER)
C0338788|T053|191805002|SNOMEDCT_US|EPISODIC ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM|EPISODIC ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM (DISORDER)
C0338788|T053|191805002|SNOMEDCT_US|EPISODIC ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM |EPISODIC ACUTE ALCOHOLIC INTOXICATION IN ALCOHOLISM (DISORDER)
C0856321|T053||SNOMEDCT_US|ALCOHOLISM (EXCLUDING PSYCHOSIS)
C0856321|T053||SNOMEDCT_US|ALCOHOLISM (EXCL PSYCHOSIS)
C0848500|T053||SNOMEDCT_US|DRINKS TOO MUCH
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF SYNDROME|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|PSYCHOSIS, KORSAKOFF|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|SYNDROME, KORSAKOFF|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|WERNICKE KORSAKOFF SYNDROME|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF'S PSYCHOSIS|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|WERNICKE-KORSAKOFF SYNDROME|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|SYNDROME, WERNICKE-KORSAKOFF|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF'S SYNDROME|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|WERNICKE ENCEPHALOPATHY|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF PSYCHOSIS|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF SYNDROME [DISEASE/FINDING]|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF PSYCHOSES|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|PSYCHOSES, KORSAKOFF|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|SYNDROMES, WERNICKE-KORSAKOFF|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|WERNICKE-KORSAKOFF SYNDROMES|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOV'S PSYCHOSIS|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOV PSYCHOSIS|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|WERNICKE-KORSAKOV SYNDROME |WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|WERNICKE-KORSAKOV SYNDROME|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOV PSYCHOSIS |WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF'S PSYCHOSIS |WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|ALCOHOL-INDUCED ENCEPHALOPATHY|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF'S DISEASE|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOV'S SYNDROME|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF'S PSYCHOSIS |WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOV; PSYCHOSIS|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOV|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFFS PSYCHOSIS|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0349464|T053|191472007|SNOMEDCT_US|KORSAKOFF'S PSYCHOSIS, ALCOHOLIC|WERNICKE-KORSAKOV SYNDROME (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC DISORDER|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC DISORDERS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC DISORDER, ALCOHOL|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC DISORDERS, ALCOHOL|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL, AMNESIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF ALCOHOL, AMNESIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC DIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL IND AMNESTIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL IND DYSMNESIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL IND KORSAKOFF SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL IND PERSISTING AMNESTIC DIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC PSYCHOSIS ALCOHOL IND|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL IND AMNESTIC PSYCHOSIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL IND DYSMNESIC PSYCHOSIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED PERSISTING AMNESTIC DISORDER |ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED PERSISTING AMNESTIC DISORDER|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL INDUCED AMNESTIC PSYCHOSIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED AMNESTIC PSYCHOSES|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC PSYCHOSES, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC PSYCHOSIS, ALCOHOL INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|PSYCHOSES, ALCOHOL-INDUCED AMNESTIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|PSYCHOSIS, ALCOHOL-INDUCED AMNESTIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL INDUCED AMNESTIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED AMNESTIC SYNDROMES|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC SYNDROME, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC SYNDROMES, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROME, ALCOHOL-INDUCED AMNESTIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROMES, ALCOHOL-INDUCED AMNESTIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC SYNDROMES|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC SYNDROME, ALCOHOL|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC SYNDROMES, ALCOHOL|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROME, ALCOHOL AMNESTIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROMES, ALCOHOL AMNESTIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL INDUCED DYSMNESIC PSYCHOSIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED DYSMNESIC PSYCHOSES|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|DYSMNESIC PSYCHOSES, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|DYSMNESIC PSYCHOSIS, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|PSYCHOSES, ALCOHOL-INDUCED DYSMNESIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|PSYCHOSIS, ALCOHOL-INDUCED DYSMNESIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL INDUCED DYSMNESIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED DYSMNESIC SYNDROMES|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|DYSMNESIC SYNDROME, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|DYSMNESIC SYNDROMES, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROME, ALCOHOL-INDUCED DYSMNESIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROMES, ALCOHOL-INDUCED DYSMNESIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL INDUCED KORSAKOFF SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED KORSAKOFF SYNDROMES|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOFF SYNDROME, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOFF SYNDROMES, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROME, ALCOHOL-INDUCED KORSAKOFF|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROMES, ALCOHOL-INDUCED KORSAKOFF|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOFF SYNDROME, ALCOHOLIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROME, ALCOHOLIC KORSAKOFF|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC DISORDR|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED DYSMNESIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOLIC KORSAKOFF SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED DYSMNESIC PSYCHOSIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED AMNESTIC PSYCHOSIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED AMNESTIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC PSYCHOSIS, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC DISORDER [DISEASE/FINDING]|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL-INDUCED KORSAKOFF SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOFFS PSYCHOSIS;ALCOHOLIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL INDUCED PERSISTING AMNESTIC DISORDER|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOLIC KORSAKOFF SYNDROMES|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOFF SYNDROMES, ALCOHOLIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROMES, ALCOHOLIC KORSAKOFF|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOFF'S PSYCHOSIS (ALCOHOLIC)|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|[X]KORSAKOV'S PSYCHOSIS, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|[X]MENTAL AND BEHAVIOURAL DISORDERS DUE TO USE OF ALCOHOL: AMNESIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: AMNESIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC SYNDROME NOS |ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|[X]MENTAL AND BEHAVIORAL DISORDERS DUE TO USE OF ALCOHOL: AMNESIC SYNDROME |ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC SYNDROME NOS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOFF'S PSYCHOSIS ALCOHOLIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOV'S PSYCHOSIS, ALCOHOLIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOLIC AMNESTIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESIC SYNDROME DUE TO ALCOHOL|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOV ALCOHOLIC PSYCHOSIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOV SYNDROME - ALCOHOLIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL AMNESTIC DISORDER |ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOV; ALCOHOLISM|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOL; AMNESTIC SYNDROME|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOLISM; KORSAKOV|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|PSYCHOSIS; KORSAKOV, ALCOHOL|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|PSYCHOSIS; ALCOHOLIC, KORSAKOV|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|PSYCHOSIS; ALCOHOLIC, POLYNEURITIC|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|AMNESTIC; SYNDROME, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROME; AMNESTIC, ALCOHOL-INDUCED|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|SYNDROME; AMNESTIC, ALCOHOL|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|ALCOHOLIC KORSAKOFF'S PSYCHOSIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0001940|T053|191473002|SNOMEDCT_US|KORSAKOFFS ALCOHOLIC PSYCHOSIS|ALCOHOL AMNESTIC SYNDROME NOS (DISORDER)
C0154474|T053||SNOMEDCT_US|OTHER AND UNSPECIFIED ALCOHOL DEPENDENCE
C0154474|T053||SNOMEDCT_US|OTHER AND UNSPECIFIED ALCOHOL DEPENDENCE, UNSPECIFIED DRINKING BEHAVIOR
C0154474|T053||SNOMEDCT_US|ALCOH DEP NEC/NOS-UNSPEC
C0154474|T053||SNOMEDCT_US|OTHER AND UNSPECIFIED ALCOHOL DEPENDENCE, UNSPECIFIED
C0683991|T053||SNOMEDCT_US|EX-ALCOHOLIC
