C0040615|T121||RXNORM|ANTIPSYCHOTIC AGENTS
C4048284|T121||RXNORM|BENZODIAZEPINE
C0005064|T121||RXNORM|BENZODIAZEPINES
C0023870|T121|6448|RXNORM|LITHIUM|LITHIUM
C3540800|T121||RXNORM|LITHIUM ANTIPSYCHOTICS
C0287163|T121|83553|RXNORM|SEROQUEL|SEROQUEL
C0072953|T121||RXNORM|RACLOPRIDE
C0072953|T121||RXNORM|BENZAMIDE, 3,5-DICHLORO-N-((1-ETHYL-2-PYRROLIDINYL)-METHYL)-2-HYDROXY-6-METHOXY-
C0072953|T121||RXNORM|RACLOPRIDE [CHEMICAL/INGREDIENT]
C0073393|T121|35636|RXNORM|RISPERIDONE|RISPERIDONE
C0073393|T121|35636|RXNORM|4H-PYRIDO(1,2-A)PYRIMIDIN-4-ONE, 3-(2-(4-(6-FLUORO-1,2-BENZISOXAZOL-3-YL)-1-PIPERIDINYL)ETHYL)-6 ,7,8,9-TETRAHYDRO-2-METHYL-|RISPERIDONE
C0073393|T121|35636|RXNORM|RISPERIDONE |RISPERIDONE
C0073393|T121|35636|RXNORM|RISPERIDONE [CHEMICAL/INGREDIENT]|RISPERIDONE
C0073393|T121|35636|RXNORM|RISPERIDONE |RISPERIDONE
C0073393|T121|35636|RXNORM|RISPERIDONE |RISPERIDONE
C0008286|T121|2403|RXNORM|CHLORPROMAZINE|CHLORPROMAZINE
C0008286|T121|2403|RXNORM|10H-PHENOTHIAZINE-10-PROPANAMINE, 2-CHLORO-N,N-DIMETHYL-|CHLORPROMAZINE
C0008286|T121|2403|RXNORM|2-CHLORO-10-(3-(DIMETHYLAMINO)PROPYL)PHENOTHIAZINE|CHLORPROMAZINE
C0008286|T121|2403|RXNORM|CHLORPROMAZINES |CHLORPROMAZINE
C0008286|T121|2403|RXNORM|CHLORPROMAZINES|CHLORPROMAZINE
C0008286|T121|2403|RXNORM|CHLORPROMAZINE [CHEMICAL/INGREDIENT]|CHLORPROMAZINE
C0008286|T121|2403|RXNORM|CPZ - CHLORPROMAZINE|CHLORPROMAZINE
C0008286|T121|2403|RXNORM|CHLORPROMAZINE |CHLORPROMAZINE
C0008286|T121|2403|RXNORM|CHLORPROMAZINE |CHLORPROMAZINE
C0016368|T121|4496|RXNORM|FLUPHENAZINE|FLUPHENAZINE
C0016368|T121|4496|RXNORM|1-PIPERAZINEETHANOL, 4-(3-(2-(TRIFLUOROMETHYL)-10H-PHENOTHIAZIN-10-YL)PROPYL)-|FLUPHENAZINE
C0016368|T121|4496|RXNORM|1-PIPERAZINEETHANOL, 4-(3-(2-(TRIFLUOROMETHYL)-10H-PHENOTHIAZIN-10-YL)PROPYL)-(9CI)|FLUPHENAZINE
C0016368|T121|4496|RXNORM|FLUPHENAZINE [CHEMICAL/INGREDIENT]|FLUPHENAZINE
C0016368|T121|4496|RXNORM|FLUFENAZIN|FLUPHENAZINE
C0016368|T121|4496|RXNORM|FLUPHENAZINE |FLUPHENAZINE
C0016368|T121|4496|RXNORM|FLUPHENAZINE |FLUPHENAZINE
C0018546|T121|5093|RXNORM|HALOPERIDOL|HALOPERIDOL
C0018546|T121|5093|RXNORM|1-BUTANONE, 4-(4-(4-CHLOROPHENYL)-4-HYDROXY-1-PIPERIDINYL)-1-(4-FLUOROPHENYL)-|HALOPERIDOL
C0018546|T121|5093|RXNORM|4-[4-(4-CHLOROPHENYL)-4-HYDROXY-1-PIPERIDINYL]-1-(4-FLUOROPHENYL)-1-BUTANONE|HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL |HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL [CHEMICAL/INGREDIENT]|HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL [ANTIPSYCHOTIC]|HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL [TICS, CHOREA] [SEE D47..]|HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL [TICS, CHOREA] [SEE D47..] |HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL [ANTIPSYCHOTIC] |HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL |HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL |HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL [ANTIPSYCHOTIC] |HALOPERIDOL
C0018546|T121|5093|RXNORM|HALOPERIDOL [TICS, CHOREA] [SEE D47..] |HALOPERIDOL
C0031935|T121|8331|RXNORM|PIMOZIDE|PIMOZIDE
C0031935|T121|8331|RXNORM|2H-BENZIMIDAZOL-2-ONE, 1-(1-(4,4-BIS(4-FLUOROPHENYL)BUTYL)-4-PIPERIDINYL)-1,3-DIHYDRO-|PIMOZIDE
C0031935|T121|8331|RXNORM|OPIRAN|PIMOZIDE
C0031935|T121|8331|RXNORM|PIMOZIDE |PIMOZIDE
C0031935|T121|8331|RXNORM|PIMOZIDE [CHEMICAL/INGREDIENT]|PIMOZIDE
C0031935|T121|8331|RXNORM|PIMOZIDE |PIMOZIDE
C0031935|T121|8331|RXNORM|PIMOZIDE |PIMOZIDE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE|PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|10H-PHENOTHIAZINE, 2-CHLORO-10-(3-(4-METHYL-1-PIPERAZINYL)PROPYL)-|PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|2-CHLORO-10-(3-(1-METHYL-4-PIPERAZINYL)PROPYL)-PHENOTHIAZINE|PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE |PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE [CHEMICAL/INGREDIENT]|PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE [NAUSEA]|PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE [NAUSEA] |PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE [ANTIPSYCH] [SEE DHE..]|PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE [ANTIPSYCH] [SEE DHE..] |PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE |PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE |PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PCPZ|PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE [ANTIPSYCH] [SEE DHE..] |PROCHLORPERAZINE
C0033229|T121|8704|RXNORM|PROCHLORPERAZINE [NAUSEA] |PROCHLORPERAZINE
C0039943|T121|10502|RXNORM|THIORIDAZINE|THIORIDAZINE
C0039943|T121|10502|RXNORM|10H-PHENOTHIAZINE, 10-(2-(1-METHYL-2-PIPERIDINYL)ETHYL)-2-(METHYLTHIO)-|THIORIDAZINE
C0039943|T121|10502|RXNORM|THIORIDAZINE (DISCONTINUED)|THIORIDAZINE
C0039943|T121|10502|RXNORM|THIORIDAZINE (DISCONTINUED) |THIORIDAZINE
C0039943|T121|10502|RXNORM|THIORIDAZINE [CHEMICAL/INGREDIENT]|THIORIDAZINE
C0039943|T121|10502|RXNORM|THIORIDAZINE |THIORIDAZINE
C0039943|T121|10502|RXNORM|THIORIDAZINE |THIORIDAZINE
C0009079|T121|2626|RXNORM|CLOZAPINE|CLOZAPINE
C0009079|T121|2626|RXNORM|5H-DIBENZO(B,E)(1,4)DIAZEPINE, 8-CHLORO-11-(4-METHYL-1-PIPERAZINYL)-|CLOZAPINE
C0009079|T121|2626|RXNORM|CLOZAPINE |CLOZAPINE
C0009079|T121|2626|RXNORM|CLOZAPINE [CHEMICAL/INGREDIENT]|CLOZAPINE
C0009079|T121|2626|RXNORM|8-CHLORO-11-(4-METHYL-1-PIPERAZINYL)-5H-DIBENZO(B,E)(1,4)DIAZEPINE|CLOZAPINE
C0009079|T121|2626|RXNORM|CLOZAPINE |CLOZAPINE
C0009079|T121|2626|RXNORM|CLOZAPINE |CLOZAPINE
C0016367|T121|4495|RXNORM|FLUPENTHIXOL|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|1-PIPERAZINEETHANOL, 4-(3-(2-(TRIFLUOROMETHYL)-9H-THIOXANTHEN-9-YLIDENE)PROPYL)-|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTIXOL|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|ALPHA-FLUPENTHIXOL|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTHIXOL [CHEMICAL/INGREDIENT]|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|CIS-FLUPENTHIXOL|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|ANTIPSYCHOTICS FLUPENTIXOL|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTIXOL |FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTIXOL [ANTIPSYCHOTIC]|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTHIXOL [ANTIPSYCHOTIC] |FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTHIXOL [ANTIDEPRESSANT]|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTHIXOL [ANTIDEPRESSANT] |FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTHIXOL [ANTIPSYCHOTIC]|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTIXOL [ANTIDEPRESSANT]|FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTIXOL |FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTIXOL |FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTHIXOL [ANTIDEPRESSANT] |FLUPENTHIXOL
C0016367|T121|4495|RXNORM|FLUPENTHIXOL [ANTIPSYCHOTIC] |FLUPENTHIXOL
C0026388|T121|7019|RXNORM|MOLINDONE|MOLINDONE
C0026388|T121|7019|RXNORM|4H-INDOL-4-ONE, 3-ETHYL-1,5,6,7-TETRAHYDRO-2-METHYL-5-(4-MORPHOLINYLMETHYL)-|MOLINDONE
C0026388|T121|7019|RXNORM|MOLINDONE [CHEMICAL/INGREDIENT]|MOLINDONE
C0026388|T121|7019|RXNORM|MOLINDONE |MOLINDONE
C0026388|T121|7019|RXNORM|MOLINDONE |MOLINDONE
C0027999|T121|7394|RXNORM|NIALAMIDE|NIALAMIDE
C0027999|T121|7394|RXNORM|4-PYRIDINECARBOXYLIC ACID, 2-(3-OXO-3-((PHENYLMETHYL)AMINO)PROPYL)HYDRAZIDE|NIALAMIDE
C0027999|T121|7394|RXNORM|1-(2-(BENZYLCARBAMOYL)ETHYL)-2-ISONICOTINOYLHYDRAZINE|NIALAMIDE
C0027999|T121|7394|RXNORM|NIALAMIDE [CHEMICAL/INGREDIENT]|NIALAMIDE
C0027999|T121|7394|RXNORM|NIALAMIDE |NIALAMIDE
C0030815|T121|7974|RXNORM|PENFLURIDOL|PENFLURIDOL
C0030815|T121|7974|RXNORM|4-PIPERIDINOL, 1-(4,4-BIS(4-FLUOROPHENYL)BUTYL)-4-(4-CHLORO-3-(TRIFLUOROMETHYL)PHENYL)-|PENFLURIDOL
C0030815|T121|7974|RXNORM|PENFLURIDOL [CHEMICAL/INGREDIENT]|PENFLURIDOL
C0030815|T121|7974|RXNORM|PENFLURIDOL |PENFLURIDOL
C0035179|T121|9260|RXNORM|RESERPINE|RESERPINE
C0035179|T121|9260|RXNORM|YOHIMBAN-16-CARBOXYLIC ACID, 11,17-DIMETHOXY-18-((3,4,5-TRIMETHOXYBENZOYL)OXY)-, METHYL ESTER, (3BETA,16BETA,17ALPHA,18BETA,20ALPHA)-|RESERPINE
C0035179|T121|9260|RXNORM|(3BETA,16BETA,17ALPHA,18BETA,20ALPHA)-11,17-DIMETHOXY-18-[(3,4,5-TRIMETHOXYBENZOYL)OXY]YOHIMBAN-16-CARBOXYLIC ACID METHYL ESTER|RESERPINE
C0035179|T121|9260|RXNORM|RESERPINE |RESERPINE
C0035179|T121|9260|RXNORM|RESERPINE [CHEMICAL/INGREDIENT]|RESERPINE
C0035179|T121|9260|RXNORM|RESERPINE - CHEMICAL|RESERPINE
C0035179|T121|9260|RXNORM|RESERPINE - CHEMICAL |RESERPINE
C0035179|T121|9260|RXNORM|RESERPINE |RESERPINE
C0035179|T121|9260|RXNORM|RESERPINE |RESERPINE
C0037956|T121||RXNORM|SPIPERONE
C0037956|T121||RXNORM|1,3,8-TRIAZASPIRO(4.5)DECAN-4-ONE, 8-(4-(4-FLUOROPHENYL)-4-OXOBUTYL)-1-PHENYL-
C0037956|T121||RXNORM|SPIROPERIDOL
C0037956|T121||RXNORM|SPIPERONE [CHEMICAL/INGREDIENT]
C0037956|T121||RXNORM|SPIROPERONE
C0037956|T121||RXNORM|SPIPERONE - CHEMICAL 
C0037956|T121||RXNORM|SPIPERONE - CHEMICAL
C0037956|T121||RXNORM|SPIPERONE 
C0038803|T121|10239|RXNORM|SULPIRIDE|SULPIRIDE
C0038803|T121|10239|RXNORM|BENZAMIDE, 5-(AMINOSULFONYL)-N-((1-ETHYL-2-PYRROLIDINYL)METHYL)-2-METHOXY-|SULPIRIDE
C0038803|T121|10239|RXNORM|SULPIRIDE [CHEMICAL/INGREDIENT]|SULPIRIDE
C0038803|T121|10239|RXNORM|SULPERIDE|SULPIRIDE
C0038803|T121|10239|RXNORM|N-((1-ETHYL-2-PYRROLIDINYL)METHYL)-5-SULFAMOYL-O-ANISAMIDE|SULPIRIDE
C0038803|T121|10239|RXNORM|ANTIDEPRESSANTS SULPIRIDE|SULPIRIDE
C0038803|T121|10239|RXNORM|SULPIRIDE |SULPIRIDE
C0038803|T121|10239|RXNORM|SULPIRIDE |SULPIRIDE
C0038803|T121|10239|RXNORM|SULPIRIDE |SULPIRIDE
C0039955|T121|10510|RXNORM|THIOTHIXENE|THIOTHIXENE
C0039955|T121|10510|RXNORM|9H-THIOXANTHENE-2-SULFONAMIDE, N,N-DIMETHYL-9-(3-(4-METHYL-1-PIPERAZINYL)PROPYLIDENE)-|THIOTHIXENE
C0039955|T121|10510|RXNORM|THIOXANTHENE-2-SULFONAMIDE, N,N-DIMETHYL-9-(3-(4-METHYL-1-PIPERAZINYL)PROPYLIDENE)-|THIOTHIXENE
C0039955|T121|10510|RXNORM|N,N-DIMETHYL-9-(3-(4-METHYLPIPERAZIN-1-YL)PROPYLIDENE)-9H-THIOXANTHENE-2-SULPHONAMIDE|THIOTHIXENE
C0039955|T121|10510|RXNORM|NAVARON|THIOTHIXENE
C0039955|T121|10510|RXNORM|ORBINAMON|THIOTHIXENE
C0039955|T121|10510|RXNORM|THIOTHIXENE |THIOTHIXENE
C0039955|T121|10510|RXNORM|THIOTHIXENE [CHEMICAL/INGREDIENT]|THIOTHIXENE
C0039955|T121|10510|RXNORM|TIOTIXENE|THIOTHIXENE
C0039955|T121|10510|RXNORM|THIOTHIXENE |THIOTHIXENE
C0039955|T121|10510|RXNORM|THIOTHIXENE |THIOTHIXENE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|10H-PHENOTHIAZINE, 10-(3-(4-METHYL-1-PIPERAZINYL)PROPYL)-2-(TRIFLUOROMETHYL)-|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|10-(3-(4-METHYL-1-PIPERAZINYL)PROPYL)-2-(TRIFLUOROMETHYL)-10H-PHENOTHIAZINE|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TFP|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE [CHEMICAL/INGREDIENT]|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOROPERAZINE|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUPERAZINE|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE [ANTIPSYCHOTIC]|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE [ANTIPSYCHOTIC] |TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE [NAUSEA] [SEE DH4..] |TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE [NAUSEA] [SEE DH4..]|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|10-[3-(4-METHYL-1-PIPERAZINYL)PROPYL]-2-(TRIFLUOROMETHYL)-10H-PHENOTHIAZINE|TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE |TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE |TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE [ANTIPSYCHOTIC] |TRIFLUOPERAZINE
C0040979|T121|10800|RXNORM|TRIFLUOPERAZINE [NAUSEA] [SEE DH4..] |TRIFLUOPERAZINE
C0871650|T121||RXNORM|ANTISCHIZOPHRENIC DRUGS
C0701357|T121||RXNORM|ICI204636
C0701357|T121||RXNORM|204636, ICI
C0701357|T121||RXNORM|204,636, ICI
C0701357|T121||RXNORM|ICI 204,636
C0701357|T121||RXNORM|ICI-204636
C0701357|T121||RXNORM|ICI 204636
C0171023|T121|61381|RXNORM|2-METHYL-4-(4-METHYL-1-PIPERAZINYL)-10H-THIENO(2,3-B)(1,5)BENZODIAZEPINE|OLANZAPINE
C0171023|T121|61381|RXNORM|OLANZAPINE|OLANZAPINE
C0171023|T121|61381|RXNORM|OLANZAPINE |OLANZAPINE
C0171023|T121|61381|RXNORM|OLANZAPINE [CHEMICAL/INGREDIENT]|OLANZAPINE
C0171023|T121|61381|RXNORM|OLANZAPINE (ZYPREXA)|OLANZAPINE
C0171023|T121|61381|RXNORM|OLANZAPINE |OLANZAPINE
C0171023|T121|61381|RXNORM|OLANZAPINE |OLANZAPINE
C0380393|T121|115698|RXNORM|5-(2-(4-(3-BENZISOTHIAZOLYL)PIPERAZINYL)ETHYL)-6-CHLORO-1,3-DIHYDRO-2H-INDOL-2-ONE|ZIPRASIDONE
C0380393|T121|115698|RXNORM|ZIPRASIDONE|ZIPRASIDONE
C0380393|T121|115698|RXNORM|2H-INDOL-2-ONE, 5-(2-(4-(1,2-BENZISOTHIAZOL-3-YL)-1-PIPERAZINYL)ETHYL)-6-CHLORO-1,3-DIHYDRO-|ZIPRASIDONE
C0380393|T121|115698|RXNORM|ZIPRASIDONE [CHEMICAL/INGREDIENT]|ZIPRASIDONE
C0380393|T121|115698|RXNORM|ZIPRAZIDONE|ZIPRASIDONE
C0380393|T121|115698|RXNORM|ZIPRASIDONE |ZIPRASIDONE
C0380393|T121|115698|RXNORM|ZIPRASIDONE |ZIPRASIDONE
C0597883|T121||RXNORM|ALENTEMOL
C0597884|T121||RXNORM|ANTISCHIZOPHRENIC
C0000959|T121|155|RXNORM|ACEPROMAZINE|ACEPROMAZINE
C0000959|T121|155|RXNORM|ETHANONE, 1-(10-(3-(DIMETHYLAMINO)PROPYL)-10H-PHENOTHIAZIN-2-YL)-|ACEPROMAZINE
C0000959|T121|155|RXNORM|ACEPROMAZINE [CHEMICAL/INGREDIENT]|ACEPROMAZINE
C0000959|T121|155|RXNORM|ACETOPROMAZINE|ACEPROMAZINE
C0000959|T121|155|RXNORM|ACETAZINE|ACEPROMAZINE
C0000959|T121|155|RXNORM|ACETYLPROMAZINE|ACEPROMAZINE
C0000959|T121|155|RXNORM|10-(3-DIMETHYLAMINOPROPYL)PHENOTHIAZINE-3-ETHYLONE|ACEPROMAZINE
C0000959|T121|155|RXNORM|ACEPROMAZINE |ACEPROMAZINE
C0004477|T121||RXNORM|AZAPERONE
C0004477|T121||RXNORM|1-BUTANONE, 1-(4-FLUOROPHENYL)-4-(4-(2-PYRIDINYL)-1-PIPERAZINYL)-
C0004477|T121||RXNORM|AZAPERONE [CHEMICAL/INGREDIENT]
C0004477|T121||RXNORM|AZAPERONE 
C0005013|T121|1373|RXNORM|BENPERIDOL|BENPERIDOL
C0005013|T121|1373|RXNORM|2H-BENZIMIDAZOL-2-ONE, 1-(1-(4-(4-FLUOROPHENYL)-4-OXOBUTYL)-4-PIPERIDINYL)-1,3-DIHYDRO-|BENPERIDOL
C0005013|T121|1373|RXNORM|BENPERIDOL |BENPERIDOL
C0005013|T121|1373|RXNORM|BENPERIDOL - CHEMICAL|BENPERIDOL
C0005013|T121|1373|RXNORM|BENPERIDOL |BENPERIDOL
C0005013|T121|1373|RXNORM|BENPERIDOL - CHEMICAL |BENPERIDOL
C0005013|T121|1373|RXNORM|BENPERIDOL [CHEMICAL/INGREDIENT]|BENPERIDOL
C0005013|T121|1373|RXNORM|BENPERIDOL |BENPERIDOL
C0006467|T121||RXNORM|BUTACLAMOL
C0006467|T121||RXNORM|BUTACLAMOL [CHEMICAL/INGREDIENT]
C0008290|T121|2406|RXNORM|CHLORPROTHIXENE|CHLORPROTHIXENE
C0008290|T121|2406|RXNORM|1-PROPANAMINE, 3-(2-CHLORO-9H-THIOXANTHEN-9-YLIDENE)-N,N-DIMETHYL-, (Z)-|CHLORPROTHIXENE
C0008290|T121|2406|RXNORM|CHLORPROTHIXENE |CHLORPROTHIXENE
C0008290|T121|2406|RXNORM|CHLORPROTIXEN|CHLORPROTHIXENE
C0008290|T121|2406|RXNORM|CHLORPROTHIXENE [CHEMICAL/INGREDIENT]|CHLORPROTHIXENE
C0008290|T121|2406|RXNORM|CHLORPROTHIXENE |CHLORPROTHIXENE
C0008290|T121|2406|RXNORM|CHLORPROTHIXENE |CHLORPROTHIXENE
C0009026|T121||RXNORM|CLOPENTHIXOL
C0009026|T121||RXNORM|1-PIPERAZINEETHANOL, 4-(3-(2-CHLORO-9H-THIOXANTHEN-9-YLIDENE)PROPYL)-
C0009026|T121||RXNORM|CLOPENTHIXOL 
C0009026|T121||RXNORM|CLOPENTHIXOL [CHEMICAL/INGREDIENT]
C0009026|T121||RXNORM|CLOPENTHIXOL, TRANS
C0009026|T121||RXNORM|CLOPENTHIXOL 
C0013136|T121|3648|RXNORM|DROPERIDOL|DROPERIDOL
C0013136|T121|3648|RXNORM|2H-BENZIMIDAZOL-2-ONE, 1-(1-(4-(4-FLUOROPHENYL)-4-OXOBUTYL)-1,2,3,6-TETRAHYDRO-4-PYRIDINYL)-1,3-DIHYDRO-|DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL |DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL [CHEMICAL/INGREDIENT]|DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL [CENTRAL NERVOUS SYSTEM USE] |DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL [CENTRAL NERVOUS SYSTEM USE]|DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL [ANESTHESIA] |DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL [ANAESTHESIA]|DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL [ANESTHESIA]|DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL |DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL |DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL [ANESTHESIA] |DROPERIDOL
C0013136|T121|3648|RXNORM|DROPERIDOL [CENTRAL NERVOUS SYSTEM USE] |DROPERIDOL
C0014958|T121||RXNORM|ETAZOLATE
C0014958|T121||RXNORM|1H-PYRAZOLO(3,4-B)PYRIDINE-5-CARBOXYLIC ACID, 1-ETHYL-4-((1-METHYLETHYLIDENE)HYDRAZINO)-, ETHYL ESTER
C0014958|T121||RXNORM|ETAZOLATE [CHEMICAL/INGREDIENT]
C0016383|T121|4507|RXNORM|FLUSPIRILENE|FLUSPIRILENE
C0016383|T121|4507|RXNORM|1,3,8-TRIAZASPIRO(4.5)DECAN-4-ONE, 8-(4,4-BIS(4-FLUOROPHENYL)BUTYL)-1-PHENYL-|FLUSPIRILENE
C0016383|T121|4507|RXNORM|SPIRODIFLAMINE|FLUSPIRILENE
C0016383|T121|4507|RXNORM|FLUSPIRILENE [CHEMICAL/INGREDIENT]|FLUSPIRILENE
C0016383|T121|4507|RXNORM|FLUSPIRILENE |FLUSPIRILENE
C0016383|T121|4507|RXNORM|FLUSPIRILENE |FLUSPIRILENE
C0024056|T121|6475|RXNORM|LOXAPINE|LOXAPINE
C0024056|T121|6475|RXNORM|DIBENZ(B,F)(1,4)OXAZEPINE, 2-CHLORO-11-(4-METHYL-1-PIPERAZINYL)-|LOXAPINE
C0024056|T121|6475|RXNORM|LOXAPINE |LOXAPINE
C0024056|T121|6475|RXNORM|OXILAPINE|LOXAPINE
C0024056|T121|6475|RXNORM|2-CHLORO-11-(4-METHYL-1-PIPERAZINYL)-DIBENZ(B,F)(1,4)OXAZEPINE|LOXAPINE
C0024056|T121|6475|RXNORM|CLOXAZEPINE|LOXAPINE
C0024056|T121|6475|RXNORM|LOXAPINE [CHEMICAL/INGREDIENT]|LOXAPINE
C0024056|T121|6475|RXNORM|LOXAPINE |LOXAPINE
C0024056|T121|6475|RXNORM|LOXAPINE |LOXAPINE
C0025497|T121|6779|RXNORM|MESORIDAZINE|MESORIDAZINE
C0025497|T121|6779|RXNORM|10H-PHENOTHIAZINE, 10-(2-(1-METHYL-2-PIPERIDINYL)ETHYL)-2-(METHYLSULFINYL)-|MESORIDAZINE
C0025497|T121|6779|RXNORM|MESORIDAZINE |MESORIDAZINE
C0025497|T121|6779|RXNORM|MESORIDAZINE [CHEMICAL/INGREDIENT]|MESORIDAZINE
C0025497|T121|6779|RXNORM|MESORIDAZINE |MESORIDAZINE
C0025497|T121|6779|RXNORM|MESORIDAZINE |MESORIDAZINE
C0025654|T121||RXNORM|METHIOTHEPIN
C0025654|T121||RXNORM|PIPERAZINE, 1-(10,11-DIHYDRO-8-(METHYLTHIO)DIBENZO(B,F)THIEPIN-10-YL)-4-METHYL-
C0025654|T121||RXNORM|METITEPINE
C0025654|T121||RXNORM|METHIOTHEPINE
C0025654|T121||RXNORM|METHIOTHEPIN [CHEMICAL/INGREDIENT]
C0025678|T121|6852|RXNORM|METHOTRIMEPRAZINE|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|10H-PHENOTHIAZINE-10-PROPANAMINE, 2-METHOXY-N,N,BETA-TRIMETHYL-, (R)-|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|METHOTRIMEPRAZINE PRODUCT|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|METHOTRIMEPRAZINE (DISCONTINUED) |METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|METHOTRIMEPRAZINE (DISCONTINUED)|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|LEVOMEPROMAZINE|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|METHOTRIMEPRAZINE [CHEMICAL/INGREDIENT]|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|LEVOMEPRAZIN|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|LEVOPROMAZINE|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|(-)-10-(3-(DIMETHYLAMINO)-2-METHYLPROPYL)-2-METHOXYPHENOTHIAZINE|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|LEVOMEPROMAZINE PRODUCT|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|METHOTRIMEPRAZINE PRODUCT |METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|LEVOMEPRAZINE|METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|METHOTRIMEPRAZINE |METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|METHOTRIMEPRAZINE |METHOTRIMEPRAZINE
C0025678|T121|6852|RXNORM|LEVOMEPROMAZINE PRODUCT |METHOTRIMEPRAZINE
C0030969|T121|8042|RXNORM|PERAZINE|PERAZINE
C0030969|T121|8042|RXNORM|10H-PHENOTHIAZINE, 10-(3-(4-METHYL-1-PIPERAZINYL)PROPYL)-|PERAZINE
C0030969|T121|8042|RXNORM|PERAZINE [CHEMICAL/INGREDIENT]|PERAZINE
C0030969|T121|8042|RXNORM|PERNAZINE|PERAZINE
C0030969|T121|8042|RXNORM|PERAZINE |PERAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE|PERPHENAZINE
C0031184|T121|8076|RXNORM|1-PIPERAZINEETHANOL, 4-(3-(2-CHLORO-10H-PHENOTHIAZIN-10-YL)PROPYL)-|PERPHENAZINE
C0031184|T121|8076|RXNORM|4-[3-(2-CHLORO-10H-PHENOTHIAZIN-10-YL)PROPYL]-1-PIPERAZINEETHANOL|PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE |PERPHENAZINE
C0031184|T121|8076|RXNORM|CHLORPIPRAZINE|PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE [CHEMICAL/INGREDIENT]|PERPHENAZINE
C0031184|T121|8076|RXNORM|PERFENAZINE|PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE [CENTRAL NERVOUS SYSTEM USE]|PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE [ANESTHESIA]|PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE [CENTRAL NERVOUS SYSTEM USE] |PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE [ANESTHESIA] |PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE [ANAESTHESIA]|PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE |PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE |PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE [ANESTHESIA] |PERPHENAZINE
C0031184|T121|8076|RXNORM|PERPHENAZINE [CENTRAL NERVOUS SYSTEM USE] |PERPHENAZINE
C0033399|T121|8742|RXNORM|PROMAZINE|PROMAZINE
C0033399|T121|8742|RXNORM|10H-PHENOTHIAZINE-10-PROPANAMINE, N,N-DIMETHYL-|PROMAZINE
C0033399|T121|8742|RXNORM|PROMAZINE [CHEMICAL/INGREDIENT]|PROMAZINE
C0033399|T121|8742|RXNORM|PROMAZINE |PROMAZINE
C0033399|T121|8742|RXNORM|PROMAZINE |PROMAZINE
C0040988|T121|10804|RXNORM|TRIFLUPERIDOL|TRIFLUPERIDOL
C0040988|T121|10804|RXNORM|1-BUTANONE, 1-(4-FLUOROPHENYL)-4-(4-HYDROXY-4-(3-(TRIFLUOROMETHYL)PHENYL)-1-PIPERIDINYL)-|TRIFLUPERIDOL
C0040988|T121|10804|RXNORM|TRIFLURIDOL|TRIFLUPERIDOL
C0040988|T121|10804|RXNORM|TRIFLUPERIDOL [CHEMICAL/INGREDIENT]|TRIFLUPERIDOL
C0040988|T121|10804|RXNORM|TRIFLUPERIDOL |TRIFLUPERIDOL
C0040988|T121|10804|RXNORM|TRIFLUPERIDOL |TRIFLUPERIDOL
C0040989|T121|10805|RXNORM|TRIFLUPROMAZINE|TRIFLUPROMAZINE
C0040989|T121|10805|RXNORM|10H-PHENOTHIAZINE-10-PROPANAMINE, N,N-DIMETHYL-2-(TRIFLUOROMETHYL)-|TRIFLUPROMAZINE
C0040989|T121|10805|RXNORM|TRIFLUPROMAZINE (DISCONTINUED) |TRIFLUPROMAZINE
C0040989|T121|10805|RXNORM|TRIFLUPROMAZINE (DISCONTINUED)|TRIFLUPROMAZINE
C0040989|T121|10805|RXNORM|TRIFLUOPROMAZINE|TRIFLUPROMAZINE
C0040989|T121|10805|RXNORM|TRIFLUPROMAZINE [CHEMICAL/INGREDIENT]|TRIFLUPROMAZINE
C0040989|T121|10805|RXNORM|FLUOPROMAZINE|TRIFLUPROMAZINE
C0040989|T121|10805|RXNORM|TRIFLUPROMAZINE |TRIFLUPROMAZINE
C0040989|T121|10805|RXNORM|TRIFLUPROMAZINE |TRIFLUPROMAZINE
C0085260|T121||RXNORM|RITANSERIN
C0085260|T121||RXNORM|5H-THIAZOLO(3,2-A)PYRIMIDIN-5-ONE, 6-(2-(4-(BIS(4-FLUOROPHENYL)METHYLENE)-1-PIPERIDINYL)ETHYL)-7-METHYL-
C0085260|T121||RXNORM|RITANSERIN [CHEMICAL/INGREDIENT]
C0085260|T121||RXNORM|6-(2-(4-(BIS(4-FLUOROPHENYL)METHYLENE)-1-PIPERIDINYL)ETHYL)-7-METHYL-5H-THIAZOLO(3,2-A)PYRIMIDIN-5-ONE
C0085260|T121||RXNORM|6-(2-(4-(BIS(P-FLUOROPHENYL)METHYLENE)-PIPERIDINO)ETHYL)-7-METHYL-5H-THIAZOLO-(3,2-A)PYRIMIDIN-5-ONE
C0061851|T121|26225|RXNORM|ONDANSETRON|ONDANSETRON
C0061851|T121|26225|RXNORM|4H-CARBAZOL-4-ONE, 1,2,3,9-TETRAHYDRO-9-METHYL-3-((2-METHYL-1H-IMIDAZOL-1-YL)METHYL)-|ONDANSETRON
C0061851|T121|26225|RXNORM|ONDANSETRON |ONDANSETRON
C0061851|T121|26225|RXNORM|ONDANSETRON [CHEMICAL/INGREDIENT]|ONDANSETRON
C0061851|T121|26225|RXNORM|ONDANSETRON, (+,-)-ISOMER|ONDANSETRON
C0061851|T121|26225|RXNORM|ONDANSETRON |ONDANSETRON
C0061851|T121|26225|RXNORM|ONDANSETRON |ONDANSETRON
C0073047|T121|35350|RXNORM|REMOXIPRIDE|REMOXIPRIDE
C0073047|T121|35350|RXNORM|BENZAMIDE, 3-BROMO-N-((1-ETHYL-2-PYRROLIDINYL)METHYL)-2,6-DIMETHOXY-, (S)-|REMOXIPRIDE
C0073047|T121|35350|RXNORM|REMOXIPRIDE [CHEMICAL/INGREDIENT]|REMOXIPRIDE
C0073047|T121|35350|RXNORM|(S)-3-BROMO-N-((1-ETHYL-2-PYRROLIDINYL)METHYL)-2,6-DIMETHOXYBENZAMIDE|REMOXIPRIDE
C0073047|T121|35350|RXNORM|REMOXIPRIDE |REMOXIPRIDE
C0073047|T121|35350|RXNORM|REMOXIPRIDE |REMOXIPRIDE
C0023870|T121|6448|RXNORM|LITHIUM|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM PRODUCT|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM |LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM [CHEMICAL/INGREDIENT]|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM METALLICUM|LITHIUM
C0023870|T121|6448|RXNORM|LI|LITHIUM
C0023870|T121|6448|RXNORM|LI ELEMENT|LITHIUM
C0023870|T121|6448|RXNORM|LI+ ELEMENT|LITHIUM
C0023870|T121|6448|RXNORM|LI - LITHIUM|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM |LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM |LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM, NOS|LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM PRODUCT |LITHIUM
C0023870|T121|6448|RXNORM|LITHIUM PRODUCT |LITHIUM
C3179399|T121||RXNORM|HYDROCHLORIDE, TIAPAMIL
C3179399|T121||RXNORM|TIAPAMIL HYDROCHLORIDE
C3179399|T121||RXNORM|TIAPAMIL HYDROCHLORIDE [CHEMICAL/INGREDIENT]
C3179399|T121||RXNORM|1,3-DITHIANE-2-PROPANAMINE, 2-(3,4-DIMETHOXYPHENYL)-N-(2-(3,4-DIMETHOXYPHENYL)ETHYL)-N-METHYL-, 1,1,3,3-TETRAOXIDE, HYDROCHLORIDE
C3179399|T121||RXNORM|N-(3,4-DIMETHOXYPHENETHYL)-2-(3,4-DIMETHOXYPHENYL)-N-METHYL-M-DITHIAN-2-PROPYLAMIN-1,1,3,3-TETROXIDE HYDROCHLORIDE
C0040615|T121||RXNORM|AGENTS, ANTIPSYCHOTIC
C0040615|T121||RXNORM|AGENTS, MAJOR TRANQUILIZING
C0040615|T121||RXNORM|AGENTS, MAJOR TRANQUILLIZING
C0040615|T121||RXNORM|ANTIPSYCHOTIC AGENTS
C0040615|T121||RXNORM|MAJOR TRANQUILIZING AGENTS
C0040615|T121||RXNORM|MAJOR TRANQUILLIZING AGENTS
C0040615|T121||RXNORM|ANTIPSYCHOTIC AGENT
C0040615|T121||RXNORM|AGENTS, NEUROLEPTIC
C0040615|T121||RXNORM|DRUGS, ANTIPSYCHOTIC
C0040615|T121||RXNORM|DRUGS, NEUROLEPTIC
C0040615|T121||RXNORM|TRANQUILIZERS, MAJOR
C0040615|T121||RXNORM|NEUROLEPTIC
C0040615|T121||RXNORM|ANTIPSYCHOTICS
C0040615|T121||RXNORM|NEUROLEPTIC AGENT
C0040615|T121||RXNORM|ANTISCHIZOPHRENIC AGENT
C0040615|T121||RXNORM|MAJOR TRANQUILIZER
C0040615|T121||RXNORM|NEUROLOGICAL AGENTS NEUROLEPTICS
C0040615|T121||RXNORM|ANTIPSYCHOTICS 
C0040615|T121||RXNORM|NEUROLEPTICS
C0040615|T121||RXNORM|NEUROLEPTICS 
C0040615|T121||RXNORM|ANTIPSYCHOTIC AGENT [TC]
C0040615|T121||RXNORM|ANTIPSYCHOTIC
C0040615|T121||RXNORM|[CN700] ANTIPSYCHOTICS
C0040615|T121||RXNORM|ANTIPSYCHOTIC DRUG
C0040615|T121||RXNORM|ANTIPSYCHOTIC DRUG 
C0040615|T121||RXNORM|ANTIPSYCHOTIC DRUGS
C0040615|T121||RXNORM|NEUROLEPTIC AGENTS
C0040615|T121||RXNORM|MAJOR TRANQUILIZERS
C0040615|T121||RXNORM|NEUROLEPTIC DRUGS
C0040615|T121||RXNORM|TRANQUILLIZING AGENTS, MAJOR
C0040615|T121||RXNORM|TRANQUILIZING AGENTS, MAJOR
C0040615|T121||RXNORM|NEUROLEPTIC DRUG
C0040615|T121||RXNORM|ANTI-PSYCHOTIC AGENT 
C0040615|T121||RXNORM|ANTI-PSYCHOTIC AGENT 
C0040615|T121||RXNORM|ANTI-PSYCHOTIC AGENT
C0040615|T121||RXNORM|ANTI-PSYCHOTIC AGENT, NOS
C0040615|T121||RXNORM|NEUROLEPTIC DRUG, NOS
C0039623|T121|10390|RXNORM|TETRABENAZINE|TETRABENAZINE
C0039623|T121|10390|RXNORM|2H-BENZO(A)QUINOLIZIN-2-ONE, 1,3,4,6,7,11B-HEXAHYDRO-9,10-DIMETHOXY-3-(2-METHYLPROPYL)-|TETRABENAZINE
C0039623|T121|10390|RXNORM|TETRABENAZINE ORPHAN BRAND|TETRABENAZINE
C0039623|T121|10390|RXNORM|2-OXO-3-ISOBUTYL-9,10-DIMETHOXY-1,3,4,6,7,11-BETA-HEXAHYDRO-|TETRABENAZINE
C0039623|T121|10390|RXNORM|ORPHAN BRAND OF TETRABENAZINE|TETRABENAZINE
C0039623|T121|10390|RXNORM|TETRABENAZINE [CHEMICAL/INGREDIENT]|TETRABENAZINE
C0039623|T121|10390|RXNORM|NEUROLOGICAL AGENTS TETRABENAZINE|TETRABENAZINE
C0039623|T121|10390|RXNORM|TETRABENAZINE |TETRABENAZINE
C0039623|T121|10390|RXNORM|TETRABENAZINE PRODUCT|TETRABENAZINE
C0039623|T121|10390|RXNORM|TETRABENAZINE |TETRABENAZINE
C0039623|T121|10390|RXNORM|TETRABENAZINE PRODUCT |TETRABENAZINE
C0039623|T121|10390|RXNORM|TETRABENAZINE PRODUCT |TETRABENAZINE
C0304370|T121||RXNORM|PHENOTHIAZINE DERIVATIVES
C0304370|T121||RXNORM|PHENOTHIAZINE DERIVATIVES 
C0304370|T121||RXNORM|PHENOTHIAZINE DERIVATIVE 
C0304370|T121||RXNORM|PHENOTHIAZINE DERIVATIVE ANTIPSYCHOTIC
C0304370|T121||RXNORM|PHENOTHIAZINE DERIVATIVE
C0304370|T121||RXNORM|PHENOTHIAZINE DERIVATIVE ANTIPSYCHOTIC 
C0304370|T121||RXNORM|PHENOTHIAZINE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304370|T121||RXNORM|PHENOTHIAZINE DERIVATIVE ANTIPSYCHOTIC AGENT
C0304370|T121||RXNORM|PHENOTHIAZINE AND/OR DERIVATIVE
C0304370|T121||RXNORM|PHENOTHIAZINE AND/OR DERIVATIVE 
C0304370|T121||RXNORM|PHENOTHIAZINE DERIVATIVE 
C0304370|T121||RXNORM|PHENOTHIAZINE AND/OR DERIVATIVE 
C0304370|T121||RXNORM|PHENOTHIAZINES
C0301410|T121||RXNORM|HYDROXYPHENAMATE
C0301410|T121||RXNORM|2-HYDROXY-2-PHENYLBUTYL CARBAMATE
C0301410|T121||RXNORM|HYDROXYPHENAMATE 
C0301410|T121||RXNORM|OXYFENAMATE
C0165561|T121||RXNORM|2-METHYL-5-(4-METHYL-1-PIPERAZINYL)-11H-(1,2,4)TRIAZOLO(1,5-C)(1,3)BENZODIAZEPINE
C0165561|T121||RXNORM|11H-(1,2,4)TRIAZOLO(1,5-C)(1,3)BENZODIAZEPINE, 2-METHYL-5-(4-METHYL-1-PIPERAZINYL)-
C0165561|T121||RXNORM|BATELAPINE
C2698335|T121||RXNORM|BATELAPINE MALEATE
C0054138|T121|19777|RXNORM|4-(4-(4-BROMOPHENYL)-4-HYDROXYPIPERIDINO)-4'-FLUOROBUTYROPHENONE|BROMPERIDOL
C0054138|T121|19777|RXNORM|BROMOPERIDOL|BROMPERIDOL
C0054138|T121|19777|RXNORM|BROMPERIDOL|BROMPERIDOL
C0054138|T121|19777|RXNORM|BROMPERIDOL |BROMPERIDOL
C1321935|T121||RXNORM|BUTAPERAZINE MALEATE 
C1321935|T121||RXNORM|BUTAPERAZINE MALEATE
C0133602|T121||RXNORM|(2-(4-(6-FLUORO-1,2-BENZISOXAZOL-3-YL)-1-PIPERIDINYL)ETHYL)-2,9-DIMETHYL-4H-PYRIDO(1,2-A)PYRIMIDIN-4-ONE
C0133602|T121||RXNORM|OCAPERIDONE
C0133602|T121||RXNORM|4H-PYRIDO(1,2-A)PYRIMIDIN-4-ONE, 3-(2-(4-(6-FLUORO-1,2-BENZISOXAZOL-3-YL)-1-PIPERIDINYL)ETHYL)-2,9-DIMETHYL-
C2698647|T121|1294588|RXNORM|OLANZAPINE PAMOATE|OLANZAPINE PAMOATE
C0137024|T121||RXNORM|BENZAMIDE, 3,5-DIMETHYL-N-(4-PYRIDINYLMETHYL)-
C0137024|T121||RXNORM|N-(4-PICOLYL)-3,5-DIMETHYLBENZAMIDE
C0137024|T121||RXNORM|PICOBENZIDE
C2699086|T121||RXNORM|RILAPINE
C0076043|T121||RXNORM|2-TRIFLUORMETHYL-6-FLUORO-9-(3-(4-(2-HYDROXYPIPERAZIN-1-YL))PROPYL)THIOXANTHENE
C0076043|T121||RXNORM|TEFLUTIXOL
C2699912|T121||RXNORM|TENILAPINE
C0076666|T121||RXNORM|TIENOCARBIN
C0076666|T121||RXNORM|TIENOCARBINE
C0076685|T121||RXNORM|10-FLUORO-1,2,3,4,4A,5-HEXAHYDRO-3-METHYL-7-(2-THIENYL)PYRAZINO(1,2-A)(1,4)BENZODIAZEPINE
C0076685|T121||RXNORM|TIMELOTEM
C2699946|T121||RXNORM|TIMIRDINE
C2699963|T121||RXNORM|TOLPIPRAZOLE
C2700075|T121||RXNORM|TRICLODAZOL
C2699390|T121||RXNORM|CLOXYPENDYL
C2698342|T121||RXNORM|BELAPERIDONE
C2698342|T121||RXNORM|(+)-3-(2-((1S,5R,6S)-6-(P-FLUOROPHENYL)-3-AZABICYCLO(3.2.0)HEPT-3-YL)ETHYL)-2,4(1H,3H)-QUINAZOLINEDIONE
C2699631|T121||RXNORM|3,5-DICHLOR-N-(2-(DIETHYLAMINO)ETHYL)-2-METHOXYBENZAMID
C2699631|T121||RXNORM|DICLOMETIDE
C2719618|T121|860647|RXNORM|ASENAPINE MALEATE|ASENAPINE MALEATE
C2719618|T121|860647|RXNORM|1H-DIBENZ(2,3:6,7)OXEPINO(4,5-C)PYRROLE, 5-CHLORO-2,3,3A,12B-TETRAHYDRO-2-METHYL-,(3AR,12BR)-REL-, (2Z)-2-BUTENEDIOATE (1:1)|ASENAPINE MALEATE
C2719618|T121|860647|RXNORM|5-CHLORO-2,3,3A,12B-TETRAHYDRO-2-METHYL-1H-DIBENZ(2,3-6,7)OXEPINO(4,5-C)PYRROLE|ASENAPINE MALEATE
C2699376|T121||RXNORM|4-(2-CHLOROXANTHEN-9-YLIDENE)-1-METHYLPIPERIDINE
C2699376|T121||RXNORM|CLOPIPAZAN
C0668910|T121||RXNORM|CARVOTROLINE
C0668910|T121||RXNORM|1H-PYRIDO(4,3-B)INDOLE, 8-FLUORO-2,3,4,5-TETRAHYDRO-2-(2-(4-PYRIDINYL)ETHYL)-
C0770896|T121||RXNORM|THIOPROPERAZINE MESYLATE
C0770896|T121||RXNORM|THIOPROPERAZINE METHANESULFONATE
C0936105|T121|282427|RXNORM|AMITRIPTYLINE + PERPHENAZINE |AMITRIPTYLINE / PERPHENAZINE
C0936105|T121|282427|RXNORM|AMITRIPTYLINE + PERPHENAZINE|AMITRIPTYLINE / PERPHENAZINE
C0936105|T121|282427|RXNORM|AMITRIPTYLINE/PERPHENAZINE|AMITRIPTYLINE / PERPHENAZINE
C0936105|T121|282427|RXNORM|AMITRIPTYLINE-PERPHENAZINE|AMITRIPTYLINE / PERPHENAZINE
C0936105|T121|282427|RXNORM|AMITRIPTYLINE, PERPHENAZINE DRUG COMBINATION|AMITRIPTYLINE / PERPHENAZINE
C0936105|T121|282427|RXNORM|AMITRIPTYLINE - PERPHENAZINE|AMITRIPTYLINE / PERPHENAZINE
C0936105|T121|282427|RXNORM|AMITRIPTYLINE-PERPHENAZINE COMBINATION|AMITRIPTYLINE / PERPHENAZINE
C0936105|T121|282427|RXNORM|AMITRIPTYLINE / PERPHENAZINE|AMITRIPTYLINE / PERPHENAZINE
C0936105|T121|282427|RXNORM|PERPHENAZINE-AMITRIPTYLINE COMBINATION|AMITRIPTYLINE / PERPHENAZINE
C0066682|T121|30129|RXNORM|FLUPHENAZINE ENANTHATE|FLUPHENAZINE ENANTHATE
C0066682|T121|30129|RXNORM|FLUOHENAZINE ENANTHATE|FLUPHENAZINE ENANTHATE
C0066682|T121|30129|RXNORM|FLUPHENAZINE ENANTHATE (DISCONTINUED) |FLUPHENAZINE ENANTHATE
C0066682|T121|30129|RXNORM|FLUPHENAZINE ENANTHATE (DISCONTINUED)|FLUPHENAZINE ENANTHATE
C0066682|T121|30129|RXNORM|FLUPHENAZINE ENANTHATE [CHEMICAL/INGREDIENT]|FLUPHENAZINE ENANTHATE
C0066682|T121|30129|RXNORM|FLUPHENAZINE ENANTHATE |FLUPHENAZINE ENANTHATE
C0066682|T121|30129|RXNORM|FLUPHENAZINE ENANTHATE |FLUPHENAZINE ENANTHATE
C0066682|T121|30129|RXNORM|FLUOPHENAZINE ENANTHATE|FLUPHENAZINE ENANTHATE
C0066682|T121|30129|RXNORM|FLUOPHENAZINE ENANTHATE |FLUPHENAZINE ENANTHATE
C0078168|T121|39468|RXNORM|VERALIPRIDE|VERALIPRIDE
C0078168|T121|39468|RXNORM|N-(1-ALLYL-2-PYRROLIDINYL)METHYL-2,3-DIMETHOXY-5-SULFAMOYLBENZAMIDE|VERALIPRIDE
C0078168|T121|39468|RXNORM|VERALIPRIDE |VERALIPRIDE
C0009071|T121|2620|RXNORM|CLOTHIAPINE|CLOTHIAPINE
C0009071|T121|2620|RXNORM|CLOTIAPINE|CLOTHIAPINE
C0009071|T121|2620|RXNORM|DIBENZO(B,F)(1,4)THIAZEPINE, 2-CHLORO-11-(4-METHYL-1-PIPERAZINYL)-|CLOTHIAPINE
C0009071|T121|2620|RXNORM|CLOTHIAPINE |CLOTHIAPINE
C0009071|T121|2620|RXNORM|CLOTIAPINE |CLOTHIAPINE
C2000088|T121|784649|RXNORM|ASENAPINE|ASENAPINE
C2000088|T121|784649|RXNORM|ASENAPINE |ASENAPINE
C2000088|T121|784649|RXNORM|ASENAPINE |ASENAPINE
C2000088|T121|784649|RXNORM|ANTIPSYCHOTICS ASENAPINE|ASENAPINE
C2000088|T121|784649|RXNORM|ASENAPINE |ASENAPINE
C0951571|T121|289326|RXNORM|CARPIPRAMINE DIHYDROCHLORIDE|CARPIPRAMINE DIHYDROCHLORIDE
C0050458|T121|16735|RXNORM|ACETOPHENAZINE|ACETOPHENAZINE
C0050458|T121|16735|RXNORM|ACETOPHENAZINE [CHEMICAL/INGREDIENT]|ACETOPHENAZINE
C0050458|T121|16735|RXNORM|ACETOPHENAZINE |ACETOPHENAZINE
C2825691|T121||RXNORM|LORPIPRAZOLE
C0033459|T121|8766|RXNORM|PERICYAZINE|PERICIAZINE
C0033459|T121|8766|RXNORM|PERICIAZINE|PERICIAZINE
C0033459|T121|8766|RXNORM|PERICYAZINE |PERICIAZINE
C0033459|T121|8766|RXNORM|PROPERICIAZINE|PERICIAZINE
C0033459|T121|8766|RXNORM|PERICYAZINE |PERICIAZINE
C0033459|T121|8766|RXNORM|PERICYAZINE |PERICIAZINE
C2825692|T121||RXNORM|CLOPIPAZAN MESYLATE
C0060479|T121||RXNORM|6,8-DIFLUORO-2,3,4,9-TETRAHYDRO-N,N-DIMETHYL-1H-CARBAZOLE-3-AMINE
C0060479|T121||RXNORM|FLUCINDOLE
C2825693|T121||RXNORM|FENIMIDE
C0772014|T121|236710|RXNORM|PROTHIPENDYL HYDROCHLORIDE|PROTHIPENDYL HYDROCHLORIDE
C2825694|T121||RXNORM|CLOTHIXAMIDE MALEATE
C2825695|T121||RXNORM|CYCLOPHENAZINE HYDROCHLORIDE
C0068168|T121||RXNORM|3-(3-HYDROXYPHENYL)-N-N-PROPYLPIPERIDINE
C0068168|T121||RXNORM|3-PPP
C0068168|T121||RXNORM|N-N-PROPYL-3(N-HYDROXYPHENYL)PIPERIDINE
C0068168|T121||RXNORM|PHENOL, 3-(1-PROPYL-3-PIPERIDINYL)-
C0068168|T121||RXNORM|PRECLAMOL
C0068168|T121||RXNORM|(-)-(S)-M-(1-PROPYL-3-PIPERIDYL)PHENOL
C0068168|T121||RXNORM|N-N-PROPYL-3-(3-HYDROXYPHENYL)PIPERIDINE
C2827084|T121||RXNORM|BENZINDOPYRINE
C0247194|T121|73178|RXNORM|ETHANONE, 1-(4-(3-(4-(6-FLUORO-1,2-BENZISOXAZOL-3-YL)-1-PIPERIDINYL)PROPOXY)-3-METHOXYPHENYL)-|ILOPERIDONE
C0247194|T121|73178|RXNORM|ILOPERIDONE|ILOPERIDONE
C0247194|T121|73178|RXNORM|ILOPERIDONE |ILOPERIDONE
C0247194|T121|73178|RXNORM|ILOPERIDONE |ILOPERIDONE
C0247194|T121|73178|RXNORM|4'-(3-(4-(6-FLUORO-1,2-BENZISOXAZOL-3-YL)PIPERIDINO)PROPOXY)-3'-METHOXYACETOPHENONE|ILOPERIDONE
C0247194|T121|73178|RXNORM|ANTIPSYCHOTICS ILOPERIDONE|ILOPERIDONE
C0247194|T121|73178|RXNORM|ILOPERIDONE |ILOPERIDONE
C0072200|T121||RXNORM|PROPIONYLPROMAZINE
C0072200|T121||RXNORM|PROPIOPROMAZINE
C0072200|T121||RXNORM|1-PROPANONE, 1-(10-(3-(DIMETHYLAMINO)PROPYL)-10H-PHENOTHIAZIN-2-YL)-
C0072200|T121||RXNORM|1-PROPANONE, 1-(10-(3-(DIMETHYLAMINO)PROPYL)PHENOTHIAZIN-2-YL)-
C0072200|T121||RXNORM|1-(10-(3-(DIMETHYLAMINO)PROPYL)-10H-PHENOTHIAZIN-2-YL)PROPAN-1-ONE
C0954036|T121||RXNORM|PROPIOPROMAZINE HYDROCHLORIDE
C0954036|T121||RXNORM|1-(10-(3-(DIMETHYLAMINO)PROPYL)-10H-PHENOTHIAZIN-2-YL)-1-PROPANONE
C0954036|T121||RXNORM|1-PROPANONE, 1-(10-(3-(DIMETHYLAMINO)PROPYL)-10H-PHENOTHIAZIN-2-YL)-, MONOHYDROCHLORIDE
C0954036|T121||RXNORM|PROPIONYLPROMAZINE HYDROCHLORIDE
C0954036|T121||RXNORM|PROPIOPROMAZINE HYDROCHLORIDE 
C0139007|T121|55244|RXNORM|PROTHIPENDYL|PROTHIPENDYL
C0139007|T121|55244|RXNORM|PROTHIPENDYL |PROTHIPENDYL
C0075591|T121||RXNORM|SULFORIDAZINE
C2026712|T121||RXNORM|CERULETIDE DIETHYLAMINE (DISCONTINUED) 
C2026712|T121||RXNORM|NEUROLEPTICS CERULETIDE DIETHYLAMINE (DISCONTINUED)
C2026712|T121||RXNORM|CERULETIDE DIETHYLAMINE (DISCONTINUED)
C2092061|T121||RXNORM|TRADITIONAL ANTIPSYCHOTICS 
C2092061|T121||RXNORM|TRADITIONAL ANTIPSYCHOTICS
C2092062|T121||RXNORM|NOVEL ANTIPSYCHOTICS
C2092062|T121||RXNORM|NOVEL ANTIPSYCHOTICS 
C1875654|T121||RXNORM|PHENOTHIAZINE/RELATED ANTIPSYCHOTICS
C1875654|T121||RXNORM|[CN701] PHENOTHIAZINE/RELATED ANTIPSYCHOTICS
C1874317|T121||RXNORM|ANTIPSYCHOTICS,OTHER
C1874317|T121||RXNORM|[CN709] ANTIPSYCHOTICS,OTHER
C2719626|T121|858045|RXNORM|PALIPERIDONE PALMITATE|PALIPERIDONE PALMITATE
C2719626|T121|858045|RXNORM|HEXADECANOIC ACID, 3-(2-(4-(6-FLUORO-1,2-BENZISOXAZOL-3-YL)-1-PIPERIDINYL)ETHYL)-6,7,8,9-TETRAHYDRO-2-METHYL-4-OXO-4H-PYRIDO(1,2-A)PYRIMIDIN-9-YL ESTER|PALIPERIDONE PALMITATE
C2719626|T121|858045|RXNORM|PALIPERIDONE PALMITATE |PALIPERIDONE PALMITATE
C2719626|T121|858045|RXNORM|PALMITATE, PALIPERIDONE|PALIPERIDONE PALMITATE
C2719626|T121|858045|RXNORM|PALIPERIDONE PALMITATE [CHEMICAL/INGREDIENT]|PALIPERIDONE PALMITATE
C2719626|T121|858045|RXNORM|ANTIPSYCHOTICS PALIPERIDONE PALMITATE|PALIPERIDONE PALMITATE
C2719626|T121|858045|RXNORM|PALIPERIDONE PALMITATE |PALIPERIDONE PALMITATE
C0031968|T121|8348|RXNORM|10H-PHENOTHIAZINE-2-SULFONAMIDE,10-(3-(4-(2-HYDROXYETHYL)-1-PIPERIDINYL)PROPYL)-N,N-DIMETHYL-|PIPOTHIAZINE
C0031968|T121|8348|RXNORM|PIPOTHIAZINE|PIPOTHIAZINE
C0031968|T121|8348|RXNORM|PIPOTIAZIN|PIPOTHIAZINE
C0031968|T121|8348|RXNORM|PIPOTIAZINE|PIPOTHIAZINE
C0031968|T121|8348|RXNORM|10-[3-[4-(2-HYDROXYETHYL)PIPERIDINO]PROPYL]-N,N-DIMETHYLPHENOTHIAZINE-2-SULFONAMIDE|PIPOTHIAZINE
C0031968|T121|8348|RXNORM|PIPOTHIAZINE |PIPOTHIAZINE
C0031968|T121|8348|RXNORM|PIPOTIAZINE |PIPOTHIAZINE
C0031968|T121|8348|RXNORM|PIPOTHIAZINE |PIPOTHIAZINE
C2983804|T121||RXNORM|CINUPERONE
C2983866|T121||RXNORM|LUSAPERIDONE
C0066451|T121||RXNORM|2-METHYL-11-(4-METHYL-1-PIPERAZINYL)-DIBENZO (B,F)(1,4)THIAZEPINE
C0066451|T121||RXNORM|METIAPINE
C0069710|T121||RXNORM|10-(3-(4-(2-(1,3-DIOXAN-2-YL)ETHYL)-1- PIPERAZINYL)PROPYL)-2-TRIFLUOROMETHYLPHENOTHIAZINE
C0069710|T121||RXNORM|OXAFLUMAZINE
C0533453|T121||RXNORM|3-(3-(4--(5-METHOXY-4-PYRIMIDINYL)-1-PIPERAZINYL)PROPYL)-N-METHYL-1H-INDOLE-5-METHANESULFONAMIDE FUMARATE
C0533453|T121||RXNORM|3-(3-(4-(5-METHOXY-4-PYRIMIDINYL)-1-PIPERAZINYL)PROPYL)-N-METHYLINDOLE-5-METHANESULFONAMIDE
C0533453|T121||RXNORM|AVITRIPTAN
C0006481|T121||RXNORM|BUTAPERAZINE
C0006481|T121||RXNORM|BUTYRYLPERAZINE
C0006481|T121||RXNORM|1-BUTANONE, 1-(10-(3-(4-METHYL-1-PIPERAZINYL)PROPYL)-10H-PHENOTHIAZIN-2-YL)-
C0006481|T121||RXNORM|BUTAPERIZINE
C0006481|T121||RXNORM|BUTAPERAZINE 
C2825448|T121||RXNORM|CLOTHIXAMIDE
C2825448|T121||RXNORM|CLOTIXAMIDE
C0770895|T121|235745|RXNORM|PIPOTHIAZIN PALMITATE|PIPOTIAZINE PALMITATE
C0770895|T121|235745|RXNORM|PIPOTHIAZINE PALMITATE|PIPOTIAZINE PALMITATE
C0770895|T121|235745|RXNORM|HEXADECANOIC ACID, 2-(1-(3-(2-((DIMETHYLAMINO)SULFONYL)-10H-PHENOTHIAZIN-10-YL)PROPYL)-4-PIPERIDINYL)ETHYL ESTER|PIPOTIAZINE PALMITATE
C0770895|T121|235745|RXNORM|PIPOTIAZINE PALMITATE|PIPOTIAZINE PALMITATE
C0770895|T121|235745|RXNORM|PIPOTIAZINE PALMITATE |PIPOTIAZINE PALMITATE
C0770895|T121|235745|RXNORM|10-(3-(4-(2-HYDROXYETHYL)PIPERIDINO)PROPYL)-N,N-DIMETHYLPHENOTHIAZINE-2-SULFONAMIDE PALMITATE (ESTER)|PIPOTIAZINE PALMITATE
C0770895|T121|235745|RXNORM|PIPOTHIAZINE PALMITATE |PIPOTIAZINE PALMITATE
C0770895|T121|235745|RXNORM|PIPOTIAZINE PALMITATE |PIPOTIAZINE PALMITATE
C0770895|T121|235745|RXNORM|PIPOTHIAZINE PALMITATE |PIPOTIAZINE PALMITATE
C0149491|T121|58338|RXNORM|CLOPENTHIXOL ACETATE ESTER|ZUCLOPENTHIXOL ACETATE
C0149491|T121|58338|RXNORM|ZUCLOPENTHIXOL ACETATE|ZUCLOPENTHIXOL ACETATE
C0149491|T121|58338|RXNORM|(Z)-4-[3-(2-CHLOROTHIOXANTHEN-9-YLIDENE)PROPYL]-1-PIPERAZINEETHANOL ACETATE|ZUCLOPENTHIXOL ACETATE
C0149491|T121|58338|RXNORM|ZUCLOPENTHIXOL ACETATE |ZUCLOPENTHIXOL ACETATE
C0149491|T121|58338|RXNORM|ZUCLOPENTHIXOL ACETATE |ZUCLOPENTHIXOL ACETATE
C0149492|T121|58339|RXNORM|ZUCLOPENTHIXOL DECANOATE|ZUCLOPENTHIXOL DECANOATE
C0149492|T121|58339|RXNORM|DECANOIC ACID, 2-(4-(3-(2-CHLORO-9H-THIOXANTHEN-9-YLIDENE)PROPYL)-1-PIPERAZINYL)ETHYL ESTER, (Z)-|ZUCLOPENTHIXOL DECANOATE
C0149492|T121|58339|RXNORM|ZUCLOPENTHIXOL DECANOATE |ZUCLOPENTHIXOL DECANOATE
C0149492|T121|58339|RXNORM|ZUCLOPENTHIXOL DECANOATE |ZUCLOPENTHIXOL DECANOATE
C0149492|T121|58339|RXNORM|ZUCLOPENTHIXOLE DECANOATE|ZUCLOPENTHIXOL DECANOATE
C0350505|T121|102546|RXNORM|ZUCLOPENTHIXOL DIHYDROCHLORIDE|ZUCLOPENTHIXOL DIHYDROCHLORIDE
C0350505|T121|102546|RXNORM|ZUCLOPENTHIXOL DIHYDROCHLORIDE |ZUCLOPENTHIXOL DIHYDROCHLORIDE
C0350505|T121|102546|RXNORM|CIS-CLOPENTHIXOL HYDROCHLORIDE|ZUCLOPENTHIXOL DIHYDROCHLORIDE
C0350505|T121|102546|RXNORM|(Z)-4-(3-(2-CHLORO-9H-THIOXANTHEN-9-YLIDENE)PROPYL)-1-PIPERAZINEETHANOL DIHYDROCHLORIDE|ZUCLOPENTHIXOL DIHYDROCHLORIDE
C0350505|T121|102546|RXNORM|ZUCLOPENTHIXOL HYDROCHLORIDE|ZUCLOPENTHIXOL DIHYDROCHLORIDE
C0350505|T121|102546|RXNORM|ZUCLOPENTHIXOL DIHYDROCHLORIDE |ZUCLOPENTHIXOL DIHYDROCHLORIDE
C0075662|T121||RXNORM|6-(7-CHLORO-1,8-NAPHTHYRIDIN-2-YL)-2,3,6,7-TETRAHYDRO-7-OXO-5H-(1,4)DITHIINO(2,3-C)PYRROL-5-YL-4-METHYLPIPERAZINE-1-CARBOXYLATE
C0075662|T121||RXNORM|SURICLONE
C0075662|T121||RXNORM|(R,S)-6-(7-CHLOR-1,8-NAPHTHYRIDIN-2-YL)-3,5,6,7-TETRAHYDRO-5-OXO-2H-(1,4)DITHIXINO(2,3-C)PYRROL-7-YL-4-METHYL-1-PIPERAZINYLCARBOXYLAT
C0075662|T121||RXNORM|4-METHYL-1-PIPERAZINECARBOXYLIC ACID ESTER WITH (+-)-6-(7-CHLORO-1,8-NAPHTHYRIDIN-2-YL)-2,3,6,7-TETRAHYDRO-7-HYDROXY-5H-P-DITHIINO(2,3-C)PYRROL-5-ONE
C0075662|T121||RXNORM|(8-(7-CHLORO(1,8)NAPHTHYRIDIN-2-YL)-7-OXO-2,5-DITHIA-8-AZABICYCLO(4.3.0)NON-10-EN-9-YL) 4-METHYLPIPERAZINE-1-CARBOXYLATE
C0006525|T121||RXNORM|BUTYROPHENONES
C0006525|T121||RXNORM|BUTYROPHENONE
C0006525|T121||RXNORM|BUTYROPHENONE 
C0006525|T121||RXNORM|BUTYROPHENONES [CHEMICAL/INGREDIENT]
C0006525|T121||RXNORM|1-PHENYLBUTAN-1-ONE
C0006525|T121||RXNORM|BUTYROPHENONE PRODUCT
C0006525|T121||RXNORM|BUTYROPHENONE 
C0886927|T121||RXNORM|TIAPRIDE HYDROCHLORIDE
C0886927|T121||RXNORM|MONOHYDROCHLORIDE, TIAPRIDE
C0886927|T121||RXNORM|HYDROCHLORIDE, TIAPRIDE
C0886927|T121||RXNORM|TIAPRIDE HYDROCHLORIDE [CHEMICAL/INGREDIENT]
C0886927|T121||RXNORM|TIAPRIDE MONOHYDROCHLORIDE
C0886927|T121||RXNORM|N,N-DIETHYL-2-((2-METHOXY-5-(METHYLSULFONYL)BENZOYL)AMINO)ETHANAMINIUM CHLORIDE
C2983907|T121||RXNORM|PENTIAPINE MALEATE
C0039961|T121||RXNORM|THIOXANTHENES
C0039961|T121||RXNORM|THIOXANTHENES [CHEMICAL/INGREDIENT]
C0039961|T121||RXNORM|THIOXANTHENE 
C0039961|T121||RXNORM|THIOXANTHENE
C0039961|T121||RXNORM|THIOXANTHENE 
C0064748|T121||RXNORM|4'-FLUORO-4-(4-(P-FLUOROBENOZYL)PIPERIDINO)BUTYROPHENONE
C0064748|T121||RXNORM|LENPERONE
C0064748|T121||RXNORM|LENPERONE 
C0175156|T121||RXNORM|AZACYCLONOL
C0175156|T121||RXNORM|DIPHENYL CARBINOL
C0175156|T121||RXNORM|AZACYCLONOL 
C0380392|T121|1294533|RXNORM|ZIPRASIDONE HYDROCHLORIDE|ZIPRASIDONE HYDROCHLORIDE
C0380392|T121|1294533|RXNORM|5-(2-(4-(1,2-BENZISOTHIAZOL-3-YL)-1-PIPERAZINYL)ETHYL)-6-CHLORO-1,3-DIHYDRO-2H-INDOL-2-ONE MONOHYDROCHLORIDE|ZIPRASIDONE HYDROCHLORIDE
C0380392|T121|1294533|RXNORM|ZIPRASIDONE HYDROCHLORIDE |ZIPRASIDONE HYDROCHLORIDE
C0380392|T121|1294533|RXNORM|ANTIPSYCHOTICS ZIPRASIDONE HYDROCHLORIDE|ZIPRASIDONE HYDROCHLORIDE
C0380392|T121|1294533|RXNORM|ZIPRASIDONE HYDROCHLORIDE |ZIPRASIDONE HYDROCHLORIDE
C0608826|T121|161203|RXNORM|ACEPROMETAZINE|ACEPROMETAZINE
C0608826|T121|161203|RXNORM|1-(10-(2-(DIMETHYLAMINO)PROPYL)-10H-PHENOTHIAZIN- 2-YL)ETHANONE|ACEPROMETAZINE
C0654391|T121|186024|RXNORM|4-(4-BROMOPHENYL)-1-(4-(4-FLUOROPHENYL)-4-OXOBUTYL)-4-PIPERIDINYL DECANOATE|BROMPERIDOL DECANOATE
C0654391|T121|186024|RXNORM|BROMPERIDOL DECANOATE|BROMPERIDOL DECANOATE
C0654391|T121|186024|RXNORM|BROMPERIDOL DECANOATE |BROMPERIDOL DECANOATE
C1981574|T121||RXNORM|ANTIPSYCHOTICS &#X7C; URINE
C1994723|T121||RXNORM|PIMOZIDE &#X7C; BLD-SER-PLAS
C0060157|T121||RXNORM|2-ETHYLAMINO-3-PHENYLNORCAMPHANE
C0060157|T121||RXNORM|BICYCLO(2.2.1)HEPTAN-2-AMINE, N-ETHYL-3-PHENYL-
C0060157|T121||RXNORM|FENCAMFAMINE
C0060157|T121||RXNORM|N-ETHYL-3-PHENYLBICYCLO(2.2.1)HEPTAN-2-AMINE
C0060157|T121||RXNORM|FENCAMFAMIN
C0060157|T121||RXNORM|2-NORBORNANAMINE, N-ETHYL-3-PHENYL-
C0060157|T121||RXNORM|3-PHENYL-N-ETHYL-2-NORBORNANAMINE
C0060157|T121||RXNORM|2-PHENYL-3-ETHYLAMINOBICYCLO(2.2.1)HEPTANE
C0060157|T121||RXNORM|2-ETHYLAMINO-3-PHENYLNORBORNANE
C0060157|T121||RXNORM|FENCAMFAMIN 
C1974051|T121||RXNORM|SULPIRIDE &#X7C; BLD-SER-PLAS
C1981573|T121||RXNORM|ANTIPSYCHOTICS &#X7C; BLD-SER-PLAS
C1980662|T121||RXNORM|ACETOPHENAZINE &#X7C; BLD-SER-PLAS
C0043513|T121|1535252|RXNORM|ZOLAZEPAM|ZOLAZEPAM
C0043513|T121|1535252|RXNORM|PYRAZOLO(3,4-E)(1,4)DIAZEPIN-7(1H)-ONE, 4-(2-FLUOROPHENYL)-6,8-DIHYDRO-1,3,8-TRIMETHYL-|ZOLAZEPAM
C0043513|T121|1535252|RXNORM|ZOLAZEPAM [CHEMICAL/INGREDIENT]|ZOLAZEPAM
C0043513|T121|1535252|RXNORM|ZOLASEPAM|ZOLAZEPAM
C1981247|T121||RXNORM|AMILSULPRIDE &#X7C; BLD-SER-PLAS
C0123091|T121|51272|RXNORM|QUETIAPINE|QUETIAPINE
C0123091|T121|51272|RXNORM|QUETIAPINE |QUETIAPINE
C0123091|T121|51272|RXNORM|2-(2-(4-DIBENZO(B,F)(1,4)THIAZEPINE-11-YL-1-PIPERAZINYL)ETHOXY)ETHANOL|QUETIAPINE
C0123091|T121|51272|RXNORM|QUETIAPINE |QUETIAPINE
C0123091|T121|51272|RXNORM|QUETIAPINE |QUETIAPINE
C0031436|T121||RXNORM|PHENOTHIAZINES
C0031436|T121||RXNORM|PHENOTHIAZINES 
C0031436|T121||RXNORM|PHENOTHIAZINES [CHEMICAL/INGREDIENT]
C1533126|T121|588250|RXNORM|CYCLOPROPANECARBOXAMIDE, 2-(AMINOMETHYL)-N,N-DIETHYL-1-PHENYL-, CIS-(+-)-|MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN|MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN |MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN |MILNACIPRAN
C1533126|T121|588250|RXNORM|MIDALCIPRAN|MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN [CHEMICAL/INGREDIENT]|MILNACIPRAN
C1533126|T121|588250|RXNORM|ANTIDEPRESSANTS SNRI MILNACIPRAN|MILNACIPRAN
C1533126|T121|588250|RXNORM|MILNACIPRAN |MILNACIPRAN
C2925168|T121||RXNORM|ILOPERIDONE &#X7C; BLD-SER-PLAS
C1994732|T121||RXNORM|PIPAMPERONE &#X7C; BLD-SER-PLAS
C1983134|T121||RXNORM|BROMPERIDOL &#X7C; BLD-SER-PLAS
C2925288|T121||RXNORM|METHOTRIMEPRAZINE METABOLITE &#X7C; URINE
C2738464|T121||RXNORM|NOROLANZAPINE &#X7C; BLD-SER-PLAS
C0770404|T121||RXNORM|CARPHENAZINE MALEATE
C0770404|T121||RXNORM|CARPHENAZINE MALEATE (DISCONTINUED) 
C0770404|T121||RXNORM|CARPHENAZINE MALEATE (DISCONTINUED)
C0770404|T121||RXNORM|CARPHENAZINE MALEATE 
C3847696|T121||RXNORM|FLUSPIRILENE &#X7C; BLD-SER-PLAS
C3871108|T121||RXNORM|ANTIPSYCHOTICS &#X7C; BLOOD OR URINE
C0299792|T121|89013|RXNORM|ARIPIPRAZOLE|ARIPIPRAZOLE
C0299792|T121|89013|RXNORM|2(1H)-QUINOLINONE, 7-(4-(4-(2,3-DICHLOROPHENYL)-1-PIPERAZINYL)BUTOXY)-3,4-DIHYDRO-|ARIPIPRAZOLE
C0299792|T121|89013|RXNORM|ARIPIPRAZOLE |ARIPIPRAZOLE
C0299792|T121|89013|RXNORM|7-(4-(4-(2,3-DICHLOROPHENYL)-1-PIPERAZINYL)BUTYLOXY)-3,4-DIHYDRO-2(1H)-QUINOLINONE|ARIPIPRAZOLE
C0299792|T121|89013|RXNORM|ARIPIPRAZOLE [CHEMICAL/INGREDIENT]|ARIPIPRAZOLE
C0299792|T121|89013|RXNORM|ARIPIPRAZOL|ARIPIPRAZOLE
C0299792|T121|89013|RXNORM|ARIPIPRAZOLE |ARIPIPRAZOLE
C0299792|T121|89013|RXNORM|ARIPIPRAZOLE |ARIPIPRAZOLE
C4038379|T121||RXNORM|7-HYDROXYQUETIAPINE &#X7C; URINE
C0724680|T121|221153|RXNORM|QUETIAPINE FUMARATE|QUETIAPINE FUMARATE
C0724680|T121|221153|RXNORM|ETHANOL, 2-(2-(4-DIBENZO(B,F)(1,4)THIAZEPIN-11-YL-1-PIPERAZINYL)ETHOXY)-,(E)-2-BUTENEDIOATE(2:1)(SALT)|QUETIAPINE FUMARATE
C0724680|T121|221153|RXNORM|FUMARATE, QUETIAPINE|QUETIAPINE FUMARATE
C0724680|T121|221153|RXNORM|ETHANOL, 2-(2-(4-DIBENZO(B,F)(1,4)THIAZEPIN-11-YL-1-PIPERAZINYL)ETHOXY)-, (E)-2-BUTENEDIOATE (2:1) (SALT)|QUETIAPINE FUMARATE
C0724680|T121|221153|RXNORM|QUETIAPINE FUMARATE [CHEMICAL/INGREDIENT]|QUETIAPINE FUMARATE
C0724680|T121|221153|RXNORM|QUETIAPINE FUMARATE |QUETIAPINE FUMARATE
C2697950|T121|1040027|RXNORM|LURASIDONE HYDROCHLORIDE|LURASIDONE HYDROCHLORIDE
C2697950|T121|1040027|RXNORM|LURASIDONE HYDROCHLORIDE |LURASIDONE HYDROCHLORIDE
C2697950|T121|1040027|RXNORM|HCL, LURASIDONE|LURASIDONE HYDROCHLORIDE
C2697950|T121|1040027|RXNORM|HYDROCHLORIDE, LURASIDONE|LURASIDONE HYDROCHLORIDE
C2697950|T121|1040027|RXNORM|LURASIDONE HCL|LURASIDONE HYDROCHLORIDE
C2697950|T121|1040027|RXNORM|LURASIDONE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|LURASIDONE HYDROCHLORIDE
C4072501|T121||RXNORM|BENPERIDOL &#X7C; BLD-SER-PLAS
C0103045|T121|46303|RXNORM|AMISULPRIDE|AMISULPRIDE
C0103045|T121|46303|RXNORM|AMISULPRIDE - CHEMICAL|AMISULPRIDE
C0103045|T121|46303|RXNORM|AMISULPRIDE |AMISULPRIDE
C0103045|T121|46303|RXNORM|AMISULPRIDE - CHEMICAL |AMISULPRIDE
C0103045|T121|46303|RXNORM|AMISULPRIDE |AMISULPRIDE
C4072058|T121||RXNORM|PENFLURIDOL &#X7C; BLD-SER-PLAS
C2003424|T121|1040028|RXNORM|LURASIDONE|LURASIDONE
C2003424|T121|1040028|RXNORM|N-(2-(4-(1,2-BENZISOTHIAZOL-3-YL)-1-PIPERAZINYLMETHYL)-1-CYCLOHEXYLMETHYL)-2,3-BICYCLO(2.2.1)HEPTANEDICARBOXIMIDE|LURASIDONE
C2003424|T121|1040028|RXNORM|LURASIDONE |LURASIDONE
C2003424|T121|1040028|RXNORM|LURASIDONE |LURASIDONE
C2003424|T121|1040028|RXNORM|ANTIPSYCHOTICS LURASIDONE|LURASIDONE
C4056439|T121|1673265|RXNORM|ARIPIPRAZOLE LAUROXIL|ARIPIPRAZOLE LAUROXIL
C4056439|T121|1673265|RXNORM|ANTIPSYCHOTICS ARIPIPRAZOLE LAUROXIL|ARIPIPRAZOLE LAUROXIL
C4056439|T121|1673265|RXNORM|ARIPIPRAZOLE LAUROXIL |ARIPIPRAZOLE LAUROXIL
C0358425|T121||RXNORM|ANXIOLYTICS AND NEUROLEPTIC PERIOPERATIVE DRUGS 
C0358425|T121||RXNORM|ANXIOLYTICS AND NEUROLEPTIC PERIOPERATIVE DRUGS
C0358425|T121||RXNORM|ANXIOLYTICS AND NEUROLEPTIC PERIOPERATIVE DRUGS 
C0030077|T121|7815|RXNORM|OXYPERTINE|OXYPERTINE
C0030077|T121|7815|RXNORM|1H-INDOLE, 5,6-DIMETHOXY-2-METHYL-3-(2-(4-PHENYL-1-PIPERAZINYL)ETHYL)-|OXYPERTINE
C0030077|T121|7815|RXNORM|5,6-DIMETHOXY-2-METHYL-3-(2-(4-PHENYL-1-PIPERAZINYL)ETHYL)INDOLE|OXYPERTINE
C0030077|T121|7815|RXNORM|WIN 18,501-2|OXYPERTINE
C0030077|T121|7815|RXNORM|OXYPERTINE |OXYPERTINE
C0030077|T121|7815|RXNORM|OXYPERTINE |OXYPERTINE
C0355185|T121||RXNORM|ANTIPSYCHOTIC DEPOT INJECTIONS 
C0355185|T121||RXNORM|ANTIPSYCHOTIC DEPOT INJECTIONS
C0355185|T121||RXNORM|ANTIPSYCHOTIC DEPOT INJECTIONS 
C0304387|T121||RXNORM|BUTYROPHENONE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304387|T121||RXNORM|BUTYROPHENONE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304387|T121||RXNORM|BUTYROPHENONE DERIVATIVE ANTIPSYCHOTIC AGENT
C0304387|T121||RXNORM|BUTYROPHENONE DERIVATIVE ANTIPSYCHOTIC AGENT, NOS
C0304389|T121||RXNORM|DIBENZOXAZEPINE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304389|T121||RXNORM|DIBENZOXAZEPINE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304389|T121||RXNORM|DIBENZOXAZEPINE DERIVATIVE ANTIPSYCHOTIC AGENT
C0304389|T121||RXNORM|DIBENZOXAZEPINE DERIVATIVE ANTIPSYCHOTIC AGENT, NOS
C0304392|T121||RXNORM|DIHYDROINDOLONE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304392|T121||RXNORM|DIHYDROINDOLONE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304392|T121||RXNORM|DIHYDROINDOLONE DERIVATIVE ANTIPSYCHOTIC AGENT
C0304392|T121||RXNORM|DIHYDROINDOLONE DERIVATIVE ANTIPSYCHOTIC AGENT, NOS
C0304393|T121||RXNORM|DIPHENYLBUTYLPIPERIDINE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304393|T121||RXNORM|DIPHENYLBUTYLPIPERIDINE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304393|T121||RXNORM|DIPHENYLBUTYLPIPERIDINE DERIVATIVE ANTIPSYCHOTIC AGENT
C0304393|T121||RXNORM|DIPHENYLBUTYLPIPERIDINE DERIVATIVE ANTIPSYCHOTIC AGENT, NOS
C1268911|T121||RXNORM|PHENYLBUTYLPIPERADINE DERIVATIVE ANTIPSYCHOTIC AGENT 
C1268911|T121||RXNORM|PHENYLBUTYLPIPERADINE DERIVATIVE ANTIPSYCHOTIC AGENT 
C1268911|T121||RXNORM|PHENYLBUTYLPIPERADINE DERIVATIVE ANTIPSYCHOTIC AGENT
C1276996|T121||RXNORM|ATYPICAL ANTIPSYCHOTIC
C1276996|T121||RXNORM|ATYPICAL ANTIPSYCHOTIC 
C1276996|T121||RXNORM|ATYPICAL ANTIPSYCHOTIC 
C0304383|T121||RXNORM|THIOXANTHENE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304383|T121||RXNORM|THIOXANTHENE DERIVATIVE ANTIPSYCHOTIC AGENT 
C0304383|T121||RXNORM|THIOXANTHENE DERIVATIVE ANTIPSYCHOTIC AGENT
C0304383|T121||RXNORM|THIOXANTHENE DERIVATIVE ANTIPSYCHOTIC AGENT, NOS
C1268910|T121||RXNORM|BENZISOXAZOLE DERIVATIVE ANTIPSYCHOTIC AGENT 
C1268910|T121||RXNORM|BENZISOXAZOLE DERIVATIVE ANTIPSYCHOTIC AGENT 
C1268910|T121||RXNORM|BENZISOXAZOLE DERIVATIVE ANTIPSYCHOTIC AGENT
C1320173|T121||RXNORM|DIHYDROCARBOSTYRIL DERIVATIVE ANTIPSYCHOTIC 
C1320173|T121||RXNORM|DIHYDROCARBOSTYRIL DERIVATIVE ANTIPSYCHOTIC AGENT 
C1320173|T121||RXNORM|DIHYDROCARBOSTYRIL DERIVATIVE ANTIPSYCHOTIC AGENT
C1320173|T121||RXNORM|DIHYDROCARBOSTYRIL DERIVATIVE ANTIPSYCHOTIC
C0100267|T121||RXNORM|8-HYDROXYLOXAPINE
C0100267|T121||RXNORM|DIBENZ(B,F)(1,4)OXAZEPIN-8-OL, 2-CHLORO-11-(4-METHYL-1-PIPERAZINYL)-
C0100267|T121||RXNORM|8-HYDROXYLOXAPINE 
C0304394|T121||RXNORM|DIMOZIDE
C0304394|T121||RXNORM|DIMOZIDE 
C0753678|T121|679314|RXNORM|PALIPERIDONE|PALIPERIDONE
C0753678|T121|679314|RXNORM|PALIPERIDONE |PALIPERIDONE
C0753678|T121|679314|RXNORM|PALIPERIDONE |PALIPERIDONE
C0753678|T121|679314|RXNORM|PALIPERIDONE |PALIPERIDONE
C0753678|T121|679314|RXNORM|9-HYDROXYRISPERIDONE|PALIPERIDONE
C0753678|T121|679314|RXNORM|4H-PYRIDO(1,2-A)PYRIMIDIN-4-ONE, 3-(2-(4-(6-FLUORO-1,2-BENZISOXAZOL-3-YL)-1-PIPERIDINYL)ETHYL)-6,7,8,9-TETRAHYDRO-9-HYDROXY-2-METHYL-|PALIPERIDONE
C0753678|T121|679314|RXNORM|9 HYDROXY RISPERIDONE|PALIPERIDONE
C0753678|T121|679314|RXNORM|9 OH RISPERIDONE|PALIPERIDONE
C0753678|T121|679314|RXNORM|9 HYDROXYRISPERIDONE|PALIPERIDONE
C0753678|T121|679314|RXNORM|9-HYDROXY-RISPERIDONE|PALIPERIDONE
C0753678|T121|679314|RXNORM|3-(2-(4-(6-FLUORO-3-(1,2-BENZISOXAZOLYL))-1-PIPERIDINYL)ETHYL)-6,7,8,9-TETRAHYDRO-9-HYDROXY-2-METHYL-4H-PYRIDO(1,2-A)PYRIMIDIN-4-ONE|PALIPERIDONE
C0753678|T121|679314|RXNORM|9-OH-RISPERIDONE|PALIPERIDONE
C0753678|T121|679314|RXNORM|9-HYDROXYRISPERIDONE |PALIPERIDONE
C0060473|T121||RXNORM|4'-FLUORO-4-(4-(O-METHOXYPHENYL)-1-PIPERAZINYL)- BUTYROPHENONE
C0060473|T121||RXNORM|FLUANISONE
C0060473|T121||RXNORM|HALOANISONE
C0060473|T121||RXNORM|HALOANIZONE
C0071098|T121|33739|RXNORM|1'-(3-(4-FLUOROBENZOYL)PROPYL)-(1,4'-BIPIPERIDINE) -4'-CARBOXAMIDE|PIPAMPERONE
C0071098|T121|33739|RXNORM|PIPAMPERONE|PIPAMPERONE
C0071098|T121|33739|RXNORM|PIPAMPERONE |PIPAMPERONE
C0071098|T121|33739|RXNORM|PIPAMPERONE |PIPAMPERONE
C0066477|T121|29961|RXNORM|4'-FLUOR-4-(4-METHYLPIPERIDINO)-BUTYROPHENONE|MELPERONE
C0066477|T121|29961|RXNORM|MELPERON|MELPERONE
C0066477|T121|29961|RXNORM|MELPERONE|MELPERONE
C0066477|T121|29961|RXNORM|METHYLPERON|MELPERONE
C0066477|T121|29961|RXNORM|METYLPERON|MELPERONE
C0066477|T121|29961|RXNORM|MELPERONE |MELPERONE
C0066477|T121|29961|RXNORM|MELPERONE |MELPERONE
C0075226|T121||RXNORM|STEPHOLIDINE
C0075630|T121|37416|RXNORM|N-(ETHYL-1-PYRROLIDINYL- 2-METHYL)METHOXY-2-ETHYLSULFONYL-5-BENZAMIDE|SULTOPRIDE
C0075630|T121|37416|RXNORM|SULTOPRIDE|SULTOPRIDE
C0075630|T121|37416|RXNORM|N-((1-ETHYL-2-PYRROLIDINYL)METHYL)-5-(ETHYLSULFONYL)-O-ANISAMIDE|SULTOPRIDE
C0074587|T121||RXNORM|2,6-METHANO-3-BENZAZOCIN-8-OL, 1,2,3,4,5,6-HEXAHYDRO-6,11-DIMETHYL-3-(2-PROPENYL)-
C0074587|T121||RXNORM|SK&F 10047
C0074587|T121||RXNORM|SKF 10047
C0074587|T121||RXNORM|SKF-10047
C0058518|T121||RXNORM|10-(2-METHYL 3-(1-HYDROXYETHOXYETHYL-4-PIPERAZINYL)PROPYL)PHENOTHIAZINE
C0058518|T121||RXNORM|DIXYRAZINE
C0076278|T121||RXNORM|5,8,13,13A-TETRAHYDRO-2,3,9,10-TETRAMETHOXY-6H-DIBENZO(A,G)QUINOLIZINE
C0076278|T121||RXNORM|TETRAHYDROPALMATINE
C0076278|T121||RXNORM|TETRAHYDROPALMITINE
C0071053|T121||RXNORM|6-FLUORO-9-(3-(4-(2-HYDROXYETHYL)PIPERIDINO) PROPYLIDENE)-2-TRIFLUOROMETHYL-THIOXANTHENE
C0071053|T121||RXNORM|PIFLUTIXOL
C0063970|T121||RXNORM|1-PIPERAZINEETHANOL, 4-(3-FLUORO-10,11-DIHYDRO-8-(1-METHYLETHYL)DIBENZO(B,F)THIEPIN-10-YL)-
C0063970|T121||RXNORM|3-FLUOR-8-ISOPROPYL-10-(4-(2-HYDROXYETHYL)PIPERAZINO)-10,11-DIHYDRODIBENZO(B,F)THIEPIN
C0063970|T121||RXNORM|ISOFLOXYTHEPIN
C0078849|T121|40003|RXNORM|2-CHLORO-11-(2-DIMETHYLAMINOETHOXY)DIBENZO(B,F)THIEPINE|ZOTEPINE
C0078849|T121|40003|RXNORM|ZOTEPINE|ZOTEPINE
C0078849|T121|40003|RXNORM|2-((8-CHLORODIBENZO(B,F)THIEPIN-10-YL)OXY)-N,N-DIMETHYLETHANAMINE|ZOTEPINE
C0078849|T121|40003|RXNORM|ZOTEPINE |ZOTEPINE
C0078849|T121|40003|RXNORM|ZOTEPINE |ZOTEPINE
C0076688|T121||RXNORM|4'-FLUORO-4-(4-(2-THIOXO-1-BENZIMIDAZOLINYL)PIPERIDINO)BUTYROPHENONE
C0076688|T121||RXNORM|4-(4-(2,3-DIHYDRO-2-THIOXO-1H-BENZIMIDAZOL-1-YL)-1-PIPERIDINYL)-1-(4-FLUOROPHENYL)-1- BUTANONE
C0076688|T121||RXNORM|TIMIPERONE
C0078761|T121||RXNORM|1-(3-CHLOROPHENYL)-3-(2-(3,3-DIMETHYL-1-AZETIDINYL)ETHYL)IMIDAZOLIDIN-2-ONE
C0078761|T121||RXNORM|2-IMIDAZOLIDINONE, 1-(3-CHLOROPHENYL)-3-(2-(3,3-DIMETHYL-1-AZETIDINYL)ETHYL)-
C0078761|T121||RXNORM|ZETIDOLINE
C0055929|T121||RXNORM|CLOPENTHIXOL DECANOATE
C0055929|T121||RXNORM|CLOPENTIXOL DECANOATE
C0058537|T121||RXNORM|DN 1417
C0058537|T121||RXNORM|DN-1417
C0058537|T121||RXNORM|L-PROLINAMIDE, N-((TETRAHYDRO-5-OXO-2-FURANYL)CARBONYL)-L-HISTIDYL-
C0217937|T121||RXNORM|BENZAMIDE, 5-CHLORO-2-METHOXY-4-(METHYLAMINO)-N-(2-METHYL-1-(PHENYLMETHYL)-3-PYRROLIDINYL)-
C0217937|T121||RXNORM|NEMONAPRIDE
C0073502|T121||RXNORM|4H-PYRROLO(2,3-G)ISOQUINOLIN-4-ONE, 3-ETHYL-1,4A,5,6,7,8,8A,9-OCTAHYDRO-2,6-DIMETHYL-, TRANS-(+-)-
C0073502|T121||RXNORM|RO 22-1319
C0073502|T121||RXNORM|RO-22-1319
C0062103|T121|26420|RXNORM|HALOPERIDOL DECANOATE|HALOPERIDOL DECANOATE
C0062103|T121|26420|RXNORM|HALOPERIDOL DECONOATE|HALOPERIDOL DECANOATE
C0062103|T121|26420|RXNORM|HALOPERIDOL DECANOATE (DISCONTINUED) |HALOPERIDOL DECANOATE
C0062103|T121|26420|RXNORM|HALOPERIDOL DECANOATE (DISCONTINUED)|HALOPERIDOL DECANOATE
C0062103|T121|26420|RXNORM|HALOPERIDOL DECANOATE [CHEMICAL/INGREDIENT]|HALOPERIDOL DECANOATE
C0062103|T121|26420|RXNORM|HALOPERIDOL DECANOATE |HALOPERIDOL DECANOATE
C0062103|T121|26420|RXNORM|HALOPERIDOL DECANOATE |HALOPERIDOL DECANOATE
C0062103|T121|26420|RXNORM|HALOPERIDOL DECONOATE |HALOPERIDOL DECANOATE
C0140593|T121||RXNORM|CIS-9-(3-(3,5-DIMETHYL-1-PIPERAZINYL)PROPYL)CARBAZOLE
C0140593|T121||RXNORM|RIMCAZOLE
C0057143|T121|22298|RXNORM|1,2,4-TRIAZOLO(4,3-A)PYRIDINE, 5,6,7,8-TETRAHYDRO-3-(2-(4-(2-METHYLPHENYL)-1-PIPERAZINYL)ETHYL)-|DAPIPRAZOLE
C0057143|T121|22298|RXNORM|DAPIPRAZOLE|DAPIPRAZOLE
C0057143|T121|22298|RXNORM|DAPIPRAZOLE [CHEMICAL/INGREDIENT]|DAPIPRAZOLE
C0057143|T121|22298|RXNORM|DAPIPRAZOLE |DAPIPRAZOLE
C0057143|T121|22298|RXNORM|DAPIPRAZOLE |DAPIPRAZOLE
C0060579|T121||RXNORM|3-FLUORO-6-(4-METHYLPIPERAZINYL)-11H-DIBENZ(B,E)AZEPINE
C0060579|T121||RXNORM|FLUPERLAPINE
C0051747|T121||RXNORM|AMPEROZIDE
C1099053|T121||RXNORM|ECOPIPAM
C1099053|T121||RXNORM|5H-BENZO(D)NAPHTH(2,1-B)AZEPIN-12-OL, 11-CHLORO-6,6A,7,8,9,13B-HEXAHYDRO-7-METHYL-, TRANS-(-)-
C0378456|T121||RXNORM|3,4,4A,10B-TETRAHYDRO-4-PROPYL-2H,5H-(1)BENZOPYRANO(4,3-B)-1,4-OXAZIN-9-OL
C0378456|T121||RXNORM|PBPO
C0378456|T121||RXNORM|PBTO
C0084572|T121||RXNORM|2-(4-(4-(1,2-BENZISOTHIAZOL-3-YL)-1-PIPERAZINYL)BUTYL)HEXAHYDRO-1H-ISOINDOLE-1,3-(2H)-DIONE
C0084572|T121||RXNORM|PEROSPIRONE
C0084528|T121|41996|RXNORM|1-(2-(4-(5-CHLORO-1-(4-FLUOROPHENYL)-1H-INDOL-3-YL)-1-PIPERIDINYL)ETHYL)-2-IMIDAZOLIDINONE|SERTINDOLE
C0084528|T121|41996|RXNORM|SERTINDOLE|SERTINDOLE
C0084528|T121|41996|RXNORM|SERTINDOLE |SERTINDOLE
C0084528|T121|41996|RXNORM|SERTINDOLE [CHEMICAL/INGREDIENT]|SERTINDOLE
C0084528|T121|41996|RXNORM|SERTINDOLE |SERTINDOLE
C0084528|T121|41996|RXNORM|SERTINDOLE |SERTINDOLE
C0526908|T121||RXNORM|2-(3-(4-(4-FLUOROPHENYL)-1-PIPERAZINYL)PROPYL)-2H-NAPHTH(1,8-CD)ISOTHIAZOLE 1,1-DIOXIDE
C0526908|T121||RXNORM|FANANSERIN
C0526908|T121||RXNORM|FANANSERINE
C0211640|T121||RXNORM|DUP-734
C0211640|T121||RXNORM|ETHANONE, 2-(1-(CYCLOPROPYLMETHYL)-4-PIPERIDINYL)-1-(4-FLUOROPHENYL)-, HYDROBROMIDE
C0211640|T121||RXNORM|DUP 734
C0248068|T121||RXNORM|BENZENEETHANAMINE, 4-METHOXY-3-(2-PHENYLETHOXY)-N,N-DIPROPYL-, HYDROCHLORIDE
C0248068|T121||RXNORM|N,N-DIPROPYL-2-(4-METHOXY-3-(2-PHENYLETHOXY)PHENYL)ETHYLAMINE MONOHYDROCHLORIDE
C0293258|T121||RXNORM|SR 142801
C0293258|T121||RXNORM|SR-142801
C0293258|T121||RXNORM|SR142801
C0389977|T121||RXNORM|3-((4-(4-CHLOROPHENYL)PIPERAZIN-1-YL)METHYL)-1H-PYRROLO(2,3-B)PYRIDINE
C0389977|T121||RXNORM|CPMPP-3
C0057820|T121||RXNORM|2,3,4,4A,5,9B-HEXAHYDRO-2,8-DIMETHYL-1H-PYRIDO(4,3-B)INDOLE
C0057820|T121||RXNORM|CARBIDINE
C0057820|T121||RXNORM|DICARBINE
C0057820|T121||RXNORM|1H-PYRIDO(4,3-B)INDOLE, 2,3,4,4A,5,9B-HEXAHYDRO-2,8-DIMETHYL-
C1443761|T121||RXNORM|BENZIMIDAZOLINONE DERIVATIVE ANTIPSYCHOTIC PREPARATION 
C1443761|T121||RXNORM|BENZIMIDAZOLINONE DERIVATIVE ANTIPSYCHOTIC PREPARATION
C1443762|T121||RXNORM|BENZIMIDAZOLINONE DERIVATIVE ANTIPSYCHOTIC AGENT 
C1443762|T121||RXNORM|BENZIMIDAZOLINONE DERIVATIVE ANTIPSYCHOTIC AGENT
C0031434|T121||RXNORM|PHENOTHIAZINE
C0031434|T121||RXNORM|PHENOSAN
C0031434|T121||RXNORM|PHENOTHIAZINE 
C0031434|T121||RXNORM|THIODIPHENYLAMINE
C0031434|T121||RXNORM|PHENOTHIAZINE 
C0031434|T121||RXNORM|PHENOTHIAZINE, NOS
C0060580|T121|25190|RXNORM|FLUPHENAZINE DECANOATE|FLUPHENAZINE DECANOATE
C0060580|T121|25190|RXNORM|FLUPHENAZINE DEPOT|FLUPHENAZINE DECANOATE
C0060580|T121|25190|RXNORM|FTORPHENAZINE DECANOATE|FLUPHENAZINE DECANOATE
C0060580|T121|25190|RXNORM|FLUFENAZINE DECANOATE|FLUPHENAZINE DECANOATE
C0060580|T121|25190|RXNORM|FLUPHENAZINE DECANOATE |FLUPHENAZINE DECANOATE
C0060580|T121|25190|RXNORM|FLUPHENAZINE DEPOT [CHEMICAL/INGREDIENT]|FLUPHENAZINE DECANOATE
C0060580|T121|25190|RXNORM|FLUOPHENAZINE DECANOATE|FLUPHENAZINE DECANOATE
C0060580|T121|25190|RXNORM|FLUOPHENAZINE DECANOATE |FLUPHENAZINE DECANOATE
C0060580|T121|25190|RXNORM|FLUPHENAZINE DECANOATE |FLUPHENAZINE DECANOATE
C0060580|T121|25190|RXNORM|FLUPHENAZINE DECANOATE |FLUPHENAZINE DECANOATE
C0304386|T121|91135|RXNORM|THIOTHIXENE HYDROCHLORIDE|THIOTHIXENE HYDROCHLORIDE
C0304386|T121|91135|RXNORM|CP 12252-1|THIOTHIXENE HYDROCHLORIDE
C0304386|T121|91135|RXNORM|9H-THIOXANTHENE-2-SULFONAMIDE, N,N-DIMETHYL-9-(3-(4-METHYL-1-PIPERAZINYL)PROPYLIDENE)-, DIHYDROCHLORIDE, DIHYDRATE|THIOTHIXENE HYDROCHLORIDE
C0304386|T121|91135|RXNORM|ANTIPSYCHOTICS THIOTHIXENE HYDROCHLORIDE|THIOTHIXENE HYDROCHLORIDE
C0304386|T121|91135|RXNORM|THIOTHIXENE HYDROCHLORIDE |THIOTHIXENE HYDROCHLORIDE
C0304386|T121|91135|RXNORM|THIOTHIXENE HYDROCHLORIDE |THIOTHIXENE HYDROCHLORIDE
C0304386|T121|91135|RXNORM|TIOTIXENE HYDROCHLORIDE|THIOTHIXENE HYDROCHLORIDE
C1170754|T121|353116|RXNORM|ZIPRASIDONE MESYLATE|ZIPRASIDONE MESYLATE
C1170754|T121|353116|RXNORM|ZIPRASIDONE MESYLATE |ZIPRASIDONE MESYLATE
C1170754|T121|353116|RXNORM|ZIPRASIDONE MESYLATE |ZIPRASIDONE MESYLATE
C0242518|T121|71529|RXNORM|THIETHYLPERAZINE MALEATE|THIETHYLPERAZINE MALATE
C0242518|T121|71529|RXNORM|THIETHYLPERAZINE MALATE|THIETHYLPERAZINE MALATE
C0242518|T121|71529|RXNORM|THIETHYLPERAZINE MALATE (DISCONTINUED)|THIETHYLPERAZINE MALATE
C0242518|T121|71529|RXNORM|THIETHYLPERAZINE MALATE (DISCONTINUED) |THIETHYLPERAZINE MALATE
C0242518|T121|71529|RXNORM|THIETHYLPERAZINE MALEATE |THIETHYLPERAZINE MALATE
C0242518|T121|71529|RXNORM|THIETHYLPERAZINE MALATE [CHEMICAL/INGREDIENT]|THIETHYLPERAZINE MALATE
C0242518|T121|71529|RXNORM|10H-PHENOTHIAZINE, 2-(ETHYLTHIO)-10-(3-(4-METHYL-1-PIPERAZINYL)PROPYL)-, (Z)-2-BUTENEDIOATE|THIETHYLPERAZINE MALATE
C0242518|T121|71529|RXNORM|THIETHYLPERAZINE MALATE |THIETHYLPERAZINE MALATE
C0242518|T121|71529|RXNORM|THIETHYLPERAZINE MALEATE |THIETHYLPERAZINE MALATE
C0033473|T121|8770|RXNORM|PROPIOMAZINE|PROPIOMAZINE
C0033473|T121|8770|RXNORM|1-PROPANONE, 1-(10-(2-(DIMETHYLAMINO)PROPYL)-10H-PHENOTHIAZIN-2-YL)-|PROPIOMAZINE
C0033473|T121|8770|RXNORM|DROPIOMAZINE|PROPIOMAZINE
C0033473|T121|8770|RXNORM|PROPIOMAZINE -RETIRED-|PROPIOMAZINE
C0033473|T121|8770|RXNORM|PROPIOMAZINE [CHEMICAL/INGREDIENT]|PROPIOMAZINE
C0033473|T121|8770|RXNORM|PROPIOMAZINE |PROPIOMAZINE
C0033473|T121|8770|RXNORM|PROPIOMAZINE |PROPIOMAZINE
C1721449|T121||RXNORM|BIFEPRUNOX
C1721449|T121||RXNORM|1-(2-OXO-BENZOXAZOLIN-7-YL)-4-(3-BIPHENYL)METHYLPIPERAZINEMESYLATE
C0601644|T121||RXNORM|IMICLOPAZINE
C0601644|T121||RXNORM|1-(2-(4-(3-(2-CHLORO-10H-PHENOTHIAZIN-10-YL)PROPYL)-1-PIPERAZINYL)ETHYL)-3- METHYL-2-IMIDAZOLIDINONE
C0601644|T121||RXNORM|1-(2-(3-(2-CHLOROPHENOTHIAZIN- 10-YL)PROPYL)-1-PIPERAZINYLETHYL)-3-METHYL-2- IMIDAZOLIDINONE
C0601644|T121||RXNORM|CHLORIMIPHENINE
C1883076|T121||RXNORM|SPICLOMAZINE
C0125997|T121|52105|RXNORM|LITHIUM CITRATE|LITHIUM CITRATE
C0125997|T121|52105|RXNORM|LITHIUM CITRATE |LITHIUM CITRATE
C0125997|T121|52105|RXNORM|LITHIUM (AS CITRATE)|LITHIUM CITRATE
C0125997|T121|52105|RXNORM|LITHIUM CITRATE [CHEMICAL/INGREDIENT]|LITHIUM CITRATE
C0125997|T121|52105|RXNORM|LITHIUM CITRATE |LITHIUM CITRATE
C0125997|T121|52105|RXNORM|LITHIUM CITRATE |LITHIUM CITRATE
C0024057|T121|6476|RXNORM|LOXAPINE SUCCINATE|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|BUTANEDIOIC ACID, COMPOUND WITH 2-CHLORO-11-(4-METHYL-1-PIPERAZINYL)DIBENZ(B,F)(1,4)OXAZEPINE(1:1)|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|2-CHLORO-11-(4-METHYL-1-PIPERAZINYL)DIBENZ(B,F)(1,4)OXAZEPINE SUCCINATE(1:1)|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|CLOXAZEPIN|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|LOXAPINE SUCCINATE |LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|LOXAPINSUCCINATE|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|DAXOLIN|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|SUCCINATE, LOXAPINE|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|LOXAPINE SUCCINATE [CHEMICAL/INGREDIENT]|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|LOXIPINE SUCCINATE|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|OXILAPINE SUCCINATE|LOXAPINE SUCCINATE
C0024057|T121|6476|RXNORM|LOXAPINE SUCCINATE |LOXAPINE SUCCINATE
C1880734|T121||RXNORM|FARAMPATOR
C1880823|T121||RXNORM|FLUSPIPERONE
C0065505|T121||RXNORM|4'-((3-(4-(2-FLUOROPHENYL)-1-PIPERAZINYL)PROPYL)OXY)-3'-METHOXYACETANILIDE
C0065505|T121||RXNORM|MAFOPRAZINE
C0700543|T121|203186|RXNORM|MESORIDAZINE BESYLATE|MESORIDAZINE BESYLATE
C0700543|T121|203186|RXNORM|MESORIDAZINE BENZENESULPHONATE|MESORIDAZINE BESYLATE
C0700543|T121|203186|RXNORM|MESORIDAZINE BENZENESULFONATE|MESORIDAZINE BESYLATE
C0700543|T121|203186|RXNORM|MESORIDAZINE BESYLATE |MESORIDAZINE BESYLATE
C0301379|T121||RXNORM|MEBUTAMATE
C0301379|T121||RXNORM|MEBUTAMATE (DISCONTINUED)
C0301379|T121||RXNORM|MEBUTAMATE (DISCONTINUED) 
C0301379|T121||RXNORM|MEBUTAMATE 
C0013015|T121|3626|RXNORM|DOMPERIDONE|DOMPERIDONE
C0013015|T121|3626|RXNORM|2H-BENZIMIDAZOL-2-ONE, 5-CHLORO-1-(1-(3-(2,3-DIHYDRO-2-OXO-1H-BENZIMIDAZOL-1-YL)PROPYL)-4-PIPERIDINYL)-1,3-DIHYDRO-|DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDON|DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDONE [CHEMICAL/INGREDIENT]|DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDONE(MOTILITY) [SEE CHAPTER D FOR PREPARATIONS] |DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDONE(MOTILITY) [SEE CHAPTER D FOR PREPARATIONS]|DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDONE [NAUSEA]|DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDONE [NAUSEA] |DOMPERIDONE
C0013015|T121|3626|RXNORM|GI PROKINETIC MOTILITY AGENTS DOMPERIDONE |DOMPERIDONE
C0013015|T121|3626|RXNORM|GI PROKINETIC MOTILITY AGENTS DOMPERIDONE|DOMPERIDONE
C0013015|T121|3626|RXNORM|ANTINAUSEANTS DOMPERIDONE |DOMPERIDONE
C0013015|T121|3626|RXNORM|ANTINAUSEANTS DOMPERIDONE|DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDONE |DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDONE |DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDONE [NAUSEA] |DOMPERIDONE
C0013015|T121|3626|RXNORM|DOMPERIDONE(MOTILITY) [SEE CHAPTER D FOR PREPARATIONS] |DOMPERIDONE
C1880846|T121||RXNORM|FOSENAZIDE
C0546875|T121|142444|RXNORM|HYDROCHLORIDE, PROMAZINE|PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|PROMAZINE HYDROCHLORIDE|PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|STARAZIN|PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|TALOFEN|PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|10-(3-(DIMETHYLAMINO)PROPYL)PHENOTHIAZINE MONOHYDROCHLORIDE|PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|10H-PHENOTHIAZINE-10-PROPANAMINE, N,N-DIMETHYL-, MONOHYDROCHLORIDE|PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|PROMAZINE HYDROCHLORIDE (DISCONTINUED) |PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|ANTIPSYCHOTICS PROMAZINE HYDROCHLORIDE (DISCONTINUED)|PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|PROMAZINE HYDROCHLORIDE (DISCONTINUED)|PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|PROMAZINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|PROMAZINE HYDROCHLORIDE |PROMAZINE HYDROCHLORIDE
C0546875|T121|142444|RXNORM|PROMAZINE HYDROCHLORIDE [DUP] |PROMAZINE HYDROCHLORIDE
C0085217|T121|42351|RXNORM|CARBONATE, LITHIUM|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|CARBONATE, DILITHIUM|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|CARBONIC ACID, DILITHIUM SALT|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE |LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE [CHEMICAL/INGREDIENT]|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|DILITHIUM CARBONATE|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE PREPARATION|LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE |LITHIUM CARBONATE
C0085217|T121|42351|RXNORM|LITHIUM CARBONATE |LITHIUM CARBONATE
C0023044|T121|6232|RXNORM|PROPIOMAZINE HYDROCHLORIDE|PROPIOMAZINE HYDROCHLORIDE
C0023044|T121|6232|RXNORM|PROPIOMAZINE HYDROCHLORIDE |PROPIOMAZINE HYDROCHLORIDE
C0066492|T121||RXNORM|2-METHYLAMINO-4-N-METHYLPIPERAZINO-5-THIOMETHYL-6-CHLOROPYRIMIDINE
C0066492|T121||RXNORM|2-PYRIDINAMINE, 4-CHLORO-N-METHYL-6-(4-METHYL-1-PIPERAZINYL)-5-(METHYLTHIO)-
C0066492|T121||RXNORM|MEZILAMINE
C0075006|T121||RXNORM|8-(3-(4-FLUOROPHENOXY)PROPYL)-1-PHENYL-1,3,8-TRIAZASPIRO(4.5)DECAN-4-ONE
C0075006|T121||RXNORM|SPIRAMIDE
C0075006|T121||RXNORM|8-(3-(4-FLUOROPHENOXY) PROPYL)-1-PHENYL-1,3,8-TRIAZASPIRO(4, 5)DECAN-4-ONE
C0058805|T121||RXNORM|(4-FLUOROPHENYL)(1-(3-(2-(TRIFLUOROMETHYL)-10H-PHENOTHIAZINE-10-YL)PROPYL)-4-PIPERIDINYL)METHANONE
C0058805|T121||RXNORM|DUOPERONE
C0304376|T121|91125|RXNORM|TRIFLUPROMAZINE HYDROCHLORIDE|TRIFLUPROMAZINE HYDROCHLORIDE
C0304376|T121|91125|RXNORM|TRIFLUPROMAZINE HYDROCHLORIDE (DISCONTINUED) |TRIFLUPROMAZINE HYDROCHLORIDE
C0304376|T121|91125|RXNORM|ANTIPSYCHOTICS TRIFLUPROMAZINE HYDROCHLORIDE (DISCONTINUED)|TRIFLUPROMAZINE HYDROCHLORIDE
C0304376|T121|91125|RXNORM|TRIFLUPROMAZINE HYDROCHLORIDE (DISCONTINUED)|TRIFLUPROMAZINE HYDROCHLORIDE
C0304376|T121|91125|RXNORM|TRIFLUPROMAZINE HYDROCHLORIDE |TRIFLUPROMAZINE HYDROCHLORIDE
C0663536|T121||RXNORM|PANAMESINE
C0663536|T121||RXNORM|(5S)-5-((4-HYDROXY-4-(3,4-(METHYLENEDIOXY)PHENYL)PIPERIDINO)METHYL)-3-(P-METHOXYPHENYL)-2-OXAZOLIDINONE
C0282249|T121|82051|RXNORM|HYDROCHLORIDE, MOLINDONE|MOLINDONE HYDROCHLORIDE
C0282249|T121|82051|RXNORM|MOLINDONE HYDROCHLORIDE|MOLINDONE HYDROCHLORIDE
C0282249|T121|82051|RXNORM|4H-INDOL-4-ONE, 3-ETHYL-1,5,6,7-TETRAHYDRO-2-METHYL-5-(4-MORPHOLINYLMETHYL)-, MONOHYDROCHLORIDE|MOLINDONE HYDROCHLORIDE
C0282249|T121|82051|RXNORM|LIDONE|MOLINDONE HYDROCHLORIDE
C0282249|T121|82051|RXNORM|MOLINDONE HYDROCHLORIDE |MOLINDONE HYDROCHLORIDE
C0282249|T121|82051|RXNORM|MOLINDONE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|MOLINDONE HYDROCHLORIDE
C0282249|T121|82051|RXNORM|MOLINDONE MONOHYDROCHLORIDE|MOLINDONE HYDROCHLORIDE
C0282249|T121|82051|RXNORM|MONOHYDROCHLORIDE, MOLINDONE|MOLINDONE HYDROCHLORIDE
C0282249|T121|82051|RXNORM|MOLINDONE HYDROCHLORIDE |MOLINDONE HYDROCHLORIDE
C0386741|T121||RXNORM|4-AMINO-2-BUTOXY-5-CHLORO-N-(1-(1,3-DIOXOLAN-2-YLMETHYL)PIPERID-4-YL)BENZAMIDE
C0386741|T121||RXNORM|DOBUPRIDE
C0376160|T121|114176|RXNORM|ZUCLOPENTHIXOL|ZUCLOPENTHIXOL
C0376160|T121|114176|RXNORM|ZUCLOPENTHIXOL |ZUCLOPENTHIXOL
C0376160|T121|114176|RXNORM|ZUCLOPENTHIXOL |ZUCLOPENTHIXOL
C0376160|T121|114176|RXNORM|CLOPENTIXOL CIS-(Z)-|ZUCLOPENTHIXOL
C0376160|T121|114176|RXNORM|(Z)-4-(3-(2-CHLOROTHIOXANTHEN-9-YLIDENE)PROPYL)-1-PIPERAZINEETHANOL|ZUCLOPENTHIXOL
C0376160|T121|114176|RXNORM|ALPHA-CLOPENTHIXOL|ZUCLOPENTHIXOL
C0376160|T121|114176|RXNORM|ALPHA CLOPENTHIXOL|ZUCLOPENTHIXOL
C1882247|T121||RXNORM|OXYPENDYL
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE|CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|2-CHLORO-10-(3-(DIMETHYLAMINO)PROPYL)PHENOTHIAZINE MONOHYDROCHLORIDE|CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE |CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|HYDROCHLORIDE, CHLORPROMAZINE|CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE (OBSOLETE)|CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE [ANESTHESIA]|CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE [ANESTHESIA] |CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE |CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE [NAUSEA] [SEE DH2..]|CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE [NAUSEA] [SEE DH2..] |CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE [ANAESTHESIA]|CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE |CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE [ANESTHESIA] |CHLORPROMAZINE HYDROCHLORIDE
C0355077|T121|104728|RXNORM|CHLORPROMAZINE HYDROCHLORIDE [NAUSEA] [SEE DH2..] |CHLORPROMAZINE HYDROCHLORIDE
C0031954|T121|8338|RXNORM|PIPERACETAZINE|PIPERACETAZINE
C0031954|T121|8338|RXNORM|1-(10-(3-(4-(2-HYDROXYETHYL)-1-PIPERIDINYL)PROPYL)-10H-PHENOTHIAZIN-2-YL)ETHANONE|PIPERACETAZINE
C0031954|T121|8338|RXNORM|PIPERACETAZINE (DISCONTINUED)|PIPERACETAZINE
C0031954|T121|8338|RXNORM|PIPERACETAZINE (DISCONTINUED) |PIPERACETAZINE
C0031954|T121|8338|RXNORM|PIPERACETAZINE [CHEMICAL/INGREDIENT]|PIPERACETAZINE
C0031954|T121|8338|RXNORM|PIPERACETAZINE |PIPERACETAZINE
C0304378|T121|91127|RXNORM|ACETOPHENAZINE MALEATE|ACETOPHENAZINE MALEATE
C0304378|T121|91127|RXNORM|ACETOPHENAZINE MALEATE (DISCONTINUED)|ACETOPHENAZINE MALEATE
C0304378|T121|91127|RXNORM|ACETOPHENAZINE MALEATE (DISCONTINUED) |ACETOPHENAZINE MALEATE
C0304378|T121|91127|RXNORM|ACETOPHENAZINE MALEATE |ACETOPHENAZINE MALEATE
C1880547|T121||RXNORM|ERIZEPINE
C1881437|T121||RXNORM|LOFENDAZAM
C0070425|T121||RXNORM|1-(3-(2-METHOXYPHENOTHIAZIN-10-YL)-2-METHYLPROPYL)-4-PIPERIDINOL
C0070425|T121||RXNORM|PERIMETAZINE
C0304381|T121|91130|RXNORM|TRIFLUOPERAZINE HYDROCHLORIDE|TRIFLUOPERAZINE HYDROCHLORIDE
C0304381|T121|91130|RXNORM|TRIFLUOPERAZINE DIHYDROCHLORIDE|TRIFLUOPERAZINE HYDROCHLORIDE
C0304381|T121|91130|RXNORM|10-(3-(4-METHYL-1-PIPERAZINYL)PROPYL)-2-(TRIFLUOROMETHYL)-10H-PHENOTHIAZINE DIHYDROCHLORIDE|TRIFLUOPERAZINE HYDROCHLORIDE
C0304381|T121|91130|RXNORM|TRIFLUOPERAZINE HYDROCHLORIDE |TRIFLUOPERAZINE HYDROCHLORIDE
C0304381|T121|91130|RXNORM|ANTIPSYCHOTICS TRIFLUOPERAZINE HYDROCHLORIDE|TRIFLUOPERAZINE HYDROCHLORIDE
C0304381|T121|91130|RXNORM|TRIFLUOPERAZINE HCL|TRIFLUOPERAZINE HYDROCHLORIDE
C0304381|T121|91130|RXNORM|TRIFLUOPERAZINE HYDROCHLORIDE |TRIFLUOPERAZINE HYDROCHLORIDE
C0304381|T121|91130|RXNORM|TRIFLUOPERAZINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|TRIFLUOPERAZINE HYDROCHLORIDE
C0304381|T121|91130|RXNORM|TRIFLUOPERAZINE HYDROCHLORIDE |TRIFLUOPERAZINE HYDROCHLORIDE
C0700499|T121|203165|RXNORM|THIORIDAZINE HYDROCHLORIDE|THIORIDAZINE HYDROCHLORIDE
C0700499|T121|203165|RXNORM|THIORIDAZINE HYDROCHLORIDE |THIORIDAZINE HYDROCHLORIDE
C0700499|T121|203165|RXNORM|ANTIPSYCHOTICS THIORIDAZINE HYDROCHLORIDE|THIORIDAZINE HYDROCHLORIDE
C0700499|T121|203165|RXNORM|THIORIDAZINE HCL|THIORIDAZINE HYDROCHLORIDE
C0700499|T121|203165|RXNORM|THIORIDAZINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|THIORIDAZINE HYDROCHLORIDE
C0700499|T121|203165|RXNORM|THIORIDAZINE HYDROCHLORIDE |THIORIDAZINE HYDROCHLORIDE
C0700499|T121|203165|RXNORM|THIORIDAZINE HYDROCHLORIDE [DUP] |THIORIDAZINE HYDROCHLORIDE
C0700567|T121|203207|RXNORM|HYDROCHLORIDE, FLUPHENAZINE|FLUPHENAZINE HYDROCHLORIDE
C0700567|T121|203207|RXNORM|FLUPHENAZINE HYDROCHLORIDE|FLUPHENAZINE HYDROCHLORIDE
C0700567|T121|203207|RXNORM|FLUPHENAZINE HYDROCHLORIDE |FLUPHENAZINE HYDROCHLORIDE
C0700567|T121|203207|RXNORM|FLUPHENAZINE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|FLUPHENAZINE HYDROCHLORIDE
C0700567|T121|203207|RXNORM|FLUPHENAZINE HYDROCHLORIDE |FLUPHENAZINE HYDROCHLORIDE
C0700567|T121|203207|RXNORM|FLUPHENAZINE HYDROCHLORIDE [DUP] |FLUPHENAZINE HYDROCHLORIDE
C0062101|T121||RXNORM|HALOPEMIDE
C0062101|T121||RXNORM|N-(2-(4-(5-CHLORO-2-OXO-1-BENZIMIDAZOLINYL)PIPERIDINO)ETHYL)-P-FLUOROBENZAMIDE
C1997166|T121||RXNORM|BENZAMIDE DERIVATIVE ANTIPSYCHOTIC AGENT 
C1997166|T121||RXNORM|BENZAMIDE DERIVATIVE ANTIPSYCHOTIC AGENT 
C1997166|T121||RXNORM|BENZAMIDE DERIVATIVE ANTIPSYCHOTIC AGENT
C1997166|T121||RXNORM|BENZAMIDE ANTIPSYCHOTIC
C0080138|T121||RXNORM|SCH 23390
C0080138|T121||RXNORM|SCH-23390
C0080138|T121||RXNORM|SCH23390
C2348790|T121||RXNORM|TILOZEPINE
C2348297|T121||RXNORM|DIMEPROZAN
C2348661|T121||RXNORM|TERBEQUINIL
C0075494|T121||RXNORM|2-((3-(2-CHLOROETHYL)TETRAHYDRO-2H-1,3,2-OXAZAPHOSPHORIN-2-YL)AMINO)ETHANOL, METHANESULFONATE (ESTER), P-OXIDE
C0075494|T121||RXNORM|3-(2-CHLOROETHYL)-2-(2-MESYLOXYETHYLAMINO)TETRAHYDRO-2H-1,3,2-OXAZAPHOSPHORINE 2-OXIDE
C0075494|T121||RXNORM|CYTIMUN
C0075494|T121||RXNORM|SUFOSFAMIDE
C2347049|T121||RXNORM|BRAZERGOLINE
C2346736|T121||RXNORM|AMICARBALIDE
C2347353|T121||RXNORM|NIFURSEMIZONE
C0762225|T121||RXNORM|ABAPERIDONE
C0762225|T121||RXNORM|7-(3-(4-(6-FLUORO-1,2-BENZISOXAZOL-3-YL)PIPERIDIN-1-YL)PROPOXY)-3-(HYDROXYMETHYL)CHROMEN-4-ONE
C2346888|T121||RXNORM|AXAMOZIDE
C0052743|T121||RXNORM|AZABUPERONE
C0052743|T121||RXNORM|AZABUTYRONE
C2346967|T121||RXNORM|BATOPRAZINE
C0771221|T121||RXNORM|CARPHENAZINE
C0039936|T121|10498|RXNORM|THIOPROPERAZINE|THIOPROPERAZINE
C0039936|T121|10498|RXNORM|10H-PHENOTHIAZINE-2-SULFONAMIDE, N,N-DIMETHYL-10-(3-(4-METHYL-1-PIPERAZINYL)PROPYL)-|THIOPROPERAZINE
C1451709|T121||RXNORM|SONEPIPRAZOLE
C1451709|T121||RXNORM|ISOCHR-ETPIP-PHSO2NH2
C1451709|T121||RXNORM|4-(4-(2-(ISOCHROMAN-1-YL)ETHYL)PIPERAZIN-1-YL)BENZENESULFONAMIDE
C1451709|T121||RXNORM|4-(4-(2-(3,4-DIHYDRO-1H-2-BENZOPYRAN-1-YL)ETHYL)-1-PIPERAZINYL)BENZENESULFONAMIDE MONOMETHANESULFONATE
C2348431|T121||RXNORM|ALPERTINE
C0256089|T121|76887|RXNORM|QUINAGOLIDE|QUINAGOLIDE
C0256089|T121|76887|RXNORM|DOPAMINE AGONISTS CV 205-502|QUINAGOLIDE
C0256089|T121|76887|RXNORM|QUINAGOLIDE |QUINAGOLIDE
C0256089|T121|76887|RXNORM|N,N-DIETHYL-N'-(1,2,3,4,4A,5,10,10A-OCTAHYDRO-6-HYDROXY-1-PROPYL-3-BENZO(G)QUINOLINYL)SULFAMIDE, (3ALPHA,4AALPHA,10ABETA)-(+-)-ISOMER|QUINAGOLIDE
C0256089|T121|76887|RXNORM|QUINAGOLIDE, (3ALPHA,4AALPHA,10ABETA)-(+-)-ISOMER|QUINAGOLIDE
C0256089|T121|76887|RXNORM|QUINAGOLIDE |QUINAGOLIDE
C0256089|T121|76887|RXNORM|QUINAGOLIDE |QUINAGOLIDE
C2348812|T121||RXNORM|TRABOXOPINE
C0071968|T121|34479|RXNORM|3-PIPERIDINO-1,1-DIPHENYLPROPANOL|PRIDINOL
C0071968|T121|34479|RXNORM|3-PIPERIDINYL-1,1-DIPHENYLPROPAN-1-OL|PRIDINOL
C0071968|T121|34479|RXNORM|ALPHA,ALPHA-DIPHENYL-1-PIPERIDINEPROPANOL|PRIDINOL
C0071968|T121|34479|RXNORM|PRIDINOL|PRIDINOL
C0071968|T121|34479|RXNORM|RIDINOL|PRIDINOL
C2347680|T121||RXNORM|PRINOMIDE TROMETHAMINE
C2346887|T121||RXNORM|AVITRIPTAN FUMARATE
C2346887|T121||RXNORM|1H-INDOLE-5-METHANESULFONAMIDE, 3-(3-(4-(5-METHOXY-4-PYRIMIDINYL)-1-PIPERAZINYL)PROPYL)-N-METHYL-, (E)-2-BUTENEDIOATE (1:1)
C2348400|T121||RXNORM|ELOPIPRAZOLE
C2346998|T121||RXNORM|BENZINDOPYRINE HYDROCHLORIDE
C2348601|T121||RXNORM|SULMEPRIDE
C2347211|T121||RXNORM|BROCLEPRIDE
C2346718|T121||RXNORM|ACAPRAZINE
C0115127|T121||RXNORM|DUOPERONE FUMARATE
C2347032|T121||RXNORM|BISORCIC
C2346745|T121||RXNORM|AMIPERONE
C2346894|T121||RXNORM|AZAQUINZOLE
C2346785|T121||RXNORM|ANISOPIROL
C0002333|T121|596|RXNORM|ALPRAZOLAM|ALPRAZOLAM
C0002333|T121|596|RXNORM|4H-(1,2,4)TRIAZOLO(4,3-A)(1,4)BENZODIAZEPINE, 8-CHLORO-1-METHYL-6-PHENYL-|ALPRAZOLAM
C0002333|T121|596|RXNORM|ALPRAZOLAM |ALPRAZOLAM
C0002333|T121|596|RXNORM|ALPRAZOLAN|ALPRAZOLAM
C0002333|T121|596|RXNORM|ALPRAZOLAM [CHEMICAL/INGREDIENT]|ALPRAZOLAM
C0002333|T121|596|RXNORM|ALPRAZOLAM - CHEMICAL|ALPRAZOLAM
C0002333|T121|596|RXNORM|ALPRAZOLAM - CHEMICAL |ALPRAZOLAM
C0002333|T121|596|RXNORM|ALPRAZOLAM |ALPRAZOLAM
C0002333|T121|596|RXNORM|ALPRAZOLAM |ALPRAZOLAM
C0008188|T121|2356|RXNORM|CHLORDIAZEPOXIDE|CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|7 CHLORO N METHYL 5 PHENYL 3H 1,4 BENZODIAZEPIN 2 AMINE 4 OXIDE|CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|3H-1,4-BENZODIAZEPIN-2-AMINE, 7-CHLORO-N-METHYL-5-PHENYL-, 4-OXIDE|CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|3H-1,4-BENZODIAZEPIN-2-AMINE, 7-CHLORO-N-METHYL-5-PHENYL, 4-OXIDE|CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|CHLORDIAZEPOXIDE (DISCONTINUED)|CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|CHLORDIAZEPOXIDE (DISCONTINUED) |CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|7-CHLORO-N-METHYL-5-PHENYL-3H-1,4-BENZODIAZEPIN-2-AMINE 4-OXIDE|CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|CHLORDIAZEPOXIDE [CHEMICAL/INGREDIENT]|CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|METHAMINODIAZEPOXIDE|CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|CHLORDIAZEPOXIDE |CHLORDIAZEPOXIDE
C0008188|T121|2356|RXNORM|CHLORDIAZEPOXIDE |CHLORDIAZEPOXIDE
C0009011|T121|2598|RXNORM|CLONAZEPAM|CLONAZEPAM
C0009011|T121|2598|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 5-(2-CHLOROPHENYL)-1,3-DIHYDRO-7-NITRO-|CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM |CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM [CHEMICAL/INGREDIENT]|CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM [STATUS EPILEPSY]|CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM [STATUS EPILEPSY] |CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM [EPILEPSY CONTROL]|CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM [EPILEPSY CONTROL] |CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM |CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM |CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM [EPILEPSY CONTROL] |CLONAZEPAM
C0009011|T121|2598|RXNORM|CLONAZEPAM [STATUS EPILEPSY] |CLONAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM|DIAZEPAM
C0012010|T121|3322|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-1,3-DIHYDRO-1-METHYL-5-PHENYL-|DIAZEPAM
C0012010|T121|3322|RXNORM|7-CHLORO-1,3-DIHYDRO-1-METHYL-5-PHENYL-2H-1,4-BENZODIAZEPIN-2-ONE|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM AS ANXIOLYTIC |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM AS ANXIOLYTIC|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [CHEMICAL/INGREDIENT]|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [ANXIOLYTIC]|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [ANESTHESIA]|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [SKELETAL MUSCLE RELAXANT] |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [ANXIOLYTIC] |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [EPILEPSY USE] |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [EPILEPSY USE]|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [SKELETAL MUSCLE RELAXANT]|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [ANAESTHESIA]|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [ANESTHESIA] |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM PRODUCT|DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [ANESTHESIA] |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [ANXIOLYTIC] |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [EPILEPSY USE] |DIAZEPAM
C0012010|T121|3322|RXNORM|DIAZEPAM [SKELETAL MUSCLE RELAXANT] |DIAZEPAM
C0016375|T121|4501|RXNORM|FLURAZEPAM|FLURAZEPAM
C0016375|T121|4501|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-1-(2-(DIETHYLAMINO)ETHYL)-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-|FLURAZEPAM
C0016375|T121|4501|RXNORM|FLURAZEPAM [CHEMICAL/INGREDIENT]|FLURAZEPAM
C0016375|T121|4501|RXNORM|7-CHLORO-1-(2-(DIETHYLAMINO)ETHYL)-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-2H-1,4-BENZODIAZEPIN-2-ONE|FLURAZEPAM
C0016375|T121|4501|RXNORM|FLURAZEPAM |FLURAZEPAM
C0016375|T121|4501|RXNORM|FLURAZEPAM |FLURAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM|LORAZEPAM
C0024002|T121|6470|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-5-(2-CHLOROPHENYL)-1,3-DIHYDRO-3-HYDROXY-|LORAZEPAM
C0024002|T121|6470|RXNORM|7-CHLORO-5-(2-CHLOROPHENYL)-1, 3-DIHYDRO-3-HYDROXY-1,4- BENZODIAZEPIN-2-ONE|LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM |LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [CHEMICAL/INGREDIENT]|LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [EPILEPSY] |LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [ANESTHESIA]|LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [ANESTHESIA] |LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [ANXIOLYTIC] |LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [ANAESTHESIA]|LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [EPILEPSY]|LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [ANXIOLYTIC]|LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM |LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM |LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [ANESTHESIA] |LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [ANXIOLYTIC] |LORAZEPAM
C0024002|T121|6470|RXNORM|LORAZEPAM [EPILEPSY] |LORAZEPAM
C0026056|T121|6960|RXNORM|MIDAZOLAM|MIDAZOLAM
C0026056|T121|6960|RXNORM|4H-IMIDAZO(1,5-A)(1,4)BENZODIAZEPINE, 8-CHLORO-6-(2-FLUOROPHENYL)-1-METHYL-|MIDAZOLAM
C0026056|T121|6960|RXNORM|8-CHLORO-6-(2-FLUOROPHENYL)-1-METHYL- 4H- IMIDAZO(1,5A)(1,4)BENZODIAZEPINE|MIDAZOLAM
C0026056|T121|6960|RXNORM|MIDAZOLAM |MIDAZOLAM
C0026056|T121|6960|RXNORM|SEDATIVES MIDAZOLAM|MIDAZOLAM
C0026056|T121|6960|RXNORM|MIDAZOLAM [CHEMICAL/INGREDIENT]|MIDAZOLAM
C0026056|T121|6960|RXNORM|MIDAZOLAM |MIDAZOLAM
C0026056|T121|6960|RXNORM|MIDAZOLAM |MIDAZOLAM
C0029997|T121|7781|RXNORM|OXAZEPAM|OXAZEPAM
C0029997|T121|7781|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-1,3-DIHYDRO-3-HYDROXY-5-PHENYL-|OXAZEPAM
C0029997|T121|7781|RXNORM|RO 5-6789|OXAZEPAM
C0029997|T121|7781|RXNORM|SERESTA|OXAZEPAM
C0029997|T121|7781|RXNORM|OXAZEPAM |OXAZEPAM
C0029997|T121|7781|RXNORM|OXAZEPAM [CHEMICAL/INGREDIENT]|OXAZEPAM
C0029997|T121|7781|RXNORM|WY-3498|OXAZEPAM
C0029997|T121|7781|RXNORM|OXAZEPAM |OXAZEPAM
C0029997|T121|7781|RXNORM|OXAZEPAM |OXAZEPAM
C0040879|T121|10767|RXNORM|TRIAZOLAM|TRIAZOLAM
C0040879|T121|10767|RXNORM|4H-(1,2,4)TRIAZOLO(4,3-A)(1,4)BENZODIAZEPINE, 8-CHLORO-6-(2-CHLOROPHENYL)-1-METHYL-|TRIAZOLAM
C0040879|T121|10767|RXNORM|CLORAZOLAM|TRIAZOLAM
C0040879|T121|10767|RXNORM|TRIAZOLAM |TRIAZOLAM
C0040879|T121|10767|RXNORM|SEDATIVES TRIAZOLAM|TRIAZOLAM
C0040879|T121|10767|RXNORM|TRIAZOLAM [CHEMICAL/INGREDIENT]|TRIAZOLAM
C0040879|T121|10767|RXNORM|8-CHLORO-6-(2-CHLOROPHENYL)-1-METHYL-4H-(1,2,4)TRIAZOLO(4,3-A)(1,4)BENZODIAZEPINE|TRIAZOLAM
C0040879|T121|10767|RXNORM|TRIAZOLAM |TRIAZOLAM
C0040879|T121|10767|RXNORM|TRIAZOLAM |TRIAZOLAM
C0055891|T121|21241|RXNORM|1-PHENYL-5-METHYL-8-CHLORO-1,2,4,5- TETRAHYDRO-2,4-DIKETO-3H-1,5-BENZODIAZEPINE|CLOBAZAM
C0055891|T121|21241|RXNORM|CLOBAZAM|CLOBAZAM
C0055891|T121|21241|RXNORM|CLOBAZAM |CLOBAZAM
C0055891|T121|21241|RXNORM|CLOBAZAM [CHEMICAL/INGREDIENT]|CLOBAZAM
C0055891|T121|21241|RXNORM|CLOBAZAM [EPILEPSY ONLY]|CLOBAZAM
C0055891|T121|21241|RXNORM|CLOBAZAM [EPILEPSY ONLY] |CLOBAZAM
C0055891|T121|21241|RXNORM|CLOBAZAM |CLOBAZAM
C0055891|T121|21241|RXNORM|CLOBAZAM |CLOBAZAM
C0055891|T121|21241|RXNORM|CLOBAZAM [EPILEPSY ONLY] |CLOBAZAM
C0682884|T121||RXNORM|SHORT-ACTING BENZODIAZEPINES
C0682884|T121||RXNORM|SHORT-ACTING BENZODIAZEPINES 
C0008174|T121|2353|RXNORM|CLORAZEPATE|CLORAZEPATE
C0008174|T121|2353|RXNORM|ANXIOLYTICS CLORAZEPATE|CLORAZEPATE
C0008174|T121|2353|RXNORM|CLORAZEPATE |CLORAZEPATE
C0008174|T121|2353|RXNORM|CLORAZEPATE |CLORAZEPATE
C0008174|T121|2353|RXNORM|CLORAZEPATE PRODUCT |CLORAZEPATE
C0008174|T121|2353|RXNORM|CLORAZEPATE PRODUCT|CLORAZEPATE
C0008174|T121|2353|RXNORM|CHLORAZEPATE|CLORAZEPATE
C0917859|T121|1999183|RXNORM|HYDROCHLORIDE, ZOLAZEPAM|ZOLAZEPAM HYDROCHLORIDE
C0917859|T121|1999183|RXNORM|ZOLAZEPAM HYDROCHLORIDE|ZOLAZEPAM HYDROCHLORIDE
C0917859|T121|1999183|RXNORM|ZOLAZEPAM HYDROCHLORIDE |ZOLAZEPAM HYDROCHLORIDE
C0552500|T121||RXNORM|HYDROXYALPRAZOLAM
C0552500|T121||RXNORM|HYDROXYALPRAZOLAM 
C0552500|T121||RXNORM|HYDROXYALPRAZOLAM 
C0064304|T121|28181|RXNORM|11-CHLORO-8,12B-DIHYDRO-2,8-DIMETHYL-12B-PHENYL-4H-(1,3)OXAZINO(3,2-D)(1,4)BENZODIAZEPINE-4,7(6H)-DIONE|KETAZOLAM
C0064304|T121|28181|RXNORM|KETAZOLAM|KETAZOLAM
C0064304|T121|28181|RXNORM|KETAZOLAM |KETAZOLAM
C0064304|T121|28181|RXNORM|KETAZOLAM |KETAZOLAM
C0064304|T121|28181|RXNORM|KETAZOLAM |KETAZOLAM
C0006213|T121|1749|RXNORM|BROMAZEPAM|BROMAZEPAM
C0006213|T121|1749|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-BROMO-1,3-DIHYDRO-5-(2-PYRIDINYL)-|BROMAZEPAM
C0006213|T121|1749|RXNORM|BROMAZEPAM |BROMAZEPAM
C0006213|T121|1749|RXNORM|BROMAZEPAM [CHEMICAL/INGREDIENT]|BROMAZEPAM
C0006213|T121|1749|RXNORM|7-BROMO-1,3-DIHYDRO-5-(2-PYRIDYL)-2H-1,4-BENZODIAZEPIN-2-ONE|BROMAZEPAM
C0006213|T121|1749|RXNORM|BROMAZEPAM - CHEMICAL|BROMAZEPAM
C0006213|T121|1749|RXNORM|BROMAZEPAM - CHEMICAL |BROMAZEPAM
C0006213|T121|1749|RXNORM|BROMAZEPAM |BROMAZEPAM
C0006213|T121|1749|RXNORM|BROMAZEPAM |BROMAZEPAM
C0065185|T121|28894|RXNORM|7-CHLORO-5-(2-CHLOROPHENYL)-1,3-DIHYDRO-3-HYDROXY-1-METHYL-2H-1,4-BENZODIAZEPIN-2-ONE|LORMETAZEPAM
C0065185|T121|28894|RXNORM|LORMETAZEPAM|LORMETAZEPAM
C0065185|T121|28894|RXNORM|SEDATIVES LORMETAZEPAM|LORMETAZEPAM
C0065185|T121|28894|RXNORM|LORMETAZEPAM |LORMETAZEPAM
C0065185|T121|28894|RXNORM|7-CHLORO-5-(O-CHLOROPHENYL)-1,3-DIHYDRO-3-HYDROXY-1-METHYL-2H-1,4-BENZODIAZEPIN-2-ONE|LORMETAZEPAM
C0065185|T121|28894|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-5-(2-CHLOROPHENYL)-1,3-DIHYDRO-3-HYDROXY-1-METHYL-|LORMETAZEPAM
C0065185|T121|28894|RXNORM|LORMETAZEPAM |LORMETAZEPAM
C0065185|T121|28894|RXNORM|LORMETAZEPAM |LORMETAZEPAM
C0072828|T121|35185|RXNORM|7-CHLORO-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-1-(2,2,2-TRIFLUOROETHYL)-2H-1,4-BENZODIAZEPINE-2-THIONE|QUAZEPAM
C0072828|T121|35185|RXNORM|QUAZEPAM|QUAZEPAM
C0072828|T121|35185|RXNORM|2H-1,4-BENZODIAZEPINE-2-THIONE, 7-CHLORO-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-1-(2,2,2-TRIFLUOROETHYL)-|QUAZEPAM
C0072828|T121|35185|RXNORM|QUAZEPAM |QUAZEPAM
C0072828|T121|35185|RXNORM|QUAZEPAM [CHEMICAL/INGREDIENT]|QUAZEPAM
C0072828|T121|35185|RXNORM|QUAZEPAM |QUAZEPAM
C0072828|T121|35185|RXNORM|QUAZEPAM PRODUCT |QUAZEPAM
C0072828|T121|35185|RXNORM|QUAZEPAM PRODUCT|QUAZEPAM
C0014892|T121|4077|RXNORM|ESTAZOLAM|ESTAZOLAM
C0014892|T121|4077|RXNORM|4H-(1,2,4)TRIAZOLO(4,3-A)(1,4)BENZODIAZEPINE, 8-CHLORO-6-PHENYL-|ESTAZOLAM
C0014892|T121|4077|RXNORM|8-CHLORO-6-PHENYL-4H-(1,2,4)TRIAZOLO-(4,3-A)(1,4)BENZODIAZEPINE|ESTAZOLAM
C0014892|T121|4077|RXNORM|SEDATIVES ESTAZOLAM|ESTAZOLAM
C0014892|T121|4077|RXNORM|ESTAZOLAM |ESTAZOLAM
C0014892|T121|4077|RXNORM|ESTAZOLAM [CHEMICAL/INGREDIENT]|ESTAZOLAM
C0014892|T121|4077|RXNORM|ESTAZOLAM |ESTAZOLAM
C0014892|T121|4077|RXNORM|ESTAZOLAM PRODUCT |ESTAZOLAM
C0014892|T121|4077|RXNORM|ESTAZOLAM PRODUCT|ESTAZOLAM
C0011279|T121|3155|RXNORM|N DESCYCLOPROPYLMETHYL PRAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|N DESCYCLOPROPYLMETHYLPRAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|N DESTRIFLUOROETHYLHALAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|NORDAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-1,3-DIHYDRO-5-PHENYL-|NORDAZEPAM
C0011279|T121|3155|RXNORM|DESMETHYLDIAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|DEMETHYLDIAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|N-DESCYCLOPROPYLMETHYL-PRAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|N-DESCYCLOPROPYLMETHYLPRAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|N-DESTRIFLUOROETHYLHALAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|NORDAZEPAM [CHEMICAL/INGREDIENT]|NORDAZEPAM
C0011279|T121|3155|RXNORM|DEOXYDEMOXEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|NORDIAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|NORPRAZEPAM|NORDAZEPAM
C0011279|T121|3155|RXNORM|7-CHLORO-1,3-DIHYDRO-5-PHENYL-2H-1,4-BENZODIAZEPIN-2-ONE|NORDAZEPAM
C0011279|T121|3155|RXNORM|NORDAZEPAM |NORDAZEPAM
C0304401|T121||RXNORM|BENZODIAZEPINE NUCLEUS
C0304401|T121||RXNORM|BENZODIAZEPINE NUCLEUS 
C0028126|T121|7440|RXNORM|NITRAZEPAM|NITRAZEPAM
C0028126|T121|7440|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 1,3-DIHYDRO-7-NITRO-5-PHENYL-|NITRAZEPAM
C0028126|T121|7440|RXNORM|NITRAZEPAM |NITRAZEPAM
C0028126|T121|7440|RXNORM|SEDATIVES NITRAZEPAM|NITRAZEPAM
C0028126|T121|7440|RXNORM|NITRAZEPAM [CHEMICAL/INGREDIENT]|NITRAZEPAM
C0028126|T121|7440|RXNORM|NITRODIAZEPAM|NITRAZEPAM
C0028126|T121|7440|RXNORM|1,3-DIHYDRO-7-NITRO-5-PHENYL-2H-1,4-BENZODIAZEPIN-2-ONE|NITRAZEPAM
C0028126|T121|7440|RXNORM|NITRAZEPAM |NITRAZEPAM
C0028126|T121|7440|RXNORM|NITRAZEPAM |NITRAZEPAM
C0525768|T121||RXNORM|7-AMINO-FLUNITRAZEPAM
C0525768|T121||RXNORM|7-AMINOFLUNITRAZEPAM
C0525768|T121||RXNORM|7-AMINOFLUNITRAZEPAM 
C0039468|T121|10355|RXNORM|TEMAZEPAM|TEMAZEPAM
C0039468|T121|10355|RXNORM|3 HYDROXYDIAZEPAM|TEMAZEPAM
C0039468|T121|10355|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-1,3-DIHYDRO-3-HYDROXY-1-METHYL-5-PHENYL-|TEMAZEPAM
C0039468|T121|10355|RXNORM|OXYDIAZEPAM|TEMAZEPAM
C0039468|T121|10355|RXNORM|10-CHLORO-4-HYDROXY-6-METHYL-2-PHENYL-3,6-DIAZABICYCLO[5.4.0]UNDECA-2,8,10,12-TETRAEN-5-ONE|TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM |TEMAZEPAM
C0039468|T121|10355|RXNORM|HYDROXYDIAZEPAM|TEMAZEPAM
C0039468|T121|10355|RXNORM|3-HYDROXYDIAZEPAM|TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM [CHEMICAL/INGREDIENT]|TEMAZEPAM
C0039468|T121|10355|RXNORM|METHYLOXAZEPAM|TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM [ANAESTHESIA]|TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM [ANESTHESIA] |TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM [ANESTHESIA]|TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM [HYPNOTIC]|TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM [HYPNOTIC] |TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM |TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM |TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM [ANESTHESIA] |TEMAZEPAM
C0039468|T121|10355|RXNORM|TEMAZEPAM [HYPNOTIC] |TEMAZEPAM
C0016296|T121|4460|RXNORM|FLUNITRAZEPAM|FLUNITRAZEPAM
C0016296|T121|4460|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 5-(2-FLUOROPHENYL)-1,3-DIHYDRO-1-METHYL-7-NITRO-|FLUNITRAZEPAM
C0016296|T121|4460|RXNORM|FLUNITRAZEPAM |FLUNITRAZEPAM
C0016296|T121|4460|RXNORM|FLURIDRAZEPAM|FLUNITRAZEPAM
C0016296|T121|4460|RXNORM|FLUNITRAZEPAM [CHEMICAL/INGREDIENT]|FLUNITRAZEPAM
C0016296|T121|4460|RXNORM|5-(O-FLUOROPHENYL)-1,3-DIHYDRO-1-METHYL-7-NITRO-2H-1,4-BENZODIAZEPIN-2-ONE|FLUNITRAZEPAM
C0016296|T121|4460|RXNORM|FLUNITRAZEPAM |FLUNITRAZEPAM
C0016296|T121|4460|RXNORM|FLUNITRAZEPAM |FLUNITRAZEPAM
C1289963|T121||RXNORM|DESMETHYLCLOBAZAM 
C1289963|T121||RXNORM|DESMETHYLCLOBAZAM
C0063132|T121||RXNORM|HYDROXYETHYLFLURAZEPAM
C0063132|T121||RXNORM|HYDROXYETHYLFLURAZEPAM 
C0077013|T121|38555|RXNORM|6-(2-CHLOROPHENYL)-2,4-DIHYDRO-2-((4-METHYL-1-PIPERAZINYL)METHYLENE)-8-NITRO-1H-IMIDAZO(1,2-A) (1,4)BENZODIAZEPIN-1-ONE|LOPRAZOLAM
C0077013|T121|38555|RXNORM|LOPRAZOLAM|LOPRAZOLAM
C0077013|T121|38555|RXNORM|TRIAZULENONE|LOPRAZOLAM
C0077013|T121|38555|RXNORM|LOPRAZOLAM |LOPRAZOLAM
C0077013|T121|38555|RXNORM|LOPRAZOLAM |LOPRAZOLAM
C0032910|T121|8627|RXNORM|PRAZEPAM|PRAZEPAM
C0032910|T121|8627|RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-1-(CYCLOPROPYLMETHYL)-1,3-DIHYDRO-5-PHENYL-|PRAZEPAM
C0032910|T121|8627|RXNORM|PRAZEPAM (DISCONTINUED) |PRAZEPAM
C0032910|T121|8627|RXNORM|PRAZEPAM (DISCONTINUED)|PRAZEPAM
C0032910|T121|8627|RXNORM|PRAZEPAM [CHEMICAL/INGREDIENT]|PRAZEPAM
C0032910|T121|8627|RXNORM|PRAZEPAM |PRAZEPAM
C0032910|T121|8627|RXNORM|PRAZEPAM |PRAZEPAM
C0025051|T121|6680|RXNORM|MEDAZEPAM|MEDAZEPAM
C0025051|T121|6680|RXNORM|1H-1,4-BENZODIAZEPINE, 7-CHLORO-2,3-DIHYDRO-1-METHYL-5-PHENYL-|MEDAZEPAM
C0025051|T121|6680|RXNORM|MEDAZAPAM|MEDAZEPAM
C0025051|T121|6680|RXNORM|MEDAZEPAM [CHEMICAL/INGREDIENT]|MEDAZEPAM
C0025051|T121|6680|RXNORM|MEDAZAPAM |MEDAZEPAM
C0025051|T121|6680|RXNORM|MEDAZEPAM |MEDAZEPAM
C0025051|T121|6680|RXNORM|MEDAZEPAM |MEDAZEPAM
C0062092|T121|26412|RXNORM|7-CHLORO-1,3-DIHYDRO-5-PHENYL-1- (2,2,2-TRIFLUOROETHYL)-2H-1,4-BENZODIAZEPIN-2-ONE|HALAZEPAM
C0062092|T121|26412|RXNORM|HALAZEPAM|HALAZEPAM
C0062092|T121|26412|RXNORM|HALAZEPAM |HALAZEPAM
C0062092|T121|26412|RXNORM|HALAZEPAM [CHEMICAL/INGREDIENT]|HALAZEPAM
C0062092|T121|26412|RXNORM|HALAZEPAM |HALAZEPAM
C0062092|T121|26412|RXNORM|HALAZEPAM PRODUCT |HALAZEPAM
C0062092|T121|26412|RXNORM|HALAZEPAM PRODUCT|HALAZEPAM
C0552501|T121||RXNORM|HYDROXYTRIAZOLAM
C0552501|T121||RXNORM|HYDROXYTRIAZOLAM 
C0057377|T121||RXNORM|7-CHLORO-1,3-DIHYDRO-5-PHENYL-2H-1,4-BENZODIAZEPIN-2-ONE 4-OXIDE
C0057377|T121||RXNORM|DEMOXEPAM
C0057377|T121||RXNORM|DEMOXEPAM 
C0690642|T121|198317|RXNORM|TRIAZOLAM 0.125 MG ORAL TABLET|TRIAZOLAM 0.125 MG ORAL TABLET
C0690642|T121|198317|RXNORM|TRIAZOLAM 0.125MG ORAL TABLET|TRIAZOLAM 0.125 MG ORAL TABLET
C0690642|T121|198317|RXNORM|TRIAZOLAM, 0.125 MG ORAL TABLET|TRIAZOLAM 0.125 MG ORAL TABLET
C0690642|T121|198317|RXNORM|TRIAZOLAM 0.125MG TAB|TRIAZOLAM 0.125 MG ORAL TABLET
C0690642|T121|198317|RXNORM|TRIAZOLAM 0.125 MILLIGRAM IN 1 TABLET ORAL TABLET|TRIAZOLAM 0.125 MG ORAL TABLET
C0690642|T121|198317|RXNORM|TRIAZOLAM TAB 0.125 MG|TRIAZOLAM 0.125 MG ORAL TABLET
C0690642|T121|198317|RXNORM|TRIAZOLAM 0.125MG TAB [VA PRODUCT]|TRIAZOLAM 0.125 MG ORAL TABLET
C0690642|T121|198317|RXNORM|TRIAZOLAM 0.125 MG ORAL TABLET [TRIAZOLAM]|TRIAZOLAM 0.125 MG ORAL TABLET
C0690642|T121|198317|RXNORM|TRIAZOLAM 0.125MG TABLET |TRIAZOLAM 0.125 MG ORAL TABLET
C0690642|T121|198317|RXNORM|TRIAZOLAM 0.125MG TABLET|TRIAZOLAM 0.125 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM 0.25 MG ORAL TABLET|TRIAZOLAM 0.25 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM 0.25MG ORAL TABLET|TRIAZOLAM 0.25 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM, 0.25 MG ORAL TABLET|TRIAZOLAM 0.25 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM 0.25MG TAB|TRIAZOLAM 0.25 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM 0.25 MILLIGRAM IN 1 TABLET ORAL TABLET|TRIAZOLAM 0.25 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM TAB 0.25 MG|TRIAZOLAM 0.25 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM 0.25MG TAB [VA PRODUCT]|TRIAZOLAM 0.25 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM 0.25 MG ORAL TABLET [TRIAZOLAM]|TRIAZOLAM 0.25 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM 0.25MG TABLET |TRIAZOLAM 0.25 MG ORAL TABLET
C0690643|T121|198318|RXNORM|TRIAZOLAM 0.25MG TABLET|TRIAZOLAM 0.25 MG ORAL TABLET
C4048284|T121||RXNORM|BENZODIAZEPINE
C4048284|T121||RXNORM|BENZODIAZEPINE 
C4048284|T121||RXNORM|BENZODIAZEPINE 
C4048284|T121||RXNORM|BENZODIAZEPINE, NOS
C0071082|T121||RXNORM|7-CHLORO-5-PHENYL-1-PROPARGYL-1,4-BENZODIAZEPIN-2- ONE
C0071082|T121||RXNORM|PINAZEPAM
C0071082|T121||RXNORM|PROPAZEPAM
C0071082|T121||RXNORM|PINAZEPAM 
C0071082|T121||RXNORM|PINAZEPAM 
C0009073|T121|2622|RXNORM|CLOTIAZEPAM|CLOTIAZEPAM
C0009073|T121|2622|RXNORM|2H-THIENO(2,3-E)-1,4-DIAZEPIN-2-ONE, 5-(2-CHLOROPHENYL)-7-ETHYL-1,3-DIHYDRO-1-METHYL-|CLOTIAZEPAM
C0009073|T121|2622|RXNORM|CLOTIAZEPAM |CLOTIAZEPAM
C0053117|T121||RXNORM|1,3,6,7,8,9-HEXAHYDRO-5-PHENYL-2H-(1)BENZOTHIENO(2,3-E)-1,4-DIAZEPIN-2-ONE
C0053117|T121||RXNORM|6,7-TETRAMETHYLENE-5-PHENYL-1,2-DIHYDRO-3H-THIENO(2,3-E)(1,4)DIAZEPIN-2-ONE
C0053117|T121||RXNORM|BENTAZEPAM
C0053117|T121||RXNORM|BENTAZEPAM 
C0076341|T121|37985|RXNORM|7-CHLORO-5-(1-CYCLOHEXEN-1- YL)-1,3-DIHYDRO-1-METHYL-2H-1,4-BENZODIAZEPIN-2-ONE|TETRAZEPAM
C0076341|T121|37985|RXNORM|TETRAZEPAM|TETRAZEPAM
C0076341|T121|37985|RXNORM|TETRAZEPAM |TETRAZEPAM
C0076341|T121|37985|RXNORM|TETRAZEPAM |TETRAZEPAM
C0054151|T121|19790|RXNORM|2-BROMO-4-(2-CHLOROPHENYL)-9-METHYL-6H-THIENO(3,2-F)(1,2,4)TRIAZOLO(4,3-A)(1,4)DIAZEPINE|BROTIZOLAM
C0054151|T121|19790|RXNORM|BROTIZOLAM|BROTIZOLAM
C0054151|T121|19790|RXNORM|SEDATIVES BROTIZOLAM|BROTIZOLAM
C0054151|T121|19790|RXNORM|BROTIZOLAM |BROTIZOLAM
C0054151|T121|19790|RXNORM|6H-THIENO(3,2-F)(1,2,4)TRIAZOLO(4,3-A)(1,4)DIAZEPINE,2-BROMO-4-(2-CHLOROPHENYL)-9-METHYL-|BROTIZOLAM
C0054151|T121|19790|RXNORM|2-BROMO-4-(O-CHLOROPHENYL)-9-METHYL-6H-THIENO(3,2-F)-S-TRIAZOLO(4,3-A)(1,4)DIAZEPINE|BROTIZOLAM
C0054151|T121|19790|RXNORM|BROTIZOLAM |BROTIZOLAM
C0005064|T121||RXNORM|BENZODIAZEPINES
C0005064|T121||RXNORM|BENZODIAZEPINE CPDS
C0005064|T121||RXNORM|BENZODIAZEPINES 
C0005064|T121||RXNORM|BENZODIAZEPINES [CHEMICAL/INGREDIENT]
C0005064|T121||RXNORM|BENZODIAZEPINE COMPOUNDS
C0005064|T121||RXNORM|BENZODIAZEPINE
C0360114|T121||RXNORM|BENZODIAZEPINE SEDATIVE
C0360114|T121||RXNORM|BENZODIAZEPINE SEDATIVE 
C0360114|T121||RXNORM|BENZODIAZEPINE SEDATIVE 
C0053218|T121||RXNORM|BENZODIAZEPINE ANTIEPILEPTIC 
C0053218|T121||RXNORM|BENZODIAZEPINE ANTIEPILEPTIC
C0242293|T121|71484|RXNORM|FLURAZEPAM HYDROCHLORIDE|FLURAZEPAM HYDROCHLORIDE
C0242293|T121|71484|RXNORM|HYDROCHLORIDE, FLURAZEPAM|FLURAZEPAM HYDROCHLORIDE
C0242293|T121|71484|RXNORM|FLURAZEPAM HYDROCHLORIDE |FLURAZEPAM HYDROCHLORIDE
C0242293|T121|71484|RXNORM|FLURAZEPAM HYDROCHLORIDE [CHEMICAL/INGREDIENT]|FLURAZEPAM HYDROCHLORIDE
C0242293|T121|71484|RXNORM|FLURAZEPAM DIHYDROCHLORIDE|FLURAZEPAM HYDROCHLORIDE
C0242293|T121|71484|RXNORM|DIHYDROCHLORIDE, FLURAZEPAM|FLURAZEPAM HYDROCHLORIDE
C0242293|T121|71484|RXNORM|INSUMIN DIHYDROCHLORIDE|FLURAZEPAM HYDROCHLORIDE
C0242293|T121|71484|RXNORM|FLURAZEPAM HCL|FLURAZEPAM HYDROCHLORIDE
C0242293|T121|71484|RXNORM|FLURAZEPAM HYDROCHLORIDE |FLURAZEPAM HYDROCHLORIDE
C0057905|T121||RXNORM|DESALKYLFLURAZEPAM
C0057905|T121||RXNORM|DESDIALKYLFLURAZEPAM
C0057905|T121||RXNORM|DIDEETHYLFLURAZEPAM
C0057905|T121||RXNORM|DIDESETHYLFLURAZEPAM
C0057905|T121||RXNORM|N-DESALKYLFLURAZEPAM
C0057905|T121||RXNORM|DESALKYLFLURAZEPAM 
C0057905|T121||RXNORM|N-1-DESALKYLFLURAZEPAM
C0005065|T121||RXNORM|BENZODIAZEPINONES
C0005065|T121||RXNORM|BENZODIAZEPINONES [CHEMICAL/INGREDIENT]
C0016293|T121|4457|RXNORM|FLUMAZENIL|FLUMAZENIL
C0016293|T121|4457|RXNORM|4H-IMIDAZO(1,5-A)(1,4)BENZODIAZEPINE-3-CARBOXYLIC ACID, 8-FLUORO-5,6-DIHYDRO-5-METHYL-6-OXO-, ETHYL ESTER|FLUMAZENIL
C0016293|T121|4457|RXNORM|FLUMAZENIL |FLUMAZENIL
C0016293|T121|4457|RXNORM|FLUMAZENIL [CHEMICAL/INGREDIENT]|FLUMAZENIL
C0016293|T121|4457|RXNORM|FLUMAZEPIL|FLUMAZENIL
C0016293|T121|4457|RXNORM|FLUMAZENIL |FLUMAZENIL
C0016293|T121|4457|RXNORM|FLUMAZENIL |FLUMAZENIL
C0031978|T121|8352|RXNORM|PIRENZEPINE|PIRENZEPINE
C0031978|T121|8352|RXNORM|6H-PYRIDO(2,3-B)(1,4)BENZODIAZEPIN-6-ONE, 5,11-DIHYDRO-11-((4-METHYL-1-PIPERAZINYL)ACETYL)-|PIRENZEPINE
C0031978|T121|8352|RXNORM|PIRENZEPIN|PIRENZEPINE
C0031978|T121|8352|RXNORM|PYRENZEPINE|PIRENZEPINE
C0031978|T121|8352|RXNORM|PIRENZEPINE [CHEMICAL/INGREDIENT]|PIRENZEPINE
C0031978|T121|8352|RXNORM|PIRENZEPINE |PIRENZEPINE
C0031978|T121|8352|RXNORM|PIRENZEPINE |PIRENZEPINE
C0536095|T121||RXNORM|RO 48-6791
C0536095|T121||RXNORM|RO-48-6791
C0701356|T121||RXNORM|WY 4036
C0701356|T121||RXNORM|WY4036
C0701356|T121||RXNORM|WY-4036
C0702213|T121||RXNORM|TAZEPAM
C0702214|T121|204360|RXNORM|SERAX|SERAX
C0702215|T121||RXNORM|ADUMBRAN
C2352304|T121||RXNORM|RS 678
C2352304|T121||RXNORM|RS678 CPD
C2352304|T121||RXNORM|RS-678
C2352305|T121||RXNORM|RS 779
C2352305|T121||RXNORM|RS779 CPD
C2352305|T121||RXNORM|RS-779
C0009033|T121|2607|RXNORM|CHLORAZEPATE, DIPOTASSIUM|POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|CLORAZEPATE DIPOTASSIUM|POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|DIPOTASSIUM, CLORAZEPATE|POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|1H-1,4-BENZODIAZEPINE-3-CARBOXYLIC ACID, 7-CHLORO-2,3-DIHYDRO-2-OXO-5-PHENYL-, MONOPOTASSIUM SALT, COMPD. WITH POTASSIUM HYDROXIDE (K(OH)) (1:1)|POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|1H-1,4-BENZODIAZEPINE-3-CARBOXYLIC ACID, 7-CHLORO-2,3-DIHYDRO-2-OXO-5-PHENYL-, MONOPOTASSIUM SALT, COMPOUND WITH POTASSIUM HYDROXIDE|POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|POTASSIUM 7-CHLORO-2,3-DIHYDRO-2-OXO-5-PHENYL-1H-1,4-BENZODIAZEPINE-3-CARBOXYLATE KOH|POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|CLORAZEPATE DIPOTASSIUM |POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|CLORAZEPATE DIPOTASSIUM [CHEMICAL/INGREDIENT]|POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|DIPOTASSIUM CHLORAZEPATE|POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|POTASSIUM CLORAZEPATE|POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|CLORAZEPATE DIPOTASSIUM |POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|CLORAZEPATE DIPOTASSIUM |POTASSIUM CLORAZEPATE
C0009033|T121|2607|RXNORM|DIPOTASSIUM CLORAZEPATE|POTASSIUM CLORAZEPATE
C2604475|T121||RXNORM|GWL78 CPD
C2604475|T121||RXNORM|GWL 78
C2604475|T121||RXNORM|GWL-78
C2604604|T121||RXNORM|COCOBOO-ACETAMIDE
C2604604|T121||RXNORM|2-(5-CYCLOHEXYL-1-(2-CYCLOPENTYL-2-OXOETHYL)-2-OXO-1,2-DIHYDRO-3H-1,3,4-BENZOTRIAZEPIN-3-YL)-N-(3-(5-OXO-2,5-DIHYDRO-(1,2,4)OXADIAZOL-3-YL)PHENYL)ACETAMIDE
C2604810|T121||RXNORM|ETHYL FNIBC
C2604810|T121||RXNORM|ETHYL 8-FLUORO-6-(3-NITROPHENYL)-4H-IMIDAZO(1,5-A)(1,4)BENZODIAZEPINE-3-CARBOXYLATE
C2606964|T121||RXNORM|PWZ-029
C2606902|T121||RXNORM|QUINO(7,8-B)BENZODIAZEPINE
C0050844|T121||RXNORM|ADINAZOLAM
C0167214|T121||RXNORM|ADINAZOLAM MESYLATE
C0009034|T121||RXNORM|MONOPOTASSIUM, CLORAZEPATE
C0009034|T121||RXNORM|CLORAZEPATE MONOPOTASSIUM
C0009034|T121||RXNORM|CLORAZEPATE MONOPOTASSIUM 
C2699536|T121||RXNORM|CYPRAZEPAM
C2697918|T121||RXNORM|LEVOTOFISOPAM
C0068774|T121||RXNORM|1-METHYL-7-NITRO-5-PHENYL-1,3-DIHYDRO-2H-1,4- BENZODIAZEPIN-2-ONE
C0068774|T121||RXNORM|NIMETAZEPAM
C2698499|T121||RXNORM|NORTETRAZEPAM
C2699964|T121||RXNORM|TOLUFAZEPAM
C2699964|T121||RXNORM|1-(4'-METHYLPHENYLSULFONYL)ETHYL-5-(2-CHLOROPHENYL)-7-CHLORO-2H-1,4-BENZODIAZEPIN-2-ONE
C2698992|T121||RXNORM|CARBURAZEPAM
C0055715|T121||RXNORM|8-BROMO-6-(ORTHO-CHLOROPHENYL)-1-CYCLOHEXYL-4H-5-TRIAZOLO(3,4-C)THIENO(2,4-E)-1,4-DIAZEPINE
C0055715|T121||RXNORM|CICLOTIZOLAM
C0164835|T121||RXNORM|7-CHLORO-5-(2-FLUOROPHENYL)-2,3-DIHYDRO-3-HYDROXY-2-OXO-1H-1,4-BENZODIAZEPINE-1-PROPIONITRILE
C0164835|T121||RXNORM|CINOLAZEPAM
C0110063|T121||RXNORM|4H-IMIDAZO(1,5-A)(1,4)BENZODIAZEPINE, 8-CHLORO-6-(2-CHLOROPHENYL)-1-METHYL-
C0110063|T121||RXNORM|8-CHLORO-6-(2-CHLOROPHENYL)-1-METHYL-4H-IMIDAZO(1,5A)(1,4)BENZODIAZEPINE
C0110063|T121||RXNORM|CLIMAZOLAM
C2714934|T121||RXNORM|7-CHLORO-4-(CYCLOHEXYLMETHYL)-1-METHYL-3,4-DIHYDRO-1H-1,4-BENZODIAZEPINE-2,5-DIONE
C2714934|T121||RXNORM|BNZ-1 CPD
C2714935|T121||RXNORM|4-CYCLOHEXYLMETHYL-1-METHYL-3,4-DIHYDRO-1H-1,4-BENZODIAZEPINE-2,5-DIONE
C2714935|T121||RXNORM|BNZ-2 CPD
C2715396|T121||RXNORM|IODOPHENYL-MOPDBDU
C2715396|T121||RXNORM|1-(3-IODOPHENYL)-3-(1-METHYL-2-OXO-5-PHENYL-2,3-DIHYDRO-1H-BENZO(E)(1,4)DIAZEPIN-3-YL)UREA
C2715729|T121||RXNORM|LIMAZEPINE B1
C2715731|T121||RXNORM|LIMAZEPINE D
C2717477|T121||RXNORM|RO4938581
C2717477|T121||RXNORM|3-BROMO-10-DIFLUOROMETHYL-9H-IMIDAZO(1,5-A)(1,2,4)TRIAZOLO(1,5-D)(1,4)BENZODIAZEPINE
C2744849|T121||RXNORM|RO 4882224
C2744849|T121||RXNORM|RO4882224
C2744849|T121||RXNORM|RO-4882224
C0604102|T121||RXNORM|7-CHLORO-2,3-DIHYDRO-1-(2,2,2-TRIFLUOROETHYL)-5-(O-FLUOROPHENYL)-1H-1,4-BENZODIA ZEPINE
C0604102|T121||RXNORM|FLETAZEPAM
C0065179|T121||RXNORM|2H-PYRIDO(3,2-E)-1,4-DIAZEPIN-2-ONE, 7-CHLORO-5-(2-CHLOROPHENYL)-1,3-DIHYDRO-3-HYDROXY-
C0065179|T121||RXNORM|3-HYDROXY-5-(O-CHLOROPHENYL)-7-CHLORO-1,2-DIHYDRO-2H-PYRIDO(3,2-E)-1,4-DIAZEPIN-2-ONE
C0065179|T121||RXNORM|LOPIRAZEPAM
C0089958|T121||RXNORM|10-CHLORO-2,3,7,11B-TETRAHYDRO-3-METHYL-11B-(2-CHLOROPHENYL)OXAZOLO(3,2-D)(1,4)BENZODIAZEPIN-6(5H)-ONE
C0089958|T121||RXNORM|MEXAZOLAM
C0089958|T121||RXNORM|10-CHLORO-11B-(2-CHLOROPHENYL)-2,3,7,11B-TETRAHYDRO-3-METHYLOXAZOLO(3,2-D)(1,4)BENZODIAZEPIN-6(5H)-ONE
C0120735|T121||RXNORM|10-BROMO-11B-(2-FLUOROPHENYL)-2,3,7,11B-TETRAHYDROOXAZOLO(3,2-D)(1,4)BENZODIAZEPIN-6(5H)-ONE
C0120735|T121||RXNORM|HALOXAZOLAM
C0065842|T121||RXNORM|3-METHYLCLONAZEPAM
C0065842|T121||RXNORM|5-(2-CHLOROPHENYL)-1,3-DIHYDRO-3-METHYL-7-NITRO- 2H-1,4-BENZODIAZEPIN-2-ONE
C0065842|T121||RXNORM|MECLONAZEPAM
C1619621|T121|614654|RXNORM|1H-1,4-BENZODIAZEPINE, 7-BROMO-5-(2-CHLOROPHENYL)-2,3-DIHYDRO-2-(METHOXYMETHYL)-1-METHYL-|METACLAZEPAM
C1619621|T121|614654|RXNORM|1H-1,4-BENZODIAZEPINE, 7-BROMO-5-(2-CHLOROPHENYL)-2,3-DIHYDRO-2-METHOXY-1-METHYL-|METACLAZEPAM
C1619621|T121|614654|RXNORM|METACLAZEPAM|METACLAZEPAM
C0066040|T121|29590|RXNORM|METACLAZEPAM HYDROCHLORIDE|METACLAZEPAM HYDROCHLORIDE
C0066040|T121|29590|RXNORM|7-BROMO-5-(O-CHLOROPHENYL)-2,3-DIHYDRO-2-(METHOXYMETHYL)-1-METHYL-1H-1,4-BENZODIAZEPINE HYDROCHLORIDE|METACLAZEPAM HYDROCHLORIDE
C0066040|T121|29590|RXNORM|7-BROMO-5-(2-CHLOROPHENYL)-2,3-DIHYDRO-2-(METHOXYMETHYL)-1-METHYL-1H-1,4-BENZODIAZEPINE HYDROCHLORIDE|METACLAZEPAM HYDROCHLORIDE
C0066040|T121|29590|RXNORM|BROMETAZEPAM HYDROCHLORIDE|METACLAZEPAM HYDROCHLORIDE
C0066040|T121|29590|RXNORM|METUCLAZEPAM HYDROCHLORIDE|METACLAZEPAM HYDROCHLORIDE
C0066040|T121|29590|RXNORM|7-BROMO-5-(2'-CHLOROPHENYL)-2,3-DIHYDRO-2-(METHOXYL)-1-METHYL-1H-1,4-BENZODIAZEPINE.HCL|METACLAZEPAM HYDROCHLORIDE
C0027556|T121|7285|RXNORM|NEFOPAM|NEFOPAM
C0027556|T121|7285|RXNORM|1H-2,5-BENZOXAZOCINE, 3,4,5,6-TETRAHYDRO-5-METHYL-1-PHENYL-|NEFOPAM
C0027556|T121|7285|RXNORM|NEFOPAM [CHEMICAL/INGREDIENT]|NEFOPAM
C0027556|T121|7285|RXNORM|BENZOXAZOCINE|NEFOPAM
C0027556|T121|7285|RXNORM|NEFOPAM |NEFOPAM
C0027556|T121|7285|RXNORM|NEFOPAM |NEFOPAM
C0015820|T121|4324|RXNORM|HYDROCHLORIDE, NEFOPAM|NEFOPAM HYDROCHLORIDE
C0015820|T121|4324|RXNORM|NEFOPAM HYDROCHLORIDE|NEFOPAM HYDROCHLORIDE
C0015820|T121|4324|RXNORM|NEFOPAM HYDROCHLORIDE |NEFOPAM HYDROCHLORIDE
C0015820|T121|4324|RXNORM|3,4,5,6-TETRAHYDRO-5-METHYL-1-PHENYL-1H-2,5-BENZOXAZOCINE HYDROCHLORIDE|NEFOPAM HYDROCHLORIDE
C0015820|T121|4324|RXNORM|NEFOPAM HYDROCHLORIDE PRODUCT |NEFOPAM HYDROCHLORIDE
C0015820|T121|4324|RXNORM|NEFOPAM HYDROCHLORIDE PRODUCT|NEFOPAM HYDROCHLORIDE
C0015820|T121|4324|RXNORM|FENAZOXINE|NEFOPAM HYDROCHLORIDE
C0015820|T121|4324|RXNORM|NEFOPAM HYDROCHLORIDE |NEFOPAM HYDROCHLORIDE
C0055964|T121|21311|RXNORM|10-CHLORO-2,3,5,6,7,11B-HEXAHYDRO-11B-(O- CHLOROPHENYL)BENZO(6,7)-1,4-DIAZEPINO-(5,4-B)-OXAZOL-6-ONE|CLOXAZOLAM
C0055964|T121|21311|RXNORM|CLOXAZOLAM|CLOXAZOLAM
C0055964|T121|21311|RXNORM|CLOXAZOLAM |CLOXAZOLAM
C0055964|T121|21311|RXNORM|BETAVEL|CLOXAZOLAM
C0055964|T121|21311|RXNORM|10-CHLORO-11B-(O-CHLOROPHENYL)-2,3,7,11B-TETRAHYDRO-OXAZOLO(3,2-D) (1,4)BENZODIAZEPIN-6(5H)-ONE|CLOXAZOLAM
C0055964|T121|21311|RXNORM|ENADEL|CLOXAZOLAM
C0055964|T121|21311|RXNORM|TOLESTAN|CLOXAZOLAM
C0059772|T121|24524|RXNORM|1H-1,4-BENZODIAZEPINE-3-CARBOXYLIC ACID, 7-CHLORO-5-(2-FLUOROPHENYL)-2,3-DIHYDRO-2-OXO-, ETHYL ESTER|ETHYL LOFLAZEPATE
C0059772|T121|24524|RXNORM|ETHYL FLUCOZEPATE|ETHYL LOFLAZEPATE
C0059772|T121|24524|RXNORM|ETHYL LOFLAZEPATE|ETHYL LOFLAZEPATE
C0059772|T121|24524|RXNORM|ETHYL LOFLAZEPATE |ETHYL LOFLAZEPATE
C0059862|T121||RXNORM|ETIZOLAM
C0059862|T121||RXNORM|ETIZOLAM 
C2932012|T121||RXNORM|4-(3,5-DIHYDROXYBENZYL)-N-(2-METHYL-4-((1-METHYL-4,10-DIHYDROPYRAZOLO(3,4-B)(1,5)BENZODIAZEPIN-5(1H)-YL)CARBONYL)BENZYL)PIPERAZINE-1-CARBOXAMIDE
C2933864|T121||RXNORM|EVT 201
C2933864|T121||RXNORM|EVT201
C2933864|T121||RXNORM|EVT-201
C2934398|T121||RXNORM|2-AMINO-PPBI
C2934398|T121||RXNORM|2-AMINO-4-(PIPERIDIN-1-YL)-11H-PYRIMIDO(4,5-B)(1,5)BENZODIAZEPIN-6-IUM
C2934400|T121||RXNORM|2-AMINO-4-(METHYL(2-METHYLPHENYL)AMINO)-11H-PYRIMIDO(4,5-B)(1,5)BENZODIAZEPIN-6-IUM
C2934400|T121||RXNORM|2-AMINO-MMAPBI
C2935069|T121||RXNORM|BENZOPYRANO(4,3-C)-1,5-BENZODIAZEPINE
C2935196|T121||RXNORM|TKM0150
C2976597|T121||RXNORM|5-(2-CHLOROPHENYL)-7-FLUORO-1,2-DIHYDRO-8-METHOXY-3-METHYLPYRAZOL(3,4B)(1,4)BENZODIAZEPINE
C1527794|T121||RXNORM|DIAZEPINOMICIN
C1527794|T121||RXNORM|11H-DIBENZO(B,E)(1,4)DIAZEPIN-11-ONE, 5,10-DIHYDRO-4,6,8-TRIHYDROXY-10-((2E,6E)-3,7,11-TRIMETHYL-2,6,10-DODECATRIEN-1-YL)-
C0117998|T121||RXNORM|7-CHLORO-1-CYCLOPROPYLMETHYL-1,3-DIHYDRO-5-(2-FLUOROPHENYL)-2H-1,4-BENZODIAZEPIN-2-ONE
C0117998|T121||RXNORM|FLUTOPRAZEPAM
C1881907|T121||RXNORM|MOTRAZEPAM
C1881907|T121||RXNORM|2,3-DIHYDRO-1-(METHOXYMETHYL)-7-NITRO-5-PHENYL-1H-1,4-BENZODIAZEPIN-2-ON
C0605583|T121||RXNORM|7-CHLORO-1,3-DIHYDRO-5-PHENYL-1H-2-OXO-3-PIVALYLOXY- 1,4-BENZODIAZEPINE
C0605583|T121||RXNORM|PIVOXAZEPAM
C0605583|T121||RXNORM|7-CHLORO-1,3-DIHYDRO-3-HYDROXY-5-PHENYL-2H-1,4-BENZODIAZEPIN-2-ONE PIVALATE (ESTER)
C2348591|T121||RXNORM|SULAZEPAM
C0059029|T121||RXNORM|7-CHLORO-1-(2-(ETHYLSULFONYL)ETHYL)-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-2H-1,4-BENZODIAZEP IN-2-ONE
C0059029|T121||RXNORM|ELFAZEPAM
C2347902|T121||RXNORM|RECLAZEPAM
C2347902|T121||RXNORM|2-(7-CHLORO-5-(O-CHLOROPHENYL)-2,3-DIHYDRO-1H-1,4-BENZODIAZEPIN-1-YL)-2-OXAZOLIN-4-ONE
C2347902|T121||RXNORM|4(5H)-OXAZOLONE, 2-(7-CHLORO-5-(2-CHLOROPHENYL)-2,3-DIHYDRO-1H-1,4-BENZODIAZEPIN-1-YL)-
C3272985|T121||RXNORM|3-(11-DIMETHYLHEPTYL)-7,8,9,10-TETRAHYDRO-6,6,9-TRIMETHYL-6H-DIBENZO(B,D)PYRAN-1-YL 4-(1-AZEPANYL)BUTYRAT
C3272985|T121||RXNORM|1H-AZEPINE-1-BUTANOIC ACID, HEXAHYDRO-, 3-(1,2-DIMETHYLHEPTYL)-7,8,9,10-TETRAHYDRO-6,6,9-TRIMETHYL-6H-DIBENZO(B,D)PYRAN-1-YL ESTER
C3272985|T121||RXNORM|SP 175
C3272985|T121||RXNORM|NABAZENIL
C3272985|T121||RXNORM|SP-175
C0006795|T121||RXNORM|CAMAZEPAM
C0006795|T121||RXNORM|CARBAMIC ACID, DIMETHYL-, 7-CHLORO-2,3-DIHYDRO-1-METHYL-2-OXO-5-PHENYL-1H-1,4-BENZODIAZEPIN-3-YL ESTER
C0006795|T121||RXNORM|3-N,N-DIMETHYLCARBAMOYLOXY-7-CHLORO-5-PHENYL-1-METHYL-1,3-DIHYDRO-2H-1,4-BENZODIAZEPIN-2-ONE
C0055353|T121||RXNORM|2'-CHLORONORDIAZEPAM
C0055353|T121||RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-5-(2-CHLOROPHENYL)-1,3-DIHYDRO-
C0055353|T121||RXNORM|7-CHLORO-5-(2-CHLOROPHENYL) 1,3-DIHYDRO-2H-1,4-BENZODIAZEPIN-2-ONE
C0055353|T121||RXNORM|CHLORDEMETHYLDIAZEPAM
C0055353|T121||RXNORM|CHLORDESMETHYLDIAZEPAM
C0055353|T121||RXNORM|CHLORODESMETHYLDIAZEPAM
C0055353|T121||RXNORM|DELORAZEPAM
C0055353|T121||RXNORM|2-CHLORONORDIAZEPAM
C0055353|T121||RXNORM|B1, BENZODIAZEPINE
C0055353|T121||RXNORM|CL-DMDZ
C0055353|T121||RXNORM|1,3-DIHYDRO-7-CHLORO-5-(O-CHLOROPHENYL)-2H-1,4-BENZODIAZEPIN-2-ONE
C3273839|T121||RXNORM|7-CHLORO-1,3-DIHYDRO-1-METHYL-5-PHENYL-2H-BENZO-1,4-DIAZEPIN-2-ONEMONOHYDROCHLORIDE
C3273839|T121||RXNORM|DIAZEPAM HYDROCHLORIDE
C3273839|T121||RXNORM|DIAZEPAM HCL
C0887259|T121||RXNORM|MONOHYDROCHLORIDE, FLURAZEPAM
C0887259|T121||RXNORM|FLURAZEPAM MONOHYDROCHLORIDE
C0887259|T121||RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-1-(2-(DIETHYLAMINO)ETHYL)-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-, MONOHYDROCHLORIDE
C0060689|T121||RXNORM|7-CHLORO-1-(DIMETHYLPHOSPHINMETHYL)-5-PHENYL-1,3- DIHYDRO-2H-1,4-BENZODIAZEPIN-2-ONE
C0060689|T121||RXNORM|FOSAZEPAM
C0060689|T121||RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-1-((DIMETHYLPHOSPHINYL)METHYL)-1,3-DIHYDRO-5-PHENYL-
C0060689|T121||RXNORM|7-CHLORO-1-((DIMETHYLPHOSPHINYL)METHYL)-1,3-DIHYDRO-5-PHENYL-2H-1,4-BENZODIAZEPIN-2-ONE
C0172965|T121||RXNORM|(1-HYDRAZINOCARBONYL)-7-BROMO-5-PHENYL-1,2-DIHYDRO-3H-1,4-BENZODIAZEPINE-2-ONE
C0172965|T121||RXNORM|GIDAZEPAM
C0069747|T121||RXNORM|BUTANEDIOIC ACID, MONO(7-CHLORO-2,3-DIHYDRO-2-OXO-5-PHENYL-1H-1,4-BENZODIAZEPIN-3-YL) ESTER
C0069747|T121||RXNORM|OXAZEPAM HEMISUCCINATE
C0069747|T121||RXNORM|(RS)-OXAZEPAM H
C0069747|T121||RXNORM|( -)-OXAZEPAM SUCCINATE
C0069747|T121||RXNORM|7-CHLORO-1,3-DIHYDRO-3-HEMISUCCINYLOXY-2H-1,4-BENZODIAZEPIN-2-ONE
C3273842|T121||RXNORM|OXAZEPAM MONOSODIUM SUCCINATE
C0070543|T121||RXNORM|7-BROMO-5-(2-CHLORPHENYL)-1,2-DIHYDRO-3H-1,4-BENZODIAZEPIN-2-ONE
C0070543|T121||RXNORM|FENAZEPAM
C0070543|T121||RXNORM|PHENAZEPAM
C0070543|T121||RXNORM|7-BROMO-5-(2-CHLOROPHENYL) 1,3-DIHYDRO-2H-1,4-BENZODIAZEPIN-2-ONE
C0070543|T121||RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 1,3-DIHYDRO-7-BROMO-5-(2-CHLOROPHENYL)-
C0073389|T121||RXNORM|1-ETHYL-4,6-DIHYDRO-3-METHYL-8-PHENYLPYRAZOLO(4,3-E)(1,4)DIAZEPIN-5(LH)-ONE
C0073389|T121||RXNORM|PYRAZAPON
C0073389|T121||RXNORM|RIPAZEPAM
C0073389|T121||RXNORM|1-ETHYL-4,6-DIHYDRO-3-METHYL-8-PHENYLPYRAZOLO(4,3-E)(1,4)DIAZEPIN-5(1H)-ONE
C0073389|T121||RXNORM|PYRAZOLO(4,3-E)(1,4)DIAZEPIN-5(1H)-ONE, 1-ETHYL-4,6-DIHYDRO-3-METHYL-8-PHENYL-
C3273843|T121||RXNORM|TUCLAZEPAM
C3273843|T121||RXNORM|7-CHLOR-5-(2-CHLORPHENYL)-2,3-DIHYDRO-1-METHYL-1H-1,4-BENZODIAZEPIN-2-METHANOL
C0077789|T121||RXNORM|2-(ALLYLOXY)AMINO 7-CHLORO-5-(O-CHLOROPHENYL)-3H-1, 4-BENZODIAZEPINE
C0077789|T121||RXNORM|ULDAZEPAM
C0077789|T121||RXNORM|2-((ALLYLOXY)AMINO)-7-CHLORO-5-(O-CHLOROPHENYL)-3H-1,4-BENZODIAZEPINE
C1982372|T121||RXNORM|BENZODIAZEPINES &#X7C; VITREOUS FLUID
C1982367|T121||RXNORM|BENZODIAZEPINES &#X7C; GASTRIC FLUID
C1982371|T121||RXNORM|BENZODIAZEPINES &#X7C; URINE
C1982364|T121||RXNORM|BENZODIAZEPINES &#X7C; BLD-SER-PLAS
C1982365|T121||RXNORM|BENZODIAZEPINES &#X7C; BODY FLUID
C2600781|T121||RXNORM|BENZODIAZEPINES.OTHER &#X7C; URINE
C3534272|T121||RXNORM|BENZODIAZEPINES &#X7C; SALIVA
C1972398|T121||RXNORM|QUAZEPAM &#X7C; BLD-SER-PLAS
C1982369|T121||RXNORM|BENZODIAZEPINES &#X7C; MECONIUM
C1982363|T121||RXNORM|BENZODIAZEPINE METABOLITES &#X7C; URINE
C1982370|T121||RXNORM|BENZODIAZEPINES &#X7C; STOOL
C1982368|T121||RXNORM|BENZODIAZEPINES &#X7C; HAIR
C1982373|T121||RXNORM|BENZODIAZEPINES &#X7C; XXX
C3711897|T121||RXNORM|R1498 COMPOUND
C3252279|T121||RXNORM|EVACETRAPIB
C3712514|T121||RXNORM|OLANZAPINE PROPAN-2-OL HEMISOLVATE MONOHYDRATE
C2975231|T121||RXNORM|I-BET COMPOUND
C2975231|T121||RXNORM|GSK525762A
C2975231|T121||RXNORM|GSK 525762A
C2975231|T121||RXNORM|GSK-525762A
C2975231|T121||RXNORM|GSK525762
C2975231|T121||RXNORM|IBET COMPOUND
C2975231|T121||RXNORM|BET INHIBITOR GSK525762
C2975231|T121||RXNORM|I-BET762
C3713096|T121||RXNORM|7-CHLORO-2-METHYLAMINO-5-PHENYL-3H-1,4-BENZODIAZEPINE-4-OXIDE
C3712513|T121||RXNORM|OLANZAPINE PROPAN-2-ONE HEMISOLVATE MONOHYDRATE
C3491461|T121||RXNORM|PF-184563
C3177676|T121||RXNORM|7-METHOXY-8-(5-(4-(1,3-BENZOTHIAZOL-2-YL)-2-METHOXYPHENOXY)PENTYL)OXY-(11AS)1,2,3,11A-TETRA-HYDRO-5H-PYRROLO(2,1-C)(1,4)BENZODIAZEPIN-5-ONE
C3177676|T121||RXNORM|7-MB-MP-PB CPD
C3712515|T121||RXNORM|2-METHYL-4-(4-METHYLPIPERAZIN-1-YL)-10H-THIENO(2,3-B)(1,5)BENZODIAZEPINE
C3181149|T121||RXNORM|8-ETHYNYL-6-(2'-PYRIDINE)-4H-2,5,10B-TRIAZABENZO(E)AZULENE-3-CARBOXYLIC ACID ETHYL ESTER
C3829073|T121||RXNORM|MIDAZOLAM-CONTAINING BUCCAL LIQUID
C3851482|T121||RXNORM|LIMAZEPINE H
C3851484|T121||RXNORM|LIMAZEPINE G
C3886229|T121||RXNORM|N-P-TOSYL-1,5-BENZODIAZEPIN-2-ONE
C3886414|T121||RXNORM|PGW5 COMPOUND
C3884716|T121||RXNORM|OXOPROTHRACARCIN
C3884297|T121||RXNORM|JM-20 COMPOUND
C3884297|T121||RXNORM|3-ETHOXYCARBONYL-2-METHYL-4-(2-NITROPHENYL)-4,11-DIHYDRO-1H-PYRIDO(2,3-B)(1,5)BENZODIAZEPINE
C3885219|T121||RXNORM|QH-II-66
C4079047|T121||RXNORM|DIETHYL-(Z)-2-(5,7-DIPHENYL-1,3,4-OXADIAZEPIN-2-YL)-2-BUTENEDIOATE
C0699927|T121||RXNORM|ROHYPNOL
C0699927|T121||RXNORM|ROHYPNOL (NOT APPROVED FOR USE IN U.S.)
C0699927|T121||RXNORM|ROHYPNOL (NOT APPROVED FOR USE IN U.S.) 
C0699927|T121||RXNORM|ROHIPNOL
C0699927|T121||RXNORM|ROCHE BRAND OF FLUNITRAZEPAM
C0699927|T121||RXNORM|NARCOZEP
C0069749|T121||RXNORM|10-CHLORO-2,3,7,11B-TETRAHYDRO-2-METHYL-11B-PHENYLBENZO(6,7)(1,4)DIAZEPINO(5,4-B) OXAZOL-6-ONE
C0069749|T121||RXNORM|OXAZOLAM
C0069749|T121||RXNORM|OXAZOLAZEPAM
C0060485|T121||RXNORM|1-METHYL-5-(2-FLUOROPHENYL)-7-CHLORO-1,3-DIHYDRO-2H-(1,4)BENZODIAZEPIN-2-ONE
C0060485|T121||RXNORM|7-CHLORO-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-1-METHYL-2H-1,4-BENZODIAZEPIN-2-ONE
C0060485|T121||RXNORM|FLUDIAZEPAM
C0060485|T121||RXNORM|FLUDIAZEPAN
C0054826|T121|20342|RXNORM|5-(3-(4-PIPERIDINO-4-CARBAMOYLPIPERIDINO)PROPYL)- 10,11-DIHYDRO-5(H)-DIBENZ(B,F)AZEPINE|CARPIPRAMINE
C0054826|T121|20342|RXNORM|CARBADIPIMIDINE|CARPIPRAMINE
C0054826|T121|20342|RXNORM|CARPIPRAMINE|CARPIPRAMINE
C0114875|T121||RXNORM|1-(2-HYDROXYETHYL)-3-HYDROXY-7-CHLORO-1,3-DIHYDRO-5-(O-FLUOROPHENYL)-2H-1,4-BENZODIAZEPIN-2-ONE
C0114875|T121||RXNORM|DOXEFAZEPAM
C0603384|T121||RXNORM|7-CHLORO-5-(2-CHLOROPHENYL)-1,3--DIHYDRO-3-HYDROXY-1-(2-HYDROXYETHYL)-2H-1,4-BENZODIAZEPIN-2-ONE
C0603384|T121||RXNORM|N-(2-HYDROXYETHYL)LORAZEPAM
C0604445|T121||RXNORM|7-CHLORO-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-1-(2-(METHYLSULFONYL)ETHYL)-2H-1,4-BENZODIAZEPIN-2-ONE
C0604445|T121||RXNORM|ID 622
C0604445|T121||RXNORM|ID-622
C0604760|T121||RXNORM|2H-1,5-BENZODIAZEPIN-2-ONE, 8-CHLORO-1,3,4,5-TETRAHYDRO-1-PHENYL-
C0604760|T121||RXNORM|8-CHLORO-1-PHENYL-2,3,4,5-TETRAHYDRO-1H-1,5-BENZODIAZEPIN-2-ONE
C0076784|T121|38365|RXNORM|1-(3,4-DIMETHOXYPHENYL)-5-ETHYL-7,8-DIMETHOXY- 4-METHYL-5H-2,3-BENZODIAZEPINE|TOFISOPAM
C0076784|T121|38365|RXNORM|TOFISOPAM|TOFISOPAM
C0076784|T121|38365|RXNORM|TOFIZOPAM|TOFISOPAM
C0076784|T121|38365|RXNORM|1-(3,4-DIMETHOXYPHENYL)-5-ETHYL-7,8-DIMETHOXY-4-METHYL-5H-2,3-BENZODIAZEPINE|TOFISOPAM
C0060593|T121||RXNORM|10-CHLORO-11B-(2'-FLUOROPHENYL)-2,3,5,6,7,11B-HEXAHYDRO-7-(2''-HYDROXYETHYL)BENZO(6,7)-1,4-DIAZEPINO(5,4-B)OXAZOL-6-ONE
C0060593|T121||RXNORM|10-CHLORO-11B-(2-FLUOROPHENYL)-2,3,7,11B-TETRAHYDRO-7-(2-HYDROXYETHYL)OXAZOLO(3,2-D)(1,4)BENZODIAZEPIN-6(5H)-ONE
C0060593|T121||RXNORM|FLUTAZOLAM
C0076658|T121||RXNORM|2-METHYLDIETHYLAMINOETHYL-4-P-PHENYLTHIOPHENYL-3H- (1,5)BENZODIAZEPINE IODIDE
C0076658|T121||RXNORM|THIABENZONIUM IODIDE
C0076658|T121||RXNORM|TIBENZONIUM IODIDE
C0076658|T121||RXNORM|TIBEZONIUM
C0076658|T121||RXNORM|DIETHYLMETHYL(2-((4-(P-(PHENYLTHIO)PHENYL)-3H-1,5-BENZODIAZEPIN-2-YL)THIO)ETHYL)AMMONIUM
C0063325|T121||RXNORM|ID 690
C0063325|T121||RXNORM|ID-690
C0606744|T121||RXNORM|7-CHLORO-5-(2-CHLOROPHENYL)-1,3-DIHYDRO-1-METHYL-3-(4-MORPHOLINYLMETHYLENE)-2H-1,4-BENZODIAZEPIN-2-ONE
C0606744|T121||RXNORM|AX-A411-BS
C0055866|T121||RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-1-(2-(CYCLOPROPYLMETHOXY)ETHYL)-1,3-DIHYDRO-5-PHENYL-
C0055866|T121||RXNORM|7-CHLORO-1,3-DIHYDRO-1-((2-CYCLOPROPYLMETHOXY)ETHYL)-5-PHENYL-2H-1,4-BENZODIAZEPIN-2-ONE
C0055866|T121||RXNORM|CLAZEPAM
C0073449|T121||RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 1,3-DIHYDRO-1-(METHOXYMETHYL)-7-NITRO-5-PHENYL-
C0073449|T121||RXNORM|RO 06-9098-000
C0132831|T121||RXNORM|N-DESALKYL-2-OXOQUAZEPAM
C0132831|T121||RXNORM|7-CHLORO-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-2H-1,4- BENZODIAZEPIN-2-ONE
C0132831|T121||RXNORM|NORFLUTOPRAZEPAM
C0132831|T121||RXNORM|NORFLUDIAZEPAM
C0132831|T121||RXNORM|NORFLURAZEPAM
C0073528|T121||RXNORM|5-(2-FLUOROPHENYL)-1,3-DIHYDRO-1-METHYL-2H-1,4- BENZODIAZEPIN-2-ONE
C0073528|T121||RXNORM|RO 5-3438
C0092802|T121||RXNORM|2-CHLORODIAZEPAM
C0092802|T121||RXNORM|2H-1,4-BENZODIAZEPIN-2-ONE, 7-CHLORO-5-(2-CHLOROPHENYL)-1,3-DIHYDRO-1-METHYL-
C0067928|T121||RXNORM|1H-1,5-BENZODIAZEPINE-2,4(3H,5H)-DIONE, 8-CHLORO-1-PHENYL-
C0067928|T121||RXNORM|DEMETHYLCLOBAZAM
C0067928|T121||RXNORM|N-DESMETHYLCLOBAZAM
C0067928|T121||RXNORM|NORCLOBAZAM
C0611677|T121||RXNORM|SAS 646
C0611797|T121||RXNORM|KA 2547
C0611797|T121||RXNORM|KA-2547
C0056431|T121||RXNORM|CP 1414 S
C0056431|T121||RXNORM|CP 1414S
C0056431|T121||RXNORM|CP-1414 S
C0616152|T121||RXNORM|4,5-DIHYDRO-2,3-DIMETHYL-4-PHENYL-3H-1,3-BENZODIAZEPINE
C0616486|T121||RXNORM|PSYTON
C0076670|T121||RXNORM|1-METHYL-2-(3-THIENYLCARBONYL)AMINOMETHYL-5-(2-FLUOROPHENYL)-H-2,3-DIHYDRO-1,4-BENZODIAZEPINE
C0076670|T121||RXNORM|3-THIOPHENECARBOXAMIDE, N-((5-(2-FLUOROPHENYL)-2,3-DIHYDRO-1-METHYL-1H-1,4-BENZODIAZEPIN-2-YL)METHYL)-
C0076670|T121||RXNORM|TIFLUADOM
C0076670|T121||RXNORM|TITFLUADOM
C0074103|T121||RXNORM|SC 32855
C0074103|T121||RXNORM|SC-32855
C0617110|T121||RXNORM|5H-PYRROLO(2,1-C)(1,4)BENZODIAZEPIN-5-ONE, 2-ETHYLIDENE-1,2,3,11A-TETRAHYDRO-, (+)-
C0617110|T121||RXNORM|PROTHRACARCIN
C0052237|T121||RXNORM|1,3,4,14B-TETRAHYDRO-2-METHYL-10H-PYRAZINO-(1,2-A)PYRROLO(2,1-C)(1,4)BENZODIAZEPINE
C0052237|T121||RXNORM|APTAZAPINE
C0052237|T121||RXNORM|2H,10H-PARAZINO(1,2-A)PYRROLO(2,1-C)(1,4)BENZODIAZEPINE,1,3,4,14B-TETRAHYDRO-2-METHYL-
C0047483|T121||RXNORM|3-HYDROXYPHENAZEPAM
C0047483|T121||RXNORM|3-OXYFENAZEPAM
C0061841|T121||RXNORM|GP 55-129
C0061841|T121||RXNORM|GP 55129
C0061841|T121||RXNORM|GP-55129
C0073469|T121||RXNORM|RO 14-7437
C0073469|T121||RXNORM|RO-14-7437
C0093602|T121||RXNORM|2-OXOQUAZEPAM
C0093602|T121||RXNORM|2OXOQUAZ
C0093602|T121||RXNORM|7-CHLORO-1-(2,2,2-TRIFLUOROETHYL)-1,3-DIHYDRO-5-(2-FLUOROPHENYL)-2H-1,4-BENZODIAZEPIN-2-ONE
C0619423|T121||RXNORM|SCH 23-324
C0619423|T121||RXNORM|SCH-23-324
C0619423|T121||RXNORM|SCH 23324
C0147987|T121||RXNORM|1-METHYL-4-CARBAMOYL-5-PHENYL-7-CHLORO-1,3,4,5-TETRAHYDRO-2H-1,4-BENZODIAZEPINE-2-ONE
C0147987|T121||RXNORM|4H-1,4-BENZODIAZEPINE-4-CARBOXAMIDE, 7-CHLORO-1,2,3,5-TETRAHYDRO-1-METHYL-2-OXO-5-PHENYL-
C0147987|T121||RXNORM|UXEPAM
C0099755|T121||RXNORM|7-CHLORO-5-(2-FLUOROPHENYL) 2,3-DIHYDRO-2-OXO-1H-1,4-BENZODIAZEPINE-3-CARBOXYLIC ACID
C0099755|T121||RXNORM|LOFLAZEPIC ACID
C0621265|T121||RXNORM|LEPIRAZEPAM
C0055302|T121||RXNORM|1,2,3,11A-TETRAHYDRO-2,8-DIHYDROXY-7-METHOXY-5H-PYRROLO(2,1-C)(1,4)-BENZODIAZEPIN-5-ONE
C0055302|T121||RXNORM|5H-PYRROLO(2,1-C)(1,4)BENZODIAZEPIN-5-ONE, 1,2,3,11A-TETRAHYDRO-2,8-DIHYDROXY-7-METHOXY-, (2S-TRANS)-
C0055302|T121||RXNORM|CHICAMYCIN B
C0055301|T121||RXNORM|1,2,3,10,11A-PENTAHYDRO-2,8-DIHYDROXY-7,11-DIMETHOXY-5H-PYRROLO(2,1-C)(1,4)-BENZODIAZEPIN-5-ONE
C0055301|T121||RXNORM|5H-PYRROLO(2,1-C)(1,4)BENZODIAZEPIN-5-ONE, 1,2,3,10,11,11A-HEXAHYDRO-2,8-DIHYDROXY-7,11-DIMETHOXY-, (2S-(2ALPHA,11ALPHA,11ABETA))-
C0055301|T121||RXNORM|CHICAMYCIN A
C0129948|T121||RXNORM|N,N-DIMETHYL-6-PHENYL-11H-PYRIDO(2,3-B)(1,4)BENZODIAZEPIN-11-PROPANAMINE
C0129948|T121||RXNORM|11H-PYRIDO(2,3-B)(1,4)BENZODIAZEPINE-11-PROPANAMINE, N,N-DIMETHYL-6-PHENYL-, (E)-2-BUTENEDIOATE (1:1)
C0129948|T121||RXNORM|TAMPRAMINE FUMARATE
C0073477|T121||RXNORM|4H-IMIDAZO(1,5-A)(1,4)BENZODIAZEPINE-3-CARBOXYLIC ACID, 8-AZIDO-5,6-DIHYDRO-5-METHYL-6-OXO-, (Z,E,E,E,E)-
C0073477|T121||RXNORM|RO 15-4513
C0073477|T121||RXNORM|RO-154513
C0073477|T121||RXNORM|RO15-4513
C0623223|T121||RXNORM|7-CHLORO 5-(2-CHLOROPHENYL)-1,3-DIHYDRO-2H-(1,4)-BENZODIAZEPINE-2-THIONE
C0623223|T121||RXNORM|7-CCDBT
C0073670|T121||RXNORM|1H-IMIDAZO(1,2-A)(1,4)BENZODIAZEPIN-1-ONE, 6-(2-CHLOROPHENYL)-2-((4-ETHYL-1-PIPERAZINYL)METHYLENE)-2,4-DIHYDRO-8-NITRO-, (R-(R*,R*))-2,3-DIHYDROXYBUTANEDIOATE (1:1)
C0073670|T121||RXNORM|RU 32007
C0073670|T121||RXNORM|RU-32007
C0623725|T121||RXNORM|PYRAZINO(1,2-A)(1,4)BENZODIAZEPINE, 1,2,3,4,4A,5-HEXAHYDRO-3-METHYL-7-(2-THIENYL)-
C0623725|T121||RXNORM|KC 5944
C0623725|T121||RXNORM|KC-5944
C0623750|T121||RXNORM|AGAROSE, ((N,N'-1,2-ETHANEDIYLBIS(N-(CARBOXYMETHYL)GLYCINATO))(4-)-N,N',O,O',ON,ON')-, (2S-TRANS)-
C0623750|T121||RXNORM|1012-S-ACETAMIDE ADIPIC HYDRAZIDE SEPHAROSE 4B
C0623750|T121||RXNORM|BAAHS
C0164299|T121||RXNORM|1-(3-CHLOROPHENYL)-4-METHYL-7,8-DIMETHOXY-5H-2,3-BENZODIAZEPINE
C0164299|T121||RXNORM|GIRISOPAM
C0060496|T121||RXNORM|7-FLUORO-2-METHYL-4(4-METHYL-1-PIPERAZINYL)-10H-THIENO(2,3B)(1,5)BENZODIAZEPINE
C0060496|T121||RXNORM|FLUMEZAPINE
C0067931|T121||RXNORM|N-DESMETHYLMETACLAZEPAM
C0073481|T121||RXNORM|RO 16-0521
C0073481|T121||RXNORM|RO-16-0521
C0073481|T121||RXNORM|UREA, N-(6-BROMO-5-(2-CHLOROPHENYL)-2,3-DIHYDRO-1,3-DIMETHYL-2-OXO-1H-1,4-BENZODIAZEPIN-7-YL)-N'-(2-HYDROXY-1-(HYDROXYMETHYL)-1-METHYLETHYL)-, (S)-
C0628287|T121||RXNORM|N-DESMETHYLQUAZEPAM
C0066721|T121||RXNORM|MONO-N-DEMETHYLADINAZOLAM
C0066721|T121||RXNORM|MONO-N-DESMETHYLADIN AZOLAM
C0066721|T121||RXNORM|N-DESMETHYLADINAZOLAM
C0066721|T121||RXNORM|N-DESMETHYLADINAZOLAM MESYLATE
C0066721|T121||RXNORM|N-DESMETHYLADINOZOLAM
C0066721|T121||RXNORM|MONO-N-DEMETHYLADINAZOLAM MESYLATE
C0073534|T121||RXNORM|RO 7-0213
C0073534|T121||RXNORM|RO-7-0213
C0049851|T121||RXNORM|7-BPDBD
C0049851|T121||RXNORM|7-BROMO-5-PHENYL-1,2-DIHYDRO-2H-1,4-BENZODIAZEPIN-2-ONE
C0085056|T121||RXNORM|ZIMET 54-79
C0085056|T121||RXNORM|ZIMET 5479
C0073510|T121||RXNORM|RO 23-0364
C0073510|T121||RXNORM|RO-23-0364
C0632104|T121||RXNORM|N-DEMETHYLTIMELOTEM
C0632104|T121||RXNORM|N-DESMETHYLTIMELOTEM
C0635312|T121||RXNORM|5H-PYRROLO(2,1-C)(1,4)BENZODIAZEPIN-5-ONE, 7-((4,6-DIDEOXY-3-C-METHYL-4-(METHYLAMINO)-ALPHA-L-MANNOPYRANOSYL)OXY)-1,2,3,11A-TETRAHYDRO-2-PROPYLIDENE-
C0635312|T121||RXNORM|SIBANOMICIN
C0636784|T121||RXNORM|AHR 11797
C0636784|T121||RXNORM|AHR-11797
C0044701|T121||RXNORM|1012S
C0044701|T121||RXNORM|COMPOUND 1012S
C0526445|T121||RXNORM|NERISOPAM
C0526445|T121||RXNORM|1-(4-AMINOPHENYL)-4-METHYL-7,8-DIMETHOXY-5H-2,3-BENZODIAZEPINE
C0638880|T121||RXNORM|6H-IMIDAZO(1,5-A)(1,4)BENZODIAZEPIN-6-ONE, 3-(5-CYCLOPROPYL-1,2,4-OXADIAZOL-3-YL)-4,5-DIHYDRO-5-METHYL-
C0638880|T121||RXNORM|FG 8119
C0638880|T121||RXNORM|FG-8119
C0062021|T121||RXNORM|BENZENAMINE, 4-(8-METHYL-9H-1,3-DIOXOLO(4,5-H)(2,3)BENZODIAZEPIN-5-YL)-
C0062021|T121||RXNORM|GYKI 52466
C0062021|T121||RXNORM|GYKI-52466
C0639138|T121||RXNORM|ACETAMIDE, 2-(7-BROMO-5-(2-FLUOROPHENYL)-1,3-DIHYDRO-1-METHYL-2H-1,4-BENZODIAZEPIN-2-YLIDENE)-, (E)-
C0639138|T121||RXNORM|KC 2846
C0639138|T121||RXNORM|KC-2846
C0072934|T121||RXNORM|R 82150
C0072934|T121||RXNORM|R-82150
C0072934|T121||RXNORM|R82150
C0083173|T121||RXNORM|6H-IMIDAZO(1,5-A)(1,4)BENZODIAZEPIN-6-ONE, 7-CHLORO-4,5-DIHYDRO-5-METHYL-3-(5-(1-METHYLETHYL)-1,2,4-OXADIAZOL-3-YL)-
C0083173|T121||RXNORM|L 663581
C0083173|T121||RXNORM|L-663581
C0641973|T121||RXNORM|GYKI 52713
C0641973|T121||RXNORM|GYKI-52713
C0643367|T121||RXNORM|2-HYDROXY-4-METHYLPYRIMIDO(4,5-B)(1,5)BENZODIAZEPIN-5-ONE
C0643367|T121||RXNORM|HMPBD
C0084281|T121||RXNORM|IMIDAZO(4,5,1-JK)(1,4)BENZODIAZEPINE-2(1H)-THIONE, 9-CHLORO-4,5,6,7-TETRAHYDRO-5-METHYL-6-(3-METHYL-2-BUTENYL)-, (S)-
C0084281|T121||RXNORM|R 82913
C0084281|T121||RXNORM|R-82913
C0084281|T121||RXNORM|R82913
C0645521|T121||RXNORM|QUINAZOLINO(3',2':1,6)PYRIDO(2,3-B)(1,4)BENZODIAZEPINE-9,16-DIONE, 6,7,7A,8-TETRAHYDRO-, (-)-
C0645521|T121||RXNORM|AURANTHINE
C0140776|T121||RXNORM|RO 24-7429
C0140776|T121||RXNORM|RO-24-7429
C0109226|T121||RXNORM|CGS 15040A
C0109226|T121||RXNORM|CGS-15040A
C0109226|T121||RXNORM|2H,10H-INDOLO(2,1-C)PYRAZINO(1,2-A)(1,4)BENZODIAZEPINE-16-CARBOXYLIC ACID, 1,3,4,16B-TETRAHYDRO-2-METHYL-, METHYL ESTER, MONOHYDROCHLORIDE
C0147541|T121||RXNORM|U-46,195
C0147541|T121||RXNORM|U46,195
C0147541|T121||RXNORM|U-46195
C0147541|T121||RXNORM|U 46195
C0649797|T121||RXNORM|7-(4-BROMOPHENYL)-8-PHENOXY-4,5-BENZO-3-AZA-2-NONEM
C0649797|T121||RXNORM|7-BPPBAN
C0168533|T121||RXNORM|BIM-18216
C0168533|T121||RXNORM|BIM 18216
C0653743|T121||RXNORM|BIOTIN-(N-(2-AMINOETHYL)-8-CHLORO-6-(2-CHLOROPHENYL)-4H(1,2,4)TRIAZOLO(3,4-A)(1,4)BENZODIAZEPINE-2-CARBOXAMIDE) CONJUGATE
C0653743|T121||RXNORM|BIOTINYLATED 1012-S CONJUGATE
C0653743|T121||RXNORM|BIOTIN-1012-S
C0656355|T121||RXNORM|12,13,14,14A-TETRAHYDRO-9H,11H-PYRAZINO(2,1-C)PYRROLO(1,2-A)(1,4)BENZODIAZEPINE
C0656355|T121||RXNORM|ISONORAPTAZEPINE
C0213386|T121||RXNORM|GYKI-53655
C0213386|T121||RXNORM|GYKI 53655
C0660404|T121||RXNORM|U-51477
C0660404|T121||RXNORM|U 51477
C0660406|T121||RXNORM|U-34599
C0660406|T121||RXNORM|U 34599
C0660406|T121||RXNORM|4H-(1,2,4)TRIAZOLO(4,3-A)(1,4)DIAZEPINE, 8-CHLORO-1,4-DIMETHYL-6-PHENYL-
C0219102|T121||RXNORM|6-(2-BROMOPHENYL)-8-FLUORO-4-H-IMIDAZO(1,5-A)(1-4)BENZODIAZEPINE-3-CARBOXAMIDE
C0219102|T121||RXNORM|IMIDAZENIL
C0661222|T121||RXNORM|4-BDBDT
C0661222|T121||RXNORM|4-(3-BROMOPHENYL)-1,3-DIHYDRO-2H-1,5-BENZODIAZEPIN-2-THIONE
C0249301|T121||RXNORM|TRIPITRAMINE
C0250723|T121||RXNORM|GYKI 53405
C0250723|T121||RXNORM|GYKI-53405
C0252422|T121||RXNORM|9A,9B,14B,14C-TETRAPHENYLBENZO(1,2-H-4,5-H')DICYCLOHEPTA(1,2,3-BC)GLYCOLURIL
C0252422|T121||RXNORM|TPB-DCHU
C0252468|T121||RXNORM|R 86183
C0252468|T121||RXNORM|R-86183
C0252468|T121||RXNORM|R86183
C0254734|T121||RXNORM|L 368935
C0254734|T121||RXNORM|L-368,935
C0254734|T121||RXNORM|UREA, N-(2,3-DIHYDRO-1-(2-METHYLPROPYL)-2-OXO-5-PHENYL-1H-1,4-BENZODIAZEPIN-3-YL)-N'-(3-(1H-TETRAZOL-5-YL)PHENYL)-, (R)-
C0254783|T121||RXNORM|YM 022
C0254783|T121||RXNORM|YM-022
C0254783|T121||RXNORM|YM022
C0254783|T121||RXNORM|UREA, N-(2,3-DIHYDRO-1-(2-(2-METHYLPHENYL)-2-OXOETHYL)-2-OXO-5-PHENYL-1H-1,4-BENZODIAZEPIN-3-YL)-N'-(3-METHYLPHENYL)-, (R)-
C0257405|T121||RXNORM|BENZOMALVIN A
C0257406|T121||RXNORM|BENZOMALVIN B
C0257407|T121||RXNORM|BENZOMALVIN C
C0289297|T121||RXNORM|1,1-BIS(((5,11-DIHYDRO-6-OXO-6H-PYRIDO(2,3-B)(1,4)BENZODIAZEPIN-11-YL)CARBONYL)METHYL)-8,17-DIMETHYL-1,8,17,24-TETRAAZATETRACOSANE
C0289297|T121||RXNORM|DIPITRAMINE
C0290224|T121||RXNORM|BZA 5B
C0290224|T121||RXNORM|BZA-5B
C0294497|T121||RXNORM|R 79882
C0294497|T121||RXNORM|R-79882
C0294497|T121||RXNORM|R79882
C0383534|T121||RXNORM|RO 14-5974
C0383534|T121||RXNORM|RO 145974
C0383534|T121||RXNORM|RO-14-5974
C0383534|T121||RXNORM|RO-145974
C0383538|T121||RXNORM|RO 19-0528
C0383538|T121||RXNORM|RO 190528
C0383538|T121||RXNORM|RO-19-0528
C0383538|T121||RXNORM|RO-190528
C0385516|T121||RXNORM|8-CHLORO-TIBO
C0385516|T121||RXNORM|8-CHLOROTETRAHYDROIMIDAZO(4,5,1-JK)(1,4)-BENZODIAZEPIN-2(1H)-THIONE
C0385516|T121||RXNORM|TIVIRAPINE
C0385516|T121||RXNORM|(S)-8-CHLORO-4,5,6,7-TETRAHYDRO-5-METHYL-6-(3-METHYL-2-BUTENYL)IMIDAZO(4,5,1-JK)(1,4)BENZODIAZEPINE-2(1H)-THIONE
C0077112|T121||RXNORM|1-METHYL-5-PHENYL-7-TRIFLUOROMETHYL-(1H)-1,5-BENZODIAZEPINE-2,4-(3H,5H)DIONE
C0077112|T121||RXNORM|TRIFLUBAZAM
C0391429|T121||RXNORM|NNC 13-8241
C0391429|T121||RXNORM|NNC-13-8241
C0531537|T121||RXNORM|9-AMINO-11-ETHYL-6-METHYLPYRIDO(2,3-B)(1,4)BENZODIAZEPIN-5-ONE
C0531537|T121||RXNORM|9-AMINONEVIRAPINE
C0532436|T121||RXNORM|SARMAZENIL
C0532436|T121||RXNORM|ETHYL 7-CHLORO-5,6-DIHYDRO-5-METHYL-6-OXO-4H-IMIDAZO-(1,5-A)(1,4)BENZODIAZEPINE-3-CARBOXYLATE
C0536423|T121||RXNORM|1-(3-(N'-(4-(2-(N-AMINOSULFONYLAMIDINO)ETHYLTHIOMETHYL)THIAZOL-2-YL)GUANIDINOMETHYL)PHENYL)-3-(1-METHYL-2-OXO-5-PHENYL-2,3-DIHYDRO-1H-1,4-BENZODIAZEPIN-3-YL)UREA
C0536423|T121||RXNORM|AETGPMOPDBU
C0537435|T121||RXNORM|GYKI 53665
C0537435|T121||RXNORM|GYKI-53665
C0538541|T121||RXNORM|EGIS 7649
C0538541|T121||RXNORM|EGIS-7649
C0538838|T121||RXNORM|S 8510
C0538838|T121||RXNORM|S-8510
C0540410|T121||RXNORM|7-CHLORO-1,3-DIHYDRO-3-HEMISUCCINYLOXY-5-PHENYL-1,4-BENZODIAZEPIN-2-ONE
C0541175|T121||RXNORM|RO 48-6792
C0541355|T121||RXNORM|4,5,6,7-TETRAHYDRO-5-METHYLIMIDAZO(4,5,1-JK)(1,4)BENZODIAZEPIN-2(1H)-ONE
C0541355|T121||RXNORM|4567-TMB
C0667114|T121||RXNORM|7-CHLORO-1,3-DIHYDRO-1-(1,1-DIMETHYLETHYL)-5-(2-FLUOROPHENYL)-2H-1,4-BENZODIAZEPIN-2-ONE
C0667114|T121||RXNORM|7-CDDFB
C0667714|T121||RXNORM|RY80
C0667714|T121||RXNORM|RY 80
C0670249|T121||RXNORM|RO 48-8684
C0670792|T121||RXNORM|BDA 452
C0670792|T121||RXNORM|BDA-452
C0670792|T121||RXNORM|BDA452
C0670796|T121||RXNORM|BDA 250
C0670796|T121||RXNORM|BDA-250
C0670796|T121||RXNORM|BDA250
C0755389|T121||RXNORM|L-364,373
C0755389|T121||RXNORM|L 364373
C0755389|T121||RXNORM|L364373
C0756415|T121||RXNORM|RY-008, IMIDAZOBENZODIAZEPINE
C0756415|T121||RXNORM|RY 008
C0756868|T121||RXNORM|1-(4'-AMINOPHENYL)-3,5-DIHYDRO-7,8-DIMETHOXY-4H-2M3-BENZODIAZEPINE-4-THIONE
C0756868|T121||RXNORM|1-NHPH-DDBT
C0759918|T121||RXNORM|RL 218
C0759918|T121||RXNORM|RL-218
C0759921|T121||RXNORM|RL 236
C0759921|T121||RXNORM|RL-236
C0760184|T121||RXNORM|TS 941
C0760184|T121||RXNORM|TS-941
C0760184|T121||RXNORM|TS941
C0760535|T121||RXNORM|L 735,821
C0760535|T121||RXNORM|L-735,821
C0760535|T121||RXNORM|L 735821
C0760535|T121||RXNORM|L-735821
C0761079|T121||RXNORM|CR 2945
C0761079|T121||RXNORM|CR-2945
C0761079|T121||RXNORM|CR2945
C0764989|T121||RXNORM|TARAZEPIDE
C0764989|T121||RXNORM|(-)-N-((S)-2,3-DIHYDRO-1-METHYL-2-OXO-5-PHENYL-1H-1,4-BENZODIAZEPIN-3-YL)-5,6-DIHYDRO-4H-PYRROLO(3,2,1-IJ)QUINOLINE-2-CARBOXAMIDE
C0765506|T121||RXNORM|DMP 406
C0765506|T121||RXNORM|DMP-406
C0766295|T121||RXNORM|GYKI 53784
C0766295|T121||RXNORM|GYKI-53784
C0768431|T121||RXNORM|LE 511
C0768431|T121||RXNORM|LE-511
C0768431|T121||RXNORM|LE511
C0907968|T121||RXNORM|1-(4'-AMINOPHENYL)-3,5-DIHYDRO-7,8--DIMETHOXY-2,3-BENZODIAZEPINE
C0907968|T121||RXNORM|2,3-BZ CPD
C0908355|T121||RXNORM|VP 339
C0908355|T121||RXNORM|VP-339
C0908356|T121||RXNORM|VP 365
C0908356|T121||RXNORM|VP-365
C0908672|T121||RXNORM|7-BROMO-5-PHENYL-DIHYDRO-3H-1,4-BENZODIAZEPINE
C0908672|T121||RXNORM|7-BROMO-PHHBDZ
C0909356|T121||RXNORM|CL 385,004
C0909356|T121||RXNORM|CL 385004
C0909356|T121||RXNORM|CL-385,004
C0909356|T121||RXNORM|CL-385004
C0914661|T121||RXNORM|TETRAZOLO(1,5-A)(1,4)BENZODIAZEPINE
C0914662|T121||RXNORM|TRIAZOLO(4,3-D)BENZODIAZEPINE
C0960422|T121||RXNORM|LOTRAFIBAN
C0961688|T121||RXNORM|4-PHENYL-2-TRICHLOROMETHYL-3H-1,5-BENZODIAZEPINE
C1306120|T121||RXNORM|7-CYANO-2,3,4,5-TETRAHYDRO-1-(1H-IMIDAZOL-4-YLMETHYL)-3-(PHENYLMETHYL)-4-(2-THIENYLSULFONYL)-1H-1,4-BENZODIAZEPINE
C0963297|T121||RXNORM|1,5-BENZODIAZEPIN-2-ONE
C0963508|T121||RXNORM|GYKI 47261
C0963508|T121||RXNORM|GYKI-47261
C0967164|T121||RXNORM|1,2,3,4-TETRAHYDROBENZO(E)(1,4)DIAZEPIN-5-ONE
C0967164|T121||RXNORM|TH-BDAO
C0969588|T121||RXNORM|8-FLUORO-12-(4-METHYLPIPERAZIN-1-YL)-6H-(1)BENZOTHIENO(2,3-B)(1,5)BENZODIAZEPINE
C0969588|T121||RXNORM|8-FLUORO-12-(4-METHYLPIPERAZIN-1-YL)-6H-(1)BENZOTHIENO(2,3-B)(1,5)BENZODIAZEPINE MALEATE
C0969588|T121||RXNORM|Y 931
C1097584|T121||RXNORM|ETHYL-8-ETHYL-5,6-DIHYDRO-5-METHYL-6-OXO-4H-IMIDAZO(1,5A)(1,4)BENZODIAZEPINE-3-CARBOXYLATE
C1097588|T121||RXNORM|ETADOAIB CPD
C1097588|T121||RXNORM|ETHYL-8-TRIMETHYLSILYL-2-ACETYL-12,12A-DIHYDRO-9-OXO-9H,11H-AZETO(2,1-C)IMIDAZO(1,5A)-1,4-BENZODIAZEPINE
C1098285|T121||RXNORM|BZA-2B
C1098285|T121||RXNORM|CYS-(N-METHYL)-3-AMINO-1-CARBOXYMETHYL-2,3-DIHYDRO-5-PHENYL-1H-1,4-BENZODIAZEPIN-2-ONE-MET
C1098621|T121||RXNORM|CIRCUMDATIN C
C1434719|T121||RXNORM|PBDS CPD
C1434719|T121||RXNORM|PYRROLO(2,1-C)(1,4)BENZODIAZEPINE
C1136832|T121||RXNORM|BD-1158
C1143145|T121||RXNORM|RY 024
C1143145|T121||RXNORM|RY024
C1143677|T121||RXNORM|3-TERT-BUTOXYCARBONYLAMINO-2-OXO-2,3,4,5-TETRAHYDRO-1,5-BENZODIAZEPINE-1-ACETIC ACID METHYL ESTER
C1143677|T121||RXNORM|BTOTBAM ESTER
C1143762|T121||RXNORM|1-M-6P-TBD
C1143762|T121||RXNORM|1-METHYL-6-PHENYL-4H-S-TRIAZO-(4,3-ALPHA)(1,4)BENZODIAZEPINONE
C1172344|T121||RXNORM|1,4-BENZODIAZEPINE
C1172344|T121||RXNORM|BZ-423
C1172477|T121||RXNORM|6-CHLORO-PPPBD
C1172477|T121||RXNORM|8-CHLORO-6-(4-PHENETHYL-1-PIPERAZINYL)-11H-PYRIDO(2,3-B)(1,4)BENZODIAZEPINE
C1173066|T121||RXNORM|INDIPLON
C1174538|T121||RXNORM|5-P-3-U-BDA
C1174538|T121||RXNORM|5-PHENYL-3-UREIDO-1,5-BENZODIAZEPINE
C1311127|T121||RXNORM|(11AS)-8-HYDROXY-7-METHOXY-1,2,3,11A-TETRAHYDRO-5H-PYRROLO(2,1-C)(1,4)BENZODIAZEPIN-5-ONE
C1311268|T121||RXNORM|TIBO CPD
C1311268|T121||RXNORM|4,5,6,7-TETRAHYDROIMIDAZO-(4,5,1- JK)(1,4)BENZODIAZEPIN-2 (1 H)-ONE
C1311387|T121||RXNORM|8,9-DIMETHOXY-6-(4-BROMOPHENYL)-11H-(1,2,4)TRIAZOLO(4,5-C)(2,3)BENZODIAZEPIN-3(2H)-ONE
C1311387|T121||RXNORM|8,9-DIMETHOXY-BTBDO
C1313512|T121||RXNORM|1-(4-DIMETHYLAMINOMETHYLPHENYL)-8,9-DIHYDRO-7H-2,7,9A-BENZO(CD)AZULEN-6-ONE
C1435117|T121||RXNORM|2,3,4,5-TETRAHYDRO-1-(1H-IMIDAZOL-4-YLMETHYL)-4-(2-BIPHENYLYLCARBONYL)-1H-1,4-BENZODIAZEPINE
C1454299|T121||RXNORM|BMS-225975
C1454299|T121||RXNORM|BMS225975
C1505431|T121||RXNORM|GI 181771X
C1505431|T121||RXNORM|GI-181771X
C1505431|T121||RXNORM|GI181771X
C1608551|T121|611247|RXNORM|FLUOXETINE/OLANZAPINE|FLUOXETINE / OLANZAPINE
C1608551|T121|611247|RXNORM|FLUOXETINE / OLANZAPINE|FLUOXETINE / OLANZAPINE
C1608551|T121|611247|RXNORM|FLUOXETINE-OLANZAPINE|FLUOXETINE / OLANZAPINE
C1608551|T121|611247|RXNORM|OLANZAPINE + FLUOXETINE |FLUOXETINE / OLANZAPINE
C1608551|T121|611247|RXNORM|OLANZAPINE + FLUOXETINE|FLUOXETINE / OLANZAPINE
C1608551|T121|611247|RXNORM|OLANZAPINE-FLUOXETINE COMBINATION|FLUOXETINE / OLANZAPINE
C1570489|T121||RXNORM|MMY-SJG COMPOUND
C1571352|T121||RXNORM|FQP-BD CPD
C1571352|T121||RXNORM|FLUOROQUINOLONE-PYRROLO(2,1-C)(1,4)BENZODIAZEPINE
C1611910|T121||RXNORM|2,3-DIMETHYL-6-PHENYL-12H-(1,3)DIOXOLO(4,5-H)IMIDAZO(1,2-C)(2,3)BENZODIAZEPINE
C1615028|T121||RXNORM|EGIS-10608
C1614477|T121||RXNORM|EGIS-8332
C1687864|T121||RXNORM|RY 023
C1686352|T121||RXNORM|6-FLUORO-10-(3-(2-METHOXYETHYL)-4-METHYLPIPERAZIN-1-YL)-2-METHYL-4H-3-THIA-4,9-DIAZABENZO(F)AZULENE
C1698804|T121||RXNORM|RWJ-351647
C1700769|T121||RXNORM|DPBDA CPD
C1700769|T121||RXNORM|5,11-DIHYDRO-PYRIDO(2,3-B)(1,5)BENZODIAZEPINE
C1721896|T121||RXNORM|ALPHA5IA-II
C1871751|T121||RXNORM|RO0281501
C1871751|T121||RXNORM|RO 0281501
C1872487|T121||RXNORM|2-HYDROXYMETHYLOLANZAPINE
C1870086|T121||RXNORM|DRH-417
C1870086|T121||RXNORM|NSC 709119
C1880572|T121||RXNORM|ETHYL CARFLUZEPATE
C1880826|T121||RXNORM|FLUTEMAZEPAM
C1882473|T121||RXNORM|PROFLAZEPAM
C0209249|T121||RXNORM|2-BENZOYL-6-ETHYL-7-METHOXY-5-METHYLIMIDAZOL(1,2-A)PYRIMIDINE
C0209249|T121||RXNORM|METHANONE, (6-ETHYL-7-METHOXY-5-METHYLIMIDAZO(1,2-A)PYRIMIDIN-2-YL)PHENYL-
C0209249|T121||RXNORM|DIVAPLON
C0700528|T121|203173|RXNORM|HYDROCHLORIDE, CHLORDIAZEPOXIDE|CHLORDIAZEPOXIDE HYDROCHLORIDE
C0700528|T121|203173|RXNORM|CHLORDIAZEPOXIDE HYDROCHLORIDE|CHLORDIAZEPOXIDE HYDROCHLORIDE
C0700528|T121|203173|RXNORM|CHLORDIAZEPOXIDE HYDROCHLORIDE |CHLORDIAZEPOXIDE HYDROCHLORIDE
C0700528|T121|203173|RXNORM|CHLORDIAZEPOXIDE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|CHLORDIAZEPOXIDE HYDROCHLORIDE
C0700528|T121|203173|RXNORM|CHLORDIAZEPOXIDE MONOHYDROCHLORIDE|CHLORDIAZEPOXIDE HYDROCHLORIDE
C0700528|T121|203173|RXNORM|MONOHYDROCHLORIDE, CHLORDIAZEPOXIDE|CHLORDIAZEPOXIDE HYDROCHLORIDE
C0700528|T121|203173|RXNORM|CHLORDIAZEPOXIDE HYDROCHLORIDE |CHLORDIAZEPOXIDE HYDROCHLORIDE
C0700528|T121|203173|RXNORM|CHLORDIAZEPOXIDE HYDROCHLORIDE |CHLORDIAZEPOXIDE HYDROCHLORIDE
C0770393|T121|235408|RXNORM|CLORAZEPIC ACID|CLORAZEPIC ACID
C1881125|T121||RXNORM|ICLAZEPAM
C1881782|T121||RXNORM|MENITRAZEPAM
C0071879|T121||RXNORM|3,7-DIHYDRO-5-PHENYL-6,7-DIMETHYLPYRROLE(3,4-E)(1,4)DIAZEPIN-2-(1H)-ONE
C0071879|T121||RXNORM|PREMAZEPAM
C0035766|T121||RXNORM|HYDROCHLORIDE, MEDAZEPAM
C0035766|T121||RXNORM|MEDAZEPAM HYDROCHLORIDE
C0035766|T121||RXNORM|MONOHYDROCHLORIDE, MEDAZEPAM
C0035766|T121||RXNORM|MEDAZEPAM MONOHYDROCHLORIDE
C1880574|T121||RXNORM|ETHYL DIRAZEPATE
C0700457|T121|203128|RXNORM|HYDROCHLORIDE, MIDAZOLAM|MIDAZOLAM HYDROCHLORIDE
C0700457|T121|203128|RXNORM|MIDAZOLAM HYDROCHLORIDE|MIDAZOLAM HYDROCHLORIDE
C0700457|T121|203128|RXNORM|ANXIOLYTICS MIDAZOLAM HYDROCHLORIDE|MIDAZOLAM HYDROCHLORIDE
C0700457|T121|203128|RXNORM|MIDAZOLAM HYDROCHLORIDE |MIDAZOLAM HYDROCHLORIDE
C0700457|T121|203128|RXNORM|MIDAZOLAM HYDROCHLORIDE [CHEMICAL/INGREDIENT]|MIDAZOLAM HYDROCHLORIDE
C0700457|T121|203128|RXNORM|MIDAZOLAM (AS HYDROCHLORIDE)|MIDAZOLAM HYDROCHLORIDE
C0700457|T121|203128|RXNORM|MIDAZOLAM HYDROCHLORIDE |MIDAZOLAM HYDROCHLORIDE
C0700457|T121|203128|RXNORM|MIDAZOLAM HYDROCHLORIDE |MIDAZOLAM HYDROCHLORIDE
C3179470|T121||RXNORM|REMIMAZOLAM
C2000107|T121||RXNORM|4-(2-HYDROXYPHENYL)-2-PHENYL-2,3-DIHYDRO-1H-1,5-BENZODIAZEPINE
C2000107|T121||RXNORM|4-(2-HYDROXYPHENYL)-PDBDZ
C0065086|T121|1310187|RXNORM|LITHIUM BROMIDE|LITHIUM BROMIDE
C0065086|T121|1310187|RXNORM|LITHIUM BROMIDE |LITHIUM BROMIDE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150 MG ORAL CAPSULE|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150MG ORAL CAPSULE|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE, 150 MG ORAL CAPSULE|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM 150 MG ORAL CAPSULE|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150MG CAP|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150MG CAP UD|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150 MILLIGRAM IN 1 CAPSULE ORAL CAPSULE|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE CAP 150 MG|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150 MG ORAL CAPSULE, GELATIN COATED|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150MG CAP,UD [VA PRODUCT]|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150MG CAP,UD|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150MG CAP [VA PRODUCT]|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150 MG ORAL CAPSULE [LITHIUM CARBONATE]|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LICO3 150 MG ORAL CAPSULE|LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150MG CAPSULE |LICO3 150 MG ORAL CAPSULE
C0978225|T121|311355|RXNORM|LITHIUM CARBONATE 150MG CAPSULE|LICO3 150 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE 300 MG ORAL CAPSULE|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE 300MG ORAL CAPSULE|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE, 300 MG ORAL CAPSULE|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM 300 MG ORAL CAPSULE|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE 300MG CAP|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE 300 MILLIGRAM IN 1 CAPSULE ORAL CAPSULE|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE CAP 300 MG|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE 300 MG ORAL CAPSULE, GELATIN COATED|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE 300MG CAP [VA PRODUCT]|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE 300 MG ORAL CAPSULE [LITHIUM CARBONATE]|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LICO3 300 MG ORAL CAPSULE|LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE 300MG CAPSULE |LICO3 300 MG ORAL CAPSULE
C0689383|T121|197889|RXNORM|LITHIUM CARBONATE 300MG CAPSULE|LICO3 300 MG ORAL CAPSULE
C0689384|T121|197890|RXNORM|LITHIUM CARBONATE 300 MG ORAL TABLET|LICO3 300 MG ORAL TABLET
C0689384|T121|197890|RXNORM|LITHIUM CARBONATE 300MG ORAL TABLET|LICO3 300 MG ORAL TABLET
C0689384|T121|197890|RXNORM|LITHIUM CARBONATE, 300 MG ORAL TABLET|LICO3 300 MG ORAL TABLET
C0689384|T121|197890|RXNORM|LITHIUM 300 MG ORAL TABLET|LICO3 300 MG ORAL TABLET
C0689384|T121|197890|RXNORM|LITHIUM CARBONATE 300MG TAB|LICO3 300 MG ORAL TABLET
C0689384|T121|197890|RXNORM|LITHIUM CARBONATE TAB 300 MG|LICO3 300 MG ORAL TABLET
C0689384|T121|197890|RXNORM|LITHIUM CARBONATE 300MG TAB [VA PRODUCT]|LICO3 300 MG ORAL TABLET
C0689384|T121|197890|RXNORM|LICO3 300 MG ORAL TABLET|LICO3 300 MG ORAL TABLET
C0689384|T121|197890|RXNORM|LITHIUM CARBONATE 300MG TABLET |LICO3 300 MG ORAL TABLET
C0689384|T121|197890|RXNORM|LITHIUM CARBONATE 300MG TABLET|LICO3 300 MG ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300 MG ORAL TABLET, EXTENDED RELEASE|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300MG ORAL TABLET, EXTENDED RELEASE|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM 300 MG ORAL TABLET, EXTENDED RELEASE|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300MG SA TAB|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE TAB CR 300 MG|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300MG SLOW RELEASE TABLET|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300 MG ORAL TABLET, FILM COATED, EXTENDED RELEASE|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300MG TAB,SA|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300MG TAB,SA [VA PRODUCT]|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300 MG ORAL TABLET, EXTENDED RELEASE [LITHIUM CARBONATE]|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300 MG ORAL TABLET, FILM COATED, EXTENDED RELEASE [LITHIUM CARBONATE]|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300 MG EXTENDED RELEASE ORAL TABLET|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LICO3 300 MG EXTENDED RELEASE ORAL TABLET|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE, 300 MG ORAL TABLET, EXTENDED RELEASE|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300MG M/R TABLET|LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689385|T121|197891|RXNORM|LITHIUM CARBONATE 300MG M/R TABLET |LICO3 300 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450 MG ORAL TABLET, EXTENDED RELEASE|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450MG ORAL TABLET, EXTENDED RELEASE|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450MG TABLET|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM 450 MG ORAL TABLET, EXTENDED RELEASE|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450MG SA TAB|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE TAB CR 450 MG|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450MG TAB,SA [VA PRODUCT]|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450MG TAB,SA|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450 MG ORAL TABLET, EXTENDED RELEASE [LITHIUM CARBONATE]|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE CR 450MG TABLET |LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE CR 450MG TABLET|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450 MG EXTENDED RELEASE ORAL TABLET|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LICO3 450 MG EXTENDED RELEASE ORAL TABLET|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450 MG ORAL TABLET [LITHIUM CARBONATE ER]|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450MG M/R TABLET|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450MG M/R TABLET |LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE, 450 MG ORAL TABLET, EXTENDED RELEASE|LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450MG M/R TABLET |LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689386|T121|197892|RXNORM|LITHIUM CARBONATE 450MG TABLET |LICO3 450 MG EXTENDED RELEASE ORAL TABLET
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE 600 MG ORAL CAPSULE|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE 600MG ORAL CAPSULE|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE, 600 MG ORAL CAPSULE|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM 600 MG ORAL CAPSULE|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE 600MG CAP|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE 600 MILLIGRAM IN 1 CAPSULE ORAL CAPSULE|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE CAP 600 MG|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE 600 MG ORAL CAPSULE, GELATIN COATED|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE 600MG CAP [VA PRODUCT]|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LICO3 600 MG ORAL CAPSULE|LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE 600MG CAPSULE |LICO3 600 MG ORAL CAPSULE
C0689387|T121|197893|RXNORM|LITHIUM CARBONATE 600MG CAPSULE|LICO3 600 MG ORAL CAPSULE
C0700189|T121|203056|RXNORM|LITHONATE|LITHONATE
C0771417|T121||RXNORM|LITHIUM SALICYLATE
C0700753|T121|203323|RXNORM|ESKALITH|ESKALITH
C0700753|T121|203323|RXNORM|ESCALITH|ESKALITH
C0700751|T121|203321|RXNORM|LITHOBID|LITHOBID
C0700752|T121|203322|RXNORM|LITHANE|LITHANE
C0065091|T121|28815|RXNORM|LITHIUM OROTATE|LITHIUM OROTATE
C2716130|T121||RXNORM|POTASSIUM LITHIUM TITANATE
C1966347|T121|746070|RXNORM|LITHIUM ASPARTATE|LITHIUM ASPARTATE
C1966347|T121|746070|RXNORM|ANTIMANICS LITHIUM ASPARTATE|LITHIUM ASPARTATE
C1966347|T121|746070|RXNORM|LITHIUM ASPARTATE |LITHIUM ASPARTATE
C0689381|T121|756059|RXNORM|LITHIUM 8 MEQ/5 ML ORAL SOLUTION|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8MEQ/5ML ORAL SOLUTION|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 60 MG/ML ORAL SOLUTION|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8MEQ/5ML SF SYRUP|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM HYDROXIDE MONOHYDRATE 8 MEQ IN 5 ML ORAL SOLUTION|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8MEQ/5ML ORAL SYRUP|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8 MEQ/5 ML ORAL SOLUTION|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8MEQ/5ML SYRUP|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8MEQ/5ML (SF) SYRUP|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8MEQ/5ML (SF) SYRUP [VA PRODUCT]|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8MEQ/5ML SYRUP [VA PRODUCT]|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CARBONATE 8 MEQ IN 5 ML ORAL SOLUTION [LITHIUM]|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8MEQ/5ML SOLUTION|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM 8MEQ/5ML ORAL SOLUTION|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM 8MEQ/5ML SOLUTION|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM 8MEQ/5ML SOLN,ORAL|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM 8MEQ/5ML ORAL SOLN|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM 8MEQ/5ML SOLN,ORAL [VA PRODUCT]|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM ION 8 MEQ PER 5 ML ORAL SYRUP|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE EQV TO LITHIUM CARBONATE 300 MG PER 5 ML (LITHIUM ION 8 MEQ PER 5 ML) ORAL SYRUP|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CARBONATE 300 MG IN 5 ML ORAL SOLUTION [LITHIUM]|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 8 MEQ IN 5 ML ORAL SOLUTION|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM ORAL SOLUTION 8 MEQ/5ML|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE 300 MG/5 ML ORAL SYRUP|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM CITRATE, 300 MG/5 ML ORAL SYRUP|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0689381|T121|756059|RXNORM|LITHIUM 300 MG/5 ML ORAL SYRUP|LITHIUM ION 8 MEQ IN 5 ML ORAL SOLUTION
C0693401|T121|199762|RXNORM|LITHIUM CARBONATE 400 MG ORAL TABLET, EXTENDED RELEASE|LICO3 400 MG EXTENDED RELEASE ORAL TABLET
C0693401|T121|199762|RXNORM|LICO3 400 MG EXTENDED RELEASE ORAL TABLET|LICO3 400 MG EXTENDED RELEASE ORAL TABLET
C0693401|T121|199762|RXNORM|LITHIUM CARBONATE 400 MG EXTENDED RELEASE ORAL TABLET|LICO3 400 MG EXTENDED RELEASE ORAL TABLET
C0693401|T121|199762|RXNORM|LITHIUM CARBONATE 400MG M/R TABLET|LICO3 400 MG EXTENDED RELEASE ORAL TABLET
C0693401|T121|199762|RXNORM|LITHIUM CARBONATE 400MG M/R TABLET |LICO3 400 MG EXTENDED RELEASE ORAL TABLET
C0693401|T121|199762|RXNORM|LITHIUM CARBONATE 400MG M/R TABLET |LICO3 400 MG EXTENDED RELEASE ORAL TABLET
C0350511|T121|102547|RXNORM|LITHIUM CARBONATE 104 MG/ML ORAL SOLUTION|LITHIUM CARBONATE 520 MG PER 5 ML ORAL SOLUTION
C0350511|T121|102547|RXNORM|LITHIUM CARBONATE 520 MG PER 5 ML ORAL SOLUTION|LITHIUM CARBONATE 520 MG PER 5 ML ORAL SOLUTION
C0350511|T121|102547|RXNORM|LICO3 104 MG/ML ORAL SOLUTION|LITHIUM CARBONATE 520 MG PER 5 ML ORAL SOLUTION
C0350511|T121|102547|RXNORM|LITHIUM CARBONATE 520MG/5ML SUGAR FREE LIQUID |LITHIUM CARBONATE 520 MG PER 5 ML ORAL SOLUTION
C0350511|T121|102547|RXNORM|LITHIUM CARBONATE 520MG/5ML SUGAR FREE LIQUID|LITHIUM CARBONATE 520 MG PER 5 ML ORAL SOLUTION
C0350511|T121|102547|RXNORM|LITHIUM CARBONATE 520MG/5ML SUGAR FREE LIQUID |LITHIUM CARBONATE 520 MG PER 5 ML ORAL SOLUTION
C0692744|T121|199324|RXNORM|LITHIUM CARBONATE 250 MG ORAL TABLET|LICO3 250 MG ORAL TABLET
C0692744|T121|199324|RXNORM|LICO3 250 MG ORAL TABLET|LICO3 250 MG ORAL TABLET
C0692744|T121|199324|RXNORM|LITHIUM CARBONATE 250MG TABLET|LICO3 250 MG ORAL TABLET
C0692744|T121|199324|RXNORM|LITHIUM CARBONATE 250MG TABLET |LICO3 250 MG ORAL TABLET
C0692744|T121|199324|RXNORM|LITHIUM CARBONATE 250MG TABLET |LICO3 250 MG ORAL TABLET
C0789694|T121|248306|RXNORM|LITHIUM CARBONATE 200 MG EXTENDED RELEASE ORAL TABLET|LICO3 200 MG EXTENDED RELEASE ORAL TABLET
C0789694|T121|248306|RXNORM|LICO3 200 MG EXTENDED RELEASE ORAL TABLET|LICO3 200 MG EXTENDED RELEASE ORAL TABLET
C0789694|T121|248306|RXNORM|LITHIUM CARBONATE 200MG M/R TABLET|LICO3 200 MG EXTENDED RELEASE ORAL TABLET
C0789694|T121|248306|RXNORM|LITHIUM CARBONATE 200MG M/R TABLET |LICO3 200 MG EXTENDED RELEASE ORAL TABLET
C0789694|T121|248306|RXNORM|LITHIUM CARBONATE 200MG M/R TABLET |LICO3 200 MG EXTENDED RELEASE ORAL TABLET
C0302213|T121||RXNORM|LITHIUM SALTS
C0302213|T121||RXNORM|[CN750] LITHIUM SALTS
C0302213|T121||RXNORM|LITHIUM SALT
C0302213|T121||RXNORM|LITHIUM SALT 
C0302213|T121||RXNORM|LITHIUM SALT, NOS
C0065093|T121|28817|RXNORM|LITHIUM SUCCINATE|LITHIUM SUCCINATE
C0065093|T121|28817|RXNORM|LITHIUM SUCCINATE |LITHIUM SUCCINATE
C0065093|T121|28817|RXNORM|LITHIUM SUCCINATE |LITHIUM SUCCINATE
C0065093|T121|28817|RXNORM|ANTIMANICS LITHIUM SUCCINATE|LITHIUM SUCCINATE
C0065093|T121|28817|RXNORM|LITHIUM SUCCINATE |LITHIUM SUCCINATE
C1991690|T121||RXNORM|LITHIUM &#X7C; BODY FLUID
C1991692|T121||RXNORM|LITHIUM &#X7C; RED BLOOD CELLS
C2738318|T121||RXNORM|LITHIUM &#X7C; GASTRIC FLUID
C0366526|T121||RXNORM|LITHIUM:MASS:PT:DOSE:QN
C0366526|T121||RXNORM|LITHIUM DOSE
C0366526|T121||RXNORM|LITHIUM [MASS] OF DOSE
C0366526|T121||RXNORM|LITHIUM:MASS:POINT IN TIME:DOSE MED OR SUBSTANCE:QUANTITATIVE
C1991694|T121||RXNORM|LITHIUM &#X7C; TISSUE AND SMEARS
C1991695|T121||RXNORM|LITHIUM &#X7C; URINE
C1991691|T121||RXNORM|LITHIUM &#X7C; HAIR
C1991696|T121||RXNORM|LITHIUM &#X7C; URINE AND SERUM OR PLASMA
C1991693|T121||RXNORM|LITHIUM &#X7C; SALIVA
C1991688|T121||RXNORM|LITHIUM &#X7C; BLD-SER-PLAS
C3495095|T121|1546265|RXNORM|LITHIUM CATION|LITHIUM CATION
C3495095|T121|1546265|RXNORM|LI+|LITHIUM CATION
C3495095|T121|1546265|RXNORM|LITHIUM ION|LITHIUM CATION
C0303507|T121||RXNORM|LITHIUM ISOTOPE
C0303507|T121||RXNORM|LITHIUM ISOTOPE 
C0078149|T121||RXNORM|VEINOBIASE
C1121051|T121||RXNORM|NOOLITH
C1122689|T121||RXNORM|DYSPROSIUM LITHIUM BORATE GLASS
C1175911|T121||RXNORM|LITAO3
C1175911|T121||RXNORM|LITHIUM TANTALATE OXIDE
C1175913|T121||RXNORM|LIFEPO4
C1311954|T121||RXNORM|LI2ZRO3
C1311954|T121||RXNORM|LITHIUM ZIRCONATE
C1455455|T121||RXNORM|LIMN2O4
C1455455|T121||RXNORM|LITHIUM MANGANESE OXIDE
C0287163|T121|83553|RXNORM|SEROQUEL|SEROQUEL
C0287163|T121|83553|RXNORM|QUETIAPINE (SEROQUEL)|SEROQUEL
