C0015879|T034|LP15568-6|LNC|FERRITIN|FERRITIN
C0373607|T034||LNC|FERRITIN MEASUREMENT
C0015879|T034|LP15568-6|LNC|FERRITIN|FERRITIN
C0015879|T034|LP15568-6|LNC|FERRITINS|FERRITIN
C0015879|T034|LP15568-6|LNC|FERRITINS [CHEMICAL/INGREDIENT]|FERRITIN
C0015879|T034|LP15568-6|LNC|FERRITIN |FERRITIN
C1987810|T034|LP43619-3|LNC|FERRITIN &#X7C; BLD-SER-PLAS|FERRITIN &#X7C; BLD-SER-PLAS
C1987811|T034|LP62244-6|LNC|FERRITIN &#X7C; RED BLOOD CELLS|FERRITIN &#X7C; RED BLOOD CELLS
C0166450|T034||LNC|HEME FERRITIN
C0166450|T034||LNC|HEMOFERRITIN
C0166450|T034||LNC|HAEMOFERRITIN
C0373607|T034||LNC|FERRITIN
C0373607|T034||LNC|FERRITIN MEASUREMENT
C0373607|T034||LNC|TEST;FERRITIN
C0373607|T034||LNC|ASSAY OF FERRITIN
C0373607|T034||LNC|FERRITIN (BLOOD PROTEIN) LEVEL
C0373607|T034||LNC|MEASUREMENT OF FERRITIN
C0373607|T034||LNC|FERRITIN LEVEL
C0373607|T034||LNC|FERRITIN MEASUREMENT 
C0373607|T034||LNC|FERRITIN TEST
C1276043|T034||LNC|PLASMA FERRITIN LEVEL
C1276043|T034||LNC|PLASMA FERRITIN MEASUREMENT 
C1276043|T034||LNC|PLASMA FERRITIN MEASUREMENT
C0696113|T034||LNC|SERUM FERRITIN
C0696113|T034||LNC|SERUM FERRITIN LEVEL 
C0696113|T034||LNC|SERUM FERRITIN LEVEL
C0696113|T034||LNC|SERUM FERRITIN LEVEL 
C0696113|T034||LNC|FERRITIN - SERUM
C0696113|T034||LNC|SERUM FERRITIN MEASUREMENT 
C0696113|T034||LNC|SERUM FERRITIN MEASUREMENT
C0696113|T034||LNC|SERUM FERRITIN EACH TEST
C0696113|T034||LNC|SERUM FERRITIN EA.TST
# C0565897|T034||LNC|IS THIS A RATIO? OR JUST BOTH BEING MEASURED. WOULD EXCLUDE IF THIS IS RETURNING A RATIO.
C0565897|T034||LNC|SERUM FERRITIN/TOTAL IRON BINDING CAPACITY MEASUREMENT
C0565897|T034||LNC|SERUM FERRITIN/TOTAL IRON BINDING CAPACITY MEASUREMENT 
C0565897|T034||LNC|SERUM FERRITIN/TIBC
C0565897|T034||LNC|SERUM FERRITIN/TIBC MEASUREMENT
