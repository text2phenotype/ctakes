C0199967|T037|74287006|SNOMEDCT_US|BLOOD TRANSFUSION|TRANSFUSION OF COAGULATION FACTORS (PROCEDURE)
C0852255|T037||SNOMEDCT_US|BLOOD AND BLOOD PRODUCT TREATMENT
C0481253|T037|216993005|SNOMEDCT_US|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED |CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED (EVENT)
C0481253|T037|216993005|SNOMEDCT_US|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED (EVENT)
C0730400|T037|313039003|SNOMEDCT_US|SOLID ORGAN TRANSPLANT|SOLID ORGAN TRANSPLANT (PROCEDURE)
C0857825|T037||SNOMEDCT_US|INFECTION IN SOLID ORGAN TRANSPLANT RECIPIENTS
C2064857|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN ALBUMIN, NORMAL SERUM 
C2064857|T037||SNOMEDCT_US|PLASMA FRACTIONS, HUMAN ALBUMIN, NORMAL SERUM
C0854629|T037||SNOMEDCT_US|ALLOGENIC BONE MARROW TRANSPLANTATION THERAPY
C0854631|T037||SNOMEDCT_US|CORD BLOOD TRANSPLANT THERAPY
C0015236|T037|39188002|SNOMEDCT_US|EXCHANGE TRANSFUSION, WHOLE BLOOD|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|BLOOD EXCHANGE TRANSFUSION|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EXCHANGE BLOOD TRANSFUSION|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EXCHANGE TRANSFUSION|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EXCHANGE TRANSFUSION |EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EXCHANGE TRANSFUSION OF BLOOD|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EXCHANGE BLOOD TRANSFUSION NOS|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EXCHANGE BLOOD TRANSFUSION NOS |EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EXCHANGE TRANSFUSION, BLOOD|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|TRANSFUSION REPLACEMENT, TOTAL|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EXSANGUINATION TRANSFUSION|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EBT - EXCHANGE BLOOD TRANSFUSION|EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|EXCHANGE TRANSFUSION |EXCHANGE TRANSFUSION (PROCEDURE)
C0015236|T037|39188002|SNOMEDCT_US|TRANSFUSION, EXSANGUINATION|EXCHANGE TRANSFUSION (PROCEDURE)
C0854634|T037||SNOMEDCT_US|MISMATCHED DONOR BONE MARROW TRANSPLANTATION THERAPY
C0371803|T037|180202002|SNOMEDCT_US|EXCHANGE TRANSFUSION, BLOOD; NEWBORN|NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0371803|T037|180202002|SNOMEDCT_US|NEONATAL EXCHANGE BLOOD TRANSFUSION|NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0371803|T037|180202002|SNOMEDCT_US|EXCHANGE TRANSFUSION OF NEWBORN |NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0371803|T037|180202002|SNOMEDCT_US|EXCHANGE TRANSFUSION OF NEWBORN|NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0371803|T037|180202002|SNOMEDCT_US|NEONATAL EXCHANGE TRANSFUSION|NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0371803|T037|180202002|SNOMEDCT_US|BL EXCHANGE/TRANSFUSE NB|NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0371803|T037|180202002|SNOMEDCT_US|EXCHNG TRANSFUSION BLOOD NEWBORN|NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0371803|T037|180202002|SNOMEDCT_US|EXCHANGE BLOOD TRANSFUSION, NEWBORN|NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0371803|T037|180202002|SNOMEDCT_US|EXCHANGE BLOOD TRANSFUSION (NEONATAL)|NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0371803|T037|180202002|SNOMEDCT_US|NEONATAL EXCHANGE TRANSFUSION |NEONATAL EXCHANGE TRANSFUSION (PROCEDURE)
C0199962|T037|71493000|SNOMEDCT_US|PACKED RED BLOOD CELL TRANSFUSION|TRANSFUSION OF PACKED RED BLOOD CELLS (PROCEDURE)
C0199962|T037|71493000|SNOMEDCT_US|TRANSFUSION OF PACKED RED BLOOD CELLS|TRANSFUSION OF PACKED RED BLOOD CELLS (PROCEDURE)
C0199962|T037|71493000|SNOMEDCT_US|RED BLOOD CELL TRANSFUSION|TRANSFUSION OF PACKED RED BLOOD CELLS (PROCEDURE)
C0199962|T037|71493000|SNOMEDCT_US|TRANSFUSION OF PRBC|TRANSFUSION OF PACKED RED BLOOD CELLS (PROCEDURE)
C0199962|T037|71493000|SNOMEDCT_US|INTRAVENOUS BLOOD TRANSFUSION OF PACKED CELLS|TRANSFUSION OF PACKED RED BLOOD CELLS (PROCEDURE)
C0199962|T037|71493000|SNOMEDCT_US|INTRAVENOUS BLOOD TRANSFUSION OF PACKED CELLS |TRANSFUSION OF PACKED RED BLOOD CELLS (PROCEDURE)
C0199962|T037|71493000|SNOMEDCT_US|TRANSFUSION OF PACKED RED BLOOD CELLS |TRANSFUSION OF PACKED RED BLOOD CELLS (PROCEDURE)
C0199962|T037|71493000|SNOMEDCT_US|PRBC TRANSFUSION|TRANSFUSION OF PACKED RED BLOOD CELLS (PROCEDURE)
C0199964|T037|288173003|SNOMEDCT_US|PLASMA EXPANDER TRANSFUSION|PLASMA EXPANDER TRANSFUSION (PROCEDURE)
C0199964|T037|288173003|SNOMEDCT_US|BLOOD EXPANDER TRANSFUS|PLASMA EXPANDER TRANSFUSION (PROCEDURE)
C0199964|T037|288173003|SNOMEDCT_US|BLOOD EXPANDER TRANSFUSION|PLASMA EXPANDER TRANSFUSION (PROCEDURE)
C0199964|T037|288173003|SNOMEDCT_US|TRANSFUSION OF BLOOD EXPANDER|PLASMA EXPANDER TRANSFUSION (PROCEDURE)
C0199964|T037|288173003|SNOMEDCT_US|PLASMA EXPANDER TRANSFUSION |PLASMA EXPANDER TRANSFUSION (PROCEDURE)
C0199964|T037|288173003|SNOMEDCT_US|TRANSFUSION OF BLOOD EXPANDER |PLASMA EXPANDER TRANSFUSION (PROCEDURE)
C0199964|T037|288173003|SNOMEDCT_US|TRANSFUSION OF PLASMA EXPANDER|PLASMA EXPANDER TRANSFUSION (PROCEDURE)
C0199964|T037|288173003|SNOMEDCT_US|TRANSFUSION OF BLOOD EXPANDER, NOS|PLASMA EXPANDER TRANSFUSION (PROCEDURE)
C0199964|T037|288173003|SNOMEDCT_US|TRANSFUSION OF PLASMA EXPANDER, NOS|PLASMA EXPANDER TRANSFUSION (PROCEDURE)
C0032134|T037|20720000|SNOMEDCT_US|CASE REPORTABLE TRANSMISSION, WILL LEAVE ON HERE|PLASMAPHERESIS (PROCEDURE)
C0032134|T037|20720000|SNOMEDCT_US|PLASMAPHERESIS|PLASMAPHERESIS (PROCEDURE)
C0032134|T037|20720000|SNOMEDCT_US|THERAPEU PLASMAPHERESIS|PLASMAPHERESIS (PROCEDURE)
C0032134|T037|20720000|SNOMEDCT_US|PLASMAPHORESIS|PLASMAPHERESIS (PROCEDURE)
C0032134|T037|20720000|SNOMEDCT_US|PLASMA EXCHANGE|PLASMAPHERESIS (PROCEDURE)
C0032134|T037|20720000|SNOMEDCT_US|PLASMAPHERESIS |PLASMAPHERESIS (PROCEDURE)
C0032134|T037|20720000|SNOMEDCT_US|THERAPEUTIC PLASMAPHERESIS|PLASMAPHERESIS (PROCEDURE)
C0032134|T037|20720000|SNOMEDCT_US|THERAPEUTIC PLASMA EXCHANGE|PLASMAPHERESIS (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|PLATELET TRANSFUSION|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|PLATELET TRANSFUSIONS|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|TRANSFUSION, PLATELET|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|TRANSFUSIONS, PLATELET|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|BLOOD PLATELET TRANSFUSIONS|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|PLATELET TRANSFUSION, BLOOD|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|PLATELET TRANSFUSIONS, BLOOD|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|TRANSFUSION, BLOOD PLATELET|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|TRANSFUSIONS, BLOOD PLATELET|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|TRANSFUSION OF PLATELETS |PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|TRANSFUSION OF PLATELETS|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|PLATELET TRANSFUSION |PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|BLOOD PLATELETS--TRANSFUSION|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|BLOOD PLATELET TRANSFUSION|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|TRANSFUSION OF THROMBOCYTES|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|INTRAVENOUS BLOOD TRANSFUSION OF PLATELETS|PLATELET TRANSFUSION (PROCEDURE)
C0086818|T037|12719002|SNOMEDCT_US|INTRAVENOUS BLOOD TRANSFUSION OF PLATELETS |PLATELET TRANSFUSION (PROCEDURE)
C0854635|T037||SNOMEDCT_US|UNRELATED DONOR BONE MARROW TRANSPLANTATION THERAPY
C0919689|T037||SNOMEDCT_US|DONOR LEUKOCYTE INFUSION
C1879316|T037|5447007|SNOMEDCT_US|TRANSFUSION|TRANSFUSION
C1879316|T037|5447007|SNOMEDCT_US|TRANSFUSION |TRANSFUSION
C1879316|T037|5447007|SNOMEDCT_US|TRANSFUSIONS|TRANSFUSION
C1879316|T037|5447007|SNOMEDCT_US|TRANSFUSIONS |TRANSFUSION
C1879316|T037|5447007|SNOMEDCT_US|TRANSFUSION, NOS|TRANSFUSION
C0852255|T037||SNOMEDCT_US|BLOOD AND BLOOD PRODUCT TREATMENT
C4049189|T037||SNOMEDCT_US|IMMUNOADSORPTION THERAPY
C0481253|T037|216993005|SNOMEDCT_US|CONTAMINATED TRANSFUSION|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED (EVENT)
C0481253|T037|216993005|SNOMEDCT_US|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED |CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED (EVENT)
C0481253|T037|216993005|SNOMEDCT_US|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED NOS |CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED (EVENT)
C0481253|T037|216993005|SNOMEDCT_US|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED (EVENT)
C0481253|T037|216993005|SNOMEDCT_US|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED NOS|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED (EVENT)
C0481253|T037|216993005|SNOMEDCT_US|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED |CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED (EVENT)
C0481253|T037|216993005|SNOMEDCT_US|CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED NOS |CONTAMINATED SUBSTANCE TRANSFUSED OR INFUSED (EVENT)
C1261338|T037|223196007|SNOMEDCT_US|CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCE, TRANSFUSED OR INFUSED|[X]CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCES, TRANSFUSED OR INFUSED (DISORDER)
C1261338|T037|223196007|SNOMEDCT_US|INJURY DUE TO CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCE, TRANSFUSED OR INFUSED|[X]CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCES, TRANSFUSED OR INFUSED (DISORDER)
C1261338|T037|223196007|SNOMEDCT_US|CONTAMINATED MED/BIOLOG SUB, TRANSFUSED OR INFUSED|[X]CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCES, TRANSFUSED OR INFUSED (DISORDER)
C1261338|T037|223196007|SNOMEDCT_US|[X]CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCES, TRANSFUSED OR INFUSED |[X]CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCES, TRANSFUSED OR INFUSED (DISORDER)
C1261338|T037|223196007|SNOMEDCT_US|[X]CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCES, TRANSFUSED OR INFUSED|[X]CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCES, TRANSFUSED OR INFUSED (DISORDER)
C1261338|T037|223196007|SNOMEDCT_US|[X]CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCES, TRANSFUSED OR INFUSED |[X]CONTAMINATED MEDICAL OR BIOLOGICAL SUBSTANCES, TRANSFUSED OR INFUSED (DISORDER)
C2108022|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH BACTERIA 
C2108022|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH BACTERIA
C2108032|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH ENDOTOXIN-PRODUCING BACTERIA 
C2108032|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH ENDOTOXIN-PRODUCING BACTERIA
C2108026|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH VIRUS 
C2108026|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH VIRUS
C2108013|T037||SNOMEDCT_US|CONTAMINATED BLOOD, FLUID, OR DRUG DURING TRANSFUSION OR INFUSION 
C2108013|T037||SNOMEDCT_US|CONTAMINATED BLOOD, FLUID, OR DRUG DURING TRANSFUSION OR INFUSION
C2108023|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH BACTERIAL PYOGENS 
C2108023|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH BACTERIAL PYOGENS
C2108024|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH HEPATOTOXIC SUBSTANCE
C2108024|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH HEPATOTOXIC SUBSTANCE 
C2108025|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH VIRAL HEPATITIS 
C2108025|T037||SNOMEDCT_US|CONTAMINATION DURING TRANSFUSION OR INFUSION WITH VIRAL HEPATITIS
C0030275|T037|149522005|SNOMEDCT_US|GRAFTINGS, PANCREAS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREAS GRAFTING|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREAS GRAFTINGS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREAS TRANSPLANTATION|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREAS TRANSPLANTATIONS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|TRANSPLANTATIONS, PANCREAS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREAS TRANSPL|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|TRANSPL PANCREAS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREATIC TRANSPLANTATION|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREATIC TRANSPLANTATION |PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREAT TRANSPLANT NOS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREAS TRANSPLANT|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|TRANSPLANTATION OF PANCREAS NOS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|TRANSPLANTATION OF PANCREAS NOS |PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREATIC TRANSPLANT|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREATIC TRANSPLANT |PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREAS TRANSPLANTATION PROCEDURES|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|GRAFTING, PANCREAS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|TRANSPLANTATION, PANCREAS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|TRANSPLANTATION OF PANCREAS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|TRANSPLANTATION OF PANCREAS |PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|TRANSPLANTATION OF PANCREAS, NOS|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|PANCREATIC TRANSPLANT, NOT OTHERWISE SPECIFIED|PANCREATIC TRANSPLANT (PROCEDURE)
C0030275|T037|149522005|SNOMEDCT_US|TRANSPLANT OF PANCREAS|PANCREATIC TRANSPLANT (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|GRAFTINGS, LUNG|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG GRAFTING|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG GRAFTINGS|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG TRANSPLANTATION|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG TRANSPLANTATIONS|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|TRANSPLANTATIONS, LUNG|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG TRANSPLANT|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG TRANSPL|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|TRANSPL LUNG|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG TRANSPLANT |TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|SURGERY LUNG TRANSPLANT|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG TRANSPLANT NOS|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|TRANSPLANT OF LUNG|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|TRANSPLANTATION OF LUNG NOS|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|TRANSPLANTATION OF LUNG NOS |TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG TRANSPLANT |TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG TRANSPLANTATION PROCEDURES|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNGS--TRANSPLANTATION|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|CARDIO/PULM: LUNG TRANSPLANT|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|GRAFTING, LUNG|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|TRANSPLANTATION, LUNG|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LTX - LUNG TRANSPLANT|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|TRANSPLANT OF LUNG |TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|TRANSPLANT OF LUNG, NOS|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|LUNG TRANSPLANTATION, NOT OTHERWISE SPECIFIED|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|EN BLOC LUNG TRANSPLANTATION|TRANSPLANT OF LUNG (PROCEDURE)
C0024128|T037|88039007|SNOMEDCT_US|TRANSPLANT;LUNG|TRANSPLANT OF LUNG (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|GRAFTING, HEART LUNG|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|GRAFTINGS, HEART-LUNG|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART LUNG TRANSPLANTATION|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART-LUNG GRAFTING|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART-LUNG GRAFTINGS|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART-LUNG TRANSPLANTATION|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART-LUNG TRANSPLANTATIONS|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|TRANSPLANTATION, HEART LUNG|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|TRANSPLANTATIONS, HEART-LUNG|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART AND LUNG TRANSPLANT|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|TRANSPL HEART LUNG|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART LUNG TRANSPL|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART-LUNG TRANSPLANT|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART-LUNG TRANSPLANT |HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART & LUNG TRANSPLANT|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|COMB HEART/LUNG TRANSPLA|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART AND HEART-LUNG TRANSPLANT|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART AND HEART-LUNG TRANSPLANT |HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|TRANSPLANTATION OF HEART AND LUNG NOS |HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|TRANSPLANTATION OF HEART AND LUNG NOS|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART AND HEART-LUNG TRANSPLANTATION|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART/LUNG TRANSPLANTATION PROCEDURES|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|GRAFTING, HEART-LUNG|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|TRANSPLANTATION, HEART-LUNG|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HLTX - HEART LUNG TRANSPLANT|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART LUNG GRAFTING|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|HEART AND LUNG TRANSPLANTATION|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0018833|T037|232971009|SNOMEDCT_US|COMBINED HEART-LUNG TRANSPLANTATION|HEART AND HEART-LUNG TRANSPLANT (PROCEDURE)
C0730400|T037|313039003|SNOMEDCT_US|SOLID ORGAN TRANSPLANT |SOLID ORGAN TRANSPLANT (PROCEDURE)
C0730400|T037|313039003|SNOMEDCT_US|SOLID ORGAN TRANSPLANT|SOLID ORGAN TRANSPLANT (PROCEDURE)
C0730400|T037|313039003|SNOMEDCT_US|SOLID ORGAN TRANSPLANT |SOLID ORGAN TRANSPLANT (PROCEDURE)
C0401176|T037|175902000|SNOMEDCT_US|RENAL TRANSPLANT CADAVERIC DONOR|CADAVERIC RENAL TRANSPLANT (PROCEDURE)
C0401176|T037|175902000|SNOMEDCT_US|CADAVERIC DONOR RENAL TRANSPLANT |CADAVERIC RENAL TRANSPLANT (PROCEDURE)
C0401176|T037|175902000|SNOMEDCT_US|CADAVERIC DONOR RENAL TRANSPLANT|CADAVERIC RENAL TRANSPLANT (PROCEDURE)
C0401176|T037|175902000|SNOMEDCT_US|CADAVER RENAL ALLOGRAFT|CADAVERIC RENAL TRANSPLANT (PROCEDURE)
C0401176|T037|175902000|SNOMEDCT_US|CADAVER RENAL ALLOTRANSPLANT|CADAVERIC RENAL TRANSPLANT (PROCEDURE)
C0401176|T037|175902000|SNOMEDCT_US|CADAVERIC RENAL TRANSPLANT|CADAVERIC RENAL TRANSPLANT (PROCEDURE)
C0401176|T037|175902000|SNOMEDCT_US|CADAVERIC RENAL TRANSPLANT |CADAVERIC RENAL TRANSPLANT (PROCEDURE)
C0194034|T037|149298002|SNOMEDCT_US|SPLEEN TRANSPLANTATION|SPLEEN TRANSPLANT (PROCEDURE)
C0194034|T037|149298002|SNOMEDCT_US|SPLEEN TRANSPLANT|SPLEEN TRANSPLANT (PROCEDURE)
C0194034|T037|149298002|SNOMEDCT_US|SPLEEN TRANSPLANT |SPLEEN TRANSPLANT (PROCEDURE)
C0194034|T037|149298002|SNOMEDCT_US|TRANSPLANTATION OF SPLEEN|SPLEEN TRANSPLANT (PROCEDURE)
C0194034|T037|149298002|SNOMEDCT_US|TRANSPLANTATION OF SPLEEN |SPLEEN TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|KIDNEY GRAFTING|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|KIDNEY TRANSPLANTATION|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|KIDNEY TRANSPLANTATIONS|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|RENAL TRANSPLANTATIONS|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANTATIONS, KIDNEY|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANTATIONS, RENAL|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|KIDNEY TRANSPLANT|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|RENAL TRANSPLANT|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|KIDNEY TRANSPL|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|RENAL TRANSPL|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPL RENAL|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPL KIDNEY|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|RENAL TRANSPLANTATION|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|RENAL TRANSPLANT |RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANTATION OF KIDNEY NOS |RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANTATION OF KIDNEY NOS|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|RENAL TRANSPLANT |RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|RENAL TRANSPLANTATION PROCEDURES|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|KIDNEYS--TRANSPLANTATION|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANTATION, KIDNEY|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANTATION, RENAL|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|GRAFTING, KIDNEY|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANT OF KIDNEY|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|RENAL GRAFT|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANTATION OF KIDNEY|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TX - KIDNEY TRANSPLANTATION|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TX - RENAL TRANSPLANTATION|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANT OF KIDNEY |RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANT OF KIDNEY, NOS|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|KIDNEY TRANSPLANTATION, NOS|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|RENAL TRANSPLANT, NOS|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|KIDNEY TRANSPLANTS|RENAL TRANSPLANT (PROCEDURE)
C0022671|T037|149586006|SNOMEDCT_US|TRANSPLANT;RENAL|RENAL TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|GRAFTINGS, LIVER|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|HEPATIC TRANSPLANTATIONS|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER GRAFTING|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER GRAFTINGS|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER TRANSPLANTATION|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER TRANSPLANTATIONS|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANTATIONS, HEPATIC|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANTATIONS, LIVER|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER TRANSPLANT|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|HEPATIC TRANSPLANTATION|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANTATION OF LIVER|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPL HEPATIC|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|HEPATIC TRANSPL|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPL LIVER|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER TRANSPL|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER TRANSPLANT |LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANTATION OF LIVER NOS|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANTATION OF LIVER NOS |LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER TRANSPLANT |LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER TRANSPLANTATION PROCEDURES|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LIVER--TRANSPLANTATION|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|GRAFTING, LIVER|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANTATION, LIVER|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANTATION, HEPATIC|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TX - LIVER TRANSPLANTATION|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|LTX - LIVER TRANSPLANT|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANTATION OF LIVER |LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANTATION OF LIVER, NOS|LIVER TRANSPLANT (PROCEDURE)
C0023911|T037|149473000|SNOMEDCT_US|TRANSPLANT;LIVER|LIVER TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|CARDIAC TRANSPLANTATIONS|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|GRAFTINGS, HEART|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HEART GRAFTING|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HEART GRAFTINGS|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HEART TRANSPLANTATION|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HEART TRANSPLANTATIONS|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPLANTATIONS, CARDIAC|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPLANTATIONS, HEART|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HEART TRANSPLANT|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPL CARDIAC|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|CARDIAC TRANSPL|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPL HEART|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HEART TRANSPL|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPLANTATION OF HEART|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPLANTATION OF HEART |HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|CARDIAC TRANSPLANTATION|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPLANT;CARDIAC|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HEART TRANSPLANT |HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HEART--TRANSPLANTATION|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|CARDIAC TRANSPLANT|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|CARDIO/PULM: HEART TRANSPLANT|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|GRAFTING, HEART|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPLANTATION, HEART|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPLANTATION, CARDIAC|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|CTX - CARDIAC TRANSPLANT|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HTX - HEART TRANSPLANT|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HTTX - HEART TRANSPLANT|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPLANTATION OF HEART |HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|TRANSPLANTATION OF HEART, NOS|HEART TRANSPLANT (PROCEDURE)
C0018823|T037|149204008|SNOMEDCT_US|HEART TRANSPLANTS|HEART TRANSPLANT (PROCEDURE)
C0857825|T037||SNOMEDCT_US|INFECTION IN SOLID ORGAN TRANSPLANT RECIPIENTS
