C0027415|T053||SNOMEDCT_US|NARCOTICS
C0202273|T053|40823001|SNOMEDCT_US|DRUG OF ABUSE, QUANTITATIVE SCREEN, INCLUDES AMPHETAMINES, BARBITURATES, BENZODIAZEPINES, CANNABINOIDS, COCAINE, METHADONE, METHAQUALONE, OPIATES, PHENCYCLIDINES AND PROPOXYPHENE|DRUG OF ABUSE, QUANTITATIVE SCREEN, INCLUDES AMPHETAMINES, BARBITURATES, BENZODIAZEPINES, CANNABINOIDS, COCAINE, METHADONE, METHAQUALONE, OPIATES, PHENCYCLIDINES AND PROPOXYPHENE (PROCEDURE)
C0086190|T053|77657003|SNOMEDCT_US|ILLICIT DRUGS|ILLEGAL DRUG (SUBSTANCE)
C2911101|T053||SNOMEDCT_US|DRUG ABUSE COUNSELING AND SURVEILLANCE OF DRUG ABUSER
C0202273|T053|40823001|SNOMEDCT_US|DRUG OF ABUSE, QUANTITATIVE SCREEN, INCLUDES AMPHETAMINES, BARBITURATES, BENZODIAZEPINES, CANNABINOIDS, COCAINE, METHADONE, METHAQUALONE, OPIATES, PHENCYCLIDINES AND PROPOXYPHENE|DRUG OF ABUSE, QUANTITATIVE SCREEN, INCLUDES AMPHETAMINES, BARBITURATES, BENZODIAZEPINES, CANNABINOIDS, COCAINE, METHADONE, METHAQUALONE, OPIATES, PHENCYCLIDINES AND PROPOXYPHENE (PROCEDURE)
C0221793|T053|395994000|SNOMEDCT_US|OPIATE ALKALOID|OPIUM ALKALOID (SUBSTANCE)
C0221793|T053|395994000|SNOMEDCT_US|ALKALOIDS, OPIATE|OPIUM ALKALOID (SUBSTANCE)
C0221793|T053|395994000|SNOMEDCT_US|OPIATE ALKALOIDS|OPIUM ALKALOID (SUBSTANCE)
C0221793|T053|395994000|SNOMEDCT_US|OPIATE ALKALOIDS [CHEMICAL/INGREDIENT]|OPIUM ALKALOID (SUBSTANCE)
C0221793|T053|395994000|SNOMEDCT_US|OPIUM ALKALOID|OPIUM ALKALOID (SUBSTANCE)
C0221793|T053|395994000|SNOMEDCT_US|OPIUM ALKALOID |OPIUM ALKALOID (SUBSTANCE)
C0221793|T053|395994000|SNOMEDCT_US|OPIUM ALKALOID |OPIUM ALKALOID (SUBSTANCE)
C0221793|T053|395994000|SNOMEDCT_US|OPIUM ALKALOIDS|OPIUM ALKALOID (SUBSTANCE)
C0025605|T053|387286002|SNOMEDCT_US|METHADONE|METHADONE (SUBSTANCE)
C0025605|T053|387286002|SNOMEDCT_US|3-HEPTANONE, 6-(DIMETHYLAMINO)-4,4-DIPHENYL-|METHADONE (SUBSTANCE)
C0025605|T053|387286002|SNOMEDCT_US|METHADONE [CHEMICAL/INGREDIENT]|METHADONE (SUBSTANCE)
C0025605|T053|387286002|SNOMEDCT_US|METHADONE |METHADONE (SUBSTANCE)
C0025605|T053|387286002|SNOMEDCT_US|METHADONE |METHADONE (SUBSTANCE)
C0030350|T053|372784001|SNOMEDCT_US|PAPAVERINE|PAPAVERINE (SUBSTANCE)
C0030350|T053|372784001|SNOMEDCT_US|ISOQUINOLINE, 1-((3,4-DIMETHOXYPHENYL)METHYL)-6,7-DIMETHOXY-|PAPAVERINE (SUBSTANCE)
C0030350|T053|372784001|SNOMEDCT_US|PAPAVERINE [CHEMICAL/INGREDIENT]|PAPAVERINE (SUBSTANCE)
C0030350|T053|372784001|SNOMEDCT_US|PAPAVERINE |PAPAVERINE (SUBSTANCE)
C0030350|T053|372784001|SNOMEDCT_US|PAPAVERINE |PAPAVERINE (SUBSTANCE)
C0030350|T053|372784001|SNOMEDCT_US|PAP|PAPAVERINE (SUBSTANCE)
C0728935|T053||SNOMEDCT_US|K 315
C0728935|T053||SNOMEDCT_US|K315
C0728935|T053||SNOMEDCT_US|K-315
C0205752|T053||SNOMEDCT_US|ENDOGENOUS OPIOIDS
C0205752|T053||SNOMEDCT_US|ENDOGENOUS OPIATE
C0205752|T053||SNOMEDCT_US|ENDOGENOUS OPIATES
C0205752|T053||SNOMEDCT_US|ENDORPHIN
C0205752|T053||SNOMEDCT_US|ENDOGENOUS OPIOID
C0205752|T053||SNOMEDCT_US|OPIOIDS (ENDOGENOUS)
C0205752|T053||SNOMEDCT_US|OPIATES, ENDOGENOUS
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHANOL TARTRATE|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|TARTRATE, LEVORPHANOL|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|L-3-HYDROXY-N-METHYLMORPHINAN BITARTRATE|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|2H-10,4A-IMINOETHANOPHENANTHREN-6-OL, 1,3,4,9,10,10A-HEXAHYDRO-11-METHYL-, TARTRATE|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEMORAN|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|MORPHINAN-3-OL, 17-METHYL-, TARTRATE(1:1)(SALT)|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|MORPHINAN-3-OL, 17-METHYL-,(2R,3R)-2,3-DIHYDROXYBUTANEDIOATE(1:1)|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|NIH 4590|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|RO 1-5431/7|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHANOL TARTRATE |LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|SYNTHETIC NARCOTICS LEVORPHANOL TARTRATE|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHANOL TARTRATE [CHEMICAL/INGREDIENT]|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHANOL TARTRATE [ANAESTH]|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHANOL TARTRATE [ANESTH]|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHANOL TARTRATE |LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHANOL TARTRATE [ANESTH] |LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHAN TARTRATE|LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHANOL TARTRATE [ANESTH] |LEVORPHANOL TARTRATE (SUBSTANCE)
C0596008|T053|67347006|SNOMEDCT_US|LEVORPHANOL TARTRATE [DUP] |LEVORPHANOL TARTRATE (SUBSTANCE)
C0376196|T053|360204007|SNOMEDCT_US|OPIATES|OPIATE (PRODUCT)
C0376196|T053|360204007|SNOMEDCT_US|OPIATE|OPIATE (PRODUCT)
C0376196|T053|360204007|SNOMEDCT_US|OPIATE |OPIATE (PRODUCT)
C0376196|T053|360204007|SNOMEDCT_US|OPIUM DERIVATIVES|OPIATE (PRODUCT)
C0002327|T053|52885008|SNOMEDCT_US|ALPHAPRODINE|ALPHAPRODINE (SUBSTANCE)
C0002327|T053|52885008|SNOMEDCT_US|4-PIPERIDINOL, 1,3-DIMETHYL-4-PHENYL-, PROPANOATE (ESTER), CIS-|ALPHAPRODINE (SUBSTANCE)
C0002327|T053|52885008|SNOMEDCT_US|ALPHAPRODINE [CHEMICAL/INGREDIENT]|ALPHAPRODINE (SUBSTANCE)
C0002327|T053|52885008|SNOMEDCT_US|ALPHAPRODINE |ALPHAPRODINE (SUBSTANCE)
C0006405|T053|387173000|SNOMEDCT_US|BUPRENORPHINE|BUPRENORPHINE (SUBSTANCE)
C0006405|T053|387173000|SNOMEDCT_US|6,14-ETHENOMORPHINAN-7-METHANOL, 17-(CYCLOPROPYLMETHYL)-ALPHA-(1,1-DIMETHYLETHYL)-4,5-EPOXY-18,19-DIHYDRO-3-HYDROXY-6-METHOXY-ALPHA-METHYL-, (5ALPHA,7ALPHA(S))-|BUPRENORPHINE (SUBSTANCE)
C0006405|T053|387173000|SNOMEDCT_US|BUPRENORPHINE [CHEMICAL/INGREDIENT]|BUPRENORPHINE (SUBSTANCE)
C0006405|T053|387173000|SNOMEDCT_US|BUPRENORPHINE PRODUCT|BUPRENORPHINE (SUBSTANCE)
C0006405|T053|387173000|SNOMEDCT_US|BUPRENORPHINE PRODUCT |BUPRENORPHINE (SUBSTANCE)
C0006405|T053|387173000|SNOMEDCT_US|BUPRENORPHINE |BUPRENORPHINE (SUBSTANCE)
C0006405|T053|387173000|SNOMEDCT_US|BUPRENORPHINE |BUPRENORPHINE (SUBSTANCE)
C0006491|T053|373467000|SNOMEDCT_US|BUTORPHANOL|BUTORPHANOL (SUBSTANCE)
C0006491|T053|373467000|SNOMEDCT_US|MORPHINAN-3,14-DIOL, 17-(CYCLOBUTYLMETHYL)-|BUTORPHANOL (SUBSTANCE)
C0006491|T053|373467000|SNOMEDCT_US|17-(CYCLOBUTYLMETHYL)MORPHINAN-3,14-DIOL|BUTORPHANOL (SUBSTANCE)
C0006491|T053|373467000|SNOMEDCT_US|BUTORPHANOL [CHEMICAL/INGREDIENT]|BUTORPHANOL (SUBSTANCE)
C0006491|T053|373467000|SNOMEDCT_US|BUTORPHANOL PRODUCT|BUTORPHANOL (SUBSTANCE)
C0006491|T053|373467000|SNOMEDCT_US|BUTORPHANOL PRODUCT |BUTORPHANOL (SUBSTANCE)
C0006491|T053|373467000|SNOMEDCT_US|BUTORPHANOL |BUTORPHANOL (SUBSTANCE)
C0006491|T053|373467000|SNOMEDCT_US|BUTORPHANOL |BUTORPHANOL (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|CODEINE|CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|N METHYLMORPHINE|CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|MORPHINAN-6-OL, 7,8-DIDEHYDRO-4,5-EPOXY-3-METHOXY-17-METHYL-, (5ALPHA,6ALPHA)-|CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|CODEINE |CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|NARCOTICS CODEINE|CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|CODEINE [CHEMICAL/INGREDIENT]|CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|N-METHYLMORPHINE|CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|METHYL MORPHINE|CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|METHYLMORPHINE|CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|CODEINE |CODEINE (SUBSTANCE)
C0009214|T053|387494007|SNOMEDCT_US|CODEINE |CODEINE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|D MORAMIDE|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|DEXTROMORAMIDE|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|PYRROLIDINE, 1-(3-METHYL-4-(4-MORPHOLINYL)-1-OXO-2,2-DIPHENYLBUTYL)-, (S)-|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|MORAMIDE D|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|PYRROLAMIDOL|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|D-MORAMIDE|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|DEXTROMORAMIDE [CHEMICAL/INGREDIENT]|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|SKF-5137|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|4-(2-METHYL-4-OXO-3,3-DIPHENYL-4-(1-PYRROLIDINYL)BUTYL)MORPHOLINE|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|R-875|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|(+)-4-(2-METHYL-4-OXO-3,3-DIPHENYL-4-(1-PYRROLIDINYL)BUTYL)MORPHOLINE|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|D-2,2-DIPHENYL-3-METHYL-4-MORPHOLINOBUTYRYLPYRROLIDINE|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|(+)-1-(3-METHYL-4-MORPHOLINO-2,2-DIPHENYLBUTYRYL)PYRROLIDINE|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|1-((3S)-3-METHYL-4-(4-MORPHOLINYL)-1-OXO-2,2-DIPHENYLBUTYL)PYRROLIDINE|DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|DEXTROMORAMIDE |DEXTROMORAMIDE (SUBSTANCE)
C0011817|T053|387561007|SNOMEDCT_US|DEXTROMORAMIDE |DEXTROMORAMIDE (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|HEROIN|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|MORPHINAN-3,6-DIOL, 7,8-DIDEHYDRO-4,5-EPOXY-17-METHYL- (5ALPHA,6ALPHA)-, DIACETATE (ESTER)|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|DIACETYLMORPHINE|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|DIAMORPHINE|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|HEROIN [CHEMICAL/INGREDIENT]|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|HEROIN (SCHEDULE I SUBSTANCE)|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|JUNK|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|SMACK|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|SKAG|HEROIN (SUBSTANCE)
# C0011892|T053|387341002|SNOMEDCT_US|H|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|ACETOMORPHINE|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|BLACK TAR|HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|HEROIN |HEROIN (SUBSTANCE)
C0011892|T053|387341002|SNOMEDCT_US|HEROIN |HEROIN (SUBSTANCE)
C0012305|T053||SNOMEDCT_US|DIHYDROMORPHINE
C0012305|T053||SNOMEDCT_US|MORPHINAN-3,6-DIOL, 4,5-EPOXY-17-METHYL-, (5ALPHA,6ALPHA)-
C0012305|T053||SNOMEDCT_US|DIHYDROMORPHINE [CHEMICAL/INGREDIENT]
C0012305|T053||SNOMEDCT_US|PARAMORPHAN
C0012305|T053||SNOMEDCT_US|PARAMORFAN
C0012306|T053|414428000|SNOMEDCT_US|HYDROMORPHONE|HYDROMORPHONE (PRODUCT)
C0012306|T053|414428000|SNOMEDCT_US|MORPHINAN-6-ONE, 4,5-EPOXY-3-HYDROXY-17-METHYL-, (5ALPHA)-|HYDROMORPHONE (PRODUCT)
C0012306|T053|414428000|SNOMEDCT_US|DIHYDROMORPHINONE|HYDROMORPHONE (PRODUCT)
C0012306|T053|414428000|SNOMEDCT_US|HYDROMORPHON|HYDROMORPHONE (PRODUCT)
C0012306|T053|414428000|SNOMEDCT_US|HYDROMORPHONE |HYDROMORPHONE (PRODUCT)
C0012306|T053|414428000|SNOMEDCT_US|HYDROMORPHONE [CHEMICAL/INGREDIENT]|HYDROMORPHONE (PRODUCT)
C0012306|T053|414428000|SNOMEDCT_US|(-)-HYDROMORPHONE|HYDROMORPHONE (PRODUCT)
C0012306|T053|414428000|SNOMEDCT_US|HYDROMORPHONE |HYDROMORPHONE (PRODUCT)
C0012306|T053|414428000|SNOMEDCT_US|HYDROMORPHONE |HYDROMORPHONE (PRODUCT)
C0015109|T053|422453004|SNOMEDCT_US|ETHYLMORPHINE|ETHYLMORPHINE (PRODUCT)
C0015109|T053|422453004|SNOMEDCT_US|MORPHINAN-6-OL, 7,8-DIDEHYDRO-4,5-EPOXY-3-ETHOXY-17-METHYL-, (5ALPHA,6ALPHA)-|ETHYLMORPHINE (PRODUCT)
C0015109|T053|422453004|SNOMEDCT_US|ETHYLMORPHINE |ETHYLMORPHINE (PRODUCT)
C0015109|T053|422453004|SNOMEDCT_US|CODETHYLINE|ETHYLMORPHINE (PRODUCT)
C0015109|T053|422453004|SNOMEDCT_US|ETHOMORPHINE|ETHYLMORPHINE (PRODUCT)
C0015109|T053|422453004|SNOMEDCT_US|ETHYLMORPHINE [CHEMICAL/INGREDIENT]|ETHYLMORPHINE (PRODUCT)
C0015109|T053|422453004|SNOMEDCT_US|(5ALPHA,6ALPHA)-7,8-DIDEHYDRO-4,5-EPOXY-3-ETHOXY-17-METHYLMORPHINAN-6-OL|ETHYLMORPHINE (PRODUCT)
C0015109|T053|422453004|SNOMEDCT_US|ETHYL MORPHINE|ETHYLMORPHINE (PRODUCT)
C0015109|T053|422453004|SNOMEDCT_US|ETHYL MORPHINE |ETHYLMORPHINE (PRODUCT)
C0015134|T053|96188003|SNOMEDCT_US|ETORPHINE|ETORPHINE (SUBSTANCE)
C0015134|T053|96188003|SNOMEDCT_US|6,14-ETHENOMORPHINAN-7-METHANOL, 4,5-EPOXY-3-HYDROXY-6-METHOXY-ALPHA,17-DIMETHYL-ALPHA-PROPYL-, (5ALPHA,7ALPHA(R))-|ETORPHINE (SUBSTANCE)
C0015134|T053|96188003|SNOMEDCT_US|ETHORPHINE|ETORPHINE (SUBSTANCE)
C0015134|T053|96188003|SNOMEDCT_US|ETORPHINE [CHEMICAL/INGREDIENT]|ETORPHINE (SUBSTANCE)
C0015134|T053|96188003|SNOMEDCT_US|ETORPHINE |ETORPHINE (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|FENTANYL|FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|PROPANAMIDE, N-PHENYL-N-(1-(2-PHENYLETHYL)-4-PIPERIDINYL)-|FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|FENTYL|FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|FENTANYL |FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|FENTANYL [CHEMICAL/INGREDIENT]|FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|PHENTANYL|FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|N-(1-PHENETHYLPIPERIDIN-4-YL)-N-PHENYLPROPIONAMIDE|FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|LOCAL ANESTHETIC FENTANYL |FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|LOCAL ANESTHETIC FENTANYL|FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|FENTANYL PRODUCT|FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|FENTANYL |FENTANYL (SUBSTANCE)
C0015846|T053|373492002|SNOMEDCT_US|FENTANYL |FENTANYL (SUBSTANCE)
C0020264|T053|372671002|SNOMEDCT_US|HYDROCODONE|HYDROCODONE (SUBSTANCE)
C0020264|T053|372671002|SNOMEDCT_US|MORPHINAN-6-ONE, 4,5-EPOXY-3-METHOXY-17-METHYL-, (5ALPHA)-|HYDROCODONE (SUBSTANCE)
C0020264|T053|372671002|SNOMEDCT_US|HYDROCODONE [CHEMICAL/INGREDIENT]|HYDROCODONE (SUBSTANCE)
C0020264|T053|372671002|SNOMEDCT_US|DIHYDROCODEINONE|HYDROCODONE (SUBSTANCE)
C0020264|T053|372671002|SNOMEDCT_US|HYDROCODON|HYDROCODONE (SUBSTANCE)
C0020264|T053|372671002|SNOMEDCT_US|HYDROCODONE |HYDROCODONE (SUBSTANCE)
C0020264|T053|372671002|SNOMEDCT_US|HYDROCODONE |HYDROCODONE (SUBSTANCE)
C0023586|T053|387275004|SNOMEDCT_US|LEVORPHANOL|LEVORPHANOL (SUBSTANCE)
C0023586|T053|387275004|SNOMEDCT_US|MORPHINAN-3-OL, 17-METHYL-|LEVORPHANOL (SUBSTANCE)
C0023586|T053|387275004|SNOMEDCT_US|LEVORPHANOL [CHEMICAL/INGREDIENT]|LEVORPHANOL (SUBSTANCE)
C0023586|T053|387275004|SNOMEDCT_US|LEVODROMAN|LEVORPHANOL (SUBSTANCE)
C0023586|T053|387275004|SNOMEDCT_US|LEVORPHAN|LEVORPHANOL (SUBSTANCE)
C0023586|T053|387275004|SNOMEDCT_US|LEVORPHANOL |LEVORPHANOL (SUBSTANCE)
C0023586|T053|387275004|SNOMEDCT_US|LEVORPHANOL |LEVORPHANOL (SUBSTANCE)
C0025376|T053|54544005|SNOMEDCT_US|MEPERIDINE|MEPERIDINE (SUBSTANCE)
C0025376|T053|54544005|SNOMEDCT_US|4-PIPERIDINECARBOXYLIC ACID, 1-METHYL-4-PHENYL-, ETHYL ESTER|MEPERIDINE (SUBSTANCE)
C0025376|T053|54544005|SNOMEDCT_US|ISONIPECAIN|MEPERIDINE (SUBSTANCE)
C0025376|T053|54544005|SNOMEDCT_US|MEPERIDINE [CHEMICAL/INGREDIENT]|MEPERIDINE (SUBSTANCE)
C0025376|T053|54544005|SNOMEDCT_US|PETHIDINE|MEPERIDINE (SUBSTANCE)
C0025376|T053|54544005|SNOMEDCT_US|NARCOTICS MEPERIDINE|MEPERIDINE (SUBSTANCE)
C0025376|T053|54544005|SNOMEDCT_US|MEPERIDINE |MEPERIDINE (SUBSTANCE)
C0025376|T053|54544005|SNOMEDCT_US|MEPERIDINE |MEPERIDINE (SUBSTANCE)
C0025376|T053|54544005|SNOMEDCT_US|MEPERIDINE |MEPERIDINE (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL|MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|PHENOL, 3-(3-ETHYLHEXAHYDRO-1-METHYL-1H-AZEPIN-3-YL)-|MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL [CHEMICAL/INGREDIENT]|MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|M-(3-ETHYLHEXAHYDRO-1-METHYL-1H-AZEPIN-3-YL)PHENOL|MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL [ANESTHESIA] |MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL [ANALGESIC] |MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL [ANAESTHESIA]|MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL [ANALGESIC]|MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL [ANESTHESIA]|MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL |MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL |MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL [ANALGESIC] |MEPTAZINOL (SUBSTANCE)
C0025387|T053|395783008|SNOMEDCT_US|MEPTAZINOL [ANESTHESIA] |MEPTAZINOL (SUBSTANCE)
C0025607|T053||SNOMEDCT_US|METHADYL ACETATE
C0025607|T053||SNOMEDCT_US|METHADYLACETATE
C0025607|T053||SNOMEDCT_US|BENZENEETHANOL, BETA-(2-(DIMETHYLAMINO)PROPYL)-ALPHA-ETHYL-BETA-PHENYL-, ACETATE (ESTER)
C0025607|T053||SNOMEDCT_US|ACETYLMETHADOL
C0025607|T053||SNOMEDCT_US|METHADYL ACETATE [CHEMICAL/INGREDIENT]
C0025607|T053||SNOMEDCT_US|6-(DIMETHYLAMINO)-4,4-DIPHENYL-3-HEPTANOL ACETATE
C0026549|T053|373529000|SNOMEDCT_US|MORPHINE|MORPHINE (SUBSTANCE)
C0026549|T053|373529000|SNOMEDCT_US|MORPHINAN-3,6-DIOL, 7,8-DIDEHYDRO-4,5-EPOXY-17-METHYL- (5ALPHA,6ALPHA)-|MORPHINE (SUBSTANCE)
C0026549|T053|373529000|SNOMEDCT_US|MORPHIA|MORPHINE (SUBSTANCE)
C0026549|T053|373529000|SNOMEDCT_US|MORPHINE [CHEMICAL/INGREDIENT]|MORPHINE (SUBSTANCE)
C0026549|T053|373529000|SNOMEDCT_US|NARCOTICS MORPHINE|MORPHINE (SUBSTANCE)
C0026549|T053|373529000|SNOMEDCT_US|MORPHINE |MORPHINE (SUBSTANCE)
C0026549|T053|373529000|SNOMEDCT_US|MORPHINE |MORPHINE (SUBSTANCE)
C0026549|T053|373529000|SNOMEDCT_US|MORPHINE |MORPHINE (SUBSTANCE)
C0026549|T053|373529000|SNOMEDCT_US|MORPH|MORPHINE (SUBSTANCE)
C0027348|T053|373539006|SNOMEDCT_US|NALBUPHINE|NALBUPHINE (SUBSTANCE)
C0027348|T053|373539006|SNOMEDCT_US|MORPHINAN-3,6,14-TRIOL, 17-(CYCLOBUTYLMETHYL)-4,5-EPOXY-, (5ALPHA,6ALPHA)-|NALBUPHINE (SUBSTANCE)
C0027348|T053|373539006|SNOMEDCT_US|NALBUPHINE [CHEMICAL/INGREDIENT]|NALBUPHINE (SUBSTANCE)
C0027348|T053|373539006|SNOMEDCT_US|NALBUPHINE PRODUCT |NALBUPHINE (SUBSTANCE)
C0027348|T053|373539006|SNOMEDCT_US|NALBUPHINE PRODUCT|NALBUPHINE (SUBSTANCE)
C0027348|T053|373539006|SNOMEDCT_US|NALBUPHINE |NALBUPHINE (SUBSTANCE)
C0027348|T053|373539006|SNOMEDCT_US|NALBUPHINE |NALBUPHINE (SUBSTANCE)
C0029112|T053|21919007|SNOMEDCT_US|OPIUM|OPIUM (SUBSTANCE)
C0029112|T053|21919007|SNOMEDCT_US|OPIUM PREPARATIONS |OPIUM (SUBSTANCE)
C0029112|T053|21919007|SNOMEDCT_US|OPIUM PREPARATIONS|OPIUM (SUBSTANCE)
C0029112|T053|21919007|SNOMEDCT_US|OPIUM [CHEMICAL/INGREDIENT]|OPIUM (SUBSTANCE)
C0029112|T053|21919007|SNOMEDCT_US|OPIUM PREPARATION|OPIUM (SUBSTANCE)
C0029112|T053|21919007|SNOMEDCT_US|OPIUM |OPIUM (SUBSTANCE)
C0029112|T053|21919007|SNOMEDCT_US|OPIUM PREPARATION |OPIUM (SUBSTANCE)
C0029112|T053|21919007|SNOMEDCT_US|OPIUM PREPARATION |OPIUM (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCODONE|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|MORPHINAN-6-ONE, 4,5-EPOXY-14-HYDROXY-3-METHOXY-17-METHYL-, (5ALPHA)-|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|4,5-EPOXY-14-HYDROXY-3-METHOXY-17-METHYLMORPHINAN-6-ONE|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCODONE |OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|SYNTHETIC NARCOTICS OXYCODONE|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|DIHYDROHYDROXYCODEINONE|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCODONE [CHEMICAL/INGREDIENT]|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCODEINON|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|DINARKON|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|DIHYDRONE|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCONE|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCODONE PRODUCT |OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCODONE PRODUCT|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|14-HYDROXYDIHYDROCODEINONE|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCODONE |OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCODONE SR|OXYCODONE (SUBSTANCE)
C0030049|T053|55452001|SNOMEDCT_US|OXYCODONE |OXYCODONE (SUBSTANCE)
C0030073|T053|24751001|SNOMEDCT_US|OXYMORPHONE|OXYMORPHONE (SUBSTANCE)
C0030073|T053|24751001|SNOMEDCT_US|MORPHINAN-6-ONE, 4,5-EPOXY-3,14-DIHYDROXY-17-METHYL-, (5ALPHA)-|OXYMORPHONE (SUBSTANCE)
C0030073|T053|24751001|SNOMEDCT_US|OXYMORPHONE [CHEMICAL/INGREDIENT]|OXYMORPHONE (SUBSTANCE)
C0030073|T053|24751001|SNOMEDCT_US|MORPHINAN-6-ONE, 4,5-EPOXY-3,14-DIHYDROXY-17-METHYL-|OXYMORPHONE (SUBSTANCE)
C0030073|T053|24751001|SNOMEDCT_US|4,5ALPHA-EPOXY-3,14-DIHYDROXY-17-METHYLMORPHINAN-6-ONE|OXYMORPHONE (SUBSTANCE)
C0030073|T053|24751001|SNOMEDCT_US|OXYMORPHONE |OXYMORPHONE (SUBSTANCE)
C0030073|T053|24751001|SNOMEDCT_US|OXYMORPHONE PRODUCT |OXYMORPHONE (SUBSTANCE)
C0030073|T053|24751001|SNOMEDCT_US|OXYMORPHONE PRODUCT|OXYMORPHONE (SUBSTANCE)
C0030873|T053|387213004|SNOMEDCT_US|PENTAZOCINE|PENTAZOCINE (SUBSTANCE)
C0030873|T053|387213004|SNOMEDCT_US|2,6-METHANO-3-BENZAZOCIN-8-OL, 1,2,3,4,5,6-HEXAHYDRO-6,11-DIMETHYL-3-(3-METHYL-2-BUTENYL)-, (2ALPHA,6ALPHA,11R*)-|PENTAZOCINE (SUBSTANCE)
C0030873|T053|387213004|SNOMEDCT_US|PENTAZOCINE |PENTAZOCINE (SUBSTANCE)
C0030873|T053|387213004|SNOMEDCT_US|SYNTHETIC NARCOTICS PENTAZOCINE|PENTAZOCINE (SUBSTANCE)
C0030873|T053|387213004|SNOMEDCT_US|PENTAZOCINE [CHEMICAL/INGREDIENT]|PENTAZOCINE (SUBSTANCE)
C0030873|T053|387213004|SNOMEDCT_US|PENTAZOCINE |PENTAZOCINE (SUBSTANCE)
C0030873|T053|387213004|SNOMEDCT_US|PENTAZOCINE |PENTAZOCINE (SUBSTANCE)
C0031376|T053|387326002|SNOMEDCT_US|PHENAZOCINE|PHENAZOCINE (SUBSTANCE)
C0031376|T053|387326002|SNOMEDCT_US|2,6-METHANO-3-BENZAZOCIN-8-OL, 1,2,3,4,5,6-HEXAHYDRO-6,11-DIMETHYL-3-(2-PHENYLETHYL)-|PHENAZOCINE (SUBSTANCE)
C0031376|T053|387326002|SNOMEDCT_US|PHENAZOCINE [CHEMICAL/INGREDIENT]|PHENAZOCINE (SUBSTANCE)
C0031376|T053|387326002|SNOMEDCT_US|PHENBENZORPHAN|PHENAZOCINE (SUBSTANCE)
C0031376|T053|387326002|SNOMEDCT_US|PHENETHYLAZOCINE|PHENAZOCINE (SUBSTANCE)
C0031376|T053|387326002|SNOMEDCT_US|PHENAZOCINE |PHENAZOCINE (SUBSTANCE)
C0031376|T053|387326002|SNOMEDCT_US|PHENAZOCINE |PHENAZOCINE (SUBSTANCE)
C0031432|T053|420076001|SNOMEDCT_US|PHENOPERIDINE|PHENOPERIDINE (SUBSTANCE)
C0031432|T053|420076001|SNOMEDCT_US|4-PIPERIDINECARBOXYLIC ACID, 1-(3-HYDROXY-3-PHENYLPROPYL)-4-PHENYL-, ETHYL ESTER|PHENOPERIDINE (SUBSTANCE)
C0031432|T053|420076001|SNOMEDCT_US|FENOPERIDINE|PHENOPERIDINE (SUBSTANCE)
C0031432|T053|420076001|SNOMEDCT_US|PHENOPERIDINE [CHEMICAL/INGREDIENT]|PHENOPERIDINE (SUBSTANCE)
C0031432|T053|420076001|SNOMEDCT_US|PHENOPERIDINE |PHENOPERIDINE (SUBSTANCE)
C0031432|T053|420076001|SNOMEDCT_US|PHENOPERIDINE |PHENOPERIDINE (SUBSTANCE)
C0031982|T053|707837002|SNOMEDCT_US|PIRINITRAMIDE|PIRITRAMIDE (SUBSTANCE)
C0031982|T053|707837002|SNOMEDCT_US|(1,4'-BIPIPERIDINE)-4'-CARBOXAMIDE, 1'-(3-CYANO-3,3-DIPHENYLPROPYL)-|PIRITRAMIDE (SUBSTANCE)
C0031982|T053|707837002|SNOMEDCT_US|PIRITRAMIDE|PIRITRAMIDE (SUBSTANCE)
C0031982|T053|707837002|SNOMEDCT_US|PIRINITRAMIDE [CHEMICAL/INGREDIENT]|PIRITRAMIDE (SUBSTANCE)
C0031982|T053|707837002|SNOMEDCT_US|PIRITRAMID|PIRITRAMIDE (SUBSTANCE)
C0031982|T053|707837002|SNOMEDCT_US|PIRITRAMIDE |PIRITRAMIDE (SUBSTANCE)
C0031982|T053|707837002|SNOMEDCT_US|1'-(3-CYANO-3,3-DIPHENYLPROPYL)-(1,4'-BIPIPERIDINE)-4'-CARBOXAMIDE|PIRITRAMIDE (SUBSTANCE)
C0031982|T053|707837002|SNOMEDCT_US|(1,4'-BIPIPERIDINE)-4'-CARBOXAMIDE, 1'-(3-CYANO-3,3-DIPHENYLPROPYL)|PIRITRAMIDE (SUBSTANCE)
C0031982|T053|707837002|SNOMEDCT_US|R 3365|PIRITRAMIDE (SUBSTANCE)
C0033400|T053||SNOMEDCT_US|PROMEDOL
C0033400|T053||SNOMEDCT_US|4-PIPERIDINOL, 1,2,5-TRIMETHYL-4-PHENYL-, PROPANOATE (ESTER)
C0033400|T053||SNOMEDCT_US|DIMETHYLMEPERIDINE
C0033400|T053||SNOMEDCT_US|PROMEDOL [CHEMICAL/INGREDIENT]
C0039746|T053|89851001|SNOMEDCT_US|THEBAINE|THEBAINE (SUBSTANCE)
C0039746|T053|89851001|SNOMEDCT_US|MORPHINAN, 6,7,8,14-TETRADEHYDRO-4,5-EPOXY-3,6-DIMETHOXY-17-METHYL-, (5ALPHA)-|THEBAINE (SUBSTANCE)
C0039746|T053|89851001|SNOMEDCT_US|THEBAINE [CHEMICAL/INGREDIENT]|THEBAINE (SUBSTANCE)
C0039746|T053|89851001|SNOMEDCT_US|3-O-METHYL-ORIPAVIN|THEBAINE (SUBSTANCE)
C0039746|T053|89851001|SNOMEDCT_US|4,5ALPHA-EPOXY-3,6-DIMETHOXY-17-METHYL-6,8-MORPHINADIEN|THEBAINE (SUBSTANCE)
C0039746|T053|89851001|SNOMEDCT_US|PARAMORPHINE|THEBAINE (SUBSTANCE)
C0039746|T053|89851001|SNOMEDCT_US|THEBAINE |THEBAINE (SUBSTANCE)
C0040219|T053|373562008|SNOMEDCT_US|TILIDINE|TILIDINE (SUBSTANCE)
C0040219|T053|373562008|SNOMEDCT_US|3-CYCLOHEXENE-1-CARBOXYLIC ACID, 2-(DIMETHYLAMINO)-1-PHENYL-, ETHYL ESTER, TRANS-(+-)-|TILIDINE (SUBSTANCE)
C0040219|T053|373562008|SNOMEDCT_US|TILIDATE|TILIDINE (SUBSTANCE)
C0040219|T053|373562008|SNOMEDCT_US|TILIDINE [CHEMICAL/INGREDIENT]|TILIDINE (SUBSTANCE)
C0040219|T053|373562008|SNOMEDCT_US|TILIDINE |TILIDINE (SUBSTANCE)
C0040219|T053|373562008|SNOMEDCT_US|TILIDINE |TILIDINE (SUBSTANCE)
C0040610|T053|386858008|SNOMEDCT_US|TRAMADOL|TRAMADOL (SUBSTANCE)
C0040610|T053|386858008|SNOMEDCT_US|CYCLOHEXANOL, 2-((DIMETHYLAMINO)METHYL)-1-(3-METHOXYPHENYL)-, CIS-(+-)-|TRAMADOL (SUBSTANCE)
C0040610|T053|386858008|SNOMEDCT_US|TRAMADOL [CHEMICAL/INGREDIENT]|TRAMADOL (SUBSTANCE)
C0040610|T053|386858008|SNOMEDCT_US|TRAMADOL |TRAMADOL (SUBSTANCE)
C0040610|T053|386858008|SNOMEDCT_US|TRAMADOL |TRAMADOL (SUBSTANCE)
C0002026|T053|387560008|SNOMEDCT_US|ALFENTANIL|ALFENTANIL (SUBSTANCE)
C0002026|T053|387560008|SNOMEDCT_US|PROPANAMIDE, N-(1-(2-(4-ETHYL-4,5-DIHYDRO-5-OXO-1H-TETRAZOL-1-YL)ETHYL)-4-(METHOXYMETHYL)-4-PIPERIDINYL)-N-PHENYL-|ALFENTANIL (SUBSTANCE)
C0002026|T053|387560008|SNOMEDCT_US|ALFENTANYL|ALFENTANIL (SUBSTANCE)
C0002026|T053|387560008|SNOMEDCT_US|ALFENTANIL [CHEMICAL/INGREDIENT]|ALFENTANIL (SUBSTANCE)
C0002026|T053|387560008|SNOMEDCT_US|ALFENTANIL - CHEMICAL|ALFENTANIL (SUBSTANCE)
C0002026|T053|387560008|SNOMEDCT_US|ALFENTANIL - CHEMICAL |ALFENTANIL (SUBSTANCE)
C0002026|T053|387560008|SNOMEDCT_US|ALFENTANIL |ALFENTANIL (SUBSTANCE)
C0002026|T053|387560008|SNOMEDCT_US|ALFENTANIL |ALFENTANIL (SUBSTANCE)
C0143993|T053|49998007|SNOMEDCT_US|SUFENTANIL|SUFENTANIL (SUBSTANCE)
C0143993|T053|49998007|SNOMEDCT_US|PROPANAMIDE, N-(4-(METHOXYMETHYL)-1-(2-(2-THIENYL)ETHYL)-4-PIPERIDINYL)-N-PHENYL-|SUFENTANIL (SUBSTANCE)
C0143993|T053|49998007|SNOMEDCT_US|SUFENTANIL [CHEMICAL/INGREDIENT]|SUFENTANIL (SUBSTANCE)
C0143993|T053|49998007|SNOMEDCT_US|SULFENTANYL|SUFENTANIL (SUBSTANCE)
C0143993|T053|49998007|SNOMEDCT_US|SULFENTANIL|SUFENTANIL (SUBSTANCE)
C0143993|T053|49998007|SNOMEDCT_US|SUFENTANIL |SUFENTANIL (SUBSTANCE)
C0143993|T053|49998007|SNOMEDCT_US|SUFENTANIL PRODUCT |SUFENTANIL (SUBSTANCE)
C0143993|T053|49998007|SNOMEDCT_US|SUFENTANIL PRODUCT|SUFENTANIL (SUBSTANCE)
C0033493|T053|117005003|SNOMEDCT_US|PROPOXYPHENE|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|D PROPOXYPHENE|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|BENZENEETHANOL, ALPHA-(2-(DIMETHYLAMINO)-1-METHYLETHYL)-ALPHA-PHENYL-, PROPANOATE (ESTER), (S-(R*,S*))-|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|PROPOXYPHENE D|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|DEXTROPROPOXYPHENE|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|PROPOXYPHENE |PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|DEXTROPROPOXYPHENE |PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|SYNTHETIC NARCOTICS PROPOXYPHENE PREPARATIONS|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|PROPOXYPHENE PREPARATIONS |PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|PROPOXYPHENE PREPARATIONS|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|D-PROPOXYPHENE|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|DEXTROPROPOXYPHENE [CHEMICAL/INGREDIENT]|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|4-DIMETHYLAMINO-3-METHYL-1,2-DIPHENYL-2-PROPOXYBUTANE|PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|PROPOXYPHENE |PROPOXYPHENE (PRODUCT)
C0033493|T053|117005003|SNOMEDCT_US|DEXTROPROPOXYPHENE |PROPOXYPHENE (PRODUCT)
C0027415|T053||SNOMEDCT_US|NARCOTICS
C0027415|T053||SNOMEDCT_US|NARCOTIC
C0027415|T053||SNOMEDCT_US|NARCOTICS 
C2193937|T053||SNOMEDCT_US|SODIUM IODIDE + NIACINAMIDE HYDROIODIDE
C2193937|T053||SNOMEDCT_US|NARCOTICS SODIUM IODIDE + NIACINAMIDE HYDROIODIDE
C2193937|T053||SNOMEDCT_US|SODIUM IODIDE + NIACINAMIDE HYDROIODIDE 
C0355546|T053|322508000|SNOMEDCT_US|DEXTROMORAMIDE TARTRATE|DEXTROMORAMIDE TARTRATE (SUBSTANCE)
C0355546|T053|322508000|SNOMEDCT_US|DEXTROMORAMIDE TARTRATE |DEXTROMORAMIDE TARTRATE (SUBSTANCE)
C0355546|T053|322508000|SNOMEDCT_US|NARCOTICS DEXTROMORAMIDE TARTRATE|DEXTROMORAMIDE TARTRATE (SUBSTANCE)
C0355546|T053|322508000|SNOMEDCT_US|DEXTROMORAMIDE TARTRATE |DEXTROMORAMIDE TARTRATE (SUBSTANCE)
C0355546|T053|322508000|SNOMEDCT_US|TARTRATE, DEXTROMORAMIDE|DEXTROMORAMIDE TARTRATE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIACETYLMORPHINE HYDROCHLORIDE|DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIACETYLMORPHINE HYDROCHLORIDE |DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|HEROIN HYDROCHLORIDE|DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIAMORPHINE HYDROCHLORIDE|DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|HEROINE HYDROCHLORIDE|DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|MORPHINAN-3,6ALPHA-DIOL, 7,8-DIDEHYDRO-4,5ALPHA-EPOXY-17-METHYL-, MORPHINE, DIACETATE (ESTER), HYDROCHLORIDE|DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|HYDROCHLORIDE, HEROIN|DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIAMORPHINE HCL [COUGH]|DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIAMORPHINE HCL [COUGH] |DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIAMORPHINE HCL [ANALGESIC] |DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIAMORPHINE HCL [ANALGESIC]|DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIAMORPHINE HYDROCHLORIDE |DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIAMORPHINE HCL [ANALGESIC] |DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|DIAMORPHINE HCL [COUGH] |DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C0282128|T053|396019002|SNOMEDCT_US|HYDROCHLORIDE, DIACETYLMORPHINE|DIAMORPHINE HYDROCHLORIDE (SUBSTANCE)
C2194296|T053||SNOMEDCT_US|NARCOTICS ASPIRIN + CAFFEINE + OPIUM
C2194296|T053||SNOMEDCT_US|ASPIRIN + CAFFEINE + OPIUM 
C2194296|T053||SNOMEDCT_US|ASPIRIN + CAFFEINE + OPIUM
C2194297|T053||SNOMEDCT_US|ASPIRIN + PHENOBARBITAL
C2194297|T053||SNOMEDCT_US|ASPIRIN + PHENOBARBITAL 
C2194297|T053||SNOMEDCT_US|PHENOBARBITAL + ASPIRIN 
C2194297|T053||SNOMEDCT_US|PHENOBARBITAL + ASPIRIN
C2194297|T053||SNOMEDCT_US|NARCOTICS ASPIRIN + PHENOBARBITAL
C2194297|T053||SNOMEDCT_US|ASPIRIN / PHENOBARBITAL
C2146622|T053||SNOMEDCT_US|ACETAMINOPHEN + IBUPROFEN + CODEINE
C2146622|T053||SNOMEDCT_US|NARCOTICS ACETAMINOPHEN + IBUPROFEN + CODEINE
C2146622|T053||SNOMEDCT_US|ACETAMINOPHEN + IBUPROFEN + CODEINE 
C2146622|T053||SNOMEDCT_US|ACETAMINOPHEN / CODEINE / IBUPROFEN
C2117853|T053||SNOMEDCT_US|ACETAMINOPHEN + ASPIRIN + MEPROBAMATE + CAFFEINE + CODEINE 
C2117853|T053||SNOMEDCT_US|ACETAMINOPHEN + ASPIRIN + MEPROBAMATE + CAFFEINE + CODEINE
C1873942|T053||SNOMEDCT_US|ACETAMINOPHEN/ASPIRIN/CAFFEINE/CODEINE/SALICYLAMIDE
C1873942|T053||SNOMEDCT_US|ACETAMINOPHEN + ASPIRIN + SALICYLAMIDE + CAFFEINE + CODEINE
C1873942|T053||SNOMEDCT_US|ACETAMINOPHEN + ASPIRIN + SALICYLAMIDE + CAFFEINE + CODEINE 
C1873942|T053||SNOMEDCT_US|ACETAMINOPHEN / ASPIRIN / CAFFEINE / CODEINE / SALICYLAMIDE
C2194298|T053||SNOMEDCT_US|ALUMINUM ASPIRIN + ACETAMINOPHEN + CHLORPHENOXAMINE + PHENOBARBITAL 
C2194298|T053||SNOMEDCT_US|ALUMINUM ASPIRIN + ACETAMINOPHEN + CHLORPHENOXAMINE + PHENOBARBITAL
C2114801|T053||SNOMEDCT_US|PROMETHAZINE + ASPIRIN-PHENACETIN-CAFFEINE + DIHYDROCODEINE
C2114801|T053||SNOMEDCT_US|PROMETHAZINE + ASPIRIN-PHENACETIN-CAFFEINE + DIHYDROCODEINE 
C2114800|T053||SNOMEDCT_US|NARCOTICS PROMETHAZINE + APAP + CAFFEINE + DIHYDROCODEINE
C2114800|T053||SNOMEDCT_US|PROMETHAZINE + APAP + CAFFEINE + DIHYDROCODEINE
C2114800|T053||SNOMEDCT_US|PROMETHAZINE + APAP + CAFFEINE + DIHYDROCODEINE 
C1874363|T053||SNOMEDCT_US|ASPIRIN/CAFFEINE/DIHYDROCODEINE/PROMETHAZINE
C1874363|T053||SNOMEDCT_US|NARCOTICS POMETHAZINE + ASPIRIN + CAFFEINE + DIHYDROCODEINE
C1874363|T053||SNOMEDCT_US|PROMETHAZINE + ASPIRIN + CAFFEINE + DIHYDROCODEINE
C1874363|T053||SNOMEDCT_US|PROMETHAZINE + ASPIRIN + CAFFEINE + DIHYDROCODEINE 
C1874363|T053||SNOMEDCT_US|ASPIRIN / CAFFEINE / DIHYDROCODEINE / PROMETHAZINE
C1302959|T053|400776001|SNOMEDCT_US|PENTAZOCINE HYDROCHLORIDE + ASPIRIN (DISCONTINUED) |ASPIRIN + PENTAZOCINE HYDROCHLORIDE (PRODUCT)
C1302959|T053|400776001|SNOMEDCT_US|PENTAZOCINE HYDROCHLORIDE + ASPIRIN (DISCONTINUED)|ASPIRIN + PENTAZOCINE HYDROCHLORIDE (PRODUCT)
C1302959|T053|400776001|SNOMEDCT_US|ASPIRIN + PENTAZOCINE HYDROCHLORIDE |ASPIRIN + PENTAZOCINE HYDROCHLORIDE (PRODUCT)
C1302959|T053|400776001|SNOMEDCT_US|ASPIRIN + PENTAZOCINE HYDROCHLORIDE|ASPIRIN + PENTAZOCINE HYDROCHLORIDE (PRODUCT)
C2052847|T053||SNOMEDCT_US|PENTAZOCINE + ASPIRIN + CAFFEINE 
C2052847|T053||SNOMEDCT_US|PENTAZOCINE + ASPIRIN + CAFFEINE
C0030131|T053||SNOMEDCT_US|P CHLOROAMPHETAMINE
C0030131|T053||SNOMEDCT_US|P-CHLOROAMPHETAMINE
C0030131|T053||SNOMEDCT_US|P CHLORAMPHETAMINE
C0030131|T053||SNOMEDCT_US|PARA CHLOROAMPHETAMINE
C0030131|T053||SNOMEDCT_US|BENZENEETHANAMINE, 4-CHLORO-ALPHA-METHYL-
C0030131|T053||SNOMEDCT_US|CHLOROAMPHETAMINE P
C0030131|T053||SNOMEDCT_US|CHLORAMPHETAMINE P
C0030131|T053||SNOMEDCT_US|PCA
C0030131|T053||SNOMEDCT_US|4-CHLOROAMPHETAMINE
C0030131|T053||SNOMEDCT_US|ALPHA-METHYL-P-CHLOROPHENETHYLAMINE
C0030131|T053||SNOMEDCT_US|NARCOTICS PATIENT CONTROLLED ANESTHESIA (PCA) 
C0030131|T053||SNOMEDCT_US|NARCOTICS PCA
C0030131|T053||SNOMEDCT_US|NARCOTICS PATIENT CONTROLLED ANESTHESIA (PCA)
C0030131|T053||SNOMEDCT_US|PARACHLOROAMPHETAMINE
C0030131|T053||SNOMEDCT_US|P-CHLORAMPHETAMINE
C0030131|T053||SNOMEDCT_US|PARA-CHLOROAMPHETAMINE
C0030131|T053||SNOMEDCT_US|P-CHLOROAMPHETAMINE [CHEMICAL/INGREDIENT]
C2047970|T053||SNOMEDCT_US|IMED PANEL LOCKED
C2047970|T053||SNOMEDCT_US|NARCOTICS IMED PANEL LOCKED
C2047970|T053||SNOMEDCT_US|IMED PANEL LOCKED 
C0770427|T053||SNOMEDCT_US|ANILERIDINE HYDROCHLORIDE
C0770427|T053||SNOMEDCT_US|ANILERIDINE HYDROCHLORIDE (DISCONTINUED)
C0770427|T053||SNOMEDCT_US|NARCOTICS ANILERIDINE HYDROCHLORIDE (DISCONTINUED)
C0770427|T053||SNOMEDCT_US|ANILERIDINE HYDROCHLORIDE (DISCONTINUED) 
C0770428|T053||SNOMEDCT_US|ANILERIDINE PHOSPHATE (DISCONTINUED) 
C0770428|T053||SNOMEDCT_US|ANILERIDINE PHOSPHATE (DISCONTINUED)
C0770428|T053||SNOMEDCT_US|NARCOTICS ANILERIDINE PHOSPHATE (DISCONTINUED)
C0770428|T053||SNOMEDCT_US|ANILERIDINE PHOSPHATE
C0700525|T053|69241001|SNOMEDCT_US|BUTORPHANOL TARTRATE|BUTORPHANOL TARTRATE (SUBSTANCE)
C0700525|T053|69241001|SNOMEDCT_US|NARCOTICS BUTORPHANOL TARTRATE|BUTORPHANOL TARTRATE (SUBSTANCE)
C0700525|T053|69241001|SNOMEDCT_US|BUTORPHANOL TARTRATE |BUTORPHANOL TARTRATE (SUBSTANCE)
C0700525|T053|69241001|SNOMEDCT_US|BUTORPHANOL TARTRATE [CHEMICAL/INGREDIENT]|BUTORPHANOL TARTRATE (SUBSTANCE)
C0700525|T053|69241001|SNOMEDCT_US|(-)-17-(CYCLOBUTYLMETHYL)MORPHINAN-3,14-DIOL D-(-)-TARTRATE (1:1) (SALT)|BUTORPHANOL TARTRATE (SUBSTANCE)
C0700525|T053|69241001|SNOMEDCT_US|BUTORPHANOL TARTRATE |BUTORPHANOL TARTRATE (SUBSTANCE)
C0700562|T053|96184001|SNOMEDCT_US|ALFENTANIL HYDROCHLORIDE|ALFENTANIL HYDROCHLORIDE (SUBSTANCE)
C0700562|T053|96184001|SNOMEDCT_US|ALFENTANIL HYDROCHLORIDE |ALFENTANIL HYDROCHLORIDE (SUBSTANCE)
C0700562|T053|96184001|SNOMEDCT_US|ALFENTANIL HYDROCHLORIDE [CHEMICAL/INGREDIENT]|ALFENTANIL HYDROCHLORIDE (SUBSTANCE)
C0700562|T053|96184001|SNOMEDCT_US|ALFENTANIL HYDROCHLORIDE - CHEMICAL|ALFENTANIL HYDROCHLORIDE (SUBSTANCE)
C0700562|T053|96184001|SNOMEDCT_US|ALFENTANIL HYDROCHLORIDE - CHEMICAL |ALFENTANIL HYDROCHLORIDE (SUBSTANCE)
C0700562|T053|96184001|SNOMEDCT_US|ALFENTANIL HYDROCHLORIDE |ALFENTANIL HYDROCHLORIDE (SUBSTANCE)
C2001271|T053|441757005|SNOMEDCT_US|TAPENTADOL|TAPENTADOL (SUBSTANCE)
C2001271|T053|441757005|SNOMEDCT_US|TAPENTADOL |TAPENTADOL (SUBSTANCE)
C2001271|T053|441757005|SNOMEDCT_US|TAPENTADOL |TAPENTADOL (SUBSTANCE)
C2001271|T053|441757005|SNOMEDCT_US|3-((1R,2R)-3-(DIMETHYLAMINO)-1-ETHYL-2-METHYLPROPYL)PHENOL|TAPENTADOL (SUBSTANCE)
C2001271|T053|441757005|SNOMEDCT_US|TAPENTADOL |TAPENTADOL (SUBSTANCE)
C2001271|T053|441757005|SNOMEDCT_US|NARCOTICS TAPENTADOL|TAPENTADOL (SUBSTANCE)
C0306074|T053||SNOMEDCT_US|EMPIRIN WITH CODEINE
C0306074|T053||SNOMEDCT_US|NARCOTICS ASPIRIN + CODEINE (EMPIRIN WITH CODEINE)
C0306074|T053||SNOMEDCT_US|ASPIRIN + CODEINE (EMPIRIN WITH CODEINE) 
C0306074|T053||SNOMEDCT_US|ASPIRIN + CODEINE (EMPIRIN WITH CODEINE)
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN/CODEINE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|PARACETAMOL +CODEINE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|PARACETAMOL +CODIENE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|CODEINE PHOSPHATE + ACETAMINOPHEN|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|CODEINE PHOSPHATE + ACETAMINOPHEN |PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|NARCOTICS ACETAMINOPHEN + CODEINE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN + CODEINE |PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN + CODEINE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN-CODEINE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN-CODEINE PHOSPHATE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|CO-CODAMOL|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN - CODEINE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN, CODEINE DRUG COMBINATION|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|COCODAMOL|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN+CODEINE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN / CODEINE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|PARACETAMOL + CODEINE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|PARACETAMOL + CODEINE PHOSPHATE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN + CODEINE PHOSPHATE |PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN + CODEINE PHOSPHATE|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|CO-CODAMOL |PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN #3|PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|CO-CODAMOL |PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN + CODEINE |PARACETAMOL +CODIENE
C2351132|T053|412556009|SNOMEDCT_US|ACETAMINOPHEN WITH CODEINE|PARACETAMOL +CODIENE
C0724655|T053|37451001|SNOMEDCT_US|LAUDANUM|LAUDANUM (SUBSTANCE)
C0724655|T053|37451001|SNOMEDCT_US|OPIUM TINCTURE|LAUDANUM (SUBSTANCE)
C0724655|T053|37451001|SNOMEDCT_US|TINCTURE OF OPIUM|LAUDANUM (SUBSTANCE)
C0724655|T053|37451001|SNOMEDCT_US|NARCOTICS TINCTURE OF OPIUM|LAUDANUM (SUBSTANCE)
C0724655|T053|37451001|SNOMEDCT_US|TINCTURE OF OPIUM |LAUDANUM (SUBSTANCE)
C0724655|T053|37451001|SNOMEDCT_US|LAUDANUM |LAUDANUM (SUBSTANCE)
C0724655|T053|37451001|SNOMEDCT_US|DTO|LAUDANUM (SUBSTANCE)
C0724655|T053|37451001|SNOMEDCT_US|DEODORIZED TINCTURE OF OPIUM|LAUDANUM (SUBSTANCE)
C2013185|T053||SNOMEDCT_US|OPIATE ALKALOID HYDROCHLORIDE (PANTOPAN INJECTABLE) 
C2013185|T053||SNOMEDCT_US|OPIATE ALKALOID HYDROCHLORIDE (PANTOPAN INJECTABLE)
C2066455|T053||SNOMEDCT_US|NARCOTIC ANTITUSSIVES
C2066455|T053||SNOMEDCT_US|NARCOTIC ANTITUSSIVES 
C0282275|T053|69899006|SNOMEDCT_US|OXYMORPHONE HYDROCHLORIDE|OXYMORPHONE HYDROCHLORIDE (SUBSTANCE)
C0282275|T053|69899006|SNOMEDCT_US|4,5-ALPHA-EPOXY-3,14-DIHYDROXY-17-METHYLMORPHINAN-6-ONE HYDROCHLORIDE|OXYMORPHONE HYDROCHLORIDE (SUBSTANCE)
C0282275|T053|69899006|SNOMEDCT_US|OXYMORPHONE HYDROCHLORIDE |OXYMORPHONE HYDROCHLORIDE (SUBSTANCE)
C0282275|T053|69899006|SNOMEDCT_US|NARCOTICS OXYMORPHONE HYDROCHLORIDE|OXYMORPHONE HYDROCHLORIDE (SUBSTANCE)
C0282275|T053|69899006|SNOMEDCT_US|OXYMORPHONE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|OXYMORPHONE HYDROCHLORIDE (SUBSTANCE)
C0282275|T053|69899006|SNOMEDCT_US|OXYMORPHONE HCL|OXYMORPHONE HYDROCHLORIDE (SUBSTANCE)
C0282275|T053|69899006|SNOMEDCT_US|OXYMORPHONE HYDROCHLORIDE |OXYMORPHONE HYDROCHLORIDE (SUBSTANCE)
C0717478|T053|400609000|SNOMEDCT_US|BELLADONNA/OPIUM|OPIUM+BELLADONNA (PRODUCT)
C0717478|T053|400609000|SNOMEDCT_US|NARCOTICS OPIUM + BELLADONNA|OPIUM+BELLADONNA (PRODUCT)
C0717478|T053|400609000|SNOMEDCT_US|OPIUM + BELLADONNA |OPIUM+BELLADONNA (PRODUCT)
C0717478|T053|400609000|SNOMEDCT_US|OPIUM + BELLADONNA|OPIUM+BELLADONNA (PRODUCT)
C0717478|T053|400609000|SNOMEDCT_US|BELLADONNA-OPIUM|OPIUM+BELLADONNA (PRODUCT)
C0717478|T053|400609000|SNOMEDCT_US|OPIUM+BELLADONNA |OPIUM+BELLADONNA (PRODUCT)
C0717478|T053|400609000|SNOMEDCT_US|OPIUM+BELLADONNA|OPIUM+BELLADONNA (PRODUCT)
C0700533|T053|83929000|SNOMEDCT_US|HYDROMORPHONE HYDROCHLORIDE|DIHYDROMORPHINONE HYDROCHLORIDE
C0700533|T053|83929000|SNOMEDCT_US|HYDROMORPHONE HYDROCHLORIDE |DIHYDROMORPHINONE HYDROCHLORIDE
C0700533|T053|83929000|SNOMEDCT_US|HYDROMORPHONE HYDROCHLORIDE [CHEMICAL/INGREDIENT]|DIHYDROMORPHINONE HYDROCHLORIDE
C0700533|T053|83929000|SNOMEDCT_US|HYDROMORPHONE HCL|DIHYDROMORPHINONE HYDROCHLORIDE
C0700533|T053|83929000|SNOMEDCT_US|NARCOTICS HYDROMORPHONE HCL|DIHYDROMORPHINONE HYDROCHLORIDE
C0700533|T053|83929000|SNOMEDCT_US|HYDROMORPHONE HCL |DIHYDROMORPHINONE HYDROCHLORIDE
C0700533|T053|83929000|SNOMEDCT_US|HYDROMORPHONE HYDROCHLORIDE |DIHYDROMORPHINONE HYDROCHLORIDE
C0700533|T053|83929000|SNOMEDCT_US|HYDROMORPHONE HYDROCHLORIDE |DIHYDROMORPHINONE HYDROCHLORIDE
C0700533|T053|83929000|SNOMEDCT_US|DIHYDROMORPHINONE HYDROCHLORIDE|DIHYDROMORPHINONE HYDROCHLORIDE
C2928489|T053||SNOMEDCT_US|ACETAMINOPHEN / CHLORPHENIRAMINE / CODEINE
C2928489|T053||SNOMEDCT_US|ACETAMINOPHEN/CHLORPHENIRAMINE/CODEINE
C2928489|T053||SNOMEDCT_US|ACETAMINOPHEN + CHLORPHENIRAMINE + CODEINE 
C2928489|T053||SNOMEDCT_US|ACETAMINOPHEN + CHLORPHENIRAMINE + CODEINE
C2928489|T053||SNOMEDCT_US|NARCOTICS ACETAMINOPHEN + CHLORPHENIRAMINE + CODEINE
C0058763|T053||SNOMEDCT_US|14-HYDROXYDIHYDRO-6 BETA-THEBAINOL 4-METHYL ETHER
C0058763|T053||SNOMEDCT_US|3,4-DIMETHOXY-17-METHYLMORPHINAN-6 BETA,14-DIOL
C0058763|T053||SNOMEDCT_US|DROTEBANOL
C0058763|T053||SNOMEDCT_US|OXYMETHEBANOL
C0002772|T053||SNOMEDCT_US|ANALGESICS, OPIOID
C0002772|T053||SNOMEDCT_US|OPIOID ANALGESICS
C0002772|T053||SNOMEDCT_US|[CN101] OPIOID ANALGESICS
C0049689|T053|118290009|SNOMEDCT_US|6-(0-ACETYL)MORPHINE|6-O-MONOACETYLMORPHINE (SUBSTANCE)
C0049689|T053|118290009|SNOMEDCT_US|6-ACETYLMORPHINE|6-O-MONOACETYLMORPHINE (SUBSTANCE)
C0049689|T053|118290009|SNOMEDCT_US|6-MONOACETYLMORPHINE|6-O-MONOACETYLMORPHINE (SUBSTANCE)
C0049689|T053|118290009|SNOMEDCT_US|6-O-MONOACETYLMORPHINE|6-O-MONOACETYLMORPHINE (SUBSTANCE)
C0049689|T053|118290009|SNOMEDCT_US|MORPHINE-6-ACETATE|6-O-MONOACETYLMORPHINE (SUBSTANCE)
C0049689|T053|118290009|SNOMEDCT_US|6-MAM CPD|6-O-MONOACETYLMORPHINE (SUBSTANCE)
C0049689|T053|118290009|SNOMEDCT_US|MONOACETYLMORPHINE|6-O-MONOACETYLMORPHINE (SUBSTANCE)
C0049689|T053|118290009|SNOMEDCT_US|6-O-MONOACETYLMORPHINE |6-O-MONOACETYLMORPHINE (SUBSTANCE)
C0049689|T053|118290009|SNOMEDCT_US|ACETYLMORPHINE|6-O-MONOACETYLMORPHINE (SUBSTANCE)
C1992537|T053||SNOMEDCT_US|METHYLFENTANYL &#X7C; BLD-SER-PLAS
C1993205|T053||SNOMEDCT_US|NARCOTICS AND OPIOIDS &#X7C; URINE
C0066619|T053|725692004|SNOMEDCT_US|16,17-DIDEHYDRO-9,17-DIMETHOXY-17,18-SECO-20-ALPHA-YOHIMBAN-16-CARBOXYLIC ACID METHYL ESTER|MITRAGYNINE (SUBSTANCE)
C0066619|T053|725692004|SNOMEDCT_US|MITRAGYNINE|MITRAGYNINE (SUBSTANCE)
C0041029|T053|96180005|SNOMEDCT_US|TRIMEPERIDINE|TRIMEPERIDINE (SUBSTANCE)
C0041029|T053|96180005|SNOMEDCT_US|TRIPETHIDINE|TRIMEPERIDINE (SUBSTANCE)
C0041029|T053|96180005|SNOMEDCT_US|TRIMEPERIDINE |TRIMEPERIDINE (SUBSTANCE)
C0058056|T053|387322000|SNOMEDCT_US|DIHYDROCODEINE|DIHYDROCODEINE (SUBSTANCE)
C0058056|T053|387322000|SNOMEDCT_US|DIHYDROCODEINE ACID|DIHYDROCODEINE (SUBSTANCE)
C0058056|T053|387322000|SNOMEDCT_US|MORPHINAN-6-ALPHA-OL, 4,5-ALPHA-EPOXY-3-METHOXY-17-METHYL-|DIHYDROCODEINE (SUBSTANCE)
C0058056|T053|387322000|SNOMEDCT_US|DIHYDROCODEINE [CHEMICAL/INGREDIENT]|DIHYDROCODEINE (SUBSTANCE)
C0058056|T053|387322000|SNOMEDCT_US|DIHYDROCODEINE |DIHYDROCODEINE (SUBSTANCE)
C0058056|T053|387322000|SNOMEDCT_US|DIHYDROCODEINE |DIHYDROCODEINE (SUBSTANCE)
C1993204|T053||SNOMEDCT_US|NARCOTICS AND OPIOIDS &#X7C; GASTRIC FLUID
C0058410|T053|387226000|SNOMEDCT_US|4,4-DIPHENYL-6-PIPERIDINO-3-HEPTANONE|DIPIPANONE (SUBSTANCE)
C0058410|T053|387226000|SNOMEDCT_US|DIPIPANONE|DIPIPANONE (SUBSTANCE)
C0058410|T053|387226000|SNOMEDCT_US|PHENYLPIPERONE|DIPIPANONE (SUBSTANCE)
C0058410|T053|387226000|SNOMEDCT_US|DIPIPANONE |DIPIPANONE (SUBSTANCE)
C0058410|T053|387226000|SNOMEDCT_US|DIPIPANONE |DIPIPANONE (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|ANTAGONISTS, NARCOTIC|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|NARCOTIC ANTAGONISTS|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|NARCOTIC ANTAGONIST|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|ANTAGONISTS, OPIOID|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|OPIOID ANTAG|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|NARCOTIC ANTAG|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|RECEPTOR ANTAGONISTS, OPIOID|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|ANTAGONISTS, OPIOID RECEPTOR|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|OPIOID ANTAGONISTS|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|OPIOID RECEPTOR ANTAGONISTS|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|OPIOID ANTAGONIST|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|OPIATE ANTAGONIST |OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|OPIATE ANTAGONIST |OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|OPIATE ANTAGONIST|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|OPIATE ANTAGONIST, NOS|OPIATE ANTAGONIST (SUBSTANCE)
C0027410|T053|14103001|SNOMEDCT_US|OPIATE ANTAGONISTS|OPIATE ANTAGONIST (SUBSTANCE)
C0068699|T053|96181009|SNOMEDCT_US|BIS(NICOTINYL)MORPHINE|NICOMORPHINE (SUBSTANCE)
C0068699|T053|96181009|SNOMEDCT_US|MORPHINE DINICOTINATE|NICOMORPHINE (SUBSTANCE)
C0068699|T053|96181009|SNOMEDCT_US|NICOMORPHINE|NICOMORPHINE (SUBSTANCE)
C0068699|T053|96181009|SNOMEDCT_US|NICOMORPHINE |NICOMORPHINE (SUBSTANCE)
C0051908|T053|55793008|SNOMEDCT_US|ANILERIDINE|ANILERIDINE (SUBSTANCE)
C0051908|T053|55793008|SNOMEDCT_US|ANILERIDINE |ANILERIDINE (SUBSTANCE)
C1993203|T053||SNOMEDCT_US|NARCOTICS AND OPIOIDS &#X7C; BLD-SER-PLAS
C1993202|T053||SNOMEDCT_US|NARCOTICS AND OPIOIDS &#124; BILE FLUID
C1993202|T053||SNOMEDCT_US|NARCOTICS AND OPIOIDS &#X7C; BILE FLUID
C3870663|T053||SNOMEDCT_US|MITRAGYNINE+7-HYDROXYMITRAGYNINE &#X7C; URINE
C3870618|T053||SNOMEDCT_US|TAPENTADOL GLUCURONIDE &#X7C; URINE
C0027409|T053|360204007|SNOMEDCT_US|NARCOTIC ANALGESICS|NARCOTIC ANALGESIC PRODUCT
C0027409|T053|360204007|SNOMEDCT_US|NARCOTIC AGONISTS |NARCOTIC ANALGESIC PRODUCT
C0027409|T053|360204007|SNOMEDCT_US|NARCOTIC AGONISTS|NARCOTIC ANALGESIC PRODUCT
C0027409|T053|360204007|SNOMEDCT_US|NARCOTIC ANALGESIC|NARCOTIC ANALGESIC PRODUCT
C0027409|T053|360204007|SNOMEDCT_US|NARCOTIC ANALGESIC PRODUCT|NARCOTIC ANALGESIC PRODUCT
C0027409|T053|360204007|SNOMEDCT_US|ANALGESICS, NARCOTIC|NARCOTIC ANALGESIC PRODUCT
C0027409|T053|360204007|SNOMEDCT_US|NARCOTIC ANALGESIC AGENT|NARCOTIC ANALGESIC PRODUCT
C0058916|T053|373563003|SNOMEDCT_US|3 BETA-HYDROXY-2 BETA-TROPANECARBOXYLIC ACID|ECGONINE (SUBSTANCE)
C0058916|T053|373563003|SNOMEDCT_US|ECGONINE|ECGONINE (SUBSTANCE)
C0058916|T053|373563003|SNOMEDCT_US|ECGONINE |ECGONINE (SUBSTANCE)
C0058916|T053|373563003|SNOMEDCT_US|ECGONINE |ECGONINE (SUBSTANCE)
C0068953|T053||SNOMEDCT_US|6-(METHYLAMINO)-4,4-DIPHENYL-3-HEPTANOL ACETATE
C0068953|T053||SNOMEDCT_US|ALPHA-ETHYL-BETA- (2-(METHYLAMINO)PROPYL)-BETA-PHENYLBENZENEETHANOL, ACETATE (ESTER)
C0068953|T053||SNOMEDCT_US|PARACYMETHADOL
C0058841|T053||SNOMEDCT_US|DYNORPHIN (1-13)
C0058917|T053||SNOMEDCT_US|ECGONINE METHYL ESTER
C0058917|T053||SNOMEDCT_US|METHYL ECGONINE
C0242402|T053|404642006|SNOMEDCT_US|OPIOIDS|OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIATE AGONIST AGENT|OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIOID|OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIATE AGONIST |OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIATE AGONIST|OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIOID PRODUCT|OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIATE AGONIST PRODUCT|OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIATE AGONIST |OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIOID |OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIATE PRODUCT|OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIATE AGONIST, NOS|OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIATE |OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIOID |OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIOID AGENT|OPIOID RECEPTOR AGONIST
C0242402|T053|404642006|SNOMEDCT_US|OPIATE AGONISTS|OPIOID RECEPTOR AGONIST
C0430053|T053|252158001|SNOMEDCT_US|OPIOID SCREENING |OPIOID SCREENING (PROCEDURE)
C0430053|T053|252158001|SNOMEDCT_US|OPIOID SCREENING|OPIOID SCREENING (PROCEDURE)
C0038388|T053||SNOMEDCT_US|DRUGS, STREET
C0038388|T053||SNOMEDCT_US|STREET DRUGS
C0086190|T053|77657003|SNOMEDCT_US|ABUSE DRUGS|ILLEGAL DRUG (SUBSTANCE)
C0086190|T053|77657003|SNOMEDCT_US|DRUGS, ILLICIT|ILLEGAL DRUG (SUBSTANCE)
C0086190|T053|77657003|SNOMEDCT_US|ILLICIT DRUGS|ILLEGAL DRUG (SUBSTANCE)
C0086190|T053|77657003|SNOMEDCT_US|DRUGS OF ABUSE|ILLEGAL DRUG (SUBSTANCE)
C0086190|T053|77657003|SNOMEDCT_US|ILLEGAL DRUG |ILLEGAL DRUG (SUBSTANCE)
C0086190|T053|77657003|SNOMEDCT_US|ILLEGAL DRUG|ILLEGAL DRUG (SUBSTANCE)
C0086190|T053|77657003|SNOMEDCT_US|ILLEGAL DRUG, NOS|ILLEGAL DRUG (SUBSTANCE)
C0086190|T053|77657003|SNOMEDCT_US|ILLEGAL DRUG |ILLEGAL DRUG (SUBSTANCE)
C2911101|T053||SNOMEDCT_US|DRUG ABUSE COUNSELING AND SURVEILLANCE OF DRUG ABUSER
