C2169446|T053||SNOMEDCT_US|SEX WITH AN HCV INFECTED PERSON
C2169446|T053||SNOMEDCT_US|SEX WITH AN HCV PARTNER
C2169446|T053||SNOMEDCT_US|SEX WITH AN HCV PERSON
