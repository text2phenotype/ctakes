C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISEASE|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C1963138|T047||SNOMEDCT_US|HYPERTENSION ADVERSE EVENT
C0085580|T047|59621000|SNOMEDCT_US|ESSENTIAL HYPERTENSION|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|PRIMARY HYPERTENSION|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|ESSENTIAL (PRIMARY) HYPERTENSION|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|HYPERTENSION, ESSENTIAL|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|IDIOPATHIC HYPERTENSION|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|ESSENTIAL HYPERTENSION |ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|HYPERTENSION NOS|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|HYPERTENSION;ESSENTIAL|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|ESSENTIAL HYPERTENSION |ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|ESSENTIAL HYPERTENSION NOS |ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|ESSENTIAL HYPERTENSION NOS|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|ESSENTIAL HYPERTENSION, UNSPECIFIED|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|UNSPECIFIED ESSENTIAL HYPERTENSION|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|SYSTEMIC PRIMARY ARTERIAL HYPERTENSION|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|ESSENTIAL HYPERTENSION, NOS|ESSENTIAL HYPERTENSION (DISORDER)
C0085580|T047|59621000|SNOMEDCT_US|PRIMARY HYPERTENSION, NOS|ESSENTIAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|HYPERTENSION, RENAL|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|HYPERTENSIONS, RENAL|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|RENAL HYPERTENSIONS|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|RENAL HYPERTENSION|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|HYPERTENSION, RENAL [DISEASE/FINDING]|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|HYPERTENSION;CARDIORENAL|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|SECONDARY HYPERTENSION TO RENAL DISORDERS|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|HYPERTENSION SECONDARY TO RENAL DISORDERS|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|HYPERTENSION SECONDARY TO RENAL DISORDERS |RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|RENAL HYPERTENSION NOS|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|HYPERTENSION RENAL|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|RENAL HYPERTENSION |RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|CARDIORENAL; HYPERTENSION|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|HYPERTENSION; RENAL|RENAL HYPERTENSION (DISORDER)
C0020544|T047|28119000|SNOMEDCT_US|RENAL; HYPERTENSION|RENAL HYPERTENSION (DISORDER)
C0264641|T047|59997006|SNOMEDCT_US|ENDOCRINE HYPERTENSION|ENDOCRINE HYPERTENSION (DISORDER)
C0264641|T047|59997006|SNOMEDCT_US|ADRENAL HYPERTENSION|ENDOCRINE HYPERTENSION (DISORDER)
C0264641|T047|59997006|SNOMEDCT_US|ENDOCRINE HYPERTENSION |ENDOCRINE HYPERTENSION (DISORDER)
C0264641|T047|59997006|SNOMEDCT_US|ENDOCRINE; DISORDER HYPERTENSION|ENDOCRINE HYPERTENSION (DISORDER)
C0264641|T047|59997006|SNOMEDCT_US|HYPERTENSION; ENDOCRINE DISORDERS|ENDOCRINE HYPERTENSION (DISORDER)
C0596515|T047||SNOMEDCT_US|ENVIRONMENT ASSOCIATED HYPERTENSION
C0598428|T047||SNOMEDCT_US|FAMILIAL HYPERTENSION
C0598428|T047||SNOMEDCT_US|CONGENITAL HYPERTENSION
C0598428|T047||SNOMEDCT_US|GENETIC HYPERTENSION
C0597048|T047||SNOMEDCT_US|NEUROGENIC HYPERTENSION
C0596088|T047||SNOMEDCT_US|ANGIOTENSIN/RENIN/ALDOSTERONE HYPERTENSION
C0810002|T047||SNOMEDCT_US|HYPERTENSION WITH COMPLICATIONS AND SECONDARY HYPERTENSION
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE|HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE |HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE NOS|HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSION;HEART DISEASE|HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE NOS |HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE |HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE, UNSPECIFIED|HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|UNSPECIFIED HYPERTENSIVE HEART DISEASE|HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSIVE CARDIOPATHY|HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSIVE CARDIOVASCULAR DISEASE|HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HHD - HYPERTENSIVE HEART DISEASE|HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HEART; HYPERTENSION|HYPERTENSIVE HEART DISEASE (DISORDER)
C0152105|T047|64715009|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE, NOS|HYPERTENSIVE HEART DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE NEPHROPATHY|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE NEPHROPATHY |HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE KIDNEY DISEASE |HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE KIDNEY DISEASE|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE NOS|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSION;RENAL DISEASE|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSION;NEPHROPATHY|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE NOS |HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE, UNSPECIFIED|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|NEPHROPATHY HYPERTENSIVE|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE |HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|RENAL DISEASE; HYPERTENSION|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE NEPHROPATHY, NOS|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE, NOS|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0848548|T047|38481006|SNOMEDCT_US|HYPERTENSION SECONDARY TO RENAL DISEASE|HYPERTENSIVE RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE NOS|HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE, UNSPECIFIED|HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|CARDIORENAL DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE |HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE NOS |HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE; WITH HYPERTENSIVE KIDNEY DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|KIDNEY; HYPERTENSION, WITH HYPERTENSIVE HEART DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|CARDIORENAL DISEASE, NOS|HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE, NOS|HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155601|T047|86234004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE [DUP] |HYPERTENSIVE HEART AND RENAL DISEASE (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|SECONDARY HYPERTENSION|SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|SECONDARY HYPERTENSION, UNSPECIFIED|SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|UNSPECIFIED SECONDARY HYPERTENSION |SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|SECONDARY HYPERTENSION |SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|UNSPECIFIED SECONDARY HYPERTENSION|SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|SECONDARY HYPERTENSION |SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|SECONDARY HYPERTENSION NOS|SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|SECONDARY HYPERTENSION NOS |SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|HYPERTENSION SECONDARY|SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|HYPERTENSION; SECONDARY|SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|SECONDARY; HYPERTENSION|SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|SECONDARY HYPERTENSION, NOS|SECONDARY HYPERTENSION (DISORDER)
C0155616|T047|31992008|SNOMEDCT_US|HYPERTENSION;SECONDARY|SECONDARY HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|HYPERTENSION, MALIGNANT|MALIGNANT HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|MALIGNANT HYPERTENSION|MALIGNANT HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|ACCELERATED HYPERTENSION|MALIGNANT HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|HYPERTENSION, MALIGNANT [DISEASE/FINDING]|MALIGNANT HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|HYPERTENSION;MALIGNANT|MALIGNANT HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|MALIGNANT HYPERTENSION |MALIGNANT HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|HYPERTENSION (SYSTEMIC) MALIGNANT|MALIGNANT HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|MALIGNANT HYPERTENSION |MALIGNANT HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|HYPERTENSION MALIGNANT|MALIGNANT HYPERTENSION (DISORDER)
C0020540|T047|70272006|SNOMEDCT_US|MALIGNANT HYPERTENSION NOS|MALIGNANT HYPERTENSION (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HIGH BLOOD PRESSURE|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSION|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISEASES|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|SYSTEMIC HYPERTENSION|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISORDER, SYSTEMIC ARTERIAL|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HTN|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERPIESIA|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERPIESIS|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISEASE|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|SYSTEMIC HTN|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|SYSTEMIC HYPERTENSION |(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HBP|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
# C0020538|T047|266287006|SNOMEDCT_US|HT|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|BLOOD PRESSURE, HIGH|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSION [DISEASE/FINDING]|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISEASES (I10-I15)|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|COMPLICATIONS AFFECTING OTHER SPECIFIED BODY SYSTEMS, NOT ELSEWHERE CLASSIFIED, HYPERTENSION|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISEASE NOS |(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISEASE NOS|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSION NOS|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISEASE |(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|(HYPERTENSIVE DISEASE) OR (HYPERTENSION)|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) |(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|[X]HYPERTENSIVE DISEASES |(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|[X]HYPERTENSIVE DISEASES|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|INCREASED BLOOD PRESSURE|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|BLOOD PRESSURE, INCREASED|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|PRESSURE, HIGH BLOOD|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|ELEVATED BLOOD PRESSURE|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSION ARTERIAL|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|BLOOD PRESSURE HIGH|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|CARDIO/PULM: HYPERTENSIVE DISORDER|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE VASCULAR DEGENERATION|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE VASCULAR DISEASE|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|BP - HIGH BLOOD PRESSURE|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HIGH BLOOD PRESSURE DISORDER|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|SYSTEMIC ARTERIAL HYPERTENSION|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HBP - HIGH BLOOD PRESSURE|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|BP+ - HYPERTENSION|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HT - HYPERTENSION|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISORDER, SYSTEMIC ARTERIAL |(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISORDER|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HTN - HYPERTENSION|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|BLOOD PRESSURE; HIGH|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HIGH; ARTERIAL TENSION|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HIGH; BLOOD PRESSURE|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSION, NOS|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HYPERTENSIVE DISEASE, NOS|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|RAISED BLOOD PRESSURE |(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|BLOOD PRESSURES, HIGH|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|HIGH BLOOD PRESSURES|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0020538|T047|266287006|SNOMEDCT_US|VASCULAR HYPERTENSIVE DISORDER|(HYPERTENSIVE DISEASE) OR (HYPERTENSION) (DISORDER)
C0745138|T047|443482000|SNOMEDCT_US|HYPERTENSIVE URGENCY |HYPERTENSIVE URGENCY (DISORDER)
C0745138|T047|443482000|SNOMEDCT_US|HYPERTENSIVE URGENCY|HYPERTENSIVE URGENCY (DISORDER)
C0745138|T047|443482000|SNOMEDCT_US|HYPERTENSIVE URGENCY |HYPERTENSIVE URGENCY (DISORDER)
C3695318|T047|104931000119100|SNOMEDCT_US|HYPERTENSIVE CHRONIC KIDNEY DISEASE|CHRONIC KIDNEY DISEASE DUE TO HYPERTENSION (DISORDER)
C3695318|T047|104931000119100|SNOMEDCT_US|HYPERTENSIVE CHRONIC KIDNEY DISEASE |CHRONIC KIDNEY DISEASE DUE TO HYPERTENSION (DISORDER)
C3695318|T047|104931000119100|SNOMEDCT_US|HYPERTENSIVE CHRONIC KIDNEY DISEASE NOS|CHRONIC KIDNEY DISEASE DUE TO HYPERTENSION (DISORDER)
C3695318|T047|104931000119100|SNOMEDCT_US|CHRONIC KIDNEY DISEASE DUE TO HYPERTENSION|CHRONIC KIDNEY DISEASE DUE TO HYPERTENSION (DISORDER)
C3695318|T047|104931000119100|SNOMEDCT_US|CHRONIC KIDNEY DISEASE DUE TO HYPERTENSION |CHRONIC KIDNEY DISEASE DUE TO HYPERTENSION (DISORDER)
C3695318|T047|104931000119100|SNOMEDCT_US|HYPERTENSIVE CHRONIC KIDNEY DISEASE |CHRONIC KIDNEY DISEASE DUE TO HYPERTENSION (DISORDER)
C1719469|T047|8501000119104|SNOMEDCT_US|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE (DISORDER)
C1719469|T047|8501000119104|SNOMEDCT_US|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE |HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE (DISORDER)
C1719469|T047|8501000119104|SNOMEDCT_US|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE |HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE (DISORDER)
C2169401|T047||SNOMEDCT_US|REACTIVE HYPERTENSION
C2169401|T047||SNOMEDCT_US|REACTIVE HYPERTENSION 
C1171349|T047||SNOMEDCT_US|KALLIKREIN ATTENUATED HYPERTENSION
C1171349|T047||SNOMEDCT_US|KALLIKREIN HYPERTENSION
C2931778|T047||SNOMEDCT_US|TACHYCARDIA HYPERTENSION MICROPHTHALMOS HYPERGLYCINURIA
C0152132|T047|6962006|SNOMEDCT_US|HYPERTENSIVE RETINOPATHY|HYPERTENSIVE RETINOPATHY (DISORDER)
C0152132|T047|6962006|SNOMEDCT_US|HYPERTENSIVE RETINOPATHY |HYPERTENSIVE RETINOPATHY (DISORDER)
C0152132|T047|6962006|SNOMEDCT_US|RETINOPATHY HYPERTENSIVE|HYPERTENSIVE RETINOPATHY (DISORDER)
C0152132|T047|6962006|SNOMEDCT_US|RETINOPATHY, HYPERTENSIVE|HYPERTENSIVE RETINOPATHY (DISORDER)
C0152132|T047|6962006|SNOMEDCT_US|HYPERTENSIVE RETINOPATHIES|HYPERTENSIVE RETINOPATHY (DISORDER)
C0152132|T047|6962006|SNOMEDCT_US|RETINOPATHIES, HYPERTENSIVE|HYPERTENSIVE RETINOPATHY (DISORDER)
C0152132|T047|6962006|SNOMEDCT_US|RETINOPATHY;HYPERTENSIVE|HYPERTENSIVE RETINOPATHY (DISORDER)
C0152132|T047|6962006|SNOMEDCT_US|HYPERTENSIVE RETINOPATHY [DISEASE/FINDING]|HYPERTENSIVE RETINOPATHY (DISORDER)
C0152132|T047|6962006|SNOMEDCT_US|HYPERTENSIVE RETINOPATHY |HYPERTENSIVE RETINOPATHY (DISORDER)
C0152132|T047|6962006|SNOMEDCT_US|HYPERTENSIVE RETINOPATHY [AMBIGUOUS]|HYPERTENSIVE RETINOPATHY (DISORDER)
C0745121|T047||SNOMEDCT_US|IATROGENIC HYPERTENSION 
C0745121|T047||SNOMEDCT_US|IATROGENIC HYPERTENSION
C3178811|T047||SNOMEDCT_US|HYPERTENSION, MASKED
C3178811|T047||SNOMEDCT_US|HYPERTENSIONS, MASKED
C3178811|T047||SNOMEDCT_US|MASKED HYPERTENSION
C3178811|T047||SNOMEDCT_US|MASKED HYPERTENSIONS
C3178811|T047||SNOMEDCT_US|MASKED HYPERTENSION [DISEASE/FINDING]
C2186383|T047||SNOMEDCT_US|REPORTED A HISTORY OF INTERMITTENT HYPERTENSION
C2186383|T047||SNOMEDCT_US|REPORTED HISTORY OF INTERMITTENT HYPERTENSION 
C2186383|T047||SNOMEDCT_US|REPORTED HISTORY OF INTERMITTENT HYPERTENSION
C2186383|T047||SNOMEDCT_US|INTERMITTENT HYPERTENSION
C0745136|T047|132721000119104|SNOMEDCT_US|HYPERTENSIVE EMERGENCY |HYPERTENSIVE EMERGENCY (DISORDER)
C0745136|T047|132721000119104|SNOMEDCT_US|HYPERTENSIVE EMERGENCY|HYPERTENSIVE EMERGENCY (DISORDER)
C0155583|T047|1201005|SNOMEDCT_US|BENIGN ESSENTIAL HYPERTENSION |BENIGN ESSENTIAL HYPERTENSION
C0155583|T047|1201005|SNOMEDCT_US|BENIGN ESSENTIAL HYPERTENSION |BENIGN ESSENTIAL HYPERTENSION
C0155583|T047|1201005|SNOMEDCT_US|BENIGN ESSENTIAL HYPERTENSION|BENIGN ESSENTIAL HYPERTENSION
C0155583|T047|1201005|SNOMEDCT_US|BENIGN HYPERTENSION|BENIGN ESSENTIAL HYPERTENSION
C0155583|T047|1201005|SNOMEDCT_US|ESSENTIAL HYPERTENSION, BENIGN|BENIGN ESSENTIAL HYPERTENSION
C0333301|T047|15614009|SNOMEDCT_US|HYPERTENSIVE ISCHEMIC ULCER -RETIRED-|HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|HYPERTENSIVE ISCHAEMIC ULCER -RETIRED-|HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|HYPERTENSIVE ISCHEMIC ULCER|HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|HYPERTENSIVE ISCHAEMIC ULCER|HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|HYPERTENSIVE ISCHEMIC ULCER |HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|ULCER OF SKIN CAUSED BY ISCHEMIA DUE TO HYPERTENSION|HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|ULCER OF SKIN CAUSED BY ISCHAEMIA DUE TO HYPERTENSION|HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|ULCER OF SKIN CAUSED BY ISCHAEMIA DUE TO HYPERTENSIVE DISEASE|HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|ULCER OF SKIN CAUSED BY ISCHEMIA DUE TO HYPERTENSIVE DISEASE |HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|ULCER OF SKIN CAUSED BY ISCHEMIA DUE TO HYPERTENSIVE DISEASE|HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0333301|T047|15614009|SNOMEDCT_US|ULCER OF SKIN CAUSED BY ISCHEMIA DUE TO HYPERTENSIVE DISEASE. DL |HYPERTENSIVE ISCHEMIC ULCER (DISORDER)
C0340272|T047|194793008|SNOMEDCT_US|OTHER SPECIFIED HYPERTENSIVE DISEASE|OTHER SPECIFIED HYPERTENSIVE DISEASE (DISORDER)
C0340272|T047|194793008|SNOMEDCT_US|OTHER SPECIFIED HYPERTENSIVE DISEASE |OTHER SPECIFIED HYPERTENSIVE DISEASE (DISORDER)
C1301626|T047|397748008|SNOMEDCT_US|HYPERTENSION WITH ALBUMINURIA|HYPERTENSION WITH ALBUMINURIA (DISORDER)
C1301626|T047|397748008|SNOMEDCT_US|HYPERTENSION WITH ALBUMINURIA |HYPERTENSION WITH ALBUMINURIA (DISORDER)
C1301626|T047|397748008|SNOMEDCT_US|HYPERTENSION WITH ALBUMINURIA |HYPERTENSION WITH ALBUMINURIA (DISORDER)
C0264637|T047|10725009|SNOMEDCT_US|BENIGN HYPERTENSION |BENIGN HYPERTENSION
C0264637|T047|10725009|SNOMEDCT_US|HYPERTENSION;BENIGN|BENIGN HYPERTENSION
C0264637|T047|10725009|SNOMEDCT_US|BENIGN HYPERTENSION|BENIGN HYPERTENSION
C0264637|T047|10725009|SNOMEDCT_US|BENIGN HYPERTENSION |BENIGN HYPERTENSION
C0264637|T047|10725009|SNOMEDCT_US|BENIGN; HYPERTENSION|BENIGN HYPERTENSION
C0264637|T047|10725009|SNOMEDCT_US|HYPERTENSION; BENIGN|BENIGN HYPERTENSION
C0235222|T047|48146000|SNOMEDCT_US|DIASTOLIC HYPERTENSION|DIASTOLIC HYPERTENSION (DISORDER)
C0235222|T047|48146000|SNOMEDCT_US|DIASTOLIC HYPERTENSION |DIASTOLIC HYPERTENSION (DISORDER)
C0235222|T047|48146000|SNOMEDCT_US|HYPERTENION DIASTOLIC|DIASTOLIC HYPERTENSION (DISORDER)
C0235222|T047|48146000|SNOMEDCT_US|HYPERTENSION DIASTOLIC|DIASTOLIC HYPERTENSION (DISORDER)
C0235222|T047|48146000|SNOMEDCT_US|DIASTOLIC HYPERTENSION |DIASTOLIC HYPERTENSION (DISORDER)
C0235222|T047|48146000|SNOMEDCT_US|DIASTOLIC HYPERTENSION, NOS|DIASTOLIC HYPERTENSION (DISORDER)
C0520539|T047|62275004|SNOMEDCT_US|HYPERTENSIVE EPISODES|HYPERTENSIVE EPISODE (DISORDER)
C1997276|T047|429198000|SNOMEDCT_US|EXERTIONAL HYPERTENSION|EXERTIONAL HYPERTENSION (DISORDER)
C1997276|T047|429198000|SNOMEDCT_US|EXERTIONAL HYPERTENSION |EXERTIONAL HYPERTENSION (DISORDER)
C1997276|T047|429198000|SNOMEDCT_US|EXERTIONAL HYPERTENSION |EXERTIONAL HYPERTENSION (DISORDER)
C0221155|T047|56218007|SNOMEDCT_US|SYSTOLIC HYPERTENSION|SYSTOLIC HYPERTENSION (DISORDER)
C0221155|T047|56218007|SNOMEDCT_US|SYSTOLIC HYPERTENSION |SYSTOLIC HYPERTENSION (DISORDER)
C0221155|T047|56218007|SNOMEDCT_US|SYSTOLIC HYPERTENSION |SYSTOLIC HYPERTENSION (DISORDER)
C0221155|T047|56218007|SNOMEDCT_US|HYPERTENSION SYSTOLIC|SYSTOLIC HYPERTENSION (DISORDER)
C0520540|T047|84094009|SNOMEDCT_US|REBOUND HYPERTENSION |REBOUND HYPERTENSION (DISORDER)
C0520540|T047|84094009|SNOMEDCT_US|REBOUND HYPERTENSION|REBOUND HYPERTENSION (DISORDER)
C0520540|T047|84094009|SNOMEDCT_US|HYPERTENSION REBOUND|REBOUND HYPERTENSION (DISORDER)
C0520540|T047|84094009|SNOMEDCT_US|REBOUND HYPERTENSION |REBOUND HYPERTENSION (DISORDER)
C3669043|T047|697929007|SNOMEDCT_US|INTERMITTENT HYPERTENSION |INTERMITTENT HYPERTENSION
C3669043|T047|697929007|SNOMEDCT_US|INTERMITTENT HYPERTENSION|INTERMITTENT HYPERTENSION
C1862170|T047|720568003|SNOMEDCT_US|HYPERTENSION WITH BRACHYDACTYLY|BRACHYDACTYLY TYPE E WITH SHORT STATURE AND HYPERTENSION
C1862170|T047|720568003|SNOMEDCT_US|BRACHYDACTYLY TYPE E WITH SHORT STATURE AND HYPERTENSION|BRACHYDACTYLY TYPE E WITH SHORT STATURE AND HYPERTENSION
C1862170|T047|720568003|SNOMEDCT_US|BRACHYDACTYLY WITH HYPERTENSION|BRACHYDACTYLY TYPE E WITH SHORT STATURE AND HYPERTENSION
C1862170|T047|720568003|SNOMEDCT_US|BRACHYDACTYLY, TYPE E, WITH SHORT STATURE AND HYPERTENSION|BRACHYDACTYLY TYPE E WITH SHORT STATURE AND HYPERTENSION
C1862170|T047|720568003|SNOMEDCT_US|HTNB|BRACHYDACTYLY TYPE E WITH SHORT STATURE AND HYPERTENSION
C1837739|T047||SNOMEDCT_US|HYPERTENSION, DIASTOLIC, RESISTANCE TO
C1839021|T047||SNOMEDCT_US|HYPOMAGNESEMIA, HYPERTENSION, AND HYPERCHOLESTEROLEMIA, MITOCHONDRIAL
C1839021|T047||SNOMEDCT_US|HYPERTENSION, HYPERCHOLESTEROLEMIA, AND HYPOMAGNESEMIA, MITOCHONDRIAL
C1833688|T047||SNOMEDCT_US|OSTEOCHONDRODYSPLASIA, RHIZOMELIC, WITH CALLOSAL AGENESIS, THROMBOCYTOPENIA, HYDROCEPHALUS, AND HYPERTENSION
C3501739|T047||SNOMEDCT_US|TACHYCARDIA, HYPERTENSION, MICROPHTHALMIA, AND HYPERGLYCINURIA
C1854631|T047||SNOMEDCT_US|HYPERTENSION, EARLY-ONSET, AUTOSOMAL DOMINANT, WITH SEVERE EXACERBATION IN PREGNANCY
C1834155|T047||SNOMEDCT_US|HYPERTENSION, RESISTANT TO CONVENTIONAL THERAPY
C1834155|T047||SNOMEDCT_US|HYPERTENSION RESISTANT TO CONVENTIONAL THERAPY
C1865267|T047|717824007|SNOMEDCT_US|ARTERIAL OCCLUSIVE DISEASE, PROGRESSIVE, WITH HYPERTENSION, HEART DEFECTS, BONE FRAGILITY, AND BRACHYSYNDACTYLY|GRANGE OCCLUSIVE ARTERIAL SYNDROME
C1865267|T047|717824007|SNOMEDCT_US|GRANGE OCCLUSIVE ARTERIAL SYNDROME|GRANGE OCCLUSIVE ARTERIAL SYNDROME
C3831106|T047||SNOMEDCT_US|CHRONIC MATERNAL HYPERTENSION WITH SUPERIMPOSED PREECLAMPSIA
C3827254|T047||SNOMEDCT_US|CHRONIC MATERNAL HYPERTENSION
C3837203|T047||SNOMEDCT_US|HYPERTENSION (SYSTEMIC) SUSCEPTIBILITY
C3837203|T047||SNOMEDCT_US|HYPERTENSION (SYSTEMIC) SUSCEPTIBILITY 
C3874846|T047|71421000119105|SNOMEDCT_US|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE 2 DIABETES MELLITUS |HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE 2 DIABETES MELLITUS (DISORDER)
C3874846|T047|71421000119105|SNOMEDCT_US|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE II DIABETES MELLITUS|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE 2 DIABETES MELLITUS (DISORDER)
C3874846|T047|71421000119105|SNOMEDCT_US|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE 2 DIABETES MELLITUS|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE 2 DIABETES MELLITUS (DISORDER)
C3874779|T047|71701000119105|SNOMEDCT_US|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE 1 DIABETES MELLITUS |HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE I DIABETES MELLITUS
C3874779|T047|71701000119105|SNOMEDCT_US|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE I DIABETES MELLITUS|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE I DIABETES MELLITUS
C3874779|T047|71701000119105|SNOMEDCT_US|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE 1 DIABETES MELLITUS|HYPERTENSION IN CHRONIC KIDNEY DISEASE DUE TO TYPE I DIABETES MELLITUS
C0020546|T047|706882009|SNOMEDCT_US|HYPERTENSIVE CRISIS|HYPERTENSIVE CRISIS (DISORDER)
C0020546|T047|706882009|SNOMEDCT_US|HYPERTENSIVE CRISIS |HYPERTENSIVE CRISIS (DISORDER)
C0020546|T047|706882009|SNOMEDCT_US|CRISIS HYPERTENSIVE|HYPERTENSIVE CRISIS (DISORDER)
C2902961|T047|367821000119106|SNOMEDCT_US|PAGE KIDNEY|HYPERTENSION DUE TO COMPRESSION OF RENAL PARENCHYMA
C2902961|T047|367821000119106|SNOMEDCT_US|PAGE KIDNEY |HYPERTENSION DUE TO COMPRESSION OF RENAL PARENCHYMA
C2902961|T047|367821000119106|SNOMEDCT_US|HYPERTENSION DUE TO COMPRESSION OF RENAL PARENCHYMA|HYPERTENSION DUE TO COMPRESSION OF RENAL PARENCHYMA
C2902961|T047|367821000119106|SNOMEDCT_US|HYPERTENSION DUE TO COMPRESSION OF RENAL PARENCHYMA |HYPERTENSION DUE TO COMPRESSION OF RENAL PARENCHYMA
C1857175|T047||SNOMEDCT_US|HYPERTENSION, EPISODIC
C1857175|T047||SNOMEDCT_US|EPISODIC HYPERTENSION
C4025693|T047||SNOMEDCT_US|HYPERTENSION ASSOCIATED WITH PHEOCHROMOCYTOMA
C0020545|T047|194790006|SNOMEDCT_US|HYPERTENSION, RENOVASCULAR|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|RENOVASCULAR HYPERTENSION|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|RENOVASCULAR HYPERTENSION |SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|SECONDARY HYPERTENSION RENOVASCULAR|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|HYPERTENSION, RENOVASCULAR [DISEASE/FINDING]|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|SECONDARY RENOVASCULAR HYPERTENSION NOS|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|SECONDARY RENOVASCULAR HYPERTENSION NOS |SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|HYPERTENSION DUE TO RENAL ARTERY HYPERPLASIA|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|HYPERTENSION DUE TO RENOVASCULAR DISEASE|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|RENOVASCULAR HYPERTENSION |SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|HYPERTENSION; RENOVASCULAR DISORDERS|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|HYPERTENSION; RENOVASCULAR|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|RENAL DISEASE; HYPERTENSION, ARTERIAL|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C0020545|T047|194790006|SNOMEDCT_US|RENOVASCULAR; HYPERTENSION|SECONDARY RENOVASCULAR HYPERTENSION NOS (DISORDER)
C4076686|T047|712832005|SNOMEDCT_US|SUPINE HYPERTENSION|SUPINE HYPERTENSION (DISORDER)
C4076686|T047|712832005|SNOMEDCT_US|SUPINE HYPERTENSION |SUPINE HYPERTENSION (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|HYPERTENSIVE ENCEPHALOPATHY|HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|HYPERTENSIVE ENCEPH|HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|ENCEPH HYPERTENSIVE|HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|HYPERTENSIVE ENCEPHALOPATHY |HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|HYPERTENS ENCEPHALOPATHY|HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|ENCEPHALOPATHY, HYPERTENSIVE|HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|HYPERTENSIVE ENCEPHALOPATHY [DISEASE/FINDING]|HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|HYPERTENSIVE ENCEPHALOPATHY |HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|ENCEPHALOPATHY HYPERTENSIVE|HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0151620|T047|50490005|SNOMEDCT_US|ENCEPHALOPATHY; HYPERTENSIVE|HYPERTENSIVE ENCEPHALOPATHY (DISORDER)
C0494575|T047|194779001|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE, UNSPECIFIED, WITH CONGESTIVE HEART FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH (CONGESTIVE) HEART FAILURE (DISORDER)
C0494575|T047|194779001|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH (CONGESTIVE) HEART FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH (CONGESTIVE) HEART FAILURE (DISORDER)
C0494575|T047|194779001|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH (CONGESTIVE) HEART FAILURE |HYPERTENSIVE HEART AND RENAL DISEASE WITH (CONGESTIVE) HEART FAILURE (DISORDER)
C0494575|T047|194779001|SNOMEDCT_US|FAILURE; CARDIORENAL, HYPERTENSIVE, WITH HEART FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH (CONGESTIVE) HEART FAILURE (DISORDER)
C0264650|T047|5148006|SNOMEDCT_US|UNSPECIFIED HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE|HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE (DISORDER)
C0264650|T047|5148006|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE WITH (CONGESTIVE) HEART FAILURE|HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE (DISORDER)
C0264650|T047|5148006|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE NOS WITH CONGESTIVE CARDIAC FAILURE |HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE (DISORDER)
C0264650|T047|5148006|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE NOS WITH CONGESTIVE CARDIAC FAILURE|HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE (DISORDER)
C0264650|T047|5148006|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE|HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE (DISORDER)
C0264650|T047|5148006|SNOMEDCT_US|HYPERTENSIVE HEART DIS WITH CONGESTIVE HEART FAILURE|HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE (DISORDER)
C0264650|T047|5148006|SNOMEDCT_US|HYPERTENSIVE HEART DIS WITH CONGESTIVE HEART FAILURE |HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE (DISORDER)
C0264650|T047|5148006|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE |HYPERTENSIVE HEART DISEASE WITH CONGESTIVE HEART FAILURE (DISORDER)
C0494574|T047||SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE WITHOUT RENAL FAILURE
C0494574|T047||SNOMEDCT_US|HY KID NOS W CR KID I-IV
C0494574|T047||SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE, UNSPECIFIED, WITHOUT MENTION OF RENAL FAILURE
C0494574|T047||SNOMEDCT_US|HYPERTENSIVE CHRONIC KIDNEY DISEASE, UNSPECIFIED, WITH CHRONIC KIDNEY DISEASE STAGE I THROUGH STAGE IV, OR UNSPECIFIED
C0348586|T047|195538006|SNOMEDCT_US|OTHER UNSPECIFIED SECONDARY HYPERTENSION|[X]OTHER SECONDARY HYPERTENSION (DISORDER)
C0348586|T047|195538006|SNOMEDCT_US|OTHER SECONDARY HYPERTENSION|[X]OTHER SECONDARY HYPERTENSION (DISORDER)
C0348586|T047|195538006|SNOMEDCT_US|SECOND HYPERTENSION NEC|[X]OTHER SECONDARY HYPERTENSION (DISORDER)
C0348586|T047|195538006|SNOMEDCT_US|[X]OTHER SECONDARY HYPERTENSION|[X]OTHER SECONDARY HYPERTENSION (DISORDER)
C0348586|T047|195538006|SNOMEDCT_US|[X]OTHER SECONDARY HYPERTENSION |[X]OTHER SECONDARY HYPERTENSION (DISORDER)
C0155591|T047|60899001|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE WITHOUT (CONGESTIVE) HEART FAILURE|HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE (DISORDER)
C0155591|T047|60899001|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE NOS WITHOUT CONGESTIVE CARDIAC FAILURE|HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE (DISORDER)
C0155591|T047|60899001|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE NOS WITHOUT CONGESTIVE CARDIAC FAILURE |HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE (DISORDER)
C0155591|T047|60899001|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE|HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE (DISORDER)
C0155591|T047|60899001|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE |HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE (DISORDER)
C0155591|T047|60899001|SNOMEDCT_US|UNSPECIFIED HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE|HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE (DISORDER)
C0155591|T047|60899001|SNOMEDCT_US|HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE |HYPERTENSIVE HEART DISEASE WITHOUT CONGESTIVE HEART FAILURE (DISORDER)
C0155620|T047|194785008|SNOMEDCT_US|SECONDARY BENIGN HYPERTENSION|SECONDARY BENIGN HYPERTENSION (DISORDER)
C0155620|T047|194785008|SNOMEDCT_US|BENIGN SECONDARY HYPERTENSION |SECONDARY BENIGN HYPERTENSION (DISORDER)
C0155620|T047|194785008|SNOMEDCT_US|BENIGN SECONDARY HYPERTENSION|SECONDARY BENIGN HYPERTENSION (DISORDER)
C0155620|T047|194785008|SNOMEDCT_US|SECONDARY HYPERTENSION BENIGN|SECONDARY BENIGN HYPERTENSION (DISORDER)
C0155620|T047|194785008|SNOMEDCT_US|SECONDARY BENIGN HYPERTENSION NOS|SECONDARY BENIGN HYPERTENSION (DISORDER)
C0155620|T047|194785008|SNOMEDCT_US|SECONDARY BENIGN HYPERTENSION NOS |SECONDARY BENIGN HYPERTENSION (DISORDER)
C0155620|T047|194785008|SNOMEDCT_US|BENIGN SECONDARY HYPERTENSION |SECONDARY BENIGN HYPERTENSION (DISORDER)
C0155620|T047|194785008|SNOMEDCT_US|SECONDARY HYPERTENSION, BENIGN|SECONDARY BENIGN HYPERTENSION (DISORDER)
C0155620|T047|194785008|SNOMEDCT_US|SECONDARY BENIGN HYPERTENSION |SECONDARY BENIGN HYPERTENSION (DISORDER)
C0544618|T047||SNOMEDCT_US|ORTHOSTATIC HYPERTENSION
C1171328|T047||SNOMEDCT_US|CATECHOLAMINE HYPERTENSION
C0597290|T047||SNOMEDCT_US|PROSTAGLANDIN HYPERTENSION
C0155622|T047||SNOMEDCT_US|OTHER BENIGN SECONDARY HYPERTENSION
C0155622|T047||SNOMEDCT_US|BENIGN SECOND HYPERT NEC
C0221154|T047|23130000|SNOMEDCT_US|PAROXYSMAL HYPERTENSION (PHYSICAL FINDING)|EPISODIC HYPERTENSION
C0221154|T047|23130000|SNOMEDCT_US|PAROXYSMAL HYPERTENSION|EPISODIC HYPERTENSION
C0221154|T047|23130000|SNOMEDCT_US|PAROXYSMAL HYPERTENSION WAS OBSERVED|EPISODIC HYPERTENSION
C0221154|T047|23130000|SNOMEDCT_US|HYPERTENSION PAROXYSMAL|EPISODIC HYPERTENSION
C0221154|T047|23130000|SNOMEDCT_US|PAROXYSMAL HYPERTENSION |EPISODIC HYPERTENSION
C0341909|T047|199013004|SNOMEDCT_US|HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH, AND THE PUERPERIUM|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C0341909|T047|199013004|SNOMEDCT_US|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM NOS|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C0341909|T047|199013004|SNOMEDCT_US|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED |UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C0341909|T047|199013004|SNOMEDCT_US|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C0341909|T047|199013004|SNOMEDCT_US|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM |UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C0341909|T047|199013004|SNOMEDCT_US|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM NOS |UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C0341909|T047|199013004|SNOMEDCT_US|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C0341909|T047|199013004|SNOMEDCT_US|HYPERTENSION COMPLICATING PREGNANCY; CHILDBIRTH AND THE PUERPERIUM|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C0341909|T047|199013004|SNOMEDCT_US|HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C0341909|T047|199013004|SNOMEDCT_US|HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM |UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH AND THE PUERPERIUM UNSPECIFIED (DISORDER)
C1171326|T047||SNOMEDCT_US|BRADYKININ HYPERTENSION
C1171351|T047||SNOMEDCT_US|KININ HYPERTENSION
C0349368|T047|194788005|SNOMEDCT_US|HYPERTENSION SECONDARY TO ENDOCRINE DISORDERS|HYPERTENSION SECONDARY TO ENDOCRINE DISORDER (DISORDER)
C0349368|T047|194788005|SNOMEDCT_US|HYPERTENSION SECONDARY TO ENDOCRINE DISORDERS |HYPERTENSION SECONDARY TO ENDOCRINE DISORDER (DISORDER)
C0349368|T047|194788005|SNOMEDCT_US|SECONDARY HYPERTENSION TO ENDOCRINE DISORDERS|HYPERTENSION SECONDARY TO ENDOCRINE DISORDER (DISORDER)
C0349368|T047|194788005|SNOMEDCT_US|HYPERTENSION; SECONDARY, DUE TO ENDOCRINE DISORDERS|HYPERTENSION SECONDARY TO ENDOCRINE DISORDER (DISORDER)
C0349368|T047|194788005|SNOMEDCT_US|SECONDARY; HYPERTENSION, DUE TO ENDOCRINE DISORDERS|HYPERTENSION SECONDARY TO ENDOCRINE DISORDER (DISORDER)
C0349368|T047|194788005|SNOMEDCT_US|HYPERTENSION SECONDARY TO ENDOCRINE DISORDER |HYPERTENSION SECONDARY TO ENDOCRINE DISORDER (DISORDER)
C0349368|T047|194788005|SNOMEDCT_US|HYPERTENSION SECONDARY TO ENDOCRINE DISORDER|HYPERTENSION SECONDARY TO ENDOCRINE DISORDER (DISORDER)
C0349368|T047|194788005|SNOMEDCT_US|HYPERTENSION SECONDARY TO ENDOCRINE DISORDERS |HYPERTENSION SECONDARY TO ENDOCRINE DISORDER (DISORDER)
C0348587|T047|195539003|SNOMEDCT_US|HYPERTENSION SECONDARY TO OTHER RENAL DISORDERS|[X]HYPERTENSION SECONDARY TO OTHER RENAL DISORDERS (DISORDER)
C0348587|T047|195539003|SNOMEDCT_US|[X]HYPERTENSION SECONDARY TO OTHER RENAL DISORDERS |[X]HYPERTENSION SECONDARY TO OTHER RENAL DISORDERS (DISORDER)
C0348587|T047|195539003|SNOMEDCT_US|[X]HYPERTENSION SECONDARY TO OTHER RENAL DISORDERS|[X]HYPERTENSION SECONDARY TO OTHER RENAL DISORDERS (DISORDER)
C0348587|T047|195539003|SNOMEDCT_US|HYPERTENSION; SECONDARY, DUE TO RENAL DISORDERS|[X]HYPERTENSION SECONDARY TO OTHER RENAL DISORDERS (DISORDER)
C0348587|T047|195539003|SNOMEDCT_US|SECONDARY; HYPERTENSION, DUE TO RENAL DISORDERS|[X]HYPERTENSION SECONDARY TO OTHER RENAL DISORDERS (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE, UNSPECIFIED, WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYP KID NOS W CR KID V|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE CHRONIC KIDNEY DISEASE, UNSPECIFIED, WITH CHRONIC KIDNEY DISEASE STAGE V OR END STAGE RENAL DISEASE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE KIDNEY DISEASE WITH RENAL FAILURE |HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE KIDNEY DISEASE WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE |HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|HYPERTENSION; RENAL DISEASE, HYPERTENSIVE, WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|INSUFFICIENCY; RENAL, CHRONIC, HYPERTENSIVE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|INSUFFICIENCY; RENAL, WITH HYPERTENSION|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348860|T047|194774006|SNOMEDCT_US|KIDNEY; HYPERTENSION, WITH RENAL FAILURE|HYPERTENSIVE RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE, UNSPECIFIED, WITH RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE |HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE WITH RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HY HT/KD NOS ST V W/O HF|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE, UNSPECIFIED, WITHOUT HEART FAILURE AND WITH CHRONIC KIDNEY DISEASE STAGE V OR END STAGE RENAL DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE |HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|FAILURE; CARDIORENAL, HYPERTENSIVE, WITH RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|INSUFFICIENCY; RENAL, WITH HYPERTENSIVE HEART DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0348879|T047|194780003|SNOMEDCT_US|KIDNEY; INSUFFICIENCY, WITH HYPERTENSIVE HEART DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE WITH RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE, UNSPECIFIED, WITH CONGESTIVE HEART FAILURE AND RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYP HT/KD NOS ST V W HF|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND CHRONIC KIDNEY DISEASE, UNSPECIFIED, WITH HEART FAILURE AND CHRONIC KIDNEY DISEASE STAGE V OR END STAGE RENAL DISEASE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE, UNSPECIFIED, WITH HEART FAILURE AND RENAL FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE |HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|INSUFFICIENCY; RENAL, WITH HYPERTENSIVE HEART DISEASE AND HEART FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0494576|T047|194781004|SNOMEDCT_US|KIDNEY; INSUFFICIENCY, WITH HYPERTENSIVE HEART DISEASE AND HEART FAILURE|HYPERTENSIVE HEART AND RENAL DISEASE WITH BOTH (CONGESTIVE) HEART FAILURE AND RENAL FAILURE (DISORDER)
C0269660|T047|69909000|SNOMEDCT_US|ECLAMPSIA ADDED TO PRE-EXISTING HYPERTENSION|ECLAMPSIA ADDED TO PRE-EXISTING HYPERTENSION (DISORDER)
C0269660|T047|69909000|SNOMEDCT_US|ECLAMPSIA ADDED TO PRE-EXISTING HYPERTENSION |ECLAMPSIA ADDED TO PRE-EXISTING HYPERTENSION (DISORDER)
C0156689|T047||SNOMEDCT_US|HYPERTENS NOS-ANTEPARTUM
C0156689|T047||SNOMEDCT_US|UNSPECIFIED HYPERTENSION COMPLICATING PREGNANCY, CHILDBIRTH, OR THE PUERPERIUM, ANTEPARTUM CONDITION OR COMPLICATION
C0156689|T047||SNOMEDCT_US|UNSPECIFIED ANTEPARTUM HYPERTENSION
C0497248|T047||SNOMEDCT_US|HYPERTENSION;UNCOMPLICATED
C0497248|T047||SNOMEDCT_US|UNCOMPLICATED HYPERTENSION
C1335457|T047||SNOMEDCT_US|POSTPARTUM HYPERTENSION
C0028840|T047|4210003|SNOMEDCT_US|HYPERTENSIONS, OCULAR|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|OCULAR HYPERTENSION|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|OCULAR HYPERTENSIONS|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|PREGLAUCOMA OCULAR HYPERTENSION |OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|PREGLAUCOMA OCULAR HYPERTENSION|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|HYPERTENSION, OCULAR|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|OCULAR HYPERTENSION [DISEASE/FINDING]|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|HYPERTENSION OCULAR|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|OH - OCULAR HYPERTENSION|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|OHT - OCULAR HYPERTENSION|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|OCULAR HYPERTENSION |OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|HYPERTENSION; OCULAR|OCULAR HYPERTENSION (DISORDER)
C0028840|T047|4210003|SNOMEDCT_US|OCULAR; HYPERTENSION|OCULAR HYPERTENSION (DISORDER)
C2227904|T047||SNOMEDCT_US|AMERICAN COLLEGE OF PHYSICIANS (ACP) STAGING STAGE 1 HYPERTENSION: 140-159/90-99 (PHYSICAL FINDING)
C2227904|T047||SNOMEDCT_US|AMERICAN COLLEGE OF PHYSICIANS (ACP) STAGING STAGE 1 HYPERTENSION: 140-159/90-99
C2227904|T047||SNOMEDCT_US|ACP STAGING STAGE 1 HYPERTENSION: 140-159 / 90-99
C2227905|T047||SNOMEDCT_US|AMERICAN COLLEGE OF PHYSICIANS (ACP) STAGING STAGE 2 HYPERTENSION: GREATER THAN EQUAL TO 160/100
C2227905|T047||SNOMEDCT_US|AMERICAN COLLEGE OF PHYSICIANS (ACP) STAGING STAGE 2 HYPERTENSION: GREATER THAN EQUAL TO 160/100 (PHYSICAL FINDING)
C2227905|T047||SNOMEDCT_US|ACP STAGING STAGE 2 HYPERTENSION: GREATER THAN OR = 160/100
C1556272|T047||SNOMEDCT_US|CTCAE GRADE 1 HYPERTENSION
C1556272|T047||SNOMEDCT_US|GRADE 1 HYPERTENSION
C1556275|T047||SNOMEDCT_US|CTCAE GRADE 4 HYPERTENSION
C1556275|T047||SNOMEDCT_US|GRADE 4 HYPERTENSION
C1556276|T047||SNOMEDCT_US|CTCAE GRADE 5 HYPERTENSION
C1556276|T047||SNOMEDCT_US|GRADE 5 HYPERTENSION
C1556274|T047||SNOMEDCT_US|CTCAE GRADE 3 HYPERTENSION
C1556274|T047||SNOMEDCT_US|GRADE 3 HYPERTENSION
C1556273|T047||SNOMEDCT_US|CTCAE GRADE 2 HYPERTENSION
C1556273|T047||SNOMEDCT_US|GRADE 2 HYPERTENSION
