C0474232|T129||CVX|PATIENT IMMUNE TO HEPATITIS B
C0474232|T129||CVX|PATIENT IMMUNE TO HEP B
C0474232|T129||CVX|PATIENT VACCINATED FOR HEP B
C0474232|T129||CVX|HEPATITIS B VACCINATION (SNOMED:16584000)
C2716397|T129|146|CVX|DIPHTHERIA AND TETANUS TOXOIDS AND ACELLULAR PERTUSSIS ADSORBED, INACTIVATED POLIOVIRUS, HAEMOPHILUS B CONJUGATE (MENINGOCOCCAL PROTEIN CONJUGATE), AND HEPATITIS B (RECOMBINANT) VACCINE.|DTAP,IPV,HIB,HEPB
C2716397|T129|146|CVX|DTAP,IPV,HIB,HEPB|DTAP,IPV,HIB,HEPB
C3644155|T129||CVX|DTAP-HEP B-IPV
C3644155|T129||CVX|DTAP-HEPATITIS B AND POLIOVIRUS VACCINE
C3644182|T129|132|CVX|DTAP-IPV-HIB-HEP B, HISTORICAL|DTAP-IPV-HIB-HEP B, HISTORICAL
C1548467|T129|102|CVX|DTAP/DTP-HIB-HEP B|DTP-HIB-HEP B
C1548467|T129|102|CVX|DTP- HAEMOPHILUS INFLUENZAE TYPE B CONJUGATE AND HEPATITIS B VACCINE|DTP-HIB-HEP B
C0694743|T129||CVX|HAEMOPHILUS INFLUENZAE TYPE B CONJUGATE AND HEPATITIS B VACCINE
C3644158|T129||CVX|HEP B, UNSPECIFIED FORMULATION
C1552908|T129|42|CVX|HEPATITIS B VACCINE, ADOLESCENT/HIGH RISK INFANT DOSAGE|HEP B, ADOLESCENT/HIGH RISK INFANT
C1552909|T129|43|CVX|HEPATITIS B VACCINE, ADULT DOSAGE|HEP B, ADULT
C0694736|T129|44|CVX|HEPATITIS B VACCINE, DIALYSIS PATIENT DOSAGE|HEP B, DIALYSIS
C0694733|T129|08|CVX|HEPATITIS B VACCINE, PEDIATRIC OR PEDIATRIC/ADOLESCENT DOSAGE|HEP B, ADOLESCENT OR PEDIATRIC
C3644158|T129||CVX|HEPATITIS B VACCINE, UNSPECIFIED FORMULATION
C0694743|T129||CVX|HIB-HEP B
C3644182|T129|132|CVX|HISTORICAL RECORD OF VACCINE CONTAINING * DIPHTHERIA, TETANUS TOXOIDS AND ACELLULAR PERTUSSIS, * POLIOVIRUS, INACTIVATED, * HAEMOPHILUS INFLUENZAE TYPE B CONJUGATE, * HEPATITIS B|DTAP-IPV-HIB-HEP B, HISTORICAL
C1170008|T129||CVX|HEP A-HEP B
C0730242|T129||CVX|COMBINED HEPATITIS A & HEPATITIS B VACCINATION
C0730242|T129||CVX|COMBINED HEPATITIS A AND HEPATITIS B VACCINATION 
C0730242|T129||CVX|COMBINED HEPATITIS A AND HEPATITIS B VACCINATION
C0730242|T129||CVX|COMBINED HEPATITIS A AND B VACCINATION
C0730242|T129||CVX|COMBINED HEPATITIS A AND B VACCINATION 
C1300747|T129||CVX|VACC COMB BACT & VIRAL ADMINISTERED DIPHTH - ACELL PERTUS - HEPB - IPV
C1300747|T129||CVX|DIPHTHERIA-ACELLULAR PERTUSSIS-HEPB-IPV VACCINATION
C1300747|T129||CVX|DIPHTHERIA-ACELLULAR PERTUSSIS-HEPB-IPV VACCINATION 
C1300747|T129||CVX|DIPHTHERIA, ACELLULAR PERTUSSIS, HEPATITIS B AND INACTIVATED POLIO VACCINATION 
C1300747|T129||CVX|DIPHTHERIA, ACELLULAR PERTUSSIS, HEPATITIS B AND INACTIVATED POLIO VACCINATION
C0474232|T129||CVX|HEPATITIS B IMMUNISATION
C0474232|T129||CVX|IMMUNISATION;HEPATITIS B
C0474232|T129||CVX|HEPATITIS B IMMUNIZATION
C0474232|T129||CVX|HEPATITIS B VACCINE (ACTIVE) ADMINISTRATION
C0474232|T129||CVX|HEPATITIS B VACCINE ADMINISTRATION 
C0474232|T129||CVX|HEPATITIS B VACCINE ADMINISTRATION
C0474232|T129||CVX|ADMINISTRATION OF HEPATITIS B VACCINE
C0474232|T129||CVX|HEP B VACCINATION
C0474232|T129||CVX|HEPATITIS B SERIES IMMUNIZATION
C0474232|T129||CVX|HEPATITIS B VACCINATION
C0474232|T129||CVX|HEPATITIS B INJECTION
C0474232|T129||CVX|HEPATITIS B SERIES IMMUNISATION
C0474232|T129||CVX|HEPATITIS B VACCINATION 
C0474232|T129||CVX|ADMIN HEPATITIS B VACCINE
C0474232|T129||CVX|IMMUNIZATION;HEPATITIS B
C0419731|T129||CVX|BOOSTER HEPATITIS B VACCINATION 
C0419731|T129||CVX|BOOSTER HEPATITIS B VACCINATION
C0419731|T129||CVX|HEPATITIS B VACCINE (ACTIVE) BOOSTER VACCINATION 
C0419731|T129||CVX|HEPATITIS B VACCINE (ACTIVE) BOOSTER VACCINATION
C0419729|T129||CVX|FOURTH HEPATITIS B VACCINATION 
C0419729|T129||CVX|FOURTH HEPATITIS B VACCINATION
C0419729|T129||CVX|HEPATITIS B VACCINE (ACTIVE) FOURTH VACCINATION
C0419729|T129||CVX|HEPATITIS B VACCINE (ACTIVE) FOURTH VACCINATION 
C0419729|T129||CVX|4TH HEPATITIS B VACCINATION
C0419727|T129||CVX|SECOND HEPATITIS B VACCINATION 
C0419727|T129||CVX|SECOND HEPATITIS B VACCINATION
C0419727|T129||CVX|HEPATITIS B VACCINE (ACTIVE) SECOND VACCINATION
C0419727|T129||CVX|HEPATITIS B VACCINE (ACTIVE) SECOND VACCINATION 
C0419727|T129||CVX|2ND HEPATITIS B VACCINATION
C0419728|T129||CVX|THIRD HEPATITIS B VACCINATION 
C0419728|T129||CVX|THIRD HEPATITIS B VACCINATION
C0419728|T129||CVX|HEPATITIS B VACCINE (ACTIVE) THIRD VACCINATION
C0419728|T129||CVX|HEPATITIS B VACCINE (ACTIVE) THIRD VACCINATION 
C0419728|T129||CVX|3RD HEPATITIS B VACCINATION
C0419726|T129||CVX|FIRST HEPATITIS B VACCINATION
C0419726|T129||CVX|FIRST HEPATITIS B VACCINATION 
C0419726|T129||CVX|HEPATITIS B VACCINE (ACTIVE) FIRST VACCINATION
C0419726|T129||CVX|HEPATITIS B VACCINE (ACTIVE) FIRST VACCINATION 
C0419726|T129||CVX|1ST HEPATITIS B VACCINATION
C0419730|T129||CVX|FIFTH HEPATITIS B VACCINATION
C0419730|T129||CVX|FIFTH HEPATITIS B VACCINATION 
C0419730|T129||CVX|5TH HEPATITIS B VACCINATION
C1562257|T129||CVX|SIXTH HEPATITIS B VACCINATION 
C1562257|T129||CVX|SIXTH HEPATITIS B VACCINATION
C3661302|T129||CVX|INFANRIX HEXA
C2716397|T129|146|CVX|DIPHTHERIA-TETANUS-ACELLULAR PERTUSSIS-INACTIVATED POLIOVIRUS-HAEMOPHILUS INFLUENZAE B CONJUGATE-HEPATITIS B VACCINE|DTAP,IPV,HIB,HEPB
C2716397|T129|146|CVX|DTAP-IPV-HIB-HBV VACCINE|DTAP,IPV,HIB,HEPB
C2716397|T129|146|CVX|DTAP-IPV-HIB-HBV CONJUGATE VACCINE|DTAP,IPV,HIB,HEPB
C2716397|T129|146|CVX|DTAP-IPV-HIB-HEPB|DTAP,IPV,HIB,HEPB
C2716397|T129|146|CVX|DTAP-IPV-HIB-HEPB |DTAP,IPV,HIB,HEPB
C2716397|T129|146|CVX|DTAP,IPV,HIB,HEPB|DTAP,IPV,HIB,HEPB
C2716397|T129|146|CVX|DIPHTHERIA AND TETANUS TOXOIDS AND ACELLULAR PERTUSSIS ADSORBED, INACTIVATED POLIOVIRUS, HAEMOPHILUS B CONJUGATE (MENINGOCOCCAL PROTEIN CONJUGATE), AND HEPATITIS B (RECOMBINANT) VACCINE.|DTAP,IPV,HIB,HEPB
C3644155|T129||CVX|DTAP-HEP B-IPV
C3644155|T129||CVX|DTAP-HEPATITIS B AND POLIOVIRUS VACCINE
C3644182|T129|132|CVX|HISTORICAL RECORD OF VACCINE CONTAINING * DIPHTHERIA, TETANUS TOXOIDS AND ACELLULAR PERTUSSIS, * POLIOVIRUS, INACTIVATED, * HAEMOPHILUS INFLUENZAE TYPE B CONJUGATE, * HEPATITIS B|DTAP-IPV-HIB-HEP B, HISTORICAL
C3644182|T129|132|CVX|DTAP-IPV-HIB-HEP B, HISTORICAL|DTAP-IPV-HIB-HEP B, HISTORICAL
C1548467|T129|102|CVX|DTAP/DTP-HIB-HEP B|DTP-HIB-HEP B
C1548467|T129|102|CVX|DTP- HAEMOPHILUS INFLUENZAE TYPE B CONJUGATE AND HEPATITIS B VACCINE|DTP-HIB-HEP B
C1548467|T129|102|CVX|DTP-HIB-HEP B|DTP-HIB-HEP B
C0694743|T129||CVX|HIB-HEP B
C0694743|T129||CVX|HAEMOPHILUS INFLUENZAE TYPE B CONJUGATE AND HEPATITIS B VACCINE
C0694733|T129|08|CVX|HEPATITIS B VACCINE, PEDIATRIC OR PEDIATRIC/ADOLESCENT DOSAGE|HEP B, ADOLESCENT OR PEDIATRIC
C0694733|T129|08|CVX|HEP B, ADOLESCENT OR PEDIATRIC|HEP B, ADOLESCENT OR PEDIATRIC
C1552908|T129|42|CVX|HEPATITIS B VACCINE, ADOLESCENT/HIGH RISK INFANT DOSAGE|HEP B, ADOLESCENT/HIGH RISK INFANT
C1552908|T129|42|CVX|HEP B, ADOLESCENT/HIGH RISK INFANT|HEP B, ADOLESCENT/HIGH RISK INFANT
C1552909|T129|43|CVX|HEPATITIS B VACCINE, ADULT DOSAGE|HEP B, ADULT
C0694736|T129|44|CVX|HEPATITIS B VACCINE, DIALYSIS PATIENT DOSAGE|HEP B, DIALYSIS
C3644158|T129||CVX|HEP B, UNSPECIFIED FORMULATION
C3644158|T129||CVX|HEPATITIS B VACCINE, UNSPECIFIED FORMULATION
C1170689|T129||CVX|TWINRIX JUNIOR
C1170008|T129||CVX|HEPATITIS A AND HEPATITIS B VACCINE
C1170008|T129||CVX|HEP A-HEP B
C1170008|T129||CVX|HEPATITIS A-HEPATITIS B VACCINE
