C0086287|T032||HL7V3.0|FEMALE
C0086287|T032||HL7V3.0|WOMAN
# C0086287|T032||HL7V3.0|COMMON BUT WILL IT GIVE YOU TOO MANY FASLE HITS?
C0086582|T032||HL7V3.0|MALE
C0086582|T032||HL7V3.0|MAN
# C0086582|T032||HL7V3.0|M
# C1550327|T032|ADMINISTRATIVEGENDER|HL7V3.0|ADMINISTRATIVE GENDER|ADMINISTRATIVEGENDER
# C0079399|T032||HL7V3.0|GENDER
# C1522384|T032||HL7V3.0|SEX
C1706180|T032||HL7V3.0|MALE GENDER, SELF REPORT
C1710069|T032||HL7V3.0|SEX OR GENDER
C3839079|T032||HL7V3.0|MASCULINE GENDER
C3839293|T032||HL7V3.0|FEMININE GENDER
C0043210|T032||HL7V3.0|WOMEN
C0043210|T032||HL7V3.0|WOMAN
C0043210|T032||HL7V3.0|WOMAN (PERSON)
C0043210|T032||HL7V3.0|HUMAN, FEMALE
C0025266|T032||HL7V3.0|MAN
C0025266|T032||HL7V3.0|MAN (PERSON)
C0025266|T032||HL7V3.0|HUMAN, MALE
C0086582|T032||HL7V3.0|MALE
# C0086582|T032||HL7V3.0|M
C0086582|T032||HL7V3.0|MALE GENDER
C0086582|T032||HL7V3.0|MALE GENDER [DISEASE/FINDING]
C0086582|T032||HL7V3.0|MALE 
C0086582|T032||HL7V3.0|MALES
C0086582|T032||HL7V3.0|MALE INDIVIDUAL
C0086582|T032||HL7V3.0|MALE INDIVIDUAL, NOS
C0086582|T032||HL7V3.0|MALE, NOS
C0086582|T032||HL7V3.0|HUMAN, MALE
C0432475|T032||HL7V3.0|XX MALE
C0432475|T032||HL7V3.0|MALE WITH 46,XX KARYOTYPE
C0432475|T032||HL7V3.0|MALE WITH 46,XX KARYOTYPE 
C0432475|T032||HL7V3.0|XX MALES
C0432475|T032||HL7V3.0|MALE WITH 46, XX KARYOTYPE
C0432475|T032||HL7V3.0|XX MALES 
C0432475|T032||HL7V3.0|KARYOTYPE; 46,XX, MALE
C1706429|T032||HL7V3.0|MALE
C1706429|T032||HL7V3.0|MALE, SELF-REPORTED
C1706429|T032||HL7V3.0|MALE, SELF-REPORT
C1706429|T032||HL7V3.0|MALE SEX, SELF REPORT
C1706428|T032||HL7V3.0|MALE
C1706428|T032||HL7V3.0|MALE PHENOTYPE
C1706180|T032||HL7V3.0|MALE
C1706180|T032||HL7V3.0|MALE GENDER, SELF REPORTED
C1706180|T032||HL7V3.0|MALE GENDER, SELF REPORT
C1706180|T032||HL7V3.0|MALE GENDER
C0419384|T032||HL7V3.0|MALE BABY
C0419384|T032||HL7V3.0|BABY MALE
C0419384|T032||HL7V3.0|BABY MALE 
C0015780|T032||HL7V3.0|FEMALE
# C0015780|T032||HL7V3.0|F
C0015780|T032||HL7V3.0|FEMALE GENDER, SELF REPORTED
C0015780|T032||HL7V3.0|FEMALE GENDER, SELF REPORT
C0015780|T032||HL7V3.0|FEMALE GENDER
C0015780|T032||HL7V3.0|FEMALE GENDER [DISEASE/FINDING]
C0015780|T032||HL7V3.0|FEMALE 
C0015780|T032||HL7V3.0|FEMALE INDIVIDUAL
C0015780|T032||HL7V3.0|FEMALE STRUCTURE 
C0015780|T032||HL7V3.0|FEMALE STRUCTURE
C0015780|T032||HL7V3.0|FEMALE INDIVIDUAL, NOS
C0015780|T032||HL7V3.0|FEMALE, NOS
C1561593|T032|UN|HL7V3.0|ADMINISTRATIVE GENDER - UNDIFFERENTIATED|UNDIFFERENTIATED
C0036866|T032||HL7V3.0|CHARACTERISTIC, SEX
C0036866|T032||HL7V3.0|CHARACTERISTICS, SEX
C0079399|T032||HL7V3.0|GENDER
C0079399|T032||HL7V3.0|GENDER [DISEASE/FINDING]
C0079399|T032||HL7V3.0|GENDER 
C0079399|T032||HL7V3.0|GENDER (OBSERVABLE ENTITY)
# C1522384|T032||HL7V3.0|SEX
# C1522384|T032||HL7V3.0|SEX OF INDIVIDUAL
# C1522384|T032||HL7V3.0|GENDER
# C1522384|T032||HL7V3.0|SEX OF INDIVIDUAL, NOS
# C1522384|T032||HL7V3.0|SEX, NOS
C1257955|T032||HL7V3.0|GENOTYPIC SEX
C1257955|T032||HL7V3.0|SEX, GENOTYPIC
C1257956|T032||HL7V3.0|PHENOTYPIC SEX
C1257956|T032||HL7V3.0|SEX, PHENOTYPIC
C0278457|T032||HL7V3.0|INDETERMINATE SEX, UNSPECIFIED
C0278457|T032||HL7V3.0|INDETERMINATE SEX
C0278457|T032||HL7V3.0|INDETERMINATE SEX 
C0278457|T032||HL7V3.0|INDETERMINATE SEX NOS
C0278457|T032||HL7V3.0|INDETERMINATE SEX NOS 
C0278457|T032||HL7V3.0|INDETERMINATE SEX 
C0278457|T032||HL7V3.0|INDETERMINATE SEX 
C0278457|T032||HL7V3.0|SEX; INDETERMINATE
C0558141|T032||HL7V3.0|TRANSSEXUAL
C0558141|T032||HL7V3.0|TRANSGENDER