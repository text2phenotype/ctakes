C0270611|T037|702632000|SNOMEDCT_US|BRAIN INJURIES|ACQUIRED BRAIN INJURY
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL INJURY|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|BRAIN DAMAGE, CHRONIC|CHRONIC BRAIN SYNDROME (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|BRAIN CONCUSSION|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|BRAIN CONCUSSIONS|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION, BRAIN|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION |CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CEREBRAL CONCUSSIONS|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION, CEREBRAL|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION NOS|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|COMMOTIO CEREBRI|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|BRAIN CONCUSSION [DISEASE/FINDING]|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CEREBRAL CONCUSSION|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION |CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION NOS |CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION INJURY OF BRAIN |CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION INJURY OF BRAIN|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|BRAIN--CONCUSSION|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|MILD TRAUMATIC BRAIN INJURY|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|MTBI - MILD TRAUMATIC BRAIN INJURY|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|NOT GREAT BUT WON'T RETURN FALSE POSITIVES|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION, UNSPECIFIED|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|NEURO: CONCUSSION|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION INJURY OF BRAIN |CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|BRAIN; COMMOTIO|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|BRAIN; CONCUSSION|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CEREBRAL; CONCUSSION|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CEREBRI; COMMOTIO|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|COMMOTIO; BRAIN|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION; BRAIN|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION; CEREBRAL|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|CONCUSSION (BRAIN)|CONCUSSION INJURY OF BRAIN
C0006107|T037|110030002|SNOMEDCT_US|INJURY;CONCUSSION;HEAD|CONCUSSION INJURY OF BRAIN
C0852861|T037||SNOMEDCT_US|BRAIN DAMAGE (EXCLUDING PERINATAL)
C0852861|T037||SNOMEDCT_US|BRAIN DAMAGE (EXCL PERINATAL)
C0014557|T037|157437008|SNOMEDCT_US|EPILEPSIES, POST-TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|EPILEPSIES, TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|EPILEPSY, POST TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|EPILEPSY, POST-TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|POST-TRAUMATIC EPILEPSIES|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|POST-TRAUMATIC EPILEPSY|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|TRAUMATIC EPILEPSIES|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|TRAUMATIC EPILEPSY|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|SEIZURE DIS POST TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|POST TRAUMATIC SEIZURE DIS|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|DISORDER, POST-TRAUMATIC SEIZURE|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|DISORDERS, POST-TRAUMATIC SEIZURE|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|POST TRAUMATIC SEIZURE DISORDER|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|POST-TRAUMATIC SEIZURE DISORDERS|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|SEIZURE DISORDER, POST TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|SEIZURE DISORDERS, POST-TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|EPILEPSY, POST-TRAUMATIC [DISEASE/FINDING]|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|POST-TRAUMATIC SEIZURE DISORDER|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|EPILEPSY, TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|SEIZURE DISORDER, POST-TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|TRAUMATIC EPILEPSY |TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|PTE - POST-TRAUMATIC EPILEPSY|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|POST-TRAUMATIC EPILEPSY |TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|EPILEPSY; TRAUMATIC|TRAUMATIC EPILEPSY (DISORDER)
C0014557|T037|157437008|SNOMEDCT_US|TRAUMATIC; EPILEPTIC|TRAUMATIC EPILEPSY (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|PNEUMOCEPHALUS|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|AIROCELE, CRANIAL|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|AIROCELES, CRANIAL|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|CRANIAL AIROCELES|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|PNEUMOCYST, CRANIAL|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|CRANIAL PNEUMOCYSTS|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|PNEUMOCYSTS, CRANIAL|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|GAS, INTRACRANIAL|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|CRANIAL AIROCELE|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|CRANIAL PNEUMOCYST|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|PNEUMOCEPHALUS [DISEASE/FINDING]|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|INTRACRANIAL GAS|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|AIROCOELE|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|AIROCELE|PNEUMOCEPHALUS (DISORDER)
C0032268|T037|14415006|SNOMEDCT_US|PNEUMOCEPHALUS |PNEUMOCEPHALUS (DISORDER)
C0751799|T037||SNOMEDCT_US|BRAIN HEMORRHAGE, TRAUMATIC
C0751799|T037||SNOMEDCT_US|BRAIN HEMORRHAGES, TRAUMATIC
C0751799|T037||SNOMEDCT_US|HEMORRHAGE, TRAUMATIC BRAIN
C0751799|T037||SNOMEDCT_US|TRAUMATIC BRAIN HEMORRHAGES
C0751799|T037||SNOMEDCT_US|BRAIN HEMORRHAGE, TRAUMATIC [DISEASE/FINDING]
C0751799|T037||SNOMEDCT_US|TRAUMATIC BRAIN HEMORRHAGE
C0751799|T037||SNOMEDCT_US|BRAIN; HEMORRHAGE, TRAUMATIC
C0751799|T037||SNOMEDCT_US|HEMORRHAGE; BRAIN, TRAUMATIC
C0751813|T037||SNOMEDCT_US|BRAIN INJ CHRONIC
C0751813|T037||SNOMEDCT_US|CHRONIC BRAIN INJ
C0751813|T037||SNOMEDCT_US|ENCEPHALOPATHY POSTTRAUMATIC CHRONIC
C0751813|T037||SNOMEDCT_US|TRAUMATIC ENCEPH CHRONIC
C0751813|T037||SNOMEDCT_US|INJ BRAIN CHRONIC
C0751813|T037||SNOMEDCT_US|ENCEPH POST TRAUMATIC CHRONIC
C0751813|T037||SNOMEDCT_US|CHRONIC POST TRAUMATIC ENCEPH
C0751813|T037||SNOMEDCT_US|BRAIN INJURIES, CHRONIC
C0751813|T037||SNOMEDCT_US|BRAIN INJURY, CHRONIC
C0751813|T037||SNOMEDCT_US|CHRONIC BRAIN INJURIES
C0751813|T037||SNOMEDCT_US|CHRONIC POST TRAUMATIC ENCEPHALOPATHY
C0751813|T037||SNOMEDCT_US|CHRONIC POST-TRAUMATIC ENCEPHALOPATHIES
C0751813|T037||SNOMEDCT_US|ENCEPHALOPATHIES, CHRONIC POST-TRAUMATIC
C0751813|T037||SNOMEDCT_US|ENCEPHALOPATHY, CHRONIC POST-TRAUMATIC
C0751813|T037||SNOMEDCT_US|POST-TRAUMATIC ENCEPHALOPATHIES, CHRONIC
C0751813|T037||SNOMEDCT_US|POST-TRAUMATIC ENCEPHALOPATHY, CHRONIC
C0751813|T037||SNOMEDCT_US|CHRONIC TRAUMATIC ENCEPHALOPATHY
C0751813|T037||SNOMEDCT_US|ENCEPHALOPATHY, CHRONIC TRAUMATIC
C0751813|T037||SNOMEDCT_US|TRAUMATIC ENCEPHALOPATHIES, CHRONIC
C0751813|T037||SNOMEDCT_US|BRAIN INJURY, CHRONIC [DISEASE/FINDING]
C0751813|T037||SNOMEDCT_US|CHRONIC BRAIN INJURY
C0751813|T037||SNOMEDCT_US|TRAUMATIC ENCEPHALOPATHY, CHRONIC
C0751813|T037||SNOMEDCT_US|CHRONIC POST-TRAUMATIC ENCEPHALOPATHY
C0751813|T037||SNOMEDCT_US|ENCEPHALOPATHY, POST-TRAUMATIC, CHRONIC
C0751813|T037||SNOMEDCT_US|INJURY, BRAIN, CHRONIC
C0751813|T037||SNOMEDCT_US|CHRONIC TRAUMATIC ENCEPHALOPATHY 
C0752219|T037||SNOMEDCT_US|DIFFUSE AXONAL INJURY
C0752219|T037||SNOMEDCT_US|DIFFUSE AXONAL INJ
C0752219|T037||SNOMEDCT_US|AXONAL INJ DIFFUSE
C0752219|T037||SNOMEDCT_US|AXONAL INJURIES, DIFFUSE
C0752219|T037||SNOMEDCT_US|DIFFUSE AXONAL INJURIES
C0752219|T037||SNOMEDCT_US|INJURIES, DIFFUSE AXONAL
C0752219|T037||SNOMEDCT_US|INJURY, DIFFUSE AXONAL
C0752219|T037||SNOMEDCT_US|DAI (DIFFUSE AXONAL INJURY)
C0752219|T037||SNOMEDCT_US|AXONAL INJURY, DIFFUSE
C0752219|T037||SNOMEDCT_US|DIFFUSE AXONAL INJURY [DISEASE/FINDING]
C0752219|T037||SNOMEDCT_US|DAIS (DIFFUSE AXONAL INJURY)
C0686721|T037|102458000|SNOMEDCT_US|SHAKEN INFANT SYNDROME |SHAKEN BABY
C0686721|T037|102458000|SNOMEDCT_US|SHAKEN INFANT SYNDROME|SHAKEN BABY
C0686721|T037|102458000|SNOMEDCT_US|SHAKEN BABY SYNDROME|SHAKEN BABY
C0686721|T037|102458000|SNOMEDCT_US|SHAKEN BABY SYNDROME [DISEASE/FINDING]|SHAKEN BABY
C0686721|T037|102458000|SNOMEDCT_US|SHAKEN BABY SYNDROME |SHAKEN BABY
C0686721|T037|102458000|SNOMEDCT_US|SHAKEN BABY SYNDROME - NON-ACCIDENTAL INJURY|SHAKEN BABY
C0686721|T037|102458000|SNOMEDCT_US|SHAKEN BABY|SHAKEN BABY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN INJURIES|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN INJURY|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|INJURY, BRAIN|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|DAMAGE, BRAIN|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN DAMAGE|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN INJ|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|INJ BRAIN|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN LESION (FROM INJURY)|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN INJURY |ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN INJURY NOS|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN INJURIES [DISEASE/FINDING]|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|INJURIES, BRAIN|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|INJURY;CEREBRAL|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|ACQUIRED BRAIN INJURY|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|INTRACEREBRAL INJURY|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|INTRACEREBRAL INJURY NOS|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN INJURY NOS |ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|CEREBRAL DAMAGE|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|ACQUIRED BRAIN INJURY |ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN DAMAGE |ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN TISSUE INJURY|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN; DAMAGE|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN; INJURY|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|CEREBRAL; INJURY|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|DAMAGE; BRAIN|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|INJURY; BRAIN|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|INJURY; CEREBRAL|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|BRAIN DAMAGE, NOS|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|INJURY;BRAIN;ACQUIRED|ACQUIRED BRAIN INJURY
C0270611|T037|702632000|SNOMEDCT_US|CEREBRAL INJURY|ACQUIRED BRAIN INJURY
C0876926|T037|51996004|SNOMEDCT_US|ENCEPH TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC BRAIN INJ|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|INJ BRAIN TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN INJ TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC ENCEPH|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC BRAIN INJURY|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC BRAIN INJURY |TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN INJURY DUE TO TRAUMA|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN TRAUMA|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN DAMAGE (TRAUMATIC)|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TBI|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN DAMAGE - TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC ENCEPHALOPATHY|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC ENCEPHALOPATHY |TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC BRAIN DAMAGE |TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC BRAIN DAMAGE|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN DAMAGE TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|ENCEPHALOPATHY, TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TBI (TRAUMATIC BRAIN INJURY)|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMA, BRAIN|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|INJURY, BRAIN, TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN DAMAGE - TRAUMATIC |TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC BRAIN INJURY |TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|ENCEPHALOPATHY; TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC; ENCEPHALOPATHY|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC ENCEPHALOPATHY  [AMBIGUOUS]|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN INJURY (TRAUMATIC)|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN INJURIES, TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN INJURY, TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|INJURIES, TRAUMATIC BRAIN|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|INJURY, TRAUMATIC BRAIN|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC BRAIN INJURIES|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|BRAIN TRAUMAS|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMAS, BRAIN|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|ENCEPHALOPATHIES, TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TRAUMATIC ENCEPHALOPATHIES|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|TBIS (TRAUMATIC BRAIN INJURY)|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C0876926|T037|51996004|SNOMEDCT_US|INJURY;BRAIN;TRAUMATIC|TRAUMATIC ENCEPHALOPATHY (DISORDER)
C1403070|T037||SNOMEDCT_US|BRAIN INJURY CICATRIX
C1403070|T037||SNOMEDCT_US|AKA BRAIN SCAR
C1403070|T037||SNOMEDCT_US|CICATRIX DUE TO BRAIN INJURY 
C1403070|T037||SNOMEDCT_US|CICATRIX DUE TO BRAIN INJURY
C1403070|T037||SNOMEDCT_US|BRAIN; CICATRIX
C1403070|T037||SNOMEDCT_US|BRAIN; SCAR
C1403070|T037||SNOMEDCT_US|SCAR; BRAIN
C1399577|T037||SNOMEDCT_US|ACQUIRED BRAIN DEFORMITY DUE TO INJURY 
C1399577|T037||SNOMEDCT_US|BRAIN INJURY ACQUIRED DEFORMITY
C1399577|T037||SNOMEDCT_US|ACQUIRED BRAIN DEFORMITY DUE TO INJURY
C1399577|T037||SNOMEDCT_US|ACQUIRED BRAIN DEFORMITY
C1399577|T037||SNOMEDCT_US|BRAIN; DEFORMITY, ACQUIRED
C1399577|T037||SNOMEDCT_US|DEFORMITY; BRAIN, ACQUIRED
C2729127|T037||SNOMEDCT_US|CEREBRAL GRANULOMA DUE TO INJURY
C2729127|T037||SNOMEDCT_US|CEREBRAL GRANULOMA DUE TO INJURY 
C2729127|T037||SNOMEDCT_US|BRAIN INJURY CEREBRAL GRANULOMA
C2729128|T037||SNOMEDCT_US|BRAIN HYPERTROPHY DUE TO INJURY 
C2729128|T037||SNOMEDCT_US|BRAIN HYPERTROPHY DUE TO INJURY
C2729128|T037||SNOMEDCT_US|BRAIN INJURY HYPERTROPHY
C2729129|T037||SNOMEDCT_US|BRAIN INDURATION DUE TO INJURY 
C2729129|T037||SNOMEDCT_US|BRAIN INJURY INDURATION
C2729129|T037||SNOMEDCT_US|BRAIN INDURATION DUE TO INJURY
C2729130|T037||SNOMEDCT_US|INTRACRANIAL PNEUMATOCELE DUE TO INJURY 
C2729130|T037||SNOMEDCT_US|INTRACRANIAL PNEUMATOCELE DUE TO INJURY
C2729130|T037||SNOMEDCT_US|BRAIN INJURY INTRACRANIAL PNEUMATOCELE
C2728325|T037||SNOMEDCT_US|MEDULLARY DEPRESSION DUE TO BRAIN INJURY 
C2728325|T037||SNOMEDCT_US|MEDULLARY DEPRESSION DUE TO BRAIN INJURY
C2728325|T037||SNOMEDCT_US|BRAIN INJURY MEDULLARY DEPRESSION
C2728507|T037||SNOMEDCT_US|MOREL-LAVALLEE LESION DUE TO BRAIN INJURY
C2728507|T037||SNOMEDCT_US|MOREL-LAVALLEE LESION DUE TO BRAIN INJURY 
C2728507|T037||SNOMEDCT_US|BRAIN INJURY MOREL-LAVALLEE LESION
C2729131|T037||SNOMEDCT_US|PNEUMOCEPHALUS DUE TO BRAIN INJURY 
C2729131|T037||SNOMEDCT_US|BRAIN INJURY PNEUMOCEPHALUS
C2729131|T037||SNOMEDCT_US|PNEUMOCEPHALUS DUE TO BRAIN INJURY
C2728280|T037||SNOMEDCT_US|BRAIN INJURY RESPIRATORY CENTER DEPRESSION
C2728280|T037||SNOMEDCT_US|RESPIRATORY CENTER DEPRESSION DUE TO BRAIN INJURY
C2728280|T037||SNOMEDCT_US|RESPIRATORY CENTER DEPRESSION DUE TO BRAIN INJURY 
C2728512|T037||SNOMEDCT_US|SPEECH IMPEDIMENT DUE TO BRAIN INJURY
C2728512|T037||SNOMEDCT_US|BRAIN INJURY SPEECH IMPEDIMENT DUE TO ORGANIC LESION
C2728512|T037||SNOMEDCT_US|SPEECH IMPEDIMENT DUE TO ORGANIC LESION
C2728512|T037||SNOMEDCT_US|SPEECH IMPEDIMENT DUE TO BRAIN INJURY 
C0433845|T037|209868002|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|CORTEX (CEREBRAL) LACER WITH OPEN INTCRAN WOUND, WITH PROLONGED LOC, W/O RTRN TO PECL|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|OPN CORTEX LAC-DEEP COMA|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433845|T037|209868002|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C3509561|T037||SNOMEDCT_US|BIRTH TRAUMA BRAIN DAMAGE
C3509561|T037||SNOMEDCT_US|BRAIN DAMAGE DUE TO BIRTH TRAUMA
C3509561|T037||SNOMEDCT_US|BRAIN DAMAGE DUE TO BIRTH TRAUMA 
C0149844|T037|34663006|SNOMEDCT_US|BRAIN CONTUSIONS|CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|CONTUSION, BRAIN|CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|CONTUSIONS, BRAIN|CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|BRAIN CONTUSION|CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|CONTUSION OF BRAIN|CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|CONTUSION OF BRAIN |CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|HEAD INJURY CONTUSION OF BRAIN|CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|CONTUSIONAL BRAIN INJURY|CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|CONTUSION OF BRAIN |CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|BRAIN; CONTUSION|CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|CONTUSION; BRAIN|CONTUSION OF BRAIN (DISORDER)
C0149844|T037|34663006|SNOMEDCT_US|CONTUSION OF BRAIN, NOS|CONTUSION OF BRAIN (DISORDER)
C0750973|T037||SNOMEDCT_US|ENCEPH POST TRAUMATIC
C0750973|T037||SNOMEDCT_US|POST TRAUMATIC ENCEPH
C0750973|T037||SNOMEDCT_US|ENCEPHALOPATHIES, POST-TRAUMATIC
C0750973|T037||SNOMEDCT_US|ENCEPHALOPATHY, POST TRAUMATIC
C0750973|T037||SNOMEDCT_US|POST TRAUMATIC ENCEPHALOPATHY
C0750973|T037||SNOMEDCT_US|POST-TRAUMATIC ENCEPHALOPATHIES
C0750973|T037||SNOMEDCT_US|POST-TRAUMATIC ENCEPHALOPATHY
C0750973|T037||SNOMEDCT_US|ENCEPHALOPATHY, POST-TRAUMATIC
C0750971|T037|262689001|SNOMEDCT_US|CEREBRAL CONTUSION|CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CEREBRAL CONTUSION |CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CONTUSION, CORTICAL|CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CONTUSIONS, CORTICAL|CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CORTICAL CONTUSIONS|CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CONTUSION;CEREBRAL|CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CORTICAL CONTUSION|CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CONTUSION OF CEREBRUM|CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CONTUSION OF CEREBRUM |CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CEREBRAL; CONTUSION|CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CONTUSION; CEREBRAL|CONTUSION OF CEREBRUM (DISORDER)
C0750971|T037|262689001|SNOMEDCT_US|CEREBRAL CONTUSION, NOS|CONTUSION OF CEREBRUM (DISORDER)
C0750972|T037||SNOMEDCT_US|POST CONCUSSIVE ENCEPH
C0750972|T037||SNOMEDCT_US|ENCEPH POST CONCUSSIVE
C0750972|T037||SNOMEDCT_US|ENCEPHALOPATHIES, POST-CONCUSSIVE
C0750972|T037||SNOMEDCT_US|ENCEPHALOPATHY, POST CONCUSSIVE
C0750972|T037||SNOMEDCT_US|POST CONCUSSIVE ENCEPHALOPATHY
C0750972|T037||SNOMEDCT_US|POST-CONCUSSIVE ENCEPHALOPATHIES
C0750972|T037||SNOMEDCT_US|POST-CONCUSSIVE ENCEPHALOPATHY
C0750972|T037||SNOMEDCT_US|ENCEPHALOPATHY, POST-CONCUSSIVE
C0452047|T037|210038008|SNOMEDCT_US|FOCAL BRAIN INJURY|FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|FOCAL BRAIN INJ|FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|BRAIN INJ FOCAL|FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|BRAIN INJURY, FOCAL|FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|INJURIES, FOCAL BRAIN|FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|INJURY, FOCAL BRAIN|FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|BRAIN INJURIES, FOCAL|FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|FOCAL BRAIN INJURIES|FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|FOCAL BRAIN INJURY |FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|BRAIN; INJURY, FOCAL|FOCAL BRAIN INJURY (DISORDER)
C0452047|T037|210038008|SNOMEDCT_US|INJURY; BRAIN, FOCAL|FOCAL BRAIN INJURY (DISORDER)
C0085742|T037||SNOMEDCT_US|ACUTE BRAIN INJURY
C0085742|T037||SNOMEDCT_US|BRAIN INJURY, ACUTE
C0085742|T037||SNOMEDCT_US|INJURY, ACUTE BRAIN
C0085742|T037||SNOMEDCT_US|INJ ACUTE BRAIN
C0085742|T037||SNOMEDCT_US|ACUTE BRAIN INJ
C0085742|T037||SNOMEDCT_US|BRAIN INJ ACUTE
C0085742|T037||SNOMEDCT_US|INJURIES, ACUTE BRAIN
C0085742|T037||SNOMEDCT_US|ACUTE BRAIN INJURIES
C0085742|T037||SNOMEDCT_US|BRAIN INJURIES, ACUTE
C0272945|T037|78914008|SNOMEDCT_US|BRAIN LACERATION|LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|LACERATION, BRAIN|LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|LACERATIONS, BRAIN|LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|LACERATION OF BRAIN |LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|LACERATING BRAIN INJURY|LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|LACERATION OF BRAIN|LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|LACERATION OF BRAIN |LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|BRAIN; LACERATION|LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|LACERATION; BRAIN|LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|LACERATION OF BRAIN, NOS|LACERATION OF BRAIN (DISORDER)
C0272945|T037|78914008|SNOMEDCT_US|BRAIN LACERATIONS|LACERATION OF BRAIN (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|DIFFUSE BRAIN INJURY|DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|BRAIN INJ DIFFUSE|DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|BRAIN INJURY, DIFFUSE|DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|DIFFUSE BRAIN INJURIES|DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|INJURIES, DIFFUSE BRAIN|DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|INJURY, DIFFUSE BRAIN|DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|DIFFUSE AXONAL BRAIN INJURY|DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|DIFFUSE BRAIN INJURY |DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|BRAIN INJURIES, DIFFUSE|DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|BRAIN; INJURY, DIFFUSE|DIFFUSE BRAIN INJURY (DISORDER)
C0433856|T037|262693007|SNOMEDCT_US|INJURY; BRAIN, DIFFUSE|DIFFUSE BRAIN INJURY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ANOXIC ENCEPHALOPATHY|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ANOXIC ENCEPH|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|BRAIN DAMAGE, ANOXIC|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|DAMAGE, ANOXIC BRAIN|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ANOXIC ENCEPHALOPATHIES|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ENCEPHALOPATHIES, ANOXIC|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ENCEPHALOPATHY, ANOXIC|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ANOXIC BRAIN DAMAGE|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ANOXIC ENCEPHALOPATHY |ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ANOXIC BRAIN INJURY|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ANOXIC BRAIN DAMAGE, NOS|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ANOXIC ENCEPHALOPATHY, NOS|ANOXIC ENCEPHALOPATHY (DISORDER)
C0003132|T037|389098007|SNOMEDCT_US|ANOXIC ENCEPHALOPATHY [DUP] |ANOXIC ENCEPHALOPATHY (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PERSISTENT VEGETATIVE STATE|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PERSISTENT VEGETATIVE STATES|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|VEGETATIVE STATES, PERSISTENT|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PERSISTENT VEGETATIVE STATE |PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PERSISTENT UNAWARENESS STATES|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|STATE, PERSISTENT UNAWARENESS|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|STATES, PERSISTENT UNAWARENESS|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|UNAWARENESS STATE, PERSISTENT|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|UNAWARENESS STATES, PERSISTENT|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|STATE, PERSISTENT VEGETATIVE|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|STATES, PERSISTENT VEGETATIVE|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PERSISTENT VEGTV STATE|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PERSISTENT UNAWARENESS STATE|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PERSISTENT VEGETATIVE STATE [DISEASE/FINDING]|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PVS (PERSISTENT VEGETATIVE STATE)|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|VEGETATIVE STATE, PERSISTENT|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PVSS (PERSISTENT VEGETATIVE STATE)|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PERSISTENT VEGETATIVE STATE |PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|CHRONIC VEGETATIVE STATE|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|VEGETATIVE STATE CHRONIC|PERSISTENT VEGETATIVE STATE (DISORDER)
C0242670|T037|24473007|SNOMEDCT_US|PVS - PERSISTENT VEGETATIVE STATE|PERSISTENT VEGETATIVE STATE (DISORDER)
C0549117|T037|192199002|SNOMEDCT_US|CAN BE DUE TO A NEURODEGENERATIVE DISEASE BUT WORTH KNOWING - IF YOU HAD A SEPERATE SECTION FOR NEURO DEGEN DZ I WOULD INCLUDE THERE AS WELL|[X]FRONTAL LOBE SYNDROME
C0549117|T037|192199002|SNOMEDCT_US|FRONTAL LOBE SYNDROME |[X]FRONTAL LOBE SYNDROME
C0549117|T037|192199002|SNOMEDCT_US|FRONTAL LOBE SYNDROME |[X]FRONTAL LOBE SYNDROME
C0549117|T037|192199002|SNOMEDCT_US|[X]FRONTAL LOBE SYNDROME|[X]FRONTAL LOBE SYNDROME
C0549117|T037|192199002|SNOMEDCT_US|FRONTAL LOBE; SYNDROME|[X]FRONTAL LOBE SYNDROME
C0549117|T037|192199002|SNOMEDCT_US|SYNDROME; FRONTAL LOBE|[X]FRONTAL LOBE SYNDROME
C0006110|T037||SNOMEDCT_US|NOT APPLICABLE TO THIS FORM, BUT MIGHT AS WELL INCLUDE
C0006110|T037||SNOMEDCT_US|CEREBRAL DEATH
C0006110|T037||SNOMEDCT_US|DEATH, BRAIN
C0006110|T037||SNOMEDCT_US|BRAIN DEATH 
C0006110|T037||SNOMEDCT_US|BRAIN DEADS
C0006110|T037||SNOMEDCT_US|BRAIN DEATH [DISEASE/FINDING]
C0006110|T037||SNOMEDCT_US|COMA DEPASSE
C0006110|T037||SNOMEDCT_US|BRAIN DEAD
C3508472|T037||SNOMEDCT_US|BRAIN INJURY TRAUMATIC MILD 
C3508472|T037||SNOMEDCT_US|BRAIN INJURY TRAUMATIC MILD
C3508472|T037||SNOMEDCT_US|MILD TRAUMATIC BRAIN INJURY
C3508472|T037||SNOMEDCT_US|INJURY, BRAIN, TRAUMATIC MILD
C0272927|T037|9015001|SNOMEDCT_US|CLOSED TRAUMATIC BRAIN INJURY|BRAIN INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0272927|T037|9015001|SNOMEDCT_US|BRAIN INJURY WITHOUT OPEN INTRACRANIAL WOUND|BRAIN INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0272927|T037|9015001|SNOMEDCT_US|BRAIN INJURY WITHOUT OPEN INTRACRANIAL WOUND |BRAIN INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0272927|T037|9015001|SNOMEDCT_US|BRAIN INJURY WITHOUT OPEN INTRACRANIAL WOUND |BRAIN INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0272927|T037|9015001|SNOMEDCT_US|BRAIN INJURY WITHOUT OPEN INTRACRANIAL WOUND, NOS|BRAIN INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0021879|T037||SNOMEDCT_US|BRAIN INJURY NEC
C0021879|T037||SNOMEDCT_US|INTCRAN INJ OF OTH AND UNSPEC NATURE, W/O MENT OF OPEN INTCRAN WOUND, WITH STATE OF CONS UNSPEC
C0021879|T037||SNOMEDCT_US|INTRACRANIAL INJURY OF OTHER AND UNSPECIFIED NATURE WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS
C1140716|T037|126944002|SNOMEDCT_US|HYPOXIC ENCEPH|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|ENCEPH HYPOXIC|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|BRAIN DAMAGE, HYPOXIC|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|DAMAGE, HYPOXIC BRAIN|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|ENCEPHALOPATHIES, HYPOXIC|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|HYPOXIC ENCEPHALOPATHIES|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|HYPOXIC BRAIN DAMAGE|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|BRAIN DAMAGE DUE TO HYPOXIA|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|HYPOXIC BRAIN INJURY|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|HYPOXIC-ISCHEMIC BRAIN INJURY|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|HYPOXIC-ISCHAEMIC BRAIN INJURY|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|HYPOXIC ENCEPHALOPATHY|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|ENCEPHALOPATHY, HYPOXIC|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C1140716|T037|126944002|SNOMEDCT_US|BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN |BRAIN DISORDER RESULTING FROM A PERIOD OF IMPAIRED OXYGEN DELIVERY TO THE BRAIN
C0338418|T037|111897007|SNOMEDCT_US|ACUTE NECROTIZING ENCEPHALITIDES|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|ACUTE NECROTIZING ENCEPHALITIS|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|ENCEPHALITIDES, ACUTE NECROTIZING|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|NECROTIZING ENCEPHALITIDES, ACUTE|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|NECROTIZING ENCEPHALITIS, ACUTE|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|ENCEPH ACUTE NECROTIZING|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|VIRAL ENCEPHALITIS ACUTE NECROTIZING|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|ACUTE NECROTIZING ENCEPHALITIS |ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|ACUTE NECROTISING ENCEPHALITIS|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|ACUTE NECROTIZING VIRAL ENCEPHALITIS|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|ACUTE NECROTISING VIRAL ENCEPHALITIS|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|ACUTE NECROTIZING ENCEPHALITIS |ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C0338418|T037|111897007|SNOMEDCT_US|ENCEPHALITIS, ACUTE NECROTIZING|ACUTE NECROTIZING ENCEPHALITIS (DISORDER)
C3897170|T037||SNOMEDCT_US|WHITE MATTER INJURY
C1456496|T037|127294003|SNOMEDCT_US|BRAIN DAMAGE|TRAUMATIC AND/OR NON-TRAUMATIC BRAIN INJURY (DISORDER)
C1456496|T037|127294003|SNOMEDCT_US|TRAUMATIC AND/OR NON-TRAUMATIC BRAIN INJURY|TRAUMATIC AND/OR NON-TRAUMATIC BRAIN INJURY (DISORDER)
C1456496|T037|127294003|SNOMEDCT_US|TRAUMATIC AND/OR NON-TRAUMATIC BRAIN INJURY |TRAUMATIC AND/OR NON-TRAUMATIC BRAIN INJURY (DISORDER)
C0149843|T037|230283005|SNOMEDCT_US|PUNCH DRUNK SYNDROME|PUNCH DRUNK SYNDROME (DISORDER)
C0149843|T037|230283005|SNOMEDCT_US|PUNCH DRUNK SYNDROME |PUNCH DRUNK SYNDROME (DISORDER)
C0149843|T037|230283005|SNOMEDCT_US|HEAD INJURY WITH DEMENTIA PUNCH DRUNK SYNDROME|PUNCH DRUNK SYNDROME (DISORDER)
C0149843|T037|230283005|SNOMEDCT_US|BOXER'S DEMENTIA|PUNCH DRUNK SYNDROME (DISORDER)
C0149843|T037|230283005|SNOMEDCT_US|DEMENTIA PUGILISTICA|PUNCH DRUNK SYNDROME (DISORDER)
C0149843|T037|230283005|SNOMEDCT_US|PUNCHDRUNK ENCEPHALOPATHY|PUNCH DRUNK SYNDROME (DISORDER)
C0149843|T037|230283005|SNOMEDCT_US|PUNCH DRUNK SYNDROME |PUNCH DRUNK SYNDROME (DISORDER)
C0160293|T037||SNOMEDCT_US|BRAIN INJURY NEC-NO COMA
C0160293|T037||SNOMEDCT_US|INTCRAN INJ OF OTH AND UNSPEC NATURE, W/O MENT OF OPEN INTCRAN WOUND, WITH NO LOC
C0160293|T037||SNOMEDCT_US|INTRACRANIAL INJURY OF OTHER AND UNSPECIFIED NATURE WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS
C0160294|T037||SNOMEDCT_US|BRAIN INJ NEC-BRIEF COMA
C0160294|T037||SNOMEDCT_US|INTCRAN INJ OF OTH AND UNSPEC NATURE, W/O MENT OF OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160294|T037||SNOMEDCT_US|INTRACRANIAL INJURY OF OTHER AND UNSPECIFIED NATURE WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160298|T037||SNOMEDCT_US|BRAIN INJ NEC-COMA NOS
C0160298|T037||SNOMEDCT_US|INTCRAN INJ OF OTH AND UNSPEC NATURE, W/O MENT OF OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURA
C0160298|T037||SNOMEDCT_US|INTRACRANIAL INJURY OF OTHER AND UNSPECIFIED NATURE WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION
C0006109|T037|78689005|SNOMEDCT_US|BRAIN DAMAGE, CHRONIC|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|CHRONIC BRAIN DAMAGE|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|ENCEPH CHRONIC|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|CHRONIC ENCEPH|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|BRAIN SYNDROME CHRONIC|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|SYNDROME BRAIN CHRONIC|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|ENCEPHALOPATHY, CHRONIC|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|BRAIN DAMAGE, CHRONIC [DISEASE/FINDING]|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|CHRONIC ENCEPHALOPATHY|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|ENCEPHALOPATHY CHRONIC|CHRONIC BRAIN SYNDROME (DISORDER)
C0006109|T037|78689005|SNOMEDCT_US|CHRONIC ENCEPHALOPATHY, NOS|CHRONIC BRAIN SYNDROME (DISORDER)
C0160292|T037||SNOMEDCT_US|INTRACRANIAL INJURY OF OTHER AND UNSPECIFIED NATURE
C0021878|T037||SNOMEDCT_US|INTRACRANIAL INJURY OF OTHER AND UNSPECIFIED NATURE WITHOUT MENTION OF OPEN INTRACRANIAL WOUND
C1321905|T037|229716009|SNOMEDCT_US|DYSFUNCTION, MINIMAL BRAIN|MINIMAL BRAIN DYSFUNCTION (DISORDER)
C1321905|T037|229716009|SNOMEDCT_US|MINIMAL BRAIN DYSFUNCTION|MINIMAL BRAIN DYSFUNCTION (DISORDER)
C1321905|T037|229716009|SNOMEDCT_US|MINIMAL BRAIN DYSFUNCTION |MINIMAL BRAIN DYSFUNCTION (DISORDER)
C1321905|T037|229716009|SNOMEDCT_US|MBD - MINIMAL BRAIN DYSFUNCTION|MINIMAL BRAIN DYSFUNCTION (DISORDER)
C1321905|T037|229716009|SNOMEDCT_US|MINIMAL BRAIN DISORDERS|MINIMAL BRAIN DYSFUNCTION (DISORDER)
C1321905|T037|229716009|SNOMEDCT_US|BRAIN DYSFUNCTION, MINIMAL|MINIMAL BRAIN DYSFUNCTION (DISORDER)
C0695222|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED
C0695222|T037||SNOMEDCT_US|OPN CEREBEL CONT-CONCUSS
C0695224|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED
C0695224|T037||SNOMEDCT_US|OPN CEREBELL LAC-CONCUSS
C0433815|T037|209835009|SNOMEDCT_US|CORTEX (CEREBRAL) CONTU W/O MENT OF OPEN INTCRAN WOUND, STATE OF CONSCIOUSNESS UNSPEC|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433815|T037|209835009|SNOMEDCT_US|CEREBRAL CORTX CONTUSION|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433815|T037|209835009|SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433815|T037|209835009|SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH UNSPECIFIED STATE OF CONSCIOUSNESS |CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433815|T037|209835009|SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH UNSPECIFIED STATE OF CONSCIOUSNESS|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433815|T037|209835009|SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, STATE OF CONSCIOUSNESS UNSPECIFIED|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433815|T037|209835009|SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, STATE OF CONSCIOUSNESS UNSPECIFIED|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433821|T037|209841002|SNOMEDCT_US|CORTEX (CEREBRAL) CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433821|T037|209841002|SNOMEDCT_US|CORTEX CONTUS-COMA NOS|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433821|T037|209841002|SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433821|T037|209841002|SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION |CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433821|T037|209841002|SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433821|T037|209841002|SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433846|T037|209853003|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND (DISORDER)
C0433846|T037|209853003|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND |CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND (DISORDER)
C0433846|T037|209853003|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND (DISORDER)
C0433846|T037|209853003|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND (DISORDER)
C0433847|T037|209854009|SNOMEDCT_US|CORTEX (CEREBRAL) LACER W/O MENT OF OPEN INTCRAN WOUND, WITH STATE OF CONSCIOUSNESS UNSPEC|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433847|T037|209854009|SNOMEDCT_US|CEREBRAL CORTEX LACERAT|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433847|T037|209854009|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433847|T037|209854009|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS |CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433847|T037|209854009|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433847|T037|209854009|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH STATE OF CONSCIOUSNESS UNSPECIFIED|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433847|T037|209854009|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH STATE OF CONSCIOUSNESS UNSPECIFIED|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433848|T037|209855005|SNOMEDCT_US|CORTEX (CEREBRAL) LACER W/O MENT OF OPEN INTCRAN WOUND, WITH NO LOC|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0433848|T037|209855005|SNOMEDCT_US|CORTEX LACERAT W/O COMA|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0433848|T037|209855005|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0433848|T037|209855005|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS |CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0433848|T037|209855005|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0433848|T037|209855005|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0433853|T037|209860009|SNOMEDCT_US|CORTEX (CEREBRAL) LACER W/O MENT OF OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433853|T037|209860009|SNOMEDCT_US|CORTEX LACERAT-COMA NOS|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433853|T037|209860009|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION |CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433853|T037|209860009|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433853|T037|209860009|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433853|T037|209860009|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433854|T037|209861008|SNOMEDCT_US|CORTEX (CEREBRAL) LACER W/O MENT OF OPEN INTCRAN WOUND, WITH CONCUSSION, UNSPEC|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0433854|T037|209861008|SNOMEDCT_US|CORTEX LACERAT-CONCUSS|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0433854|T037|209861008|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED |CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0433854|T037|209861008|SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0433854|T037|209861008|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0433854|T037|209861008|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0859613|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH NO LOC
C0160131|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160131|T037||SNOMEDCT_US|CORTEX CONTUS-BRIEF COMA
C0160131|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160131|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF LOSS OF CONSCIOUSNESS
C0160131|T037||SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF LOSS OF CONSCIOUSNESS
C0272955|T037|209838006|SNOMEDCT_US|CORTEX CONTUSION WITHOUT OPEN INTRACRANIAL WOUND AND WITH MODERATE LOSS OF CONSCIOUSNESS (1-24 HOURS) |CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX CONTUSION WITHOUT OPEN INTRACRANIAL WOUND AND WITH MODERATE LOSS OF CONSCIOUSNESS (1-24 HOURS)|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX (CEREBRAL) CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH MODERATE LOC|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX CONTUS-MOD COMA|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS |CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CONTUSION OF CORTEX W/O OPEN INTRACRANIAL WOUND, WITH MODERATE LOC (1-24 HOURS)|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX CONTUSION WITHOUT OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS (1-24 HOURS)|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX CONTUSION WITHOUT OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS (1-24 HOURS) |CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272955|T037|209838006|SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITHOUT MENTION OF INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0160133|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH PROLONGED LOC AND RTRN TO PECL
C0160133|T037||SNOMEDCT_US|CORTX CONTUS-PROLNG COMA
C0160133|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160133|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160133|T037||SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160134|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH PROLONGED LOC, W/O RTRN TO PECL
C0160134|T037||SNOMEDCT_US|CORTEX CONTUS-DEEP COMA
C0160134|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160134|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160134|T037||SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0695217|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH CONCUSSION, UNSPEC
C0695217|T037||SNOMEDCT_US|CORTEX CONTUS-CONCUS NOS
C0695217|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED
C0695217|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED
C0695217|T037||SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED
C0160138|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU WITH OPEN INTCRAN WOUND, W/O MENT OF SPECIFIC STATE OF CONSCIOUSNESS
C0160138|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH STATE OF CONSCIOUSNESS UNSPECIFIED
C0160138|T037||SNOMEDCT_US|CORTEX CONTUSION/OPN WND
C0160138|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND, WITHOUT MENTION OF SPECIFIC STATE OF CONSCIOUSNESS
C0160138|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS
C0160138|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITHOUT MENTION OF SPECIFIC STATE OF CONSCIOUSNESS
C0160138|T037||SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITHOUT MENTION OF SPECIFIC STATE OF CONSCIOUSNESS
C0160140|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU WITH OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160140|T037||SNOMEDCT_US|OPN CORT CONTUS-BRF COMA
C0160140|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160140|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH BRIEF LOSS OF CONSCIOUSNESS
C0160140|T037||SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH BRIEF LOSS OF CONSCIOUSNESS
C0160141|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU WITH OPEN INTCRAN WOUND, WITH MODERATE LOC
C0160141|T037||SNOMEDCT_US|OPN CORT CONTUS-MOD COMA
C0160141|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS
C0160141|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS
C0160141|T037||SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS
C0160142|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU WITH OPEN INTCRAN WOUND, WITH PROLONGED LOC AND RTRN TO PECL
C0160142|T037||SNOMEDCT_US|OPN CORT CONTU-PROL COMA
C0160142|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160142|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160142|T037||SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160143|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU WITH OPEN INTCRAN WOUND, WITH PROLONGED LOC, W/O RTRN TO PECL
C0160143|T037||SNOMEDCT_US|OPN CORT CONTU-DEEP COMA
C0160143|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160143|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160143|T037||SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0859614|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTU WITH OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION
C0160149|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACER W/O MENT OF OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160149|T037||SNOMEDCT_US|CORTEX LACERA-BRIEF COMA
C0160149|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160149|T037||SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF LOSS OF CONSCIOUSNESS
C0160149|T037||SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF LOSS OF CONSCIOUSNESS
C0160150|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACER W/O MENT OF OPEN INTCRAN WOUND, WITH MODERATE LOC
C0160150|T037||SNOMEDCT_US|CORTEX LACERAT-MOD COMA
C0160150|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS
C0160150|T037||SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS
C0160150|T037||SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS
C0160151|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACER W/O MENT OF OPEN INTCRAN WOUND, WITH PROLONGED LOC AND RTRN TO PECL
C0160151|T037||SNOMEDCT_US|CORTEX LACERAT-PROL COMA
C0160151|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160151|T037||SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160151|T037||SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160152|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACER W/O MENT OF OPEN INTCRAN WOUND, WITH PROLONGED LOC, W/O RTRN TO PECL
C0160152|T037||SNOMEDCT_US|CORTEX LACERAT-DEEP COMA
C0160152|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160152|T037||SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160152|T037||SNOMEDCT_US|CORTEX LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS, WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160158|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACER WITH OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160158|T037||SNOMEDCT_US|OPN CORTX LAC-BRIEF COMA
C0160158|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITH OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160158|T037||SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH BRIEF LOSS OF CONSCIOUSNESS
C0160158|T037||SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH BRIEF LOSS OF CONSCIOUSNESS
C0160159|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACER WITH OPEN INTCRAN WOUND, WITH MODERATE LOC
C0160159|T037||SNOMEDCT_US|OPN CORTX LACER-MOD COMA
C0160159|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS
C0160159|T037||SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS
C0160159|T037||SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MODERATE LOSS OF CONSCIOUSNESS
C0160160|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACER WITH OPEN INTCRAN WOUND, WITH PROLONGED LOC AND RTRN TO PECL
C0160160|T037||SNOMEDCT_US|OPN CORTX LAC-PROLN COMA
C0160160|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160160|T037||SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160160|T037||SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0859615|T037||SNOMEDCT_US|CORTEX (CEREBRAL) LACER WITH OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION
C0160165|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH STATE OF CONS UNSPEC
C0160165|T037||SNOMEDCT_US|CEREBEL/BRAIN STM CONTUS
C0160165|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS
C0160166|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH NO LOC
C0160166|T037||SNOMEDCT_US|CEREBELL CONTUS W/O COMA
C0160166|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS
C0160167|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160167|T037||SNOMEDCT_US|CEREBELL CONTUS-BRF COMA
C0160167|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160168|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH MODERATE LOC
C0160168|T037||SNOMEDCT_US|CEREBELL CONTUS-MOD COMA
C0160168|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS
C0160170|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH PROLONGED LOC, W/O RTRN TO PECL
C0160170|T037||SNOMEDCT_US|CEREBEL CONTUS-DEEP COMA
C0160170|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160171|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION
C0160171|T037||SNOMEDCT_US|CEREBELL CONTUS-COMA NOS
C0160171|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION
C0695221|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH CONCUSSION, UNSPEC
C0695221|T037||SNOMEDCT_US|CEREBELL CONTUS-CONCUSS
C0695221|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED
C0160174|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU WITH OPEN INTCRAN WOUND, WITH STATE OF CONSCIOUSNESS UNSPEC
C0160174|T037||SNOMEDCT_US|CEREBEL CONTUS W OPN WND
C0160174|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITH OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS
C0160176|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU WITH OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160176|T037||SNOMEDCT_US|OPN CEREBE CONT-BRF COMA
C0160176|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160177|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS
C0160177|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU WITH OPEN INTCRAN WOUND, WITH MODERATE LOC
C0160177|T037||SNOMEDCT_US|OPN CEREBE CONT-MOD COMA
C0160178|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU WITH OPEN INTCRAN WOUND, WITH PROLONGED LOC AND RETURN TO PECL
C0160178|T037||SNOMEDCT_US|OPN CEREBE CONT-PROL COM
C0160178|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160179|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU WITH OPEN INTCRAN WOUND, WITH PROLONGED LOC, W/O RETURN TO PECL
C0160179|T037||SNOMEDCT_US|OPN CEREBE CONT-DEEP COM
C0160179|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160180|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU WITH OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION
C0160180|T037||SNOMEDCT_US|OPN CEREBE CONT-COMA NOS
C0160180|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION
C0160183|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER W/O MENT OF OPEN INTCRAN WOUND, WITH STATE OF CONSCIOUSNESS UNSPEC
C0160183|T037||SNOMEDCT_US|CEREBEL/BRAIN STEM LACER
C0160183|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS
C0160184|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER W/O MENT OF OPEN INTCRAN WOUND, WITH NO LOC
C0160184|T037||SNOMEDCT_US|CEREBEL LACERAT W/O COMA
C0160184|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS
C0160185|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER W/O MENT OF OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160185|T037||SNOMEDCT_US|CEREBEL LACER-BRIEF COMA
C0160185|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN 1 HOUR] LOSS OF CONSCIOUSNESS
C0160186|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER W/O MENT OF OPEN INTCRAN WOUND, WITH MODERATE LOC
C0160186|T037||SNOMEDCT_US|CEREBEL LACERAT-MOD COMA
C0160186|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS
C0160187|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER W/O MENT OF OPEN INTCRAN WOUND, WITH PROLONGED LOC AND RTRN TO PECL
C0160187|T037||SNOMEDCT_US|CEREBEL LACER-PROLN COMA
C0160187|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160188|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER W/O MENT OF OPEN INTCRAN WOUND, WITH PROLONGED LOC, W/O RTRN TO PECL
C0160188|T037||SNOMEDCT_US|CEREBELL LACER-DEEP COMA
C0160188|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160189|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER W/O MENT OF OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION
C0160189|T037||SNOMEDCT_US|CEREBEL LACERAT-COMA NOS
C0160189|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION
C0695223|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER W/O MENT OF OPEN INTCRAN WOUND, WITH CONCUSSION, UNSPEC
C0695223|T037||SNOMEDCT_US|CEREBEL LACER-CONCUSSION
C0695223|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED
C0160192|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER WITH OPEN INTCRAN WOUND, WITH STATE OF CONSCIOUSNESS UNSPEC
C0160192|T037||SNOMEDCT_US|CEREBEL LACER W OPEN WND
C0160192|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITH OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS
C0160194|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER WITH OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160194|T037||SNOMEDCT_US|OPN CEREBEL LAC-BRF COMA
C0160194|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITH OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160195|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER WITH OPEN INTCRAN WOUND, WITH MODERATE LOC
C0160195|T037||SNOMEDCT_US|OPN CEREBEL LAC-MOD COMA
C0160195|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITH OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS
C0160196|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER WITH OPEN INTCRAN WOUND, WITH PROLONGED LOC AND RETURN TO PECL
C0160196|T037||SNOMEDCT_US|OPN CEREBE LAC-PROL COMA
C0160196|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160197|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER WITH OPEN INTCRAN WOUND, WITH PROLONGED LOC, W/O RETURN TO PECL
C0160197|T037||SNOMEDCT_US|OPN CEREBE LAC-DEEP COMA
C0160197|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160198|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACER WITH OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION
C0160198|T037||SNOMEDCT_US|OPN CEREBEL LAC-COMA NOS
C0160198|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITH OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION
C0160201|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, W/O MENT OF OPEN INTCRAN WOUND, WITH STATE OF CONS UNSPEC
C0160201|T037||SNOMEDCT_US|BRAIN LACERATION NEC
C0160201|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS
C0160202|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, W/O MENT OF OPEN INTCRAN WOUND, WITH NO LOC
C0160202|T037||SNOMEDCT_US|BRAIN LACER NEC W/O COMA
C0160202|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS
C0160203|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, W/O MENT OF OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160203|T037||SNOMEDCT_US|BRAIN LAC NEC-BRIEF COMA
C0160203|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160204|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, W/O MENT OF OPEN INTCRAN WOUND, WITH MODERATE LOC
C0160204|T037||SNOMEDCT_US|BRAIN LACER NEC-MOD COMA
C0160204|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS
C0160205|T037||SNOMEDCT_US|OTH AND UNSPEC CEREB LACER AND CONTU, W/O MENT OF OPEN INTCRAN WOUND, PROL LOC AND RTRN TO PECL
C0160205|T037||SNOMEDCT_US|BRAIN LAC NEC-PROLN COMA
C0160205|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS AND RETURN TO PRE- EXISTING CONSCIOUS LEVEL
C0160206|T037||SNOMEDCT_US|OTH AND UNSPEC CEREB LACER AND CONTU, W/O MENT OF OPEN INTCRAN WOUND, PROL LOC, W/O RTRN TO PECL
C0160206|T037||SNOMEDCT_US|BRAIN LAC NEC-DEEP COMA
C0160206|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160207|T037||SNOMEDCT_US|OTH AND UNSPEC CEREB LACER AND CONTU, W/O MENT OF OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION
C0160207|T037||SNOMEDCT_US|BRAIN LACER NEC-COMA NOS
C0160207|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION
C0695225|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, W/O MENT OF OPEN INTCRAN WOUND, WITH CONCUS, UNSPEC
C0695225|T037||SNOMEDCT_US|BRAIN LACER NEC-CONCUSS
C0695225|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED
C0160210|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, WITH OPEN INTCRAN WOUND, WITH STATE OF CONS UNSPEC
C0160210|T037||SNOMEDCT_US|BRAIN LAC NEC W OPEN WND
C0160210|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITH OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS
C0160211|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, WITH OPEN INTCRAN WOUND, WITH NO LOC
C0160211|T037||SNOMEDCT_US|OPN BRAIN LACER W/O COMA
C0160211|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS
C0160212|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, WITH OPEN INTCRAN WOUND, WITH BRIEF LOC
C0160212|T037||SNOMEDCT_US|OPN BRAIN LAC-BRIEF COMA
C0160212|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITH OPEN INTRACRANIAL WOUND, WITH BRIEF [LESS THAN ONE HOUR] LOSS OF CONSCIOUSNESS
C0160213|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, WITH OPEN INTCRAN WOUND, WITH MODERATE LOC
C0160213|T037||SNOMEDCT_US|OPN BRAIN LACER-MOD COMA
C0160213|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITH OPEN INTRACRANIAL WOUND, WITH MODERATE [1-24 HOURS] LOSS OF CONSCIOUSNESS
C0160214|T037||SNOMEDCT_US|OTH AND UNSPEC CEREB LACER AND CONTU, WITH OPEN INTCRAN WOUND, WITH PROL LOC AND RTRN TO PECL
C0160214|T037||SNOMEDCT_US|OPN BRAIN LAC-PROLN COMA
C0160214|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160215|T037||SNOMEDCT_US|OTH AND UNSPEC CEREB LACER AND CONTU, WITH OPEN INTCRAN WOUND, WITH PROL LOC, W/O RTRN TO PECL
C0160215|T037||SNOMEDCT_US|OPEN BRAIN LAC-DEEP COMA
C0160215|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C0160216|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, WITH OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION
C0160216|T037||SNOMEDCT_US|OPN BRAIN LACER-COMA NOS
C0160216|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITH OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION
C0695226|T037||SNOMEDCT_US|OTH AND UNSPEC CEREBRAL LACER AND CONTU, WITH OPEN INTCRAN WOUND, WITH CONCUSSION, UNSPEC
C0695226|T037||SNOMEDCT_US|OPEN BRAIN LACER-CONCUSS
C0695226|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED
C0859744|T037||SNOMEDCT_US|CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND
C0859745|T037||SNOMEDCT_US|CEREBRAL LACERATION & CONTUSION WITH OPEN INTRACRANIAL WOUND
C0859782|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH PROL LOSS CONS AND RTRN TO PECL
C0859782|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTU W/O MENT OF OPEN INTCRAN WOUND, WITH PROL LOC AND RETURN TO PECL
C0160128|T037||SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND
C0160128|T037||SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND
C0160128|T037||SNOMEDCT_US|CORTEX CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND
C0160164|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND
C0160173|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITH OPEN INTRACRANIAL WOUND
C0160182|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITHOUT MENTION OF OPEN INTRACRANIAL WOUND
C0160191|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITH OPEN INTRACRANIAL WOUND
C0160200|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITHOUT MENTION OF OPEN INTRACRANIAL WOUND
C0160209|T037||SNOMEDCT_US|OTHER AND UNSPECIFIED CEREBRAL LACERATION AND CONTUSION, WITH OPEN INTRACRANIAL WOUND
C0160137|T037|87888006|SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160137|T037|87888006|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160137|T037|87888006|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND |CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160137|T037|87888006|SNOMEDCT_US|CONTUSION OF CORTEX WITH OPEN INTRACRANIAL WOUND|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160137|T037|87888006|SNOMEDCT_US|CONTUSION OF CEREBRAL CORTEX WITH OPEN INTRACRANIAL WOUND|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160137|T037|87888006|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND |CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160137|T037|87888006|SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160127|T037|269144002|SNOMEDCT_US|CEREBRAL LACERATION AND CONTUSION|CEREBRAL LACERATION AND CONTUSION (DISORDER)
C0160127|T037|269144002|SNOMEDCT_US|CEREBRAL LACERATION AND CONTUSION |CEREBRAL LACERATION AND CONTUSION (DISORDER)
C0160127|T037|269144002|SNOMEDCT_US|CEREBRAL LACERATION AND CONTUSION NOS|CEREBRAL LACERATION AND CONTUSION (DISORDER)
C0160127|T037|269144002|SNOMEDCT_US|CEREBRAL LACERATION AND CONTUSION |CEREBRAL LACERATION AND CONTUSION (DISORDER)
C0160127|T037|269144002|SNOMEDCT_US|CEREBRAL LACERATION AND CONTUSION NOS |CEREBRAL LACERATION AND CONTUSION (DISORDER)
C0160127|T037|269144002|SNOMEDCT_US|BRAIN LACERATION AND CONTUSION NOS|CEREBRAL LACERATION AND CONTUSION (DISORDER)
C0274278|T037|74472004|SNOMEDCT_US|LATE EFFECT OF INTRACRANIAL INJURY WITHOUT MENTION OF SKULL FRACTURE|LATE EFFECT OF INTRACRANIAL INJURY WITHOUT SKULL FRACTURE (DISORDER)
C0274278|T037|74472004|SNOMEDCT_US|SEQUELAE OF INTRACRANIAL INJURY|LATE EFFECT OF INTRACRANIAL INJURY WITHOUT SKULL FRACTURE (DISORDER)
C0274278|T037|74472004|SNOMEDCT_US|LT EFF INTRACRANIAL INJ|LATE EFFECT OF INTRACRANIAL INJURY WITHOUT SKULL FRACTURE (DISORDER)
C0274278|T037|74472004|SNOMEDCT_US|LATE EFFECT OF INTRACRANIAL INJURY WITHOUT SKULL FRACTURE |LATE EFFECT OF INTRACRANIAL INJURY WITHOUT SKULL FRACTURE (DISORDER)
C0274278|T037|74472004|SNOMEDCT_US|LATE EFFECT OF INTRACRANIAL INJURY WITHOUT SKULL FRACTURE|LATE EFFECT OF INTRACRANIAL INJURY WITHOUT SKULL FRACTURE (DISORDER)
C0274278|T037|74472004|SNOMEDCT_US|LATE EFFECT OF INTRACRANIAL INJURY WITHOUT SKULL FRACTURE |LATE EFFECT OF INTRACRANIAL INJURY WITHOUT SKULL FRACTURE (DISORDER)
C0272961|T037|209845006|SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272961|T037|209845006|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND NO LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272961|T037|209845006|SNOMEDCT_US|CEREBRAL CONTUSION WITH OPEN INTRACRANIAL WOUND WITH NO LOSS OF CONSCIOUSNESS |CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272961|T037|209845006|SNOMEDCT_US|CEREBRAL CONTUSION WITH OPEN INTRACRANIAL WOUND WITH NO LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272961|T037|209845006|SNOMEDCT_US|OPN CORTX CONTUS-NO COMA|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272961|T037|209845006|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND NO LOSS OF CONSCIOUSNESS |CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272961|T037|209845006|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272961|T037|209845006|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS |CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272961|T037|209845006|SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0160175|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS
C0160175|T037||SNOMEDCT_US|OPN CEREBE CONT W/O COMA
C0160193|T037||SNOMEDCT_US|CEREBELLAR OR BRAIN STEM LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS
C0160193|T037||SNOMEDCT_US|OPN CEREBEL LAC W/O COMA
C0272967|T037|73413009|SNOMEDCT_US|CEREBRAL CONTUSION WITH OPEN INTRACRANIAL WOUND WITH CONCUSSION |CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|CEREBRAL CONTUSION W/ OPEN INTRACRANIAL WOUND W/ CONCUSSION|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|CEREBRAL CONTUSION WITH OPEN INTRACRANIAL WOUND WITH CONCUSSION|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|CORTEX (CEREBRAL) CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|OPN CORTX CONTUS-CONCUSS|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED |CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION |CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED CONCUSSION|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272967|T037|73413009|SNOMEDCT_US|CEREBRAL CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|CORTEX CONTUSION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272977|T037|209862001|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITH OPEN INTRACRANIAL WOUND|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND (FINDING)
C0272977|T037|209862001|SNOMEDCT_US|LACERATION OF CEREBRUM WITH OPEN INTRACRANIAL WOUND|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND (FINDING)
C0272977|T037|209862001|SNOMEDCT_US|LACERATION OF CEREBRUM WITH OPEN INTRACRANIAL WOUND |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND (FINDING)
C0272977|T037|209862001|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND (FINDING)
C0272977|T037|209862001|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND (FINDING)
C0272977|T037|209862001|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND (FINDING)
C0272977|T037|209862001|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND (FINDING)
C0272978|T037|111659005|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITH OPEN INTRACRANIAL WOUND, WITH STATE OF CONSCIOUSNESS UNSPECIFIED|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272978|T037|111659005|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272978|T037|111659005|SNOMEDCT_US|CORTEX LACER W OPN WOUND|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272978|T037|111659005|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITH OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272978|T037|111659005|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272978|T037|111659005|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272978|T037|111659005|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272978|T037|111659005|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272978|T037|111659005|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH STATE OF CONSCIOUSNESS UNSPECIFIED|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272978|T037|111659005|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH STATE OF CONSCIOUSNESS UNSPECIFIED|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-
C0272979|T037|209864000|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272979|T037|209864000|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND NO LOSS OF CONSCIOUSNESS|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272979|T037|209864000|SNOMEDCT_US|LACERATION OF CEREBRUM WITH OPEN INTRACRANIAL WOUND WITH NO LOSS OF CONSCIOUSNESS|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272979|T037|209864000|SNOMEDCT_US|LACERATION OF CEREBRUM WITH OPEN INTRACRANIAL WOUND WITH NO LOSS OF CONSCIOUSNESS |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272979|T037|209864000|SNOMEDCT_US|OPN CORTEX LACER-NO COMA|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272979|T037|209864000|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND NO LOSS OF CONSCIOUSNESS |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272979|T037|209864000|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272979|T037|209864000|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272979|T037|209864000|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|CORTEX (CEREBRAL) LACERATION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|LACERATION OF CEREBRUM WITH OPEN INTRACRANIAL WOUND WITH CONCUSSION|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|LACERATION OF CEREBRUM WITH OPEN INTRACRANIAL WOUND WITH CONCUSSION |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|OPN CORTX LACER-CONCUSS|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION |CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED CONCUSSION|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0272985|T037|69875006|SNOMEDCT_US|CEREBRAL CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|CORTEX LACERATION WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C1708044|T037||SNOMEDCT_US|FETAL BRAIN INJURY
C0270088|T037|206192007|SNOMEDCT_US|TENTORIAL TEAR|TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|TENTORIAL TEAR DUE TO BIRTH INJURY|TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|TENTORIAL TEAR DUE TO BIRTH TRAUMA|TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|TENTORIAL TEAR DUE TO BIRTH TRAUMA |TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|TEARS, TENTORIAL|TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|TENTORIAL TEARS|TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|TENTORIAL LACERATION DUE TO BIRTH TRAUMA|TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|TENTORIAL TEAR AS BIRTH TRAUMA|TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|TENTORIAL TEAR AS BIRTH TRAUMA |TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|TENTORIAL TEAR DUE TO BIRTH TRAUMA |TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|BIRTH; INJURY, TENTORIAL TEAR|TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C0270088|T037|206192007|SNOMEDCT_US|INJURY; BIRTH, TENTORIAL TEAR|TENTORIAL TEAR DUE TO BIRTH TRAUMA (DISORDER)
C2347482|T037||SNOMEDCT_US|PERINATAL BRAIN INJURY
C0478211|T037|213406009|SNOMEDCT_US|OTHER INTRACRANIAL INJURIES|[X]OTHER INTRACRANIAL INJURIES (DISORDER)
C0478211|T037|213406009|SNOMEDCT_US|OTHER INTRACRANIAL INJURY|[X]OTHER INTRACRANIAL INJURIES (DISORDER)
C0478211|T037|213406009|SNOMEDCT_US|[X]OTHER INTRACRANIAL INJURIES |[X]OTHER INTRACRANIAL INJURIES (DISORDER)
C0478211|T037|213406009|SNOMEDCT_US|[X]OTHER INTRACRANIAL INJURIES|[X]OTHER INTRACRANIAL INJURIES (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HAEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HAEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HEMORRHAGE NOS|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HEMORRHAGE, CRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMA, EPIDURAL, INTRACRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HEMATOMA, CRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMA, EPIDURAL, CRANIAL [DISEASE/FINDING]|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMORRHAGE, CRANIAL EPIDURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|CRANIAL EPIDURAL HEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMA, EPIDURAL, CRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|INTRACRANIAL EPIDURAL HEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMORRHAGE, CRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HAEMORRHAGE;EPIDURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HAEMORRHAGE;EPIDURAL;TRAUMATIC|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HAEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMORRHAGE NOS|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMATOMA |EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL INTRACRANIAL HEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL INTRACRANIAL HEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL INTRACRANIAL HEMORRHAGE |EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL INTRACRANIAL HAEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMORRHAGE |EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL INTRACRANIAL HEMATOMA |EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL INTRACRANIAL HAEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HAEMATOMA |EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL INTRACRANIAL HAEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL INTRACRANIAL HEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMORRHAGE, EXTRADURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|INTRACRANIAL EPIDURAL HAEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL BLEEDING|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HAEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EDH - EXTRADURAL HAEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EDH - EXTRADURAL HEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL; HEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL; HEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMA; EPIDURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMORRHAGE; EXTRADURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMORRHAGE, NOS|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HEMORRHAGE, NOS|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMORRHAGE [DUP] |EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|CRANIAL EPIDURAL HEMATOMAS|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|CRANIAL EPIDURAL HEMORRHAGES|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|CRANIAL EPIDURAL HEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|CRANIAL EXTRADURAL HEMATOMAS|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|CRANIAL EXTRADURAL HEMATOMA|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|CRANIAL EXTRADURAL HEMORRHAGES|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|CRANIAL EXTRADURAL HEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMATOMA, CRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMATOMA, INTRACRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMATOMAS, CRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMATOMAS, INTRACRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EPIDURAL HEMORRHAGES, CRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HEMATOMAS, CRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|EXTRADURAL HEMORRHAGES, CRANIAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMA, CRANIAL EPIDURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMA, CRANIAL EXTRADURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMA, INTRACRANIAL EPIDURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMAS, CRANIAL EPIDURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMAS, CRANIAL EXTRADURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMATOMAS, INTRACRANIAL EPIDURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMORRHAGE, CRANIAL EXTRADURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMORRHAGES, CRANIAL EPIDURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMORRHAGES, CRANIAL EXTRADURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|INTRACRANIAL EPIDURAL HEMATOMAS|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMORRHAGE;EPIDURAL|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|HEMORRHAGE;EPIDURAL;TRAUMATIC|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|TRAUMATIC EPIDURAL HEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0238154|T037|155392004|SNOMEDCT_US|TRAUMATIC EPIDURAL HAEMORRHAGE|EXTRADURAL HAEMATOMA (DISORDER)
C0452048|T037|210039000|SNOMEDCT_US|INTRACRANIAL INJURY WITH PROLONGED COMA|INTRACRANIAL INJURY WITH PROLONGED COMA (DISORDER)
C0452048|T037|210039000|SNOMEDCT_US|INTRACRANIAL INJURY WITH PROLONGED COMA |INTRACRANIAL INJURY WITH PROLONGED COMA (DISORDER)
C0452048|T037|210039000|SNOMEDCT_US|INTRACRANIAL INJURY UNSPECIFIED NATURE WITH PROLONGED COMA|INTRACRANIAL INJURY WITH PROLONGED COMA (DISORDER)
C0452048|T037|210039000|SNOMEDCT_US|INTRACRANIAL INJURY WITH PROLONGED COMA |INTRACRANIAL INJURY WITH PROLONGED COMA (DISORDER)
C0452048|T037|210039000|SNOMEDCT_US|INJURY; INTRACRANIAL, WITH PROLONGED COMA|INTRACRANIAL INJURY WITH PROLONGED COMA (DISORDER)
C0452048|T037|210039000|SNOMEDCT_US|INTRACRANIAL; INJURY, WITH PROLONGED COMA|INTRACRANIAL INJURY WITH PROLONGED COMA (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL INJURY|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL INJURY, UNSPECIFIED|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL INJURY OF UNSPECIFIED NATURE|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL INJURY OF UNSPECIFIED NATURE |[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY |[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INJURY;INTRACRANIAL|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL INJURY |[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL INJURY NOS|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL INJURY NOS |[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|[X]INTRACRANIAL INJURY, UNSPECIFIED|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|[X]INTRACRANIAL INJURY, UNSPECIFIED |[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INJURY; INTRACRANIAL|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL; INJURY|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0347535|T037|213407000|SNOMEDCT_US|INTRACRANIAL INJURY [AMBIGUOUS]|[X]INTRACRANIAL INJURY, UNSPECIFIED (DISORDER)
C0472391|T037|230763008|SNOMEDCT_US|TRAUMATIC CEREBRAL EDEMA|TRAUMATIC CEREBRAL EDEMA (DISORDER)
C0472391|T037|230763008|SNOMEDCT_US|TRAUMATIC CEREBRAL OEDEMA|TRAUMATIC CEREBRAL EDEMA (DISORDER)
C0472391|T037|230763008|SNOMEDCT_US|TRAUMATIC CEREBRAL EDEMA NOS|TRAUMATIC CEREBRAL EDEMA (DISORDER)
C0472391|T037|230763008|SNOMEDCT_US|CEREBRAL EDEMA TRAUMATIC|TRAUMATIC CEREBRAL EDEMA (DISORDER)
C0472391|T037|230763008|SNOMEDCT_US|TRAUMATIC CEREBRAL EDEMA |TRAUMATIC CEREBRAL EDEMA (DISORDER)
C0472391|T037|230763008|SNOMEDCT_US|TRAUMATIC CEREBRAL OEDEMA |TRAUMATIC CEREBRAL EDEMA (DISORDER)
C0472391|T037|230763008|SNOMEDCT_US|TRAUMATIC CEREBRAL EDEMA |TRAUMATIC CEREBRAL EDEMA (DISORDER)
C0472391|T037|230763008|SNOMEDCT_US|EDEMA; BRAIN, TRAUMATIC|TRAUMATIC CEREBRAL EDEMA (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|TRAUMATIC SUBARACHNOID HAEMORRHAGE|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|TRAUMATIC SUBARACHNOID HEMORRHAGE|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|HEMORRHAGE, POST-TRAUMATIC SUBARACHNOID|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|HEMORRHAGES, POST-TRAUMATIC SUBARACHNOID|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|POST TRAUMATIC SUBARACHNOID HEMORRHAGE|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|POST-TRAUMATIC SUBARACHNOID HEMORRHAGES|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE, POST-TRAUMATIC|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|SUBARACHNOID HEMORRHAGES, POST-TRAUMATIC|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|HEMORRHAGE, TRAUMATIC SUBARACHNOID|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE, TRAUMATIC|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|SUBARACHNOID HEMORRHAGES, TRAUMATIC|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|TRAUMATIC SUBARACHNOID HEMORRHAGES|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|POST-TRAUMATIC SUBARACHNOID HEMORRHAGE|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE, TRAUMATIC [DISEASE/FINDING]|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|TRAUMATIC SUBARACHNOID HEMORRHAGE NOS|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|TRAUMATIC SUBARACHNOID HEMORRHAGE |TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|TRAUMATIC SUBARACHNOID INTRACRANIAL HEMORRHAGE |TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|SUBARACHNOID HAEMORRHAGE FOLLOWING INJURY|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|TRAUMATIC SUBARACHNOID HAEMORRHAGE |TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|TRAUMATIC SUBARACHNOID INTRACRANIAL HAEMORRHAGE|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|TRAUMATIC SUBARACHNOID INTRACRANIAL HEMORRHAGE|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|HEMORRHAGE; SUBARACHNOID, TRAUMATIC|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C0475073|T037|157323000|SNOMEDCT_US|SUBARACHNOID; HEMORRHAGE, TRAUMATIC|TRAUMATIC SUBARACHNOID HAEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|TRAUMATIC SUBDURAL HAEMORRHAGE|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|TRAUMATIC SUBDURAL HEMORRHAGE|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|HEAD INJURY WITH SUBDURAL HEMORRHAGE|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|HEAD INJURY WITH SUBDURAL HEMORRHAGE |TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|HAEMORRHAGE;SUBDURAL;TRAUMATIC|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|TRAUMATIC SUBDURAL HEMORRHAGE NOS|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|TRAUMATIC SUBDURAL INTRACRANIAL HEMORRHAGE|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|TRAUMATIC SUBDURAL INTRACRANIAL HAEMORRHAGE|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|TRAUMATIC SUBDURAL INTRACRANIAL HEMORRHAGE |TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|TRAUMATIC SUBDURAL HEMORRHAGE |TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|SUBDURAL HAEMORRHAGE FOLLOWING INJURY|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|SUBDURAL HEMORRHAGE FOLLOWING INJURY|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|HEMORRHAGE; SUBDURAL, TRAUMATIC|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|SUBDURAL; HEMORRHAGE, TRAUMATIC|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C1367166|T037|209987007|SNOMEDCT_US|HEMORRHAGE;SUBDURAL;TRAUMATIC|TRAUMATIC SUBDURAL HEMORRHAGE (DISORDER)
C2832047|T037||SNOMEDCT_US|DIFFUSE TRAUMATIC BRAIN INJURY
C2832047|T037||SNOMEDCT_US|DIFFUSE TRAUMATIC BRAIN INJURY NOS
C2832047|T037||SNOMEDCT_US|BRAIN INJURY TRAUMATIC DIFFUSE
C2832047|T037||SNOMEDCT_US|DIFFUSE TRAUMATIC BRAIN INJURY 
C2832052|T037||SNOMEDCT_US|FOCAL TRAUMATIC BRAIN INJURY
C2832052|T037||SNOMEDCT_US|FOCAL TRAUMATIC BRAIN INJURY 
C2832052|T037||SNOMEDCT_US|BRAIN INJURY TRAUMATIC FOCAL
C2977736|T037||SNOMEDCT_US|OTHER SPECIFIED INTRACRANIAL INJURIES
C0272936|T037|28188001|SNOMEDCT_US|INTRACRANIAL INJURY UNSPECIFIED NATURE WITH OPEN INTRACRANIAL WOUND |BRAIN INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0272936|T037|28188001|SNOMEDCT_US|INTRACRANIAL INJURY UNSPECIFIED NATURE WITH OPEN INTRACRANIAL WOUND|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0272936|T037|28188001|SNOMEDCT_US|INTRACRANIAL INJURY OF UNSPECIFIED NATURE WITH OPEN INTRACRANIAL WOUND|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0272936|T037|28188001|SNOMEDCT_US|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND |BRAIN INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0272936|T037|28188001|SNOMEDCT_US|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0272936|T037|28188001|SNOMEDCT_US|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND, NOS|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C2118964|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH NO LOSS OF CONSCIOUSNESS 
C2118964|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH NO LOSS OF CONSCIOUSNESS
C2118964|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH NO LOC
C2118965|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH BRIEF (< 1 HR) LOSS OF CONSCIOUSNESS 
C2118965|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY BRIEF (UNDER 1 HR) UNCONSCIOUSNESS
C2118965|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH BRIEF (< 1 HR) LOSS OF CONSCIOUSNESS
C2118965|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH BRIEF (< 1 HR) LOC
C2118965|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH BRIEF (UNDER 1 HR) UNCONSCIOUSNESS
C2118966|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH MODERATE (1-24 HRS) LOSS OF CONSCIOUSNESS 
C2118966|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY MODERATE (1-24 HRS) UNCONSCIOUSNESS
C2118966|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH MODERATE (1-24 HRS) LOSS OF CONSCIOUSNESS
C2118966|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH MODERATE (1-24 HRS) LOC
C2118966|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH MODERATE (1-24 HRS) UNCONSCIOUSNESS
C2118967|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH PROLONGED (> 24 HRS) LOSS OF CONSCIOUSNESS WITH RETURN TO PRIOR LEVEL OF CONSCIOUSNESS 
C2118967|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY LOSS OF CONSCIOUSNESS >24 HR THEN RETURN TO PRIOR LEVEL
C2118967|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH PROLONGED (> 24 HRS) LOSS OF CONSCIOUSNESS WITH RETURN TO PRIOR LEVEL OF CONSCIOUSNESS
C2118967|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOC OVER 24 HR, THEN RETURN TO PRIOR LEVEL
C2118968|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH PROLONGED (> 24 HRS) LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRIOR LEVEL OF CONSCIOUSNESS
C2118968|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY LOSS OF CONSCIOUSNESS > 24 HR WITHOUT RETURN TO PRIOR LEVEL
C2118968|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH PROLONGED (> 24 HRS) LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRIOR LEVEL OF CONSCIOUSNESS 
C2118968|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOC OVER 24 HOURS WITHOUT RETURN TO PRIOR LEVEL
C2118969|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH UNCONSCIOUSNESS OF UNSPECIFIED DURATION 
C2118969|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH UNCONSCIOUSNESS OF UNSPECIFIED DURATION
C2118970|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH CONCUSSION 
C2118970|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH CONCUSSION
C2832671|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITHOUT LOSS OF CONSCIOUSNESS
C2832675|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 30 MINUTES OR LESS
C2832679|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 31 MINUTES TO 59 MINUTES
C2832683|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 1 HOUR TO 5 HOURS 59 MINUTES
C2832687|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF 6 HOURS TO 24 HOURS
C2832691|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITH RETURN TO PRE-EXISTING CONSCIOUS LEVEL
C2832695|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL WITH PATIENT SURVIVING
C2832699|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF ANY DURATION WITH DEATH DUE TO BRAIN INJURY PRIOR TO REGAINING CONSCIOUSNESS
C2832703|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF ANY DURATION WITH DEATH DUE TO OTHER CAUSE PRIOR TO REGAINING CONSCIOUSNESS
C2832707|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION
C0435306|T037|111617009|SNOMEDCT_US|OPEN FRACTURE OF SKULL WITH INTRACRANIAL INJURY |OPEN SKULL FRACTURE WITH INTRACRANIAL INJURY (DISORDER)
C0435306|T037|111617009|SNOMEDCT_US|OPEN SKULL FRACTURE WITH INTRACRANIAL INJURY|OPEN SKULL FRACTURE WITH INTRACRANIAL INJURY (DISORDER)
C0435306|T037|111617009|SNOMEDCT_US|OPEN FRACTURE OF SKULL WITH INTRACRANIAL INJURY|OPEN SKULL FRACTURE WITH INTRACRANIAL INJURY (DISORDER)
C0435306|T037|111617009|SNOMEDCT_US|OPEN FRACTURE OF SKULL NOS WITH INTRACRANIAL INJURY|OPEN SKULL FRACTURE WITH INTRACRANIAL INJURY (DISORDER)
C0435306|T037|111617009|SNOMEDCT_US|OPEN FRACTURE OF SKULL NOS WITH INTRACRANIAL INJURY |OPEN SKULL FRACTURE WITH INTRACRANIAL INJURY (DISORDER)
C0435306|T037|111617009|SNOMEDCT_US|OPEN SKULL FRACTURE WITH INTRACRANIAL INJURY |OPEN SKULL FRACTURE WITH INTRACRANIAL INJURY (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|CLOSED HEAD INJURY|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|HEAD INJURIES, CLOSED|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|HEAD INJURY, CLOSED|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|CLOSED HEAD INJURIES|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|HEAD INJ NONPENETRATING|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|INJ CLOSED HEAD|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|CLOSED HEAD INJ|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|HEAD INJ CLOSED|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|CLOSED HEAD TRAUMA|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|CLOSED HEAD TRAUMAS|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|HEAD TRAUMAS, CLOSED|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|TRAUMA, CLOSED HEAD|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|TRAUMAS, CLOSED HEAD|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|NONPENETRATING HEAD INJURIES|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|NONPENETRATING HEAD INJURY|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|HEAD INJURIES, NONPENETRATING|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|HEAD TRAUMA, CLOSED|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|HEAD INJURIES, CLOSED [DISEASE/FINDING]|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|INJURIES, CLOSED HEAD|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|HEAD INJURY, NONPENETRATING|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|CLOSED INJURY OF HEAD|CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|CLOSED INJURY OF HEAD |CLOSED INJURY OF HEAD (DISORDER)
C0085094|T037|451000119106|SNOMEDCT_US|INJURY;CLOSED HEAD|CLOSED INJURY OF HEAD (DISORDER)
C3506613|T037||SNOMEDCT_US|INJURY OF INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION 
C3506613|T037||SNOMEDCT_US|INJURY OF INTERNAL CAROTID ARTERY, INTRACRANIAL PORTION
C3506613|T037||SNOMEDCT_US|INJURY INTERNAL CAROTID ARTERY INTRACRANIAL PORTION
C3506611|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOC WITH DEATH DUE TO BRAIN INJURY PRIOR TO REGAINING CONSCIOUSNESS 
C3506611|T037||SNOMEDCT_US|UNSPECIFIED INTRACRANIAL INJURY WITH LOC WITH DEATH DUE TO BRAIN INJURY PRIOR TO REGAINING CONSCIOUSNESS
C3506611|T037||SNOMEDCT_US|UNSPEC INTRACRANIAL INJURY LOC W/ DEATH D/T BRAIN INJURY PRIOR TO REGAIN CONSC
C3506612|T037||SNOMEDCT_US|UNSPEC INTRACRANIAL INJURY LOC W/ DEATH D/T OTHER CAUSE PRIOR TO REGAIN CONSC 
C3506612|T037||SNOMEDCT_US|UNSPEC INTRACRANIAL INJURY LOC W/ DEATH D/T OTHER CAUSE PRIOR TO REGAIN CONSC
C0161401|T037|56311003|SNOMEDCT_US|INJURY OF VISUAL CORTEX|TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|INJURY OF VISUAL CORTEX |TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|INJURY TO THE VISUAL CORTEX|TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|INJURY TO VISUAL CORTEX|TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|INJURY OF VISUAL CORTEX NOS|TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|TRAUMATIC INJURY OF VISUAL CORTEX|TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|TRAUMATIC INJURY OF VISUAL CORTEX |TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|VISUAL CORTEX INJURY|TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|VISUAL CORTEX INJURY |TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|CORTEX; INJURY, VISUAL|TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|INJURY; CORTEX, VISUAL|TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|INJURY; VISUAL CORTEX|TRAUMATIC INJURY OF VISUAL CORTEX
C0161401|T037|56311003|SNOMEDCT_US|VISUAL CORTEX; INJURY|TRAUMATIC INJURY OF VISUAL CORTEX
C0270802|T037|28534004|SNOMEDCT_US|SPASTIC PARALYSIS DUE TO INTRACRANIAL BIRTH INJURY|SPASTIC PARALYSIS DUE TO INTRACRANIAL BIRTH INJURY (DISORDER)
C0270802|T037|28534004|SNOMEDCT_US|SPASTIC PARALYSIS DUE TO INTRACRANIAL BIRTH INJURY |SPASTIC PARALYSIS DUE TO INTRACRANIAL BIRTH INJURY (DISORDER)
C0475075|T037|269146000|SNOMEDCT_US|CLOSED TRAUMATIC SUBARACHNOID HAEMORRHAGE|CLOSED TRAUMATIC SUBARACHNOID HEMORRHAGE (DISORDER)
C0475075|T037|269146000|SNOMEDCT_US|CLOSED TRAUMATIC SUBARACHNOID HEMORRHAGE|CLOSED TRAUMATIC SUBARACHNOID HEMORRHAGE (DISORDER)
C0475075|T037|269146000|SNOMEDCT_US|CLOSED TRAUMATIC SUBARACHNOID HEMORRHAGE |CLOSED TRAUMATIC SUBARACHNOID HEMORRHAGE (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL HAEMORRHAGE DUE TO BIRTH INJURY|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL HEMORRHAGE DUE TO BIRTH INJURY|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL HEMORRHAGE DUE TO BIRTH TRAUMA|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL HEMORRHAGE DUE TO BIRTH TRAUMA |SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL INTRACRANIAL HEMORRHAGE DUE TO BIRTH TRAUMA |SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL INTRACRANIAL HAEMORRHAGE DUE TO BIRTH TRAUMA|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL INTRACRANIAL HEMORRHAGE DUE TO BIRTH TRAUMA|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL HEMORRHAGE DUE TO BIRTH TRAUMA |SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL HAEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA |SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0473821|T037|206190004|SNOMEDCT_US|SUBDURAL HAEMORRHAGE DUE TO BIRTH TRAUMA|SUBDURAL HEMORRHAGE UNSPECIFIED, DUE TO BIRTH TRAUMA (DISORDER)
C0475054|T037|209976004|SNOMEDCT_US|OPEN TRAUMATIC EXTRADURAL HAEMORRHAGE|OPEN TRAUMATIC EXTRADURAL HEMORRHAGE (DISORDER)
C0475054|T037|209976004|SNOMEDCT_US|OPEN TRAUMATIC EXTRADURAL HEMORRHAGE|OPEN TRAUMATIC EXTRADURAL HEMORRHAGE (DISORDER)
C0475054|T037|209976004|SNOMEDCT_US|OPEN TRAUMATIC EXTRADURAL HEMORRHAGE |OPEN TRAUMATIC EXTRADURAL HEMORRHAGE (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|CLOSED TRAUMATIC SUBDURAL INTRACRANIAL HAEMORRHAGE|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|CLOSED TRAUMATIC SUBDURAL INTRACRANIAL HEMORRHAGE|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|CLOSED TRAUMATIC SUBDURAL INTRACRANIAL HEMORRHAGE |SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|CLOSED TRAUMATIC SUBDURAL HEMORRHAGE |SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|SUBDURAL HAEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND |SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|HEAD INJURY - SUBDURAL HEMORRHAGE WITHOUT OPEN INTRACRANIAL WOUND|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|SUBDURAL HEMORRHAGE FOLLOWING HEAD INJURY WITHOUT OPEN INTRACRANIAL WOUND |SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|SUBDURAL HEMORRHAGE FOLLOWING HEAD INJURY WITHOUT OPEN INTRACRANIAL WOUND|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|CLOSED TRAUMATIC SUBDURAL HAEMORRHAGE|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475061|T037|7602002|SNOMEDCT_US|CLOSED TRAUMATIC SUBDURAL HEMORRHAGE|SUBDURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|HEMATOMA, TRAUMATIC SUBDURAL|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|HEMATOMAS, TRAUMATIC SUBDURAL|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|SUBDURAL HEMATOMAS, TRAUMATIC|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|TRAUMATIC SUBDURAL HEMATOMA|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|TRAUMATIC SUBDURAL HEMATOMAS|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|HAEMATOMA;SUBDURAL;TRAUMATIC|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|SUBDURAL HEMATOMA, TRAUMATIC|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|TRAUMATIC SUBDURAL HAEMATOMA|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|TRAUMATIC SUBDURAL HAEMATOMA |TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|TRAUMATIC SUBDURAL HEMATOMA |TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|TRAUMATIC SUBDURAL HEMATOMA |TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|SUBDURAL HEMATOMA - TRAUMATIC|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|SUBDURAL HEMATOMA (TRAUMATIC)|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|SUBDURAL HAEMATOMA (TRAUMATIC)|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0475059|T037|262951009|SNOMEDCT_US|HEMATOMA;SUBDURAL;TRAUMATIC|TRAUMATIC SUBDURAL HEMATOMA (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY NERVE INJURY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMATIC OLFACTORY NERVE INJURY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY NERVE INJURY |INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMATIC OLFACTORY NERVE INJURY |INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY OF OLFACTORY [1ST ] NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURIES, OLFACTORY NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|NERVE TRAUMA, OLFACTORY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMA, OLFACTORY NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMATIC OLFACTORY NEUROPATHIES|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|FIRST NERVE PALSY, TRAUMATIC|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|PALSY, TRAUMATIC FIRST-NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY NERVE INJURIES|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|FIRST-NERVE TRAUMAS|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|PALSIES, TRAUMATIC FIRST-NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMATIC FIRST-NERVE PALSIES|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMAS, FIRST-NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|NERVE INJURY, OLFACTORY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|NERVE TRAUMAS, OLFACTORY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|NEUROPATHY, TRAUMATIC OLFACTORY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMATIC FIRST NERVE PALSY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|FIRST NERVE TRAUMA|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY NEUROPATHIES, TRAUMATIC|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMATIC OLFACTORY NEUROPATHY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY, OLFACTORY NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|NERVE INJURIES, OLFACTORY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMA, FIRST-NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMAS, OLFACTORY NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|FIRST-NERVE PALSIES, TRAUMATIC|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY NERVE TRAUMAS|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|NEUROPATHIES, TRAUMATIC OLFACTORY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|CRANIAL NERVE I INJURY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|FIRST CRANIAL NERVE INJURY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY, FIRST CRANIAL NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY NEUROPATHY, TRAUMATIC|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|FIRST-NERVE TRAUMA|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY NERVE INJURIES [DISEASE/FINDING]|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|TRAUMATIC FIRST-NERVE PALSY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY NERVE TRAUMA|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|FIRST CRANIAL NERVE INJURIES|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|FIRST-NERVE PALSY, TRAUMATIC|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY, CRANIAL NERVE I|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY (1ST) NERVE INJURY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|OLFACTORY NERVE INJURY |INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY OF FIRST CRANIAL NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY OF OLFACTORY NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY TO OLFACTORY NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY OF OLFACTORY NERVE |INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY; OLFACTORY NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|N.OLFACTORIUS; INJURY|INJURY OF OLFACTORY NERVE (DISORDER)
C0273487|T037|72758005|SNOMEDCT_US|INJURY TO 1ST CRANIAL NERVE|INJURY OF OLFACTORY NERVE (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|SUBARACHNOID HAEMORRHAGE DUE TO BIRTH INJURY|SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY|SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|INTRACRANIAL SUBARACHNOID HAEMORRHAGE DUE TO BIRTH INJURY|SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY |SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|INTRACRANIAL SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY|SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|INTRACRANIAL SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY |SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|BIRTH TRAUMA SUBARACHNOID HEMORRHAGE|SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE DUE TO BIRTH TRAUMA|SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE DUE TO BIRTH TRAUMA |SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0475592|T037|206399009|SNOMEDCT_US|BIRTH; INJURY, SUBARACHNOID HEMORRHAGE|SUBARACHNOID HEMORRHAGE DUE TO BIRTH INJURY (DISORDER)
C0474996|T037|262719002|SNOMEDCT_US|TRAUMATIC SPINAL SUBARACHNOID HEMORRHAGE|TRAUMATIC SPINAL SUBARACHNOID HEMORRHAGE (DISORDER)
C0474996|T037|262719002|SNOMEDCT_US|HEMORRHAGE SUBARACHNOID TRAUMATIC SPINAL|TRAUMATIC SPINAL SUBARACHNOID HEMORRHAGE (DISORDER)
C0474996|T037|262719002|SNOMEDCT_US|TRAUMATIC SPINAL SUBARACHNOID HEMORRHAGE |TRAUMATIC SPINAL SUBARACHNOID HEMORRHAGE (DISORDER)
C0474996|T037|262719002|SNOMEDCT_US|TRAUMATIC SPINAL SUBARACHNOID HAEMORRHAGE|TRAUMATIC SPINAL SUBARACHNOID HEMORRHAGE (DISORDER)
C0474996|T037|262719002|SNOMEDCT_US|TRAUMATIC SPINAL SUBARACHNOID HEMORRHAGE |TRAUMATIC SPINAL SUBARACHNOID HEMORRHAGE (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|CRUSHING INJURY OF HEAD|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|CRUSHING INJURY OF HEAD, PART UNSPECIFIED|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|CRUSHING INJURY OF SKULL AND INTRACRANIAL CONTENTS|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|CRUSH INJURY OF HEAD |[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|CRUSH INJURY HEAD|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|CRUSH INJURY OF HEAD|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED |[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|CRUSHING INJURY OF SKULL AND INTRACRANIAL CONTENTS |[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|CRUSHING INJURY; HEAD|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0433070|T037|213409002|SNOMEDCT_US|HEAD; CRUSHING INJURY|[X]CRUSHING INJURY OF HEAD, PART UNSPECIFIED (DISORDER)
C0272937|T037|111655004|SNOMEDCT_US|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS -RETIRED-|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0272937|T037|111655004|SNOMEDCT_US|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0272937|T037|111655004|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS |BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0272937|T037|111655004|SNOMEDCT_US|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS |BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0272937|T037|111655004|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433774|T037|210030001|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433774|T037|210030001|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433783|T037|210021009|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433783|T037|210021009|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL |INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433769|T037|210025000|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0433769|T037|210025000|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0433776|T037|210032009|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433776|T037|210032009|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433784|T037|210022002|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS STATE|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS STATE (DISORDER)
C0433784|T037|210022002|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS STATE |INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS STATE (DISORDER)
C0433786|T037|210024001|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0433786|T037|210024001|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED |INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0433780|T037|269150007|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS |INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0433780|T037|269150007|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0433785|T037|210023007|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION |INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433785|T037|210023007|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION (DISORDER)
C0433775|T037|210031002|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433775|T037|210031002|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0433782|T037|210020005|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS |INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0433782|T037|210020005|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0433773|T037|210029006|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0433773|T037|210029006|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0433779|T037|210017002|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS |INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0433779|T037|210017002|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, UNSPECIFIED STATE OF CONSCIOUSNESS (DISORDER)
C0272938|T037|210027008|SNOMEDCT_US|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND NO LOSS OF CONSCIOUSNESS|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272938|T037|210027008|SNOMEDCT_US|HEAD INJURY WITH OPEN INTRACRANIAL WOUND WITH NO LOSS OF CONSCIOUSNESS |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272938|T037|210027008|SNOMEDCT_US|HEAD INJURY WITH OPEN INTRACRANIAL WOUND WITH NO LOSS OF CONSCIOUSNESS|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272938|T037|210027008|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272938|T037|210027008|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0272938|T037|210027008|SNOMEDCT_US|BRAIN INJURY WITH OPEN INTRACRANIAL WOUND AND NO LOSS OF CONSCIOUSNESS |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH NO LOSS OF CONSCIOUSNESS (DISORDER)
C0433778|T037|210016006|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND |INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND (DISORDER)
C0433778|T037|210016006|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND (DISORDER)
C0433781|T037|210019004|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS (DISORDER)
C0433781|T037|210019004|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS |INTRACRANIAL INJURY NOS WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS (DISORDER)
C0433777|T037|210033004|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0433777|T037|210033004|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED (DISORDER)
C0433772|T037|210028003|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOURS LOSS OF CONSCIOUSNESS |INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0433772|T037|210028003|SNOMEDCT_US|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOURS LOSS OF CONSCIOUSNESS|INTRACRANIAL INJURY NOS WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0272925|T037|54355006|SNOMEDCT_US|INTRACRANIAL INJURY WITHOUT SKULL FRACTURE|INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE (DISORDER)
C0272925|T037|54355006|SNOMEDCT_US|HEAD INJURY UNSPECIFIED INTRACRANIAL INJURY WITHOUT SKULL FRACTURE|INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE (DISORDER)
C0272925|T037|54355006|SNOMEDCT_US|INTRACRANIAL INJURY WITHOUT SKULL FRACTURE |INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE (DISORDER)
C0272925|T037|54355006|SNOMEDCT_US|HEAD INJURY, WITHOUT SKULL FRACTURE|INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE (DISORDER)
C0272925|T037|54355006|SNOMEDCT_US|INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE |INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE (DISORDER)
C0272925|T037|54355006|SNOMEDCT_US|INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE|INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE (DISORDER)
C0272925|T037|54355006|SNOMEDCT_US|HEAD INJURY, NOS, WITHOUT SKULL FRACTURE|INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE (DISORDER)
C0272925|T037|54355006|SNOMEDCT_US|INTRACRANIAL INJURY, NOS, WITHOUT SKULL FRACTURE|INTRACRANIAL INJURY, WITHOUT SKULL FRACTURE (DISORDER)
C0558400|T037|269338005|SNOMEDCT_US|H'GE - CEREBRAL TRAUMA|H'GE - CEREBRAL TRAUMA
C0558400|T037|269338005|SNOMEDCT_US|CEREBRAL TRAUMA|H'GE - CEREBRAL TRAUMA
C0558400|T037|269338005|SNOMEDCT_US|CEREBRAL TRAUMA |H'GE - CEREBRAL TRAUMA
C0558400|T037|269338005|SNOMEDCT_US|CEREBRAL TRAUMA |H'GE - CEREBRAL TRAUMA
C0411045|T037|240312009|SNOMEDCT_US|CEREBRAL INJURY DUE TO BIRTH TRAUMA|CEREBRAL INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0411045|T037|240312009|SNOMEDCT_US|CEREBRAL INJURY DUE TO BIRTH TRAUMA |CEREBRAL INJURY DUE TO BIRTH TRAUMA (DISORDER)
C0433855|T037|262692002|SNOMEDCT_US|BRAIN INJURY TRAUMATIC BURST LOBE|BURST LOBE OF BRAIN (DISORDER)
C0433855|T037|262692002|SNOMEDCT_US|BURST LOBE OF BRAIN|BURST LOBE OF BRAIN (DISORDER)
C0433855|T037|262692002|SNOMEDCT_US|BURST LOBE OF BRAIN |BURST LOBE OF BRAIN (DISORDER)
C0433855|T037|262692002|SNOMEDCT_US|BURST LOBE OF BRAIN |BURST LOBE OF BRAIN (DISORDER)
C0442857|T037|264534009|SNOMEDCT_US|HYPOTHALAMIC INJURY|HYPOTHALAMIC INJURY (DISORDER)
C0442857|T037|264534009|SNOMEDCT_US|HYPOTHALAMIC INJURY |HYPOTHALAMIC INJURY (DISORDER)
C0442857|T037|264534009|SNOMEDCT_US|HYPOTHALAMIC INJURY |HYPOTHALAMIC INJURY (DISORDER)
C0456045|T037|275361004|SNOMEDCT_US|BRAIN LACERATION TENTORIAL|TENTORIAL LACERATION (DISORDER)
C0456045|T037|275361004|SNOMEDCT_US|TENTORIAL BRAIN LACERATION|TENTORIAL LACERATION (DISORDER)
C0456045|T037|275361004|SNOMEDCT_US|TENTORIAL BRAIN LACERATION |TENTORIAL LACERATION (DISORDER)
C0456045|T037|275361004|SNOMEDCT_US|TENTORIAL LACERATION|TENTORIAL LACERATION (DISORDER)
C0456045|T037|275361004|SNOMEDCT_US|TENTORIAL LACERATION |TENTORIAL LACERATION (DISORDER)
C0435236|T037|207687004|SNOMEDCT_US|CLOSED FRACTURE OF SKULL VAULT WITH INTRACRANIAL INJURY|CLOSED FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435236|T037|207687004|SNOMEDCT_US|CLOSED FRACTURE OF SKULL VAULT WITH INTRACRANIAL INJURY |CLOSED FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435236|T037|207687004|SNOMEDCT_US|CLOSED FRACTURE OF VAULT OF SKULL WITH INTRACRANIAL INJURY |CLOSED FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435236|T037|207687004|SNOMEDCT_US|CLOSED FRACTURE OF VAULT OF SKULL WITH INTRACRANIAL INJURY|CLOSED FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435236|T037|207687004|SNOMEDCT_US|FRACTURE OF VAULT OF SKULL, CLOSED WITH INTRACRANIAL INJURY|CLOSED FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435236|T037|207687004|SNOMEDCT_US|CLOSED FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY|CLOSED FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435236|T037|207687004|SNOMEDCT_US|CLOSED FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY |CLOSED FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435223|T037|207705002|SNOMEDCT_US|OPEN FRACTURE OF SKULL VAULT WITH INTRACRANIAL INJURY|OPEN FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435223|T037|207705002|SNOMEDCT_US|OPEN FRACTURE OF SKULL VAULT WITH INTRACRANIAL INJURY |OPEN FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435223|T037|207705002|SNOMEDCT_US|OPEN FRACTURE OF VAULT OF SKULL WITH INTRACRANIAL INJURY|OPEN FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435223|T037|207705002|SNOMEDCT_US|OPEN FRACTURE OF VAULT OF SKULL WITH INTRACRANIAL INJURY |OPEN FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435223|T037|207705002|SNOMEDCT_US|FRACTURE OF VAULT OF SKULL, OPEN WITH INTRACRANIAL INJURY|OPEN FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435223|T037|207705002|SNOMEDCT_US|OPEN FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY|OPEN FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435223|T037|207705002|SNOMEDCT_US|OPEN FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY |OPEN FRACTURE VAULT OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|HEAD INJURY WITH INTRACRANIAL HEMORRHAGE|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|HEAD INJURY WITH INTRACRANIAL HEMORRHAGE |TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|HEMORRHAGE, TRAUMATIC INTRACRANIAL|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|HEMORRHAGES, TRAUMATIC INTRACRANIAL|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|INTRACRANIAL HEMORRHAGE, TRAUMATIC|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|INTRACRANIAL HEMORRHAGES, TRAUMATIC|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|TRAUMATIC INTRACRANIAL HEMORRHAGES|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|INTRACRANIAL HEMORRHAGE, TRAUMATIC [DISEASE/FINDING]|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|TRAUMATIC INTRACRANIAL HEMORRHAGE|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|HEMORRHAGE, INTRACRANIAL, TRAUMATIC|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|INTRACRANIAL HEMORRHAGE FOLLOWING INJURY|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|TRAUMATIC INTRACRANIAL HAEMORRHAGE |TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|INTRACRANIAL HEMORRHAGE FOLLOWING INJURY |TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|TRAUMATIC INTRACRANIAL HEMORRHAGE |TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|TRAUMATIC INTRACRANIAL HAEMORRHAGE|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|INTRACRANIAL HAEMORRHAGE FOLLOWING INJURY|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|TRAUMATIC INTRACRANIAL BLEEDING|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|TRAUMATIC INTRACRANIAL HAEMORRHAGE NOS|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|TRAUMATIC INTRACRANIAL HEMORRHAGE NOS|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|HEMORRHAGE; INTRACRANIAL, TRAUMATIC|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|HEMORRHAGE; TRAUMATIC, INTRACRANIAL|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|INTRACRANIAL; HEMORRHAGE, TRAUMATIC|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|TRAUMATIC; HEMORRHAGE, INTRACRANIAL|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C0273058|T037|269145001|SNOMEDCT_US|INTRACRANIAL HEMORRHAGE FOLLOWING INJURY, NOS|TRAUMATIC INTRACRANIAL HEMORRHAGE (DISORDER)
C1264285|T037|127297005|SNOMEDCT_US|INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS |INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS (DISORDER)
C1264285|T037|127297005|SNOMEDCT_US|INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS|INTRACRANIAL INJURY WITH LOSS OF CONSCIOUSNESS (DISORDER)
C0435249|T037|111607004|SNOMEDCT_US|OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY |OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435249|T037|111607004|SNOMEDCT_US|OPEN BASILAR SKULL FRACTURE WITH INTRACRANIAL INJURY|OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435249|T037|111607004|SNOMEDCT_US|OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY|OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435249|T037|111607004|SNOMEDCT_US|OPEN FRACTURE BASE OF SKULL WITH INTRACRANIAL INJURY |OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435249|T037|111607004|SNOMEDCT_US|OPEN FRACTURE BASE OF SKULL WITH INTRACRANIAL INJURY|OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435249|T037|111607004|SNOMEDCT_US|FRACTURE OF BASE OF SKULL, OPEN WITH INTRACRANIAL INJURY|OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435249|T037|111607004|SNOMEDCT_US|OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY |OPEN FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435262|T037|111603000|SNOMEDCT_US|CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY |CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435262|T037|111603000|SNOMEDCT_US|CLOSED BASILAR SKULL FRACTURE WITH INTRACRANIAL INJURY|CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435262|T037|111603000|SNOMEDCT_US|CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY|CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435262|T037|111603000|SNOMEDCT_US|CLOSED FRACTURE BASE OF SKULL WITH INTRACRANIAL INJURY |CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435262|T037|111603000|SNOMEDCT_US|CLOSED FRACTURE BASE OF SKULL WITH INTRACRANIAL INJURY|CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435262|T037|111603000|SNOMEDCT_US|FRACTURE OF BASE OF SKULL, CLOSED WITH INTRACRANIAL INJURY|CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0435262|T037|111603000|SNOMEDCT_US|CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY |CLOSED FRACTURE OF BASE OF SKULL WITH INTRACRANIAL INJURY (DISORDER)
C0273098|T037|43216008|SNOMEDCT_US|CLOSED TRAUMATIC EXTRADURAL HEMORRHAGE|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0273098|T037|43216008|SNOMEDCT_US|CLOSED TRAUMATIC EXTRADURAL HAEMORRHAGE|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0273098|T037|43216008|SNOMEDCT_US|CLOSED TRAUMATIC EXTRADURAL HEMORRHAGE |EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0273098|T037|43216008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND |EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0273098|T037|43216008|SNOMEDCT_US|HEAD INJURY - WITH EXTRADURAL HEMORRHAGE, WITHOUT OPEN INTRACRANIAL WOUND|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0273098|T037|43216008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0273098|T037|43216008|SNOMEDCT_US|EXTRADURAL HAEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0273098|T037|43216008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND |EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND (DISORDER)
C0272499|T037|61642003|SNOMEDCT_US|MULTIPLE OPEN FRACTURES OF SKULL OR FACE WITH SUBARACHNOID, SUBDURAL, OR EXTRADURAL HEMORRHAGE |MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HEMORRHAGE (DISORDER)
C0272499|T037|61642003|SNOMEDCT_US|MULTI SKULL/FACE FRACTURES OPEN W/ SUBARACHNOID, SUBDURAL, EXTRADURAL HEMORRHAGE|MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HEMORRHAGE (DISORDER)
C0272499|T037|61642003|SNOMEDCT_US|MULTIPLE OPEN FRACTURES OF SKULL OR FACE WITH SUBARACHNOID, SUBDURAL, OR EXTRADURAL HEMORRHAGE|MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HEMORRHAGE (DISORDER)
C0272499|T037|61642003|SNOMEDCT_US|MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HAEMORRHAGE|MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HEMORRHAGE (DISORDER)
C0272499|T037|61642003|SNOMEDCT_US|MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HEMORRHAGE |MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HEMORRHAGE (DISORDER)
C0272499|T037|61642003|SNOMEDCT_US|MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HEMORRHAGE|MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HEMORRHAGE (DISORDER)
C0272499|T037|61642003|SNOMEDCT_US|MULTIPLE OPEN FRACTURES OF SKULL AND FACE WITH SUBARACHNOID, SUBDURAL AND EXTRADURAL HEMORRHAGE|MULTIPLE OPEN FRACTURES OF SKULL AND/OR FACE WITH SUBARACHNOID, SUBDURAL AND/OR EXTRADURAL HEMORRHAGE (DISORDER)
C0161399|T037|69820004|SNOMEDCT_US|INJURY OF OPTIC CHIASM|INJURY OF OPTIC CHIASM (DISORDER)
C0161399|T037|69820004|SNOMEDCT_US|INJURY OF OPTIC CHIASM |INJURY OF OPTIC CHIASM (DISORDER)
C0161399|T037|69820004|SNOMEDCT_US|INJURY TO THE OPTIC CHIASM|INJURY OF OPTIC CHIASM (DISORDER)
C0161399|T037|69820004|SNOMEDCT_US|INJURY TO OPTIC CHIASM|INJURY OF OPTIC CHIASM (DISORDER)
C0161399|T037|69820004|SNOMEDCT_US|INJURY OF OPTIC CHIASM |INJURY OF OPTIC CHIASM (DISORDER)
C0161399|T037|69820004|SNOMEDCT_US|OPTIC CHIASM INJURY|INJURY OF OPTIC CHIASM (DISORDER)
C0751814|T037||SNOMEDCT_US|INJ VASCULAR BRAIN
C0751814|T037||SNOMEDCT_US|VASCULAR INJ BRAIN
C0751814|T037||SNOMEDCT_US|BRAIN INJ VASCULAR
C0751814|T037||SNOMEDCT_US|BRAIN VASCULAR INJURY
C0751814|T037||SNOMEDCT_US|INJURY, BRAIN VASCULAR
C0751814|T037||SNOMEDCT_US|INJURY, VASCULAR BRAIN
C0751814|T037||SNOMEDCT_US|VASCULAR BRAIN INJURIES
C0751814|T037||SNOMEDCT_US|VASCULAR BRAIN INJURY
C0751814|T037||SNOMEDCT_US|BRAIN VASCULAR TRAUMA
C0751814|T037||SNOMEDCT_US|TRAUMA, BRAIN VASCULAR
C0751814|T037||SNOMEDCT_US|VASCULAR TRAUMAS, BRAIN
C0751814|T037||SNOMEDCT_US|CEREBROVASCULAR TRAUMA
C0751814|T037||SNOMEDCT_US|TRAUMA, CEREBROVASCULAR
C0751814|T037||SNOMEDCT_US|BRAIN INJURY, VASCULAR
C0751814|T037||SNOMEDCT_US|CEREBROVASCULAR TRAUMA [DISEASE/FINDING]
C0751814|T037||SNOMEDCT_US|INJURY, VASCULAR, BRAIN
C0751814|T037||SNOMEDCT_US|VASCULAR INJURY, BRAIN
C0751814|T037||SNOMEDCT_US|VASCULAR TRAUMA, BRAIN
C0751814|T037||SNOMEDCT_US|CEREBRAL VESSELS; INJURY
C0751814|T037||SNOMEDCT_US|INJURY; CEREBRAL VESSELS
C0273106|T037|28155008|SNOMEDCT_US|OPEN INTRACRANIAL WOUND AND EXTRADURAL HEMORRHAGE WITH CONCUSSION |EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|OPEN INTRACRANIAL WOUND AND EXTRADURAL HEMORRHAGE WITH CONCUSSION|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|HEAD INJURY WITH OPEN INTRACRANIAL WOUND AND EXTRADURAL HEMORRHAGE WITH CONCUSSION|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|EXTRADURAL HEM-CONCUSS|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|EXTRADURAL HAEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED |EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY, WITH OPEN INTRACRANIAL WOUND, WITH CONCUSSION, UNSPECIFIED|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|EXTRADURAL HAEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION |EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0273106|T037|28155008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND UNSPECIFIED CONCUSSION|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND CONCUSSION (DISORDER)
C0475077|T037|209933001|SNOMEDCT_US|HEAD INJURY WITH SUBARACHNOID HEMORRHAGE WITH MODERATE (1-24 HRS) LOSS OF CONSCIOUSNESS|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0475077|T037|209933001|SNOMEDCT_US|HEAD INJURY WITH SUBARACHNOID HEMORRHAGE WITH MODERATE (1-24 HRS) LOSS OF CONSCIOUSNESS |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0475077|T037|209933001|SNOMEDCT_US|HEAD INJURY WITH SUBARACHNOID HEMORRHAGE MODERATE (1-24 HR) LOSS OF CONSCIOUSNESS|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0475077|T037|209933001|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0475077|T037|209933001|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0475077|T037|209933001|SNOMEDCT_US|SUBARACHNOID HAEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0273070|T037|77768006|SNOMEDCT_US|HEAD INJURY WITH OPEN INTRACRANIAL WOUND AND INTRACRANIAL HEMORRHAGE|INTRACRANIAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0273070|T037|77768006|SNOMEDCT_US|OPEN INTRACRANIAL WOUND AND HEMORRHAGE |INTRACRANIAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0273070|T037|77768006|SNOMEDCT_US|OPEN INTRACRANIAL WOUND AND HEMORRHAGE|INTRACRANIAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0273070|T037|77768006|SNOMEDCT_US|INTRACRANIAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND|INTRACRANIAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0273070|T037|77768006|SNOMEDCT_US|INTRACRANIAL HAEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND|INTRACRANIAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0273070|T037|77768006|SNOMEDCT_US|INTRACRANIAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND |INTRACRANIAL HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0273087|T037|30400005|SNOMEDCT_US|MIDDLE MENINGEAL HEMORRHAGE FOLLOWING INJURY|MIDDLE MENINGEAL HEMORRHAGE FOLLOWING INJURY (DISORDER)
C0273087|T037|30400005|SNOMEDCT_US|MIDDLE MENINGEAL HEMORRHAGE FOLLOWING INJURY |MIDDLE MENINGEAL HEMORRHAGE FOLLOWING INJURY (DISORDER)
C0273087|T037|30400005|SNOMEDCT_US|MIDDLE MENINGEAL HAEMORRHAGE FOLLOWING INJURY|MIDDLE MENINGEAL HEMORRHAGE FOLLOWING INJURY (DISORDER)
C0273087|T037|30400005|SNOMEDCT_US|MIDDLE MENINGEAL HEMORRHAGE FOLLOWING INJURY [DUP] |MIDDLE MENINGEAL HEMORRHAGE FOLLOWING INJURY (DISORDER)
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEM FOLLOWING INJ, W/O MENT OF OPEN INTCRAN WOUND, WITH LOC OF UNSPEC DURATION|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEM FOLLOWING INJ, W/O MENT OF OPEN INTCRAN WOUND, WITH PROL LOC, W/O RTRN TO PECL|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEM-DEEP COMA|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEM-COMA NOS|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS] LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION |EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HAEMORRHAGE FOLLOWING INJURY WITHOUT MENTION OF OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS |EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND, WITH LOSS OF CONSCIOUSNESS|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|HEAD INJ - W/ EXTRADURAL HEMORRHAGE, W/O OPEN INTRACRANIAL WOUND W/ LOC|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HAEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS |EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0273104|T037|90178008|SNOMEDCT_US|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS OF UNSPECIFIED DURATION|EXTRADURAL HEMORRHAGE FOLLOWING INJURY WITHOUT OPEN INTRACRANIAL WOUND AND WITH LOSS OF CONSCIOUSNESS
C0475083|T037|209942008|SNOMEDCT_US|SUBARACHNOID HAEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0475083|T037|209942008|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0475083|T037|209942008|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH 1-24 HOURS LOSS OF CONSCIOUSNESS (DISORDER)
C0475082|T037|209941001|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS (DISORDER)
C0475082|T037|209941001|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS (DISORDER)
C0475082|T037|209941001|SNOMEDCT_US|SUBARACHNOID HAEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH LESS THAN 1 HOUR LOSS OF CONSCIOUSNESS (DISORDER)
C0475085|T037|209944009|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0475085|T037|209944009|SNOMEDCT_US|SUBARACHNOID HAEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0475085|T037|209944009|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS WITHOUT RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160228|T037|5251007|SNOMEDCT_US|HEAD INJURY WITH OPEN INTRACRANIAL WOUND AND SUBARACHNOID HEMORRHAGE |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160228|T037|5251007|SNOMEDCT_US|HEAD INJURY WITH OPEN INTRACRANIAL WOUND AND SUBARACHNOID HEMORRHAGE|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160228|T037|5251007|SNOMEDCT_US|OPEN INTRACRANIAL WOUND AND SUBARACHNOID HEMORRHAGE|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160228|T037|5251007|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160228|T037|5251007|SNOMEDCT_US|SUBARACHNOID HAEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160228|T037|5251007|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|OPEN INTRACRANIAL WOUND AND SUBARACHNOID HEMORRHAGE LOSS OF CONSCIOUSNESS GREATER THAN 24 HOURS THEN RETURN TO PREVIOUS LEVEL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|OPEN INTRACRANIAL WOUND AND SUBARACHNOID HEMORRHAGE WITH PROLONGED (> 24 HRS) LOSS OF CONSCIOUSNESS WITH RETURN TO PRIOR LEVEL OF CONSCIOUSNESS |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|OPEN INTRACRANIAL WOUND AND SUBARACHNOID HEMORRHAGE WITH PROLONGED (> 24 HRS) LOSS OF CONSCIOUSNESS WITH RETURN TO PRIOR LEVEL OF CONSCIOUSNESS|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|HEAD INJURY WITH OPEN INTRACRANIAL WOUND AND SUBARACHNOID HEMORRHAGE WITH LOC OVER 24 HR, THEN RETURN TO PRIOR LEVEL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|SUBARAC HEM FOLLOWING INJ, WITH OPEN INTCRAN WOUND, WITH PROLONGED LOC AND RETURN TO PECL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|OP SUBARACH HEM-PROL COM|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH PROLONGED [MORE THAN 24 HOURS) LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|SUBARACHNOID HAEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND, WITH MORE THAN 24 HOURS LOSS OF CONSCIOUSNESS AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|SUBARACHNOID HAEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0160233|T037|73439007|SNOMEDCT_US|SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL |SUBARACHNOID HEMORRHAGE FOLLOWING INJURY WITH OPEN INTRACRANIAL WOUND AND PROLONGED LOSS OF CONSCIOUSNESS (MORE THAN 24 HOURS) AND RETURN TO PRE-EXISTING CONSCIOUS LEVEL (DISORDER)
C0541931|T037||SNOMEDCT_US|ENCEPHALITIS TOXIC CHRONIC
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PALSY|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PALSY NOS|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PALSY, UNSPECIFIED|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CP (CEREBRAL PALSY)|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PALSY [DISEASE/FINDING]|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PALSY |CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|PALSY;CEREBRAL|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CP|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PALSY (CP)|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PALSY |CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CONGENITAL CEREBRAL PALSY|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|INFANTILE CEREBRAL PALSY|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PARALYSIS|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|PALSY CEREBRAL|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CP - CEREBRAL PALSY|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL; PARALYSIS|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|PARALYSIS; CEREBRAL|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PALSY, NOS|CEREBRAL PALSY (DISORDER)
C0007789|T037|128188000|SNOMEDCT_US|CEREBRAL PALSY [AMBIGUOUS]|CEREBRAL PALSY (DISORDER)
C0553767|T037|275466008|SNOMEDCT_US|CONGEN CEREBRAL PALSY|CONGENITAL CEREBRAL PALSY (DISORDER)
C0553767|T037|275466008|SNOMEDCT_US|CONGENITAL CEREBRAL PALSY NOS |CONGENITAL CEREBRAL PALSY (DISORDER)
C0553767|T037|275466008|SNOMEDCT_US|CONGENITAL CEREBRAL PALSY|CONGENITAL CEREBRAL PALSY (DISORDER)
C0553767|T037|275466008|SNOMEDCT_US|CONGENITAL CEREBRAL PALSY NOS|CONGENITAL CEREBRAL PALSY (DISORDER)
C0553767|T037|275466008|SNOMEDCT_US|CEREBRAL PALSY CONGENITAL|CONGENITAL CEREBRAL PALSY (DISORDER)
C0553767|T037|275466008|SNOMEDCT_US|CONGENITAL CEREBRAL PALSY |CONGENITAL CEREBRAL PALSY (DISORDER)
C0553767|T037|275466008|SNOMEDCT_US|CONGENITAL CEREBRAL PALSY |CONGENITAL CEREBRAL PALSY (DISORDER)
C0553767|T037|275466008|SNOMEDCT_US|CEREBRAL PALSY, CONGENITAL|CONGENITAL CEREBRAL PALSY (DISORDER)
C0270719|T037|15139001|SNOMEDCT_US|CHATTER-BOX SYNDROME|CHRONIC BRAIN-HYDROCEPHALUS SYNDROME (DISORDER)
C0270719|T037|15139001|SNOMEDCT_US|CHRONIC BRAIN-HYDROCEPHALUS SYNDROME|CHRONIC BRAIN-HYDROCEPHALUS SYNDROME (DISORDER)
C0270719|T037|15139001|SNOMEDCT_US|COCKTAIL PARTY SYNDROME|CHRONIC BRAIN-HYDROCEPHALUS SYNDROME (DISORDER)
C0270719|T037|15139001|SNOMEDCT_US|CHRONIC BRAIN-HYDROCEPHALUS SYNDROME |CHRONIC BRAIN-HYDROCEPHALUS SYNDROME (DISORDER)
C0270674|T037|27195007|SNOMEDCT_US|CHRONIC NON-PSYCHOTIC BRAIN SYNDROME|CHRONIC NON-PSYCHOTIC BRAIN SYNDROME (DISORDER)
C0270674|T037|27195007|SNOMEDCT_US|CHRONIC NON-PSYCHOTIC BRAIN SYNDROME |CHRONIC NON-PSYCHOTIC BRAIN SYNDROME (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOL-INDUCED PERSISTENT DEMENTIA |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOL-INDUCED PERSISTENT DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH DEMENTIA |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOL DEPENDENCE WITH DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOL INDUCED PERSISTING DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOL PERSIST DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|DEMENTIA;ALCOHOLIC|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOLIC DEMENTIA NOS|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|[X]ALCOHOLIC DEMENTIA NOS|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|[X]CHRONIC ALCOHOLIC BRAIN SYNDROME|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOLIC DEMENTIA NOS |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|CHRONIC ORGANIC MENTAL DISORDER ALCOHOLIC BRAIN SYNDROME|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|CHRONIC ALCOHOLIC BRAIN SYNDROME|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|CHRONIC ALCOHOLIC BRAIN SYNDROME |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|DEMENTIA ASSOCIATED WITH ALCOHOLISM|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOL-INDUCED PERSISTING DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOLIC DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|CHRONIC ALCOHOLIC BRAIN SYNDROME |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|DEMENTIA ASSOCIATED WITH ALCOHOLISM |DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|BRAIN; SYNDROME, ALCOHOLIC (CHRONIC)|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|DEMENTIA; ALCOHOLIC|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|DEMENTIA; ALCOHOL|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOL; DEMENTIA|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|SYNDROME; BRAIN, ALCOHOLIC (CHRONIC)|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0236656|T037|281004|SNOMEDCT_US|ALCOHOLISM ASSOCIATED WITH DEMENTIA NOS|DEMENTIA ASSOCIATED WITH ALCOHOLISM (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|THIS IS POTENTIALLY REVERSIBLE AND SO MIGHT DELIVER FALSE POSITIVES, HOWEVER WITH A LIVER SPECIFIC INTAKE FORM I THINK THESE FALSE POSITIVES ARE ACCEPTABLE/VALUABLE|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHIES, PORTOSYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHIES|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|PORTOSYSTEMIC ENCEPHALOPATHIES|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPH HEPATOCEREBRAL|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPH PORTAL SYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC ENCEPH|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|PORTOSYSTEMIC ENCEPH|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPH PORTOSYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|PORTAL SYSTEMIC ENCEPH|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPH|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPH HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY |HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPHALOPATHY -RETIRED-|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHIES, HEPATOCEREBRAL|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPHALOPATHIES|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHIES, PORTAL-SYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|PORTAL SYSTEMIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|PORTAL-SYSTEMIC ENCEPHALOPATHIES|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY NOS|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|PORTOSYSTEMIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHY, HEPATOCEREBRAL|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY [DISEASE/FINDING]|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|PORTAL-SYSTEMIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHY, HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHY, PORTAL-SYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHY, PORTOSYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC COMA/ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHY, PORTAL SYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|GAUSTAD'S SYNDROME|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|PORTAL SYSTEMIC ENCEPHALOPATHY |HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|TRANSIENT HEPATARGY SYNDROME|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHY - HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATOCEREBRAL ENCEPHALOPATHY |HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHY HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HE - HEPATIC ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY |HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHY; HEPATIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|ENCEPHALOPATHY; PORTOSYSTEMIC|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|HEPATIC; ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C0019151|T037|123049003|SNOMEDCT_US|PORTOSYSTEMIC; ENCEPHALOPATHY|HEPATOCEREBRAL ENCEPHALOPATHY (DISORDER)
C2729507|T037||SNOMEDCT_US|HEPATIC ENCEPHALOPATHY WITH COMA 
C2729507|T037||SNOMEDCT_US|HEPATIC ENCEPHALOPATHY WITH COMA
C0019147|T037|72836002|SNOMEDCT_US|COMAS, HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|HEPATIC COMAS|HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|COMA, HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|HEPATIC COMA|HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|COMA HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|HEPATIC COMA NOS|HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|COMA;HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|HEPATIC COMA |HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|HEPATOCEREBRAL INTOXICATION|HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|COMA; HEPATIC|HEPATIC COMA (DISORDER)
C0019147|T037|72836002|SNOMEDCT_US|HEPATIC; COMA|HEPATIC COMA (DISORDER)
C3266165|T037|449901005|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE|HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE (DISORDER)
C3266165|T037|449901005|SNOMEDCT_US|HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE |HEPATIC ENCEPHALOPATHY IN FULMINANT HEPATIC FAILURE (DISORDER)
C0751198|T037||SNOMEDCT_US|HEPATIC STUPORS
C0751198|T037||SNOMEDCT_US|STUPOR, HEPATIC
C0751198|T037||SNOMEDCT_US|STUPORS, HEPATIC
C0751198|T037||SNOMEDCT_US|HEPATIC STUPOR
C1836797|T037||SNOMEDCT_US|COMBINED OXIDATIVE PHOSPHORYLATION DEFICIENCY 1
C1836797|T037||SNOMEDCT_US|HEPATOENCEPHALOPATHY, EARLY FATAL PROGRESSIVE
C4024937|T037||SNOMEDCT_US|CHRONIC HEPATIC ENCEPHALOPATHY
