# C0003467|T048|139476005|SNOMEDCT_US|ANXIETY|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DISORDERS|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0860603|T048||SNOMEDCT_US|ANXIETY SYMPTOMS
C1963064|T048||SNOMEDCT_US|ANXIETY ADVERSE EVENT
C4050613|T048||SNOMEDCT_US|ANXIETY SCALE (BASC-2)
C0085380|T048|191731009|SNOMEDCT_US|ANXIETIES, DENTAL|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENTAL ANXIETIES|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENTAL ANXIETY|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENTAL FEARS|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENTAL PHOBIAS|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|FEARS, DENTAL|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|ODONTOPHOBIAS|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|PHOBIAS, DENTAL|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENT ANXIETY|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|ANXIETY DENT|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENT PHOBIA|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|PHOBIA DENT|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|FEAR DENT|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENT FEAR|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENTAL PHOBIA |DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENTAL PHOBIA|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENTAL FEAR|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|ODONTOPHOBIA|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|FEAR, DENTAL|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|ANXIETY, DENTAL|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|PHOBIA, DENTAL|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|FEAR OF DENTIST|DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|DENTAL PHOBIA |DENTAL PHOBIA (DISORDER)
C0085380|T048|191731009|SNOMEDCT_US|FEAR OF DENTIST |DENTAL PHOBIA (DISORDER)
C0003476|T048|304896009|SNOMEDCT_US|ANXIETY, CASTRATION|CASTRATION ANXIETY COMPLEX (FINDING)
C0003476|T048|304896009|SNOMEDCT_US|CASTRATION ANXIETY|CASTRATION ANXIETY COMPLEX (FINDING)
C0003476|T048|304896009|SNOMEDCT_US|CASTRATION COMPLICES|CASTRATION ANXIETY COMPLEX (FINDING)
C0003476|T048|304896009|SNOMEDCT_US|COMPLICES, CASTRATION|CASTRATION ANXIETY COMPLEX (FINDING)
C0003476|T048|304896009|SNOMEDCT_US|COMPLEX, CASTRATION|CASTRATION ANXIETY COMPLEX (FINDING)
C0003476|T048|304896009|SNOMEDCT_US|CASTRATION COMPLEX|CASTRATION ANXIETY COMPLEX (FINDING)
C0003476|T048|304896009|SNOMEDCT_US|CASTRATION ANXIETY COMPLEX|CASTRATION ANXIETY COMPLEX (FINDING)
C0003476|T048|304896009|SNOMEDCT_US|CASTRATION ANXIETY COMPLEX |CASTRATION ANXIETY COMPLEX (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|ANXIETIES|ANXIOUSNESS (& SYMPTOM) (FINDING)
# C0003467|T048|139476005|SNOMEDCT_US|ANXIETY|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|ANXIETY REACTION|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|RNDX ANXIETY |ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|RNDX ANXIETY|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|FEELING;ANXIOUS|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|ANXIOUSNESS|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|ANXIOUSNESS (& SYMPTOM) |ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|ANXIOUSNESS (& SYMPTOM)|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|ANXIOUSNESS - SYMPTOM|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|ANXIOUS BEHAVIOR|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|-- ANXIETY|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|REACTION ANXIETY|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|ANXIETY |ANXIOUSNESS (& SYMPTOM) (FINDING)
C0003467|T048|139476005|SNOMEDCT_US|ANXIOUS; SENSATION|ANXIOUSNESS (& SYMPTOM) (FINDING)
C0563150|T048|285247003|SNOMEDCT_US|CATASTROPHIZATION|CATASTROPHIZATION (FINDING)
C0563150|T048|285247003|SNOMEDCT_US|CATASTROPHIZING|CATASTROPHIZATION (FINDING)
C0563150|T048|285247003|SNOMEDCT_US|CATASTROPHISATION|CATASTROPHIZATION (FINDING)
C0563150|T048|285247003|SNOMEDCT_US|CATASTROPHIZATION |CATASTROPHIZATION (FINDING)
C0458631|T048|279622009|SNOMEDCT_US|PERFORMANCE FEAR|PERFORMANCE ANXIETY (FINDING)
C0458631|T048|279622009|SNOMEDCT_US|ANXIETY, PERFORMANCE|PERFORMANCE ANXIETY (FINDING)
C0458631|T048|279622009|SNOMEDCT_US|PERFORMANCE ANXIETY|PERFORMANCE ANXIETY (FINDING)
C0458631|T048|279622009|SNOMEDCT_US|ANXIETIES, PERFORMANCE|PERFORMANCE ANXIETY (FINDING)
C0458631|T048|279622009|SNOMEDCT_US|PERFORMANCE ANXIETIES|PERFORMANCE ANXIETY (FINDING)
C0458631|T048|279622009|SNOMEDCT_US|PERFORMANCE ANXIETY |PERFORMANCE ANXIETY (FINDING)
C2077827|T048||SNOMEDCT_US|ANXIETY WHICH COMES AND GOES
C2077827|T048||SNOMEDCT_US|ANXIETY EPISODIC
C2077827|T048||SNOMEDCT_US|INTERMITTENT ANXIETY 
C2077827|T048||SNOMEDCT_US|ANXIETY WHICH COMES AND GOES (EPISODIC)
C2077827|T048||SNOMEDCT_US|INTERMITTENT ANXIETY
C0549259|T048||SNOMEDCT_US|ANXIETY AGGRAVATED
C0262376|T048||SNOMEDCT_US|GENERALIZED; ANXIETY
C0262376|T048||SNOMEDCT_US|ANXIETY; GENERALIZED
C0262377|T048||SNOMEDCT_US|SITUATIONAL ANXIETY
C0235111|T048||SNOMEDCT_US|ANXIETY COMPLEX
C0457041|T048|277838008|SNOMEDCT_US|ANXIETY ABOUT APPEARING RIDICULOUS|ANXIETY ABOUT APPEARING RIDICULOUS (FINDING)
C0457041|T048|277838008|SNOMEDCT_US|ANXIETY ABOUT APPEARING RIDICULOUS |ANXIETY ABOUT APPEARING RIDICULOUS (FINDING)
C0231397|T048|35429005|SNOMEDCT_US|ANTICIPATORY ANXIETY|ANTICIPATORY ANXIETY (FINDING)
C0231397|T048|35429005|SNOMEDCT_US|ANTICIPATORY ANXIETY |ANTICIPATORY ANXIETY (FINDING)
C0231397|T048|35429005|SNOMEDCT_US|ANTICIPATORY ANXIETY, NOS|ANTICIPATORY ANXIETY (FINDING)
C0231398|T048|11458009|SNOMEDCT_US|ANTICIPATORY ANXIETY, MILD|ANTICIPATORY ANXIETY, MILD (FINDING)
C0231398|T048|11458009|SNOMEDCT_US|ANTICIPATORY ANXIETY, MILD |ANTICIPATORY ANXIETY, MILD (FINDING)
C0231400|T048|5874002|SNOMEDCT_US|ANTICIPATORY ANXIETY, SEVERE|ANTICIPATORY ANXIETY, SEVERE (FINDING)
C0231400|T048|5874002|SNOMEDCT_US|ANTICIPATORY ANXIETY, SEVERE |ANTICIPATORY ANXIETY, SEVERE (FINDING)
C0154455|T048||SNOMEDCT_US|OTHER ANXIETY STATES
C0154455|T048||SNOMEDCT_US|ANXIETY STATE NEC
C0030319|T048|268627007|SNOMEDCT_US|DISORDERS, PANIC|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC DISORDER|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC DISORDERS|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|DISORDER, PANIC|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC DISORDER [EPISODIC PAROXYSMAL ANXIETY]|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC DIS|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC ANXIETY SYNDROME|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC DISORDER [DISEASE/FINDING]|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|DISORDER;PANIC|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|[X]PANIC DISORDER [EPISODIC PAROXYSMAL ANXIETY] |PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|[X]PANIC DISORDER [EPISODIC PAROXYSMAL ANXIETY]|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC DISORDER |PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC DISORDER |PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|-- PANIC DISORDER|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC DISORDER NOS|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|EPISODIC PAROXYSMAL ANXIETY DISORDER|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC DISORDER |PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|DISORDER; PANIC|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|PANIC; DISORDER|PANIC DISORDER (FINDING)
C0030319|T048|268627007|SNOMEDCT_US|[X]PANIC DISORDER [EPISODIC PAROXYSMAL ANXIETY] |PANIC DISORDER (FINDING)
C2128827|T048||SNOMEDCT_US|ANXIOUS ON A DAILY BASIS
C2128827|T048||SNOMEDCT_US|ANXIETY DAILY
C2128827|T048||SNOMEDCT_US|ANXIOUS EVERY DAY
C2128827|T048||SNOMEDCT_US|DAILY ANXIETY 
C2128827|T048||SNOMEDCT_US|DAILY ANXIETY
C2219855|T048||SNOMEDCT_US|ANXIETY WITH FEAR OF DYING 
C2219855|T048||SNOMEDCT_US|ANXIETY WITH FEAR OF DYING
C2219855|T048||SNOMEDCT_US|ANXIETY WITH A FEAR OF DYING
C2219861|T048||SNOMEDCT_US|ANXIETY WITH FEELINGS OF UNREALITY
C2219861|T048||SNOMEDCT_US|ANXIETY WITH FEELINGS OF UNREALITY 
C0522179|T048|191732002|SNOMEDCT_US|FEAR OF DEATH|FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|THANATOPHOBIA|FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|FEAR (OF);DEATH|FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|FEAR (OF);DYING|FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|DEATH ANXIETY|FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|FEAR ABOUT DEATH|FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|FEAR OF DYING|FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|FEAR OF DYING |FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|FEAR OF DEATH |FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|DEATH ANXIETY |FEAR OF DEATH (DISORDER)
C0522179|T048|191732002|SNOMEDCT_US|FEAR OF DEATH |FEAR OF DEATH (DISORDER)
C2219860|T048||SNOMEDCT_US|ANXIETY WITH DIZZINESS OR UNSTEADY FEELINGS 
C2219860|T048||SNOMEDCT_US|ANXIETY WITH DIZZINESS OR UNSTEADY FEELINGS
C1854339|T048||SNOMEDCT_US|ANXIETY (WITH PHEOCHROMOCYTOMA)
C0700613|T048|191704006|SNOMEDCT_US|ANXIETY STATES|ANXIETY STATE UNSPECIFIED (FINDING)
C0700613|T048|191704006|SNOMEDCT_US|ANXIETY STATE|ANXIETY STATE UNSPECIFIED (FINDING)
C0700613|T048|191704006|SNOMEDCT_US|ANXIETY STATE NOS|ANXIETY STATE UNSPECIFIED (FINDING)
C0700613|T048|191704006|SNOMEDCT_US|ANXIETY STATE UNSPECIFIED |ANXIETY STATE UNSPECIFIED (FINDING)
C0700613|T048|191704006|SNOMEDCT_US|ANXIETY STATE NOS |ANXIETY STATE UNSPECIFIED (FINDING)
C0700613|T048|191704006|SNOMEDCT_US|ANXIETY STATE UNSPECIFIED|ANXIETY STATE UNSPECIFIED (FINDING)
C0700613|T048|191704006|SNOMEDCT_US|ANXIETY STATE, UNSPECIFIED|ANXIETY STATE UNSPECIFIED (FINDING)
C0700613|T048|191704006|SNOMEDCT_US|ANXIETY STATE |ANXIETY STATE UNSPECIFIED (FINDING)
C0700613|T048|191704006|SNOMEDCT_US|STATE; ANXIETY|ANXIETY STATE UNSPECIFIED (FINDING)
C0700613|T048|191704006|SNOMEDCT_US|ANXIETY; STATE|ANXIETY STATE UNSPECIFIED (FINDING)
C0474385|T048|247825008|SNOMEDCT_US|ANXIETY ABOUT BEHAVIOR OR PERFORMANCE|ANXIETY ABOUT BEHAVIOR OR PERFORMANCE (FINDING)
C0474385|T048|247825008|SNOMEDCT_US|ANXIETY ABOUT BEHAVIOUR OR PERFORMANCE|ANXIETY ABOUT BEHAVIOR OR PERFORMANCE (FINDING)
C0474385|T048|247825008|SNOMEDCT_US|ANXIETY ABOUT SOCIAL FUNCTIONING|ANXIETY ABOUT BEHAVIOR OR PERFORMANCE (FINDING)
C0474385|T048|247825008|SNOMEDCT_US|ANXIETY ABOUT BEHAVIOR OR PERFORMANCE |ANXIETY ABOUT BEHAVIOR OR PERFORMANCE (FINDING)
C0424145|T048|247808006|SNOMEDCT_US|ANXIETY ABOUT BODY FUNCTION OR HEALTH|ANXIETY ABOUT BODY FUNCTION OR HEALTH (FINDING)
C0424145|T048|247808006|SNOMEDCT_US|ANXIETY ABOUT HEALTH|ANXIETY ABOUT BODY FUNCTION OR HEALTH (FINDING)
C0424145|T048|247808006|SNOMEDCT_US|ANXIETY ABOUT BODY FUNCTION OR HEALTH |ANXIETY ABOUT BODY FUNCTION OR HEALTH (FINDING)
C0558210|T048|225637002|SNOMEDCT_US|ANXIETY ABOUT LOSS OF CONTROL|ANXIETY ABOUT LOSS OF CONTROL (FINDING)
C0558210|T048|225637002|SNOMEDCT_US|ANXIETY ABOUT LOSS OF CONTROL |ANXIETY ABOUT LOSS OF CONTROL (FINDING)
C0558209|T048|225636006|SNOMEDCT_US|ANXIETY ABOUT FORCED DEPENDENCE|ANXIETY ABOUT FORCED DEPENDENCE (FINDING)
C0558209|T048|225636006|SNOMEDCT_US|ANXIETY ABOUT FORCED DEPENDENCE |ANXIETY ABOUT FORCED DEPENDENCE (FINDING)
C0558208|T048|225635005|SNOMEDCT_US|ANXIETY ABOUT TREATMENT|ANXIETY ABOUT TREATMENT (FINDING)
C0558208|T048|225635005|SNOMEDCT_US|ANXIETY ABOUT TREATMENT |ANXIETY ABOUT TREATMENT (FINDING)
C0870858|T048||SNOMEDCT_US|MATHEMATICS ANXIETY
C0424166|T048|247832004|SNOMEDCT_US|SOCIAL FEAR|SOCIAL FEAR (FINDING)
C0424166|T048|247832004|SNOMEDCT_US|SOCIAL FEAR |SOCIAL FEAR (FINDING)
C0424166|T048|247832004|SNOMEDCT_US|SOCIAL ANXIETY|SOCIAL FEAR (FINDING)
C0424169|T048|247835002|SNOMEDCT_US|FEAR OF PUBLIC SPEAKING|FEAR OF PUBLIC SPEAKING (FINDING)
C0424169|T048|247835002|SNOMEDCT_US|FEAR OF PUBLIC SPEAKING |FEAR OF PUBLIC SPEAKING (FINDING)
C0424169|T048|247835002|SNOMEDCT_US|SPEECH ANXIETY|FEAR OF PUBLIC SPEAKING (FINDING)
C0424169|T048|247835002|SNOMEDCT_US|COMMUNICATION APPREHENSION|FEAR OF PUBLIC SPEAKING (FINDING)
C0871504|T048||SNOMEDCT_US|TEST ANXIETY
C0935548|T048||SNOMEDCT_US|COMPUTER ANXIETY
C0577602|T048|300894000|SNOMEDCT_US|ANXIOUS PARENT|PARENTAL ANXIETY (FINDING)
C0577602|T048|300894000|SNOMEDCT_US|ANXIETY;PARENTAL|PARENTAL ANXIETY (FINDING)
C0577602|T048|300894000|SNOMEDCT_US|PARENTAL ANXIETY|PARENTAL ANXIETY (FINDING)
C0577602|T048|300894000|SNOMEDCT_US|ANXIOUS PARENTS|PARENTAL ANXIETY (FINDING)
C0577602|T048|300894000|SNOMEDCT_US|PARENTAL ANXIETY |PARENTAL ANXIETY (FINDING)
C0700031|T048|300895004|SNOMEDCT_US|ANXIETY ATTACKS|ANXIETY ATTACK (FINDING)
C0700031|T048|300895004|SNOMEDCT_US|ANXIETY ATTACK|ANXIETY ATTACK (FINDING)
C0700031|T048|300895004|SNOMEDCT_US|ANXIETY ATTACK |ANXIETY ATTACK (FINDING)
C0700031|T048|300895004|SNOMEDCT_US|ATTACK(S);ANXIETY|ANXIETY ATTACK (FINDING)
C0231402|T048|61387006|SNOMEDCT_US|MODERATE ANXIETY|MODERATE ANXIETY (FINDING)
C0231402|T048|61387006|SNOMEDCT_US|MODERATE ANXIETY |MODERATE ANXIETY (FINDING)
C0231401|T048|70997004|SNOMEDCT_US|MILD ANXIETY|MILD ANXIETY (FINDING)
C0231401|T048|70997004|SNOMEDCT_US|MILD ANXIETY |MILD ANXIETY (FINDING)
C0030318|T048|79823003|SNOMEDCT_US|PANIC|PANIC (FINDING)
C0030318|T048|79823003|SNOMEDCT_US|PANICS|PANIC (FINDING)
C0030318|T048|79823003|SNOMEDCT_US|PANIC REACTION|PANIC (FINDING)
C0030318|T048|79823003|SNOMEDCT_US|PANIC STATE|PANIC (FINDING)
C0030318|T048|79823003|SNOMEDCT_US|REACTION PANIC|PANIC (FINDING)
C0030318|T048|79823003|SNOMEDCT_US|PANIC |PANIC (FINDING)
C0030318|T048|79823003|SNOMEDCT_US|PANIC; STATE|PANIC (FINDING)
C0030318|T048|79823003|SNOMEDCT_US|STATE; PANIC|PANIC (FINDING)
C0030318|T048|79823003|SNOMEDCT_US|PANIC [AMBIGUOUS]|PANIC (FINDING)
C0233483|T048|81350009|SNOMEDCT_US|FREE-FLOATING ANXIETY|FREE-FLOATING ANXIETY (FINDING)
C0233483|T048|81350009|SNOMEDCT_US|FREE-FLOATING ANXIETY |FREE-FLOATING ANXIETY (FINDING)
C0860603|T048||SNOMEDCT_US|ANXIETY 
C0860603|T048||SNOMEDCT_US|ANXIETY
C0860603|T048||SNOMEDCT_US|ANXIETY SYMPTOMS
C0860603|T048||SNOMEDCT_US|ANXIETY SYMPTOMS NOS
C0860603|T048||SNOMEDCT_US|ANXIETY; COMPLAINT
C0028768|T048|192411009|SNOMEDCT_US|DISORDERS, OBSESSIVE-COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE DISORDER|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE DISORDERS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|DISORDER, OBSESSIVE-COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE COMPULSIVE DISORDER|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OCD|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE COMPULSIVE DIS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE COMPULSIVE DISORDER |[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OCD (OBSESSIVE COMPULSIVE DISORDER)|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|NEUROSES, OBSESSIVE-COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|NEUROSIS, OBSESSIVE COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE NEUROSIS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|ANANKASTIC PERSONALITIES|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|PERSONALITIES, ANANKASTIC|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|PERSONALITY, ANANKASTIC|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE NEUROSES|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE DIS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE DISORDER [DISEASE/FINDING]|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|NEUROSIS, OBSESSIVE-COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|ANANKASTIC PERSONALITY|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|DISORDER;OBSESSIVE-COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|ANANCASTIC NEUROSIS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED |[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE DISORDER |[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OCD - OBSESSIVE-COMPULSIVE DISORDER|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|ANANKASTIC NEUROSIS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE COMPULSIVE DISORDER |[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE COMPULSIVE NEUROSIS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE DISORDER NOS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE DISORDER NOS |[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|-- OBSESSIVE COMPULSIVE DISORDER|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|REACTION OBSESSIVE-COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE REACTION|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|DISORDER; OBSESSIVE-COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|NEUROSIS; ANANKASTIC|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|NEUROSIS; OBSESSIVE-COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE NEUROSIS OR REACTION|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE; DISORDER|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE; NEUROSIS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE-COMPULSIVE; REACTION|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|REACTION; OBSESSIVE-COMPULSIVE|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|ANANKASTIC; NEUROSIS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0028768|T048|192411009|SNOMEDCT_US|OBSESSIVE COMPULSIVE DISORDER, NOS|[X]OBSESSIVE-COMPULSIVE DISORDER, UNSPECIFIED (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIA|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|DISORDER, PHOBIC|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|DISORDERS, PHOBIC|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC DISORDER|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC DISORDERS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC ANXIETY DISORDER, UNSPECIFIED|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC ANXIETY DISORDERS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC STATE|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC DIS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC ANXIETY DISORDER|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIA |PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIA NOS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC STATE NOS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|NEUROSES, PHOBIC|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC DISORDERS [DISEASE/FINDING]|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIAS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC NEUROSES|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIAS NOS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|[X]PHOBIC ANXIETY DISORDER, UNSPECIFIED |PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIA |PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|[X]PHOBIC ANXIETY DISORDERS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC DISORDER NOS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC DISORDER NOS |PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC ANXIETY|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|[X]PHOBIC ANXIETY DISORDER, UNSPECIFIED|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIA UNSPECIFIED|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC ANXIETY DISORDER |PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|[X]PHOBIC ANXIETY DISORDERS |PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC NEUROSIS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|ABNORMAL FEAR|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIA UNSPECIFIED |PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIA, UNSPECIFIED|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC DISORDER |PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|NEUROSIS; PHOBIC|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIA; STATE|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC; ANXIETY DISORDER|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC; NEUROSIS|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIC; STATE|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|STATE; PHOBIA|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|STATE; PHOBIC|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|ANXIETY DISORDER; PHOBIC|PHOBIC ANXIETY DISORDER (DISORDER)
C0349231|T048|154884005|SNOMEDCT_US|PHOBIA, NOS|PHOBIC ANXIETY DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST-TRAUMATIC STRESS DISORDER|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|NEUROSES, POST TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST TRAUMATIC STRESS DISORDERS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST-TRAUMATIC NEUROSES|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POSTTRAUMATIC NEUROSES|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POSTTRAUMATIC STRESS DISORDER|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|PTSD|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS DISORDER, POST-TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS DISORDER, POSTTRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS DISORDERS, POST TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS DISORDERS, POST-TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST-TRAUMATIC STRESS DISORDER (PTSD)|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POSTTRAUMATIC STRESS DISORDERS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST TRAUMATIC STRESS DIS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POSTTRAUMATIC STRESS DIS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS DIS POSTTRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS DIS POST TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|COMBAT FATIGUE|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|TRAUMATIC NEUROSIS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST-TRAUMATIC STRESS DISORDER |POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST-TRAUMATIC STRESS DISORDER, UNSPECIFIED|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS DISORDER, POST TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST-TRAUMATIC STRESS DISORDERS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|NEUROSES, POSTTRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS DISORDERS, POST-TRAUMATIC [DISEASE/FINDING]|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS DISORDERS, POSTTRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|NEUROSES, POST-TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|DISORDER;POST TRAUMATIC STRESS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST-TRAUMATIC STRESS DISORDER |POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|-- POST TRAUMATIC STRESS DISORDER|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|PTSD - POST-TRAUMATIC STRESS DISORDER|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST-TRAUMATIC STRESS SYNDROME|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POSTTRAUMATIC STRESS DISORDER |POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|DISORDER, POST-TRAUMATIC STRESS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|DISORDER; POST-TRAUMATIC STRESS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|DISORDER; STRESS, POST-TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|NEUROSIS; TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST-TRAUMATIC STRESS; DISORDER|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|STRESS; DISORDER, POST-TRAUMATIC|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|TRAUMATIC; NEUROSIS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POSTTRAUMATIC STRESS DISORDER, NOS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POSTTRAUMATIC STRESS DISORDER NOS|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0038436|T048|192415000|SNOMEDCT_US|POST TRAUMATIC STRESS DISORDER|POST-TRAUMATIC STRESS DISORDER (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|ASTHENIAS, NEUROCIRCULATORY|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CARDIAC NEUROSES|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|NEUROCIRCULATORY ASTHENIA|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|NEUROCIRCULATORY ASTHENIAS|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|NEUROSES, CARDIAC|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|ASTHENIA, NEUROCIRCULATORY|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|NEUROSIS, CARDIAC|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|SYNDROME, EFFORT|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CARDIAC NEUROSIS |CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CARDIAC NEUROSIS|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|PSYCHOGEN CARDIOVASC DIS|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|NEUROCIRCULATORY ASTHENIA [DISEASE/FINDING]|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|EFFORT SYNDROME|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|NEUROSIS;CARDIAC|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|[X]NEUROCIRCULATORY ASTHENIA|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|[X]CARDIAC NEUROSIS|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|[X]DA COSTA'S SYNDROME|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CARDIOVASCULAR DISORDER, PSYCHOGENIC|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CARDIAC NEUROSIS |CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|DA COSTA'S SYNDROME|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CARDIOVASCULAR NEUROSIS|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CEREBROCARDIAC NEUROSIS|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|NEUROCIRCULATORY ASTHENIA |CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CEREBROCARDIAC NEUROSIS |CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CEREBROCARDIAC SYNDROME|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|IRRITABLE HEART SYNDROME|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CARDIONEUROSIS|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|KRISHABER'S DISEASE|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|SYNDROME EFFORT|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|NEUROSIS CARDIOVASCULAR|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|CARDIOVASCULAR MALFUNCTION ARISING FROM MENTAL FACTORS|CEREBROCARDIAC NEUROSIS (DISORDER)
C0027821|T048|72994002|SNOMEDCT_US|NEUROCIRCULATORY ASTHENIA |CEREBROCARDIAC NEUROSIS (DISORDER)
C0856254|T048|191775008|SNOMEDCT_US|NEUROTIC PERSONALITY|NEUROTIC PERSONALITY
C0860602|T048||SNOMEDCT_US|ANXIOUS PERSONALITY
C0236121|T048||SNOMEDCT_US|NEUROSIS GI
C0236121|T048||SNOMEDCT_US|GASTROINTESTINAL NEUROSIS
C0270549|T048|21897009|SNOMEDCT_US|GENERALIZED ANXIETY DISORDER|GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GENERALISED ANXIETY DISORDER|GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GENERALIZED ANXIETY DISORDER |GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GAD|GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GENERALIZED ANXIETY DIS|GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GENERALISED ANXIETY DISORDER |GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GAD - GENERALISED ANXIETY DISORDER|GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GAD - GENERALIZED ANXIETY DISORDER|GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GENERALIZED ANXIETY DISORDER |GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GENERALIZED; ANXIETY DISORDER|GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|ANXIETY DISORDER; GENERALIZED|GENERALIZED ANXIETY DISORDER (DISORDER)
C0270549|T048|21897009|SNOMEDCT_US|GENERALISED ANXIETY DISORDER [AMBIGUOUS]|GENERALIZED ANXIETY DISORDER (DISORDER)
C0001818|T048|247830007|SNOMEDCT_US|AGORAPHOBIA|FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|AGORAPHOBIAS|FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|FEAR OF OPEN SPACES|FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|AGORAPHOBIA, UNSPECIFIED|FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|AGORAPHOBIA [DISEASE/FINDING]|FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|AGORAPHOBIA |FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|[X]AGORAPHOBIA|FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|AGORAPHOBIA |FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|FEAR OF OPEN PLACES|FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|PHOBIA OF GOING OUT|FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|FEAR OF OPEN SPACES |FEAR OF OPEN SPACES (FINDING)
C0001818|T048|247830007|SNOMEDCT_US|AGORAPHOBIA, NOS|FEAR OF OPEN SPACES (FINDING)
C0038441|T048||SNOMEDCT_US|TRAUMATIC STRESS DIS
C0038441|T048||SNOMEDCT_US|STRESS DISORDERS
C0038441|T048||SNOMEDCT_US|STRESS DISORDERS, TRAUMATIC [DISEASE/FINDING]
C0038441|T048||SNOMEDCT_US|STRESS DISORDERS, TRAUMATIC
C0038441|T048||SNOMEDCT_US|STRESS DISORDER 
C0038441|T048||SNOMEDCT_US|STRESS DISORDER
C0038441|T048||SNOMEDCT_US|STRESS DISORDER, TRAUMATIC
C0038441|T048||SNOMEDCT_US|TRAUMATIC STRESS DISORDER
C0038441|T048||SNOMEDCT_US|TRAUMATIC STRESS DISORDERS
C0038441|T048||SNOMEDCT_US|DISORDER; STRESS
C0038441|T048||SNOMEDCT_US|STRESS; DISORDER
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DISORDER|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DISORDERS|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|DISORDER, ANXIETY|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|DISORDERS, ANXIETY|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DISORDER, UNSPECIFIED|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DIS|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DISORDER |[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY NOS|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DISORDERS [DISEASE/FINDING]|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DISORDER |[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|[X]ANXIETY DISORDER, UNSPECIFIED|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|[X]ANXIETY DISORDER, UNSPECIFIED |[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
# C0003469|T048|192405006|SNOMEDCT_US|ANXIETY|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DISORDER, NOS|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|ANXIETY DISORDER [AMBIGUOUS]|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0003469|T048|192405006|SNOMEDCT_US|DISORDER;ANXIETY|[X]ANXIETY DISORDER, UNSPECIFIED (DISORDER)
C0376280|T048||SNOMEDCT_US|ANXIETY STATE, NEUROTIC
C0376280|T048||SNOMEDCT_US|NEUROTIC ANXIETY STATE
C0376280|T048||SNOMEDCT_US|NEUROTIC ANXIETY STATES
C0376280|T048||SNOMEDCT_US|STATE, NEUROTIC ANXIETY
C0376280|T048||SNOMEDCT_US|STATES, NEUROTIC ANXIETY
C0376280|T048||SNOMEDCT_US|ANXIETY STATES, NEUROTIC
C0086769|T048|225624000|SNOMEDCT_US|ATTACKS, PANIC|PANIC ATTACK (FINDING)
C0086769|T048|225624000|SNOMEDCT_US|PANIC ATTACK|PANIC ATTACK (FINDING)
C0086769|T048|225624000|SNOMEDCT_US|ATTACK, PANIC|PANIC ATTACK (FINDING)
C0086769|T048|225624000|SNOMEDCT_US|PANIC ATTACKS|PANIC ATTACK (FINDING)
C0086769|T048|225624000|SNOMEDCT_US|ATTACK(S);PANIC|PANIC ATTACK (FINDING)
C0086769|T048|225624000|SNOMEDCT_US|PANIC ATTACK |PANIC ATTACK (FINDING)
C0086769|T048|225624000|SNOMEDCT_US|ATTACK; PANIC|PANIC ATTACK (FINDING)
C0086769|T048|225624000|SNOMEDCT_US|PANIC; ATTACK|PANIC ATTACK (FINDING)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE STRESS DISORDER|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE STRESS REACTION|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|STRESS DIS ACUTE|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|STRESS DIS TRAUMATIC ACUTE|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE STRESS DIS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE STRESS DISORDER |PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE REACTION TO STRESS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE REACTION TO STRESS |PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|GROSS STRESS REACTION, NOS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE STRESS REACT NOS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE CRISIS REACTION|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|PSYCHIC SHOCK|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|STRESS DISORDERS, ACUTE|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|STRESS DISORDERS, TRAUMATIC, ACUTE|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE STRESS DISORDERS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|STRESS DISORDERS, TRAUMATIC, ACUTE [DISEASE/FINDING]|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|REACTION AFTER;ACUTE STRESS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE STRESS REACTION NOS |PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|POST-TRAUMATIC STRESS - ACUTE|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|[X]ACUTE REACTION TO STRESS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE STRESS REACTION NOS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|GROSS STRESS REACTION |PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|GROSS STRESS REACTION|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|[X]PSYCHIC SHOCK|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|PSYCHIC SHOCK |PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|[X]ACUTE CRISIS REACTION|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|(EXAMINATION FEAR) OR (FLYING PHOBIA) OR (STAGE FRIGHT) OR (ACUTE STRESS REACTION NOS) |PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|(EXAMINATION FEAR) OR (FLYING PHOBIA) OR (STAGE FRIGHT) OR (ACUTE STRESS REACTION NOS)|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|[X]ACUTE STRESS REACTION|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|STRESS DISORDER, ACUTE|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE REACTION TO STRESS, UNSPECIFIED|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|UNSPECIFIED ACUTE REACTION TO STRESS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE STRESS DISORDER |PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|CRISIS; ACUTE REACTION|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|DISORDER; ACUTE STRESS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE REACTION; CRISIS|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE; STRESS DISORDER|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|ACUTE; STRESS REACTION|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|PSYCHIC; SHOCK|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|SHOCK; PSYCHIC|PSYCHIC SHOCK (DISORDER)
C0236816|T048|41897001|SNOMEDCT_US|STRESS REACTION; ACUTE|PSYCHIC SHOCK (DISORDER)
C2985218|T048||SNOMEDCT_US|SUBSTANCE-INDUCED ANXIETY DISORDER
C1279420|T048|207363009|SNOMEDCT_US|ANXIETY NEUROSIS|ANXIETY NEUROSIS (FINDING)
C1279420|T048|207363009|SNOMEDCT_US|ANXIETY NEUROSES|ANXIETY NEUROSIS (FINDING)
C1279420|T048|207363009|SNOMEDCT_US|ANXIETY NEUROSIS |ANXIETY NEUROSIS (FINDING)
C1279420|T048|207363009|SNOMEDCT_US|NEUROSIS; ANXIETY|ANXIETY NEUROSIS (FINDING)
C1279420|T048|207363009|SNOMEDCT_US|ANXIETY; NEUROSIS|ANXIETY NEUROSIS (FINDING)
C1279420|T048|207363009|SNOMEDCT_US|NEUROSES, ANXIETY|ANXIETY NEUROSIS (FINDING)
C0236794|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITHOUT AGORAPHOBIA |[X]AGORAPHOBIA WITHOUT HISTORY OF PANIC DISORDER
C0236794|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITHOUT AGORAPHOBIA|[X]AGORAPHOBIA WITHOUT HISTORY OF PANIC DISORDER
C0236794|T048|192394003|SNOMEDCT_US|PANIC DIS W/O AGORPHOBIA|[X]AGORAPHOBIA WITHOUT HISTORY OF PANIC DISORDER
C0236794|T048|192394003|SNOMEDCT_US|PANIC DISORDER [EPISODIC PAROXYSMAL ANXIETY] WITHOUT AGORAPHOBIA|[X]AGORAPHOBIA WITHOUT HISTORY OF PANIC DISORDER
C0236794|T048|192394003|SNOMEDCT_US|[X]AGORAPHOBIA WITHOUT HISTORY OF PANIC DISORDER|[X]AGORAPHOBIA WITHOUT HISTORY OF PANIC DISORDER
C0236794|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITHOUT AGORAPHOBIA |[X]AGORAPHOBIA WITHOUT HISTORY OF PANIC DISORDER
C0236794|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITHOUT AGORAPHOBIA, NOS|[X]AGORAPHOBIA WITHOUT HISTORY OF PANIC DISORDER
C0236800|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITH AGORAPHOBIA|[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITH AGORAPHOBIA |[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|AGORAPHOBIA W PANIC DIS|[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|AGORAPHOBIA WITH PANIC DISORDER|[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|[X]PANIC DISORDER WITH AGORAPHOBIA|[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITH AGORAPHOBIA AND PANIC ATTACKS|[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITH AGORAPHOBIA AND PANIC ATTACKS |[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITH AGORAPHOBIA |[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|DISORDER; PANIC, WITH AGORAPHOBIA|[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|PANIC; DISORDER, WITH AGORAPHOBIA|[X]PANIC DISORDER WITH AGORAPHOBIA
C0236800|T048|192394003|SNOMEDCT_US|PANIC DISORDER WITH AGORAPHOBIA, NOS|[X]PANIC DISORDER WITH AGORAPHOBIA
C1387823|T048||SNOMEDCT_US|MIXED ANXIETY DISORDER
C1387823|T048||SNOMEDCT_US|ANXIETY DISORDER MIXED
C1387823|T048||SNOMEDCT_US|MIXED ANXIETY DISORDER 
C1387823|T048||SNOMEDCT_US|MIXED; ANXIETY DISORDER
C1387823|T048||SNOMEDCT_US|ANXIETY DISORDER; MIXED
C0236730|T048|1686006|SNOMEDCT_US|SEDATIVE, HYPNOTIC AND/OR ANXIOLYTIC-INDUCED ANXIETY DISORDER |SEDATIVE, HYPNOTIC AND/OR ANXIOLYTIC-INDUCED ANXIETY DISORDER (DISORDER)
C0236730|T048|1686006|SNOMEDCT_US|SEDATIVE, HYPNOTIC AND/OR ANXIOLYTIC-INDUCED ANXIETY DISORDER|SEDATIVE, HYPNOTIC AND/OR ANXIOLYTIC-INDUCED ANXIETY DISORDER (DISORDER)
C0236730|T048|1686006|SNOMEDCT_US|SEDATIVE, HYPNOTIC OR ANXIOLYTIC-INDUCED ANXIETY DISORDER|SEDATIVE, HYPNOTIC AND/OR ANXIOLYTIC-INDUCED ANXIETY DISORDER (DISORDER)
C0236715|T048|51493001|SNOMEDCT_US|COCAINE INDUCED ANXIETY DISORDER |COCAINE-INDUCED ANXIETY DISORDER (DISORDER)
C0236715|T048|51493001|SNOMEDCT_US|COCAINE INDUCED ANXIETY DISORDER|COCAINE-INDUCED ANXIETY DISORDER (DISORDER)
C0236715|T048|51493001|SNOMEDCT_US|COCAINE-INDUCED ANXIETY DISORDER|COCAINE-INDUCED ANXIETY DISORDER (DISORDER)
C0236715|T048|51493001|SNOMEDCT_US|COCAINE-INDUCED ANXIETY DISORDER |COCAINE-INDUCED ANXIETY DISORDER (DISORDER)
C0236715|T048|51493001|SNOMEDCT_US|COCAINE; ANXIETY DISORDER|COCAINE-INDUCED ANXIETY DISORDER (DISORDER)
C0236715|T048|51493001|SNOMEDCT_US|ANXIETY DISORDER; DUE TO COCAINE|COCAINE-INDUCED ANXIETY DISORDER (DISORDER)
C0236801|T048|192396001|SNOMEDCT_US|SPECIFIC (ISOLATED) PHOBIAS|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|PHOBIA, SPECIFIC|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|SPECIFIC PHOBIAS|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|PHOBIA, SIMPLE|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|[X]SPECIFIC (ISOLATED) PHOBIAS|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|[X]SIMPLE PHOBIA|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|SPECIFIC PHOBIA|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|SIMPLE PHOBIA|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|SPECIFIC PHOBIA |[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|SIMPLE (SPECIFIC) PHOBIA|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|ISOLATED PHOBIA|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|SIMPLE PHOBIA |[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|PHOBIA; SIMPLE|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|PHOBIA; SPECIFIC|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|SIMPLE; PHOBIA|[X]SIMPLE PHOBIA
C0236801|T048|192396001|SNOMEDCT_US|SPECIFIC; PHOBIA|[X]SIMPLE PHOBIA
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL PHOBIA|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|PHOBIAS, SOCIAL|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL PHOBIAS|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL PHOBIA |SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL PHOBIA, UNSPECIFIED|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL NEUROSIS|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL PHOBIA |SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL PHOBIC DISORDERS|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL ANXIETY DISORDER|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|-- SOCIAL PHOBIA|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|NEUROSIS; SOCIAL|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|PHOBIA; SOCIAL|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL; NEUROSIS|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL; PHOBIA|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|ANXIETY DISORDER; SOCIAL|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|SOCIAL PHOBIA, NOS|SOCIAL PHOBIC DISORDERS
C0031572|T048|191720001|SNOMEDCT_US|PHOBIA, SOCIAL|SOCIAL PHOBIC DISORDERS
C0003477|T048||SNOMEDCT_US|SEPARATION ANXIETY DISORDER
C0003477|T048||SNOMEDCT_US|SEPARATION ANXIETY
C0003477|T048||SNOMEDCT_US|ANXIETY SEPARATION
C0003477|T048||SNOMEDCT_US|SEPARATION ANXIETY 
C0003477|T048||SNOMEDCT_US|SEPARATION ANXIETY 
C0003477|T048||SNOMEDCT_US|DISORDER; SEPARATION ANXIETY
C0003477|T048||SNOMEDCT_US|SEPARATION ANXIETY; DISORDER
C0003471|T048|109006|SNOMEDCT_US|ANXIETY DISORDER OF CHILDHOOD OR ADOLESCENCE|ANXIETY DISORDER OF CHILDHOOD OR ADOLESCENCE (DISORDER)
C0003471|T048|109006|SNOMEDCT_US|ANXIETY DISORDER OF CHILDHOOD OR ADOLESCENCE |ANXIETY DISORDER OF CHILDHOOD OR ADOLESCENCE (DISORDER)
C0003471|T048|109006|SNOMEDCT_US|ANXIETY DISORDER OF CHILDHOOD OR ADOLESCENCE |ANXIETY DISORDER OF CHILDHOOD OR ADOLESCENCE (DISORDER)
C0003471|T048|109006|SNOMEDCT_US|ANXIETY DISORDER OF CHILDHOOD OR ADOLESCENCE, NOS|ANXIETY DISORDER OF CHILDHOOD OR ADOLESCENCE (DISORDER)
C0270590|T048|69479009|SNOMEDCT_US|ANXIETY HYPERVENTILATION |ANXIETY HYPERVENTILATION (DISORDER)
C0270590|T048|69479009|SNOMEDCT_US|ANXIETY HYPERVENTILATION|ANXIETY HYPERVENTILATION (DISORDER)
C0270590|T048|69479009|SNOMEDCT_US|ANXIETY HYPERVENTILATION |ANXIETY HYPERVENTILATION (DISORDER)
C0236748|T048|52910006|SNOMEDCT_US|ORGANIC ANXIETY DISORDER|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ANXIETY DISORDER DUE TO SPECIFIED MEDICAL CONDITION|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ANXIETY DISORDER DUE TO A GENERAL MEDICAL CONDITION|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION |ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ANXIETY DISORDER DUE TO MEDICAL DISORDER|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ORGANIC ANXIETY DISORDER |ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ANXIETY DISORDER ORGANIC|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ORGANIC ANXIETY DISORDER |ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ORGANIC ANXIETY SYNDROME|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ANXIETY DISORDER DUE TO A GENERAL MEDICAL CONDITION |ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|DISORDER; ANXIETY, ORGANIC|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|DISORDER; ORGANIC, ANXIETY|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|MEDICAL CONDITION; CAUSING ANXIETY DISORDER|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ORGANIC; ANXIETY DISORDER|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ORGANIC; DISORDER, ANXIETY|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ANXIETY DISORDER; DUE TO GENERAL MEDICAL CONDITION|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C0236748|T048|52910006|SNOMEDCT_US|ANXIETY DISORDER; ORGANIC|ANXIETY DISORDER DUE TO GENERAL MEDICAL CONDITION
C1842981|T048||SNOMEDCT_US|NEUROTICISM
C3840205|T048|10743001000119103|SNOMEDCT_US|ANXIETY IN CHILDBIRTH|ANXIETY DISORDER IN MOTHER COMPLICATING CHILDBIRTH (DISORDER)
C3840205|T048|10743001000119103|SNOMEDCT_US|ANXIETY DISORDER IN MOTHER COMPLICATING CHILDBIRTH |ANXIETY DISORDER IN MOTHER COMPLICATING CHILDBIRTH (DISORDER)
C3840205|T048|10743001000119103|SNOMEDCT_US|ANXIETY DISORDER IN MOTHER COMPLICATING CHILDBIRTH|ANXIETY DISORDER IN MOTHER COMPLICATING CHILDBIRTH (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROSIS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|DISORDERS, NEUROTIC|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC DISORDER|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC DISORDERS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|DISORDER, NEUROTIC|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|PSYCHONEUROSIS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC DISORDER, UNSPECIFIED|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC DIS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROSIS NOS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROSES|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|PSYCHONEUROSES|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC DISORDERS [DISEASE/FINDING]|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|[X]NEUROTIC DISORDER, UNSPECIFIED |NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|[X] NEUROSIS NOS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|[X]NEUROSIS NOS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|[X]NEUROTIC DISORDER, UNSPECIFIED|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC DISORDER NOS |NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC DISORDER NOS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC DISORDER |NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|PSYCHIATRIC DISORDERS NEUROSIS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROSIS |NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|UNSPECIFIED NEUROTIC DISORDER|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROSIS |NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NONPSYCHOTIC MENTAL DISORDER|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|DISEASE (OR DISORDER); NEUROTIC|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|DISORDER; MENTAL, NEUROTIC|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|DISORDER; NEUROTIC|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|MENTAL; DISORDER, NEUROTIC|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROSIS; STATE|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC; DISORDER|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC; STATE|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|STATE; NEUROSIS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|STATE; NEUROTIC|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROSIS, NOS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NONPSYCHOTIC MENTAL DISORDER, NOS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|PSYCHONEUROSIS NOS|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|DISORDER;NEUROTIC|NEUROSIS (DISORDER)
C0027932|T048|111475002|SNOMEDCT_US|NEUROTIC|NEUROSIS (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|ANXIETY, SEPARATION|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|SEPARATION ANXIETY|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|SEPARATION ANXIETY DISORDER OF CHILDHOOD|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|SEPARATION ANXIETY DISORDER OF CHILDHOOD |[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|ANXIETY DISORDER, SEPARATION|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|SEPARATION ANXIETY DIS|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|ANXIETY, SEPARATION [DISEASE/FINDING]|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|SEPARATION ANXIETY DISORDER|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD |[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD|[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C1527281|T048|192610003|SNOMEDCT_US|SEPARATION ANXIETY DISORDER OF CHILDHOOD |[X]SEPARATION ANXIETY DISORDER OF CHILDHOOD (DISORDER)
C4042925|T048||SNOMEDCT_US|TRAUMA AND STRESSOR RELATED DISORDERS
C4042925|T048||SNOMEDCT_US|TRAUMA AND STRESSOR RELATED DISORDERS [DISEASE/FINDING]
C4042925|T048||SNOMEDCT_US|TRAUMA AND STRESSOR-RELATED DISORDER
C4042925|T048||SNOMEDCT_US|OTHER PSYCHIATRIC DISORDERS TRAUMA AND STRESSOR-RELATED
C4042925|T048||SNOMEDCT_US|TRAUMA AND STRESSOR-RELATED DISORDER 
C3887605|T048|192459009|SNOMEDCT_US|NIGHTMARE DISORDER|[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|NIGHTMARE DISORDER |[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|DREAM ANXIETY DISORDER|[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|[X]DREAM ANXIETY DISORDER|[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|[X] NIGHTMARES OR DREAM ANXIETY DISORDER|[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|[X] NIGHTMARES OR DREAM ANXIETY DISORDER |[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|PARONIRIA|[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|NIGHTMARE|[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|DREAM ANXIETY DISORDER |[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|NIGHTMARE, NOS|[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|NIGHTMARES|[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C3887605|T048|192459009|SNOMEDCT_US|NIGHTMARES NOS|[X] NIGHTMARES OR DREAM ANXIETY DISORDER (DISORDER)
C0338908|T048|192402009|SNOMEDCT_US|MIXED ANXIETY AND DEPRESSIVE DISORDER|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|DEPRESSION WITH ANXIETY|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|DEPRESSION WITH ANXIETY |[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIETY/DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIETY WITH DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|MIXED ANXIETY AND DEPRESSIVE DISORDER |[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIETY DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIOUS DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|MIXED ANXIETY & DEPRESSIVE|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|DEPRESSION; ANXIETY|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|DISORDER; MIXED, ANXIETY AND DEPRESSIVE|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|MIXED; DISORDER, ANXIETY AND DEPRESSIVE|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0338908|T048|192402009|SNOMEDCT_US|ANXIETY; DEPRESSION|[X]MIXED ANXIETY AND DEPRESSIVE DISORDER
C0236708|T048|82339009|SNOMEDCT_US|AMPHETAMINE-INDUCED ANXIETY DISORDER |AMPHETAMINE-INDUCED ANXIETY DISORDER (DISORDER)
C0236708|T048|82339009|SNOMEDCT_US|AMPHETAMINE-INDUCED ANXIETY DISORDER|AMPHETAMINE-INDUCED ANXIETY DISORDER (DISORDER)
C0236708|T048|82339009|SNOMEDCT_US|AMPHETAMINE INDUCED ANXIETY DISORDER|AMPHETAMINE-INDUCED ANXIETY DISORDER (DISORDER)
C0236708|T048|82339009|SNOMEDCT_US|AMPHETAMINE-INDUCED ANXIETY DISORDER |AMPHETAMINE-INDUCED ANXIETY DISORDER (DISORDER)
C0520683|T048|10586006|SNOMEDCT_US|OCCUPATION-RELATED STRESS DISORDER|OCCUPATION-RELATED STRESS DISORDER (DISORDER)
C0520683|T048|10586006|SNOMEDCT_US|OCCUPATION-RELATED STRESS DISORDER |OCCUPATION-RELATED STRESS DISORDER (DISORDER)
C0520683|T048|10586006|SNOMEDCT_US|OCCUPATION-RELATED STRESS DISORDER |OCCUPATION-RELATED STRESS DISORDER (DISORDER)
C0520683|T048|10586006|SNOMEDCT_US|WORK-RELATED STRESS DISORDER|OCCUPATION-RELATED STRESS DISORDER (DISORDER)
C0520683|T048|10586006|SNOMEDCT_US|OCCUPATION-RELATED STRESS DISORDER, NOS|OCCUPATION-RELATED STRESS DISORDER (DISORDER)
C0520683|T048|10586006|SNOMEDCT_US|WORK-RELATED STRESS DISORDER, NOS|OCCUPATION-RELATED STRESS DISORDER (DISORDER)
C0476644|T048|58535001|SNOMEDCT_US|PHYSICAL AND EMOTIONAL EXHAUSTION STATE|PHYSICAL AND EMOTIONAL EXHAUSTION STATE (DISORDER)
C0476644|T048|58535001|SNOMEDCT_US|BURNOUT|PHYSICAL AND EMOTIONAL EXHAUSTION STATE (DISORDER)
C0476644|T048|58535001|SNOMEDCT_US|BURNT OUT|PHYSICAL AND EMOTIONAL EXHAUSTION STATE (DISORDER)
C0476644|T048|58535001|SNOMEDCT_US|BURNT OUT (QUALIFIER VALUE)|PHYSICAL AND EMOTIONAL EXHAUSTION STATE (DISORDER)
C0476644|T048|58535001|SNOMEDCT_US|PHYSICAL AND EMOTIONAL EXHAUSTION STATE |PHYSICAL AND EMOTIONAL EXHAUSTION STATE (DISORDER)
C0476644|T048|58535001|SNOMEDCT_US|BURN-OUT|PHYSICAL AND EMOTIONAL EXHAUSTION STATE (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|OBSESSIONAL NEUROSIS|OBSESSIONAL NEUROSIS (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|NEUROSIS;OBSESSIVE|OBSESSIONAL NEUROSIS (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|OBSESSIONAL NEUROSIS |OBSESSIONAL NEUROSIS (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|OBSESSIONAL NEUROSIS |OBSESSIONAL NEUROSIS (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|OBSESSIVE REACTION|OBSESSIONAL NEUROSIS (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|NEUROSIS; OBSESSIONAL|OBSESSIONAL NEUROSIS (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|NEUROSIS; OBSESSION|OBSESSIONAL NEUROSIS (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|OBSESSION; NEUROSIS|OBSESSIONAL NEUROSIS (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|OBSESSIONAL; NEUROSIS|OBSESSIONAL NEUROSIS (DISORDER)
C0302832|T048|191738003|SNOMEDCT_US|OBSESSIVE NEUROSIS|OBSESSIONAL NEUROSIS (DISORDER)
C1879354|T048||SNOMEDCT_US|SEPARATION ANXIETY
C1879354|T048||SNOMEDCT_US|SEPARATION ANXIETY 
C1879354|T048||SNOMEDCT_US|SEPARATION; ANXIETY
C1879354|T048||SNOMEDCT_US|ANXIETY; SEPARATION
C1879354|T048||SNOMEDCT_US|ANXIETY;SEPARATION
C1408583|T048||SNOMEDCT_US|APPREHENSIVENESS; ABNORMAL
C0850602|T048|426174008|SNOMEDCT_US|CHRONIC STRESS DISORDER|CHRONIC STRESS DISORDER (DISORDER)
C0850602|T048|426174008|SNOMEDCT_US|CHRONIC STRESS DISORDER |CHRONIC STRESS DISORDER (DISORDER)
C0850602|T048|426174008|SNOMEDCT_US|CHRONIC STRESS DISORDER |CHRONIC STRESS DISORDER (DISORDER)
C0850602|T048|426174008|SNOMEDCT_US|DISORDER;CHRONIC STRESS|CHRONIC STRESS DISORDER (DISORDER)
C2063171|T048||SNOMEDCT_US|ANXIETY DISORDER OF UNKNOWN (AXIS III) ETIOLOGY 
C2063171|T048||SNOMEDCT_US|ANXIETY DISORDER OF UNKNOWN (AXIS III) ETIOLOGY
C1112506|T048||SNOMEDCT_US|PSEUDOANGINA
C1112506|T048||SNOMEDCT_US|ANGINA PECTORIS FALSA
C1868709|T048||SNOMEDCT_US|ACTIVATION SYNDROME
C2128829|T048||SNOMEDCT_US|ANXIETY RELIEVED BY MEDICATION 
C2128829|T048||SNOMEDCT_US|ANXIETY RELIEVED BY MEDICATION
C2128830|T048||SNOMEDCT_US|ANXIETY WITH FEAR OF GOING CRAZY 
C2128830|T048||SNOMEDCT_US|ANXIETY WITH FEAR OF GOING CRAZY
C2128830|T048||SNOMEDCT_US|ANXIETY WITH A FEAR OF GOING CRAZY
C2128831|T048||SNOMEDCT_US|ANXIETY WITH FEAR OF LOSING SELF-CONTROL 
C2128831|T048||SNOMEDCT_US|ANXIETY WITH FEAR OF LOSING SELF-CONTROL
C2128831|T048||SNOMEDCT_US|ANXIETY WITH A FEAR OF LOSING SELF-CONTROL
C2219852|T048||SNOMEDCT_US|ANXIETY WITH PERSISTENT WORRY 
C2219852|T048||SNOMEDCT_US|ANXIETY WITH A PERSISTENT WORRY
C2219852|T048||SNOMEDCT_US|ANXIETY WITH PERSISTENT WORRY
C2219854|T048||SNOMEDCT_US|ANXIETY WITH ANTICIPATION OF MISFORTUNE
C2219854|T048||SNOMEDCT_US|ANXIETY WITH ANTICIPATION OF MISFORTUNE 
C2219854|T048||SNOMEDCT_US|ANXIETY WITH AN ANTICIPATION OF MISFORTUNE TO SELF OR OTHERS
C2219856|T048||SNOMEDCT_US|ANXIETY WITH DIFFICULTY BREATHING 
C2219856|T048||SNOMEDCT_US|ANXIETY WITH DIFFICULTY BREATHING
C2219857|T048||SNOMEDCT_US|ANXIETY WITH CHEST PAIN OR DISCOMFORT 
C2219857|T048||SNOMEDCT_US|ANXIETY WITH CHEST PAIN OR DISCOMFORT
C2219858|T048||SNOMEDCT_US|ANXIETY WITH RAPID HEARTBEAT 
C2219858|T048||SNOMEDCT_US|ANXIETY WITH RAPID HEARTBEAT
C2219859|T048||SNOMEDCT_US|ANXIETY WITH CHOKING OR SMOTHERING SENSATIONS
C2219859|T048||SNOMEDCT_US|ANXIETY WITH CHOKING OR SMOTHERING SENSATIONS 
C2219862|T048||SNOMEDCT_US|ANXIETY WITH TINGLING IN HANDS AND FEET 
C2219862|T048||SNOMEDCT_US|ANXIETY WITH TINGLING IN HANDS AND FEET
C2219863|T048||SNOMEDCT_US|ANXIETY WITH MUSCLE TENSION, JITTERS 
C2219863|T048||SNOMEDCT_US|ANXIETY WITH MUSCLE TENSION, JITTERS
C2219864|T048||SNOMEDCT_US|ANXIETY WITH STOMACH DISCOMFORT
C2219864|T048||SNOMEDCT_US|ANXIETY WITH STOMACH DISCOMFORT 
C2219865|T048||SNOMEDCT_US|ANXIETY WITH FREQUENT URINATION OR DIARRHEA
C2219865|T048||SNOMEDCT_US|ANXIETY WITH FREQUENT URINATION OR DIARRHEA 
C2219866|T048||SNOMEDCT_US|ANXIETY WITH HOT AND COLD FLASHES
C2219866|T048||SNOMEDCT_US|ANXIETY WITH HOT AND COLD FLASHES 
C2219867|T048||SNOMEDCT_US|ANXIETY WITH EXCESSIVE SWEATING
C2219867|T048||SNOMEDCT_US|ANXIETY WITH EXCESSIVE SWEATING 
C2219869|T048||SNOMEDCT_US|ANXIETY UNRELATED TO EXERTION OR DANGEROUS SITUATION
C2219869|T048||SNOMEDCT_US|ANXIETY UNRELATED TO EXERTION OR DANGEROUS SITUATION 
C2219869|T048||SNOMEDCT_US|ANXIETY UNRELATED TO EXERTION OR DANGER SITUATION
C2219871|T048||SNOMEDCT_US|CONTINUOUS ANXIETY FOR A MONTH OR MORE
C2219871|T048||SNOMEDCT_US|ANXIETY CONTINUOUSLY FOR A MONTH OR MORE
C2219871|T048||SNOMEDCT_US|ANXIETY CONTINUOUSLY FOR A MONTH OR MORE 
C2219905|T048||SNOMEDCT_US|ANXIETY WITH UNREALISTIC FEAR OF DISEASE 
C2219905|T048||SNOMEDCT_US|ANXIETY WITH UNREALISTIC FEAR OF DISEASE
C2219939|T048||SNOMEDCT_US|ANXIETY FROM ANTICIPATION OF SEPARATION 
C2219939|T048||SNOMEDCT_US|ANXIETY FROM ANTICIPATION OF SEPARATION
C2219951|T048||SNOMEDCT_US|ANXIETY WHICH INTERFERES WITH SOCIAL ACTIVITIES 
C2219951|T048||SNOMEDCT_US|ANXIETY WHICH INTERFERES WITH SOCIAL ACTIVITIES
C2219951|T048||SNOMEDCT_US|ANXIETY INTERFERES WITH SOCIAL ACTIVITIES
C2219952|T048||SNOMEDCT_US|ANXIETY WHICH INTERFERES WITH WORK 
C2219952|T048||SNOMEDCT_US|ANXIETY WHICH INTERFERES WITH WORK
C2219952|T048||SNOMEDCT_US|ANXIETY INTERFERES WITH WORK
C2219955|T048||SNOMEDCT_US|ANXIETY RELIEVED BY CHECKING 
C2219955|T048||SNOMEDCT_US|ANXIETY RELIEVED BY CHECKING
C2219956|T048||SNOMEDCT_US|ANXIETY RELIEVED BY WASHING
C2219956|T048||SNOMEDCT_US|ANXIETY RELIEVED BY WASHING 
C2219957|T048||SNOMEDCT_US|ANXIETY RELIEVED BY A RITUAL 
C2219957|T048||SNOMEDCT_US|ANXIETY RELIEVED BY A RITUAL
C3162298|T048||SNOMEDCT_US|ANXIETY ABOUT MEDICAL CONDITION 
C3162298|T048||SNOMEDCT_US|ANXIETY ABOUT MEDICAL CONDITION
C3162299|T048||SNOMEDCT_US|ANXIETY ABOUT MEDICAL REGIMEN
C3162299|T048||SNOMEDCT_US|ANXIETY ABOUT MEDICAL REGIMEN 
C3854439|T048||SNOMEDCT_US|PROCEDURAL ANXIETY
C3854440|T048||SNOMEDCT_US|IMMUNISATION ANXIETY RELATED REACTION
C3854440|T048||SNOMEDCT_US|IMMUNIZATION ANXIETY RELATED REACTION
C3864091|T048||SNOMEDCT_US|ANXIETY ABOUT PLANNED SURGERY
C3864091|T048||SNOMEDCT_US|ANXIETY ABOUT PLANNED SURGERY 
C1561362|T048||SNOMEDCT_US|CTCAE GRADE 2 ANXIETY
C1561362|T048||SNOMEDCT_US|GRADE 2 ANXIETY
C1561364|T048||SNOMEDCT_US|CTCAE GRADE 4 ANXIETY
C1561364|T048||SNOMEDCT_US|GRADE 4 ANXIETY
C1561361|T048||SNOMEDCT_US|CTCAE GRADE 1 ANXIETY
C1561361|T048||SNOMEDCT_US|GRADE 1 ANXIETY
C1561365|T048||SNOMEDCT_US|CTCAE GRADE 5 ANXIETY
C1561365|T048||SNOMEDCT_US|GRADE 5 ANXIETY
C1561363|T048||SNOMEDCT_US|CTCAE GRADE 3 ANXIETY
C1561363|T048||SNOMEDCT_US|GRADE 3 ANXIETY
